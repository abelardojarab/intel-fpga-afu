// (C) 2001-2017 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


//
//              ALTERA CORPORATION
//
//
//


`timescale 1 ps/1 ps
// altera message_off 10036


module twentynm_pcs_rev_20nm1
	#(
	//PARAM_LIST_START
		parameter xcvr_native_mode = "mode_duplex",  // mode_duplex, mode_rx_only, mode_tx_only
		
		// parameters for twentynm_hssi_10g_rx_pcs
		parameter hssi_10g_rx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_align_del = "align_del_en", // align_del_dis|align_del_en
		parameter hssi_10g_rx_pcs_ber_bit_err_total_cnt = "bit_err_total_cnt_10g", // bit_err_total_cnt_10g
		parameter hssi_10g_rx_pcs_ber_clken = "ber_clk_dis", // ber_clk_dis|ber_clk_en
		parameter hssi_10g_rx_pcs_ber_xus_timer_window = 21'b100110001001010,
		parameter hssi_10g_rx_pcs_bitslip_mode = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_rx_pcs_blksync_bitslip_type = "bitslip_comb", // bitslip_comb|bitslip_reg
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_cnt = 3'b1,
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_type = "bitslip_match", // bitslip_match|bitslip_cnt
		parameter hssi_10g_rx_pcs_blksync_bypass = "blksync_bypass_dis", // blksync_bypass_dis|blksync_bypass_en
		parameter hssi_10g_rx_pcs_blksync_clken = "blksync_clk_dis", // blksync_clk_dis|blksync_clk_en
		parameter hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt = "enum_invalid_sh_cnt_10g", // enum_invalid_sh_cnt_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock = "knum_sh_cnt_postlock_10g", // knum_sh_cnt_postlock_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock = "knum_sh_cnt_prelock_10g", // knum_sh_cnt_prelock_10g
		parameter hssi_10g_rx_pcs_blksync_pipeln = "blksync_pipeln_dis", // blksync_pipeln_dis|blksync_pipeln_en
		parameter hssi_10g_rx_pcs_clr_errblk_cnt_en = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_control_del = "control_del_all", // control_del_all|control_del_none
		parameter hssi_10g_rx_pcs_crcchk_bypass = "crcchk_bypass_dis", // crcchk_bypass_dis|crcchk_bypass_en
		parameter hssi_10g_rx_pcs_crcchk_clken = "crcchk_clk_dis", // crcchk_clk_dis|crcchk_clk_en
		parameter hssi_10g_rx_pcs_crcchk_inv = "crcchk_inv_dis", // crcchk_inv_dis|crcchk_inv_en
		parameter hssi_10g_rx_pcs_crcchk_pipeln = "crcchk_pipeln_dis", // crcchk_pipeln_dis|crcchk_pipeln_en
		parameter hssi_10g_rx_pcs_crcflag_pipeln = "crcflag_pipeln_dis", // crcflag_pipeln_dis|crcflag_pipeln_en
		parameter hssi_10g_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_rx_pcs_dec64b66b_clken = "dec64b66b_clk_dis", // dec64b66b_clk_dis|dec64b66b_clk_en
		parameter hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass = "dec_64b66b_rxsm_bypass_dis", // dec_64b66b_rxsm_bypass_dis|dec_64b66b_rxsm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_bypass = "descrm_bypass_en", // descrm_bypass_dis|descrm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_clken = "descrm_clk_dis", // descrm_clk_dis|descrm_clk_en
		parameter hssi_10g_rx_pcs_descrm_mode = "async", // async|sync
		parameter hssi_10g_rx_pcs_descrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_dft_clk_out_sel = "rx_master_clk", // rx_master_clk|rx_gbexp_clk|rx_blksync_clk|rx_descrm_clk|rx_frmsync_clk|rx_64b66bdec_clk|rx_ber_clk|rx_rand_clk|rx_crcchk_clk|rx_wrfifo_clk|rx_rdfifo_clk|rx_fec_clk
		parameter hssi_10g_rx_pcs_dis_signal_ok = "dis_signal_ok_dis", // dis_signal_ok_dis|dis_signal_ok_en
		parameter hssi_10g_rx_pcs_dispchk_bypass = "dispchk_bypass_dis", // dispchk_bypass_dis|dispchk_bypass_en
		parameter hssi_10g_rx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_rx_pcs_fast_path = "fast_path_dis", // fast_path_dis|fast_path_en
		parameter hssi_10g_rx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_rx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_rx_pcs_fifo_double_read = "fifo_double_read_dis", // fifo_double_read_dis|fifo_double_read_en
		parameter hssi_10g_rx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_rx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_rx_pcs_force_align = "force_align_dis", // force_align_dis|force_align_en
		parameter hssi_10g_rx_pcs_frmsync_bypass = "frmsync_bypass_dis", // frmsync_bypass_dis|frmsync_bypass_en
		parameter hssi_10g_rx_pcs_frmsync_clken = "frmsync_clk_dis", // frmsync_clk_dis|frmsync_clk_en
		parameter hssi_10g_rx_pcs_frmsync_enum_scrm = "enum_scrm_default", // enum_scrm_default
		parameter hssi_10g_rx_pcs_frmsync_enum_sync = "enum_sync_default", // enum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_flag_type = "all_framing_words", // all_framing_words|location_only
		parameter hssi_10g_rx_pcs_frmsync_knum_sync = "knum_sync_default", // knum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_mfrm_length = 16'b100000000000,
		parameter hssi_10g_rx_pcs_frmsync_pipeln = "frmsync_pipeln_dis", // frmsync_pipeln_dis|frmsync_pipeln_en
		parameter hssi_10g_rx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_rx_pcs_gb_rx_idwidth = "width_32", // width_40|width_32|width_64
		parameter hssi_10g_rx_pcs_gb_rx_odwidth = "width_66", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_rx_pcs_gbexp_clken = "gbexp_clk_dis", // gbexp_clk_dis|gbexp_clk_en
		parameter hssi_10g_rx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_10g_rx_pcs_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_rx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_rx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_rx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_rx_pcs_pld_if_type = "fifo", // fifo|reg
		parameter hssi_10g_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_rx_pcs_rand_clken = "rand_clk_dis", // rand_clk_dis|rand_clk_en
		parameter hssi_10g_rx_pcs_rd_clk_sel = "rd_rx_pma_clk", // rd_rx_pld_clk|rd_rx_pma_clk|rd_refclk_dig
		parameter hssi_10g_rx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_rx_pcs_rx_fifo_write_ctrl = "blklock_stops", // blklock_stops|blklock_ignore
		parameter hssi_10g_rx_pcs_rx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_rx_pcs_rx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_rx_pcs_rx_signal_ok_sel = "synchronized_ver", // synchronized_ver|nonsync_ver
		parameter hssi_10g_rx_pcs_rx_sm_bypass = "rx_sm_bypass_dis", // rx_sm_bypass_dis|rx_sm_bypass_en
		parameter hssi_10g_rx_pcs_rx_sm_hiber = "rx_sm_hiber_en", // rx_sm_hiber_en|rx_sm_hiber_dis
		parameter hssi_10g_rx_pcs_rx_sm_pipeln = "rx_sm_pipeln_dis", // rx_sm_pipeln_dis|rx_sm_pipeln_en
		parameter hssi_10g_rx_pcs_rx_testbus_sel = "crc32_chk_testbus1", // crc32_chk_testbus1|crc32_chk_testbus2|frame_sync_testbus1|frame_sync_testbus2|dec64b66b_testbus|rxsm_testbus|ber_testbus|blksync_testbus1|blksync_testbus2|gearbox_exp_testbus|random_ver_testbus|descramble_testbus|blank_testbus|rx_fifo_testbus1|rx_fifo_testbus2
		parameter hssi_10g_rx_pcs_rx_true_b2b = "b2b", // single|b2b
		parameter hssi_10g_rx_pcs_rxfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_rx_pcs_rxfifo_full = "full_default", // full_default
		parameter hssi_10g_rx_pcs_rxfifo_mode = "phase_comp", // register_mode|clk_comp_10g|generic_interlaken|generic_basic|phase_comp|phase_comp_dv
		parameter hssi_10g_rx_pcs_rxfifo_pempty = 5'b10,
		parameter hssi_10g_rx_pcs_rxfifo_pfull = 5'b10111,
		parameter hssi_10g_rx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_rx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_rx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_10g_tx_pcs
		parameter hssi_10g_tx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_bitslip_en = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_10g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_10g_tx_pcs_comp_cnt = 8'b0,
		parameter hssi_10g_tx_pcs_compin_sel = "compin_master", // compin_master|compin_slave_top|compin_slave_bot|compin_default
		parameter hssi_10g_tx_pcs_crcgen_bypass = "crcgen_bypass_dis", // crcgen_bypass_dis|crcgen_bypass_en
		parameter hssi_10g_tx_pcs_crcgen_clken = "crcgen_clk_dis", // crcgen_clk_dis|crcgen_clk_en
		parameter hssi_10g_tx_pcs_crcgen_err = "crcgen_err_dis", // crcgen_err_dis|crcgen_err_en
		parameter hssi_10g_tx_pcs_crcgen_inv = "crcgen_inv_dis", // crcgen_inv_dis|crcgen_inv_en
		parameter hssi_10g_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_tx_pcs_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_10g_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_tx_pcs_dft_clk_out_sel = "tx_master_clk", // tx_master_clk|tx_rdfifo_clk|tx_frmgen_clk|tx_crcgen_clk|tx_64b66benc_txsm_clk|tx_scrm_clk|tx_dispgen_clk|tx_gbred_clk|tx_wrfifo_clk|tx_fec_clk
		parameter hssi_10g_tx_pcs_dispgen_bypass = "dispgen_bypass_dis", // dispgen_bypass_dis|dispgen_bypass_en
		parameter hssi_10g_tx_pcs_dispgen_clken = "dispgen_clk_dis", // dispgen_clk_dis|dispgen_clk_en
		parameter hssi_10g_tx_pcs_dispgen_err = "dispgen_err_dis", // dispgen_err_dis|dispgen_err_en
		parameter hssi_10g_tx_pcs_dispgen_pipeln = "dispgen_pipeln_dis", // dispgen_pipeln_dis|dispgen_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_bypass_pipeln = "distdwn_bypass_pipeln_dis", // distdwn_bypass_pipeln_dis|distdwn_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_master = "distdwn_master_en", // distdwn_master_en|distdwn_master_dis
		parameter hssi_10g_tx_pcs_distup_bypass_pipeln = "distup_bypass_pipeln_dis", // distup_bypass_pipeln_dis|distup_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distup_master = "distup_master_en", // distup_master_en|distup_master_dis
		parameter hssi_10g_tx_pcs_dv_bond = "dv_bond_dis", // dv_bond_en|dv_bond_dis
		parameter hssi_10g_tx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_tx_pcs_enc64b66b_txsm_clken = "enc64b66b_txsm_clk_dis", // enc64b66b_txsm_clk_dis|enc64b66b_txsm_clk_en
		parameter hssi_10g_tx_pcs_enc_64b66b_txsm_bypass = "enc_64b66b_txsm_bypass_dis", // enc_64b66b_txsm_bypass_dis|enc_64b66b_txsm_bypass_en
		parameter hssi_10g_tx_pcs_fastpath = "fastpath_dis", // fastpath_dis|fastpath_en
		parameter hssi_10g_tx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_tx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_tx_pcs_fifo_double_write = "fifo_double_write_dis", // fifo_double_write_dis|fifo_double_write_en
		parameter hssi_10g_tx_pcs_fifo_reg_fast = "fifo_reg_fast_dis", // fifo_reg_fast_dis|fifo_reg_fast_en
		parameter hssi_10g_tx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_tx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_tx_pcs_frmgen_burst = "frmgen_burst_dis", // frmgen_burst_dis|frmgen_burst_en
		parameter hssi_10g_tx_pcs_frmgen_bypass = "frmgen_bypass_dis", // frmgen_bypass_dis|frmgen_bypass_en
		parameter hssi_10g_tx_pcs_frmgen_clken = "frmgen_clk_dis", // frmgen_clk_dis|frmgen_clk_en
		parameter hssi_10g_tx_pcs_frmgen_mfrm_length = 16'b100000000000,
		parameter hssi_10g_tx_pcs_frmgen_pipeln = "frmgen_pipeln_dis", // frmgen_pipeln_dis|frmgen_pipeln_en
		parameter hssi_10g_tx_pcs_frmgen_pyld_ins = "frmgen_pyld_ins_dis", // frmgen_pyld_ins_dis|frmgen_pyld_ins_en
		parameter hssi_10g_tx_pcs_frmgen_wordslip = "frmgen_wordslip_dis", // frmgen_wordslip_dis|frmgen_wordslip_en
		parameter hssi_10g_tx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_tx_pcs_gb_pipeln_bypass = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_gb_tx_idwidth = "width_50", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_tx_pcs_gb_tx_odwidth = "width_32", // width_32|width_40|width_64
		parameter hssi_10g_tx_pcs_gbred_clken = "gbred_clk_dis", // gbred_clk_dis|gbred_clk_en
		parameter hssi_10g_tx_pcs_indv = "indv_en", // indv_en|indv_dis
		parameter hssi_10g_tx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_tx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_tx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_tx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del6|phcomp_rd_del5|phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_tx_pcs_pld_if_type = "fifo", // fifo|reg|fastreg
		parameter hssi_10g_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_tx_pcs_pseudo_random = "all_0", // two_lf|all_0
		parameter hssi_10g_tx_pcs_pseudo_seed_a = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_pseudo_seed_b = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_random_disp = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_tx_pcs_scrm_bypass = "scrm_bypass_dis", // scrm_bypass_dis|scrm_bypass_en
		parameter hssi_10g_tx_pcs_scrm_clken = "scrm_clk_dis", // scrm_clk_dis|scrm_clk_en
		parameter hssi_10g_tx_pcs_scrm_mode = "async", // async|sync
		parameter hssi_10g_tx_pcs_scrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_sh_err = "sh_err_dis", // sh_err_dis|sh_err_en
		parameter hssi_10g_tx_pcs_sop_mark = "sop_mark_dis", // sop_mark_en|sop_mark_dis
		parameter hssi_10g_tx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_tx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_tx_pcs_tx_scrm_err = "scrm_err_dis", // scrm_err_dis|scrm_err_en
		parameter hssi_10g_tx_pcs_tx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_tx_pcs_tx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_tx_pcs_tx_sm_bypass = "tx_sm_bypass_dis", // tx_sm_bypass_dis|tx_sm_bypass_en
		parameter hssi_10g_tx_pcs_tx_sm_pipeln = "tx_sm_pipeln_dis", // tx_sm_pipeln_dis|tx_sm_pipeln_en
		parameter hssi_10g_tx_pcs_tx_testbus_sel = "crc32_gen_testbus1", // crc32_gen_testbus1|crc32_gen_testbus2|disp_gen_testbus1|disp_gen_testbus2|frame_gen_testbus1|frame_gen_testbus2|enc64b66b_testbus|txsm_testbus|tx_cp_bond_testbus|gearbox_red_testbus|scramble_testbus|blank_testbus|tx_fifo_testbus1|tx_fifo_testbus2
		parameter hssi_10g_tx_pcs_txfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_tx_pcs_txfifo_full = "full_default", // full_default
		parameter hssi_10g_tx_pcs_txfifo_mode = "phase_comp", // register_mode|interlaken_generic|basic_generic|phase_comp
		parameter hssi_10g_tx_pcs_txfifo_pempty = 4'b10,
		parameter hssi_10g_tx_pcs_txfifo_pfull = 4'b1011,
		parameter hssi_10g_tx_pcs_wr_clk_sel = "wr_tx_pma_clk", // wr_tx_pld_clk|wr_tx_pma_clk|wr_refclk_dig
		parameter hssi_10g_tx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_8g_rx_pcs
		parameter hssi_8g_rx_pcs_auto_error_replacement = "dis_err_replace", // dis_err_replace|en_err_replace
		parameter hssi_8g_rx_pcs_auto_speed_nego = "dis_asn", // dis_asn|en_asn_g2_freq_scal
		parameter hssi_8g_rx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_rx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_rx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_rx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_rx_pcs_byte_deserializer = "dis_bds", // dis_bds|en_bds_by_2|en_bds_by_4|en_bds_by_2_det
		parameter hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask = "dis_rxvalid_mask", // dis_rxvalid_mask|en_rxvalid_mask
		parameter hssi_8g_rx_pcs_clkcmp_pattern_n = 20'b0,
		parameter hssi_8g_rx_pcs_clkcmp_pattern_p = 20'b0,
		parameter hssi_8g_rx_pcs_clock_gate_bds_dec_asn = "dis_bds_dec_asn_clk_gating", // dis_bds_dec_asn_clk_gating|en_bds_dec_asn_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_cdr_eidle = "dis_cdr_eidle_clk_gating", // dis_cdr_eidle_clk_gating|en_cdr_eidle_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk = "dis_dw_pc_wrclk_gating", // dis_dw_pc_wrclk_gating|en_dw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_rd = "dis_dw_rm_rdclk_gating", // dis_dw_rm_rdclk_gating|en_dw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_wr = "dis_dw_rm_wrclk_gating", // dis_dw_rm_wrclk_gating|en_dw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_wa = "dis_dw_wa_clk_gating", // dis_dw_wa_clk_gating|en_dw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_pc_rdclk = "dis_pc_rdclk_gating", // dis_pc_rdclk_gating|en_pc_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk = "dis_sw_pc_wrclk_gating", // dis_sw_pc_wrclk_gating|en_sw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_rd = "dis_sw_rm_rdclk_gating", // dis_sw_rm_rdclk_gating|en_sw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_wr = "dis_sw_rm_wrclk_gating", // dis_sw_rm_wrclk_gating|en_sw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_wa = "dis_sw_wa_clk_gating", // dis_sw_wa_clk_gating|en_sw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_observation_in_pld_core = "internal_sw_wa_clk", // internal_sw_wa_clk|internal_dw_wa_clk|internal_cdr_eidle_clk|internal_sm_rm_wr_clk|internal_dw_rm_wr_clk|internal_clk_2_b|internal_sw_rm_rd_clk|internal_dw_rm_rd_clk|internal_sw_rx_wr_clk|internal_dw_rx_wr_clk|internal_rx_rd_clk|internal_rx_pma_clk_gen3|internal_rx_rcvd_clk_gen3
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_rx_pcs_eidle_entry_eios = "dis_eidle_eios", // dis_eidle_eios|en_eidle_eios
		parameter hssi_8g_rx_pcs_eidle_entry_iei = "dis_eidle_iei", // dis_eidle_iei|en_eidle_iei
		parameter hssi_8g_rx_pcs_eidle_entry_sd = "dis_eidle_sd", // dis_eidle_sd|en_eidle_sd
		parameter hssi_8g_rx_pcs_eightb_tenb_decoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_rx_pcs_err_flags_sel = "err_flags_wa", // err_flags_wa|err_flags_8b10b
		parameter hssi_8g_rx_pcs_fixed_pat_det = "dis_fixed_patdet", // dis_fixed_patdet|en_fixed_patdet
		parameter hssi_8g_rx_pcs_fixed_pat_num = 4'b1111,
		parameter hssi_8g_rx_pcs_force_signal_detect = "en_force_signal_detect", // en_force_signal_detect|dis_force_signal_detect
		parameter hssi_8g_rx_pcs_gen3_clk_en = "disable_clk", // disable_clk|enable_clk
		parameter hssi_8g_rx_pcs_gen3_rx_clk_sel = "rcvd_clk", // en_dig_clk1_8g|rcvd_clk
		parameter hssi_8g_rx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // en_dig_clk2_8g|tx_pma_clk
		parameter hssi_8g_rx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_rx_pcs_ibm_invalid_code = "dis_ibm_invalid_code", // dis_ibm_invalid_code|en_ibm_invalid_code
		parameter hssi_8g_rx_pcs_invalid_code_flag_only = "dis_invalid_code_only", // dis_invalid_code_only|en_invalid_code_only
		parameter hssi_8g_rx_pcs_pad_or_edb_error_replace = "replace_edb", // replace_edb|replace_edb_dynamic|replace_pad
		parameter hssi_8g_rx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_rx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_rx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_rx_pcs_pipe_if_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_8g_rx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_rx_pcs_polinv_8b10b_dec = "dis_polinv_8b10b_dec", // dis_polinv_8b10b_dec|en_polinv_8b10b_dec
		parameter hssi_8g_rx_pcs_prot_mode = "gige", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic_rm_enable|basic_rm_disable|disabled_prot_mode
		parameter hssi_8g_rx_pcs_rate_match = "dis_rm", // dis_rm|gige_rm|pipe_rm|pipe_rm_0ppm|sw_basic_rm|dw_basic_rm
		parameter hssi_8g_rx_pcs_rate_match_del_thres = "dis_rm_del_thres", // dis_rm_del_thres|gige_rm_del_thres|pipe_rm_del_thres|pipe_rm_0ppm_del_thres|sw_basic_rm_del_thres|dw_basic_rm_del_thres
		parameter hssi_8g_rx_pcs_rate_match_empty_thres = "dis_rm_empty_thres", // dis_rm_empty_thres|gige_rm_empty_thres|pipe_rm_empty_thres|pipe_rm_0ppm_empty_thres|sw_basic_rm_empty_thres|dw_basic_rm_empty_thres
		parameter hssi_8g_rx_pcs_rate_match_full_thres = "dis_rm_full_thres", // dis_rm_full_thres|gige_rm_full_thres|pipe_rm_full_thres|pipe_rm_0ppm_full_thres|sw_basic_rm_full_thres|dw_basic_rm_full_thres
		parameter hssi_8g_rx_pcs_rate_match_ins_thres = "dis_rm_ins_thres", // dis_rm_ins_thres|gige_rm_ins_thres|pipe_rm_ins_thres|pipe_rm_0ppm_ins_thres|sw_basic_rm_ins_thres|dw_basic_rm_ins_thres
		parameter hssi_8g_rx_pcs_rate_match_start_thres = "dis_rm_start_thres", // dis_rm_start_thres|gige_rm_start_thres|pipe_rm_start_thres|pipe_rm_0ppm_start_thres|sw_basic_rm_start_thres|dw_basic_rm_start_thres
		parameter hssi_8g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_rx_pcs_rx_clk2 = "rcvd_clk_clk2", // rcvd_clk_clk2|tx_pma_clock_clk2|refclk_dig2_clk2
		parameter hssi_8g_rx_pcs_rx_clk_free_running = "en_rx_clk_free_run", // dis_rx_clk_free_run|en_rx_clk_free_run
		parameter hssi_8g_rx_pcs_rx_pcs_urst = "en_rx_pcs_urst", // dis_rx_pcs_urst|en_rx_pcs_urst
		parameter hssi_8g_rx_pcs_rx_rcvd_clk = "rcvd_clk_rcvd_clk", // rcvd_clk_rcvd_clk|tx_pma_clock_rcvd_clk
		parameter hssi_8g_rx_pcs_rx_rd_clk = "pld_rx_clk", // pld_rx_clk|rx_clk
		parameter hssi_8g_rx_pcs_rx_refclk = "dis_refclk_sel", // dis_refclk_sel|en_refclk_sel
		parameter hssi_8g_rx_pcs_rx_wr_clk = "rx_clk2_div_1_2_4", // rx_clk2_div_1_2_4|txfifo_rd_clk
		parameter hssi_8g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_rx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_rx_pcs_sync_sm_idle_eios = "dis_syncsm_idle", // dis_syncsm_idle|en_syncsm_idle
		parameter hssi_8g_rx_pcs_test_bus_sel = "tx_testbus", // tx_testbus|tx_ctrl_plane_testbus|wa_testbus|rm_testbus|rx_ctrl_testbus|pcie_ctrl_testbus|rx_ctrl_plane_testbus
		parameter hssi_8g_rx_pcs_tx_rx_parallel_loopback = "dis_plpbk", // dis_plpbk|en_plpbk
		parameter hssi_8g_rx_pcs_wa_boundary_lock_ctrl = "bit_slip", // bit_slip|sync_sm|deterministic_latency|auto_align_pld_ctrl
		parameter hssi_8g_rx_pcs_wa_clk_slip_spacing = 10'b10000,
		parameter hssi_8g_rx_pcs_wa_det_latency_sync_status_beh = "assert_sync_status_non_imm", // assert_sync_status_imm|assert_sync_status_non_imm|dont_care_assert_sync
		parameter hssi_8g_rx_pcs_wa_disp_err_flag = "dis_disp_err_flag", // dis_disp_err_flag|en_disp_err_flag
		parameter hssi_8g_rx_pcs_wa_kchar = "dis_kchar", // dis_kchar|en_kchar
		parameter hssi_8g_rx_pcs_wa_pd = "wa_pd_10", // wa_pd_7|wa_pd_10|wa_pd_20|wa_pd_40|wa_pd_8_sw|wa_pd_8_dw|wa_pd_16_sw|wa_pd_16_dw|wa_pd_32
		parameter hssi_8g_rx_pcs_wa_pd_data = 40'b0,
		parameter hssi_8g_rx_pcs_wa_pd_polarity = "dis_pd_both_pol", // dis_pd_both_pol|en_pd_both_pol|dont_care_both_pol
		parameter hssi_8g_rx_pcs_wa_pld_controlled = "dis_pld_ctrl", // dis_pld_ctrl|pld_ctrl_sw|rising_edge_sensitive_dw|level_sensitive_dw
		parameter hssi_8g_rx_pcs_wa_renumber_data = 6'b0,
		parameter hssi_8g_rx_pcs_wa_rgnumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rknumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rosnumber_data = 2'b0,
		parameter hssi_8g_rx_pcs_wa_rvnumber_data = 13'b0,
		parameter hssi_8g_rx_pcs_wa_sync_sm_ctrl = "gige_sync_sm", // gige_sync_sm|pipe_sync_sm|sw_basic_sync_sm|dw_basic_sync_sm|fibre_channel_sync_sm
		parameter hssi_8g_rx_pcs_wait_cnt = 12'b0,
		
		// parameters for twentynm_hssi_8g_tx_pcs
		parameter hssi_8g_tx_pcs_auto_speed_nego_gen2 = "dis_asn_g2", // dis_asn_g2|en_asn_g2_freq_scal
		parameter hssi_8g_tx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_tx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_tx_pcs_byte_serializer = "dis_bs", // dis_bs|en_bs_by_2|en_bs_by_4
		parameter hssi_8g_tx_pcs_clock_gate_bs_enc = "dis_bs_enc_clk_gating", // dis_bs_enc_clk_gating|en_bs_enc_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_dw_fifowr = "dis_dw_fifowr_clk_gating", // dis_dw_fifowr_clk_gating|en_dw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_fiford = "dis_fiford_clk_gating", // dis_fiford_clk_gating|en_fiford_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_sw_fifowr = "dis_sw_fifowr_clk_gating", // dis_sw_fifowr_clk_gating|en_sw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_observation_in_pld_core = "internal_refclk_b", // internal_refclk_b|internal_fifo_rd_clk|internal_sw_fifo_wr_clk|internal_dw_fifo_wr_clk|internal_tx_clk_out_gen3|internal_pipe_tx_clk_out_gen3
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_tx_pcs_data_selection_8b10b_encoder_input = "normal_data_path", // normal_data_path|gige_idle_conversion
		parameter hssi_8g_tx_pcs_dynamic_clk_switch = "dis_dyn_clk_switch", // dis_dyn_clk_switch|en_dyn_clk_switch
		parameter hssi_8g_tx_pcs_eightb_tenb_disp_ctrl = "dis_disp_ctrl", // dis_disp_ctrl|en_disp_ctrl|en_ib_disp_ctrl
		parameter hssi_8g_tx_pcs_eightb_tenb_encoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_tx_pcs_force_echar = "dis_force_echar", // dis_force_echar|en_force_echar
		parameter hssi_8g_tx_pcs_force_kchar = "dis_force_kchar", // dis_force_kchar|en_force_kchar
		parameter hssi_8g_tx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // dis_tx_clk|tx_pma_clk
		parameter hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel = "func_clk", // dis_tx_pipe_clk|func_clk
		parameter hssi_8g_tx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_tx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_tx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_tx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_tx_pcs_phfifo_write_clk_sel = "pld_tx_clk", // pld_tx_clk|tx_clk
		parameter hssi_8g_tx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_tx_pcs_prot_mode = "basic", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic|disabled_prot_mode
		parameter hssi_8g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_tx_pcs_refclk_b_clk_sel = "tx_pma_clock", // tx_pma_clock|refclk_dig
		parameter hssi_8g_tx_pcs_revloop_back_rm = "dis_rev_loopback_rx_rm", // dis_rev_loopback_rx_rm|en_rev_loopback_rx_rm
		parameter hssi_8g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_tx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_tx_pcs_tx_bitslip = "dis_tx_bitslip", // dis_tx_bitslip|en_tx_bitslip
		parameter hssi_8g_tx_pcs_tx_compliance_controlled_disparity = "dis_txcompliance", // dis_txcompliance|en_txcompliance_pipe2p0|en_txcompliance_pipe3p0
		parameter hssi_8g_tx_pcs_tx_fast_pld_reg = "dis_tx_fast_pld_reg", // dis_tx_fast_pld_reg|en_tx_fast_pld_reg
		parameter hssi_8g_tx_pcs_txclk_freerun = "dis_freerun_tx", // dis_freerun_tx|en_freerun_tx
		parameter hssi_8g_tx_pcs_txpcs_urst = "en_txpcs_urst", // dis_txpcs_urst|en_txpcs_urst
		
		// parameters for twentynm_hssi_common_pcs_pma_interface
		parameter hssi_common_pcs_pma_interface_asn_clk_enable = "false", // false|true
		parameter hssi_common_pcs_pma_interface_asn_enable = "dis_asn", // dis_asn|en_asn
		parameter hssi_common_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|pcie_gen3
		parameter hssi_common_pcs_pma_interface_bypass_early_eios = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pcie_switch = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_ltr = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_sw_done = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_ppm_lock = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_txdetectrx = "false", // false|true
		parameter hssi_common_pcs_pma_interface_cdr_control = "en_cdr_ctrl", // dis_cdr_ctrl|en_cdr_ctrl
		parameter hssi_common_pcs_pma_interface_cid_enable = "en_cid_mode", // dis_cid_mode|en_cid_mode
		parameter hssi_common_pcs_pma_interface_cp_cons_sel = "cp_cons_default", // cp_cons_master|cp_cons_slave_abv|cp_cons_slave_blw|cp_cons_default
		parameter hssi_common_pcs_pma_interface_cp_dwn_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_cp_up_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_blw|ctrl_slave_abv
		parameter hssi_common_pcs_pma_interface_data_mask_count = 16'b100111000100,
		parameter hssi_common_pcs_pma_interface_data_mask_count_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_dft_observation_clock_selection = "dft_clk_obsrv_tx0", // dft_clk_obsrv_tx0|dft_clk_obsrv_tx1|dft_clk_obsrv_tx2|dft_clk_obsrv_tx3|dft_clk_obsrv_tx4|dft_clk_obsrv_rx|dft_clk_obsrv_hclk|dft_clk_obsrv_fref|dft_clk_obsrv_clklow|dft_clk_obsrv_asn0|dft_clk_obsrv_asn1
		parameter hssi_common_pcs_pma_interface_early_eios_counter = 8'b110010,
		parameter hssi_common_pcs_pma_interface_force_freqdet = "force_freqdet_dis", // force_freqdet_dis|force1_freqdet_en|force0_freqdet_en
		parameter hssi_common_pcs_pma_interface_free_run_clk_enable = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ignore_sigdet_g23 = "false", // false|true
		parameter hssi_common_pcs_pma_interface_pc_en_counter = 7'b110111,
		parameter hssi_common_pcs_pma_interface_pc_rst_counter = 5'b10111,
		parameter hssi_common_pcs_pma_interface_pcie_hip_mode = "hip_disable", // hip_enable|hip_disable
		parameter hssi_common_pcs_pma_interface_ph_fifo_reg_mode = "phfifo_reg_mode_dis", // phfifo_reg_mode_dis|phfifo_reg_mode_en
		parameter hssi_common_pcs_pma_interface_phfifo_flush_wait = 6'b100100,
		parameter hssi_common_pcs_pma_interface_pipe_if_g3pcs = "pipe_if_8gpcs", // pipe_if_g3pcs|pipe_if_8gpcs
		parameter hssi_common_pcs_pma_interface_pma_done_counter = 18'b101010101110011000,
		parameter hssi_common_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_common_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_common_pcs_pma_interface_ppm_cnt_rst = "ppm_cnt_rst_dis", // ppm_cnt_rst_dis|ppm_cnt_rst_en
		parameter hssi_common_pcs_pma_interface_ppm_deassert_early = "deassert_early_dis", // deassert_early_dis|deassert_early_en
		parameter hssi_common_pcs_pma_interface_ppm_det_buckets = "ppm_100_bucket", // disable_prot|ppm_300_bucket|ppm_100_bucket|ppm_300_100_bucket
		parameter hssi_common_pcs_pma_interface_ppm_gen1_2_cnt = "cnt_32k", // cnt_32k|cnt_64k
		parameter hssi_common_pcs_pma_interface_ppm_post_eidle_delay = "cnt_200_cycles", // cnt_200_cycles|cnt_400_cycles
		parameter hssi_common_pcs_pma_interface_ppmsel = "ppmsel_300", // ppmsel_disable|ppmsel_5000|ppmsel_2500|ppmsel_1000|ppmsel_500|ppmsel_300|ppmsel_250|ppmsel_200|ppmsel_125|ppmsel_100|ppmsel_62p5|ppm_other
		parameter hssi_common_pcs_pma_interface_prot_mode = "disable_prot_mode", // disable_prot_mode|pipe_g12|pipe_g3|other_protocols
		parameter hssi_common_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_common_pcs_pma_interface_rxvalid_mask = "rxvalid_mask_en", // rxvalid_mask_dis|rxvalid_mask_en
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter = 12'b100111000100,
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_sim_mode = "disable", // disable|enable
		parameter hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en = "true", // false|true
		parameter hssi_common_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_common_pcs_pma_interface_testout_sel = "ppm_det_test", // ppm_det_test|asn_test|pma_pll_test|rxpmaif_test|prbs_gen_test|prbs_ver_test|uhsif_1_test|uhsif_2_test|uhsif_3_test
		parameter hssi_common_pcs_pma_interface_wait_clk_on_off_timer = 4'b100,
		parameter hssi_common_pcs_pma_interface_wait_pipe_synchronizing = 5'b10111,
		parameter hssi_common_pcs_pma_interface_wait_send_syncp_fbkp = 11'b11111010,
		
		// parameters for twentynm_hssi_common_pld_pcs_interface
		parameter hssi_common_pld_pcs_interface_dft_clk_out_en = "dft_clk_out_disable", // dft_clk_out_disable|dft_clk_out_enable
		parameter hssi_common_pld_pcs_interface_dft_clk_out_sel = "teng_rx_dft_clk", // teng_rx_dft_clk|teng_tx_dft_clk|eightg_rx_dft_clk|eightg_tx_dft_clk|pmaif_dft_clk
		parameter hssi_common_pld_pcs_interface_hrdrstctrl_en = "hrst_dis", // hrst_dis|hrst_en
		parameter hssi_common_pld_pcs_interface_pcs_testbus_block_sel = "eightg", // eightg|g3pcs|teng|krfec|pma_if
		parameter hssi_common_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_fifo_rx_pcs
		parameter hssi_fifo_rx_pcs_double_read_mode = "double_read_dis", // double_read_en|double_read_dis
		parameter hssi_fifo_rx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_fifo_tx_pcs
		parameter hssi_fifo_tx_pcs_double_write_mode = "double_write_dis", // double_write_en|double_write_dis
		parameter hssi_fifo_tx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_gen3_rx_pcs
		parameter hssi_gen3_rx_pcs_block_sync = "enable_block_sync", // bypass_block_sync|enable_block_sync
		parameter hssi_gen3_rx_pcs_block_sync_sm = "enable_blk_sync_sm", // disable_blk_sync_sm|enable_blk_sync_sm
		parameter hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn = "enable", // disable|enable
		parameter hssi_gen3_rx_pcs_lpbk_force = "lpbk_frce_dis", // lpbk_frce_dis|lpbk_frce_en
		parameter hssi_gen3_rx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_rx_pcs_rate_match_fifo = "enable_rm_fifo_600ppm", // bypass_rm_fifo|enable_rm_fifo_600ppm|enable_rm_fifo_0ppm
		parameter hssi_gen3_rx_pcs_rate_match_fifo_latency = "regular_latency", // regular_latency|low_latency
		parameter hssi_gen3_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_gen3_rx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_b4gb_par_lpbk = "b4gb_par_lpbk_dis", // b4gb_par_lpbk_dis|b4gb_par_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_force_balign = "en_force_balign", // en_force_balign|dis_force_balign
		parameter hssi_gen3_rx_pcs_rx_ins_del_one_skip = "ins_del_one_skip_en", // ins_del_one_skip_dis|ins_del_one_skip_en
		parameter hssi_gen3_rx_pcs_rx_num_fixed_pat = 4'b1000,
		parameter hssi_gen3_rx_pcs_rx_test_out_sel = "rx_test_out0", // rx_test_out0|rx_test_out1
		parameter hssi_gen3_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_gen3_tx_pcs
		parameter hssi_gen3_tx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_tx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_gen3_tx_pcs_tx_bitslip = 5'b0,
		parameter hssi_gen3_tx_pcs_tx_gbox_byp = "bypass_gbox", // bypass_gbox|enable_gbox
		
		// parameters for twentynm_hssi_krfec_rx_pcs
		parameter hssi_krfec_rx_pcs_blksync_cor_en = "detect", // detect|correct
		parameter hssi_krfec_rx_pcs_bypass_gb = "bypass_dis", // bypass_dis|bypass_en
		parameter hssi_krfec_rx_pcs_clr_ctrl = "both_enabled", // both_enabled|corr_cnt_only|uncorr_cnt_only
		parameter hssi_krfec_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_rx_pcs_dv_start = "with_blklock", // with_blksync|with_blklock
		parameter hssi_krfec_rx_pcs_err_mark_type = "err_mark_10g", // err_mark_10g|err_mark_40g
		parameter hssi_krfec_rx_pcs_error_marking_en = "err_mark_dis", // err_mark_dis|err_mark_en
		parameter hssi_krfec_rx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_krfec_rx_pcs_parity_invalid_enum = 8'b1000,
		parameter hssi_krfec_rx_pcs_parity_valid_num = 4'b100,
		parameter hssi_krfec_rx_pcs_pipeln_blksync = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_descrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errcorrect = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_ind = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_lfsr = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_loc = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_pat = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_gearbox = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_syndrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_trans_dec = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_rx_pcs_receive_order = "receive_lsb", // receive_lsb|receive_msb
		parameter hssi_krfec_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_krfec_rx_pcs_rx_testbus_sel = "overall", // overall|fast_search|fast_search_cntrs|blksync|blksync_cntrs|decoder_master_sm|decoder_master_sm_cntrs|syndrm_sm|syndrm1|syndrm2|errtrap_sm|errtrap_ind1|errtrap_ind2|errtrap_ind3|errtrap_ind4|errtrap_ind5|errtrap_loc|errtrap_pat1|errtrap_pat2|errtrap_pat3|errtrap_pat4|decoder_rd_sm|gb_and_trans
		parameter hssi_krfec_rx_pcs_signal_ok_en = "sig_ok_dis", // sig_ok_dis|sig_ok_en
		parameter hssi_krfec_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_krfec_tx_pcs
		parameter hssi_krfec_tx_pcs_burst_err = "burst_err_dis", // burst_err_dis|burst_err_en
		parameter hssi_krfec_tx_pcs_burst_err_len = "burst_err_len1", // burst_err_len1|burst_err_len2|burst_err_len3|burst_err_len4|burst_err_len5|burst_err_len6|burst_err_len7|burst_err_len8|burst_err_len9|burst_err_len10|burst_err_len11|burst_err_len12|burst_err_len13|burst_err_len14|burst_err_len15|burst_err_len16
		parameter hssi_krfec_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_tx_pcs_enc_frame_query = "enc_query_dis", // enc_query_dis|enc_query_en
		parameter hssi_krfec_tx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_encoder = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_scrambler = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_krfec_tx_pcs_transcode_err = "trans_err_dis", // trans_err_dis|trans_err_en
		parameter hssi_krfec_tx_pcs_transmit_order = "transmit_lsb", // transmit_lsb|transmit_msb
		parameter hssi_krfec_tx_pcs_tx_testbus_sel = "overall", // overall|encoder1|encoder2|scramble1|scramble2|scramble3|gearbox
		
		// parameters for twentynm_hssi_pipe_gen1_2
		parameter hssi_pipe_gen1_2_elec_idle_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_error_replace_pad = "replace_edb", // replace_edb|replace_pad
		parameter hssi_pipe_gen1_2_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_pipe_gen1_2_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen1_2_phystatus_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_phystatus_rst_toggle = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen1_2_pipe_byte_de_serializer_en = "dont_care_bds", // dis_bds|en_bds_by_2|dont_care_bds
		parameter hssi_pipe_gen1_2_prot_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|basic|disabled_prot_mode
		parameter hssi_pipe_gen1_2_reconfig_settings = "{}", // 
		parameter hssi_pipe_gen1_2_rx_pipe_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_pipe_gen1_2_rxdetect_bypass = "dis_rxdetect_bypass", // dis_rxdetect_bypass|en_rxdetect_bypass
		parameter hssi_pipe_gen1_2_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen1_2_tx_pipe_enable = "dis_pipe_tx", // dis_pipe_tx|en_pipe_tx|en_pipe3_tx
		parameter hssi_pipe_gen1_2_txswing = "dis_txswing", // dis_txswing|en_txswing
		
		// parameters for twentynm_hssi_pipe_gen3
		parameter hssi_pipe_gen3_bypass_rx_detection_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_rx_preset = 3'b0,
		parameter hssi_pipe_gen3_bypass_rx_preset_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_tx_coefficent = 18'b0,
		parameter hssi_pipe_gen3_bypass_tx_coefficent_enable = "false", // false|true
		parameter hssi_pipe_gen3_elecidle_delay_g3 = 3'b110,
		parameter hssi_pipe_gen3_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen3_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|disable_pcs
		parameter hssi_pipe_gen3_phy_status_delay_g12 = 3'b101,
		parameter hssi_pipe_gen3_phy_status_delay_g3 = 3'b101,
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g12 = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g3 = "dis_phystatus_rst_toggle_g3", // dis_phystatus_rst_toggle_g3|en_phystatus_rst_toggle_g3
		parameter hssi_pipe_gen3_rate_match_pad_insertion = "dis_rm_fifo_pad_ins", // dis_rm_fifo_pad_ins|en_rm_fifo_pad_ins
		parameter hssi_pipe_gen3_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen3_test_out_sel = "disable_test_out", // tx_test_out|rx_test_out|pipe_test_out1|pipe_test_out2|pipe_test_out3|pipe_ctrl_test_out|disable_test_out
		
		// parameters for twentynm_hssi_rx_pcs_pma_interface
		parameter hssi_rx_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|ten_g_pcs|direct_pld
		parameter hssi_rx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pcs_pma_interface_clkslip_sel = "pld", // pld|slip_eight_g_pcs
		parameter hssi_rx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pcs_pma_interface_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_rx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_rx_pcs_pma_interface_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_rx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_rx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_rx_pcs_pma_interface_prbs_ver = "prbs_off", // prbs_off|prbs_31|prbs_15|prbs_23|prbs_9|prbs_7
		parameter hssi_rx_pcs_pma_interface_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion = "rx_dyn_polinv_dis", // rx_dyn_polinv_dis|rx_dyn_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_lpbk_en = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok = "unforce_sig_ok", // unforce_sig_ok|force_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mask = "prbsmask128", // prbsmask128|prbsmask256|prbsmask512|prbsmask1024
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mode = "teng_mode", // teng_mode|eightg_mode
		parameter hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel = "sel_sig_det", // sel_sig_det|sel_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_static_polarity_inversion = "rx_stat_polinv_dis", // rx_stat_polinv_dis|rx_stat_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en = "uhsif_lpbk_dis", // uhsif_lpbk_dis|uhsif_lpbk_en
		parameter hssi_rx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_rx_pld_pcs_interface
		parameter hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx = "enable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx = "pma_64b_rx", // pma_32b_rx|pma_40b_rx|pma_64b_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_baser_mode_rx|interlaken_mode_rx|sfis_mode_rx|teng_sdi_mode_rx|basic_mode_rx|test_prp_mode_rx|test_prp_krfec_mode_rx|teng_1588_mode_rx|teng_baser_krfec_mode_rx|teng_1588_krfec_mode_rx|basic_krfec_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx = "disabled_prot_mode_rx", // pipe_g1_rx|pipe_g2_rx|pipe_g3_rx|cpri_rx|cpri_rx_tx_rx|gige_rx|gige_1588_rx|basic_rm_enable_rx|basic_rm_disable_rx|disabled_prot_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcie_g1_capable_rx|pcie_g2_capable_rx|pcie_g3_capable_rx|gige_rx|teng_baser_rx|teng_basekr_krfec_rx|fortyg_basekr_krfec_rx|cpri_8b10b_rx|interlaken_rx|sfis_rx|teng_sdi_rx|gige_1588_rx|teng_1588_baser_rx|teng_1588_basekr_krfec_rx|basic_8gpcs_rm_enable_rx|basic_8gpcs_rm_disable_rx|basic_10gpcs_rx|basic_10gpcs_krfec_rx|pcs_direct_rx|prp_rx|prp_krfec_rx|prbs_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx = "teng_mode_rx", // teng_mode_rx|non_teng_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_basekr_mode_rx|fortyg_basekr_mode_rx|teng_1588_basekr_mode_rx|basic_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|eightg_and_g3_pld_fifo_mode_rx|eightg_and_g3_reg_mode_rx|eightg_and_g3_reg_mode_hip_rx|teng_pld_fifo_mode_rx|teng_reg_mode_rx|teng_and_krfec_pld_fifo_mode_rx|teng_and_krfec_reg_mode_rx|pcs_direct_reg_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_block_sel = "pcs_direct", // eightg|teng|pcs_direct
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_rx_clk|pma_rx_clk_user
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_sel = "pld_rx_clk", // pld_rx_clk|pcs_rx_clk
		parameter hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en = "hip_rx_enable", // hip_rx_enable|hip_rx_disable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_rx_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_tx_pcs_pma_interface
		parameter hssi_tx_pcs_pma_interface_bypass_pma_txelecidle = "false", // false|true
		parameter hssi_tx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pcs_pma_interface_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx = "other_prot_mode", // pipe_g12|pipe_g3|other_prot_mode
		parameter hssi_tx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_tx_pcs_pma_interface_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_tx_pcs_pma_interface_pmagate_en = "pmagate_dis", // pmagate_dis|pmagate_en
		parameter hssi_tx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_tx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_tx_pcs_pma_interface_prbs_gen_pat = "prbs_gen_dis", // prbs_gen_dis|prbs_31|prbs_23|prbs_15|prbs_9|prbs_7
		parameter hssi_tx_pcs_pma_interface_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_tx_pcs_pma_interface_sq_wave_num = "sq_wave_4", // sq_wave_1|sq_wave_4|sq_wave_8|sq_wave_6|sq_wave_default
		parameter hssi_tx_pcs_pma_interface_sqwgen_clken = "sqwgen_clk_dis", // sqwgen_clk_dis|sqwgen_clk_en
		parameter hssi_tx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion = "tx_dyn_polinv_dis", // tx_dyn_polinv_dis|tx_dyn_polinv_en
		parameter hssi_tx_pcs_pma_interface_tx_pma_data_sel = "pld_dir", // pld_dir|pcie_gen3|eight_g_pcs|ten_g_pcs|prbs_pat|sq_wave_pat|block_sel_default|registered_uhsif_dat|directed_uhsif_dat
		parameter hssi_tx_pcs_pma_interface_tx_static_polarity_inversion = "tx_stat_polinv_dis", // tx_stat_polinv_dis|tx_stat_polinv_en
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock = "uhsif_filt_stepsz_b4lock_4", // uhsif_filt_stepsz_b4lock_2|uhsif_filt_stepsz_b4lock_4|uhsif_filt_stepsz_b4lock_6|uhsif_filt_stepsz_b4lock_8
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value = 4'b1011,
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock = "uhsif_filt_cntthr_b4lock_16", // uhsif_filt_cntthr_b4lock_8|uhsif_filt_cntthr_b4lock_16|uhsif_filt_cntthr_b4lock_24|uhsif_filt_cntthr_b4lock_32
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period = "uhsif_dcn_test_period_4", // uhsif_dcn_test_period_4|uhsif_dcn_test_period_8|uhsif_dcn_test_period_12|uhsif_dcn_test_period_16
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable = "uhsif_dcn_test_mode_disable", // uhsif_dcn_test_mode_enable|uhsif_dcn_test_mode_disable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh = "uhsif_dzt_cnt_thr_4", // uhsif_dzt_cnt_thr_2|uhsif_dzt_cnt_thr_4|uhsif_dzt_cnt_thr_6|uhsif_dzt_cnt_thr_8
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable = "uhsif_dzt_enable", // uhsif_dzt_disable|uhsif_dzt_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window = "uhsif_dzt_obr_win_32", // uhsif_dzt_obr_win_16|uhsif_dzt_obr_win_32|uhsif_dzt_obr_win_48|uhsif_dzt_obr_win_64
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size = "uhsif_dzt_skipsz_8", // uhsif_dzt_skipsz_4|uhsif_dzt_skipsz_8|uhsif_dzt_skipsz_12|uhsif_dzt_skipsz_16
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel = "uhsif_index_internal", // uhsif_index_internal|uhsif_index_cram
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin = "uhsif_dcn_margin_4", // uhsif_dcn_margin_2|uhsif_dcn_margin_3|uhsif_dcn_margin_4|uhsif_dcn_margin_5
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value = 8'b10000000,
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control = "uhsif_dft_dz_det_val_0", // uhsif_dft_dz_det_val_0|uhsif_dft_dz_det_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control = "uhsif_dft_up_val_0", // uhsif_dft_up_val_0|uhsif_dft_up_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_enable = "uhsif_disable", // uhsif_disable|uhsif_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock = "uhsif_lkd_segsz_aflock_2048", // uhsif_lkd_segsz_aflock_512|uhsif_lkd_segsz_aflock_1024|uhsif_lkd_segsz_aflock_2048|uhsif_lkd_segsz_aflock_4096
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock = "uhsif_lkd_segsz_b4lock_32", // uhsif_lkd_segsz_b4lock_16|uhsif_lkd_segsz_b4lock_32|uhsif_lkd_segsz_b4lock_64|uhsif_lkd_segsz_b4lock_128
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value = 4'b11,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value = 4'b11,
		
		// parameters for twentynm_hssi_tx_pld_pcs_interface
		parameter hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx = "enable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx = "pma_64b_tx", // pma_32b_tx|pma_40b_tx|pma_64b_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_baser_mode_tx|interlaken_mode_tx|sfis_mode_tx|teng_sdi_mode_tx|basic_mode_tx|test_prp_mode_tx|test_prp_krfec_mode_tx|teng_1588_mode_tx|teng_baser_krfec_mode_tx|teng_1588_krfec_mode_tx|basic_krfec_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx = "disabled_prot_mode_tx", // pipe_g1_tx|pipe_g2_tx|pipe_g3_tx|cpri_tx|cpri_rx_tx_tx|gige_tx|gige_1588_tx|basic_tx|disabled_prot_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcie_g1_capable_tx|pcie_g2_capable_tx|pcie_g3_capable_tx|gige_tx|teng_baser_tx|teng_basekr_krfec_tx|fortyg_basekr_krfec_tx|cpri_8b10b_tx|interlaken_tx|sfis_tx|teng_sdi_tx|gige_1588_tx|teng_1588_baser_tx|teng_1588_basekr_krfec_tx|basic_8gpcs_tx|basic_10gpcs_tx|basic_10gpcs_krfec_tx|pcs_direct_tx|uhsif_tx|prp_tx|prp_krfec_tx|prbs_tx|sqwave_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx = "teng_mode_tx", // teng_mode_tx|non_teng_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_basekr_mode_tx|fortyg_basekr_mode_tx|teng_1588_basekr_mode_tx|basic_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|eightg_and_g3_pld_fifo_mode_tx|eightg_and_g3_reg_mode_tx|eightg_and_g3_reg_mode_hip_tx|eightg_and_g3_fastreg_mode_tx|teng_pld_fifo_mode_tx|teng_reg_mode_tx|teng_fastreg_mode_tx|teng_and_krfec_pld_fifo_mode_tx|teng_and_krfec_reg_mode_tx|teng_and_krfec_fastreg_mode_tx|pcs_direct_fastreg_mode_tx|uhsif_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_tx_clk|pma_tx_clk_user
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_source = "teng", // eightg|teng|pma_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_data_source = "hip_disable", // hip_disable|hip_enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en = "delay1_clk_disable", // delay1_clk_enable|delay1_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel = "pld_tx_clk", // pld_tx_clk|pcs_tx_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl = "delay1_path0", // delay1_path0|delay1_path1|delay1_path2|delay1_path3|delay1_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel = "one_ff_delay", // one_ff_delay|two_ff_delay
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en = "delay2_clk_disable", // delay2_clk_enable|delay2_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl = "delay2_path0", // delay2_path0|delay2_path1|delay2_path2|delay2_path3|delay2_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_tx_pld_pcs_interface_reconfig_settings = "{}" // 
	//PARAM_LIST_END
	)
	(
	//PORT_LIST_START
		input wire	[8:0]	in_avmmaddress,
		input wire		in_avmmclk,
		input wire		in_avmmread,
		input wire		in_avmmrstn,
		input wire		in_avmmwrite,
		input wire	[7:0]	in_avmmwritedata,
		input wire	[4:0]	in_bond_pcs10g_in_bot,
		input wire	[4:0]	in_bond_pcs10g_in_top,
		input wire	[12:0]	in_bond_pcs8g_in_bot,
		input wire	[12:0]	in_bond_pcs8g_in_top,
		input wire	[11:0]	in_bond_pmaif_in_bot,
		input wire	[11:0]	in_bond_pmaif_in_top,
		input wire	[63:0]	in_hip_tx_data,
		input wire		in_iocsr_clk,
		input wire	[5:0]	in_iocsr_config,
		input wire		in_iocsr_rdy,
		input wire		in_iocsr_rdy_dly,
		input wire		in_pld_10g_krfec_rx_clr_errblk_cnt,
		input wire		in_pld_10g_krfec_rx_pld_rst_n,
		input wire		in_pld_10g_krfec_tx_pld_rst_n,
		input wire		in_pld_10g_rx_align_clr,
		input wire		in_pld_10g_rx_clr_ber_count,
		input wire		in_pld_10g_rx_rd_en,
		input wire	[6:0]	in_pld_10g_tx_bitslip,
		input wire		in_pld_10g_tx_burst_en,
		input wire		in_pld_10g_tx_data_valid,
		input wire	[1:0]	in_pld_10g_tx_diag_status,
		input wire		in_pld_10g_tx_wordslip,
		input wire		in_pld_8g_a1a2_size,
		input wire		in_pld_8g_bitloc_rev_en,
		input wire		in_pld_8g_byte_rev_en,
		input wire	[2:0]	in_pld_8g_eidleinfersel,
		input wire		in_pld_8g_encdt,
		input wire		in_pld_8g_g3_rx_pld_rst_n,
		input wire		in_pld_8g_g3_tx_pld_rst_n,
		input wire		in_pld_8g_rddisable_tx,
		input wire		in_pld_8g_rdenable_rx,
		input wire		in_pld_8g_refclk_dig2,
		input wire		in_pld_8g_rxpolarity,
		input wire	[4:0]	in_pld_8g_tx_boundary_sel,
		input wire		in_pld_8g_wrdisable_rx,
		input wire		in_pld_8g_wrenable_tx,
		input wire		in_pld_atpg_los_en_n,
		input wire		in_pld_bitslip,
		input wire	[17:0]	in_pld_g3_current_coeff,
		input wire	[2:0]	in_pld_g3_current_rxpreset,
		input wire		in_pld_ltr,
		input wire		in_pld_mem_krfec_atpg_rst_n,
		input wire		in_pld_partial_reconfig,
		input wire		in_pld_pcs_refclk_dig,
		input wire		in_pld_pma_adapt_start,
		input wire		in_pld_pma_csr_test_dis,
		input wire		in_pld_pma_early_eios,
		input wire	[5:0]	in_pld_pma_eye_monitor,
		input wire		in_pld_pma_ltd_b,
		input wire		in_pld_pma_nrpi_freeze,
		input wire	[1:0]	in_pld_pma_pcie_switch,
		input wire		in_pld_pma_ppm_lock,
		input wire	[4:0]	in_pld_pma_reserved_out,
		input wire		in_pld_pma_rs_lpbk_b,
		input wire		in_pld_pma_rx_qpi_pullup,
		input wire		in_pld_pma_rxpma_rstb,
		input wire		in_pld_pma_tx_bitslip,
		input wire		in_pld_pma_tx_bonding_rstb,
		input wire		in_pld_pma_tx_qpi_pulldn,
		input wire		in_pld_pma_tx_qpi_pullup,
		input wire		in_pld_pma_txdetectrx,
		input wire		in_pld_pma_txpma_rstb,
		input wire		in_pld_pmaif_rx_pld_rst_n,
		input wire		in_pld_pmaif_rxclkslip,
		input wire		in_pld_pmaif_tx_pld_rst_n,
		input wire		in_pld_polinv_rx,
		input wire		in_pld_polinv_tx,
		input wire	[1:0]	in_pld_rate,
		input wire	[9:0]	in_pld_reserved_in,
		input wire		in_pld_rx_clk,
		input wire		in_pld_rx_prbs_err_clr,
		input wire		in_pld_scan_mode_n,
		input wire		in_pld_scan_shift_n,
		input wire		in_pld_syncsm_en,
		input wire		in_pld_tx_clk,
		input wire	[17:0]	in_pld_tx_control,
		input wire	[127:0]	in_pld_tx_data,
		input wire		in_pld_txelecidle,
		input wire		in_pld_uhsif_tx_clk,
		input wire		in_pma_adapt_done,
		input wire		in_pma_clklow,
		input wire		in_pma_fref,
		input wire		in_pma_hclk,
		input wire	[1:0]	in_pma_pcie_sw_done,
		input wire		in_pma_pfdmode_lock,
		input wire	[4:0]	in_pma_reserved_in,
		input wire		in_pma_rx_clkdiv_user,
		input wire		in_pma_rx_detect_valid,
		input wire		in_pma_rx_found,
		input wire		in_pma_rx_pma_clk,
		input wire	[63:0]	in_pma_rx_pma_data,
		input wire		in_pma_rx_signal_ok,
		input wire		in_pma_rxpll_lock,
		input wire		in_pma_signal_det,
		input wire	[7:0]	in_pma_testbus,
		input wire		in_pma_tx_clkdiv_user,
		input wire		in_pma_tx_pma_clk,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen1_2,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen3,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pld_pcs_interface,
		output wire		out_blockselect_hssi_10g_rx_pcs,
		output wire		out_blockselect_hssi_10g_tx_pcs,
		output wire		out_blockselect_hssi_8g_rx_pcs,
		output wire		out_blockselect_hssi_8g_tx_pcs,
		output wire		out_blockselect_hssi_common_pcs_pma_interface,
		output wire		out_blockselect_hssi_common_pld_pcs_interface,
		output wire		out_blockselect_hssi_fifo_rx_pcs,
		output wire		out_blockselect_hssi_fifo_tx_pcs,
		output wire		out_blockselect_hssi_gen3_rx_pcs,
		output wire		out_blockselect_hssi_gen3_tx_pcs,
		output wire		out_blockselect_hssi_krfec_rx_pcs,
		output wire		out_blockselect_hssi_krfec_tx_pcs,
		output wire		out_blockselect_hssi_pipe_gen1_2,
		output wire		out_blockselect_hssi_pipe_gen3,
		output wire		out_blockselect_hssi_rx_pcs_pma_interface,
		output wire		out_blockselect_hssi_rx_pld_pcs_interface,
		output wire		out_blockselect_hssi_tx_pcs_pma_interface,
		output wire		out_blockselect_hssi_tx_pld_pcs_interface,
		output wire	[4:0]	out_bond_pcs10g_out_bot,
		output wire	[4:0]	out_bond_pcs10g_out_top,
		output wire	[12:0]	out_bond_pcs8g_out_bot,
		output wire	[12:0]	out_bond_pcs8g_out_top,
		output wire	[11:0]	out_bond_pmaif_out_bot,
		output wire	[11:0]	out_bond_pmaif_out_top,
		output wire	[2:0]	out_hip_clk_out,
		output wire	[7:0]	out_hip_ctrl_out,
		output wire		out_hip_iocsr_rdy,
		output wire		out_hip_iocsr_rdy_dly,
		output wire		out_hip_nfrzdrv,
		output wire		out_hip_npor,
		output wire	[50:0]	out_hip_rx_data,
		output wire		out_hip_usermode,
		output wire		out_pld_10g_krfec_rx_blk_lock,
		output wire	[1:0]	out_pld_10g_krfec_rx_diag_data_status,
		output wire		out_pld_10g_krfec_rx_frame,
		output wire		out_pld_10g_krfec_tx_frame,
		output wire		out_pld_10g_rx_align_val,
		output wire		out_pld_10g_rx_crc32_err,
		output wire		out_pld_10g_rx_data_valid,
		output wire		out_pld_10g_rx_empty,
		output wire		out_pld_10g_rx_fifo_del,
		output wire		out_pld_10g_rx_fifo_insert,
		output wire	[4:0]	out_pld_10g_rx_fifo_num,
		output wire		out_pld_10g_rx_frame_lock,
		output wire		out_pld_10g_rx_hi_ber,
		output wire		out_pld_10g_rx_oflw_err,
		output wire		out_pld_10g_rx_pempty,
		output wire		out_pld_10g_rx_pfull,
		output wire		out_pld_10g_tx_burst_en_exe,
		output wire		out_pld_10g_tx_empty,
		output wire	[3:0]	out_pld_10g_tx_fifo_num,
		output wire		out_pld_10g_tx_full,
		output wire		out_pld_10g_tx_pempty,
		output wire		out_pld_10g_tx_pfull,
		output wire		out_pld_10g_tx_wordslip_exe,
		output wire	[3:0]	out_pld_8g_a1a2_k1k2_flag,
		output wire		out_pld_8g_empty_rmf,
		output wire		out_pld_8g_empty_rx,
		output wire		out_pld_8g_empty_tx,
		output wire		out_pld_8g_full_rmf,
		output wire		out_pld_8g_full_rx,
		output wire		out_pld_8g_full_tx,
		output wire		out_pld_8g_rxelecidle,
		output wire		out_pld_8g_signal_detect_out,
		output wire	[4:0]	out_pld_8g_wa_boundary,
		output wire		out_pld_krfec_tx_alignment,
		output wire		out_pld_pcs_rx_clk_out,
		output wire		out_pld_pcs_tx_clk_out,
		output wire		out_pld_pma_adapt_done,
		output wire		out_pld_pma_clkdiv_rx_user,
		output wire		out_pld_pma_clkdiv_tx_user,
		output wire		out_pld_pma_clklow,
		output wire		out_pld_pma_fref,
		output wire		out_pld_pma_hclk,
		output wire	[1:0]	out_pld_pma_pcie_sw_done,
		output wire		out_pld_pma_pfdmode_lock,
		output wire	[4:0]	out_pld_pma_reserved_in,
		output wire		out_pld_pma_rx_clk_out,
		output wire		out_pld_pma_rx_detect_valid,
		output wire		out_pld_pma_rx_found,
		output wire		out_pld_pma_rxpll_lock,
		output wire		out_pld_pma_signal_ok,
		output wire	[7:0]	out_pld_pma_testbus,
		output wire		out_pld_pma_tx_clk_out,
		output wire		out_pld_pmaif_mask_tx_pll,
		output wire	[9:0]	out_pld_reserved_out,
		output wire	[19:0]	out_pld_rx_control,
		output wire	[127:0]	out_pld_rx_data,
		output wire		out_pld_rx_prbs_done,
		output wire		out_pld_rx_prbs_err,
		output wire	[19:0]	out_pld_test_data,
		output wire		out_pld_uhsif_lock,
		output wire		out_pld_uhsif_tx_clk_out,
		output wire		out_pma_adapt_start,
		output wire		out_pma_atpg_los_en_n,
		output wire		out_pma_csr_test_dis,
		output wire	[17:0]	out_pma_current_coeff,
		output wire	[2:0]	out_pma_current_rxpreset,
		output wire		out_pma_early_eios,
		output wire	[5:0]	out_pma_eye_monitor,
		output wire	[1:0]	out_pma_interface_select,
		output wire		out_pma_ltd_b,
		output wire		out_pma_ltr,
		output wire		out_pma_nfrzdrv,
		output wire		out_pma_nrpi_freeze,
		output wire	[1:0]	out_pma_pcie_switch,
		output wire		out_pma_ppm_lock,
		output wire	[4:0]	out_pma_reserved_out,
		output wire		out_pma_rs_lpbk_b,
		output wire		out_pma_rx_clkslip,
		output wire		out_pma_rx_qpi_pullup,
		output wire		out_pma_rxpma_rstb,
		output wire		out_pma_scan_mode_n,
		output wire		out_pma_scan_shift_n,
		output wire		out_pma_tx_bitslip,
		output wire		out_pma_tx_bonding_rstb,
		output wire		out_pma_tx_elec_idle,
		output wire	[63:0]	out_pma_tx_pma_data,
		output wire		out_pma_tx_qpi_pulldn,
		output wire		out_pma_tx_qpi_pullup,
		output wire		out_pma_tx_txdetectrx,
		output wire		out_pma_txpma_rstb
	//PORT_LIST_END
	);
	//wire declarations
	
	// wires for module twentynm_hssi_fifo_tx_pcs
	wire	[7:0]	w_hssi_fifo_tx_pcs_avmmreaddata;
	wire		w_hssi_fifo_tx_pcs_blockselect;
	wire	[72:0]	w_hssi_fifo_tx_pcs_data_out_10g;
	wire	[63:0]	w_hssi_fifo_tx_pcs_data_out_8g_phase_comp;
	
	// wires for module twentynm_hssi_gen3_rx_pcs
	wire	[7:0]	w_hssi_gen3_rx_pcs_avmmreaddata;
	wire		w_hssi_gen3_rx_pcs_blk_algnd_int;
	wire		w_hssi_gen3_rx_pcs_blk_start;
	wire		w_hssi_gen3_rx_pcs_blockselect;
	wire		w_hssi_gen3_rx_pcs_clkcomp_delete_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_insert_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_overfl_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_undfl_int;
	wire	[31:0]	w_hssi_gen3_rx_pcs_data_out;
	wire		w_hssi_gen3_rx_pcs_data_valid;
	wire		w_hssi_gen3_rx_pcs_ei_det_int;
	wire		w_hssi_gen3_rx_pcs_ei_partial_det_int;
	wire		w_hssi_gen3_rx_pcs_err_decode_int;
	wire		w_hssi_gen3_rx_pcs_i_det_int;
	wire		w_hssi_gen3_rx_pcs_lpbk_blk_start;
	wire	[33:0]	w_hssi_gen3_rx_pcs_lpbk_data;
	wire		w_hssi_gen3_rx_pcs_lpbk_data_valid;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk;
	wire	[39:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n;
	wire		w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int;
	wire	[19:0]	w_hssi_gen3_rx_pcs_rx_test_out;
	wire	[1:0]	w_hssi_gen3_rx_pcs_sync_hdr;
	
	// wires for module twentynm_hssi_krfec_tx_pcs
	wire	[7:0]	w_hssi_krfec_tx_pcs_avmmreaddata;
	wire		w_hssi_krfec_tx_pcs_blockselect;
	wire		w_hssi_krfec_tx_pcs_tx_alignment;
	wire	[63:0]	w_hssi_krfec_tx_pcs_tx_data_out;
	wire		w_hssi_krfec_tx_pcs_tx_frame;
	wire	[19:0]	w_hssi_krfec_tx_pcs_tx_test_data;
	
	// wires for module twentynm_hssi_krfec_rx_pcs
	wire	[7:0]	w_hssi_krfec_rx_pcs_avmmreaddata;
	wire		w_hssi_krfec_rx_pcs_blockselect;
	wire		w_hssi_krfec_rx_pcs_rx_block_lock;
	wire	[9:0]	w_hssi_krfec_rx_pcs_rx_control_out;
	wire	[63:0]	w_hssi_krfec_rx_pcs_rx_data_out;
	wire	[1:0]	w_hssi_krfec_rx_pcs_rx_data_status;
	wire		w_hssi_krfec_rx_pcs_rx_data_valid_out;
	wire		w_hssi_krfec_rx_pcs_rx_frame;
	wire		w_hssi_krfec_rx_pcs_rx_signal_ok_out;
	
	// wires for module twentynm_hssi_rx_pld_pcs_interface
	wire	[7:0]	w_hssi_rx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_rx_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_hip_rx_ctrl;
	wire	[50:0]	w_hssi_rx_pld_pcs_interface_hip_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
	wire	[3:0]	w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary;
	wire		w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_pld_rx_control;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_pld_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
	
	// wires for module twentynm_hssi_common_pld_pcs_interface
	wire	[7:0]	w_hssi_common_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_common_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_hip_cmn_clk;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_hip_cmn_ctrl;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
	wire		w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_hip_npor;
	wire		w_hssi_common_pld_pcs_interface_hip_usermode;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n;
	wire	[17:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel;
	wire		w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_clklow;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_fref;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_hclk;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_pld_pma_reserved_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
	wire	[7:0]	w_hssi_common_pld_pcs_interface_pld_pma_testbus;
	wire		w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
	wire	[9:0]	w_hssi_common_pld_pcs_interface_pld_reserved_out;
	wire	[19:0]	w_hssi_common_pld_pcs_interface_pld_test_data;
	wire		w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
	wire		w_hssi_common_pld_pcs_interface_scan_mode_n;
	
	// wires for module twentynm_hssi_10g_rx_pcs
	wire	[7:0]	w_hssi_10g_rx_pcs_avmmreaddata;
	wire		w_hssi_10g_rx_pcs_blockselect;
	wire		w_hssi_10g_rx_pcs_rx_align_val;
	wire		w_hssi_10g_rx_pcs_rx_blk_lock;
	wire		w_hssi_10g_rx_pcs_rx_clk_out;
	wire		w_hssi_10g_rx_pcs_rx_clk_out_pld_if;
	wire	[19:0]	w_hssi_10g_rx_pcs_rx_control;
	wire		w_hssi_10g_rx_pcs_rx_crc32_err;
	wire	[127:0]	w_hssi_10g_rx_pcs_rx_data;
	wire		w_hssi_10g_rx_pcs_rx_data_valid;
	wire		w_hssi_10g_rx_pcs_rx_dft_clk_out;
	wire	[1:0]	w_hssi_10g_rx_pcs_rx_diag_status;
	wire		w_hssi_10g_rx_pcs_rx_empty;
	wire		w_hssi_10g_rx_pcs_rx_fec_clk;
	wire		w_hssi_10g_rx_pcs_rx_fifo_del;
	wire		w_hssi_10g_rx_pcs_rx_fifo_insert;
	wire	[4:0]	w_hssi_10g_rx_pcs_rx_fifo_num;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_clk;
	wire	[73:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_data;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_en;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_ptr;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_frame_lock;
	wire		w_hssi_10g_rx_pcs_rx_hi_ber;
	wire		w_hssi_10g_rx_pcs_rx_master_clk;
	wire		w_hssi_10g_rx_pcs_rx_master_clk_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_oflw_err;
	wire		w_hssi_10g_rx_pcs_rx_pempty;
	wire		w_hssi_10g_rx_pcs_rx_pfull;
	wire		w_hssi_10g_rx_pcs_rx_random_err;
	wire		w_hssi_10g_rx_pcs_rx_rx_frame;
	
	// wires for module twentynm_hssi_tx_pld_pcs_interface
	wire	[7:0]	w_hssi_tx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_tx_pld_pcs_interface_blockselect;
	wire		w_hssi_tx_pld_pcs_interface_hip_tx_clk;
	wire	[6:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en;
	wire	[17:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control;
	wire	[8:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg;
	wire	[127:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start;
	wire	[4:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle;
	wire	[2:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
	wire		w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
	
	// wires for module twentynm_hssi_tx_pcs_pma_interface
	wire	[7:0]	w_hssi_tx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_tx_pcs_pma_interface_blockselect;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out;
	wire	[4:0]	w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk;
	wire		w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_pma_tx_pma_data;
	wire		w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_1;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_2;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_3;
	
	// wires for module twentynm_hssi_rx_pcs_pma_interface
	wire	[7:0]	w_hssi_rx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_rx_pcs_pma_interface_blockselect;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni;
	wire	[31:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok;
	wire		w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk;
	wire	[5:0]	w_hssi_rx_pcs_pma_interface_pma_eye_monitor;
	wire		w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
	wire		w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test;
	
	// wires for module twentynm_hssi_10g_tx_pcs
	wire	[7:0]	w_hssi_10g_tx_pcs_avmmreaddata;
	wire		w_hssi_10g_tx_pcs_blockselect;
	wire		w_hssi_10g_tx_pcs_distdwn_out_dv;
	wire		w_hssi_10g_tx_pcs_distdwn_out_rden;
	wire		w_hssi_10g_tx_pcs_distdwn_out_wren;
	wire		w_hssi_10g_tx_pcs_distup_out_dv;
	wire		w_hssi_10g_tx_pcs_distup_out_rden;
	wire		w_hssi_10g_tx_pcs_distup_out_wren;
	wire		w_hssi_10g_tx_pcs_tx_burst_en_exe;
	wire		w_hssi_10g_tx_pcs_tx_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pma_if;
	wire	[8:0]	w_hssi_10g_tx_pcs_tx_control_out_krfec;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_data_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_data_valid_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_dft_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_empty;
	wire		w_hssi_10g_tx_pcs_tx_fec_clk;
	wire	[3:0]	w_hssi_10g_tx_pcs_tx_fifo_num;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_rd_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_clk;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_en;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_frame;
	wire		w_hssi_10g_tx_pcs_tx_full;
	wire		w_hssi_10g_tx_pcs_tx_master_clk;
	wire		w_hssi_10g_tx_pcs_tx_master_clk_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_pempty;
	wire		w_hssi_10g_tx_pcs_tx_pfull;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_data;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_gating_val;
	wire	[19:0]	w_hssi_10g_tx_pcs_tx_test_data;
	wire		w_hssi_10g_tx_pcs_tx_wordslip_exe;
	
	// wires for module twentynm_hssi_8g_tx_pcs
	wire	[7:0]	w_hssi_8g_tx_pcs_avmmreaddata;
	wire		w_hssi_8g_tx_pcs_blockselect;
	wire		w_hssi_8g_tx_pcs_clk_out;
	wire		w_hssi_8g_tx_pcs_clk_out_gen3;
	wire	[19:0]	w_hssi_8g_tx_pcs_dataout;
	wire		w_hssi_8g_tx_pcs_dyn_clk_switch_n;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn;
	wire		w_hssi_8g_tx_pcs_g3_tx_pma_rstn;
	wire	[2:0]	w_hssi_8g_tx_pcs_non_gray_eidleinfersel;
	wire		w_hssi_8g_tx_pcs_ph_fifo_overflow;
	wire		w_hssi_8g_tx_pcs_ph_fifo_underflow;
	wire		w_hssi_8g_tx_pcs_phfifo_txdeemph;
	wire	[2:0]	w_hssi_8g_tx_pcs_phfifo_txmargin;
	wire		w_hssi_8g_tx_pcs_phfifo_txswing;
	wire		w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out;
	wire	[1:0]	w_hssi_8g_tx_pcs_pipe_power_down_out;
	wire		w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3;
	wire		w_hssi_8g_tx_pcs_pmaif_asn_rstn;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_refclk_b;
	wire		w_hssi_8g_tx_pcs_refclk_b_reset;
	wire		w_hssi_8g_tx_pcs_rxpolarity_int;
	wire		w_hssi_8g_tx_pcs_soft_reset_wclk1_n;
	wire		w_hssi_8g_tx_pcs_sw_fifo_wr_clk;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_blk_start_out;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_ctrlplane_testbus;
	wire	[31:0]	w_hssi_8g_tx_pcs_tx_data_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_data_valid_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_datak_out;
	wire		w_hssi_8g_tx_pcs_tx_detect_rxloopback_int;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_tx_pipe_clk;
	wire		w_hssi_8g_tx_pcs_tx_pipe_electidle;
	wire		w_hssi_8g_tx_pcs_tx_pipe_soft_reset;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_sync_hdr_out;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_testbus;
	wire		w_hssi_8g_tx_pcs_txcompliance_out;
	wire		w_hssi_8g_tx_pcs_txelecidle_out;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk;
	wire	[63:0]	w_hssi_8g_tx_pcs_wr_data_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_en_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo;
	
	// wires for module twentynm_hssi_pipe_gen3
	wire	[7:0]	w_hssi_pipe_gen3_avmmreaddata;
	wire		w_hssi_pipe_gen3_blockselect;
	wire		w_hssi_pipe_gen3_gen3_clk_sel;
	wire		w_hssi_pipe_gen3_pcs_rst;
	wire		w_hssi_pipe_gen3_phystatus;
	wire	[17:0]	w_hssi_pipe_gen3_pma_current_coeff;
	wire	[2:0]	w_hssi_pipe_gen3_pma_current_rxpreset;
	wire		w_hssi_pipe_gen3_pma_tx_elec_idle;
	wire		w_hssi_pipe_gen3_pma_txdetectrx;
	wire		w_hssi_pipe_gen3_rev_lpbk_8gpcs_out;
	wire		w_hssi_pipe_gen3_rev_lpbk_int;
	wire	[3:0]	w_hssi_pipe_gen3_rx_blk_start;
	wire	[1:0]	w_hssi_pipe_gen3_rx_sync_hdr;
	wire	[63:0]	w_hssi_pipe_gen3_rxd_8gpcs_out;
	wire	[3:0]	w_hssi_pipe_gen3_rxdataskip;
	wire		w_hssi_pipe_gen3_rxelecidle;
	wire		w_hssi_pipe_gen3_rxpolarity_8gpcs_out;
	wire		w_hssi_pipe_gen3_rxpolarity_int;
	wire	[2:0]	w_hssi_pipe_gen3_rxstatus;
	wire		w_hssi_pipe_gen3_rxvalid;
	wire		w_hssi_pipe_gen3_shutdown_clk;
	wire	[19:0]	w_hssi_pipe_gen3_test_out;
	wire		w_hssi_pipe_gen3_tx_blk_start_int;
	wire	[1:0]	w_hssi_pipe_gen3_tx_sync_hdr_int;
	wire	[31:0]	w_hssi_pipe_gen3_txdata_int;
	wire	[3:0]	w_hssi_pipe_gen3_txdatak_int;
	wire		w_hssi_pipe_gen3_txdataskip_int;
	
	// wires for module twentynm_hssi_pipe_gen1_2
	wire	[7:0]	w_hssi_pipe_gen1_2_avmmreaddata;
	wire		w_hssi_pipe_gen1_2_blockselect;
	wire	[17:0]	w_hssi_pipe_gen1_2_current_coeff;
	wire		w_hssi_pipe_gen1_2_phystatus;
	wire		w_hssi_pipe_gen1_2_polarity_inversion_rx;
	wire		w_hssi_pipe_gen1_2_rev_loopbk;
	wire		w_hssi_pipe_gen1_2_rxelecidle;
	wire		w_hssi_pipe_gen1_2_rxelectricalidle_out;
	wire	[2:0]	w_hssi_pipe_gen1_2_rxstatus;
	wire		w_hssi_pipe_gen1_2_rxvalid;
	wire		w_hssi_pipe_gen1_2_tx_elec_idle_out;
	wire		w_hssi_pipe_gen1_2_txdetectrx;
	
	// wires for module twentynm_hssi_gen3_tx_pcs
	wire	[7:0]	w_hssi_gen3_tx_pcs_avmmreaddata;
	wire		w_hssi_gen3_tx_pcs_blockselect;
	wire	[31:0]	w_hssi_gen3_tx_pcs_data_out;
	wire	[35:0]	w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out;
	wire	[31:0]	w_hssi_gen3_tx_pcs_par_lpbk_out;
	wire	[19:0]	w_hssi_gen3_tx_pcs_tx_test_out;
	
	// wires for module twentynm_hssi_8g_rx_pcs
	wire	[3:0]	w_hssi_8g_rx_pcs_a1a2k1k2flag;
	wire	[7:0]	w_hssi_8g_rx_pcs_avmmreaddata;
	wire		w_hssi_8g_rx_pcs_blockselect;
	wire	[19:0]	w_hssi_8g_rx_pcs_chnl_test_bus_out;
	wire		w_hssi_8g_rx_pcs_clock_to_pld;
	wire	[63:0]	w_hssi_8g_rx_pcs_dataout;
	wire		w_hssi_8g_rx_pcs_dis_pc_byte;
	wire		w_hssi_8g_rx_pcs_eidle_detected;
	wire	[2:0]	w_hssi_8g_rx_pcs_eios_det_cdr_ctrl;
	wire		w_hssi_8g_rx_pcs_g3_rx_pma_rstn;
	wire		w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn;
	wire		w_hssi_8g_rx_pcs_gen2ngen1;
	wire	[19:0]	w_hssi_8g_rx_pcs_parallel_rev_loopback;
	wire		w_hssi_8g_rx_pcs_pc_fifo_empty;
	wire		w_hssi_8g_rx_pcs_pcfifofull;
	wire		w_hssi_8g_rx_pcs_phystatus;
	wire	[63:0]	w_hssi_8g_rx_pcs_pipe_data;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_up;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo;
	wire	[7:0]	w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rm_fifo_empty;
	wire		w_hssi_8g_rx_pcs_rm_fifo_full;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_blk_start;
	wire		w_hssi_8g_rx_pcs_rx_clk_out_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clkslip;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_data_valid;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rx_pipe_clk;
	wire		w_hssi_8g_rx_pcs_rx_pipe_soft_reset;
	wire		w_hssi_8g_rx_pcs_rx_pma_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_sync_hdr;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_up;
	wire	[2:0]	w_hssi_8g_rx_pcs_rxstatus;
	wire		w_hssi_8g_rx_pcs_rxvalid;
	wire		w_hssi_8g_rx_pcs_signal_detect_out;
	wire	[4:0]	w_hssi_8g_rx_pcs_word_align_boundary;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk;
	wire	[79:0]	w_hssi_8g_rx_pcs_wr_data_rx_phfifo;
	wire	[31:0]	w_hssi_8g_rx_pcs_wr_data_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo;
	
	// wires for module twentynm_hssi_fifo_rx_pcs
	wire	[7:0]	w_hssi_fifo_rx_pcs_avmmreaddata;
	wire		w_hssi_fifo_rx_pcs_blockselect;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out2_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out_8g_clock_comp;
	wire	[79:0]	w_hssi_fifo_rx_pcs_data_out_8g_phase_comp;
	wire	[39:0]	w_hssi_fifo_rx_pcs_data_out_gen3;
	
	// wires for module twentynm_hssi_common_pcs_pma_interface
	wire	[7:0]	w_hssi_common_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_common_pcs_pma_interface_blockselect;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in;
	wire	[19:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out;
	wire	[7:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus;
	wire		w_hssi_common_pcs_pma_interface_pma_adapt_start;
	wire		w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
	wire		w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
	wire	[17:0]	w_hssi_common_pcs_pma_interface_pma_current_coeff;
	wire	[2:0]	w_hssi_common_pcs_pma_interface_pma_current_rxpreset;
	wire		w_hssi_common_pcs_pma_interface_pma_early_eios;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_interface_select;
	wire		w_hssi_common_pcs_pma_interface_pma_ltd_b;
	wire		w_hssi_common_pcs_pma_interface_pma_ltr;
	wire		w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
	wire		w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_pcie_switch;
	wire		w_hssi_common_pcs_pma_interface_pma_ppm_lock;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_pma_reserved_out;
	wire		w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
	wire		w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up;
	
	
	generate
		
		//module instantiations
		
		// instantiating twentynm_hssi_10g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_rx_pcs
			twentynm_hssi_10g_rx_pcs #(
				.advanced_user_mode(hssi_10g_rx_pcs_advanced_user_mode),
				.align_del(hssi_10g_rx_pcs_align_del),
				.ber_bit_err_total_cnt(hssi_10g_rx_pcs_ber_bit_err_total_cnt),
				.ber_clken(hssi_10g_rx_pcs_ber_clken),
				.ber_xus_timer_window(hssi_10g_rx_pcs_ber_xus_timer_window),
				.bitslip_mode(hssi_10g_rx_pcs_bitslip_mode),
				.blksync_bitslip_type(hssi_10g_rx_pcs_blksync_bitslip_type),
				.blksync_bitslip_wait_cnt(hssi_10g_rx_pcs_blksync_bitslip_wait_cnt),
				.blksync_bitslip_wait_type(hssi_10g_rx_pcs_blksync_bitslip_wait_type),
				.blksync_bypass(hssi_10g_rx_pcs_blksync_bypass),
				.blksync_clken(hssi_10g_rx_pcs_blksync_clken),
				.blksync_enum_invalid_sh_cnt(hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt),
				.blksync_knum_sh_cnt_postlock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock),
				.blksync_knum_sh_cnt_prelock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock),
				.blksync_pipeln(hssi_10g_rx_pcs_blksync_pipeln),
				.clr_errblk_cnt_en(hssi_10g_rx_pcs_clr_errblk_cnt_en),
				.control_del(hssi_10g_rx_pcs_control_del),
				.crcchk_bypass(hssi_10g_rx_pcs_crcchk_bypass),
				.crcchk_clken(hssi_10g_rx_pcs_crcchk_clken),
				.crcchk_inv(hssi_10g_rx_pcs_crcchk_inv),
				.crcchk_pipeln(hssi_10g_rx_pcs_crcchk_pipeln),
				.crcflag_pipeln(hssi_10g_rx_pcs_crcflag_pipeln),
				.ctrl_bit_reverse(hssi_10g_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_10g_rx_pcs_data_bit_reverse),
				.dec64b66b_clken(hssi_10g_rx_pcs_dec64b66b_clken),
				.dec_64b66b_rxsm_bypass(hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass),
				.descrm_bypass(hssi_10g_rx_pcs_descrm_bypass),
				.descrm_clken(hssi_10g_rx_pcs_descrm_clken),
				.descrm_mode(hssi_10g_rx_pcs_descrm_mode),
				.descrm_pipeln(hssi_10g_rx_pcs_descrm_pipeln),
				.dft_clk_out_sel(hssi_10g_rx_pcs_dft_clk_out_sel),
				.dis_signal_ok(hssi_10g_rx_pcs_dis_signal_ok),
				.dispchk_bypass(hssi_10g_rx_pcs_dispchk_bypass),
				.empty_flag_type(hssi_10g_rx_pcs_empty_flag_type),
				.fast_path(hssi_10g_rx_pcs_fast_path),
				.fec_clken(hssi_10g_rx_pcs_fec_clken),
				.fec_enable(hssi_10g_rx_pcs_fec_enable),
				.fifo_double_read(hssi_10g_rx_pcs_fifo_double_read),
				.fifo_stop_rd(hssi_10g_rx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_rx_pcs_fifo_stop_wr),
				.force_align(hssi_10g_rx_pcs_force_align),
				.frmsync_bypass(hssi_10g_rx_pcs_frmsync_bypass),
				.frmsync_clken(hssi_10g_rx_pcs_frmsync_clken),
				.frmsync_enum_scrm(hssi_10g_rx_pcs_frmsync_enum_scrm),
				.frmsync_enum_sync(hssi_10g_rx_pcs_frmsync_enum_sync),
				.frmsync_flag_type(hssi_10g_rx_pcs_frmsync_flag_type),
				.frmsync_knum_sync(hssi_10g_rx_pcs_frmsync_knum_sync),
				.frmsync_mfrm_length(hssi_10g_rx_pcs_frmsync_mfrm_length),
				.frmsync_pipeln(hssi_10g_rx_pcs_frmsync_pipeln),
				.full_flag_type(hssi_10g_rx_pcs_full_flag_type),
				.gb_rx_idwidth(hssi_10g_rx_pcs_gb_rx_idwidth),
				.gb_rx_odwidth(hssi_10g_rx_pcs_gb_rx_odwidth),
				.gbexp_clken(hssi_10g_rx_pcs_gbexp_clken),
				.low_latency_en(hssi_10g_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_10g_rx_pcs_lpbk_mode),
				.master_clk_sel(hssi_10g_rx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_rx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_rx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_rx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_rx_pcs_pld_if_type),
				.prot_mode(hssi_10g_rx_pcs_prot_mode),
				.rand_clken(hssi_10g_rx_pcs_rand_clken),
				.rd_clk_sel(hssi_10g_rx_pcs_rd_clk_sel),
				.rdfifo_clken(hssi_10g_rx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_rx_pcs_reconfig_settings),
				.rx_fifo_write_ctrl(hssi_10g_rx_pcs_rx_fifo_write_ctrl),
				.rx_scrm_width(hssi_10g_rx_pcs_rx_scrm_width),
				.rx_sh_location(hssi_10g_rx_pcs_rx_sh_location),
				.rx_signal_ok_sel(hssi_10g_rx_pcs_rx_signal_ok_sel),
				.rx_sm_bypass(hssi_10g_rx_pcs_rx_sm_bypass),
				.rx_sm_hiber(hssi_10g_rx_pcs_rx_sm_hiber),
				.rx_sm_pipeln(hssi_10g_rx_pcs_rx_sm_pipeln),
				.rx_testbus_sel(hssi_10g_rx_pcs_rx_testbus_sel),
				.rx_true_b2b(hssi_10g_rx_pcs_rx_true_b2b),
				.rxfifo_empty(hssi_10g_rx_pcs_rxfifo_empty),
				.rxfifo_full(hssi_10g_rx_pcs_rxfifo_full),
				.rxfifo_mode(hssi_10g_rx_pcs_rxfifo_mode),
				.rxfifo_pempty(hssi_10g_rx_pcs_rxfifo_pempty),
				.rxfifo_pfull(hssi_10g_rx_pcs_rxfifo_pfull),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.stretch_num_stages(hssi_10g_rx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_rx_pcs_sup_mode),
				.test_mode(hssi_10g_rx_pcs_test_mode),
				.wrfifo_clken(hssi_10g_rx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_rx_pcs_blockselect),
				.rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.rx_control(w_hssi_10g_rx_pcs_rx_control),
				.rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.rx_data(w_hssi_10g_rx_pcs_rx_data),
				.rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.rx_diag_status(w_hssi_10g_rx_pcs_rx_diag_status),
				.rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.rx_fec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.rx_fifo_num(w_hssi_10g_rx_pcs_rx_fifo_num),
				.rx_fifo_rd_ptr(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr),
				.rx_fifo_rd_ptr2(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2),
				.rx_fifo_wr_clk(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.rx_fifo_wr_data(w_hssi_10g_rx_pcs_rx_fifo_wr_data),
				.rx_fifo_wr_en(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.rx_fifo_wr_ptr(w_hssi_10g_rx_pcs_rx_fifo_wr_ptr),
				.rx_fifo_wr_rst_n(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.rx_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_rx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_rx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.rx_control_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0]}),
				.rx_control_in_krfec({w_hssi_krfec_rx_pcs_rx_control_out[9], w_hssi_krfec_rx_pcs_rx_control_out[8], w_hssi_krfec_rx_pcs_rx_control_out[7], w_hssi_krfec_rx_pcs_rx_control_out[6], w_hssi_krfec_rx_pcs_rx_control_out[5], w_hssi_krfec_rx_pcs_rx_control_out[4], w_hssi_krfec_rx_pcs_rx_control_out[3], w_hssi_krfec_rx_pcs_rx_control_out[2], w_hssi_krfec_rx_pcs_rx_control_out[1], w_hssi_krfec_rx_pcs_rx_control_out[0]}),
				.rx_data_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0]}),
				.rx_data_in_krfec({w_hssi_krfec_rx_pcs_rx_data_out[63], w_hssi_krfec_rx_pcs_rx_data_out[62], w_hssi_krfec_rx_pcs_rx_data_out[61], w_hssi_krfec_rx_pcs_rx_data_out[60], w_hssi_krfec_rx_pcs_rx_data_out[59], w_hssi_krfec_rx_pcs_rx_data_out[58], w_hssi_krfec_rx_pcs_rx_data_out[57], w_hssi_krfec_rx_pcs_rx_data_out[56], w_hssi_krfec_rx_pcs_rx_data_out[55], w_hssi_krfec_rx_pcs_rx_data_out[54], w_hssi_krfec_rx_pcs_rx_data_out[53], w_hssi_krfec_rx_pcs_rx_data_out[52], w_hssi_krfec_rx_pcs_rx_data_out[51], w_hssi_krfec_rx_pcs_rx_data_out[50], w_hssi_krfec_rx_pcs_rx_data_out[49], w_hssi_krfec_rx_pcs_rx_data_out[48], w_hssi_krfec_rx_pcs_rx_data_out[47], w_hssi_krfec_rx_pcs_rx_data_out[46], w_hssi_krfec_rx_pcs_rx_data_out[45], w_hssi_krfec_rx_pcs_rx_data_out[44], w_hssi_krfec_rx_pcs_rx_data_out[43], w_hssi_krfec_rx_pcs_rx_data_out[42], w_hssi_krfec_rx_pcs_rx_data_out[41], w_hssi_krfec_rx_pcs_rx_data_out[40], w_hssi_krfec_rx_pcs_rx_data_out[39], w_hssi_krfec_rx_pcs_rx_data_out[38], w_hssi_krfec_rx_pcs_rx_data_out[37], w_hssi_krfec_rx_pcs_rx_data_out[36], w_hssi_krfec_rx_pcs_rx_data_out[35], w_hssi_krfec_rx_pcs_rx_data_out[34], w_hssi_krfec_rx_pcs_rx_data_out[33], w_hssi_krfec_rx_pcs_rx_data_out[32], w_hssi_krfec_rx_pcs_rx_data_out[31], w_hssi_krfec_rx_pcs_rx_data_out[30], w_hssi_krfec_rx_pcs_rx_data_out[29], w_hssi_krfec_rx_pcs_rx_data_out[28], w_hssi_krfec_rx_pcs_rx_data_out[27], w_hssi_krfec_rx_pcs_rx_data_out[26], w_hssi_krfec_rx_pcs_rx_data_out[25], w_hssi_krfec_rx_pcs_rx_data_out[24], w_hssi_krfec_rx_pcs_rx_data_out[23], w_hssi_krfec_rx_pcs_rx_data_out[22], w_hssi_krfec_rx_pcs_rx_data_out[21], w_hssi_krfec_rx_pcs_rx_data_out[20], w_hssi_krfec_rx_pcs_rx_data_out[19], w_hssi_krfec_rx_pcs_rx_data_out[18], w_hssi_krfec_rx_pcs_rx_data_out[17], w_hssi_krfec_rx_pcs_rx_data_out[16], w_hssi_krfec_rx_pcs_rx_data_out[15], w_hssi_krfec_rx_pcs_rx_data_out[14], w_hssi_krfec_rx_pcs_rx_data_out[13], w_hssi_krfec_rx_pcs_rx_data_out[12], w_hssi_krfec_rx_pcs_rx_data_out[11], w_hssi_krfec_rx_pcs_rx_data_out[10], w_hssi_krfec_rx_pcs_rx_data_out[9], w_hssi_krfec_rx_pcs_rx_data_out[8], w_hssi_krfec_rx_pcs_rx_data_out[7], w_hssi_krfec_rx_pcs_rx_data_out[6], w_hssi_krfec_rx_pcs_rx_data_out[5], w_hssi_krfec_rx_pcs_rx_data_out[4], w_hssi_krfec_rx_pcs_rx_data_out[3], w_hssi_krfec_rx_pcs_rx_data_out[2], w_hssi_krfec_rx_pcs_rx_data_out[1], w_hssi_krfec_rx_pcs_rx_data_out[0]}),
				.rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.rx_data_valid_in_krfec(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_10g[73], w_hssi_fifo_rx_pcs_data_out_10g[72], w_hssi_fifo_rx_pcs_data_out_10g[71], w_hssi_fifo_rx_pcs_data_out_10g[70], w_hssi_fifo_rx_pcs_data_out_10g[69], w_hssi_fifo_rx_pcs_data_out_10g[68], w_hssi_fifo_rx_pcs_data_out_10g[67], w_hssi_fifo_rx_pcs_data_out_10g[66], w_hssi_fifo_rx_pcs_data_out_10g[65], w_hssi_fifo_rx_pcs_data_out_10g[64], w_hssi_fifo_rx_pcs_data_out_10g[63], w_hssi_fifo_rx_pcs_data_out_10g[62], w_hssi_fifo_rx_pcs_data_out_10g[61], w_hssi_fifo_rx_pcs_data_out_10g[60], w_hssi_fifo_rx_pcs_data_out_10g[59], w_hssi_fifo_rx_pcs_data_out_10g[58], w_hssi_fifo_rx_pcs_data_out_10g[57], w_hssi_fifo_rx_pcs_data_out_10g[56], w_hssi_fifo_rx_pcs_data_out_10g[55], w_hssi_fifo_rx_pcs_data_out_10g[54], w_hssi_fifo_rx_pcs_data_out_10g[53], w_hssi_fifo_rx_pcs_data_out_10g[52], w_hssi_fifo_rx_pcs_data_out_10g[51], w_hssi_fifo_rx_pcs_data_out_10g[50], w_hssi_fifo_rx_pcs_data_out_10g[49], w_hssi_fifo_rx_pcs_data_out_10g[48], w_hssi_fifo_rx_pcs_data_out_10g[47], w_hssi_fifo_rx_pcs_data_out_10g[46], w_hssi_fifo_rx_pcs_data_out_10g[45], w_hssi_fifo_rx_pcs_data_out_10g[44], w_hssi_fifo_rx_pcs_data_out_10g[43], w_hssi_fifo_rx_pcs_data_out_10g[42], w_hssi_fifo_rx_pcs_data_out_10g[41], w_hssi_fifo_rx_pcs_data_out_10g[40], w_hssi_fifo_rx_pcs_data_out_10g[39], w_hssi_fifo_rx_pcs_data_out_10g[38], w_hssi_fifo_rx_pcs_data_out_10g[37], w_hssi_fifo_rx_pcs_data_out_10g[36], w_hssi_fifo_rx_pcs_data_out_10g[35], w_hssi_fifo_rx_pcs_data_out_10g[34], w_hssi_fifo_rx_pcs_data_out_10g[33], w_hssi_fifo_rx_pcs_data_out_10g[32], w_hssi_fifo_rx_pcs_data_out_10g[31], w_hssi_fifo_rx_pcs_data_out_10g[30], w_hssi_fifo_rx_pcs_data_out_10g[29], w_hssi_fifo_rx_pcs_data_out_10g[28], w_hssi_fifo_rx_pcs_data_out_10g[27], w_hssi_fifo_rx_pcs_data_out_10g[26], w_hssi_fifo_rx_pcs_data_out_10g[25], w_hssi_fifo_rx_pcs_data_out_10g[24], w_hssi_fifo_rx_pcs_data_out_10g[23], w_hssi_fifo_rx_pcs_data_out_10g[22], w_hssi_fifo_rx_pcs_data_out_10g[21], w_hssi_fifo_rx_pcs_data_out_10g[20], w_hssi_fifo_rx_pcs_data_out_10g[19], w_hssi_fifo_rx_pcs_data_out_10g[18], w_hssi_fifo_rx_pcs_data_out_10g[17], w_hssi_fifo_rx_pcs_data_out_10g[16], w_hssi_fifo_rx_pcs_data_out_10g[15], w_hssi_fifo_rx_pcs_data_out_10g[14], w_hssi_fifo_rx_pcs_data_out_10g[13], w_hssi_fifo_rx_pcs_data_out_10g[12], w_hssi_fifo_rx_pcs_data_out_10g[11], w_hssi_fifo_rx_pcs_data_out_10g[10], w_hssi_fifo_rx_pcs_data_out_10g[9], w_hssi_fifo_rx_pcs_data_out_10g[8], w_hssi_fifo_rx_pcs_data_out_10g[7], w_hssi_fifo_rx_pcs_data_out_10g[6], w_hssi_fifo_rx_pcs_data_out_10g[5], w_hssi_fifo_rx_pcs_data_out_10g[4], w_hssi_fifo_rx_pcs_data_out_10g[3], w_hssi_fifo_rx_pcs_data_out_10g[2], w_hssi_fifo_rx_pcs_data_out_10g[1], w_hssi_fifo_rx_pcs_data_out_10g[0]}),
				.rx_fifo_rd_data_dw({w_hssi_fifo_rx_pcs_data_out2_10g[73], w_hssi_fifo_rx_pcs_data_out2_10g[72], w_hssi_fifo_rx_pcs_data_out2_10g[71], w_hssi_fifo_rx_pcs_data_out2_10g[70], w_hssi_fifo_rx_pcs_data_out2_10g[69], w_hssi_fifo_rx_pcs_data_out2_10g[68], w_hssi_fifo_rx_pcs_data_out2_10g[67], w_hssi_fifo_rx_pcs_data_out2_10g[66], w_hssi_fifo_rx_pcs_data_out2_10g[65], w_hssi_fifo_rx_pcs_data_out2_10g[64], w_hssi_fifo_rx_pcs_data_out2_10g[63], w_hssi_fifo_rx_pcs_data_out2_10g[62], w_hssi_fifo_rx_pcs_data_out2_10g[61], w_hssi_fifo_rx_pcs_data_out2_10g[60], w_hssi_fifo_rx_pcs_data_out2_10g[59], w_hssi_fifo_rx_pcs_data_out2_10g[58], w_hssi_fifo_rx_pcs_data_out2_10g[57], w_hssi_fifo_rx_pcs_data_out2_10g[56], w_hssi_fifo_rx_pcs_data_out2_10g[55], w_hssi_fifo_rx_pcs_data_out2_10g[54], w_hssi_fifo_rx_pcs_data_out2_10g[53], w_hssi_fifo_rx_pcs_data_out2_10g[52], w_hssi_fifo_rx_pcs_data_out2_10g[51], w_hssi_fifo_rx_pcs_data_out2_10g[50], w_hssi_fifo_rx_pcs_data_out2_10g[49], w_hssi_fifo_rx_pcs_data_out2_10g[48], w_hssi_fifo_rx_pcs_data_out2_10g[47], w_hssi_fifo_rx_pcs_data_out2_10g[46], w_hssi_fifo_rx_pcs_data_out2_10g[45], w_hssi_fifo_rx_pcs_data_out2_10g[44], w_hssi_fifo_rx_pcs_data_out2_10g[43], w_hssi_fifo_rx_pcs_data_out2_10g[42], w_hssi_fifo_rx_pcs_data_out2_10g[41], w_hssi_fifo_rx_pcs_data_out2_10g[40], w_hssi_fifo_rx_pcs_data_out2_10g[39], w_hssi_fifo_rx_pcs_data_out2_10g[38], w_hssi_fifo_rx_pcs_data_out2_10g[37], w_hssi_fifo_rx_pcs_data_out2_10g[36], w_hssi_fifo_rx_pcs_data_out2_10g[35], w_hssi_fifo_rx_pcs_data_out2_10g[34], w_hssi_fifo_rx_pcs_data_out2_10g[33], w_hssi_fifo_rx_pcs_data_out2_10g[32], w_hssi_fifo_rx_pcs_data_out2_10g[31], w_hssi_fifo_rx_pcs_data_out2_10g[30], w_hssi_fifo_rx_pcs_data_out2_10g[29], w_hssi_fifo_rx_pcs_data_out2_10g[28], w_hssi_fifo_rx_pcs_data_out2_10g[27], w_hssi_fifo_rx_pcs_data_out2_10g[26], w_hssi_fifo_rx_pcs_data_out2_10g[25], w_hssi_fifo_rx_pcs_data_out2_10g[24], w_hssi_fifo_rx_pcs_data_out2_10g[23], w_hssi_fifo_rx_pcs_data_out2_10g[22], w_hssi_fifo_rx_pcs_data_out2_10g[21], w_hssi_fifo_rx_pcs_data_out2_10g[20], w_hssi_fifo_rx_pcs_data_out2_10g[19], w_hssi_fifo_rx_pcs_data_out2_10g[18], w_hssi_fifo_rx_pcs_data_out2_10g[17], w_hssi_fifo_rx_pcs_data_out2_10g[16], w_hssi_fifo_rx_pcs_data_out2_10g[15], w_hssi_fifo_rx_pcs_data_out2_10g[14], w_hssi_fifo_rx_pcs_data_out2_10g[13], w_hssi_fifo_rx_pcs_data_out2_10g[12], w_hssi_fifo_rx_pcs_data_out2_10g[11], w_hssi_fifo_rx_pcs_data_out2_10g[10], w_hssi_fifo_rx_pcs_data_out2_10g[9], w_hssi_fifo_rx_pcs_data_out2_10g[8], w_hssi_fifo_rx_pcs_data_out2_10g[7], w_hssi_fifo_rx_pcs_data_out2_10g[6], w_hssi_fifo_rx_pcs_data_out2_10g[5], w_hssi_fifo_rx_pcs_data_out2_10g[4], w_hssi_fifo_rx_pcs_data_out2_10g[3], w_hssi_fifo_rx_pcs_data_out2_10g[2], w_hssi_fifo_rx_pcs_data_out2_10g[1], w_hssi_fifo_rx_pcs_data_out2_10g[0]}),
				.rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.rx_pma_data({w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0]}),
				.rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.signal_ok_krfec(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_10g_reg(),
				.pld_10g_krfec_rx_blk_lock_10g_txclk_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_txclk_reg(),
				.pld_10g_krfec_rx_frame_10g_reg(),
				.pld_10g_krfec_rx_frame_10g_txclk_reg(),
				.pld_10g_krfec_rx_pld_rst_n_fifo(),
				.pld_10g_krfec_rx_pld_rst_n_reg(),
				.pld_10g_krfec_rx_pld_rst_n_txclk_reg(),
				.pld_10g_rx_align_clr_fifo(),
				.pld_10g_rx_align_clr_reg(),
				.pld_10g_rx_align_clr_txclk_reg(),
				.pld_10g_rx_align_val_fifo(),
				.pld_10g_rx_align_val_reg(),
				.pld_10g_rx_align_val_txclk_reg(),
				.pld_10g_rx_clr_ber_count_reg(),
				.pld_10g_rx_clr_ber_count_txclk_reg(),
				.pld_10g_rx_crc32_err_reg(),
				.pld_10g_rx_crc32_err_txclk_reg(),
				.pld_10g_rx_data_valid_10g_reg(),
				.pld_10g_rx_data_valid_fifo(),
				.pld_10g_rx_data_valid_pcsdirect_reg(),
				.pld_10g_rx_data_valid_txclk_reg(),
				.pld_10g_rx_empty_fifo(),
				.pld_10g_rx_fifo_del_reg(),
				.pld_10g_rx_fifo_del_txclk_reg(),
				.pld_10g_rx_fifo_insert_fifo(),
				.pld_10g_rx_fifo_num_reg(),
				.pld_10g_rx_fifo_num_txclk_reg(),
				.pld_10g_rx_frame_lock_reg(),
				.pld_10g_rx_frame_lock_txclk_reg(),
				.pld_10g_rx_hi_ber_reg(),
				.pld_10g_rx_hi_ber_txclk_reg(),
				.pld_10g_rx_oflw_err_reg(),
				.pld_10g_rx_oflw_err_txclk_reg(),
				.pld_10g_rx_pempty_fifo(),
				.pld_10g_rx_pfull_reg(),
				.pld_10g_rx_pfull_txclk_reg(),
				.pld_10g_rx_rd_en_fifo(),
				.pld_pcs_rx_clk_out_10g_txclk_wire(),
				.pld_pcs_rx_clk_out_10g_wire(),
				.pld_rx_control_10g_reg(),
				.pld_rx_control_10g_txclk_reg(),
				.pld_rx_data_10g_reg(),
				.pld_rx_data_10g_txclk_reg(),
				.pld_rx_prbs_err_10g_txclk_reg(),
				.pld_rx_prbs_err_clr_10g_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_10g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_align_val = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_blk_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_control[19:0] = 20'b0;
				assign w_hssi_10g_rx_pcs_rx_crc32_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_data[127:0] = 128'b0;
				assign w_hssi_10g_rx_pcs_rx_data_valid = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_dft_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_diag_status[1:0] = 2'b0;
				assign w_hssi_10g_rx_pcs_rx_empty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fec_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_del = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_insert = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_data[73:0] = 74'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_frame_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_hi_ber = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_oflw_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pempty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pfull = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_random_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_rx_frame = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_10g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_tx_pcs
			twentynm_hssi_10g_tx_pcs #(
				.advanced_user_mode(hssi_10g_tx_pcs_advanced_user_mode),
				.bitslip_en(hssi_10g_tx_pcs_bitslip_en),
				.bonding_dft_en(hssi_10g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_10g_tx_pcs_bonding_dft_val),
				.comp_cnt(hssi_10g_tx_pcs_comp_cnt),
				.compin_sel(hssi_10g_tx_pcs_compin_sel),
				.crcgen_bypass(hssi_10g_tx_pcs_crcgen_bypass),
				.crcgen_clken(hssi_10g_tx_pcs_crcgen_clken),
				.crcgen_err(hssi_10g_tx_pcs_crcgen_err),
				.crcgen_inv(hssi_10g_tx_pcs_crcgen_inv),
				.ctrl_bit_reverse(hssi_10g_tx_pcs_ctrl_bit_reverse),
				.ctrl_plane_bonding(hssi_10g_tx_pcs_ctrl_plane_bonding),
				.data_bit_reverse(hssi_10g_tx_pcs_data_bit_reverse),
				.dft_clk_out_sel(hssi_10g_tx_pcs_dft_clk_out_sel),
				.dispgen_bypass(hssi_10g_tx_pcs_dispgen_bypass),
				.dispgen_clken(hssi_10g_tx_pcs_dispgen_clken),
				.dispgen_err(hssi_10g_tx_pcs_dispgen_err),
				.dispgen_pipeln(hssi_10g_tx_pcs_dispgen_pipeln),
				.distdwn_bypass_pipeln(hssi_10g_tx_pcs_distdwn_bypass_pipeln),
				.distdwn_master(hssi_10g_tx_pcs_distdwn_master),
				.distup_bypass_pipeln(hssi_10g_tx_pcs_distup_bypass_pipeln),
				.distup_master(hssi_10g_tx_pcs_distup_master),
				.dv_bond(hssi_10g_tx_pcs_dv_bond),
				.empty_flag_type(hssi_10g_tx_pcs_empty_flag_type),
				.enc64b66b_txsm_clken(hssi_10g_tx_pcs_enc64b66b_txsm_clken),
				.enc_64b66b_txsm_bypass(hssi_10g_tx_pcs_enc_64b66b_txsm_bypass),
				.fastpath(hssi_10g_tx_pcs_fastpath),
				.fec_clken(hssi_10g_tx_pcs_fec_clken),
				.fec_enable(hssi_10g_tx_pcs_fec_enable),
				.fifo_double_write(hssi_10g_tx_pcs_fifo_double_write),
				.fifo_reg_fast(hssi_10g_tx_pcs_fifo_reg_fast),
				.fifo_stop_rd(hssi_10g_tx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_tx_pcs_fifo_stop_wr),
				.frmgen_burst(hssi_10g_tx_pcs_frmgen_burst),
				.frmgen_bypass(hssi_10g_tx_pcs_frmgen_bypass),
				.frmgen_clken(hssi_10g_tx_pcs_frmgen_clken),
				.frmgen_mfrm_length(hssi_10g_tx_pcs_frmgen_mfrm_length),
				.frmgen_pipeln(hssi_10g_tx_pcs_frmgen_pipeln),
				.frmgen_pyld_ins(hssi_10g_tx_pcs_frmgen_pyld_ins),
				.frmgen_wordslip(hssi_10g_tx_pcs_frmgen_wordslip),
				.full_flag_type(hssi_10g_tx_pcs_full_flag_type),
				.gb_pipeln_bypass(hssi_10g_tx_pcs_gb_pipeln_bypass),
				.gb_tx_idwidth(hssi_10g_tx_pcs_gb_tx_idwidth),
				.gb_tx_odwidth(hssi_10g_tx_pcs_gb_tx_odwidth),
				.gbred_clken(hssi_10g_tx_pcs_gbred_clken),
				.indv(hssi_10g_tx_pcs_indv),
				.low_latency_en(hssi_10g_tx_pcs_low_latency_en),
				.master_clk_sel(hssi_10g_tx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_tx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_tx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_tx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_tx_pcs_pld_if_type),
				.prot_mode(hssi_10g_tx_pcs_prot_mode),
				.pseudo_random(hssi_10g_tx_pcs_pseudo_random),
				.pseudo_seed_a(hssi_10g_tx_pcs_pseudo_seed_a),
				.pseudo_seed_b(hssi_10g_tx_pcs_pseudo_seed_b),
				.random_disp(hssi_10g_tx_pcs_random_disp),
				.rdfifo_clken(hssi_10g_tx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_tx_pcs_reconfig_settings),
				.scrm_bypass(hssi_10g_tx_pcs_scrm_bypass),
				.scrm_clken(hssi_10g_tx_pcs_scrm_clken),
				.scrm_mode(hssi_10g_tx_pcs_scrm_mode),
				.scrm_pipeln(hssi_10g_tx_pcs_scrm_pipeln),
				.sh_err(hssi_10g_tx_pcs_sh_err),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sop_mark(hssi_10g_tx_pcs_sop_mark),
				.stretch_num_stages(hssi_10g_tx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_tx_pcs_sup_mode),
				.test_mode(hssi_10g_tx_pcs_test_mode),
				.tx_scrm_err(hssi_10g_tx_pcs_tx_scrm_err),
				.tx_scrm_width(hssi_10g_tx_pcs_tx_scrm_width),
				.tx_sh_location(hssi_10g_tx_pcs_tx_sh_location),
				.tx_sm_bypass(hssi_10g_tx_pcs_tx_sm_bypass),
				.tx_sm_pipeln(hssi_10g_tx_pcs_tx_sm_pipeln),
				.tx_testbus_sel(hssi_10g_tx_pcs_tx_testbus_sel),
				.txfifo_empty(hssi_10g_tx_pcs_txfifo_empty),
				.txfifo_full(hssi_10g_tx_pcs_txfifo_full),
				.txfifo_mode(hssi_10g_tx_pcs_txfifo_mode),
				.txfifo_pempty(hssi_10g_tx_pcs_txfifo_pempty),
				.txfifo_pfull(hssi_10g_tx_pcs_txfifo_pfull),
				.wr_clk_sel(hssi_10g_tx_pcs_wr_clk_sel),
				.wrfifo_clken(hssi_10g_tx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_tx_pcs_blockselect),
				.distdwn_out_dv(w_hssi_10g_tx_pcs_distdwn_out_dv),
				.distdwn_out_rden(w_hssi_10g_tx_pcs_distdwn_out_rden),
				.distdwn_out_wren(w_hssi_10g_tx_pcs_distdwn_out_wren),
				.distup_out_dv(w_hssi_10g_tx_pcs_distup_out_dv),
				.distup_out_rden(w_hssi_10g_tx_pcs_distup_out_rden),
				.distup_out_wren(w_hssi_10g_tx_pcs_distup_out_wren),
				.tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pma_if(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.tx_control_out_krfec(w_hssi_10g_tx_pcs_tx_control_out_krfec),
				.tx_data_out_krfec(w_hssi_10g_tx_pcs_tx_data_out_krfec),
				.tx_data_valid_out_krfec(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.tx_fec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_fifo_num(w_hssi_10g_tx_pcs_tx_fifo_num),
				.tx_fifo_rd_ptr(w_hssi_10g_tx_pcs_tx_fifo_rd_ptr),
				.tx_fifo_wr_clk(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.tx_fifo_wr_data(w_hssi_10g_tx_pcs_tx_fifo_wr_data),
				.tx_fifo_wr_data_dw(w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw),
				.tx_fifo_wr_en(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.tx_fifo_wr_ptr(w_hssi_10g_tx_pcs_tx_fifo_wr_ptr),
				.tx_fifo_wr_rst_n(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.tx_full(w_hssi_10g_tx_pcs_tx_full),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				.tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.tx_pma_data(w_hssi_10g_tx_pcs_tx_pma_data),
				.tx_pma_gating_val(w_hssi_10g_tx_pcs_tx_pma_gating_val),
				.tx_test_data(w_hssi_10g_tx_pcs_tx_test_data),
				.tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.distdwn_in_dv(in_bond_pcs10g_in_bot[2]),
				.distdwn_in_rden(in_bond_pcs10g_in_bot[4]),
				.distdwn_in_wren(in_bond_pcs10g_in_bot[3]),
				.distup_in_dv(in_bond_pcs10g_in_top[2]),
				.distup_in_rden(in_bond_pcs10g_in_top[4]),
				.distup_in_wren(in_bond_pcs10g_in_top[3]),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_tx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_tx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.tx_bitslip({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0]}),
				.tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.tx_control({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0]}),
				.tx_control_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0]}),
				.tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0]}),
				.tx_data_in_krfec({w_hssi_krfec_tx_pcs_tx_data_out[63], w_hssi_krfec_tx_pcs_tx_data_out[62], w_hssi_krfec_tx_pcs_tx_data_out[61], w_hssi_krfec_tx_pcs_tx_data_out[60], w_hssi_krfec_tx_pcs_tx_data_out[59], w_hssi_krfec_tx_pcs_tx_data_out[58], w_hssi_krfec_tx_pcs_tx_data_out[57], w_hssi_krfec_tx_pcs_tx_data_out[56], w_hssi_krfec_tx_pcs_tx_data_out[55], w_hssi_krfec_tx_pcs_tx_data_out[54], w_hssi_krfec_tx_pcs_tx_data_out[53], w_hssi_krfec_tx_pcs_tx_data_out[52], w_hssi_krfec_tx_pcs_tx_data_out[51], w_hssi_krfec_tx_pcs_tx_data_out[50], w_hssi_krfec_tx_pcs_tx_data_out[49], w_hssi_krfec_tx_pcs_tx_data_out[48], w_hssi_krfec_tx_pcs_tx_data_out[47], w_hssi_krfec_tx_pcs_tx_data_out[46], w_hssi_krfec_tx_pcs_tx_data_out[45], w_hssi_krfec_tx_pcs_tx_data_out[44], w_hssi_krfec_tx_pcs_tx_data_out[43], w_hssi_krfec_tx_pcs_tx_data_out[42], w_hssi_krfec_tx_pcs_tx_data_out[41], w_hssi_krfec_tx_pcs_tx_data_out[40], w_hssi_krfec_tx_pcs_tx_data_out[39], w_hssi_krfec_tx_pcs_tx_data_out[38], w_hssi_krfec_tx_pcs_tx_data_out[37], w_hssi_krfec_tx_pcs_tx_data_out[36], w_hssi_krfec_tx_pcs_tx_data_out[35], w_hssi_krfec_tx_pcs_tx_data_out[34], w_hssi_krfec_tx_pcs_tx_data_out[33], w_hssi_krfec_tx_pcs_tx_data_out[32], w_hssi_krfec_tx_pcs_tx_data_out[31], w_hssi_krfec_tx_pcs_tx_data_out[30], w_hssi_krfec_tx_pcs_tx_data_out[29], w_hssi_krfec_tx_pcs_tx_data_out[28], w_hssi_krfec_tx_pcs_tx_data_out[27], w_hssi_krfec_tx_pcs_tx_data_out[26], w_hssi_krfec_tx_pcs_tx_data_out[25], w_hssi_krfec_tx_pcs_tx_data_out[24], w_hssi_krfec_tx_pcs_tx_data_out[23], w_hssi_krfec_tx_pcs_tx_data_out[22], w_hssi_krfec_tx_pcs_tx_data_out[21], w_hssi_krfec_tx_pcs_tx_data_out[20], w_hssi_krfec_tx_pcs_tx_data_out[19], w_hssi_krfec_tx_pcs_tx_data_out[18], w_hssi_krfec_tx_pcs_tx_data_out[17], w_hssi_krfec_tx_pcs_tx_data_out[16], w_hssi_krfec_tx_pcs_tx_data_out[15], w_hssi_krfec_tx_pcs_tx_data_out[14], w_hssi_krfec_tx_pcs_tx_data_out[13], w_hssi_krfec_tx_pcs_tx_data_out[12], w_hssi_krfec_tx_pcs_tx_data_out[11], w_hssi_krfec_tx_pcs_tx_data_out[10], w_hssi_krfec_tx_pcs_tx_data_out[9], w_hssi_krfec_tx_pcs_tx_data_out[8], w_hssi_krfec_tx_pcs_tx_data_out[7], w_hssi_krfec_tx_pcs_tx_data_out[6], w_hssi_krfec_tx_pcs_tx_data_out[5], w_hssi_krfec_tx_pcs_tx_data_out[4], w_hssi_krfec_tx_pcs_tx_data_out[3], w_hssi_krfec_tx_pcs_tx_data_out[2], w_hssi_krfec_tx_pcs_tx_data_out[1], w_hssi_krfec_tx_pcs_tx_data_out[0]}),
				.tx_data_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0]}),
				.tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.tx_diag_status({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0]}),
				.tx_fifo_rd_data({w_hssi_fifo_tx_pcs_data_out_10g[72], w_hssi_fifo_tx_pcs_data_out_10g[71], w_hssi_fifo_tx_pcs_data_out_10g[70], w_hssi_fifo_tx_pcs_data_out_10g[69], w_hssi_fifo_tx_pcs_data_out_10g[68], w_hssi_fifo_tx_pcs_data_out_10g[67], w_hssi_fifo_tx_pcs_data_out_10g[66], w_hssi_fifo_tx_pcs_data_out_10g[65], w_hssi_fifo_tx_pcs_data_out_10g[64], w_hssi_fifo_tx_pcs_data_out_10g[63], w_hssi_fifo_tx_pcs_data_out_10g[62], w_hssi_fifo_tx_pcs_data_out_10g[61], w_hssi_fifo_tx_pcs_data_out_10g[60], w_hssi_fifo_tx_pcs_data_out_10g[59], w_hssi_fifo_tx_pcs_data_out_10g[58], w_hssi_fifo_tx_pcs_data_out_10g[57], w_hssi_fifo_tx_pcs_data_out_10g[56], w_hssi_fifo_tx_pcs_data_out_10g[55], w_hssi_fifo_tx_pcs_data_out_10g[54], w_hssi_fifo_tx_pcs_data_out_10g[53], w_hssi_fifo_tx_pcs_data_out_10g[52], w_hssi_fifo_tx_pcs_data_out_10g[51], w_hssi_fifo_tx_pcs_data_out_10g[50], w_hssi_fifo_tx_pcs_data_out_10g[49], w_hssi_fifo_tx_pcs_data_out_10g[48], w_hssi_fifo_tx_pcs_data_out_10g[47], w_hssi_fifo_tx_pcs_data_out_10g[46], w_hssi_fifo_tx_pcs_data_out_10g[45], w_hssi_fifo_tx_pcs_data_out_10g[44], w_hssi_fifo_tx_pcs_data_out_10g[43], w_hssi_fifo_tx_pcs_data_out_10g[42], w_hssi_fifo_tx_pcs_data_out_10g[41], w_hssi_fifo_tx_pcs_data_out_10g[40], w_hssi_fifo_tx_pcs_data_out_10g[39], w_hssi_fifo_tx_pcs_data_out_10g[38], w_hssi_fifo_tx_pcs_data_out_10g[37], w_hssi_fifo_tx_pcs_data_out_10g[36], w_hssi_fifo_tx_pcs_data_out_10g[35], w_hssi_fifo_tx_pcs_data_out_10g[34], w_hssi_fifo_tx_pcs_data_out_10g[33], w_hssi_fifo_tx_pcs_data_out_10g[32], w_hssi_fifo_tx_pcs_data_out_10g[31], w_hssi_fifo_tx_pcs_data_out_10g[30], w_hssi_fifo_tx_pcs_data_out_10g[29], w_hssi_fifo_tx_pcs_data_out_10g[28], w_hssi_fifo_tx_pcs_data_out_10g[27], w_hssi_fifo_tx_pcs_data_out_10g[26], w_hssi_fifo_tx_pcs_data_out_10g[25], w_hssi_fifo_tx_pcs_data_out_10g[24], w_hssi_fifo_tx_pcs_data_out_10g[23], w_hssi_fifo_tx_pcs_data_out_10g[22], w_hssi_fifo_tx_pcs_data_out_10g[21], w_hssi_fifo_tx_pcs_data_out_10g[20], w_hssi_fifo_tx_pcs_data_out_10g[19], w_hssi_fifo_tx_pcs_data_out_10g[18], w_hssi_fifo_tx_pcs_data_out_10g[17], w_hssi_fifo_tx_pcs_data_out_10g[16], w_hssi_fifo_tx_pcs_data_out_10g[15], w_hssi_fifo_tx_pcs_data_out_10g[14], w_hssi_fifo_tx_pcs_data_out_10g[13], w_hssi_fifo_tx_pcs_data_out_10g[12], w_hssi_fifo_tx_pcs_data_out_10g[11], w_hssi_fifo_tx_pcs_data_out_10g[10], w_hssi_fifo_tx_pcs_data_out_10g[9], w_hssi_fifo_tx_pcs_data_out_10g[8], w_hssi_fifo_tx_pcs_data_out_10g[7], w_hssi_fifo_tx_pcs_data_out_10g[6], w_hssi_fifo_tx_pcs_data_out_10g[5], w_hssi_fifo_tx_pcs_data_out_10g[4], w_hssi_fifo_tx_pcs_data_out_10g[3], w_hssi_fifo_tx_pcs_data_out_10g[2], w_hssi_fifo_tx_pcs_data_out_10g[1], w_hssi_fifo_tx_pcs_data_out_10g[0]}),
				.tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_10g_reg(),
				.pld_10g_krfec_tx_pld_rst_n_fifo(),
				.pld_10g_krfec_tx_pld_rst_n_reg(),
				.pld_10g_tx_bitslip_reg(),
				.pld_10g_tx_burst_en_exe_reg(),
				.pld_10g_tx_data_valid_10g_reg(),
				.pld_10g_tx_data_valid_fifo(),
				.pld_10g_tx_data_valid_reg(),
				.pld_10g_tx_diag_status_reg(),
				.pld_10g_tx_empty_reg(),
				.pld_10g_tx_fifo_num_reg(),
				.pld_10g_tx_full_fifo(),
				.pld_10g_tx_full_reg(),
				.pld_10g_tx_pempty_reg(),
				.pld_10g_tx_pfull_fifo(),
				.pld_10g_tx_wordslip_exe_reg(),
				.pld_10g_tx_wordslip_reg(),
				.pld_pcs_tx_clk_out_10g_wire(),
				.pld_tx_burst_en_reg(),
				.pld_tx_control_lo_10g_reg(),
				.pld_tx_data_10g_fifo(),
				.pld_tx_data_lo_10g_reg()
			);
		end // if generate
		else begin
				assign w_hssi_10g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_burst_en_exe = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pma_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_control_out_krfec[8:0] = 9'b0;
				assign w_hssi_10g_tx_pcs_tx_data_out_krfec[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_data_valid_out_krfec = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_dft_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_empty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fec_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_full = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_pempty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pfull = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_gating_val[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_test_data[19:0] = 20'b0;
				assign w_hssi_10g_tx_pcs_tx_wordslip_exe = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_rx_pcs
			twentynm_hssi_8g_rx_pcs #(
				.auto_error_replacement(hssi_8g_rx_pcs_auto_error_replacement),
				.auto_speed_nego(hssi_8g_rx_pcs_auto_speed_nego),
				.bit_reversal(hssi_8g_rx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_rx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_rx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_rx_pcs_bypass_pipeline_reg),
				.byte_deserializer(hssi_8g_rx_pcs_byte_deserializer),
				.cdr_ctrl_rxvalid_mask(hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask),
				.clkcmp_pattern_n(hssi_8g_rx_pcs_clkcmp_pattern_n),
				.clkcmp_pattern_p(hssi_8g_rx_pcs_clkcmp_pattern_p),
				.clock_gate_bds_dec_asn(hssi_8g_rx_pcs_clock_gate_bds_dec_asn),
				.clock_gate_cdr_eidle(hssi_8g_rx_pcs_clock_gate_cdr_eidle),
				.clock_gate_dw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk),
				.clock_gate_dw_rm_rd(hssi_8g_rx_pcs_clock_gate_dw_rm_rd),
				.clock_gate_dw_rm_wr(hssi_8g_rx_pcs_clock_gate_dw_rm_wr),
				.clock_gate_dw_wa(hssi_8g_rx_pcs_clock_gate_dw_wa),
				.clock_gate_pc_rdclk(hssi_8g_rx_pcs_clock_gate_pc_rdclk),
				.clock_gate_sw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk),
				.clock_gate_sw_rm_rd(hssi_8g_rx_pcs_clock_gate_sw_rm_rd),
				.clock_gate_sw_rm_wr(hssi_8g_rx_pcs_clock_gate_sw_rm_wr),
				.clock_gate_sw_wa(hssi_8g_rx_pcs_clock_gate_sw_wa),
				.clock_observation_in_pld_core(hssi_8g_rx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_rx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_rx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_rx_pcs_ctrl_plane_bonding_distribution),
				.eidle_entry_eios(hssi_8g_rx_pcs_eidle_entry_eios),
				.eidle_entry_iei(hssi_8g_rx_pcs_eidle_entry_iei),
				.eidle_entry_sd(hssi_8g_rx_pcs_eidle_entry_sd),
				.eightb_tenb_decoder(hssi_8g_rx_pcs_eightb_tenb_decoder),
				.err_flags_sel(hssi_8g_rx_pcs_err_flags_sel),
				.fixed_pat_det(hssi_8g_rx_pcs_fixed_pat_det),
				.fixed_pat_num(hssi_8g_rx_pcs_fixed_pat_num),
				.force_signal_detect(hssi_8g_rx_pcs_force_signal_detect),
				.gen3_clk_en(hssi_8g_rx_pcs_gen3_clk_en),
				.gen3_rx_clk_sel(hssi_8g_rx_pcs_gen3_rx_clk_sel),
				.gen3_tx_clk_sel(hssi_8g_rx_pcs_gen3_tx_clk_sel),
				.hip_mode(hssi_8g_rx_pcs_hip_mode),
				.ibm_invalid_code(hssi_8g_rx_pcs_ibm_invalid_code),
				.invalid_code_flag_only(hssi_8g_rx_pcs_invalid_code_flag_only),
				.pad_or_edb_error_replace(hssi_8g_rx_pcs_pad_or_edb_error_replace),
				.pcs_bypass(hssi_8g_rx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_rx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_rx_pcs_phase_compensation_fifo),
				.pipe_if_enable(hssi_8g_rx_pcs_pipe_if_enable),
				.pma_dw(hssi_8g_rx_pcs_pma_dw),
				.polinv_8b10b_dec(hssi_8g_rx_pcs_polinv_8b10b_dec),
				.prot_mode(hssi_8g_rx_pcs_prot_mode),
				.rate_match(hssi_8g_rx_pcs_rate_match),
				.rate_match_del_thres(hssi_8g_rx_pcs_rate_match_del_thres),
				.rate_match_empty_thres(hssi_8g_rx_pcs_rate_match_empty_thres),
				.rate_match_full_thres(hssi_8g_rx_pcs_rate_match_full_thres),
				.rate_match_ins_thres(hssi_8g_rx_pcs_rate_match_ins_thres),
				.rate_match_start_thres(hssi_8g_rx_pcs_rate_match_start_thres),
				.reconfig_settings(hssi_8g_rx_pcs_reconfig_settings),
				.rx_clk2(hssi_8g_rx_pcs_rx_clk2),
				.rx_clk_free_running(hssi_8g_rx_pcs_rx_clk_free_running),
				.rx_pcs_urst(hssi_8g_rx_pcs_rx_pcs_urst),
				.rx_rcvd_clk(hssi_8g_rx_pcs_rx_rcvd_clk),
				.rx_rd_clk(hssi_8g_rx_pcs_rx_rd_clk),
				.rx_refclk(hssi_8g_rx_pcs_rx_refclk),
				.rx_wr_clk(hssi_8g_rx_pcs_rx_wr_clk),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_rx_pcs_sup_mode),
				.symbol_swap(hssi_8g_rx_pcs_symbol_swap),
				.sync_sm_idle_eios(hssi_8g_rx_pcs_sync_sm_idle_eios),
				.test_bus_sel(hssi_8g_rx_pcs_test_bus_sel),
				.tx_rx_parallel_loopback(hssi_8g_rx_pcs_tx_rx_parallel_loopback),
				.wa_boundary_lock_ctrl(hssi_8g_rx_pcs_wa_boundary_lock_ctrl),
				.wa_clk_slip_spacing(hssi_8g_rx_pcs_wa_clk_slip_spacing),
				.wa_det_latency_sync_status_beh(hssi_8g_rx_pcs_wa_det_latency_sync_status_beh),
				.wa_disp_err_flag(hssi_8g_rx_pcs_wa_disp_err_flag),
				.wa_kchar(hssi_8g_rx_pcs_wa_kchar),
				.wa_pd(hssi_8g_rx_pcs_wa_pd),
				.wa_pd_data(hssi_8g_rx_pcs_wa_pd_data),
				.wa_pd_polarity(hssi_8g_rx_pcs_wa_pd_polarity),
				.wa_pld_controlled(hssi_8g_rx_pcs_wa_pld_controlled),
				.wa_renumber_data(hssi_8g_rx_pcs_wa_renumber_data),
				.wa_rgnumber_data(hssi_8g_rx_pcs_wa_rgnumber_data),
				.wa_rknumber_data(hssi_8g_rx_pcs_wa_rknumber_data),
				.wa_rosnumber_data(hssi_8g_rx_pcs_wa_rosnumber_data),
				.wa_rvnumber_data(hssi_8g_rx_pcs_wa_rvnumber_data),
				.wa_sync_sm_ctrl(hssi_8g_rx_pcs_wa_sync_sm_ctrl),
				.wait_cnt(hssi_8g_rx_pcs_wait_cnt)
			) inst_twentynm_hssi_8g_rx_pcs (
				// OUTPUTS
				.a1a2k1k2flag(w_hssi_8g_rx_pcs_a1a2k1k2flag),
				.avmmreaddata(w_hssi_8g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_rx_pcs_blockselect),
				.chnl_test_bus_out(w_hssi_8g_rx_pcs_chnl_test_bus_out),
				.clock_to_pld(w_hssi_8g_rx_pcs_clock_to_pld),
				.dataout(w_hssi_8g_rx_pcs_dataout),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidle_detected(w_hssi_8g_rx_pcs_eidle_detected),
				.eios_det_cdr_ctrl(w_hssi_8g_rx_pcs_eios_det_cdr_ctrl),
				.g3_rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.g3_rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.gen2ngen1(w_hssi_8g_rx_pcs_gen2ngen1),
				.parallel_rev_loopback(w_hssi_8g_rx_pcs_parallel_rev_loopback),
				.pc_fifo_empty(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.pcfifofull(w_hssi_8g_rx_pcs_pcfifofull),
				.phystatus(w_hssi_8g_rx_pcs_phystatus),
				.pipe_data(w_hssi_8g_rx_pcs_pipe_data),
				.rd_enable_out_chnl_down(w_hssi_8g_rx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_rx_pcs_rd_enable_out_chnl_up),
				.rd_ptr1_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo),
				.rd_ptr2_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo),
				.rd_ptr_rx_phfifo(w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.reset_pc_ptrs_out_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down),
				.reset_pc_ptrs_out_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up),
				.rm_fifo_empty(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.rm_fifo_full(w_hssi_8g_rx_pcs_rm_fifo_full),
				.rx_blk_start(w_hssi_8g_rx_pcs_rx_blk_start),
				.rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.rx_data_valid(w_hssi_8g_rx_pcs_rx_data_valid),
				.rx_div_sync_out_chnl_down(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down),
				.rx_div_sync_out_chnl_up(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up),
				.rx_pipe_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.rx_pipe_soft_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rx_pma_clk_gen3(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_rcvd_clk_gen3(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_rstn_sync2wrfifo_8g(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.rx_sync_hdr(w_hssi_8g_rx_pcs_rx_sync_hdr),
				.rx_we_out_chnl_down(w_hssi_8g_rx_pcs_rx_we_out_chnl_down),
				.rx_we_out_chnl_up(w_hssi_8g_rx_pcs_rx_we_out_chnl_up),
				.rxstatus(w_hssi_8g_rx_pcs_rxstatus),
				.rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.word_align_boundary(w_hssi_8g_rx_pcs_word_align_boundary),
				.wr_clk_rx_phfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_rx_phfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_rx_rmfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_rx_rmfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_data_rx_phfifo(w_hssi_8g_rx_pcs_wr_data_rx_phfifo),
				.wr_data_rx_rmfifo(w_hssi_8g_rx_pcs_wr_data_rx_rmfifo),
				.wr_en_rx_phfifo(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_rx_rmfifo(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_rx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_rx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_rx_phfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo),
				.wr_ptr_rx_rmfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo),
				.wr_rst_n_rx_phfifo(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_rx_rmfifo(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				// INPUTS
				.a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bit_reversal_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.datain({w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0]}),
				.disable_pc_fifo_byte_serdes(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4]),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.eidleinfersel({w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0]}),
				.eios_detected_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.enable_comma_detect(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.gen3_clk_sel(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.hrd_rst(1'b0),
				.inferred_rxvalid_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.pc_fifo_rd_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.pc_fifo_wrdisable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.phystatus_int(w_hssi_pipe_gen1_2_phystatus),
				.phystatus_pcs_gen3(w_hssi_pipe_gen3_phystatus),
				.pipe_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.polarity_inversion(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.rd_data1_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0]}),
				.rd_data2_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0]}),
				.rd_data_rx_phfifo({w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[3]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[3]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.reset_pc_ptrs_asn(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5]),
				.reset_pc_ptrs_in_chnl_down(in_bond_pcs8g_in_bot[12]),
				.reset_pc_ptrs_in_chnl_up(in_bond_pcs8g_in_top[12]),
				.reset_ppm_cntrs_pcs_pma(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7]),
				.rm_fifo_read_enable(1'b0),
				.rm_fifo_write_enable(1'b0),
				.rx_blk_start_pcs_gen3({w_hssi_pipe_gen3_rx_blk_start[3], w_hssi_pipe_gen3_rx_blk_start[2], w_hssi_pipe_gen3_rx_blk_start[1], w_hssi_pipe_gen3_rx_blk_start[0]}),
				.rx_data_pcs_gen3({w_hssi_pipe_gen3_rxd_8gpcs_out[63], w_hssi_pipe_gen3_rxd_8gpcs_out[62], w_hssi_pipe_gen3_rxd_8gpcs_out[61], w_hssi_pipe_gen3_rxd_8gpcs_out[60], w_hssi_pipe_gen3_rxd_8gpcs_out[59], w_hssi_pipe_gen3_rxd_8gpcs_out[58], w_hssi_pipe_gen3_rxd_8gpcs_out[57], w_hssi_pipe_gen3_rxd_8gpcs_out[56], w_hssi_pipe_gen3_rxd_8gpcs_out[55], w_hssi_pipe_gen3_rxd_8gpcs_out[54], w_hssi_pipe_gen3_rxd_8gpcs_out[53], w_hssi_pipe_gen3_rxd_8gpcs_out[52], w_hssi_pipe_gen3_rxd_8gpcs_out[51], w_hssi_pipe_gen3_rxd_8gpcs_out[50], w_hssi_pipe_gen3_rxd_8gpcs_out[49], w_hssi_pipe_gen3_rxd_8gpcs_out[48], w_hssi_pipe_gen3_rxd_8gpcs_out[47], w_hssi_pipe_gen3_rxd_8gpcs_out[46], w_hssi_pipe_gen3_rxd_8gpcs_out[45], w_hssi_pipe_gen3_rxd_8gpcs_out[44], w_hssi_pipe_gen3_rxd_8gpcs_out[43], w_hssi_pipe_gen3_rxd_8gpcs_out[42], w_hssi_pipe_gen3_rxd_8gpcs_out[41], w_hssi_pipe_gen3_rxd_8gpcs_out[40], w_hssi_pipe_gen3_rxd_8gpcs_out[39], w_hssi_pipe_gen3_rxd_8gpcs_out[38], w_hssi_pipe_gen3_rxd_8gpcs_out[37], w_hssi_pipe_gen3_rxd_8gpcs_out[36], w_hssi_pipe_gen3_rxd_8gpcs_out[35], w_hssi_pipe_gen3_rxd_8gpcs_out[34], w_hssi_pipe_gen3_rxd_8gpcs_out[33], w_hssi_pipe_gen3_rxd_8gpcs_out[32], w_hssi_pipe_gen3_rxd_8gpcs_out[31], w_hssi_pipe_gen3_rxd_8gpcs_out[30], w_hssi_pipe_gen3_rxd_8gpcs_out[29], w_hssi_pipe_gen3_rxd_8gpcs_out[28], w_hssi_pipe_gen3_rxd_8gpcs_out[27], w_hssi_pipe_gen3_rxd_8gpcs_out[26], w_hssi_pipe_gen3_rxd_8gpcs_out[25], w_hssi_pipe_gen3_rxd_8gpcs_out[24], w_hssi_pipe_gen3_rxd_8gpcs_out[23], w_hssi_pipe_gen3_rxd_8gpcs_out[22], w_hssi_pipe_gen3_rxd_8gpcs_out[21], w_hssi_pipe_gen3_rxd_8gpcs_out[20], w_hssi_pipe_gen3_rxd_8gpcs_out[19], w_hssi_pipe_gen3_rxd_8gpcs_out[18], w_hssi_pipe_gen3_rxd_8gpcs_out[17], w_hssi_pipe_gen3_rxd_8gpcs_out[16], w_hssi_pipe_gen3_rxd_8gpcs_out[15], w_hssi_pipe_gen3_rxd_8gpcs_out[14], w_hssi_pipe_gen3_rxd_8gpcs_out[13], w_hssi_pipe_gen3_rxd_8gpcs_out[12], w_hssi_pipe_gen3_rxd_8gpcs_out[11], w_hssi_pipe_gen3_rxd_8gpcs_out[10], w_hssi_pipe_gen3_rxd_8gpcs_out[9], w_hssi_pipe_gen3_rxd_8gpcs_out[8], w_hssi_pipe_gen3_rxd_8gpcs_out[7], w_hssi_pipe_gen3_rxd_8gpcs_out[6], w_hssi_pipe_gen3_rxd_8gpcs_out[5], w_hssi_pipe_gen3_rxd_8gpcs_out[4], w_hssi_pipe_gen3_rxd_8gpcs_out[3], w_hssi_pipe_gen3_rxd_8gpcs_out[2], w_hssi_pipe_gen3_rxd_8gpcs_out[1], w_hssi_pipe_gen3_rxd_8gpcs_out[0]}),
				.rx_data_valid_pcs_gen3({w_hssi_pipe_gen3_rxdataskip[3], w_hssi_pipe_gen3_rxdataskip[2], w_hssi_pipe_gen3_rxdataskip[1], w_hssi_pipe_gen3_rxdataskip[0]}),
				.rx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[1], in_bond_pcs8g_in_bot[0]}),
				.rx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[1], in_bond_pcs8g_in_top[0]}),
				.rx_pcs_rst(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.rx_sync_hdr_pcs_gen3({w_hssi_pipe_gen3_rx_sync_hdr[1], w_hssi_pipe_gen3_rx_sync_hdr[0]}),
				.rx_we_in_chnl_down({in_bond_pcs8g_in_bot[5], in_bond_pcs8g_in_bot[4]}),
				.rx_we_in_chnl_up({in_bond_pcs8g_in_top[5], in_bond_pcs8g_in_top[4]}),
				.rxstatus_int({w_hssi_pipe_gen1_2_rxstatus[2], w_hssi_pipe_gen1_2_rxstatus[1], w_hssi_pipe_gen1_2_rxstatus[0]}),
				.rxstatus_pcs_gen3({w_hssi_pipe_gen3_rxstatus[2], w_hssi_pipe_gen3_rxstatus[1], w_hssi_pipe_gen3_rxstatus[0]}),
				.rxvalid_int(w_hssi_pipe_gen1_2_rxvalid),
				.rxvalid_pcs_gen3(w_hssi_pipe_gen3_rxvalid),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.sig_det_from_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_ctrlplane_testbus({w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0]}),
				.tx_div_sync({w_hssi_8g_tx_pcs_tx_div_sync[1], w_hssi_8g_tx_pcs_tx_div_sync[0]}),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.tx_testbus({w_hssi_8g_tx_pcs_tx_testbus[19], w_hssi_8g_tx_pcs_tx_testbus[18], w_hssi_8g_tx_pcs_tx_testbus[17], w_hssi_8g_tx_pcs_tx_testbus[16], w_hssi_8g_tx_pcs_tx_testbus[15], w_hssi_8g_tx_pcs_tx_testbus[14], w_hssi_8g_tx_pcs_tx_testbus[13], w_hssi_8g_tx_pcs_tx_testbus[12], w_hssi_8g_tx_pcs_tx_testbus[11], w_hssi_8g_tx_pcs_tx_testbus[10], w_hssi_8g_tx_pcs_tx_testbus[9], w_hssi_8g_tx_pcs_tx_testbus[8], w_hssi_8g_tx_pcs_tx_testbus[7], w_hssi_8g_tx_pcs_tx_testbus[6], w_hssi_8g_tx_pcs_tx_testbus[5], w_hssi_8g_tx_pcs_tx_testbus[4], w_hssi_8g_tx_pcs_tx_testbus[3], w_hssi_8g_tx_pcs_tx_testbus[2], w_hssi_8g_tx_pcs_tx_testbus[1], w_hssi_8g_tx_pcs_tx_testbus[0]}),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[2]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[2]),
				
				// UNUSED
				.byte_deserializer_pcs_clk_div_by_2_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_wire(),
				.byte_deserializer_pcs_clk_div_by_2_wire(),
				.byte_deserializer_pcs_clk_div_by_4_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_2_reg(),
				.byte_deserializer_pld_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_4_txclk_reg(),
				.pld_8g_a1a2_k1k2_flag_reg(),
				.pld_8g_a1a2_k1k2_flag_txclk_reg(),
				.pld_8g_a1a2_size_reg(),
				.pld_8g_a1a2_size_txclk_reg(),
				.pld_8g_bitloc_rev_en_reg(),
				.pld_8g_bitloc_rev_en_txclk_reg(),
				.pld_8g_byte_rev_en_reg(),
				.pld_8g_byte_rev_en_txclk_reg(),
				.pld_8g_elecidle_reg(),
				.pld_8g_empty_rmf_lowlatency_reg(),
				.pld_8g_empty_rmf_lowlatency_txclk_reg(),
				.pld_8g_empty_rmf_reg(),
				.pld_8g_empty_rmf_txclk_reg(),
				.pld_8g_empty_rx_fifo(),
				.pld_8g_empty_rx_reg(),
				.pld_8g_empty_rx_txclk_reg(),
				.pld_8g_encdt_reg(),
				.pld_8g_encdt_txclk_reg(),
				.pld_8g_full_rmf_reg(),
				.pld_8g_full_rmf_txclk_reg(),
				.pld_8g_full_rx_fifo(),
				.pld_8g_full_rx_reg(),
				.pld_8g_full_rx_txclk_reg(),
				.pld_8g_g3_rx_pld_rst_n_reg(),
				.pld_8g_g3_rx_pld_rst_n_txclk_reg(),
				.pld_8g_rxelecidle_txclk_reg(),
				.pld_8g_rxpolarity_reg(),
				.pld_8g_rxpolarity_txclk_reg(),
				.pld_8g_wa_boundary_reg(),
				.pld_8g_wrdisable_rx_reg(),
				.pld_8g_wrdisable_rx_txclk_reg(),
				.pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_rx_clk_out_8g_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_wire(),
				.pld_rx_control_8g_reg(),
				.pld_rx_control_8g_txclk_reg(),
				.pld_rx_data_8g_reg(),
				.pld_rx_data_8g_txclk_reg(),
				.pld_syncsm_en_reg(),
				.pld_syncsm_en_txclk_reg(),
				.rm_fifo_partial_empty(),
				.rm_fifo_partial_full(),
				.sta_rx_clk2_by2_1(),
				.sta_rx_clk2_by2_1_out(),
				.sta_rx_clk2_by2_2(),
				.sta_rx_clk2_by2_2_out(),
				.sta_rx_clk2_by4_1(),
				.sta_rx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_rx_pcs_a1a2k1k2flag[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_rx_pcs_chnl_test_bus_out[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_clock_to_pld = 1'b0;
				assign w_hssi_8g_rx_pcs_dataout[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_dis_pc_byte = 1'b0;
				assign w_hssi_8g_rx_pcs_eidle_detected = 1'b0;
				assign w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_pma_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_gen2ngen1 = 1'b0;
				assign w_hssi_8g_rx_pcs_parallel_rev_loopback[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_pc_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_pcfifofull = 1'b0;
				assign w_hssi_8g_rx_pcs_phystatus = 1'b0;
				assign w_hssi_8g_rx_pcs_pipe_data[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_full = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clkslip = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_data_valid[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pma_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rxstatus[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_rxvalid = 1'b0;
				assign w_hssi_8g_rx_pcs_signal_detect_out = 1'b0;
				assign w_hssi_8g_rx_pcs_word_align_boundary[4:0] = 5'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79:0] = 80'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31:0] = 32'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_rmfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_tx_pcs
			twentynm_hssi_8g_tx_pcs #(
				.auto_speed_nego_gen2(hssi_8g_tx_pcs_auto_speed_nego_gen2),
				.bit_reversal(hssi_8g_tx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_tx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_tx_pcs_bypass_pipeline_reg),
				.byte_serializer(hssi_8g_tx_pcs_byte_serializer),
				.clock_gate_bs_enc(hssi_8g_tx_pcs_clock_gate_bs_enc),
				.clock_gate_dw_fifowr(hssi_8g_tx_pcs_clock_gate_dw_fifowr),
				.clock_gate_fiford(hssi_8g_tx_pcs_clock_gate_fiford),
				.clock_gate_sw_fifowr(hssi_8g_tx_pcs_clock_gate_sw_fifowr),
				.clock_observation_in_pld_core(hssi_8g_tx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_tx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_tx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_tx_pcs_ctrl_plane_bonding_distribution),
				.data_selection_8b10b_encoder_input(hssi_8g_tx_pcs_data_selection_8b10b_encoder_input),
				.dynamic_clk_switch(hssi_8g_tx_pcs_dynamic_clk_switch),
				.eightb_tenb_disp_ctrl(hssi_8g_tx_pcs_eightb_tenb_disp_ctrl),
				.eightb_tenb_encoder(hssi_8g_tx_pcs_eightb_tenb_encoder),
				.force_echar(hssi_8g_tx_pcs_force_echar),
				.force_kchar(hssi_8g_tx_pcs_force_kchar),
				.gen3_tx_clk_sel(hssi_8g_tx_pcs_gen3_tx_clk_sel),
				.gen3_tx_pipe_clk_sel(hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel),
				.hip_mode(hssi_8g_tx_pcs_hip_mode),
				.pcs_bypass(hssi_8g_tx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_tx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_tx_pcs_phase_compensation_fifo),
				.phfifo_write_clk_sel(hssi_8g_tx_pcs_phfifo_write_clk_sel),
				.pma_dw(hssi_8g_tx_pcs_pma_dw),
				.prot_mode(hssi_8g_tx_pcs_prot_mode),
				.reconfig_settings(hssi_8g_tx_pcs_reconfig_settings),
				.refclk_b_clk_sel(hssi_8g_tx_pcs_refclk_b_clk_sel),
				.revloop_back_rm(hssi_8g_tx_pcs_revloop_back_rm),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_tx_pcs_sup_mode),
				.symbol_swap(hssi_8g_tx_pcs_symbol_swap),
				.tx_bitslip(hssi_8g_tx_pcs_tx_bitslip),
				.tx_compliance_controlled_disparity(hssi_8g_tx_pcs_tx_compliance_controlled_disparity),
				.tx_fast_pld_reg(hssi_8g_tx_pcs_tx_fast_pld_reg),
				.txclk_freerun(hssi_8g_tx_pcs_txclk_freerun),
				.txpcs_urst(hssi_8g_tx_pcs_txpcs_urst)
			) inst_twentynm_hssi_8g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_8g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_tx_pcs_blockselect),
				.clk_out(w_hssi_8g_tx_pcs_clk_out),
				.clk_out_gen3(w_hssi_8g_tx_pcs_clk_out_gen3),
				.dataout(w_hssi_8g_tx_pcs_dataout),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.fifo_select_out_chnl_down(w_hssi_8g_tx_pcs_fifo_select_out_chnl_down),
				.fifo_select_out_chnl_up(w_hssi_8g_tx_pcs_fifo_select_out_chnl_up),
				.g3_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.g3_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
				.non_gray_eidleinfersel(w_hssi_8g_tx_pcs_non_gray_eidleinfersel),
				.ph_fifo_overflow(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.ph_fifo_underflow(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.phfifo_txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.phfifo_txmargin(w_hssi_8g_tx_pcs_phfifo_txmargin),
				.phfifo_txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				.pipe_en_rev_parallel_lpbk_out(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.pipe_power_down_out(w_hssi_8g_tx_pcs_pipe_power_down_out),
				.pipe_tx_clk_out_gen3(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pmaif_asn_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.rd_enable_out_chnl_down(w_hssi_8g_tx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_tx_pcs_rd_enable_out_chnl_up),
				.rd_ptr_tx_phfifo(w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rxpolarity_int(w_hssi_8g_tx_pcs_rxpolarity_int),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.tx_blk_start_out(w_hssi_8g_tx_pcs_tx_blk_start_out),
				.tx_clk_out_8g_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.tx_ctrlplane_testbus(w_hssi_8g_tx_pcs_tx_ctrlplane_testbus),
				.tx_data_out(w_hssi_8g_tx_pcs_tx_data_out),
				.tx_data_valid_out(w_hssi_8g_tx_pcs_tx_data_valid_out),
				.tx_datak_out(w_hssi_8g_tx_pcs_tx_datak_out),
				.tx_detect_rxloopback_int(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.tx_div_sync(w_hssi_8g_tx_pcs_tx_div_sync),
				.tx_div_sync_out_chnl_down(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down),
				.tx_div_sync_out_chnl_up(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up),
				.tx_pipe_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.tx_pipe_electidle(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_soft_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.tx_sync_hdr_out(w_hssi_8g_tx_pcs_tx_sync_hdr_out),
				.tx_testbus(w_hssi_8g_tx_pcs_tx_testbus),
				.txcompliance_out(w_hssi_8g_tx_pcs_txcompliance_out),
				.txelecidle_out(w_hssi_8g_tx_pcs_txelecidle_out),
				.wr_clk_tx_phfifo_dw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_tx_phfifo_sw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_data_tx_phfifo(w_hssi_8g_tx_pcs_wr_data_tx_phfifo),
				.wr_en_tx_phfifo(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_tx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_tx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_tx_phfifo(w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo),
				.wr_rst_n_tx_phfifo(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bitslip_boundary_select({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0]}),
				.clk_sel_gen3(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.coreclk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.datain({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.detectrxloopin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidleinfersel({w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0]}),
				.en_rev_parallel_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.fifo_select_in_chnl_down({in_bond_pcs8g_in_bot[11], in_bond_pcs8g_in_bot[10]}),
				.fifo_select_in_chnl_up({in_bond_pcs8g_in_top[11], in_bond_pcs8g_in_top[10]}),
				.hrdrst(1'b0),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.ph_fifo_rd_disable(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.pipe_en_rev_parallel_lpbk_in(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.pipe_tx_deemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.pipe_tx_margin({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0]}),
				.powerdn({w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0]}),
				.rate_switch(w_hssi_8g_rx_pcs_gen2ngen1),
				.rd_data_tx_phfifo({w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[9]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[9]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.rev_parallel_lpbk_data({w_hssi_8g_rx_pcs_parallel_rev_loopback[19], w_hssi_8g_rx_pcs_parallel_rev_loopback[18], w_hssi_8g_rx_pcs_parallel_rev_loopback[17], w_hssi_8g_rx_pcs_parallel_rev_loopback[16], w_hssi_8g_rx_pcs_parallel_rev_loopback[15], w_hssi_8g_rx_pcs_parallel_rev_loopback[14], w_hssi_8g_rx_pcs_parallel_rev_loopback[13], w_hssi_8g_rx_pcs_parallel_rev_loopback[12], w_hssi_8g_rx_pcs_parallel_rev_loopback[11], w_hssi_8g_rx_pcs_parallel_rev_loopback[10], w_hssi_8g_rx_pcs_parallel_rev_loopback[9], w_hssi_8g_rx_pcs_parallel_rev_loopback[8], w_hssi_8g_rx_pcs_parallel_rev_loopback[7], w_hssi_8g_rx_pcs_parallel_rev_loopback[6], w_hssi_8g_rx_pcs_parallel_rev_loopback[5], w_hssi_8g_rx_pcs_parallel_rev_loopback[4], w_hssi_8g_rx_pcs_parallel_rev_loopback[3], w_hssi_8g_rx_pcs_parallel_rev_loopback[2], w_hssi_8g_rx_pcs_parallel_rev_loopback[1], w_hssi_8g_rx_pcs_parallel_rev_loopback[0]}),
				.rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.tx_blk_start({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0]}),
				.tx_data_valid({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0]}),
				.tx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[7], in_bond_pcs8g_in_bot[6]}),
				.tx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[7], in_bond_pcs8g_in_top[6]}),
				.tx_pcs_reset(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.tx_sync_hdr({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0]}),
				.txd_fast_reg({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0]}),
				.txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[8]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[8]),
				.wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				
				// UNUSED
				.byte_serializer_pcs_clk_div_by_2_reg(),
				.byte_serializer_pcs_clk_div_by_2_wire(),
				.byte_serializer_pcs_clk_div_by_4_reg(),
				.byte_serializer_pld_clk_div_by_2_reg(),
				.byte_serializer_pld_clk_div_by_4_reg(),
				.pld_8g_empty_tx_fifo(),
				.pld_8g_empty_tx_reg(),
				.pld_8g_full_tx_fifo(),
				.pld_8g_full_tx_reg(),
				.pld_8g_g3_tx_pld_rst_n_reg(),
				.pld_8g_rddisable_tx_reg(),
				.pld_8g_tx_boundary_sel_reg(),
				.pld_pcs_tx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_tx_clk_out_8g_wire(),
				.pld_tx_data_8g_fifo(),
				.pld_tx_data_lo_8g_reg(),
				.sta_tx_clk2_by2_1(),
				.sta_tx_clk2_by2_1_out(),
				.sta_tx_clk2_by4_1(),
				.sta_tx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_dataout[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_dyn_clk_switch_n = 1'b1;		// Override default tieoff
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_g3_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_overflow = 1'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_underflow = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txdeemph = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txmargin[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txswing = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_power_down_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_pmaif_asn_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_refclk_b = 1'b0;
				assign w_hssi_8g_tx_pcs_refclk_b_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_rxpolarity_int = 1'b0;
				assign w_hssi_8g_tx_pcs_soft_reset_wclk1_n = 1'b0;
				assign w_hssi_8g_tx_pcs_sw_fifo_wr_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_blk_start_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_tx_data_out[31:0] = 32'b0;
				assign w_hssi_8g_tx_pcs_tx_data_valid_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_datak_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_detect_rxloopback_int = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_electidle = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_sync_hdr_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_txcompliance_out = 1'b0;
				assign w_hssi_8g_tx_pcs_txelecidle_out = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63:0] = 64'b0;
				assign w_hssi_8g_tx_pcs_wr_en_tx_phfifo = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pcs_pma_interface
			twentynm_hssi_common_pcs_pma_interface #(
				.asn_clk_enable(hssi_common_pcs_pma_interface_asn_clk_enable),
				.asn_enable(hssi_common_pcs_pma_interface_asn_enable),
				.block_sel(hssi_common_pcs_pma_interface_block_sel),
				.bypass_early_eios(hssi_common_pcs_pma_interface_bypass_early_eios),
				.bypass_pcie_switch(hssi_common_pcs_pma_interface_bypass_pcie_switch),
				.bypass_pma_ltr(hssi_common_pcs_pma_interface_bypass_pma_ltr),
				.bypass_pma_sw_done(hssi_common_pcs_pma_interface_bypass_pma_sw_done),
				.bypass_ppm_lock(hssi_common_pcs_pma_interface_bypass_ppm_lock),
				.bypass_send_syncp_fbkp(hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp),
				.bypass_txdetectrx(hssi_common_pcs_pma_interface_bypass_txdetectrx),
				.cdr_control(hssi_common_pcs_pma_interface_cdr_control),
				.cid_enable(hssi_common_pcs_pma_interface_cid_enable),
				.cp_cons_sel(hssi_common_pcs_pma_interface_cp_cons_sel),
				.cp_dwn_mstr(hssi_common_pcs_pma_interface_cp_dwn_mstr),
				.cp_up_mstr(hssi_common_pcs_pma_interface_cp_up_mstr),
				.ctrl_plane_bonding(hssi_common_pcs_pma_interface_ctrl_plane_bonding),
				.data_mask_count(hssi_common_pcs_pma_interface_data_mask_count),
				.data_mask_count_multi(hssi_common_pcs_pma_interface_data_mask_count_multi),
				.dft_observation_clock_selection(hssi_common_pcs_pma_interface_dft_observation_clock_selection),
				.early_eios_counter(hssi_common_pcs_pma_interface_early_eios_counter),
				.force_freqdet(hssi_common_pcs_pma_interface_force_freqdet),
				.free_run_clk_enable(hssi_common_pcs_pma_interface_free_run_clk_enable),
				.ignore_sigdet_g23(hssi_common_pcs_pma_interface_ignore_sigdet_g23),
				.pc_en_counter(hssi_common_pcs_pma_interface_pc_en_counter),
				.pc_rst_counter(hssi_common_pcs_pma_interface_pc_rst_counter),
				.pcie_hip_mode(hssi_common_pcs_pma_interface_pcie_hip_mode),
				.ph_fifo_reg_mode(hssi_common_pcs_pma_interface_ph_fifo_reg_mode),
				.phfifo_flush_wait(hssi_common_pcs_pma_interface_phfifo_flush_wait),
				.pipe_if_g3pcs(hssi_common_pcs_pma_interface_pipe_if_g3pcs),
				.pma_done_counter(hssi_common_pcs_pma_interface_pma_done_counter),
				.pma_if_dft_en(hssi_common_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_common_pcs_pma_interface_pma_if_dft_val),
				.ppm_cnt_rst(hssi_common_pcs_pma_interface_ppm_cnt_rst),
				.ppm_deassert_early(hssi_common_pcs_pma_interface_ppm_deassert_early),
				.ppm_det_buckets(hssi_common_pcs_pma_interface_ppm_det_buckets),
				.ppm_gen1_2_cnt(hssi_common_pcs_pma_interface_ppm_gen1_2_cnt),
				.ppm_post_eidle_delay(hssi_common_pcs_pma_interface_ppm_post_eidle_delay),
				.ppmsel(hssi_common_pcs_pma_interface_ppmsel),
				.prot_mode(hssi_common_pcs_pma_interface_prot_mode),
				.reconfig_settings(hssi_common_pcs_pma_interface_reconfig_settings),
				.rxvalid_mask(hssi_common_pcs_pma_interface_rxvalid_mask),
				.sigdet_wait_counter(hssi_common_pcs_pma_interface_sigdet_wait_counter),
				.sigdet_wait_counter_multi(hssi_common_pcs_pma_interface_sigdet_wait_counter_multi),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sim_mode(hssi_common_pcs_pma_interface_sim_mode),
				.spd_chg_rst_wait_cnt_en(hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en),
				.sup_mode(hssi_common_pcs_pma_interface_sup_mode),
				.testout_sel(hssi_common_pcs_pma_interface_testout_sel),
				.wait_clk_on_off_timer(hssi_common_pcs_pma_interface_wait_clk_on_off_timer),
				.wait_pipe_synchronizing(hssi_common_pcs_pma_interface_wait_pipe_synchronizing),
				.wait_send_syncp_fbkp(hssi_common_pcs_pma_interface_wait_send_syncp_fbkp)
			) inst_twentynm_hssi_common_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_common_pcs_pma_interface_blockselect),
				.int_pmaif_8g_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in),
				.int_pmaif_8g_eios_detected(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.int_pmaif_8g_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.int_pmaif_8g_power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.int_pmaif_g3_pcs_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in),
				.int_pmaif_pldif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pmaif_pldif_pcie_sw_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done),
				.int_pmaif_pldif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pmaif_pldif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pmaif_pldif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pmaif_pldif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pmaif_pldif_pma_reserved_in(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in),
				.int_pmaif_pldif_test_out(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out),
				.int_pmaif_pldif_testbus(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus),
				.pma_adapt_start(w_hssi_common_pcs_pma_interface_pma_adapt_start),
				.pma_atpg_los_en_n(w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n),
				.pma_csr_test_dis(w_hssi_common_pcs_pma_interface_pma_csr_test_dis),
				.pma_current_coeff(w_hssi_common_pcs_pma_interface_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_common_pcs_pma_interface_pma_current_rxpreset),
				.pma_early_eios(w_hssi_common_pcs_pma_interface_pma_early_eios),
				.pma_interface_select(w_hssi_common_pcs_pma_interface_pma_interface_select),
				.pma_ltd_b(w_hssi_common_pcs_pma_interface_pma_ltd_b),
				.pma_ltr(w_hssi_common_pcs_pma_interface_pma_ltr),
				.pma_nfrzdrv(w_hssi_common_pcs_pma_interface_pma_nfrzdrv),
				.pma_nrpi_freeze(w_hssi_common_pcs_pma_interface_pma_nrpi_freeze),
				.pma_pcie_switch(w_hssi_common_pcs_pma_interface_pma_pcie_switch),
				.pma_ppm_lock(w_hssi_common_pcs_pma_interface_pma_ppm_lock),
				.pma_reserved_out(w_hssi_common_pcs_pma_interface_pma_reserved_out),
				.pma_rs_lpbk_b(w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b),
				.pma_rx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup),
				.pma_scan_mode_n(w_hssi_common_pcs_pma_interface_pma_scan_mode_n),
				.pma_scan_shift_n(w_hssi_common_pcs_pma_interface_pma_scan_shift_n),
				.pma_tx_bitslip(w_hssi_common_pcs_pma_interface_pma_tx_bitslip),
				.pma_tx_bonding_rstb(w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb),
				.pma_tx_qpi_pulldn(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn),
				.pma_tx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup),
				.pma_tx_txdetectrx(w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx),
				.pmaif_bundling_out_down(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down),
				.pmaif_bundling_out_up(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_8g_current_coeff({w_hssi_pipe_gen1_2_current_coeff[17], w_hssi_pipe_gen1_2_current_coeff[16], w_hssi_pipe_gen1_2_current_coeff[15], w_hssi_pipe_gen1_2_current_coeff[14], w_hssi_pipe_gen1_2_current_coeff[13], w_hssi_pipe_gen1_2_current_coeff[12], w_hssi_pipe_gen1_2_current_coeff[11], w_hssi_pipe_gen1_2_current_coeff[10], w_hssi_pipe_gen1_2_current_coeff[9], w_hssi_pipe_gen1_2_current_coeff[8], w_hssi_pipe_gen1_2_current_coeff[7], w_hssi_pipe_gen1_2_current_coeff[6], w_hssi_pipe_gen1_2_current_coeff[5], w_hssi_pipe_gen1_2_current_coeff[4], w_hssi_pipe_gen1_2_current_coeff[3], w_hssi_pipe_gen1_2_current_coeff[2], w_hssi_pipe_gen1_2_current_coeff[1], w_hssi_pipe_gen1_2_current_coeff[0]}),
				.int_pmaif_8g_eios_det({w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0]}),
				.int_pmaif_8g_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.int_pmaif_8g_rev_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.int_pmaif_8g_tx_clk_out_gen3(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.int_pmaif_8g_txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				.int_pmaif_g3_eios_det({w_hssi_gen3_rx_pcs_ei_det_int, w_hssi_gen3_rx_pcs_ei_partial_det_int, w_hssi_gen3_rx_pcs_i_det_int}),
				.int_pmaif_g3_pma_current_coeff({w_hssi_pipe_gen3_pma_current_coeff[17], w_hssi_pipe_gen3_pma_current_coeff[16], w_hssi_pipe_gen3_pma_current_coeff[15], w_hssi_pipe_gen3_pma_current_coeff[14], w_hssi_pipe_gen3_pma_current_coeff[13], w_hssi_pipe_gen3_pma_current_coeff[12], w_hssi_pipe_gen3_pma_current_coeff[11], w_hssi_pipe_gen3_pma_current_coeff[10], w_hssi_pipe_gen3_pma_current_coeff[9], w_hssi_pipe_gen3_pma_current_coeff[8], w_hssi_pipe_gen3_pma_current_coeff[7], w_hssi_pipe_gen3_pma_current_coeff[6], w_hssi_pipe_gen3_pma_current_coeff[5], w_hssi_pipe_gen3_pma_current_coeff[4], w_hssi_pipe_gen3_pma_current_coeff[3], w_hssi_pipe_gen3_pma_current_coeff[2], w_hssi_pipe_gen3_pma_current_coeff[1], w_hssi_pipe_gen3_pma_current_coeff[0]}),
				.int_pmaif_g3_pma_current_rxpreset({w_hssi_pipe_gen3_pma_current_rxpreset[2], w_hssi_pipe_gen3_pma_current_rxpreset[1], w_hssi_pipe_gen3_pma_current_rxpreset[0]}),
				.int_pmaif_g3_pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.int_pmaif_g3_rev_lpbk(w_hssi_pipe_gen3_rev_lpbk_int),
				.int_pmaif_pldif_8g_tx_pld_rstn(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pmaif_pldif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pmaif_pldif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pmaif_pldif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pmaif_pldif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pmaif_pldif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pmaif_pldif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pmaif_pldif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pmaif_pldif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pmaif_pldif_pcie_switch({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0]}),
				.int_pmaif_pldif_pma_reserved_out({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0]}),
				.int_pmaif_pldif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pmaif_pldif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pmaif_pldif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pmaif_pldif_rate({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0]}),
				.int_pmaif_pldif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pmaif_pldif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pmaif_pldif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.int_pmaif_pldif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pmaif_pldif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pmaif_pldif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pmaif_pldif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pmaif_pldif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pmaif_pldif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.int_tx_dft_obsrv_clk({w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0]}),
				.iocsr_clk(in_iocsr_clk),
				.iocsr_config({in_iocsr_config[5], in_iocsr_config[4], in_iocsr_config[3], in_iocsr_config[2], in_iocsr_config[1], in_iocsr_config[0]}),
				.iocsr_rdy(in_iocsr_rdy),
				.iocsr_rdy_dly(in_iocsr_rdy_dly),
				.pma_adapt_done(in_pma_adapt_done),
				.pma_clklow(in_pma_clklow),
				.pma_fref(in_pma_fref),
				.pma_hclk(in_pma_hclk),
				.pma_pcie_sw_done({in_pma_pcie_sw_done[1], in_pma_pcie_sw_done[0]}),
				.pma_pfdmode_lock(in_pma_pfdmode_lock),
				.pma_reserved_in({in_pma_reserved_in[4], in_pma_reserved_in[3], in_pma_reserved_in[2], in_pma_reserved_in[1], in_pma_reserved_in[0]}),
				.pma_signal_det(in_pma_signal_det),
				.pma_testbus({in_pma_testbus[7], in_pma_testbus[6], in_pma_testbus[5], in_pma_testbus[4], in_pma_testbus[3], in_pma_testbus[2], in_pma_testbus[1], in_pma_testbus[0]}),
				.pmaif_bundling_in_down({in_bond_pmaif_in_bot[11], in_bond_pmaif_in_bot[10], in_bond_pmaif_in_bot[9], in_bond_pmaif_in_bot[8], in_bond_pmaif_in_bot[7], in_bond_pmaif_in_bot[6], in_bond_pmaif_in_bot[5], in_bond_pmaif_in_bot[4], in_bond_pmaif_in_bot[3], in_bond_pmaif_in_bot[2], in_bond_pmaif_in_bot[1], in_bond_pmaif_in_bot[0]}),
				.pmaif_bundling_in_up({in_bond_pmaif_in_top[11], in_bond_pmaif_in_top[10], in_bond_pmaif_in_top[9], in_bond_pmaif_in_top[8], in_bond_pmaif_in_top[7], in_bond_pmaif_in_top[6], in_bond_pmaif_in_top[5], in_bond_pmaif_in_top[4], in_bond_pmaif_in_top[3], in_bond_pmaif_in_top[2], in_bond_pmaif_in_top[1], in_bond_pmaif_in_top[0]}),
				.rx_pmaif_test_out({w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0]}),
				.rx_prbs_ver_test({w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0]}),
				.tx_prbs_gen_test({w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0]}),
				.uhsif_test_out_1({w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0]}),
				.uhsif_test_out_2({w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0]}),
				.uhsif_test_out_3({w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0]}),
				
				// UNUSED
				.int_pmaif_avmm_iocsr_clk(),
				.int_pmaif_avmm_iocsr_config(),
				.int_pmaif_avmm_iocsr_rdy(),
				.int_pmaif_avmm_iocsr_rdy_dly(),
				.int_pmaif_pldif_interface_select(),
				.pma_tx_pma_syncp(),
				.sta_pma_hclk_by2()
			);
		end // if generate
		else begin
				assign w_hssi_common_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19:0] = 20'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_pma_adapt_start = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_csr_test_dis = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pcs_pma_interface_pma_early_eios = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_interface_select[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltd_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltr = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nfrzdrv = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nrpi_freeze = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ppm_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_tx_bitslip = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx = in_pld_pma_txdetectrx;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11:0] = 12'b0;
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11:0] = 12'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pld_pcs_interface
			twentynm_hssi_common_pld_pcs_interface #(
				.dft_clk_out_en(hssi_common_pld_pcs_interface_dft_clk_out_en),
				.dft_clk_out_sel(hssi_common_pld_pcs_interface_dft_clk_out_sel),
				.hrdrstctrl_en(hssi_common_pld_pcs_interface_hrdrstctrl_en),
				.pcs_testbus_block_sel(hssi_common_pld_pcs_interface_pcs_testbus_block_sel),
				.reconfig_settings(hssi_common_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm1" )       //PARAM_HIDE
			) inst_twentynm_hssi_common_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_common_pld_pcs_interface_blockselect),
				.hip_cmn_clk(w_hssi_common_pld_pcs_interface_hip_cmn_clk),
				.hip_cmn_ctrl(w_hssi_common_pld_pcs_interface_hip_cmn_ctrl),
				.hip_iocsr_rdy(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy),
				.hip_iocsr_rdy_dly(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly),
				.hip_nfrzdrv(w_hssi_common_pld_pcs_interface_hip_nfrzdrv),
				.hip_npor(w_hssi_common_pld_pcs_interface_hip_npor),
				.hip_usermode(w_hssi_common_pld_pcs_interface_hip_usermode),
				.int_pldif_10g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.int_pldif_10g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.int_pldif_8g_eidleinfersel(w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel),
				.int_pldif_8g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.int_pldif_8g_refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.int_pldif_8g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.int_pldif_g3_current_coeff(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff),
				.int_pldif_g3_current_rxpreset(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset),
				.int_pldif_krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.int_pldif_krfec_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.int_pldif_krfec_scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				.int_pldif_mem_atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.int_pldif_mem_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.int_pldif_pmaif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pldif_pmaif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pldif_pmaif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pldif_pmaif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pldif_pmaif_eye_monitor(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor),
				.int_pldif_pmaif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pldif_pmaif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pldif_pmaif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pldif_pmaif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pldif_pmaif_pcie_switch(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch),
				.int_pldif_pmaif_pma_reserved_out(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out),
				.int_pldif_pmaif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pldif_pmaif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pldif_pmaif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pldif_pmaif_rate(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate),
				.int_pldif_pmaif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pldif_pmaif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pldif_pmaif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pldif_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_pldif_pmaif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pldif_pmaif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pldif_pmaif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pldif_pmaif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pldif_pmaif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pldif_pmaif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pldif_pmaif_uhsif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.pld_pma_adapt_done(w_hssi_common_pld_pcs_interface_pld_pma_adapt_done),
				.pld_pma_clklow(w_hssi_common_pld_pcs_interface_pld_pma_clklow),
				.pld_pma_fref(w_hssi_common_pld_pcs_interface_pld_pma_fref),
				.pld_pma_hclk(w_hssi_common_pld_pcs_interface_pld_pma_hclk),
				.pld_pma_pcie_sw_done(w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done),
				.pld_pma_pfdmode_lock(w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock),
				.pld_pma_reserved_in(w_hssi_common_pld_pcs_interface_pld_pma_reserved_in),
				.pld_pma_rx_detect_valid(w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid),
				.pld_pma_rx_found(w_hssi_common_pld_pcs_interface_pld_pma_rx_found),
				.pld_pma_rxpll_lock(w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock),
				.pld_pma_testbus(w_hssi_common_pld_pcs_interface_pld_pma_testbus),
				.pld_pmaif_mask_tx_pll(w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll),
				.pld_reserved_out(w_hssi_common_pld_pcs_interface_pld_reserved_out),
				.pld_test_data(w_hssi_common_pld_pcs_interface_pld_test_data),
				.pld_uhsif_lock(w_hssi_common_pld_pcs_interface_pld_uhsif_lock),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.int_pldif_10g_test_data({w_hssi_10g_tx_pcs_tx_test_data[19], w_hssi_10g_tx_pcs_tx_test_data[18], w_hssi_10g_tx_pcs_tx_test_data[17], w_hssi_10g_tx_pcs_tx_test_data[16], w_hssi_10g_tx_pcs_tx_test_data[15], w_hssi_10g_tx_pcs_tx_test_data[14], w_hssi_10g_tx_pcs_tx_test_data[13], w_hssi_10g_tx_pcs_tx_test_data[12], w_hssi_10g_tx_pcs_tx_test_data[11], w_hssi_10g_tx_pcs_tx_test_data[10], w_hssi_10g_tx_pcs_tx_test_data[9], w_hssi_10g_tx_pcs_tx_test_data[8], w_hssi_10g_tx_pcs_tx_test_data[7], w_hssi_10g_tx_pcs_tx_test_data[6], w_hssi_10g_tx_pcs_tx_test_data[5], w_hssi_10g_tx_pcs_tx_test_data[4], w_hssi_10g_tx_pcs_tx_test_data[3], w_hssi_10g_tx_pcs_tx_test_data[2], w_hssi_10g_tx_pcs_tx_test_data[1], w_hssi_10g_tx_pcs_tx_test_data[0]}),
				.int_pldif_10g_tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.int_pldif_8g_chnl_test_bus_out({w_hssi_8g_rx_pcs_chnl_test_bus_out[19], w_hssi_8g_rx_pcs_chnl_test_bus_out[18], w_hssi_8g_rx_pcs_chnl_test_bus_out[17], w_hssi_8g_rx_pcs_chnl_test_bus_out[16], w_hssi_8g_rx_pcs_chnl_test_bus_out[15], w_hssi_8g_rx_pcs_chnl_test_bus_out[14], w_hssi_8g_rx_pcs_chnl_test_bus_out[13], w_hssi_8g_rx_pcs_chnl_test_bus_out[12], w_hssi_8g_rx_pcs_chnl_test_bus_out[11], w_hssi_8g_rx_pcs_chnl_test_bus_out[10], w_hssi_8g_rx_pcs_chnl_test_bus_out[9], w_hssi_8g_rx_pcs_chnl_test_bus_out[8], w_hssi_8g_rx_pcs_chnl_test_bus_out[7], w_hssi_8g_rx_pcs_chnl_test_bus_out[6], w_hssi_8g_rx_pcs_chnl_test_bus_out[5], w_hssi_8g_rx_pcs_chnl_test_bus_out[4], w_hssi_8g_rx_pcs_chnl_test_bus_out[3], w_hssi_8g_rx_pcs_chnl_test_bus_out[2], w_hssi_8g_rx_pcs_chnl_test_bus_out[1], w_hssi_8g_rx_pcs_chnl_test_bus_out[0]}),
				.int_pldif_8g_rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.int_pldif_8g_tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.int_pldif_g3_test_out({w_hssi_pipe_gen3_test_out[19], w_hssi_pipe_gen3_test_out[18], w_hssi_pipe_gen3_test_out[17], w_hssi_pipe_gen3_test_out[16], w_hssi_pipe_gen3_test_out[15], w_hssi_pipe_gen3_test_out[14], w_hssi_pipe_gen3_test_out[13], w_hssi_pipe_gen3_test_out[12], w_hssi_pipe_gen3_test_out[11], w_hssi_pipe_gen3_test_out[10], w_hssi_pipe_gen3_test_out[9], w_hssi_pipe_gen3_test_out[8], w_hssi_pipe_gen3_test_out[7], w_hssi_pipe_gen3_test_out[6], w_hssi_pipe_gen3_test_out[5], w_hssi_pipe_gen3_test_out[4], w_hssi_pipe_gen3_test_out[3], w_hssi_pipe_gen3_test_out[2], w_hssi_pipe_gen3_test_out[1], w_hssi_pipe_gen3_test_out[0]}),
				.int_pldif_krfec_test_data({w_hssi_krfec_tx_pcs_tx_test_data[19], w_hssi_krfec_tx_pcs_tx_test_data[18], w_hssi_krfec_tx_pcs_tx_test_data[17], w_hssi_krfec_tx_pcs_tx_test_data[16], w_hssi_krfec_tx_pcs_tx_test_data[15], w_hssi_krfec_tx_pcs_tx_test_data[14], w_hssi_krfec_tx_pcs_tx_test_data[13], w_hssi_krfec_tx_pcs_tx_test_data[12], w_hssi_krfec_tx_pcs_tx_test_data[11], w_hssi_krfec_tx_pcs_tx_test_data[10], w_hssi_krfec_tx_pcs_tx_test_data[9], w_hssi_krfec_tx_pcs_tx_test_data[8], w_hssi_krfec_tx_pcs_tx_test_data[7], w_hssi_krfec_tx_pcs_tx_test_data[6], w_hssi_krfec_tx_pcs_tx_test_data[5], w_hssi_krfec_tx_pcs_tx_test_data[4], w_hssi_krfec_tx_pcs_tx_test_data[3], w_hssi_krfec_tx_pcs_tx_test_data[2], w_hssi_krfec_tx_pcs_tx_test_data[1], w_hssi_krfec_tx_pcs_tx_test_data[0]}),
				.int_pldif_pmaif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pldif_pmaif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pldif_pmaif_pcie_sw_done({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0]}),
				.int_pldif_pmaif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pldif_pmaif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pldif_pmaif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pldif_pmaif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pldif_pmaif_pma_reserved_in({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0]}),
				.int_pldif_pmaif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pldif_pmaif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_test_out({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0]}),
				.int_pldif_pmaif_testbus({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0]}),
				.int_pldif_pmaif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.pld_8g_eidleinfersel({in_pld_8g_eidleinfersel[2], in_pld_8g_eidleinfersel[1], in_pld_8g_eidleinfersel[0]}),
				.pld_8g_refclk_dig2(in_pld_8g_refclk_dig2),
				.pld_atpg_los_en_n(in_pld_atpg_los_en_n),
				.pld_g3_current_coeff({in_pld_g3_current_coeff[17], in_pld_g3_current_coeff[16], in_pld_g3_current_coeff[15], in_pld_g3_current_coeff[14], in_pld_g3_current_coeff[13], in_pld_g3_current_coeff[12], in_pld_g3_current_coeff[11], in_pld_g3_current_coeff[10], in_pld_g3_current_coeff[9], in_pld_g3_current_coeff[8], in_pld_g3_current_coeff[7], in_pld_g3_current_coeff[6], in_pld_g3_current_coeff[5], in_pld_g3_current_coeff[4], in_pld_g3_current_coeff[3], in_pld_g3_current_coeff[2], in_pld_g3_current_coeff[1], in_pld_g3_current_coeff[0]}),
				.pld_g3_current_rxpreset({in_pld_g3_current_rxpreset[2], in_pld_g3_current_rxpreset[1], in_pld_g3_current_rxpreset[0]}),
				.pld_ltr(in_pld_ltr),
				.pld_mem_krfec_atpg_rst_n(in_pld_mem_krfec_atpg_rst_n),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pcs_refclk_dig(in_pld_pcs_refclk_dig),
				.pld_pma_adapt_start(in_pld_pma_adapt_start),
				.pld_pma_csr_test_dis(in_pld_pma_csr_test_dis),
				.pld_pma_early_eios(in_pld_pma_early_eios),
				.pld_pma_eye_monitor({in_pld_pma_eye_monitor[5], in_pld_pma_eye_monitor[4], in_pld_pma_eye_monitor[3], in_pld_pma_eye_monitor[2], in_pld_pma_eye_monitor[1], in_pld_pma_eye_monitor[0]}),
				.pld_pma_ltd_b(in_pld_pma_ltd_b),
				.pld_pma_nrpi_freeze(in_pld_pma_nrpi_freeze),
				.pld_pma_pcie_switch({in_pld_pma_pcie_switch[1], in_pld_pma_pcie_switch[0]}),
				.pld_pma_ppm_lock(in_pld_pma_ppm_lock),
				.pld_pma_reserved_out({in_pld_pma_reserved_out[4], in_pld_pma_reserved_out[3], in_pld_pma_reserved_out[2], in_pld_pma_reserved_out[1], in_pld_pma_reserved_out[0]}),
				.pld_pma_rs_lpbk_b(in_pld_pma_rs_lpbk_b),
				.pld_pma_rx_qpi_pullup(in_pld_pma_rx_qpi_pullup),
				.pld_pma_tx_bitslip(in_pld_pma_tx_bitslip),
				.pld_pma_tx_bonding_rstb(in_pld_pma_tx_bonding_rstb),
				.pld_pma_tx_qpi_pulldn(in_pld_pma_tx_qpi_pulldn),
				.pld_pma_tx_qpi_pullup(in_pld_pma_tx_qpi_pullup),
				.pld_pma_txdetectrx(in_pld_pma_txdetectrx),
				.pld_rate({in_pld_rate[1], in_pld_rate[0]}),
				.pld_reserved_in({in_pld_reserved_in[9], in_pld_reserved_in[8], in_pld_reserved_in[7], in_pld_reserved_in[6], in_pld_reserved_in[5], in_pld_reserved_in[4], in_pld_reserved_in[3], in_pld_reserved_in[2], in_pld_reserved_in[1], in_pld_reserved_in[0]}),
				.pld_scan_mode_n(in_pld_scan_mode_n),
				.pld_scan_shift_n(in_pld_scan_shift_n),
				
				// UNUSED
				.int_pldif_8g_ltr(),
				.int_pldif_avmm_pld_avmm1_request(),
				.int_pldif_avmm_pld_avmm2_request(),
				.int_pldif_avmm_refclk_dig_en(),
				.int_pldif_g3_scan_mode_n(),
				.pld_8g_eidleinfersel_fifo(),
				.pld_8g_eidleinfersel_reg(),
				.pld_partial_reconfig_fifo(),
				.pld_partial_reconfig_rx_div_by_2_rxclk_wire(),
				.pld_partial_reconfig_rx_div_by_2_txclk_wire(),
				.pld_partial_reconfig_rxclk_reg(),
				.pld_partial_reconfig_tx_div_by_2_wire(),
				.pld_partial_reconfig_txclk_reg(),
				.pld_rate_reg(),
				.pld_test_data_reg()
			);
		end // if generate
		else begin
				assign w_hssi_common_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_clk[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_npor = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_usermode = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2 = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_adapt_done = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_clklow = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_fref = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_hclk = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_found = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_testbus[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_reserved_out[9:0] = 10'b0;
				assign w_hssi_common_pld_pcs_interface_pld_test_data[19:0] = 20'b0;
				assign w_hssi_common_pld_pcs_interface_pld_uhsif_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_scan_mode_n = 1'b1;		// Override default tieoff
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_rx_pcs
			twentynm_hssi_fifo_rx_pcs #(
				.double_read_mode(hssi_fifo_rx_pcs_double_read_mode),
				.prot_mode(hssi_fifo_rx_pcs_prot_mode),
				.silicon_rev( "20nm1" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_rx_pcs_blockselect),
				.data_out2_10g(w_hssi_fifo_rx_pcs_data_out2_10g),
				.data_out2_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp),
				.data_out_10g(w_hssi_fifo_rx_pcs_data_out_10g),
				.data_out_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out_8g_clock_comp),
				.data_out_8g_phase_comp(w_hssi_fifo_rx_pcs_data_out_8g_phase_comp),
				.data_out_gen3(w_hssi_fifo_rx_pcs_data_out_gen3),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_data[73], w_hssi_10g_rx_pcs_rx_fifo_wr_data[72], w_hssi_10g_rx_pcs_rx_fifo_wr_data[71], w_hssi_10g_rx_pcs_rx_fifo_wr_data[70], w_hssi_10g_rx_pcs_rx_fifo_wr_data[69], w_hssi_10g_rx_pcs_rx_fifo_wr_data[68], w_hssi_10g_rx_pcs_rx_fifo_wr_data[67], w_hssi_10g_rx_pcs_rx_fifo_wr_data[66], w_hssi_10g_rx_pcs_rx_fifo_wr_data[65], w_hssi_10g_rx_pcs_rx_fifo_wr_data[64], w_hssi_10g_rx_pcs_rx_fifo_wr_data[63], w_hssi_10g_rx_pcs_rx_fifo_wr_data[62], w_hssi_10g_rx_pcs_rx_fifo_wr_data[61], w_hssi_10g_rx_pcs_rx_fifo_wr_data[60], w_hssi_10g_rx_pcs_rx_fifo_wr_data[59], w_hssi_10g_rx_pcs_rx_fifo_wr_data[58], w_hssi_10g_rx_pcs_rx_fifo_wr_data[57], w_hssi_10g_rx_pcs_rx_fifo_wr_data[56], w_hssi_10g_rx_pcs_rx_fifo_wr_data[55], w_hssi_10g_rx_pcs_rx_fifo_wr_data[54], w_hssi_10g_rx_pcs_rx_fifo_wr_data[53], w_hssi_10g_rx_pcs_rx_fifo_wr_data[52], w_hssi_10g_rx_pcs_rx_fifo_wr_data[51], w_hssi_10g_rx_pcs_rx_fifo_wr_data[50], w_hssi_10g_rx_pcs_rx_fifo_wr_data[49], w_hssi_10g_rx_pcs_rx_fifo_wr_data[48], w_hssi_10g_rx_pcs_rx_fifo_wr_data[47], w_hssi_10g_rx_pcs_rx_fifo_wr_data[46], w_hssi_10g_rx_pcs_rx_fifo_wr_data[45], w_hssi_10g_rx_pcs_rx_fifo_wr_data[44], w_hssi_10g_rx_pcs_rx_fifo_wr_data[43], w_hssi_10g_rx_pcs_rx_fifo_wr_data[42], w_hssi_10g_rx_pcs_rx_fifo_wr_data[41], w_hssi_10g_rx_pcs_rx_fifo_wr_data[40], w_hssi_10g_rx_pcs_rx_fifo_wr_data[39], w_hssi_10g_rx_pcs_rx_fifo_wr_data[38], w_hssi_10g_rx_pcs_rx_fifo_wr_data[37], w_hssi_10g_rx_pcs_rx_fifo_wr_data[36], w_hssi_10g_rx_pcs_rx_fifo_wr_data[35], w_hssi_10g_rx_pcs_rx_fifo_wr_data[34], w_hssi_10g_rx_pcs_rx_fifo_wr_data[33], w_hssi_10g_rx_pcs_rx_fifo_wr_data[32], w_hssi_10g_rx_pcs_rx_fifo_wr_data[31], w_hssi_10g_rx_pcs_rx_fifo_wr_data[30], w_hssi_10g_rx_pcs_rx_fifo_wr_data[29], w_hssi_10g_rx_pcs_rx_fifo_wr_data[28], w_hssi_10g_rx_pcs_rx_fifo_wr_data[27], w_hssi_10g_rx_pcs_rx_fifo_wr_data[26], w_hssi_10g_rx_pcs_rx_fifo_wr_data[25], w_hssi_10g_rx_pcs_rx_fifo_wr_data[24], w_hssi_10g_rx_pcs_rx_fifo_wr_data[23], w_hssi_10g_rx_pcs_rx_fifo_wr_data[22], w_hssi_10g_rx_pcs_rx_fifo_wr_data[21], w_hssi_10g_rx_pcs_rx_fifo_wr_data[20], w_hssi_10g_rx_pcs_rx_fifo_wr_data[19], w_hssi_10g_rx_pcs_rx_fifo_wr_data[18], w_hssi_10g_rx_pcs_rx_fifo_wr_data[17], w_hssi_10g_rx_pcs_rx_fifo_wr_data[16], w_hssi_10g_rx_pcs_rx_fifo_wr_data[15], w_hssi_10g_rx_pcs_rx_fifo_wr_data[14], w_hssi_10g_rx_pcs_rx_fifo_wr_data[13], w_hssi_10g_rx_pcs_rx_fifo_wr_data[12], w_hssi_10g_rx_pcs_rx_fifo_wr_data[11], w_hssi_10g_rx_pcs_rx_fifo_wr_data[10], w_hssi_10g_rx_pcs_rx_fifo_wr_data[9], w_hssi_10g_rx_pcs_rx_fifo_wr_data[8], w_hssi_10g_rx_pcs_rx_fifo_wr_data[7], w_hssi_10g_rx_pcs_rx_fifo_wr_data[6], w_hssi_10g_rx_pcs_rx_fifo_wr_data[5], w_hssi_10g_rx_pcs_rx_fifo_wr_data[4], w_hssi_10g_rx_pcs_rx_fifo_wr_data[3], w_hssi_10g_rx_pcs_rx_fifo_wr_data[2], w_hssi_10g_rx_pcs_rx_fifo_wr_data[1], w_hssi_10g_rx_pcs_rx_fifo_wr_data[0]}),
				.data_in_8g_clock_comp({w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0]}),
				.data_in_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr2_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0]}),
				.rd_ptr2_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0]}),
				.rd_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0]}),
				.rd_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.wr_clk_8g_clock_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_8g_clock_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.wr_en_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.wr_en_8g_clock_comp(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_en_8g_phase_comp(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.wr_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0]}),
				.wr_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0]}),
				.wr_rst_n_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.wr_rst_n_8g_clock_comp(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_n_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_rx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79:0] = 80'b0;
				assign w_hssi_fifo_rx_pcs_data_out_gen3[39:0] = 40'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_tx_pcs
			twentynm_hssi_fifo_tx_pcs #(
				.double_write_mode(hssi_fifo_tx_pcs_double_write_mode),
				.prot_mode(hssi_fifo_tx_pcs_prot_mode),
				.silicon_rev( "20nm1" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_tx_pcs_blockselect),
				.data_out_10g(w_hssi_fifo_tx_pcs_data_out_10g),
				.data_out_8g_phase_comp(w_hssi_fifo_tx_pcs_data_out_8g_phase_comp),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in2_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0]}),
				.data_in_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_en_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.wr_en_8g_phase_comp(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0]}),
				.wr_rst_n_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_tx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_tx_pcs_data_out_10g[72:0] = 73'b0;
				assign w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63:0] = 64'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_rx_pcs
			twentynm_hssi_gen3_rx_pcs #(
				.block_sync(hssi_gen3_rx_pcs_block_sync),
				.block_sync_sm(hssi_gen3_rx_pcs_block_sync_sm),
				.cdr_ctrl_force_unalgn(hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn),
				.lpbk_force(hssi_gen3_rx_pcs_lpbk_force),
				.mode(hssi_gen3_rx_pcs_mode),
				.rate_match_fifo(hssi_gen3_rx_pcs_rate_match_fifo),
				.rate_match_fifo_latency(hssi_gen3_rx_pcs_rate_match_fifo_latency),
				.reconfig_settings(hssi_gen3_rx_pcs_reconfig_settings),
				.reverse_lpbk(hssi_gen3_rx_pcs_reverse_lpbk),
				.rx_b4gb_par_lpbk(hssi_gen3_rx_pcs_rx_b4gb_par_lpbk),
				.rx_force_balign(hssi_gen3_rx_pcs_rx_force_balign),
				.rx_ins_del_one_skip(hssi_gen3_rx_pcs_rx_ins_del_one_skip),
				.rx_num_fixed_pat(hssi_gen3_rx_pcs_rx_num_fixed_pat),
				.rx_test_out_sel(hssi_gen3_rx_pcs_rx_test_out_sel),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_rx_pcs_sup_mode)
			) inst_twentynm_hssi_gen3_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_rx_pcs_avmmreaddata),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.blk_start(w_hssi_gen3_rx_pcs_blk_start),
				.blockselect(w_hssi_gen3_rx_pcs_blockselect),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.data_out(w_hssi_gen3_rx_pcs_data_out),
				.data_valid(w_hssi_gen3_rx_pcs_data_valid),
				.ei_det_int(w_hssi_gen3_rx_pcs_ei_det_int),
				.ei_partial_det_int(w_hssi_gen3_rx_pcs_ei_partial_det_int),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.i_det_int(w_hssi_gen3_rx_pcs_i_det_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data(w_hssi_gen3_rx_pcs_lpbk_data),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.mem_rx_fifo_rd_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr),
				.mem_rx_fifo_wr_clk(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.mem_rx_fifo_wr_data(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data),
				.mem_rx_fifo_wr_en(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.mem_rx_fifo_wr_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr),
				.mem_rx_fifo_wr_rst_n(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_test_out(w_hssi_gen3_rx_pcs_rx_test_out),
				.sync_hdr(w_hssi_gen3_rx_pcs_sync_hdr),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0]}),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.mem_rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_gen3[39], w_hssi_fifo_rx_pcs_data_out_gen3[38], w_hssi_fifo_rx_pcs_data_out_gen3[37], w_hssi_fifo_rx_pcs_data_out_gen3[36], w_hssi_fifo_rx_pcs_data_out_gen3[35], w_hssi_fifo_rx_pcs_data_out_gen3[34], w_hssi_fifo_rx_pcs_data_out_gen3[33], w_hssi_fifo_rx_pcs_data_out_gen3[32], w_hssi_fifo_rx_pcs_data_out_gen3[31], w_hssi_fifo_rx_pcs_data_out_gen3[30], w_hssi_fifo_rx_pcs_data_out_gen3[29], w_hssi_fifo_rx_pcs_data_out_gen3[28], w_hssi_fifo_rx_pcs_data_out_gen3[27], w_hssi_fifo_rx_pcs_data_out_gen3[26], w_hssi_fifo_rx_pcs_data_out_gen3[25], w_hssi_fifo_rx_pcs_data_out_gen3[24], w_hssi_fifo_rx_pcs_data_out_gen3[23], w_hssi_fifo_rx_pcs_data_out_gen3[22], w_hssi_fifo_rx_pcs_data_out_gen3[21], w_hssi_fifo_rx_pcs_data_out_gen3[20], w_hssi_fifo_rx_pcs_data_out_gen3[19], w_hssi_fifo_rx_pcs_data_out_gen3[18], w_hssi_fifo_rx_pcs_data_out_gen3[17], w_hssi_fifo_rx_pcs_data_out_gen3[16], w_hssi_fifo_rx_pcs_data_out_gen3[15], w_hssi_fifo_rx_pcs_data_out_gen3[14], w_hssi_fifo_rx_pcs_data_out_gen3[13], w_hssi_fifo_rx_pcs_data_out_gen3[12], w_hssi_fifo_rx_pcs_data_out_gen3[11], w_hssi_fifo_rx_pcs_data_out_gen3[10], w_hssi_fifo_rx_pcs_data_out_gen3[9], w_hssi_fifo_rx_pcs_data_out_gen3[8], w_hssi_fifo_rx_pcs_data_out_gen3[7], w_hssi_fifo_rx_pcs_data_out_gen3[6], w_hssi_fifo_rx_pcs_data_out_gen3[5], w_hssi_fifo_rx_pcs_data_out_gen3[4], w_hssi_fifo_rx_pcs_data_out_gen3[3], w_hssi_fifo_rx_pcs_data_out_gen3[2], w_hssi_fifo_rx_pcs_data_out_gen3[1], w_hssi_fifo_rx_pcs_data_out_gen3[0]}),
				.par_lpbk_b4gb_in({w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0]}),
				.par_lpbk_in({w_hssi_gen3_tx_pcs_par_lpbk_out[31], w_hssi_gen3_tx_pcs_par_lpbk_out[30], w_hssi_gen3_tx_pcs_par_lpbk_out[29], w_hssi_gen3_tx_pcs_par_lpbk_out[28], w_hssi_gen3_tx_pcs_par_lpbk_out[27], w_hssi_gen3_tx_pcs_par_lpbk_out[26], w_hssi_gen3_tx_pcs_par_lpbk_out[25], w_hssi_gen3_tx_pcs_par_lpbk_out[24], w_hssi_gen3_tx_pcs_par_lpbk_out[23], w_hssi_gen3_tx_pcs_par_lpbk_out[22], w_hssi_gen3_tx_pcs_par_lpbk_out[21], w_hssi_gen3_tx_pcs_par_lpbk_out[20], w_hssi_gen3_tx_pcs_par_lpbk_out[19], w_hssi_gen3_tx_pcs_par_lpbk_out[18], w_hssi_gen3_tx_pcs_par_lpbk_out[17], w_hssi_gen3_tx_pcs_par_lpbk_out[16], w_hssi_gen3_tx_pcs_par_lpbk_out[15], w_hssi_gen3_tx_pcs_par_lpbk_out[14], w_hssi_gen3_tx_pcs_par_lpbk_out[13], w_hssi_gen3_tx_pcs_par_lpbk_out[12], w_hssi_gen3_tx_pcs_par_lpbk_out[11], w_hssi_gen3_tx_pcs_par_lpbk_out[10], w_hssi_gen3_tx_pcs_par_lpbk_out[9], w_hssi_gen3_tx_pcs_par_lpbk_out[8], w_hssi_gen3_tx_pcs_par_lpbk_out[7], w_hssi_gen3_tx_pcs_par_lpbk_out[6], w_hssi_gen3_tx_pcs_par_lpbk_out[5], w_hssi_gen3_tx_pcs_par_lpbk_out[4], w_hssi_gen3_tx_pcs_par_lpbk_out[3], w_hssi_gen3_tx_pcs_par_lpbk_out[2], w_hssi_gen3_tx_pcs_par_lpbk_out[1], w_hssi_gen3_tx_pcs_par_lpbk_out[0]}),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.rcvd_clk(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_pma_clk(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.rxpolarity(w_hssi_pipe_gen3_rxpolarity_int),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.sync_sm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.txdatak_in({w_hssi_pipe_gen3_txdatak_int[3], w_hssi_pipe_gen3_txdatak_int[2], w_hssi_pipe_gen3_txdatak_int[1], w_hssi_pipe_gen3_txdatak_int[0]}),
				
				// UNUSED
				.blk_lockd_int(),
				.skp_det_int()
			);
		end // if generate
		else begin
				assign w_hssi_gen3_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_rx_pcs_blk_algnd_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_delete_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_insert_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_overfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_undfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_rx_pcs_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_partial_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_err_decode_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_i_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data[33:0] = 34'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39:0] = 40'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_rx_test_out[19:0] = 20'b0;
				assign w_hssi_gen3_rx_pcs_sync_hdr[1:0] = 2'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_tx_pcs
			twentynm_hssi_gen3_tx_pcs #(
				.mode(hssi_gen3_tx_pcs_mode),
				.reverse_lpbk(hssi_gen3_tx_pcs_reverse_lpbk),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_tx_pcs_sup_mode),
				.tx_bitslip(hssi_gen3_tx_pcs_tx_bitslip),
				.tx_gbox_byp(hssi_gen3_tx_pcs_tx_gbox_byp)
			) inst_twentynm_hssi_gen3_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_gen3_tx_pcs_blockselect),
				.data_out(w_hssi_gen3_tx_pcs_data_out),
				.par_lpbk_b4gb_out(w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out),
				.par_lpbk_out(w_hssi_gen3_tx_pcs_par_lpbk_out),
				.tx_test_out(w_hssi_gen3_tx_pcs_tx_test_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_start_in(w_hssi_pipe_gen3_tx_blk_start_int),
				.data_in({w_hssi_pipe_gen3_txdata_int[31], w_hssi_pipe_gen3_txdata_int[30], w_hssi_pipe_gen3_txdata_int[29], w_hssi_pipe_gen3_txdata_int[28], w_hssi_pipe_gen3_txdata_int[27], w_hssi_pipe_gen3_txdata_int[26], w_hssi_pipe_gen3_txdata_int[25], w_hssi_pipe_gen3_txdata_int[24], w_hssi_pipe_gen3_txdata_int[23], w_hssi_pipe_gen3_txdata_int[22], w_hssi_pipe_gen3_txdata_int[21], w_hssi_pipe_gen3_txdata_int[20], w_hssi_pipe_gen3_txdata_int[19], w_hssi_pipe_gen3_txdata_int[18], w_hssi_pipe_gen3_txdata_int[17], w_hssi_pipe_gen3_txdata_int[16], w_hssi_pipe_gen3_txdata_int[15], w_hssi_pipe_gen3_txdata_int[14], w_hssi_pipe_gen3_txdata_int[13], w_hssi_pipe_gen3_txdata_int[12], w_hssi_pipe_gen3_txdata_int[11], w_hssi_pipe_gen3_txdata_int[10], w_hssi_pipe_gen3_txdata_int[9], w_hssi_pipe_gen3_txdata_int[8], w_hssi_pipe_gen3_txdata_int[7], w_hssi_pipe_gen3_txdata_int[6], w_hssi_pipe_gen3_txdata_int[5], w_hssi_pipe_gen3_txdata_int[4], w_hssi_pipe_gen3_txdata_int[3], w_hssi_pipe_gen3_txdata_int[2], w_hssi_pipe_gen3_txdata_int[1], w_hssi_pipe_gen3_txdata_int[0]}),
				.data_valid(w_hssi_pipe_gen3_txdataskip_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data_in({w_hssi_gen3_rx_pcs_lpbk_data[33], w_hssi_gen3_rx_pcs_lpbk_data[32], w_hssi_gen3_rx_pcs_lpbk_data[31], w_hssi_gen3_rx_pcs_lpbk_data[30], w_hssi_gen3_rx_pcs_lpbk_data[29], w_hssi_gen3_rx_pcs_lpbk_data[28], w_hssi_gen3_rx_pcs_lpbk_data[27], w_hssi_gen3_rx_pcs_lpbk_data[26], w_hssi_gen3_rx_pcs_lpbk_data[25], w_hssi_gen3_rx_pcs_lpbk_data[24], w_hssi_gen3_rx_pcs_lpbk_data[23], w_hssi_gen3_rx_pcs_lpbk_data[22], w_hssi_gen3_rx_pcs_lpbk_data[21], w_hssi_gen3_rx_pcs_lpbk_data[20], w_hssi_gen3_rx_pcs_lpbk_data[19], w_hssi_gen3_rx_pcs_lpbk_data[18], w_hssi_gen3_rx_pcs_lpbk_data[17], w_hssi_gen3_rx_pcs_lpbk_data[16], w_hssi_gen3_rx_pcs_lpbk_data[15], w_hssi_gen3_rx_pcs_lpbk_data[14], w_hssi_gen3_rx_pcs_lpbk_data[13], w_hssi_gen3_rx_pcs_lpbk_data[12], w_hssi_gen3_rx_pcs_lpbk_data[11], w_hssi_gen3_rx_pcs_lpbk_data[10], w_hssi_gen3_rx_pcs_lpbk_data[9], w_hssi_gen3_rx_pcs_lpbk_data[8], w_hssi_gen3_rx_pcs_lpbk_data[7], w_hssi_gen3_rx_pcs_lpbk_data[6], w_hssi_gen3_rx_pcs_lpbk_data[5], w_hssi_gen3_rx_pcs_lpbk_data[4], w_hssi_gen3_rx_pcs_lpbk_data[3], w_hssi_gen3_rx_pcs_lpbk_data[2], w_hssi_gen3_rx_pcs_lpbk_data[1], w_hssi_gen3_rx_pcs_lpbk_data[0]}),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.sync_in({w_hssi_pipe_gen3_tx_sync_hdr_int[1], w_hssi_pipe_gen3_tx_sync_hdr_int[0]}),
				.tx_pma_clk(w_hssi_8g_tx_pcs_clk_out_gen3),
				.tx_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn)
			);
		end // if generate
		else begin
				assign w_hssi_gen3_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_tx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_tx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35:0] = 36'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_tx_test_out[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_rx_pcs
			twentynm_hssi_krfec_rx_pcs #(
				.blksync_cor_en(hssi_krfec_rx_pcs_blksync_cor_en),
				.bypass_gb(hssi_krfec_rx_pcs_bypass_gb),
				.clr_ctrl(hssi_krfec_rx_pcs_clr_ctrl),
				.ctrl_bit_reverse(hssi_krfec_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_rx_pcs_data_bit_reverse),
				.dv_start(hssi_krfec_rx_pcs_dv_start),
				.err_mark_type(hssi_krfec_rx_pcs_err_mark_type),
				.error_marking_en(hssi_krfec_rx_pcs_error_marking_en),
				.low_latency_en(hssi_krfec_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_krfec_rx_pcs_lpbk_mode),
				.parity_invalid_enum(hssi_krfec_rx_pcs_parity_invalid_enum),
				.parity_valid_num(hssi_krfec_rx_pcs_parity_valid_num),
				.pipeln_blksync(hssi_krfec_rx_pcs_pipeln_blksync),
				.pipeln_descrm(hssi_krfec_rx_pcs_pipeln_descrm),
				.pipeln_errcorrect(hssi_krfec_rx_pcs_pipeln_errcorrect),
				.pipeln_errtrap_ind(hssi_krfec_rx_pcs_pipeln_errtrap_ind),
				.pipeln_errtrap_lfsr(hssi_krfec_rx_pcs_pipeln_errtrap_lfsr),
				.pipeln_errtrap_loc(hssi_krfec_rx_pcs_pipeln_errtrap_loc),
				.pipeln_errtrap_pat(hssi_krfec_rx_pcs_pipeln_errtrap_pat),
				.pipeln_gearbox(hssi_krfec_rx_pcs_pipeln_gearbox),
				.pipeln_syndrm(hssi_krfec_rx_pcs_pipeln_syndrm),
				.pipeln_trans_dec(hssi_krfec_rx_pcs_pipeln_trans_dec),
				.prot_mode(hssi_krfec_rx_pcs_prot_mode),
				.receive_order(hssi_krfec_rx_pcs_receive_order),
				.reconfig_settings(hssi_krfec_rx_pcs_reconfig_settings),
				.rx_testbus_sel(hssi_krfec_rx_pcs_rx_testbus_sel),
				.signal_ok_en(hssi_krfec_rx_pcs_signal_ok_en),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_rx_pcs_sup_mode)
			) inst_twentynm_hssi_krfec_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_rx_pcs_blockselect),
				.rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.rx_control_out(w_hssi_krfec_rx_pcs_rx_control_out),
				.rx_data_out(w_hssi_krfec_rx_pcs_rx_data_out),
				.rx_data_status(w_hssi_krfec_rx_pcs_rx_data_status),
				.rx_data_valid_out(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.rx_signal_ok_out(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.rx_data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0]}),
				.rx_krfec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_krfec_reg(),
				.pld_10g_krfec_rx_blk_lock_krfec_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg(),
				.pld_10g_krfec_rx_frame_krfec_reg(),
				.pld_10g_krfec_rx_frame_krfec_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_rx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_block_lock = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_control_out[9:0] = 10'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_status[1:0] = 2'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_valid_out = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_frame = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_signal_ok_out = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_tx_pcs
			twentynm_hssi_krfec_tx_pcs #(
				.burst_err(hssi_krfec_tx_pcs_burst_err),
				.burst_err_len(hssi_krfec_tx_pcs_burst_err_len),
				.ctrl_bit_reverse(hssi_krfec_tx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_tx_pcs_data_bit_reverse),
				.enc_frame_query(hssi_krfec_tx_pcs_enc_frame_query),
				.low_latency_en(hssi_krfec_tx_pcs_low_latency_en),
				.pipeln_encoder(hssi_krfec_tx_pcs_pipeln_encoder),
				.pipeln_scrambler(hssi_krfec_tx_pcs_pipeln_scrambler),
				.prot_mode(hssi_krfec_tx_pcs_prot_mode),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_tx_pcs_sup_mode),
				.transcode_err(hssi_krfec_tx_pcs_transcode_err),
				.transmit_order(hssi_krfec_tx_pcs_transmit_order),
				.tx_testbus_sel(hssi_krfec_tx_pcs_tx_testbus_sel)
			) inst_twentynm_hssi_krfec_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_tx_pcs_blockselect),
				.tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.tx_data_out(w_hssi_krfec_tx_pcs_tx_data_out),
				.tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.tx_test_data(w_hssi_krfec_tx_pcs_tx_test_data),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.tx_control_in({w_hssi_10g_tx_pcs_tx_control_out_krfec[8], w_hssi_10g_tx_pcs_tx_control_out_krfec[7], w_hssi_10g_tx_pcs_tx_control_out_krfec[6], w_hssi_10g_tx_pcs_tx_control_out_krfec[5], w_hssi_10g_tx_pcs_tx_control_out_krfec[4], w_hssi_10g_tx_pcs_tx_control_out_krfec[3], w_hssi_10g_tx_pcs_tx_control_out_krfec[2], w_hssi_10g_tx_pcs_tx_control_out_krfec[1], w_hssi_10g_tx_pcs_tx_control_out_krfec[0]}),
				.tx_data_in({w_hssi_10g_tx_pcs_tx_data_out_krfec[63], w_hssi_10g_tx_pcs_tx_data_out_krfec[62], w_hssi_10g_tx_pcs_tx_data_out_krfec[61], w_hssi_10g_tx_pcs_tx_data_out_krfec[60], w_hssi_10g_tx_pcs_tx_data_out_krfec[59], w_hssi_10g_tx_pcs_tx_data_out_krfec[58], w_hssi_10g_tx_pcs_tx_data_out_krfec[57], w_hssi_10g_tx_pcs_tx_data_out_krfec[56], w_hssi_10g_tx_pcs_tx_data_out_krfec[55], w_hssi_10g_tx_pcs_tx_data_out_krfec[54], w_hssi_10g_tx_pcs_tx_data_out_krfec[53], w_hssi_10g_tx_pcs_tx_data_out_krfec[52], w_hssi_10g_tx_pcs_tx_data_out_krfec[51], w_hssi_10g_tx_pcs_tx_data_out_krfec[50], w_hssi_10g_tx_pcs_tx_data_out_krfec[49], w_hssi_10g_tx_pcs_tx_data_out_krfec[48], w_hssi_10g_tx_pcs_tx_data_out_krfec[47], w_hssi_10g_tx_pcs_tx_data_out_krfec[46], w_hssi_10g_tx_pcs_tx_data_out_krfec[45], w_hssi_10g_tx_pcs_tx_data_out_krfec[44], w_hssi_10g_tx_pcs_tx_data_out_krfec[43], w_hssi_10g_tx_pcs_tx_data_out_krfec[42], w_hssi_10g_tx_pcs_tx_data_out_krfec[41], w_hssi_10g_tx_pcs_tx_data_out_krfec[40], w_hssi_10g_tx_pcs_tx_data_out_krfec[39], w_hssi_10g_tx_pcs_tx_data_out_krfec[38], w_hssi_10g_tx_pcs_tx_data_out_krfec[37], w_hssi_10g_tx_pcs_tx_data_out_krfec[36], w_hssi_10g_tx_pcs_tx_data_out_krfec[35], w_hssi_10g_tx_pcs_tx_data_out_krfec[34], w_hssi_10g_tx_pcs_tx_data_out_krfec[33], w_hssi_10g_tx_pcs_tx_data_out_krfec[32], w_hssi_10g_tx_pcs_tx_data_out_krfec[31], w_hssi_10g_tx_pcs_tx_data_out_krfec[30], w_hssi_10g_tx_pcs_tx_data_out_krfec[29], w_hssi_10g_tx_pcs_tx_data_out_krfec[28], w_hssi_10g_tx_pcs_tx_data_out_krfec[27], w_hssi_10g_tx_pcs_tx_data_out_krfec[26], w_hssi_10g_tx_pcs_tx_data_out_krfec[25], w_hssi_10g_tx_pcs_tx_data_out_krfec[24], w_hssi_10g_tx_pcs_tx_data_out_krfec[23], w_hssi_10g_tx_pcs_tx_data_out_krfec[22], w_hssi_10g_tx_pcs_tx_data_out_krfec[21], w_hssi_10g_tx_pcs_tx_data_out_krfec[20], w_hssi_10g_tx_pcs_tx_data_out_krfec[19], w_hssi_10g_tx_pcs_tx_data_out_krfec[18], w_hssi_10g_tx_pcs_tx_data_out_krfec[17], w_hssi_10g_tx_pcs_tx_data_out_krfec[16], w_hssi_10g_tx_pcs_tx_data_out_krfec[15], w_hssi_10g_tx_pcs_tx_data_out_krfec[14], w_hssi_10g_tx_pcs_tx_data_out_krfec[13], w_hssi_10g_tx_pcs_tx_data_out_krfec[12], w_hssi_10g_tx_pcs_tx_data_out_krfec[11], w_hssi_10g_tx_pcs_tx_data_out_krfec[10], w_hssi_10g_tx_pcs_tx_data_out_krfec[9], w_hssi_10g_tx_pcs_tx_data_out_krfec[8], w_hssi_10g_tx_pcs_tx_data_out_krfec[7], w_hssi_10g_tx_pcs_tx_data_out_krfec[6], w_hssi_10g_tx_pcs_tx_data_out_krfec[5], w_hssi_10g_tx_pcs_tx_data_out_krfec[4], w_hssi_10g_tx_pcs_tx_data_out_krfec[3], w_hssi_10g_tx_pcs_tx_data_out_krfec[2], w_hssi_10g_tx_pcs_tx_data_out_krfec[1], w_hssi_10g_tx_pcs_tx_data_out_krfec[0]}),
				.tx_data_valid_in(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_krfec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_krfec_reg(),
				.pld_krfec_tx_alignment_plddirect_reg(),
				.pld_krfec_tx_alignment_reg()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_tx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_alignment = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_test_data[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen1_2
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen1_2
			twentynm_hssi_pipe_gen1_2 #(
				.elec_idle_delay_val(hssi_pipe_gen1_2_elec_idle_delay_val),
				.error_replace_pad(hssi_pipe_gen1_2_error_replace_pad),
				.hip_mode(hssi_pipe_gen1_2_hip_mode),
				.ind_error_reporting(hssi_pipe_gen1_2_ind_error_reporting),
				.phystatus_delay_val(hssi_pipe_gen1_2_phystatus_delay_val),
				.phystatus_rst_toggle(hssi_pipe_gen1_2_phystatus_rst_toggle),
				.pipe_byte_de_serializer_en(hssi_pipe_gen1_2_pipe_byte_de_serializer_en),
				.prot_mode(hssi_pipe_gen1_2_prot_mode),
				.reconfig_settings(hssi_pipe_gen1_2_reconfig_settings),
				.rx_pipe_enable(hssi_pipe_gen1_2_rx_pipe_enable),
				.rxdetect_bypass(hssi_pipe_gen1_2_rxdetect_bypass),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen1_2_sup_mode),
				.tx_pipe_enable(hssi_pipe_gen1_2_tx_pipe_enable),
				.txswing(hssi_pipe_gen1_2_txswing)
			) inst_twentynm_hssi_pipe_gen1_2 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen1_2_avmmreaddata),
				.blockselect(w_hssi_pipe_gen1_2_blockselect),
				.current_coeff(w_hssi_pipe_gen1_2_current_coeff),
				.phystatus(w_hssi_pipe_gen1_2_phystatus),
				.polarity_inversion_rx(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rev_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.rxelectricalidle_out(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxstatus(w_hssi_pipe_gen1_2_rxstatus),
				.rxvalid(w_hssi_pipe_gen1_2_rxvalid),
				.tx_elec_idle_out(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pipe_rx_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.power_state_transition_done_ena(1'b0),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rev_loopbk_pcs_gen3(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.revloopback(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.rx_pipe_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rxd({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxelectricalidle(w_hssi_8g_rx_pcs_eidle_detected),
				.rxelectricalidle_pcs_gen3(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.rxpolarity_pcs_gen3(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.tx_elec_idle_comp(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.txd_ch({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswingport(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.pld_8g_rxpolarity_pipe3_reg(),
				.rxd_ch(),
				.txd()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen1_2_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen1_2_blockselect = 1'b0;
				assign w_hssi_pipe_gen1_2_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen1_2_phystatus = 1'b0;
				assign w_hssi_pipe_gen1_2_polarity_inversion_rx = 1'b0;
				assign w_hssi_pipe_gen1_2_rev_loopbk = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelectricalidle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen1_2_rxvalid = 1'b0;
				assign w_hssi_pipe_gen1_2_tx_elec_idle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_txdetectrx = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen3
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen3
			twentynm_hssi_pipe_gen3 #(
				.bypass_rx_detection_enable(hssi_pipe_gen3_bypass_rx_detection_enable),
				.bypass_rx_preset(hssi_pipe_gen3_bypass_rx_preset),
				.bypass_rx_preset_enable(hssi_pipe_gen3_bypass_rx_preset_enable),
				.bypass_tx_coefficent(hssi_pipe_gen3_bypass_tx_coefficent),
				.bypass_tx_coefficent_enable(hssi_pipe_gen3_bypass_tx_coefficent_enable),
				.elecidle_delay_g3(hssi_pipe_gen3_elecidle_delay_g3),
				.ind_error_reporting(hssi_pipe_gen3_ind_error_reporting),
				.mode(hssi_pipe_gen3_mode),
				.phy_status_delay_g12(hssi_pipe_gen3_phy_status_delay_g12),
				.phy_status_delay_g3(hssi_pipe_gen3_phy_status_delay_g3),
				.phystatus_rst_toggle_g12(hssi_pipe_gen3_phystatus_rst_toggle_g12),
				.phystatus_rst_toggle_g3(hssi_pipe_gen3_phystatus_rst_toggle_g3),
				.rate_match_pad_insertion(hssi_pipe_gen3_rate_match_pad_insertion),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen3_sup_mode),
				.test_out_sel(hssi_pipe_gen3_test_out_sel)
			) inst_twentynm_hssi_pipe_gen3 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen3_avmmreaddata),
				.blockselect(w_hssi_pipe_gen3_blockselect),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.phystatus(w_hssi_pipe_gen3_phystatus),
				.pma_current_coeff(w_hssi_pipe_gen3_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_pipe_gen3_pma_current_rxpreset),
				.pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.rev_lpbk_8gpcs_out(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.rev_lpbk_int(w_hssi_pipe_gen3_rev_lpbk_int),
				.rx_blk_start(w_hssi_pipe_gen3_rx_blk_start),
				.rx_sync_hdr(w_hssi_pipe_gen3_rx_sync_hdr),
				.rxd_8gpcs_out(w_hssi_pipe_gen3_rxd_8gpcs_out),
				.rxdataskip(w_hssi_pipe_gen3_rxdataskip),
				.rxelecidle(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity_8gpcs_out(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.rxpolarity_int(w_hssi_pipe_gen3_rxpolarity_int),
				.rxstatus(w_hssi_pipe_gen3_rxstatus),
				.rxvalid(w_hssi_pipe_gen3_rxvalid),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.test_out(w_hssi_pipe_gen3_test_out),
				.tx_blk_start_int(w_hssi_pipe_gen3_tx_blk_start_int),
				.tx_sync_hdr_int(w_hssi_pipe_gen3_tx_sync_hdr_int),
				.txdata_int(w_hssi_pipe_gen3_txdata_int),
				.txdatak_int(w_hssi_pipe_gen3_txdatak_int),
				.txdataskip_int(w_hssi_pipe_gen3_txdataskip_int),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.current_coeff({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0]}),
				.current_rxpreset({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0]}),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.pcs_asn_bundling_in({w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0]}),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pipe_tx_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_blk_start_int(w_hssi_gen3_rx_pcs_blk_start),
				.rx_sync_hdr_int({w_hssi_gen3_rx_pcs_sync_hdr[1], w_hssi_gen3_rx_pcs_sync_hdr[0]}),
				.rx_test_out({w_hssi_gen3_rx_pcs_rx_test_out[19], w_hssi_gen3_rx_pcs_rx_test_out[18], w_hssi_gen3_rx_pcs_rx_test_out[17], w_hssi_gen3_rx_pcs_rx_test_out[16], w_hssi_gen3_rx_pcs_rx_test_out[15], w_hssi_gen3_rx_pcs_rx_test_out[14], w_hssi_gen3_rx_pcs_rx_test_out[13], w_hssi_gen3_rx_pcs_rx_test_out[12], w_hssi_gen3_rx_pcs_rx_test_out[11], w_hssi_gen3_rx_pcs_rx_test_out[10], w_hssi_gen3_rx_pcs_rx_test_out[9], w_hssi_gen3_rx_pcs_rx_test_out[8], w_hssi_gen3_rx_pcs_rx_test_out[7], w_hssi_gen3_rx_pcs_rx_test_out[6], w_hssi_gen3_rx_pcs_rx_test_out[5], w_hssi_gen3_rx_pcs_rx_test_out[4], w_hssi_gen3_rx_pcs_rx_test_out[3], w_hssi_gen3_rx_pcs_rx_test_out[2], w_hssi_gen3_rx_pcs_rx_test_out[1], w_hssi_gen3_rx_pcs_rx_test_out[0]}),
				.rxd_8gpcs_in({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxdata_int({w_hssi_gen3_rx_pcs_data_out[31], w_hssi_gen3_rx_pcs_data_out[30], w_hssi_gen3_rx_pcs_data_out[29], w_hssi_gen3_rx_pcs_data_out[28], w_hssi_gen3_rx_pcs_data_out[27], w_hssi_gen3_rx_pcs_data_out[26], w_hssi_gen3_rx_pcs_data_out[25], w_hssi_gen3_rx_pcs_data_out[24], w_hssi_gen3_rx_pcs_data_out[23], w_hssi_gen3_rx_pcs_data_out[22], w_hssi_gen3_rx_pcs_data_out[21], w_hssi_gen3_rx_pcs_data_out[20], w_hssi_gen3_rx_pcs_data_out[19], w_hssi_gen3_rx_pcs_data_out[18], w_hssi_gen3_rx_pcs_data_out[17], w_hssi_gen3_rx_pcs_data_out[16], w_hssi_gen3_rx_pcs_data_out[15], w_hssi_gen3_rx_pcs_data_out[14], w_hssi_gen3_rx_pcs_data_out[13], w_hssi_gen3_rx_pcs_data_out[12], w_hssi_gen3_rx_pcs_data_out[11], w_hssi_gen3_rx_pcs_data_out[10], w_hssi_gen3_rx_pcs_data_out[9], w_hssi_gen3_rx_pcs_data_out[8], w_hssi_gen3_rx_pcs_data_out[7], w_hssi_gen3_rx_pcs_data_out[6], w_hssi_gen3_rx_pcs_data_out[5], w_hssi_gen3_rx_pcs_data_out[4], w_hssi_gen3_rx_pcs_data_out[3], w_hssi_gen3_rx_pcs_data_out[2], w_hssi_gen3_rx_pcs_data_out[1], w_hssi_gen3_rx_pcs_data_out[0]}),
				.rxdatak_int({1'b0, 1'b0, 1'b0, 1'b0}),
				.rxdataskip_int(w_hssi_gen3_rx_pcs_data_valid),
				.rxelecidle_8gpcs_in(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.tx_blk_start(w_hssi_8g_tx_pcs_tx_blk_start_out[0]),
				.tx_sync_hdr({w_hssi_8g_tx_pcs_tx_sync_hdr_out[1], w_hssi_8g_tx_pcs_tx_sync_hdr_out[0]}),
				.tx_test_out({w_hssi_gen3_tx_pcs_tx_test_out[19], w_hssi_gen3_tx_pcs_tx_test_out[18], w_hssi_gen3_tx_pcs_tx_test_out[17], w_hssi_gen3_tx_pcs_tx_test_out[16], w_hssi_gen3_tx_pcs_tx_test_out[15], w_hssi_gen3_tx_pcs_tx_test_out[14], w_hssi_gen3_tx_pcs_tx_test_out[13], w_hssi_gen3_tx_pcs_tx_test_out[12], w_hssi_gen3_tx_pcs_tx_test_out[11], w_hssi_gen3_tx_pcs_tx_test_out[10], w_hssi_gen3_tx_pcs_tx_test_out[9], w_hssi_gen3_tx_pcs_tx_test_out[8], w_hssi_gen3_tx_pcs_tx_test_out[7], w_hssi_gen3_tx_pcs_tx_test_out[6], w_hssi_gen3_tx_pcs_tx_test_out[5], w_hssi_gen3_tx_pcs_tx_test_out[4], w_hssi_gen3_tx_pcs_tx_test_out[3], w_hssi_gen3_tx_pcs_tx_test_out[2], w_hssi_gen3_tx_pcs_tx_test_out[1], w_hssi_gen3_tx_pcs_tx_test_out[0]}),
				.txcompliance(w_hssi_8g_tx_pcs_txcompliance_out),
				.txdata({w_hssi_8g_tx_pcs_tx_data_out[31], w_hssi_8g_tx_pcs_tx_data_out[30], w_hssi_8g_tx_pcs_tx_data_out[29], w_hssi_8g_tx_pcs_tx_data_out[28], w_hssi_8g_tx_pcs_tx_data_out[27], w_hssi_8g_tx_pcs_tx_data_out[26], w_hssi_8g_tx_pcs_tx_data_out[25], w_hssi_8g_tx_pcs_tx_data_out[24], w_hssi_8g_tx_pcs_tx_data_out[23], w_hssi_8g_tx_pcs_tx_data_out[22], w_hssi_8g_tx_pcs_tx_data_out[21], w_hssi_8g_tx_pcs_tx_data_out[20], w_hssi_8g_tx_pcs_tx_data_out[19], w_hssi_8g_tx_pcs_tx_data_out[18], w_hssi_8g_tx_pcs_tx_data_out[17], w_hssi_8g_tx_pcs_tx_data_out[16], w_hssi_8g_tx_pcs_tx_data_out[15], w_hssi_8g_tx_pcs_tx_data_out[14], w_hssi_8g_tx_pcs_tx_data_out[13], w_hssi_8g_tx_pcs_tx_data_out[12], w_hssi_8g_tx_pcs_tx_data_out[11], w_hssi_8g_tx_pcs_tx_data_out[10], w_hssi_8g_tx_pcs_tx_data_out[9], w_hssi_8g_tx_pcs_tx_data_out[8], w_hssi_8g_tx_pcs_tx_data_out[7], w_hssi_8g_tx_pcs_tx_data_out[6], w_hssi_8g_tx_pcs_tx_data_out[5], w_hssi_8g_tx_pcs_tx_data_out[4], w_hssi_8g_tx_pcs_tx_data_out[3], w_hssi_8g_tx_pcs_tx_data_out[2], w_hssi_8g_tx_pcs_tx_data_out[1], w_hssi_8g_tx_pcs_tx_data_out[0]}),
				.txdatak({w_hssi_8g_tx_pcs_tx_datak_out[3], w_hssi_8g_tx_pcs_tx_datak_out[2], w_hssi_8g_tx_pcs_tx_datak_out[1], w_hssi_8g_tx_pcs_tx_datak_out[0]}),
				.txdataskip(w_hssi_8g_tx_pcs_tx_data_valid_out[0]),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_8g_tx_pcs_txelecidle_out),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.dis_pc_byte(),
				.pma_rx_det_pd(),
				.pma_txdeemph(),
				.pma_txmargin(),
				.pma_txswing(),
				.reset_pc_prts()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen3_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen3_blockselect = 1'b0;
				assign w_hssi_pipe_gen3_gen3_clk_sel = 1'b0;
				assign w_hssi_pipe_gen3_pcs_rst = 1'b0;
				assign w_hssi_pipe_gen3_phystatus = 1'b0;
				assign w_hssi_pipe_gen3_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen3_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_pma_tx_elec_idle = 1'b0;
				assign w_hssi_pipe_gen3_pma_txdetectrx = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_int = 1'b0;
				assign w_hssi_pipe_gen3_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_rxd_8gpcs_out[63:0] = 64'b0;
				assign w_hssi_pipe_gen3_rxdataskip[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_int = 1'b0;
				assign w_hssi_pipe_gen3_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_rxvalid = 1'b0;
				assign w_hssi_pipe_gen3_shutdown_clk = 1'b0;
				assign w_hssi_pipe_gen3_test_out[19:0] = 20'b0;
				assign w_hssi_pipe_gen3_tx_blk_start_int = 1'b0;
				assign w_hssi_pipe_gen3_tx_sync_hdr_int[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_txdata_int[31:0] = 32'b0;
				assign w_hssi_pipe_gen3_txdatak_int[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_txdataskip_int = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pcs_pma_interface
			twentynm_hssi_rx_pcs_pma_interface #(
				.block_sel(hssi_rx_pcs_pma_interface_block_sel),
				.channel_operation_mode(hssi_rx_pcs_pma_interface_channel_operation_mode),
				.clkslip_sel(hssi_rx_pcs_pma_interface_clkslip_sel),
				.lpbk_en(hssi_rx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_rx_pcs_pma_interface_master_clk_sel),
				.pldif_datawidth_mode(hssi_rx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_rx(hssi_rx_pcs_pma_interface_pma_dw_rx),
				.pma_if_dft_en(hssi_rx_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_rx_pcs_pma_interface_pma_if_dft_val),
				.prbs9_dwidth(hssi_rx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_rx_pcs_pma_interface_prbs_clken),
				.prbs_ver(hssi_rx_pcs_pma_interface_prbs_ver),
				.prot_mode_rx(hssi_rx_pcs_pma_interface_prot_mode_rx),
				.reconfig_settings(hssi_rx_pcs_pma_interface_reconfig_settings),
				.rx_dyn_polarity_inversion(hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion),
				.rx_lpbk_en(hssi_rx_pcs_pma_interface_rx_lpbk_en),
				.rx_prbs_force_signal_ok(hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok),
				.rx_prbs_mask(hssi_rx_pcs_pma_interface_rx_prbs_mask),
				.rx_prbs_mode(hssi_rx_pcs_pma_interface_rx_prbs_mode),
				.rx_signalok_signaldet_sel(hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel),
				.rx_static_polarity_inversion(hssi_rx_pcs_pma_interface_rx_static_polarity_inversion),
				.rx_uhsif_lpbk_en(hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sup_mode(hssi_rx_pcs_pma_interface_sup_mode)
			) inst_twentynm_hssi_rx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.int_pmaif_10g_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data),
				.int_pmaif_10g_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.int_pmaif_8g_pudi(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi),
				.int_pmaif_8g_rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.int_pmaif_8g_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.int_pmaif_8g_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.int_pmaif_8g_sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.int_pmaif_g3_pma_data_in(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in),
				.int_pmaif_g3_pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.int_pmaif_g3_pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.int_pmaif_g3_pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.int_pmaif_krfec_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data),
				.int_pmaif_krfec_rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.int_pmaif_pldif_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pmaif_pldif_prbs_err_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pmaif_pldif_rx_clkdiv(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pmaif_pldif_rx_clkdiv_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pmaif_pldif_rx_data(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data),
				.int_pmaif_pldif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pmaif_pldif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pmaif_pldif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pmaif_pldif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.pma_eye_monitor(w_hssi_rx_pcs_pma_interface_pma_eye_monitor),
				.pma_rx_clkslip(w_hssi_rx_pcs_pma_interface_pma_rx_clkslip),
				.pma_rxpma_rstb(w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb),
				.rx_pmaif_test_out(w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out),
				.rx_prbs_ver_test(w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.int_pmaif_8g_rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.int_pmaif_pldif_eye_monitor({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0]}),
				.int_pmaif_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pmaif_pldif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pmaif_pldif_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pmaif_pldif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pma_rx_clkdiv_user(in_pma_rx_clkdiv_user),
				.pma_rx_detect_valid(in_pma_rx_detect_valid),
				.pma_rx_found(in_pma_rx_found),
				.pma_rx_pma_clk(in_pma_rx_pma_clk),
				.pma_rx_pma_data({in_pma_rx_pma_data[63], in_pma_rx_pma_data[62], in_pma_rx_pma_data[61], in_pma_rx_pma_data[60], in_pma_rx_pma_data[59], in_pma_rx_pma_data[58], in_pma_rx_pma_data[57], in_pma_rx_pma_data[56], in_pma_rx_pma_data[55], in_pma_rx_pma_data[54], in_pma_rx_pma_data[53], in_pma_rx_pma_data[52], in_pma_rx_pma_data[51], in_pma_rx_pma_data[50], in_pma_rx_pma_data[49], in_pma_rx_pma_data[48], in_pma_rx_pma_data[47], in_pma_rx_pma_data[46], in_pma_rx_pma_data[45], in_pma_rx_pma_data[44], in_pma_rx_pma_data[43], in_pma_rx_pma_data[42], in_pma_rx_pma_data[41], in_pma_rx_pma_data[40], in_pma_rx_pma_data[39], in_pma_rx_pma_data[38], in_pma_rx_pma_data[37], in_pma_rx_pma_data[36], in_pma_rx_pma_data[35], in_pma_rx_pma_data[34], in_pma_rx_pma_data[33], in_pma_rx_pma_data[32], in_pma_rx_pma_data[31], in_pma_rx_pma_data[30], in_pma_rx_pma_data[29], in_pma_rx_pma_data[28], in_pma_rx_pma_data[27], in_pma_rx_pma_data[26], in_pma_rx_pma_data[25], in_pma_rx_pma_data[24], in_pma_rx_pma_data[23], in_pma_rx_pma_data[22], in_pma_rx_pma_data[21], in_pma_rx_pma_data[20], in_pma_rx_pma_data[19], in_pma_rx_pma_data[18], in_pma_rx_pma_data[17], in_pma_rx_pma_data[16], in_pma_rx_pma_data[15], in_pma_rx_pma_data[14], in_pma_rx_pma_data[13], in_pma_rx_pma_data[12], in_pma_rx_pma_data[11], in_pma_rx_pma_data[10], in_pma_rx_pma_data[9], in_pma_rx_pma_data[8], in_pma_rx_pma_data[7], in_pma_rx_pma_data[6], in_pma_rx_pma_data[5], in_pma_rx_pma_data[4], in_pma_rx_pma_data[3], in_pma_rx_pma_data[2], in_pma_rx_pma_data[1], in_pma_rx_pma_data[0]}),
				.pma_rx_signal_ok(in_pma_rx_signal_ok),
				.pma_rxpll_lock(in_pma_rxpll_lock),
				.pma_signal_det(in_pma_signal_det),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.tx_pma_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0]}),
				.tx_pma_uhsif_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0]}),
				
				// UNUSED
				.int_pmaif_g3_rcvd_clk(),
				.prbs_err_lt()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31:0] = 32'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5:0] = 6'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rx_clkslip = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pld_pcs_interface
			twentynm_hssi_rx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx),
				.hd_10g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx),
				.hd_10g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx),
				.hd_10g_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx),
				.hd_10g_lpbk_en(hssi_rx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx),
				.hd_10g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx),
				.hd_10g_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx),
				.hd_10g_test_bus_mode(hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode),
				.hd_8g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx),
				.hd_8g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx),
				.hd_8g_hip_mode(hssi_rx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_rx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx),
				.hd_8g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx),
				.hd_chnl_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_clklow_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz),
				.hd_chnl_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx),
				.hd_chnl_fref_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz),
				.hd_chnl_frequency_rules_en(hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_rx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_rx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx),
				.hd_chnl_lpbk_en(hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx),
				.hd_chnl_pld_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz),
				.hd_chnl_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx),
				.hd_chnl_pma_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz),
				.hd_chnl_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx),
				.hd_chnl_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx),
				.hd_chnl_transparent_pcs_rx(hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx),
				.hd_fifo_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx),
				.hd_fifo_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx),
				.hd_g3_prot_mode(hssi_rx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx),
				.hd_krfec_lpbk_en(hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx),
				.hd_krfec_test_bus_mode(hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode),
				.hd_pldif_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx),
				.hd_pmaif_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_lpbk_en(hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx),
				.hd_pmaif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx),
				.hd_pmaif_sim_mode(hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_rx_block_sel(hssi_rx_pld_pcs_interface_pcs_rx_block_sel),
				.pcs_rx_clk_out_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel),
				.pcs_rx_clk_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_sel),
				.pcs_rx_hip_clk_en(hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en),
				.pcs_rx_output_sel(hssi_rx_pld_pcs_interface_pcs_rx_output_sel),
				.reconfig_settings(hssi_rx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm1" )       //PARAM_HIDE
			) inst_twentynm_hssi_rx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pld_pcs_interface_blockselect),
				.hip_rx_ctrl(w_hssi_rx_pld_pcs_interface_hip_rx_ctrl),
				.hip_rx_data(w_hssi_rx_pld_pcs_interface_hip_rx_data),
				.int_pldif_10g_rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.int_pldif_10g_rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.int_pldif_10g_rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.int_pldif_10g_rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.int_pldif_10g_rx_control_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb),
				.int_pldif_10g_rx_data_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb),
				.int_pldif_10g_rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.int_pldif_10g_rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.int_pldif_10g_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.int_pldif_10g_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.int_pldif_10g_rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.int_pldif_8g_a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.int_pldif_8g_bitloc_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.int_pldif_8g_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.int_pldif_8g_byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.int_pldif_8g_encdt(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.int_pldif_8g_pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.int_pldif_8g_rdenable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.int_pldif_8g_rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.int_pldif_8g_rxurstpcs_n(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.int_pldif_8g_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.int_pldif_8g_wrdisable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.int_pldif_g3_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.int_pldif_krfec_rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.int_pldif_pmaif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pldif_pmaif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pldif_pmaif_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pldif_pmaif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pld_10g_krfec_rx_blk_lock(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock),
				.pld_10g_krfec_rx_diag_data_status(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status),
				.pld_10g_krfec_rx_frame(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame),
				.pld_10g_rx_align_val(w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val),
				.pld_10g_rx_crc32_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err),
				.pld_10g_rx_data_valid(w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid),
				.pld_10g_rx_empty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty),
				.pld_10g_rx_fifo_del(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del),
				.pld_10g_rx_fifo_insert(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert),
				.pld_10g_rx_fifo_num(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num),
				.pld_10g_rx_frame_lock(w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock),
				.pld_10g_rx_hi_ber(w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber),
				.pld_10g_rx_oflw_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err),
				.pld_10g_rx_pempty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty),
				.pld_10g_rx_pfull(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull),
				.pld_8g_a1a2_k1k2_flag(w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag),
				.pld_8g_empty_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf),
				.pld_8g_empty_rx(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx),
				.pld_8g_full_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf),
				.pld_8g_full_rx(w_hssi_rx_pld_pcs_interface_pld_8g_full_rx),
				.pld_8g_rxelecidle(w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle),
				.pld_8g_signal_detect_out(w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out),
				.pld_8g_wa_boundary(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary),
				.pld_pcs_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out),
				.pld_pma_clkdiv_rx_user(w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user),
				.pld_pma_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out),
				.pld_pma_signal_ok(w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok),
				.pld_rx_control(w_hssi_rx_pld_pcs_interface_pld_rx_control),
				.pld_rx_data(w_hssi_rx_pld_pcs_interface_pld_rx_data),
				.pld_rx_prbs_done(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done),
				.pld_rx_prbs_err(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.int_pldif_10g_rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.int_pldif_10g_rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.int_pldif_10g_rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_10g_rx_control({w_hssi_10g_rx_pcs_rx_control[19], w_hssi_10g_rx_pcs_rx_control[18], w_hssi_10g_rx_pcs_rx_control[17], w_hssi_10g_rx_pcs_rx_control[16], w_hssi_10g_rx_pcs_rx_control[15], w_hssi_10g_rx_pcs_rx_control[14], w_hssi_10g_rx_pcs_rx_control[13], w_hssi_10g_rx_pcs_rx_control[12], w_hssi_10g_rx_pcs_rx_control[11], w_hssi_10g_rx_pcs_rx_control[10], w_hssi_10g_rx_pcs_rx_control[9], w_hssi_10g_rx_pcs_rx_control[8], w_hssi_10g_rx_pcs_rx_control[7], w_hssi_10g_rx_pcs_rx_control[6], w_hssi_10g_rx_pcs_rx_control[5], w_hssi_10g_rx_pcs_rx_control[4], w_hssi_10g_rx_pcs_rx_control[3], w_hssi_10g_rx_pcs_rx_control[2], w_hssi_10g_rx_pcs_rx_control[1], w_hssi_10g_rx_pcs_rx_control[0]}),
				.int_pldif_10g_rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.int_pldif_10g_rx_data({w_hssi_10g_rx_pcs_rx_data[127], w_hssi_10g_rx_pcs_rx_data[126], w_hssi_10g_rx_pcs_rx_data[125], w_hssi_10g_rx_pcs_rx_data[124], w_hssi_10g_rx_pcs_rx_data[123], w_hssi_10g_rx_pcs_rx_data[122], w_hssi_10g_rx_pcs_rx_data[121], w_hssi_10g_rx_pcs_rx_data[120], w_hssi_10g_rx_pcs_rx_data[119], w_hssi_10g_rx_pcs_rx_data[118], w_hssi_10g_rx_pcs_rx_data[117], w_hssi_10g_rx_pcs_rx_data[116], w_hssi_10g_rx_pcs_rx_data[115], w_hssi_10g_rx_pcs_rx_data[114], w_hssi_10g_rx_pcs_rx_data[113], w_hssi_10g_rx_pcs_rx_data[112], w_hssi_10g_rx_pcs_rx_data[111], w_hssi_10g_rx_pcs_rx_data[110], w_hssi_10g_rx_pcs_rx_data[109], w_hssi_10g_rx_pcs_rx_data[108], w_hssi_10g_rx_pcs_rx_data[107], w_hssi_10g_rx_pcs_rx_data[106], w_hssi_10g_rx_pcs_rx_data[105], w_hssi_10g_rx_pcs_rx_data[104], w_hssi_10g_rx_pcs_rx_data[103], w_hssi_10g_rx_pcs_rx_data[102], w_hssi_10g_rx_pcs_rx_data[101], w_hssi_10g_rx_pcs_rx_data[100], w_hssi_10g_rx_pcs_rx_data[99], w_hssi_10g_rx_pcs_rx_data[98], w_hssi_10g_rx_pcs_rx_data[97], w_hssi_10g_rx_pcs_rx_data[96], w_hssi_10g_rx_pcs_rx_data[95], w_hssi_10g_rx_pcs_rx_data[94], w_hssi_10g_rx_pcs_rx_data[93], w_hssi_10g_rx_pcs_rx_data[92], w_hssi_10g_rx_pcs_rx_data[91], w_hssi_10g_rx_pcs_rx_data[90], w_hssi_10g_rx_pcs_rx_data[89], w_hssi_10g_rx_pcs_rx_data[88], w_hssi_10g_rx_pcs_rx_data[87], w_hssi_10g_rx_pcs_rx_data[86], w_hssi_10g_rx_pcs_rx_data[85], w_hssi_10g_rx_pcs_rx_data[84], w_hssi_10g_rx_pcs_rx_data[83], w_hssi_10g_rx_pcs_rx_data[82], w_hssi_10g_rx_pcs_rx_data[81], w_hssi_10g_rx_pcs_rx_data[80], w_hssi_10g_rx_pcs_rx_data[79], w_hssi_10g_rx_pcs_rx_data[78], w_hssi_10g_rx_pcs_rx_data[77], w_hssi_10g_rx_pcs_rx_data[76], w_hssi_10g_rx_pcs_rx_data[75], w_hssi_10g_rx_pcs_rx_data[74], w_hssi_10g_rx_pcs_rx_data[73], w_hssi_10g_rx_pcs_rx_data[72], w_hssi_10g_rx_pcs_rx_data[71], w_hssi_10g_rx_pcs_rx_data[70], w_hssi_10g_rx_pcs_rx_data[69], w_hssi_10g_rx_pcs_rx_data[68], w_hssi_10g_rx_pcs_rx_data[67], w_hssi_10g_rx_pcs_rx_data[66], w_hssi_10g_rx_pcs_rx_data[65], w_hssi_10g_rx_pcs_rx_data[64], w_hssi_10g_rx_pcs_rx_data[63], w_hssi_10g_rx_pcs_rx_data[62], w_hssi_10g_rx_pcs_rx_data[61], w_hssi_10g_rx_pcs_rx_data[60], w_hssi_10g_rx_pcs_rx_data[59], w_hssi_10g_rx_pcs_rx_data[58], w_hssi_10g_rx_pcs_rx_data[57], w_hssi_10g_rx_pcs_rx_data[56], w_hssi_10g_rx_pcs_rx_data[55], w_hssi_10g_rx_pcs_rx_data[54], w_hssi_10g_rx_pcs_rx_data[53], w_hssi_10g_rx_pcs_rx_data[52], w_hssi_10g_rx_pcs_rx_data[51], w_hssi_10g_rx_pcs_rx_data[50], w_hssi_10g_rx_pcs_rx_data[49], w_hssi_10g_rx_pcs_rx_data[48], w_hssi_10g_rx_pcs_rx_data[47], w_hssi_10g_rx_pcs_rx_data[46], w_hssi_10g_rx_pcs_rx_data[45], w_hssi_10g_rx_pcs_rx_data[44], w_hssi_10g_rx_pcs_rx_data[43], w_hssi_10g_rx_pcs_rx_data[42], w_hssi_10g_rx_pcs_rx_data[41], w_hssi_10g_rx_pcs_rx_data[40], w_hssi_10g_rx_pcs_rx_data[39], w_hssi_10g_rx_pcs_rx_data[38], w_hssi_10g_rx_pcs_rx_data[37], w_hssi_10g_rx_pcs_rx_data[36], w_hssi_10g_rx_pcs_rx_data[35], w_hssi_10g_rx_pcs_rx_data[34], w_hssi_10g_rx_pcs_rx_data[33], w_hssi_10g_rx_pcs_rx_data[32], w_hssi_10g_rx_pcs_rx_data[31], w_hssi_10g_rx_pcs_rx_data[30], w_hssi_10g_rx_pcs_rx_data[29], w_hssi_10g_rx_pcs_rx_data[28], w_hssi_10g_rx_pcs_rx_data[27], w_hssi_10g_rx_pcs_rx_data[26], w_hssi_10g_rx_pcs_rx_data[25], w_hssi_10g_rx_pcs_rx_data[24], w_hssi_10g_rx_pcs_rx_data[23], w_hssi_10g_rx_pcs_rx_data[22], w_hssi_10g_rx_pcs_rx_data[21], w_hssi_10g_rx_pcs_rx_data[20], w_hssi_10g_rx_pcs_rx_data[19], w_hssi_10g_rx_pcs_rx_data[18], w_hssi_10g_rx_pcs_rx_data[17], w_hssi_10g_rx_pcs_rx_data[16], w_hssi_10g_rx_pcs_rx_data[15], w_hssi_10g_rx_pcs_rx_data[14], w_hssi_10g_rx_pcs_rx_data[13], w_hssi_10g_rx_pcs_rx_data[12], w_hssi_10g_rx_pcs_rx_data[11], w_hssi_10g_rx_pcs_rx_data[10], w_hssi_10g_rx_pcs_rx_data[9], w_hssi_10g_rx_pcs_rx_data[8], w_hssi_10g_rx_pcs_rx_data[7], w_hssi_10g_rx_pcs_rx_data[6], w_hssi_10g_rx_pcs_rx_data[5], w_hssi_10g_rx_pcs_rx_data[4], w_hssi_10g_rx_pcs_rx_data[3], w_hssi_10g_rx_pcs_rx_data[2], w_hssi_10g_rx_pcs_rx_data[1], w_hssi_10g_rx_pcs_rx_data[0]}),
				.int_pldif_10g_rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.int_pldif_10g_rx_diag_status({w_hssi_10g_rx_pcs_rx_diag_status[1], w_hssi_10g_rx_pcs_rx_diag_status[0]}),
				.int_pldif_10g_rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.int_pldif_10g_rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.int_pldif_10g_rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.int_pldif_10g_rx_fifo_num({w_hssi_10g_rx_pcs_rx_fifo_num[4], w_hssi_10g_rx_pcs_rx_fifo_num[3], w_hssi_10g_rx_pcs_rx_fifo_num[2], w_hssi_10g_rx_pcs_rx_fifo_num[1], w_hssi_10g_rx_pcs_rx_fifo_num[0]}),
				.int_pldif_10g_rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.int_pldif_10g_rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.int_pldif_10g_rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.int_pldif_10g_rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.int_pldif_10g_rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.int_pldif_10g_rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				.int_pldif_8g_a1a2_k1k2_flag({w_hssi_8g_rx_pcs_a1a2k1k2flag[3], w_hssi_8g_rx_pcs_a1a2k1k2flag[2], w_hssi_8g_rx_pcs_a1a2k1k2flag[1], w_hssi_8g_rx_pcs_a1a2k1k2flag[0]}),
				.int_pldif_8g_empty_rmf(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.int_pldif_8g_empty_rx(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.int_pldif_8g_full_rmf(w_hssi_8g_rx_pcs_rm_fifo_full),
				.int_pldif_8g_full_rx(w_hssi_8g_rx_pcs_pcfifofull),
				.int_pldif_8g_phystatus(w_hssi_8g_rx_pcs_phystatus),
				.int_pldif_8g_rx_blk_start({w_hssi_8g_rx_pcs_rx_blk_start[3], w_hssi_8g_rx_pcs_rx_blk_start[2], w_hssi_8g_rx_pcs_rx_blk_start[1], w_hssi_8g_rx_pcs_rx_blk_start[0]}),
				.int_pldif_8g_rx_clk(w_hssi_8g_rx_pcs_clock_to_pld),
				.int_pldif_8g_rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_8g_rx_data_valid({w_hssi_8g_rx_pcs_rx_data_valid[3], w_hssi_8g_rx_pcs_rx_data_valid[2], w_hssi_8g_rx_pcs_rx_data_valid[1], w_hssi_8g_rx_pcs_rx_data_valid[0]}),
				.int_pldif_8g_rx_rstn_sync2wrfifo(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.int_pldif_8g_rx_sync_hdr({w_hssi_8g_rx_pcs_rx_sync_hdr[1], w_hssi_8g_rx_pcs_rx_sync_hdr[0]}),
				.int_pldif_8g_rxd({w_hssi_8g_rx_pcs_dataout[63], w_hssi_8g_rx_pcs_dataout[62], w_hssi_8g_rx_pcs_dataout[61], w_hssi_8g_rx_pcs_dataout[60], w_hssi_8g_rx_pcs_dataout[59], w_hssi_8g_rx_pcs_dataout[58], w_hssi_8g_rx_pcs_dataout[57], w_hssi_8g_rx_pcs_dataout[56], w_hssi_8g_rx_pcs_dataout[55], w_hssi_8g_rx_pcs_dataout[54], w_hssi_8g_rx_pcs_dataout[53], w_hssi_8g_rx_pcs_dataout[52], w_hssi_8g_rx_pcs_dataout[51], w_hssi_8g_rx_pcs_dataout[50], w_hssi_8g_rx_pcs_dataout[49], w_hssi_8g_rx_pcs_dataout[48], w_hssi_8g_rx_pcs_dataout[47], w_hssi_8g_rx_pcs_dataout[46], w_hssi_8g_rx_pcs_dataout[45], w_hssi_8g_rx_pcs_dataout[44], w_hssi_8g_rx_pcs_dataout[43], w_hssi_8g_rx_pcs_dataout[42], w_hssi_8g_rx_pcs_dataout[41], w_hssi_8g_rx_pcs_dataout[40], w_hssi_8g_rx_pcs_dataout[39], w_hssi_8g_rx_pcs_dataout[38], w_hssi_8g_rx_pcs_dataout[37], w_hssi_8g_rx_pcs_dataout[36], w_hssi_8g_rx_pcs_dataout[35], w_hssi_8g_rx_pcs_dataout[34], w_hssi_8g_rx_pcs_dataout[33], w_hssi_8g_rx_pcs_dataout[32], w_hssi_8g_rx_pcs_dataout[31], w_hssi_8g_rx_pcs_dataout[30], w_hssi_8g_rx_pcs_dataout[29], w_hssi_8g_rx_pcs_dataout[28], w_hssi_8g_rx_pcs_dataout[27], w_hssi_8g_rx_pcs_dataout[26], w_hssi_8g_rx_pcs_dataout[25], w_hssi_8g_rx_pcs_dataout[24], w_hssi_8g_rx_pcs_dataout[23], w_hssi_8g_rx_pcs_dataout[22], w_hssi_8g_rx_pcs_dataout[21], w_hssi_8g_rx_pcs_dataout[20], w_hssi_8g_rx_pcs_dataout[19], w_hssi_8g_rx_pcs_dataout[18], w_hssi_8g_rx_pcs_dataout[17], w_hssi_8g_rx_pcs_dataout[16], w_hssi_8g_rx_pcs_dataout[15], w_hssi_8g_rx_pcs_dataout[14], w_hssi_8g_rx_pcs_dataout[13], w_hssi_8g_rx_pcs_dataout[12], w_hssi_8g_rx_pcs_dataout[11], w_hssi_8g_rx_pcs_dataout[10], w_hssi_8g_rx_pcs_dataout[9], w_hssi_8g_rx_pcs_dataout[8], w_hssi_8g_rx_pcs_dataout[7], w_hssi_8g_rx_pcs_dataout[6], w_hssi_8g_rx_pcs_dataout[5], w_hssi_8g_rx_pcs_dataout[4], w_hssi_8g_rx_pcs_dataout[3], w_hssi_8g_rx_pcs_dataout[2], w_hssi_8g_rx_pcs_dataout[1], w_hssi_8g_rx_pcs_dataout[0]}),
				.int_pldif_8g_rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.int_pldif_8g_rxstatus({w_hssi_8g_rx_pcs_rxstatus[2], w_hssi_8g_rx_pcs_rxstatus[1], w_hssi_8g_rx_pcs_rxstatus[0]}),
				.int_pldif_8g_rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.int_pldif_8g_signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.int_pldif_8g_wa_boundary({w_hssi_8g_rx_pcs_word_align_boundary[4], w_hssi_8g_rx_pcs_word_align_boundary[3], w_hssi_8g_rx_pcs_word_align_boundary[2], w_hssi_8g_rx_pcs_word_align_boundary[1], w_hssi_8g_rx_pcs_word_align_boundary[0]}),
				.int_pldif_krfec_rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.int_pldif_krfec_rx_data_status({w_hssi_krfec_rx_pcs_rx_data_status[1], w_hssi_krfec_rx_pcs_rx_data_status[0]}),
				.int_pldif_krfec_rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.int_pldif_pmaif_clkdiv_rx(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pldif_pmaif_clkdiv_rx_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pldif_pmaif_rx_data({w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0]}),
				.int_pldif_pmaif_rx_prbs_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pldif_pmaif_rx_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.pld_10g_krfec_rx_clr_errblk_cnt(in_pld_10g_krfec_rx_clr_errblk_cnt),
				.pld_10g_krfec_rx_pld_rst_n(in_pld_10g_krfec_rx_pld_rst_n),
				.pld_10g_rx_align_clr(in_pld_10g_rx_align_clr),
				.pld_10g_rx_clr_ber_count(in_pld_10g_rx_clr_ber_count),
				.pld_10g_rx_rd_en(in_pld_10g_rx_rd_en),
				.pld_8g_a1a2_size(in_pld_8g_a1a2_size),
				.pld_8g_bitloc_rev_en(in_pld_8g_bitloc_rev_en),
				.pld_8g_byte_rev_en(in_pld_8g_byte_rev_en),
				.pld_8g_encdt(in_pld_8g_encdt),
				.pld_8g_g3_rx_pld_rst_n(in_pld_8g_g3_rx_pld_rst_n),
				.pld_8g_rdenable_rx(in_pld_8g_rdenable_rx),
				.pld_8g_rxpolarity(in_pld_8g_rxpolarity),
				.pld_8g_wrdisable_rx(in_pld_8g_wrdisable_rx),
				.pld_bitslip(in_pld_bitslip),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_rxpma_rstb(in_pld_pma_rxpma_rstb),
				.pld_pmaif_rx_pld_rst_n(in_pld_pmaif_rx_pld_rst_n),
				.pld_pmaif_rxclkslip(in_pld_pmaif_rxclkslip),
				.pld_polinv_rx(in_pld_polinv_rx),
				.pld_rx_clk(in_pld_rx_clk),
				.pld_rx_prbs_err_clr(in_pld_rx_prbs_err_clr),
				.pld_syncsm_en(in_pld_syncsm_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.int_pldif_pmaif_rx_pld_clk(),
				.pld_8g_wa_boundary_txclk_fastreg(),
				.pld_8g_wa_boundary_txclk_reg(),
				.pld_bitslip_10g_txclk_reg(),
				.pld_bitslip_8g_txclk_reg(),
				.pld_bitslip_rxclk_parallel_loopback_reg(),
				.pld_bitslip_rxclk_reg(),
				.pld_pcs_rx_clk_out_pcsdirect_wire(),
				.pld_pma_rx_clk_out_10g_or_pcsdirect_wire(),
				.pld_pma_rx_clk_out_8g_wire(),
				.pld_pmaif_rx_pld_rst_n_reg(),
				.pld_pmaif_tx_pld_rst_n_txclk_reg(),
				.pld_polinv_rx_reg(),
				.pld_rx_clk_fifo(),
				.pld_rx_control_fifo(),
				.pld_rx_control_pcsdirect_reg(),
				.pld_rx_data_fifo(),
				.pld_rx_data_pcsdirect_reg(),
				.pld_rx_prbs_done_reg(),
				.pld_rx_prbs_done_txclk_reg(),
				.pld_rx_prbs_err_clr_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_clr_reg(),
				.pld_rx_prbs_err_disprbs_reg(),
				.pld_rx_prbs_err_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_reg(),
				.pma_rx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_data[50:0] = 51'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3:0] = 4'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_control[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_data[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pcs_pma_interface
			twentynm_hssi_tx_pcs_pma_interface #(
				.bypass_pma_txelecidle(hssi_tx_pcs_pma_interface_bypass_pma_txelecidle),
				.channel_operation_mode(hssi_tx_pcs_pma_interface_channel_operation_mode),
				.lpbk_en(hssi_tx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_tx_pcs_pma_interface_master_clk_sel),
				.pcie_sub_prot_mode_tx(hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx),
				.pldif_datawidth_mode(hssi_tx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_tx(hssi_tx_pcs_pma_interface_pma_dw_tx),
				.pma_if_dft_en(hssi_tx_pcs_pma_interface_pma_if_dft_en),
				.pmagate_en(hssi_tx_pcs_pma_interface_pmagate_en),
				.prbs9_dwidth(hssi_tx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_tx_pcs_pma_interface_prbs_clken),
				.prbs_gen_pat(hssi_tx_pcs_pma_interface_prbs_gen_pat),
				.prot_mode_tx(hssi_tx_pcs_pma_interface_prot_mode_tx),
				.reconfig_settings(hssi_tx_pcs_pma_interface_reconfig_settings),
				.silicon_rev( "20nm1" ),       //PARAM_HIDE
				.sq_wave_num(hssi_tx_pcs_pma_interface_sq_wave_num),
				.sqwgen_clken(hssi_tx_pcs_pma_interface_sqwgen_clken),
				.sup_mode(hssi_tx_pcs_pma_interface_sup_mode),
				.tx_dyn_polarity_inversion(hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion),
				.tx_pma_data_sel(hssi_tx_pcs_pma_interface_tx_pma_data_sel),
				.tx_static_polarity_inversion(hssi_tx_pcs_pma_interface_tx_static_polarity_inversion),
				.uhsif_cnt_step_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock),
				.uhsif_cnt_thresh_filt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value),
				.uhsif_cnt_thresh_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock),
				.uhsif_dcn_test_update_period(hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period),
				.uhsif_dcn_testmode_enable(hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable),
				.uhsif_dead_zone_count_thresh(hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh),
				.uhsif_dead_zone_detection_enable(hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable),
				.uhsif_dead_zone_obser_window(hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window),
				.uhsif_dead_zone_skip_size(hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size),
				.uhsif_delay_cell_index_sel(hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel),
				.uhsif_delay_cell_margin(hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin),
				.uhsif_delay_cell_static_index_value(hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value),
				.uhsif_dft_dead_zone_control(hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control),
				.uhsif_dft_up_filt_control(hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control),
				.uhsif_enable(hssi_tx_pcs_pma_interface_uhsif_enable),
				.uhsif_lock_det_segsz_after_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock),
				.uhsif_lock_det_segsz_before_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock),
				.uhsif_lock_det_thresh_cnt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value),
				.uhsif_lock_det_thresh_cnt_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value),
				.uhsif_lock_det_thresh_diff_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value),
				.uhsif_lock_det_thresh_diff_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value)
			) inst_twentynm_hssi_tx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.int_pmaif_8g_txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.int_pmaif_pldif_tx_clkdiv(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pmaif_pldif_tx_clkdiv_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pmaif_pldif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.int_pmaif_pldif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.int_tx_dft_obsrv_clk(w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk),
				.pma_tx_elec_idle(w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle),
				.pma_tx_pma_data(w_hssi_tx_pcs_pma_interface_pma_tx_pma_data),
				.pma_txpma_rstb(w_hssi_tx_pcs_pma_interface_pma_txpma_rstb),
				.tx_pma_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback),
				.tx_pma_uhsif_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback),
				.tx_prbs_gen_test(w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test),
				.uhsif_test_out_1(w_hssi_tx_pcs_pma_interface_uhsif_test_out_1),
				.uhsif_test_out_2(w_hssi_tx_pcs_pma_interface_uhsif_test_out_2),
				.uhsif_test_out_3(w_hssi_tx_pcs_pma_interface_uhsif_test_out_3),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.int_pmaif_10g_tx_pma_data({w_hssi_10g_tx_pcs_tx_pma_data[63], w_hssi_10g_tx_pcs_tx_pma_data[62], w_hssi_10g_tx_pcs_tx_pma_data[61], w_hssi_10g_tx_pcs_tx_pma_data[60], w_hssi_10g_tx_pcs_tx_pma_data[59], w_hssi_10g_tx_pcs_tx_pma_data[58], w_hssi_10g_tx_pcs_tx_pma_data[57], w_hssi_10g_tx_pcs_tx_pma_data[56], w_hssi_10g_tx_pcs_tx_pma_data[55], w_hssi_10g_tx_pcs_tx_pma_data[54], w_hssi_10g_tx_pcs_tx_pma_data[53], w_hssi_10g_tx_pcs_tx_pma_data[52], w_hssi_10g_tx_pcs_tx_pma_data[51], w_hssi_10g_tx_pcs_tx_pma_data[50], w_hssi_10g_tx_pcs_tx_pma_data[49], w_hssi_10g_tx_pcs_tx_pma_data[48], w_hssi_10g_tx_pcs_tx_pma_data[47], w_hssi_10g_tx_pcs_tx_pma_data[46], w_hssi_10g_tx_pcs_tx_pma_data[45], w_hssi_10g_tx_pcs_tx_pma_data[44], w_hssi_10g_tx_pcs_tx_pma_data[43], w_hssi_10g_tx_pcs_tx_pma_data[42], w_hssi_10g_tx_pcs_tx_pma_data[41], w_hssi_10g_tx_pcs_tx_pma_data[40], w_hssi_10g_tx_pcs_tx_pma_data[39], w_hssi_10g_tx_pcs_tx_pma_data[38], w_hssi_10g_tx_pcs_tx_pma_data[37], w_hssi_10g_tx_pcs_tx_pma_data[36], w_hssi_10g_tx_pcs_tx_pma_data[35], w_hssi_10g_tx_pcs_tx_pma_data[34], w_hssi_10g_tx_pcs_tx_pma_data[33], w_hssi_10g_tx_pcs_tx_pma_data[32], w_hssi_10g_tx_pcs_tx_pma_data[31], w_hssi_10g_tx_pcs_tx_pma_data[30], w_hssi_10g_tx_pcs_tx_pma_data[29], w_hssi_10g_tx_pcs_tx_pma_data[28], w_hssi_10g_tx_pcs_tx_pma_data[27], w_hssi_10g_tx_pcs_tx_pma_data[26], w_hssi_10g_tx_pcs_tx_pma_data[25], w_hssi_10g_tx_pcs_tx_pma_data[24], w_hssi_10g_tx_pcs_tx_pma_data[23], w_hssi_10g_tx_pcs_tx_pma_data[22], w_hssi_10g_tx_pcs_tx_pma_data[21], w_hssi_10g_tx_pcs_tx_pma_data[20], w_hssi_10g_tx_pcs_tx_pma_data[19], w_hssi_10g_tx_pcs_tx_pma_data[18], w_hssi_10g_tx_pcs_tx_pma_data[17], w_hssi_10g_tx_pcs_tx_pma_data[16], w_hssi_10g_tx_pcs_tx_pma_data[15], w_hssi_10g_tx_pcs_tx_pma_data[14], w_hssi_10g_tx_pcs_tx_pma_data[13], w_hssi_10g_tx_pcs_tx_pma_data[12], w_hssi_10g_tx_pcs_tx_pma_data[11], w_hssi_10g_tx_pcs_tx_pma_data[10], w_hssi_10g_tx_pcs_tx_pma_data[9], w_hssi_10g_tx_pcs_tx_pma_data[8], w_hssi_10g_tx_pcs_tx_pma_data[7], w_hssi_10g_tx_pcs_tx_pma_data[6], w_hssi_10g_tx_pcs_tx_pma_data[5], w_hssi_10g_tx_pcs_tx_pma_data[4], w_hssi_10g_tx_pcs_tx_pma_data[3], w_hssi_10g_tx_pcs_tx_pma_data[2], w_hssi_10g_tx_pcs_tx_pma_data[1], w_hssi_10g_tx_pcs_tx_pma_data[0]}),
				.int_pmaif_10g_tx_pma_data_gate_val({w_hssi_10g_tx_pcs_tx_pma_gating_val[63], w_hssi_10g_tx_pcs_tx_pma_gating_val[62], w_hssi_10g_tx_pcs_tx_pma_gating_val[61], w_hssi_10g_tx_pcs_tx_pma_gating_val[60], w_hssi_10g_tx_pcs_tx_pma_gating_val[59], w_hssi_10g_tx_pcs_tx_pma_gating_val[58], w_hssi_10g_tx_pcs_tx_pma_gating_val[57], w_hssi_10g_tx_pcs_tx_pma_gating_val[56], w_hssi_10g_tx_pcs_tx_pma_gating_val[55], w_hssi_10g_tx_pcs_tx_pma_gating_val[54], w_hssi_10g_tx_pcs_tx_pma_gating_val[53], w_hssi_10g_tx_pcs_tx_pma_gating_val[52], w_hssi_10g_tx_pcs_tx_pma_gating_val[51], w_hssi_10g_tx_pcs_tx_pma_gating_val[50], w_hssi_10g_tx_pcs_tx_pma_gating_val[49], w_hssi_10g_tx_pcs_tx_pma_gating_val[48], w_hssi_10g_tx_pcs_tx_pma_gating_val[47], w_hssi_10g_tx_pcs_tx_pma_gating_val[46], w_hssi_10g_tx_pcs_tx_pma_gating_val[45], w_hssi_10g_tx_pcs_tx_pma_gating_val[44], w_hssi_10g_tx_pcs_tx_pma_gating_val[43], w_hssi_10g_tx_pcs_tx_pma_gating_val[42], w_hssi_10g_tx_pcs_tx_pma_gating_val[41], w_hssi_10g_tx_pcs_tx_pma_gating_val[40], w_hssi_10g_tx_pcs_tx_pma_gating_val[39], w_hssi_10g_tx_pcs_tx_pma_gating_val[38], w_hssi_10g_tx_pcs_tx_pma_gating_val[37], w_hssi_10g_tx_pcs_tx_pma_gating_val[36], w_hssi_10g_tx_pcs_tx_pma_gating_val[35], w_hssi_10g_tx_pcs_tx_pma_gating_val[34], w_hssi_10g_tx_pcs_tx_pma_gating_val[33], w_hssi_10g_tx_pcs_tx_pma_gating_val[32], w_hssi_10g_tx_pcs_tx_pma_gating_val[31], w_hssi_10g_tx_pcs_tx_pma_gating_val[30], w_hssi_10g_tx_pcs_tx_pma_gating_val[29], w_hssi_10g_tx_pcs_tx_pma_gating_val[28], w_hssi_10g_tx_pcs_tx_pma_gating_val[27], w_hssi_10g_tx_pcs_tx_pma_gating_val[26], w_hssi_10g_tx_pcs_tx_pma_gating_val[25], w_hssi_10g_tx_pcs_tx_pma_gating_val[24], w_hssi_10g_tx_pcs_tx_pma_gating_val[23], w_hssi_10g_tx_pcs_tx_pma_gating_val[22], w_hssi_10g_tx_pcs_tx_pma_gating_val[21], w_hssi_10g_tx_pcs_tx_pma_gating_val[20], w_hssi_10g_tx_pcs_tx_pma_gating_val[19], w_hssi_10g_tx_pcs_tx_pma_gating_val[18], w_hssi_10g_tx_pcs_tx_pma_gating_val[17], w_hssi_10g_tx_pcs_tx_pma_gating_val[16], w_hssi_10g_tx_pcs_tx_pma_gating_val[15], w_hssi_10g_tx_pcs_tx_pma_gating_val[14], w_hssi_10g_tx_pcs_tx_pma_gating_val[13], w_hssi_10g_tx_pcs_tx_pma_gating_val[12], w_hssi_10g_tx_pcs_tx_pma_gating_val[11], w_hssi_10g_tx_pcs_tx_pma_gating_val[10], w_hssi_10g_tx_pcs_tx_pma_gating_val[9], w_hssi_10g_tx_pcs_tx_pma_gating_val[8], w_hssi_10g_tx_pcs_tx_pma_gating_val[7], w_hssi_10g_tx_pcs_tx_pma_gating_val[6], w_hssi_10g_tx_pcs_tx_pma_gating_val[5], w_hssi_10g_tx_pcs_tx_pma_gating_val[4], w_hssi_10g_tx_pcs_tx_pma_gating_val[3], w_hssi_10g_tx_pcs_tx_pma_gating_val[2], w_hssi_10g_tx_pcs_tx_pma_gating_val[1], w_hssi_10g_tx_pcs_tx_pma_gating_val[0]}),
				.int_pmaif_8g_pudr({w_hssi_8g_tx_pcs_dataout[19], w_hssi_8g_tx_pcs_dataout[18], w_hssi_8g_tx_pcs_dataout[17], w_hssi_8g_tx_pcs_dataout[16], w_hssi_8g_tx_pcs_dataout[15], w_hssi_8g_tx_pcs_dataout[14], w_hssi_8g_tx_pcs_dataout[13], w_hssi_8g_tx_pcs_dataout[12], w_hssi_8g_tx_pcs_dataout[11], w_hssi_8g_tx_pcs_dataout[10], w_hssi_8g_tx_pcs_dataout[9], w_hssi_8g_tx_pcs_dataout[8], w_hssi_8g_tx_pcs_dataout[7], w_hssi_8g_tx_pcs_dataout[6], w_hssi_8g_tx_pcs_dataout[5], w_hssi_8g_tx_pcs_dataout[4], w_hssi_8g_tx_pcs_dataout[3], w_hssi_8g_tx_pcs_dataout[2], w_hssi_8g_tx_pcs_dataout[1], w_hssi_8g_tx_pcs_dataout[0]}),
				.int_pmaif_8g_tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.int_pmaif_8g_tx_elec_idle(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_pma_data_out({w_hssi_gen3_tx_pcs_data_out[31], w_hssi_gen3_tx_pcs_data_out[30], w_hssi_gen3_tx_pcs_data_out[29], w_hssi_gen3_tx_pcs_data_out[28], w_hssi_gen3_tx_pcs_data_out[27], w_hssi_gen3_tx_pcs_data_out[26], w_hssi_gen3_tx_pcs_data_out[25], w_hssi_gen3_tx_pcs_data_out[24], w_hssi_gen3_tx_pcs_data_out[23], w_hssi_gen3_tx_pcs_data_out[22], w_hssi_gen3_tx_pcs_data_out[21], w_hssi_gen3_tx_pcs_data_out[20], w_hssi_gen3_tx_pcs_data_out[19], w_hssi_gen3_tx_pcs_data_out[18], w_hssi_gen3_tx_pcs_data_out[17], w_hssi_gen3_tx_pcs_data_out[16], w_hssi_gen3_tx_pcs_data_out[15], w_hssi_gen3_tx_pcs_data_out[14], w_hssi_gen3_tx_pcs_data_out[13], w_hssi_gen3_tx_pcs_data_out[12], w_hssi_gen3_tx_pcs_data_out[11], w_hssi_gen3_tx_pcs_data_out[10], w_hssi_gen3_tx_pcs_data_out[9], w_hssi_gen3_tx_pcs_data_out[8], w_hssi_gen3_tx_pcs_data_out[7], w_hssi_gen3_tx_pcs_data_out[6], w_hssi_gen3_tx_pcs_data_out[5], w_hssi_gen3_tx_pcs_data_out[4], w_hssi_gen3_tx_pcs_data_out[3], w_hssi_gen3_tx_pcs_data_out[2], w_hssi_gen3_tx_pcs_data_out[1], w_hssi_gen3_tx_pcs_data_out[0]}),
				.int_pmaif_g3_pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.int_pmaif_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pmaif_pldif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pmaif_pldif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0]}),
				.int_pmaif_pldif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pmaif_pldif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.int_pmaif_pldif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pmaif_pldif_uhsif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0]}),
				.pma_tx_clkdiv_user(in_pma_tx_clkdiv_user),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.refclk_dig_uhsif(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.uhsif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.uhsif_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				
				// UNUSED
				.avmm_user_dataout(),
				.write_en(),
				.write_en_ack()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4:0] = 5'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_txpma_rstb = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pld_pcs_interface
			twentynm_hssi_tx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx),
				.hd_10g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx),
				.hd_10g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx),
				.hd_10g_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx),
				.hd_10g_lpbk_en(hssi_tx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx),
				.hd_10g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx),
				.hd_10g_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx),
				.hd_8g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx),
				.hd_8g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx),
				.hd_8g_hip_mode(hssi_tx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_tx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx),
				.hd_8g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx),
				.hd_chnl_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx),
				.hd_chnl_frequency_rules_en(hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_tx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_tx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx),
				.hd_chnl_lpbk_en(hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx),
				.hd_chnl_pld_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz),
				.hd_chnl_pld_uhsif_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz),
				.hd_chnl_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx),
				.hd_chnl_pma_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz),
				.hd_chnl_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx),
				.hd_chnl_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx),
				.hd_fifo_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx),
				.hd_fifo_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx),
				.hd_g3_prot_mode(hssi_tx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx),
				.hd_krfec_lpbk_en(hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx),
				.hd_pldif_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx),
				.hd_pmaif_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_ctrl_plane_bonding(hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding),
				.hd_pmaif_lpbk_en(hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx),
				.hd_pmaif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx),
				.hd_pmaif_sim_mode(hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_tx_clk_out_sel(hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel),
				.pcs_tx_clk_source(hssi_tx_pld_pcs_interface_pcs_tx_clk_source),
				.pcs_tx_data_source(hssi_tx_pld_pcs_interface_pcs_tx_data_source),
				.pcs_tx_delay1_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en),
				.pcs_tx_delay1_clk_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel),
				.pcs_tx_delay1_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl),
				.pcs_tx_delay1_data_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel),
				.pcs_tx_delay2_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en),
				.pcs_tx_delay2_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl),
				.pcs_tx_output_sel(hssi_tx_pld_pcs_interface_pcs_tx_output_sel),
				.reconfig_settings(hssi_tx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm1" )       //PARAM_HIDE
			) inst_twentynm_hssi_tx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pld_pcs_interface_blockselect),
				.hip_tx_clk(w_hssi_tx_pld_pcs_interface_hip_tx_clk),
				.int_pldif_10g_tx_bitslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip),
				.int_pldif_10g_tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.int_pldif_10g_tx_control(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control),
				.int_pldif_10g_tx_control_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg),
				.int_pldif_10g_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data),
				.int_pldif_10g_tx_data_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg),
				.int_pldif_10g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.int_pldif_10g_tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.int_pldif_10g_tx_diag_status(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status),
				.int_pldif_10g_tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.int_pldif_10g_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.int_pldif_10g_tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				.int_pldif_8g_pld_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.int_pldif_8g_powerdown(w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown),
				.int_pldif_8g_rddisable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.int_pldif_8g_rev_loopbk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.int_pldif_8g_tx_blk_start(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start),
				.int_pldif_8g_tx_boundary_sel(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel),
				.int_pldif_8g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid),
				.int_pldif_8g_tx_sync_hdr(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr),
				.int_pldif_8g_txd(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd),
				.int_pldif_8g_txd_fast_reg(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg),
				.int_pldif_8g_txdeemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.int_pldif_8g_txdetectrxloopback(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.int_pldif_8g_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.int_pldif_8g_txmargin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin),
				.int_pldif_8g_txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.int_pldif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.int_pldif_8g_wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				.int_pldif_pmaif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pldif_pmaif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pldif_pmaif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data),
				.int_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pldif_pmaif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pldif_pmaif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pldif_pmaif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pldif_pmaif_uhsif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data),
				.pld_10g_krfec_tx_frame(w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame),
				.pld_10g_tx_burst_en_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe),
				.pld_10g_tx_empty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty),
				.pld_10g_tx_fifo_num(w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num),
				.pld_10g_tx_full(w_hssi_tx_pld_pcs_interface_pld_10g_tx_full),
				.pld_10g_tx_pempty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty),
				.pld_10g_tx_pfull(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull),
				.pld_10g_tx_wordslip_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe),
				.pld_8g_empty_tx(w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx),
				.pld_8g_full_tx(w_hssi_tx_pld_pcs_interface_pld_8g_full_tx),
				.pld_krfec_tx_alignment(w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment),
				.pld_pcs_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out),
				.pld_pma_clkdiv_tx_user(w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user),
				.pld_pma_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out),
				.pld_uhsif_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.hip_tx_data({in_hip_tx_data[63], in_hip_tx_data[62], in_hip_tx_data[61], in_hip_tx_data[60], in_hip_tx_data[59], in_hip_tx_data[58], in_hip_tx_data[57], in_hip_tx_data[56], in_hip_tx_data[55], in_hip_tx_data[54], in_hip_tx_data[53], in_hip_tx_data[52], in_hip_tx_data[51], in_hip_tx_data[50], in_hip_tx_data[49], in_hip_tx_data[48], in_hip_tx_data[47], in_hip_tx_data[46], in_hip_tx_data[45], in_hip_tx_data[44], in_hip_tx_data[43], in_hip_tx_data[42], in_hip_tx_data[41], in_hip_tx_data[40], in_hip_tx_data[39], in_hip_tx_data[38], in_hip_tx_data[37], in_hip_tx_data[36], in_hip_tx_data[35], in_hip_tx_data[34], in_hip_tx_data[33], in_hip_tx_data[32], in_hip_tx_data[31], in_hip_tx_data[30], in_hip_tx_data[29], in_hip_tx_data[28], in_hip_tx_data[27], in_hip_tx_data[26], in_hip_tx_data[25], in_hip_tx_data[24], in_hip_tx_data[23], in_hip_tx_data[22], in_hip_tx_data[21], in_hip_tx_data[20], in_hip_tx_data[19], in_hip_tx_data[18], in_hip_tx_data[17], in_hip_tx_data[16], in_hip_tx_data[15], in_hip_tx_data[14], in_hip_tx_data[13], in_hip_tx_data[12], in_hip_tx_data[11], in_hip_tx_data[10], in_hip_tx_data[9], in_hip_tx_data[8], in_hip_tx_data[7], in_hip_tx_data[6], in_hip_tx_data[5], in_hip_tx_data[4], in_hip_tx_data[3], in_hip_tx_data[2], in_hip_tx_data[1], in_hip_tx_data[0]}),
				.int_pldif_10g_tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.int_pldif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.int_pldif_10g_tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_10g_tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.int_pldif_10g_tx_fifo_num({w_hssi_10g_tx_pcs_tx_fifo_num[3], w_hssi_10g_tx_pcs_tx_fifo_num[2], w_hssi_10g_tx_pcs_tx_fifo_num[1], w_hssi_10g_tx_pcs_tx_fifo_num[0]}),
				.int_pldif_10g_tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.int_pldif_10g_tx_full(w_hssi_10g_tx_pcs_tx_full),
				.int_pldif_10g_tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.int_pldif_10g_tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.int_pldif_10g_tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				.int_pldif_8g_empty_tx(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.int_pldif_8g_full_tx(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.int_pldif_8g_tx_clk_out(w_hssi_8g_tx_pcs_clk_out),
				.int_pldif_8g_tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_krfec_tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.int_pldif_krfec_tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.int_pldif_pmaif_clkdiv_tx(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pldif_pmaif_clkdiv_tx_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pldif_pmaif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.pld_10g_krfec_tx_pld_rst_n(in_pld_10g_krfec_tx_pld_rst_n),
				.pld_10g_tx_bitslip({in_pld_10g_tx_bitslip[6], in_pld_10g_tx_bitslip[5], in_pld_10g_tx_bitslip[4], in_pld_10g_tx_bitslip[3], in_pld_10g_tx_bitslip[2], in_pld_10g_tx_bitslip[1], in_pld_10g_tx_bitslip[0]}),
				.pld_10g_tx_burst_en(in_pld_10g_tx_burst_en),
				.pld_10g_tx_data_valid(in_pld_10g_tx_data_valid),
				.pld_10g_tx_diag_status({in_pld_10g_tx_diag_status[1], in_pld_10g_tx_diag_status[0]}),
				.pld_10g_tx_wordslip(in_pld_10g_tx_wordslip),
				.pld_8g_g3_tx_pld_rst_n(in_pld_8g_g3_tx_pld_rst_n),
				.pld_8g_rddisable_tx(in_pld_8g_rddisable_tx),
				.pld_8g_tx_boundary_sel({in_pld_8g_tx_boundary_sel[4], in_pld_8g_tx_boundary_sel[3], in_pld_8g_tx_boundary_sel[2], in_pld_8g_tx_boundary_sel[1], in_pld_8g_tx_boundary_sel[0]}),
				.pld_8g_wrenable_tx(in_pld_8g_wrenable_tx),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_txpma_rstb(in_pld_pma_txpma_rstb),
				.pld_pmaif_tx_pld_rst_n(in_pld_pmaif_tx_pld_rst_n),
				.pld_polinv_tx(in_pld_polinv_tx),
				.pld_tx_clk(in_pld_tx_clk),
				.pld_tx_control({in_pld_tx_control[17], in_pld_tx_control[16], in_pld_tx_control[15], in_pld_tx_control[14], in_pld_tx_control[13], in_pld_tx_control[12], in_pld_tx_control[11], in_pld_tx_control[10], in_pld_tx_control[9], in_pld_tx_control[8], in_pld_tx_control[7], in_pld_tx_control[6], in_pld_tx_control[5], in_pld_tx_control[4], in_pld_tx_control[3], in_pld_tx_control[2], in_pld_tx_control[1], in_pld_tx_control[0]}),
				.pld_tx_data({in_pld_tx_data[127], in_pld_tx_data[126], in_pld_tx_data[125], in_pld_tx_data[124], in_pld_tx_data[123], in_pld_tx_data[122], in_pld_tx_data[121], in_pld_tx_data[120], in_pld_tx_data[119], in_pld_tx_data[118], in_pld_tx_data[117], in_pld_tx_data[116], in_pld_tx_data[115], in_pld_tx_data[114], in_pld_tx_data[113], in_pld_tx_data[112], in_pld_tx_data[111], in_pld_tx_data[110], in_pld_tx_data[109], in_pld_tx_data[108], in_pld_tx_data[107], in_pld_tx_data[106], in_pld_tx_data[105], in_pld_tx_data[104], in_pld_tx_data[103], in_pld_tx_data[102], in_pld_tx_data[101], in_pld_tx_data[100], in_pld_tx_data[99], in_pld_tx_data[98], in_pld_tx_data[97], in_pld_tx_data[96], in_pld_tx_data[95], in_pld_tx_data[94], in_pld_tx_data[93], in_pld_tx_data[92], in_pld_tx_data[91], in_pld_tx_data[90], in_pld_tx_data[89], in_pld_tx_data[88], in_pld_tx_data[87], in_pld_tx_data[86], in_pld_tx_data[85], in_pld_tx_data[84], in_pld_tx_data[83], in_pld_tx_data[82], in_pld_tx_data[81], in_pld_tx_data[80], in_pld_tx_data[79], in_pld_tx_data[78], in_pld_tx_data[77], in_pld_tx_data[76], in_pld_tx_data[75], in_pld_tx_data[74], in_pld_tx_data[73], in_pld_tx_data[72], in_pld_tx_data[71], in_pld_tx_data[70], in_pld_tx_data[69], in_pld_tx_data[68], in_pld_tx_data[67], in_pld_tx_data[66], in_pld_tx_data[65], in_pld_tx_data[64], in_pld_tx_data[63], in_pld_tx_data[62], in_pld_tx_data[61], in_pld_tx_data[60], in_pld_tx_data[59], in_pld_tx_data[58], in_pld_tx_data[57], in_pld_tx_data[56], in_pld_tx_data[55], in_pld_tx_data[54], in_pld_tx_data[53], in_pld_tx_data[52], in_pld_tx_data[51], in_pld_tx_data[50], in_pld_tx_data[49], in_pld_tx_data[48], in_pld_tx_data[47], in_pld_tx_data[46], in_pld_tx_data[45], in_pld_tx_data[44], in_pld_tx_data[43], in_pld_tx_data[42], in_pld_tx_data[41], in_pld_tx_data[40], in_pld_tx_data[39], in_pld_tx_data[38], in_pld_tx_data[37], in_pld_tx_data[36], in_pld_tx_data[35], in_pld_tx_data[34], in_pld_tx_data[33], in_pld_tx_data[32], in_pld_tx_data[31], in_pld_tx_data[30], in_pld_tx_data[29], in_pld_tx_data[28], in_pld_tx_data[27], in_pld_tx_data[26], in_pld_tx_data[25], in_pld_tx_data[24], in_pld_tx_data[23], in_pld_tx_data[22], in_pld_tx_data[21], in_pld_tx_data[20], in_pld_tx_data[19], in_pld_tx_data[18], in_pld_tx_data[17], in_pld_tx_data[16], in_pld_tx_data[15], in_pld_tx_data[14], in_pld_tx_data[13], in_pld_tx_data[12], in_pld_tx_data[11], in_pld_tx_data[10], in_pld_tx_data[9], in_pld_tx_data[8], in_pld_tx_data[7], in_pld_tx_data[6], in_pld_tx_data[5], in_pld_tx_data[4], in_pld_tx_data[3], in_pld_tx_data[2], in_pld_tx_data[1], in_pld_tx_data[0]}),
				.pld_txelecidle(in_pld_txelecidle),
				.pld_uhsif_tx_clk(in_pld_uhsif_tx_clk),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.hip_clk_out_div_by_2_wire(),
				.hip_clk_out_wire(),
				.int_pldif_pmaif_tx_pld_clk(),
				.pld_10g_tx_burst_en_exe_10g_fastreg(),
				.pld_10g_tx_burst_en_exe_plddirect_reg(),
				.pld_10g_tx_data_valid_2ff_delay1_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay3_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg(),
				.pld_10g_tx_data_valid_fastreg(),
				.pld_10g_tx_data_valid_plddirect_fastreg(),
				.pld_pcs_tx_clk_out_pma_wire(),
				.pld_pma_tx_clk_out_wire(),
				.pld_pmaif_tx_pld_rst_n_reg(),
				.pld_polinv_tx_10g_pcsdirect_reg(),
				.pld_polinv_tx_8g_reg(),
				.pld_polinv_tx_pat_reg(),
				.pld_tx_clk_fifo(),
				.pld_tx_control_fifo(),
				.pld_tx_control_hi_10g_reg(),
				.pld_tx_control_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_10g_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_8g_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_control_lo_plddirect_fastreg(),
				.pld_tx_control_lo_plddirect_reg(),
				.pld_tx_data_hi_reg(),
				.pld_tx_data_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_10g_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_8g_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_data_lo_plddirect_fastreg(),
				.pld_tx_data_lo_plddirect_reg(),
				.pld_uhsif_reg(),
				.pma_tx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_hip_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6:0] = 7'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17:0] = 18'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8:0] = 9'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127:0] = 128'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4:0] = 5'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2:0] = 3'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_full = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_full_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out = 1'b0;
		end // if not generate
		
		//output assignments
		assign out_avmmreaddata_hssi_10g_rx_pcs = {w_hssi_10g_rx_pcs_avmmreaddata[7], w_hssi_10g_rx_pcs_avmmreaddata[6], w_hssi_10g_rx_pcs_avmmreaddata[5], w_hssi_10g_rx_pcs_avmmreaddata[4], w_hssi_10g_rx_pcs_avmmreaddata[3], w_hssi_10g_rx_pcs_avmmreaddata[2], w_hssi_10g_rx_pcs_avmmreaddata[1], w_hssi_10g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_10g_tx_pcs = {w_hssi_10g_tx_pcs_avmmreaddata[7], w_hssi_10g_tx_pcs_avmmreaddata[6], w_hssi_10g_tx_pcs_avmmreaddata[5], w_hssi_10g_tx_pcs_avmmreaddata[4], w_hssi_10g_tx_pcs_avmmreaddata[3], w_hssi_10g_tx_pcs_avmmreaddata[2], w_hssi_10g_tx_pcs_avmmreaddata[1], w_hssi_10g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_rx_pcs = {w_hssi_8g_rx_pcs_avmmreaddata[7], w_hssi_8g_rx_pcs_avmmreaddata[6], w_hssi_8g_rx_pcs_avmmreaddata[5], w_hssi_8g_rx_pcs_avmmreaddata[4], w_hssi_8g_rx_pcs_avmmreaddata[3], w_hssi_8g_rx_pcs_avmmreaddata[2], w_hssi_8g_rx_pcs_avmmreaddata[1], w_hssi_8g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_tx_pcs = {w_hssi_8g_tx_pcs_avmmreaddata[7], w_hssi_8g_tx_pcs_avmmreaddata[6], w_hssi_8g_tx_pcs_avmmreaddata[5], w_hssi_8g_tx_pcs_avmmreaddata[4], w_hssi_8g_tx_pcs_avmmreaddata[3], w_hssi_8g_tx_pcs_avmmreaddata[2], w_hssi_8g_tx_pcs_avmmreaddata[1], w_hssi_8g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pcs_pma_interface = {w_hssi_common_pcs_pma_interface_avmmreaddata[7], w_hssi_common_pcs_pma_interface_avmmreaddata[6], w_hssi_common_pcs_pma_interface_avmmreaddata[5], w_hssi_common_pcs_pma_interface_avmmreaddata[4], w_hssi_common_pcs_pma_interface_avmmreaddata[3], w_hssi_common_pcs_pma_interface_avmmreaddata[2], w_hssi_common_pcs_pma_interface_avmmreaddata[1], w_hssi_common_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pld_pcs_interface = {w_hssi_common_pld_pcs_interface_avmmreaddata[7], w_hssi_common_pld_pcs_interface_avmmreaddata[6], w_hssi_common_pld_pcs_interface_avmmreaddata[5], w_hssi_common_pld_pcs_interface_avmmreaddata[4], w_hssi_common_pld_pcs_interface_avmmreaddata[3], w_hssi_common_pld_pcs_interface_avmmreaddata[2], w_hssi_common_pld_pcs_interface_avmmreaddata[1], w_hssi_common_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_rx_pcs = {w_hssi_fifo_rx_pcs_avmmreaddata[7], w_hssi_fifo_rx_pcs_avmmreaddata[6], w_hssi_fifo_rx_pcs_avmmreaddata[5], w_hssi_fifo_rx_pcs_avmmreaddata[4], w_hssi_fifo_rx_pcs_avmmreaddata[3], w_hssi_fifo_rx_pcs_avmmreaddata[2], w_hssi_fifo_rx_pcs_avmmreaddata[1], w_hssi_fifo_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_tx_pcs = {w_hssi_fifo_tx_pcs_avmmreaddata[7], w_hssi_fifo_tx_pcs_avmmreaddata[6], w_hssi_fifo_tx_pcs_avmmreaddata[5], w_hssi_fifo_tx_pcs_avmmreaddata[4], w_hssi_fifo_tx_pcs_avmmreaddata[3], w_hssi_fifo_tx_pcs_avmmreaddata[2], w_hssi_fifo_tx_pcs_avmmreaddata[1], w_hssi_fifo_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_rx_pcs = {w_hssi_gen3_rx_pcs_avmmreaddata[7], w_hssi_gen3_rx_pcs_avmmreaddata[6], w_hssi_gen3_rx_pcs_avmmreaddata[5], w_hssi_gen3_rx_pcs_avmmreaddata[4], w_hssi_gen3_rx_pcs_avmmreaddata[3], w_hssi_gen3_rx_pcs_avmmreaddata[2], w_hssi_gen3_rx_pcs_avmmreaddata[1], w_hssi_gen3_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_tx_pcs = {w_hssi_gen3_tx_pcs_avmmreaddata[7], w_hssi_gen3_tx_pcs_avmmreaddata[6], w_hssi_gen3_tx_pcs_avmmreaddata[5], w_hssi_gen3_tx_pcs_avmmreaddata[4], w_hssi_gen3_tx_pcs_avmmreaddata[3], w_hssi_gen3_tx_pcs_avmmreaddata[2], w_hssi_gen3_tx_pcs_avmmreaddata[1], w_hssi_gen3_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_rx_pcs = {w_hssi_krfec_rx_pcs_avmmreaddata[7], w_hssi_krfec_rx_pcs_avmmreaddata[6], w_hssi_krfec_rx_pcs_avmmreaddata[5], w_hssi_krfec_rx_pcs_avmmreaddata[4], w_hssi_krfec_rx_pcs_avmmreaddata[3], w_hssi_krfec_rx_pcs_avmmreaddata[2], w_hssi_krfec_rx_pcs_avmmreaddata[1], w_hssi_krfec_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_tx_pcs = {w_hssi_krfec_tx_pcs_avmmreaddata[7], w_hssi_krfec_tx_pcs_avmmreaddata[6], w_hssi_krfec_tx_pcs_avmmreaddata[5], w_hssi_krfec_tx_pcs_avmmreaddata[4], w_hssi_krfec_tx_pcs_avmmreaddata[3], w_hssi_krfec_tx_pcs_avmmreaddata[2], w_hssi_krfec_tx_pcs_avmmreaddata[1], w_hssi_krfec_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen1_2 = {w_hssi_pipe_gen1_2_avmmreaddata[7], w_hssi_pipe_gen1_2_avmmreaddata[6], w_hssi_pipe_gen1_2_avmmreaddata[5], w_hssi_pipe_gen1_2_avmmreaddata[4], w_hssi_pipe_gen1_2_avmmreaddata[3], w_hssi_pipe_gen1_2_avmmreaddata[2], w_hssi_pipe_gen1_2_avmmreaddata[1], w_hssi_pipe_gen1_2_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen3 = {w_hssi_pipe_gen3_avmmreaddata[7], w_hssi_pipe_gen3_avmmreaddata[6], w_hssi_pipe_gen3_avmmreaddata[5], w_hssi_pipe_gen3_avmmreaddata[4], w_hssi_pipe_gen3_avmmreaddata[3], w_hssi_pipe_gen3_avmmreaddata[2], w_hssi_pipe_gen3_avmmreaddata[1], w_hssi_pipe_gen3_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pcs_pma_interface = {w_hssi_rx_pcs_pma_interface_avmmreaddata[7], w_hssi_rx_pcs_pma_interface_avmmreaddata[6], w_hssi_rx_pcs_pma_interface_avmmreaddata[5], w_hssi_rx_pcs_pma_interface_avmmreaddata[4], w_hssi_rx_pcs_pma_interface_avmmreaddata[3], w_hssi_rx_pcs_pma_interface_avmmreaddata[2], w_hssi_rx_pcs_pma_interface_avmmreaddata[1], w_hssi_rx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pld_pcs_interface = {w_hssi_rx_pld_pcs_interface_avmmreaddata[7], w_hssi_rx_pld_pcs_interface_avmmreaddata[6], w_hssi_rx_pld_pcs_interface_avmmreaddata[5], w_hssi_rx_pld_pcs_interface_avmmreaddata[4], w_hssi_rx_pld_pcs_interface_avmmreaddata[3], w_hssi_rx_pld_pcs_interface_avmmreaddata[2], w_hssi_rx_pld_pcs_interface_avmmreaddata[1], w_hssi_rx_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pcs_pma_interface = {w_hssi_tx_pcs_pma_interface_avmmreaddata[7], w_hssi_tx_pcs_pma_interface_avmmreaddata[6], w_hssi_tx_pcs_pma_interface_avmmreaddata[5], w_hssi_tx_pcs_pma_interface_avmmreaddata[4], w_hssi_tx_pcs_pma_interface_avmmreaddata[3], w_hssi_tx_pcs_pma_interface_avmmreaddata[2], w_hssi_tx_pcs_pma_interface_avmmreaddata[1], w_hssi_tx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pld_pcs_interface = {w_hssi_tx_pld_pcs_interface_avmmreaddata[7], w_hssi_tx_pld_pcs_interface_avmmreaddata[6], w_hssi_tx_pld_pcs_interface_avmmreaddata[5], w_hssi_tx_pld_pcs_interface_avmmreaddata[4], w_hssi_tx_pld_pcs_interface_avmmreaddata[3], w_hssi_tx_pld_pcs_interface_avmmreaddata[2], w_hssi_tx_pld_pcs_interface_avmmreaddata[1], w_hssi_tx_pld_pcs_interface_avmmreaddata[0]};
		assign out_blockselect_hssi_10g_rx_pcs = w_hssi_10g_rx_pcs_blockselect;
		assign out_blockselect_hssi_10g_tx_pcs = w_hssi_10g_tx_pcs_blockselect;
		assign out_blockselect_hssi_8g_rx_pcs = w_hssi_8g_rx_pcs_blockselect;
		assign out_blockselect_hssi_8g_tx_pcs = w_hssi_8g_tx_pcs_blockselect;
		assign out_blockselect_hssi_common_pcs_pma_interface = w_hssi_common_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_common_pld_pcs_interface = w_hssi_common_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_fifo_rx_pcs = w_hssi_fifo_rx_pcs_blockselect;
		assign out_blockselect_hssi_fifo_tx_pcs = w_hssi_fifo_tx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_rx_pcs = w_hssi_gen3_rx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_tx_pcs = w_hssi_gen3_tx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_rx_pcs = w_hssi_krfec_rx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_tx_pcs = w_hssi_krfec_tx_pcs_blockselect;
		assign out_blockselect_hssi_pipe_gen1_2 = w_hssi_pipe_gen1_2_blockselect;
		assign out_blockselect_hssi_pipe_gen3 = w_hssi_pipe_gen3_blockselect;
		assign out_blockselect_hssi_rx_pcs_pma_interface = w_hssi_rx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_rx_pld_pcs_interface = w_hssi_rx_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_tx_pcs_pma_interface = w_hssi_tx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_tx_pld_pcs_interface = w_hssi_tx_pld_pcs_interface_blockselect;
		assign out_bond_pcs10g_out_bot = {w_hssi_10g_tx_pcs_distdwn_out_rden, w_hssi_10g_tx_pcs_distdwn_out_wren, w_hssi_10g_tx_pcs_distdwn_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs10g_out_top = {w_hssi_10g_tx_pcs_distup_out_rden, w_hssi_10g_tx_pcs_distup_out_wren, w_hssi_10g_tx_pcs_distup_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs8g_out_bot = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down, w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_down, w_hssi_8g_tx_pcs_wr_enable_out_chnl_down, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_down, w_hssi_8g_rx_pcs_wr_enable_out_chnl_down, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[0]};
		assign out_bond_pcs8g_out_top = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up, w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_up, w_hssi_8g_tx_pcs_wr_enable_out_chnl_up, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_up, w_hssi_8g_rx_pcs_wr_enable_out_chnl_up, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[0]};
		assign out_bond_pmaif_out_bot = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[0]};
		assign out_bond_pmaif_out_top = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[0]};
		assign out_hip_clk_out = {w_hssi_common_pld_pcs_interface_hip_cmn_clk[1], w_hssi_common_pld_pcs_interface_hip_cmn_clk[0], w_hssi_tx_pld_pcs_interface_hip_tx_clk};
		assign out_hip_ctrl_out = {w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[4], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[3], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[2], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[1], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[0], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[0]};
		assign out_hip_iocsr_rdy = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
		assign out_hip_iocsr_rdy_dly = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
		assign out_hip_nfrzdrv = w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
		assign out_hip_npor = w_hssi_common_pld_pcs_interface_hip_npor;
		assign out_hip_rx_data = {w_hssi_rx_pld_pcs_interface_hip_rx_data[50], w_hssi_rx_pld_pcs_interface_hip_rx_data[49], w_hssi_rx_pld_pcs_interface_hip_rx_data[48], w_hssi_rx_pld_pcs_interface_hip_rx_data[47], w_hssi_rx_pld_pcs_interface_hip_rx_data[46], w_hssi_rx_pld_pcs_interface_hip_rx_data[45], w_hssi_rx_pld_pcs_interface_hip_rx_data[44], w_hssi_rx_pld_pcs_interface_hip_rx_data[43], w_hssi_rx_pld_pcs_interface_hip_rx_data[42], w_hssi_rx_pld_pcs_interface_hip_rx_data[41], w_hssi_rx_pld_pcs_interface_hip_rx_data[40], w_hssi_rx_pld_pcs_interface_hip_rx_data[39], w_hssi_rx_pld_pcs_interface_hip_rx_data[38], w_hssi_rx_pld_pcs_interface_hip_rx_data[37], w_hssi_rx_pld_pcs_interface_hip_rx_data[36], w_hssi_rx_pld_pcs_interface_hip_rx_data[35], w_hssi_rx_pld_pcs_interface_hip_rx_data[34], w_hssi_rx_pld_pcs_interface_hip_rx_data[33], w_hssi_rx_pld_pcs_interface_hip_rx_data[32], w_hssi_rx_pld_pcs_interface_hip_rx_data[31], w_hssi_rx_pld_pcs_interface_hip_rx_data[30], w_hssi_rx_pld_pcs_interface_hip_rx_data[29], w_hssi_rx_pld_pcs_interface_hip_rx_data[28], w_hssi_rx_pld_pcs_interface_hip_rx_data[27], w_hssi_rx_pld_pcs_interface_hip_rx_data[26], w_hssi_rx_pld_pcs_interface_hip_rx_data[25], w_hssi_rx_pld_pcs_interface_hip_rx_data[24], w_hssi_rx_pld_pcs_interface_hip_rx_data[23], w_hssi_rx_pld_pcs_interface_hip_rx_data[22], w_hssi_rx_pld_pcs_interface_hip_rx_data[21], w_hssi_rx_pld_pcs_interface_hip_rx_data[20], w_hssi_rx_pld_pcs_interface_hip_rx_data[19], w_hssi_rx_pld_pcs_interface_hip_rx_data[18], w_hssi_rx_pld_pcs_interface_hip_rx_data[17], w_hssi_rx_pld_pcs_interface_hip_rx_data[16], w_hssi_rx_pld_pcs_interface_hip_rx_data[15], w_hssi_rx_pld_pcs_interface_hip_rx_data[14], w_hssi_rx_pld_pcs_interface_hip_rx_data[13], w_hssi_rx_pld_pcs_interface_hip_rx_data[12], w_hssi_rx_pld_pcs_interface_hip_rx_data[11], w_hssi_rx_pld_pcs_interface_hip_rx_data[10], w_hssi_rx_pld_pcs_interface_hip_rx_data[9], w_hssi_rx_pld_pcs_interface_hip_rx_data[8], w_hssi_rx_pld_pcs_interface_hip_rx_data[7], w_hssi_rx_pld_pcs_interface_hip_rx_data[6], w_hssi_rx_pld_pcs_interface_hip_rx_data[5], w_hssi_rx_pld_pcs_interface_hip_rx_data[4], w_hssi_rx_pld_pcs_interface_hip_rx_data[3], w_hssi_rx_pld_pcs_interface_hip_rx_data[2], w_hssi_rx_pld_pcs_interface_hip_rx_data[1], w_hssi_rx_pld_pcs_interface_hip_rx_data[0]};
		assign out_hip_usermode = w_hssi_common_pld_pcs_interface_hip_usermode;
		assign out_pld_10g_krfec_rx_blk_lock = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
		assign out_pld_10g_krfec_rx_diag_data_status = {w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1], w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[0]};
		assign out_pld_10g_krfec_rx_frame = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
		assign out_pld_10g_krfec_tx_frame = w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
		assign out_pld_10g_rx_align_val = w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
		assign out_pld_10g_rx_crc32_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
		assign out_pld_10g_rx_data_valid = w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
		assign out_pld_10g_rx_empty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
		assign out_pld_10g_rx_fifo_del = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
		assign out_pld_10g_rx_fifo_insert = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
		assign out_pld_10g_rx_fifo_num = {w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[3], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[2], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[1], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[0]};
		assign out_pld_10g_rx_frame_lock = w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
		assign out_pld_10g_rx_hi_ber = w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
		assign out_pld_10g_rx_oflw_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
		assign out_pld_10g_rx_pempty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
		assign out_pld_10g_rx_pfull = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
		assign out_pld_10g_tx_burst_en_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
		assign out_pld_10g_tx_empty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
		assign out_pld_10g_tx_fifo_num = {w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[2], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[1], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[0]};
		assign out_pld_10g_tx_full = w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
		assign out_pld_10g_tx_pempty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
		assign out_pld_10g_tx_pfull = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
		assign out_pld_10g_tx_wordslip_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
		assign out_pld_8g_a1a2_k1k2_flag = {w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[2], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[1], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[0]};
		assign out_pld_8g_empty_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
		assign out_pld_8g_empty_rx = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
		assign out_pld_8g_empty_tx = w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
		assign out_pld_8g_full_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
		assign out_pld_8g_full_rx = w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
		assign out_pld_8g_full_tx = w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
		assign out_pld_8g_rxelecidle = w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
		assign out_pld_8g_signal_detect_out = w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
		assign out_pld_8g_wa_boundary = {w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0]};
		assign out_pld_krfec_tx_alignment = w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
		assign out_pld_pcs_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
		assign out_pld_pcs_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
		assign out_pld_pma_adapt_done = w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
		assign out_pld_pma_clkdiv_rx_user = w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
		assign out_pld_pma_clkdiv_tx_user = w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
		assign out_pld_pma_clklow = w_hssi_common_pld_pcs_interface_pld_pma_clklow;
		assign out_pld_pma_fref = w_hssi_common_pld_pcs_interface_pld_pma_fref;
		assign out_pld_pma_hclk = w_hssi_common_pld_pcs_interface_pld_pma_hclk;
		assign out_pld_pma_pcie_sw_done = {w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1], w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[0]};
		assign out_pld_pma_pfdmode_lock = w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
		assign out_pld_pma_reserved_in = {w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[3], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[2], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[1], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[0]};
		assign out_pld_pma_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
		assign out_pld_pma_rx_detect_valid = w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
		assign out_pld_pma_rx_found = w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
		assign out_pld_pma_rxpll_lock = w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
		assign out_pld_pma_signal_ok = w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
		assign out_pld_pma_testbus = {w_hssi_common_pld_pcs_interface_pld_pma_testbus[7], w_hssi_common_pld_pcs_interface_pld_pma_testbus[6], w_hssi_common_pld_pcs_interface_pld_pma_testbus[5], w_hssi_common_pld_pcs_interface_pld_pma_testbus[4], w_hssi_common_pld_pcs_interface_pld_pma_testbus[3], w_hssi_common_pld_pcs_interface_pld_pma_testbus[2], w_hssi_common_pld_pcs_interface_pld_pma_testbus[1], w_hssi_common_pld_pcs_interface_pld_pma_testbus[0]};
		assign out_pld_pma_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
		assign out_pld_pmaif_mask_tx_pll = w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
		assign out_pld_reserved_out = {w_hssi_common_pld_pcs_interface_pld_reserved_out[9], w_hssi_common_pld_pcs_interface_pld_reserved_out[8], w_hssi_common_pld_pcs_interface_pld_reserved_out[7], w_hssi_common_pld_pcs_interface_pld_reserved_out[6], w_hssi_common_pld_pcs_interface_pld_reserved_out[5], w_hssi_common_pld_pcs_interface_pld_reserved_out[4], w_hssi_common_pld_pcs_interface_pld_reserved_out[3], w_hssi_common_pld_pcs_interface_pld_reserved_out[2], w_hssi_common_pld_pcs_interface_pld_reserved_out[1], w_hssi_common_pld_pcs_interface_pld_reserved_out[0]};
		assign out_pld_rx_control = {w_hssi_rx_pld_pcs_interface_pld_rx_control[19], w_hssi_rx_pld_pcs_interface_pld_rx_control[18], w_hssi_rx_pld_pcs_interface_pld_rx_control[17], w_hssi_rx_pld_pcs_interface_pld_rx_control[16], w_hssi_rx_pld_pcs_interface_pld_rx_control[15], w_hssi_rx_pld_pcs_interface_pld_rx_control[14], w_hssi_rx_pld_pcs_interface_pld_rx_control[13], w_hssi_rx_pld_pcs_interface_pld_rx_control[12], w_hssi_rx_pld_pcs_interface_pld_rx_control[11], w_hssi_rx_pld_pcs_interface_pld_rx_control[10], w_hssi_rx_pld_pcs_interface_pld_rx_control[9], w_hssi_rx_pld_pcs_interface_pld_rx_control[8], w_hssi_rx_pld_pcs_interface_pld_rx_control[7], w_hssi_rx_pld_pcs_interface_pld_rx_control[6], w_hssi_rx_pld_pcs_interface_pld_rx_control[5], w_hssi_rx_pld_pcs_interface_pld_rx_control[4], w_hssi_rx_pld_pcs_interface_pld_rx_control[3], w_hssi_rx_pld_pcs_interface_pld_rx_control[2], w_hssi_rx_pld_pcs_interface_pld_rx_control[1], w_hssi_rx_pld_pcs_interface_pld_rx_control[0]};
		assign out_pld_rx_data = {w_hssi_rx_pld_pcs_interface_pld_rx_data[127], w_hssi_rx_pld_pcs_interface_pld_rx_data[126], w_hssi_rx_pld_pcs_interface_pld_rx_data[125], w_hssi_rx_pld_pcs_interface_pld_rx_data[124], w_hssi_rx_pld_pcs_interface_pld_rx_data[123], w_hssi_rx_pld_pcs_interface_pld_rx_data[122], w_hssi_rx_pld_pcs_interface_pld_rx_data[121], w_hssi_rx_pld_pcs_interface_pld_rx_data[120], w_hssi_rx_pld_pcs_interface_pld_rx_data[119], w_hssi_rx_pld_pcs_interface_pld_rx_data[118], w_hssi_rx_pld_pcs_interface_pld_rx_data[117], w_hssi_rx_pld_pcs_interface_pld_rx_data[116], w_hssi_rx_pld_pcs_interface_pld_rx_data[115], w_hssi_rx_pld_pcs_interface_pld_rx_data[114], w_hssi_rx_pld_pcs_interface_pld_rx_data[113], w_hssi_rx_pld_pcs_interface_pld_rx_data[112], w_hssi_rx_pld_pcs_interface_pld_rx_data[111], w_hssi_rx_pld_pcs_interface_pld_rx_data[110], w_hssi_rx_pld_pcs_interface_pld_rx_data[109], w_hssi_rx_pld_pcs_interface_pld_rx_data[108], w_hssi_rx_pld_pcs_interface_pld_rx_data[107], w_hssi_rx_pld_pcs_interface_pld_rx_data[106], w_hssi_rx_pld_pcs_interface_pld_rx_data[105], w_hssi_rx_pld_pcs_interface_pld_rx_data[104], w_hssi_rx_pld_pcs_interface_pld_rx_data[103], w_hssi_rx_pld_pcs_interface_pld_rx_data[102], w_hssi_rx_pld_pcs_interface_pld_rx_data[101], w_hssi_rx_pld_pcs_interface_pld_rx_data[100], w_hssi_rx_pld_pcs_interface_pld_rx_data[99], w_hssi_rx_pld_pcs_interface_pld_rx_data[98], w_hssi_rx_pld_pcs_interface_pld_rx_data[97], w_hssi_rx_pld_pcs_interface_pld_rx_data[96], w_hssi_rx_pld_pcs_interface_pld_rx_data[95], w_hssi_rx_pld_pcs_interface_pld_rx_data[94], w_hssi_rx_pld_pcs_interface_pld_rx_data[93], w_hssi_rx_pld_pcs_interface_pld_rx_data[92], w_hssi_rx_pld_pcs_interface_pld_rx_data[91], w_hssi_rx_pld_pcs_interface_pld_rx_data[90], w_hssi_rx_pld_pcs_interface_pld_rx_data[89], w_hssi_rx_pld_pcs_interface_pld_rx_data[88], w_hssi_rx_pld_pcs_interface_pld_rx_data[87], w_hssi_rx_pld_pcs_interface_pld_rx_data[86], w_hssi_rx_pld_pcs_interface_pld_rx_data[85], w_hssi_rx_pld_pcs_interface_pld_rx_data[84], w_hssi_rx_pld_pcs_interface_pld_rx_data[83], w_hssi_rx_pld_pcs_interface_pld_rx_data[82], w_hssi_rx_pld_pcs_interface_pld_rx_data[81], w_hssi_rx_pld_pcs_interface_pld_rx_data[80], w_hssi_rx_pld_pcs_interface_pld_rx_data[79], w_hssi_rx_pld_pcs_interface_pld_rx_data[78], w_hssi_rx_pld_pcs_interface_pld_rx_data[77], w_hssi_rx_pld_pcs_interface_pld_rx_data[76], w_hssi_rx_pld_pcs_interface_pld_rx_data[75], w_hssi_rx_pld_pcs_interface_pld_rx_data[74], w_hssi_rx_pld_pcs_interface_pld_rx_data[73], w_hssi_rx_pld_pcs_interface_pld_rx_data[72], w_hssi_rx_pld_pcs_interface_pld_rx_data[71], w_hssi_rx_pld_pcs_interface_pld_rx_data[70], w_hssi_rx_pld_pcs_interface_pld_rx_data[69], w_hssi_rx_pld_pcs_interface_pld_rx_data[68], w_hssi_rx_pld_pcs_interface_pld_rx_data[67], w_hssi_rx_pld_pcs_interface_pld_rx_data[66], w_hssi_rx_pld_pcs_interface_pld_rx_data[65], w_hssi_rx_pld_pcs_interface_pld_rx_data[64], w_hssi_rx_pld_pcs_interface_pld_rx_data[63], w_hssi_rx_pld_pcs_interface_pld_rx_data[62], w_hssi_rx_pld_pcs_interface_pld_rx_data[61], w_hssi_rx_pld_pcs_interface_pld_rx_data[60], w_hssi_rx_pld_pcs_interface_pld_rx_data[59], w_hssi_rx_pld_pcs_interface_pld_rx_data[58], w_hssi_rx_pld_pcs_interface_pld_rx_data[57], w_hssi_rx_pld_pcs_interface_pld_rx_data[56], w_hssi_rx_pld_pcs_interface_pld_rx_data[55], w_hssi_rx_pld_pcs_interface_pld_rx_data[54], w_hssi_rx_pld_pcs_interface_pld_rx_data[53], w_hssi_rx_pld_pcs_interface_pld_rx_data[52], w_hssi_rx_pld_pcs_interface_pld_rx_data[51], w_hssi_rx_pld_pcs_interface_pld_rx_data[50], w_hssi_rx_pld_pcs_interface_pld_rx_data[49], w_hssi_rx_pld_pcs_interface_pld_rx_data[48], w_hssi_rx_pld_pcs_interface_pld_rx_data[47], w_hssi_rx_pld_pcs_interface_pld_rx_data[46], w_hssi_rx_pld_pcs_interface_pld_rx_data[45], w_hssi_rx_pld_pcs_interface_pld_rx_data[44], w_hssi_rx_pld_pcs_interface_pld_rx_data[43], w_hssi_rx_pld_pcs_interface_pld_rx_data[42], w_hssi_rx_pld_pcs_interface_pld_rx_data[41], w_hssi_rx_pld_pcs_interface_pld_rx_data[40], w_hssi_rx_pld_pcs_interface_pld_rx_data[39], w_hssi_rx_pld_pcs_interface_pld_rx_data[38], w_hssi_rx_pld_pcs_interface_pld_rx_data[37], w_hssi_rx_pld_pcs_interface_pld_rx_data[36], w_hssi_rx_pld_pcs_interface_pld_rx_data[35], w_hssi_rx_pld_pcs_interface_pld_rx_data[34], w_hssi_rx_pld_pcs_interface_pld_rx_data[33], w_hssi_rx_pld_pcs_interface_pld_rx_data[32], w_hssi_rx_pld_pcs_interface_pld_rx_data[31], w_hssi_rx_pld_pcs_interface_pld_rx_data[30], w_hssi_rx_pld_pcs_interface_pld_rx_data[29], w_hssi_rx_pld_pcs_interface_pld_rx_data[28], w_hssi_rx_pld_pcs_interface_pld_rx_data[27], w_hssi_rx_pld_pcs_interface_pld_rx_data[26], w_hssi_rx_pld_pcs_interface_pld_rx_data[25], w_hssi_rx_pld_pcs_interface_pld_rx_data[24], w_hssi_rx_pld_pcs_interface_pld_rx_data[23], w_hssi_rx_pld_pcs_interface_pld_rx_data[22], w_hssi_rx_pld_pcs_interface_pld_rx_data[21], w_hssi_rx_pld_pcs_interface_pld_rx_data[20], w_hssi_rx_pld_pcs_interface_pld_rx_data[19], w_hssi_rx_pld_pcs_interface_pld_rx_data[18], w_hssi_rx_pld_pcs_interface_pld_rx_data[17], w_hssi_rx_pld_pcs_interface_pld_rx_data[16], w_hssi_rx_pld_pcs_interface_pld_rx_data[15], w_hssi_rx_pld_pcs_interface_pld_rx_data[14], w_hssi_rx_pld_pcs_interface_pld_rx_data[13], w_hssi_rx_pld_pcs_interface_pld_rx_data[12], w_hssi_rx_pld_pcs_interface_pld_rx_data[11], w_hssi_rx_pld_pcs_interface_pld_rx_data[10], w_hssi_rx_pld_pcs_interface_pld_rx_data[9], w_hssi_rx_pld_pcs_interface_pld_rx_data[8], w_hssi_rx_pld_pcs_interface_pld_rx_data[7], w_hssi_rx_pld_pcs_interface_pld_rx_data[6], w_hssi_rx_pld_pcs_interface_pld_rx_data[5], w_hssi_rx_pld_pcs_interface_pld_rx_data[4], w_hssi_rx_pld_pcs_interface_pld_rx_data[3], w_hssi_rx_pld_pcs_interface_pld_rx_data[2], w_hssi_rx_pld_pcs_interface_pld_rx_data[1], w_hssi_rx_pld_pcs_interface_pld_rx_data[0]};
		assign out_pld_rx_prbs_done = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
		assign out_pld_rx_prbs_err = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
		assign out_pld_test_data = {w_hssi_common_pld_pcs_interface_pld_test_data[19], w_hssi_common_pld_pcs_interface_pld_test_data[18], w_hssi_common_pld_pcs_interface_pld_test_data[17], w_hssi_common_pld_pcs_interface_pld_test_data[16], w_hssi_common_pld_pcs_interface_pld_test_data[15], w_hssi_common_pld_pcs_interface_pld_test_data[14], w_hssi_common_pld_pcs_interface_pld_test_data[13], w_hssi_common_pld_pcs_interface_pld_test_data[12], w_hssi_common_pld_pcs_interface_pld_test_data[11], w_hssi_common_pld_pcs_interface_pld_test_data[10], w_hssi_common_pld_pcs_interface_pld_test_data[9], w_hssi_common_pld_pcs_interface_pld_test_data[8], w_hssi_common_pld_pcs_interface_pld_test_data[7], w_hssi_common_pld_pcs_interface_pld_test_data[6], w_hssi_common_pld_pcs_interface_pld_test_data[5], w_hssi_common_pld_pcs_interface_pld_test_data[4], w_hssi_common_pld_pcs_interface_pld_test_data[3], w_hssi_common_pld_pcs_interface_pld_test_data[2], w_hssi_common_pld_pcs_interface_pld_test_data[1], w_hssi_common_pld_pcs_interface_pld_test_data[0]};
		assign out_pld_uhsif_lock = w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
		assign out_pld_uhsif_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
		assign out_pma_adapt_start = w_hssi_common_pcs_pma_interface_pma_adapt_start;
		assign out_pma_atpg_los_en_n = w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
		assign out_pma_csr_test_dis = w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
		assign out_pma_current_coeff = {w_hssi_common_pcs_pma_interface_pma_current_coeff[17], w_hssi_common_pcs_pma_interface_pma_current_coeff[16], w_hssi_common_pcs_pma_interface_pma_current_coeff[15], w_hssi_common_pcs_pma_interface_pma_current_coeff[14], w_hssi_common_pcs_pma_interface_pma_current_coeff[13], w_hssi_common_pcs_pma_interface_pma_current_coeff[12], w_hssi_common_pcs_pma_interface_pma_current_coeff[11], w_hssi_common_pcs_pma_interface_pma_current_coeff[10], w_hssi_common_pcs_pma_interface_pma_current_coeff[9], w_hssi_common_pcs_pma_interface_pma_current_coeff[8], w_hssi_common_pcs_pma_interface_pma_current_coeff[7], w_hssi_common_pcs_pma_interface_pma_current_coeff[6], w_hssi_common_pcs_pma_interface_pma_current_coeff[5], w_hssi_common_pcs_pma_interface_pma_current_coeff[4], w_hssi_common_pcs_pma_interface_pma_current_coeff[3], w_hssi_common_pcs_pma_interface_pma_current_coeff[2], w_hssi_common_pcs_pma_interface_pma_current_coeff[1], w_hssi_common_pcs_pma_interface_pma_current_coeff[0]};
		assign out_pma_current_rxpreset = {w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[1], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[0]};
		assign out_pma_early_eios = w_hssi_common_pcs_pma_interface_pma_early_eios;
		assign out_pma_eye_monitor = {w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0]};
		assign out_pma_interface_select = {w_hssi_common_pcs_pma_interface_pma_interface_select[1], w_hssi_common_pcs_pma_interface_pma_interface_select[0]};
		assign out_pma_ltd_b = w_hssi_common_pcs_pma_interface_pma_ltd_b;
		assign out_pma_ltr = w_hssi_common_pcs_pma_interface_pma_ltr;
		assign out_pma_nfrzdrv = w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
		assign out_pma_nrpi_freeze = w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
		assign out_pma_pcie_switch = {w_hssi_common_pcs_pma_interface_pma_pcie_switch[1], w_hssi_common_pcs_pma_interface_pma_pcie_switch[0]};
		assign out_pma_ppm_lock = w_hssi_common_pcs_pma_interface_pma_ppm_lock;
		assign out_pma_reserved_out = {w_hssi_common_pcs_pma_interface_pma_reserved_out[4], w_hssi_common_pcs_pma_interface_pma_reserved_out[3], w_hssi_common_pcs_pma_interface_pma_reserved_out[2], w_hssi_common_pcs_pma_interface_pma_reserved_out[1], w_hssi_common_pcs_pma_interface_pma_reserved_out[0]};
		assign out_pma_rs_lpbk_b = w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
		assign out_pma_rx_clkslip = w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
		assign out_pma_rx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
		assign out_pma_rxpma_rstb = w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
		assign out_pma_scan_mode_n = w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
		assign out_pma_scan_shift_n = w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
		assign out_pma_tx_bitslip = w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
		assign out_pma_tx_bonding_rstb = w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
		assign out_pma_tx_elec_idle = w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
		assign out_pma_tx_pma_data = {w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0]};
		assign out_pma_tx_qpi_pulldn = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
		assign out_pma_tx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
		assign out_pma_tx_txdetectrx = w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
		assign out_pma_txpma_rstb = w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	endgenerate
endmodule
module twentynm_pcs_rev_20nm2
	#(
	//PARAM_LIST_START
		parameter xcvr_native_mode = "mode_duplex",  // mode_duplex, mode_rx_only, mode_tx_only
		
		// parameters for twentynm_hssi_10g_rx_pcs
		parameter hssi_10g_rx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_align_del = "align_del_en", // align_del_dis|align_del_en
		parameter hssi_10g_rx_pcs_ber_bit_err_total_cnt = "bit_err_total_cnt_10g", // bit_err_total_cnt_10g
		parameter hssi_10g_rx_pcs_ber_clken = "ber_clk_dis", // ber_clk_dis|ber_clk_en
		parameter hssi_10g_rx_pcs_ber_xus_timer_window = 21'b100110001001010,
		parameter hssi_10g_rx_pcs_bitslip_mode = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_rx_pcs_blksync_bitslip_type = "bitslip_comb", // bitslip_comb|bitslip_reg
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_cnt = 3'b1,
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_type = "bitslip_match", // bitslip_match|bitslip_cnt
		parameter hssi_10g_rx_pcs_blksync_bypass = "blksync_bypass_dis", // blksync_bypass_dis|blksync_bypass_en
		parameter hssi_10g_rx_pcs_blksync_clken = "blksync_clk_dis", // blksync_clk_dis|blksync_clk_en
		parameter hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt = "enum_invalid_sh_cnt_10g", // enum_invalid_sh_cnt_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock = "knum_sh_cnt_postlock_10g", // knum_sh_cnt_postlock_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock = "knum_sh_cnt_prelock_10g", // knum_sh_cnt_prelock_10g
		parameter hssi_10g_rx_pcs_blksync_pipeln = "blksync_pipeln_dis", // blksync_pipeln_dis|blksync_pipeln_en
		parameter hssi_10g_rx_pcs_clr_errblk_cnt_en = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_control_del = "control_del_all", // control_del_all|control_del_none
		parameter hssi_10g_rx_pcs_crcchk_bypass = "crcchk_bypass_dis", // crcchk_bypass_dis|crcchk_bypass_en
		parameter hssi_10g_rx_pcs_crcchk_clken = "crcchk_clk_dis", // crcchk_clk_dis|crcchk_clk_en
		parameter hssi_10g_rx_pcs_crcchk_inv = "crcchk_inv_dis", // crcchk_inv_dis|crcchk_inv_en
		parameter hssi_10g_rx_pcs_crcchk_pipeln = "crcchk_pipeln_dis", // crcchk_pipeln_dis|crcchk_pipeln_en
		parameter hssi_10g_rx_pcs_crcflag_pipeln = "crcflag_pipeln_dis", // crcflag_pipeln_dis|crcflag_pipeln_en
		parameter hssi_10g_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_rx_pcs_dec64b66b_clken = "dec64b66b_clk_dis", // dec64b66b_clk_dis|dec64b66b_clk_en
		parameter hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass = "dec_64b66b_rxsm_bypass_dis", // dec_64b66b_rxsm_bypass_dis|dec_64b66b_rxsm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_bypass = "descrm_bypass_en", // descrm_bypass_dis|descrm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_clken = "descrm_clk_dis", // descrm_clk_dis|descrm_clk_en
		parameter hssi_10g_rx_pcs_descrm_mode = "async", // async|sync
		parameter hssi_10g_rx_pcs_descrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_dft_clk_out_sel = "rx_master_clk", // rx_master_clk|rx_gbexp_clk|rx_blksync_clk|rx_descrm_clk|rx_frmsync_clk|rx_64b66bdec_clk|rx_ber_clk|rx_rand_clk|rx_crcchk_clk|rx_wrfifo_clk|rx_rdfifo_clk|rx_fec_clk
		parameter hssi_10g_rx_pcs_dis_signal_ok = "dis_signal_ok_dis", // dis_signal_ok_dis|dis_signal_ok_en
		parameter hssi_10g_rx_pcs_dispchk_bypass = "dispchk_bypass_dis", // dispchk_bypass_dis|dispchk_bypass_en
		parameter hssi_10g_rx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_rx_pcs_fast_path = "fast_path_dis", // fast_path_dis|fast_path_en
		parameter hssi_10g_rx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_rx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_rx_pcs_fifo_double_read = "fifo_double_read_dis", // fifo_double_read_dis|fifo_double_read_en
		parameter hssi_10g_rx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_rx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_rx_pcs_force_align = "force_align_dis", // force_align_dis|force_align_en
		parameter hssi_10g_rx_pcs_frmsync_bypass = "frmsync_bypass_dis", // frmsync_bypass_dis|frmsync_bypass_en
		parameter hssi_10g_rx_pcs_frmsync_clken = "frmsync_clk_dis", // frmsync_clk_dis|frmsync_clk_en
		parameter hssi_10g_rx_pcs_frmsync_enum_scrm = "enum_scrm_default", // enum_scrm_default
		parameter hssi_10g_rx_pcs_frmsync_enum_sync = "enum_sync_default", // enum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_flag_type = "all_framing_words", // all_framing_words|location_only
		parameter hssi_10g_rx_pcs_frmsync_knum_sync = "knum_sync_default", // knum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_mfrm_length = 16'b100000000000,
		parameter hssi_10g_rx_pcs_frmsync_pipeln = "frmsync_pipeln_dis", // frmsync_pipeln_dis|frmsync_pipeln_en
		parameter hssi_10g_rx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_rx_pcs_gb_rx_idwidth = "width_32", // width_40|width_32|width_64
		parameter hssi_10g_rx_pcs_gb_rx_odwidth = "width_66", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_rx_pcs_gbexp_clken = "gbexp_clk_dis", // gbexp_clk_dis|gbexp_clk_en
		parameter hssi_10g_rx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_10g_rx_pcs_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_rx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_rx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_rx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_rx_pcs_pld_if_type = "fifo", // fifo|reg
		parameter hssi_10g_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_rx_pcs_rand_clken = "rand_clk_dis", // rand_clk_dis|rand_clk_en
		parameter hssi_10g_rx_pcs_rd_clk_sel = "rd_rx_pma_clk", // rd_rx_pld_clk|rd_rx_pma_clk|rd_refclk_dig
		parameter hssi_10g_rx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_rx_pcs_rx_fifo_write_ctrl = "blklock_stops", // blklock_stops|blklock_ignore
		parameter hssi_10g_rx_pcs_rx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_rx_pcs_rx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_rx_pcs_rx_signal_ok_sel = "synchronized_ver", // synchronized_ver|nonsync_ver
		parameter hssi_10g_rx_pcs_rx_sm_bypass = "rx_sm_bypass_dis", // rx_sm_bypass_dis|rx_sm_bypass_en
		parameter hssi_10g_rx_pcs_rx_sm_hiber = "rx_sm_hiber_en", // rx_sm_hiber_en|rx_sm_hiber_dis
		parameter hssi_10g_rx_pcs_rx_sm_pipeln = "rx_sm_pipeln_dis", // rx_sm_pipeln_dis|rx_sm_pipeln_en
		parameter hssi_10g_rx_pcs_rx_testbus_sel = "crc32_chk_testbus1", // crc32_chk_testbus1|crc32_chk_testbus2|frame_sync_testbus1|frame_sync_testbus2|dec64b66b_testbus|rxsm_testbus|ber_testbus|blksync_testbus1|blksync_testbus2|gearbox_exp_testbus|random_ver_testbus|descramble_testbus|blank_testbus|rx_fifo_testbus1|rx_fifo_testbus2
		parameter hssi_10g_rx_pcs_rx_true_b2b = "b2b", // single|b2b
		parameter hssi_10g_rx_pcs_rxfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_rx_pcs_rxfifo_full = "full_default", // full_default
		parameter hssi_10g_rx_pcs_rxfifo_mode = "phase_comp", // register_mode|clk_comp_10g|generic_interlaken|generic_basic|phase_comp|phase_comp_dv
		parameter hssi_10g_rx_pcs_rxfifo_pempty = 5'b10,
		parameter hssi_10g_rx_pcs_rxfifo_pfull = 5'b10111,
		parameter hssi_10g_rx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_rx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_rx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_10g_tx_pcs
		parameter hssi_10g_tx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_bitslip_en = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_10g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_10g_tx_pcs_comp_cnt = 8'b0,
		parameter hssi_10g_tx_pcs_compin_sel = "compin_master", // compin_master|compin_slave_top|compin_slave_bot|compin_default
		parameter hssi_10g_tx_pcs_crcgen_bypass = "crcgen_bypass_dis", // crcgen_bypass_dis|crcgen_bypass_en
		parameter hssi_10g_tx_pcs_crcgen_clken = "crcgen_clk_dis", // crcgen_clk_dis|crcgen_clk_en
		parameter hssi_10g_tx_pcs_crcgen_err = "crcgen_err_dis", // crcgen_err_dis|crcgen_err_en
		parameter hssi_10g_tx_pcs_crcgen_inv = "crcgen_inv_dis", // crcgen_inv_dis|crcgen_inv_en
		parameter hssi_10g_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_tx_pcs_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_10g_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_tx_pcs_dft_clk_out_sel = "tx_master_clk", // tx_master_clk|tx_rdfifo_clk|tx_frmgen_clk|tx_crcgen_clk|tx_64b66benc_txsm_clk|tx_scrm_clk|tx_dispgen_clk|tx_gbred_clk|tx_wrfifo_clk|tx_fec_clk
		parameter hssi_10g_tx_pcs_dispgen_bypass = "dispgen_bypass_dis", // dispgen_bypass_dis|dispgen_bypass_en
		parameter hssi_10g_tx_pcs_dispgen_clken = "dispgen_clk_dis", // dispgen_clk_dis|dispgen_clk_en
		parameter hssi_10g_tx_pcs_dispgen_err = "dispgen_err_dis", // dispgen_err_dis|dispgen_err_en
		parameter hssi_10g_tx_pcs_dispgen_pipeln = "dispgen_pipeln_dis", // dispgen_pipeln_dis|dispgen_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_bypass_pipeln = "distdwn_bypass_pipeln_dis", // distdwn_bypass_pipeln_dis|distdwn_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_master = "distdwn_master_en", // distdwn_master_en|distdwn_master_dis
		parameter hssi_10g_tx_pcs_distup_bypass_pipeln = "distup_bypass_pipeln_dis", // distup_bypass_pipeln_dis|distup_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distup_master = "distup_master_en", // distup_master_en|distup_master_dis
		parameter hssi_10g_tx_pcs_dv_bond = "dv_bond_dis", // dv_bond_en|dv_bond_dis
		parameter hssi_10g_tx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_tx_pcs_enc64b66b_txsm_clken = "enc64b66b_txsm_clk_dis", // enc64b66b_txsm_clk_dis|enc64b66b_txsm_clk_en
		parameter hssi_10g_tx_pcs_enc_64b66b_txsm_bypass = "enc_64b66b_txsm_bypass_dis", // enc_64b66b_txsm_bypass_dis|enc_64b66b_txsm_bypass_en
		parameter hssi_10g_tx_pcs_fastpath = "fastpath_dis", // fastpath_dis|fastpath_en
		parameter hssi_10g_tx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_tx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_tx_pcs_fifo_double_write = "fifo_double_write_dis", // fifo_double_write_dis|fifo_double_write_en
		parameter hssi_10g_tx_pcs_fifo_reg_fast = "fifo_reg_fast_dis", // fifo_reg_fast_dis|fifo_reg_fast_en
		parameter hssi_10g_tx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_tx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_tx_pcs_frmgen_burst = "frmgen_burst_dis", // frmgen_burst_dis|frmgen_burst_en
		parameter hssi_10g_tx_pcs_frmgen_bypass = "frmgen_bypass_dis", // frmgen_bypass_dis|frmgen_bypass_en
		parameter hssi_10g_tx_pcs_frmgen_clken = "frmgen_clk_dis", // frmgen_clk_dis|frmgen_clk_en
		parameter hssi_10g_tx_pcs_frmgen_mfrm_length = 16'b100000000000,
		parameter hssi_10g_tx_pcs_frmgen_pipeln = "frmgen_pipeln_dis", // frmgen_pipeln_dis|frmgen_pipeln_en
		parameter hssi_10g_tx_pcs_frmgen_pyld_ins = "frmgen_pyld_ins_dis", // frmgen_pyld_ins_dis|frmgen_pyld_ins_en
		parameter hssi_10g_tx_pcs_frmgen_wordslip = "frmgen_wordslip_dis", // frmgen_wordslip_dis|frmgen_wordslip_en
		parameter hssi_10g_tx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_tx_pcs_gb_pipeln_bypass = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_gb_tx_idwidth = "width_50", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_tx_pcs_gb_tx_odwidth = "width_32", // width_32|width_40|width_64
		parameter hssi_10g_tx_pcs_gbred_clken = "gbred_clk_dis", // gbred_clk_dis|gbred_clk_en
		parameter hssi_10g_tx_pcs_indv = "indv_en", // indv_en|indv_dis
		parameter hssi_10g_tx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_tx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_tx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_tx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del6|phcomp_rd_del5|phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_tx_pcs_pld_if_type = "fifo", // fifo|reg|fastreg
		parameter hssi_10g_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_tx_pcs_pseudo_random = "all_0", // two_lf|all_0
		parameter hssi_10g_tx_pcs_pseudo_seed_a = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_pseudo_seed_b = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_random_disp = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_tx_pcs_scrm_bypass = "scrm_bypass_dis", // scrm_bypass_dis|scrm_bypass_en
		parameter hssi_10g_tx_pcs_scrm_clken = "scrm_clk_dis", // scrm_clk_dis|scrm_clk_en
		parameter hssi_10g_tx_pcs_scrm_mode = "async", // async|sync
		parameter hssi_10g_tx_pcs_scrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_sh_err = "sh_err_dis", // sh_err_dis|sh_err_en
		parameter hssi_10g_tx_pcs_sop_mark = "sop_mark_dis", // sop_mark_en|sop_mark_dis
		parameter hssi_10g_tx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_tx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_tx_pcs_tx_scrm_err = "scrm_err_dis", // scrm_err_dis|scrm_err_en
		parameter hssi_10g_tx_pcs_tx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_tx_pcs_tx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_tx_pcs_tx_sm_bypass = "tx_sm_bypass_dis", // tx_sm_bypass_dis|tx_sm_bypass_en
		parameter hssi_10g_tx_pcs_tx_sm_pipeln = "tx_sm_pipeln_dis", // tx_sm_pipeln_dis|tx_sm_pipeln_en
		parameter hssi_10g_tx_pcs_tx_testbus_sel = "crc32_gen_testbus1", // crc32_gen_testbus1|crc32_gen_testbus2|disp_gen_testbus1|disp_gen_testbus2|frame_gen_testbus1|frame_gen_testbus2|enc64b66b_testbus|txsm_testbus|tx_cp_bond_testbus|gearbox_red_testbus|scramble_testbus|blank_testbus|tx_fifo_testbus1|tx_fifo_testbus2
		parameter hssi_10g_tx_pcs_txfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_tx_pcs_txfifo_full = "full_default", // full_default
		parameter hssi_10g_tx_pcs_txfifo_mode = "phase_comp", // register_mode|interlaken_generic|basic_generic|phase_comp
		parameter hssi_10g_tx_pcs_txfifo_pempty = 4'b10,
		parameter hssi_10g_tx_pcs_txfifo_pfull = 4'b1011,
		parameter hssi_10g_tx_pcs_wr_clk_sel = "wr_tx_pma_clk", // wr_tx_pld_clk|wr_tx_pma_clk|wr_refclk_dig
		parameter hssi_10g_tx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_8g_rx_pcs
		parameter hssi_8g_rx_pcs_auto_error_replacement = "dis_err_replace", // dis_err_replace|en_err_replace
		parameter hssi_8g_rx_pcs_auto_speed_nego = "dis_asn", // dis_asn|en_asn_g2_freq_scal
		parameter hssi_8g_rx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_rx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_rx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_rx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_rx_pcs_byte_deserializer = "dis_bds", // dis_bds|en_bds_by_2|en_bds_by_4|en_bds_by_2_det
		parameter hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask = "dis_rxvalid_mask", // dis_rxvalid_mask|en_rxvalid_mask
		parameter hssi_8g_rx_pcs_clkcmp_pattern_n = 20'b0,
		parameter hssi_8g_rx_pcs_clkcmp_pattern_p = 20'b0,
		parameter hssi_8g_rx_pcs_clock_gate_bds_dec_asn = "dis_bds_dec_asn_clk_gating", // dis_bds_dec_asn_clk_gating|en_bds_dec_asn_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_cdr_eidle = "dis_cdr_eidle_clk_gating", // dis_cdr_eidle_clk_gating|en_cdr_eidle_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk = "dis_dw_pc_wrclk_gating", // dis_dw_pc_wrclk_gating|en_dw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_rd = "dis_dw_rm_rdclk_gating", // dis_dw_rm_rdclk_gating|en_dw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_wr = "dis_dw_rm_wrclk_gating", // dis_dw_rm_wrclk_gating|en_dw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_wa = "dis_dw_wa_clk_gating", // dis_dw_wa_clk_gating|en_dw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_pc_rdclk = "dis_pc_rdclk_gating", // dis_pc_rdclk_gating|en_pc_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk = "dis_sw_pc_wrclk_gating", // dis_sw_pc_wrclk_gating|en_sw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_rd = "dis_sw_rm_rdclk_gating", // dis_sw_rm_rdclk_gating|en_sw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_wr = "dis_sw_rm_wrclk_gating", // dis_sw_rm_wrclk_gating|en_sw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_wa = "dis_sw_wa_clk_gating", // dis_sw_wa_clk_gating|en_sw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_observation_in_pld_core = "internal_sw_wa_clk", // internal_sw_wa_clk|internal_dw_wa_clk|internal_cdr_eidle_clk|internal_sm_rm_wr_clk|internal_dw_rm_wr_clk|internal_clk_2_b|internal_sw_rm_rd_clk|internal_dw_rm_rd_clk|internal_sw_rx_wr_clk|internal_dw_rx_wr_clk|internal_rx_rd_clk|internal_rx_pma_clk_gen3|internal_rx_rcvd_clk_gen3
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_rx_pcs_eidle_entry_eios = "dis_eidle_eios", // dis_eidle_eios|en_eidle_eios
		parameter hssi_8g_rx_pcs_eidle_entry_iei = "dis_eidle_iei", // dis_eidle_iei|en_eidle_iei
		parameter hssi_8g_rx_pcs_eidle_entry_sd = "dis_eidle_sd", // dis_eidle_sd|en_eidle_sd
		parameter hssi_8g_rx_pcs_eightb_tenb_decoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_rx_pcs_err_flags_sel = "err_flags_wa", // err_flags_wa|err_flags_8b10b
		parameter hssi_8g_rx_pcs_fixed_pat_det = "dis_fixed_patdet", // dis_fixed_patdet|en_fixed_patdet
		parameter hssi_8g_rx_pcs_fixed_pat_num = 4'b1111,
		parameter hssi_8g_rx_pcs_force_signal_detect = "en_force_signal_detect", // en_force_signal_detect|dis_force_signal_detect
		parameter hssi_8g_rx_pcs_gen3_clk_en = "disable_clk", // disable_clk|enable_clk
		parameter hssi_8g_rx_pcs_gen3_rx_clk_sel = "rcvd_clk", // en_dig_clk1_8g|rcvd_clk
		parameter hssi_8g_rx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // en_dig_clk2_8g|tx_pma_clk
		parameter hssi_8g_rx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_rx_pcs_ibm_invalid_code = "dis_ibm_invalid_code", // dis_ibm_invalid_code|en_ibm_invalid_code
		parameter hssi_8g_rx_pcs_invalid_code_flag_only = "dis_invalid_code_only", // dis_invalid_code_only|en_invalid_code_only
		parameter hssi_8g_rx_pcs_pad_or_edb_error_replace = "replace_edb", // replace_edb|replace_edb_dynamic|replace_pad
		parameter hssi_8g_rx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_rx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_rx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_rx_pcs_pipe_if_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_8g_rx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_rx_pcs_polinv_8b10b_dec = "dis_polinv_8b10b_dec", // dis_polinv_8b10b_dec|en_polinv_8b10b_dec
		parameter hssi_8g_rx_pcs_prot_mode = "gige", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic_rm_enable|basic_rm_disable|disabled_prot_mode
		parameter hssi_8g_rx_pcs_rate_match = "dis_rm", // dis_rm|gige_rm|pipe_rm|pipe_rm_0ppm|sw_basic_rm|dw_basic_rm
		parameter hssi_8g_rx_pcs_rate_match_del_thres = "dis_rm_del_thres", // dis_rm_del_thres|gige_rm_del_thres|pipe_rm_del_thres|pipe_rm_0ppm_del_thres|sw_basic_rm_del_thres|dw_basic_rm_del_thres
		parameter hssi_8g_rx_pcs_rate_match_empty_thres = "dis_rm_empty_thres", // dis_rm_empty_thres|gige_rm_empty_thres|pipe_rm_empty_thres|pipe_rm_0ppm_empty_thres|sw_basic_rm_empty_thres|dw_basic_rm_empty_thres
		parameter hssi_8g_rx_pcs_rate_match_full_thres = "dis_rm_full_thres", // dis_rm_full_thres|gige_rm_full_thres|pipe_rm_full_thres|pipe_rm_0ppm_full_thres|sw_basic_rm_full_thres|dw_basic_rm_full_thres
		parameter hssi_8g_rx_pcs_rate_match_ins_thres = "dis_rm_ins_thres", // dis_rm_ins_thres|gige_rm_ins_thres|pipe_rm_ins_thres|pipe_rm_0ppm_ins_thres|sw_basic_rm_ins_thres|dw_basic_rm_ins_thres
		parameter hssi_8g_rx_pcs_rate_match_start_thres = "dis_rm_start_thres", // dis_rm_start_thres|gige_rm_start_thres|pipe_rm_start_thres|pipe_rm_0ppm_start_thres|sw_basic_rm_start_thres|dw_basic_rm_start_thres
		parameter hssi_8g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_rx_pcs_rx_clk2 = "rcvd_clk_clk2", // rcvd_clk_clk2|tx_pma_clock_clk2|refclk_dig2_clk2
		parameter hssi_8g_rx_pcs_rx_clk_free_running = "en_rx_clk_free_run", // dis_rx_clk_free_run|en_rx_clk_free_run
		parameter hssi_8g_rx_pcs_rx_pcs_urst = "en_rx_pcs_urst", // dis_rx_pcs_urst|en_rx_pcs_urst
		parameter hssi_8g_rx_pcs_rx_rcvd_clk = "rcvd_clk_rcvd_clk", // rcvd_clk_rcvd_clk|tx_pma_clock_rcvd_clk
		parameter hssi_8g_rx_pcs_rx_rd_clk = "pld_rx_clk", // pld_rx_clk|rx_clk
		parameter hssi_8g_rx_pcs_rx_refclk = "dis_refclk_sel", // dis_refclk_sel|en_refclk_sel
		parameter hssi_8g_rx_pcs_rx_wr_clk = "rx_clk2_div_1_2_4", // rx_clk2_div_1_2_4|txfifo_rd_clk
		parameter hssi_8g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_rx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_rx_pcs_sync_sm_idle_eios = "dis_syncsm_idle", // dis_syncsm_idle|en_syncsm_idle
		parameter hssi_8g_rx_pcs_test_bus_sel = "tx_testbus", // tx_testbus|tx_ctrl_plane_testbus|wa_testbus|rm_testbus|rx_ctrl_testbus|pcie_ctrl_testbus|rx_ctrl_plane_testbus
		parameter hssi_8g_rx_pcs_tx_rx_parallel_loopback = "dis_plpbk", // dis_plpbk|en_plpbk
		parameter hssi_8g_rx_pcs_wa_boundary_lock_ctrl = "bit_slip", // bit_slip|sync_sm|deterministic_latency|auto_align_pld_ctrl
		parameter hssi_8g_rx_pcs_wa_clk_slip_spacing = 10'b10000,
		parameter hssi_8g_rx_pcs_wa_det_latency_sync_status_beh = "assert_sync_status_non_imm", // assert_sync_status_imm|assert_sync_status_non_imm|dont_care_assert_sync
		parameter hssi_8g_rx_pcs_wa_disp_err_flag = "dis_disp_err_flag", // dis_disp_err_flag|en_disp_err_flag
		parameter hssi_8g_rx_pcs_wa_kchar = "dis_kchar", // dis_kchar|en_kchar
		parameter hssi_8g_rx_pcs_wa_pd = "wa_pd_10", // wa_pd_7|wa_pd_10|wa_pd_20|wa_pd_40|wa_pd_8_sw|wa_pd_8_dw|wa_pd_16_sw|wa_pd_16_dw|wa_pd_32
		parameter hssi_8g_rx_pcs_wa_pd_data = 40'b0,
		parameter hssi_8g_rx_pcs_wa_pd_polarity = "dis_pd_both_pol", // dis_pd_both_pol|en_pd_both_pol|dont_care_both_pol
		parameter hssi_8g_rx_pcs_wa_pld_controlled = "dis_pld_ctrl", // dis_pld_ctrl|pld_ctrl_sw|rising_edge_sensitive_dw|level_sensitive_dw
		parameter hssi_8g_rx_pcs_wa_renumber_data = 6'b0,
		parameter hssi_8g_rx_pcs_wa_rgnumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rknumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rosnumber_data = 2'b0,
		parameter hssi_8g_rx_pcs_wa_rvnumber_data = 13'b0,
		parameter hssi_8g_rx_pcs_wa_sync_sm_ctrl = "gige_sync_sm", // gige_sync_sm|pipe_sync_sm|sw_basic_sync_sm|dw_basic_sync_sm|fibre_channel_sync_sm
		parameter hssi_8g_rx_pcs_wait_cnt = 12'b0,
		
		// parameters for twentynm_hssi_8g_tx_pcs
		parameter hssi_8g_tx_pcs_auto_speed_nego_gen2 = "dis_asn_g2", // dis_asn_g2|en_asn_g2_freq_scal
		parameter hssi_8g_tx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_tx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_tx_pcs_byte_serializer = "dis_bs", // dis_bs|en_bs_by_2|en_bs_by_4
		parameter hssi_8g_tx_pcs_clock_gate_bs_enc = "dis_bs_enc_clk_gating", // dis_bs_enc_clk_gating|en_bs_enc_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_dw_fifowr = "dis_dw_fifowr_clk_gating", // dis_dw_fifowr_clk_gating|en_dw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_fiford = "dis_fiford_clk_gating", // dis_fiford_clk_gating|en_fiford_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_sw_fifowr = "dis_sw_fifowr_clk_gating", // dis_sw_fifowr_clk_gating|en_sw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_observation_in_pld_core = "internal_refclk_b", // internal_refclk_b|internal_fifo_rd_clk|internal_sw_fifo_wr_clk|internal_dw_fifo_wr_clk|internal_tx_clk_out_gen3|internal_pipe_tx_clk_out_gen3
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_tx_pcs_data_selection_8b10b_encoder_input = "normal_data_path", // normal_data_path|gige_idle_conversion
		parameter hssi_8g_tx_pcs_dynamic_clk_switch = "dis_dyn_clk_switch", // dis_dyn_clk_switch|en_dyn_clk_switch
		parameter hssi_8g_tx_pcs_eightb_tenb_disp_ctrl = "dis_disp_ctrl", // dis_disp_ctrl|en_disp_ctrl|en_ib_disp_ctrl
		parameter hssi_8g_tx_pcs_eightb_tenb_encoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_tx_pcs_force_echar = "dis_force_echar", // dis_force_echar|en_force_echar
		parameter hssi_8g_tx_pcs_force_kchar = "dis_force_kchar", // dis_force_kchar|en_force_kchar
		parameter hssi_8g_tx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // dis_tx_clk|tx_pma_clk
		parameter hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel = "func_clk", // dis_tx_pipe_clk|func_clk
		parameter hssi_8g_tx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_tx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_tx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_tx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_tx_pcs_phfifo_write_clk_sel = "pld_tx_clk", // pld_tx_clk|tx_clk
		parameter hssi_8g_tx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_tx_pcs_prot_mode = "basic", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic|disabled_prot_mode
		parameter hssi_8g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_tx_pcs_refclk_b_clk_sel = "tx_pma_clock", // tx_pma_clock|refclk_dig
		parameter hssi_8g_tx_pcs_revloop_back_rm = "dis_rev_loopback_rx_rm", // dis_rev_loopback_rx_rm|en_rev_loopback_rx_rm
		parameter hssi_8g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_tx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_tx_pcs_tx_bitslip = "dis_tx_bitslip", // dis_tx_bitslip|en_tx_bitslip
		parameter hssi_8g_tx_pcs_tx_compliance_controlled_disparity = "dis_txcompliance", // dis_txcompliance|en_txcompliance_pipe2p0|en_txcompliance_pipe3p0
		parameter hssi_8g_tx_pcs_tx_fast_pld_reg = "dis_tx_fast_pld_reg", // dis_tx_fast_pld_reg|en_tx_fast_pld_reg
		parameter hssi_8g_tx_pcs_txclk_freerun = "dis_freerun_tx", // dis_freerun_tx|en_freerun_tx
		parameter hssi_8g_tx_pcs_txpcs_urst = "en_txpcs_urst", // dis_txpcs_urst|en_txpcs_urst
		
		// parameters for twentynm_hssi_common_pcs_pma_interface
		parameter hssi_common_pcs_pma_interface_asn_clk_enable = "false", // false|true
		parameter hssi_common_pcs_pma_interface_asn_enable = "dis_asn", // dis_asn|en_asn
		parameter hssi_common_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|pcie_gen3
		parameter hssi_common_pcs_pma_interface_bypass_early_eios = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pcie_switch = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_ltr = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_sw_done = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_ppm_lock = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_txdetectrx = "false", // false|true
		parameter hssi_common_pcs_pma_interface_cdr_control = "en_cdr_ctrl", // dis_cdr_ctrl|en_cdr_ctrl
		parameter hssi_common_pcs_pma_interface_cid_enable = "en_cid_mode", // dis_cid_mode|en_cid_mode
		parameter hssi_common_pcs_pma_interface_cp_cons_sel = "cp_cons_default", // cp_cons_master|cp_cons_slave_abv|cp_cons_slave_blw|cp_cons_default
		parameter hssi_common_pcs_pma_interface_cp_dwn_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_cp_up_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_blw|ctrl_slave_abv
		parameter hssi_common_pcs_pma_interface_data_mask_count = 16'b100111000100,
		parameter hssi_common_pcs_pma_interface_data_mask_count_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_dft_observation_clock_selection = "dft_clk_obsrv_tx0", // dft_clk_obsrv_tx0|dft_clk_obsrv_tx1|dft_clk_obsrv_tx2|dft_clk_obsrv_tx3|dft_clk_obsrv_tx4|dft_clk_obsrv_rx|dft_clk_obsrv_hclk|dft_clk_obsrv_fref|dft_clk_obsrv_clklow|dft_clk_obsrv_asn0|dft_clk_obsrv_asn1
		parameter hssi_common_pcs_pma_interface_early_eios_counter = 8'b110010,
		parameter hssi_common_pcs_pma_interface_force_freqdet = "force_freqdet_dis", // force_freqdet_dis|force1_freqdet_en|force0_freqdet_en
		parameter hssi_common_pcs_pma_interface_free_run_clk_enable = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ignore_sigdet_g23 = "false", // false|true
		parameter hssi_common_pcs_pma_interface_pc_en_counter = 7'b110111,
		parameter hssi_common_pcs_pma_interface_pc_rst_counter = 5'b10111,
		parameter hssi_common_pcs_pma_interface_pcie_hip_mode = "hip_disable", // hip_enable|hip_disable
		parameter hssi_common_pcs_pma_interface_ph_fifo_reg_mode = "phfifo_reg_mode_dis", // phfifo_reg_mode_dis|phfifo_reg_mode_en
		parameter hssi_common_pcs_pma_interface_phfifo_flush_wait = 6'b100100,
		parameter hssi_common_pcs_pma_interface_pipe_if_g3pcs = "pipe_if_8gpcs", // pipe_if_g3pcs|pipe_if_8gpcs
		parameter hssi_common_pcs_pma_interface_pma_done_counter = 18'b101010101110011000,
		parameter hssi_common_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_common_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_common_pcs_pma_interface_ppm_cnt_rst = "ppm_cnt_rst_dis", // ppm_cnt_rst_dis|ppm_cnt_rst_en
		parameter hssi_common_pcs_pma_interface_ppm_deassert_early = "deassert_early_dis", // deassert_early_dis|deassert_early_en
		parameter hssi_common_pcs_pma_interface_ppm_det_buckets = "ppm_100_bucket", // disable_prot|ppm_300_bucket|ppm_100_bucket|ppm_300_100_bucket
		parameter hssi_common_pcs_pma_interface_ppm_gen1_2_cnt = "cnt_32k", // cnt_32k|cnt_64k
		parameter hssi_common_pcs_pma_interface_ppm_post_eidle_delay = "cnt_200_cycles", // cnt_200_cycles|cnt_400_cycles
		parameter hssi_common_pcs_pma_interface_ppmsel = "ppmsel_300", // ppmsel_disable|ppmsel_5000|ppmsel_2500|ppmsel_1000|ppmsel_500|ppmsel_300|ppmsel_250|ppmsel_200|ppmsel_125|ppmsel_100|ppmsel_62p5|ppm_other
		parameter hssi_common_pcs_pma_interface_prot_mode = "disable_prot_mode", // disable_prot_mode|pipe_g12|pipe_g3|other_protocols
		parameter hssi_common_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_common_pcs_pma_interface_rxvalid_mask = "rxvalid_mask_en", // rxvalid_mask_dis|rxvalid_mask_en
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter = 12'b100111000100,
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_sim_mode = "disable", // disable|enable
		parameter hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en = "true", // false|true
		parameter hssi_common_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_common_pcs_pma_interface_testout_sel = "ppm_det_test", // ppm_det_test|asn_test|pma_pll_test|rxpmaif_test|prbs_gen_test|prbs_ver_test|uhsif_1_test|uhsif_2_test|uhsif_3_test
		parameter hssi_common_pcs_pma_interface_wait_clk_on_off_timer = 4'b100,
		parameter hssi_common_pcs_pma_interface_wait_pipe_synchronizing = 5'b10111,
		parameter hssi_common_pcs_pma_interface_wait_send_syncp_fbkp = 11'b11111010,
		
		// parameters for twentynm_hssi_common_pld_pcs_interface
		parameter hssi_common_pld_pcs_interface_dft_clk_out_en = "dft_clk_out_disable", // dft_clk_out_disable|dft_clk_out_enable
		parameter hssi_common_pld_pcs_interface_dft_clk_out_sel = "teng_rx_dft_clk", // teng_rx_dft_clk|teng_tx_dft_clk|eightg_rx_dft_clk|eightg_tx_dft_clk|pmaif_dft_clk
		parameter hssi_common_pld_pcs_interface_hrdrstctrl_en = "hrst_dis", // hrst_dis|hrst_en
		parameter hssi_common_pld_pcs_interface_pcs_testbus_block_sel = "eightg", // eightg|g3pcs|teng|krfec|pma_if
		parameter hssi_common_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_fifo_rx_pcs
		parameter hssi_fifo_rx_pcs_double_read_mode = "double_read_dis", // double_read_en|double_read_dis
		parameter hssi_fifo_rx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_fifo_tx_pcs
		parameter hssi_fifo_tx_pcs_double_write_mode = "double_write_dis", // double_write_en|double_write_dis
		parameter hssi_fifo_tx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_gen3_rx_pcs
		parameter hssi_gen3_rx_pcs_block_sync = "enable_block_sync", // bypass_block_sync|enable_block_sync
		parameter hssi_gen3_rx_pcs_block_sync_sm = "enable_blk_sync_sm", // disable_blk_sync_sm|enable_blk_sync_sm
		parameter hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn = "enable", // disable|enable
		parameter hssi_gen3_rx_pcs_lpbk_force = "lpbk_frce_dis", // lpbk_frce_dis|lpbk_frce_en
		parameter hssi_gen3_rx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_rx_pcs_rate_match_fifo = "enable_rm_fifo_600ppm", // bypass_rm_fifo|enable_rm_fifo_600ppm|enable_rm_fifo_0ppm
		parameter hssi_gen3_rx_pcs_rate_match_fifo_latency = "regular_latency", // regular_latency|low_latency
		parameter hssi_gen3_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_gen3_rx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_b4gb_par_lpbk = "b4gb_par_lpbk_dis", // b4gb_par_lpbk_dis|b4gb_par_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_force_balign = "en_force_balign", // en_force_balign|dis_force_balign
		parameter hssi_gen3_rx_pcs_rx_ins_del_one_skip = "ins_del_one_skip_en", // ins_del_one_skip_dis|ins_del_one_skip_en
		parameter hssi_gen3_rx_pcs_rx_num_fixed_pat = 4'b1000,
		parameter hssi_gen3_rx_pcs_rx_test_out_sel = "rx_test_out0", // rx_test_out0|rx_test_out1
		parameter hssi_gen3_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_gen3_tx_pcs
		parameter hssi_gen3_tx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_tx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_gen3_tx_pcs_tx_bitslip = 5'b0,
		parameter hssi_gen3_tx_pcs_tx_gbox_byp = "bypass_gbox", // bypass_gbox|enable_gbox
		
		// parameters for twentynm_hssi_krfec_rx_pcs
		parameter hssi_krfec_rx_pcs_blksync_cor_en = "detect", // detect|correct
		parameter hssi_krfec_rx_pcs_bypass_gb = "bypass_dis", // bypass_dis|bypass_en
		parameter hssi_krfec_rx_pcs_clr_ctrl = "both_enabled", // both_enabled|corr_cnt_only|uncorr_cnt_only
		parameter hssi_krfec_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_rx_pcs_dv_start = "with_blklock", // with_blksync|with_blklock
		parameter hssi_krfec_rx_pcs_err_mark_type = "err_mark_10g", // err_mark_10g|err_mark_40g
		parameter hssi_krfec_rx_pcs_error_marking_en = "err_mark_dis", // err_mark_dis|err_mark_en
		parameter hssi_krfec_rx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_krfec_rx_pcs_parity_invalid_enum = 8'b1000,
		parameter hssi_krfec_rx_pcs_parity_valid_num = 4'b100,
		parameter hssi_krfec_rx_pcs_pipeln_blksync = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_descrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errcorrect = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_ind = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_lfsr = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_loc = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_pat = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_gearbox = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_syndrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_trans_dec = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_rx_pcs_receive_order = "receive_lsb", // receive_lsb|receive_msb
		parameter hssi_krfec_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_krfec_rx_pcs_rx_testbus_sel = "overall", // overall|fast_search|fast_search_cntrs|blksync|blksync_cntrs|decoder_master_sm|decoder_master_sm_cntrs|syndrm_sm|syndrm1|syndrm2|errtrap_sm|errtrap_ind1|errtrap_ind2|errtrap_ind3|errtrap_ind4|errtrap_ind5|errtrap_loc|errtrap_pat1|errtrap_pat2|errtrap_pat3|errtrap_pat4|decoder_rd_sm|gb_and_trans
		parameter hssi_krfec_rx_pcs_signal_ok_en = "sig_ok_dis", // sig_ok_dis|sig_ok_en
		parameter hssi_krfec_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_krfec_tx_pcs
		parameter hssi_krfec_tx_pcs_burst_err = "burst_err_dis", // burst_err_dis|burst_err_en
		parameter hssi_krfec_tx_pcs_burst_err_len = "burst_err_len1", // burst_err_len1|burst_err_len2|burst_err_len3|burst_err_len4|burst_err_len5|burst_err_len6|burst_err_len7|burst_err_len8|burst_err_len9|burst_err_len10|burst_err_len11|burst_err_len12|burst_err_len13|burst_err_len14|burst_err_len15|burst_err_len16
		parameter hssi_krfec_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_tx_pcs_enc_frame_query = "enc_query_dis", // enc_query_dis|enc_query_en
		parameter hssi_krfec_tx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_encoder = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_scrambler = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_krfec_tx_pcs_transcode_err = "trans_err_dis", // trans_err_dis|trans_err_en
		parameter hssi_krfec_tx_pcs_transmit_order = "transmit_lsb", // transmit_lsb|transmit_msb
		parameter hssi_krfec_tx_pcs_tx_testbus_sel = "overall", // overall|encoder1|encoder2|scramble1|scramble2|scramble3|gearbox
		
		// parameters for twentynm_hssi_pipe_gen1_2
		parameter hssi_pipe_gen1_2_elec_idle_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_error_replace_pad = "replace_edb", // replace_edb|replace_pad
		parameter hssi_pipe_gen1_2_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_pipe_gen1_2_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen1_2_phystatus_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_phystatus_rst_toggle = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen1_2_pipe_byte_de_serializer_en = "dont_care_bds", // dis_bds|en_bds_by_2|dont_care_bds
		parameter hssi_pipe_gen1_2_prot_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|basic|disabled_prot_mode
		parameter hssi_pipe_gen1_2_reconfig_settings = "{}", // 
		parameter hssi_pipe_gen1_2_rx_pipe_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_pipe_gen1_2_rxdetect_bypass = "dis_rxdetect_bypass", // dis_rxdetect_bypass|en_rxdetect_bypass
		parameter hssi_pipe_gen1_2_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen1_2_tx_pipe_enable = "dis_pipe_tx", // dis_pipe_tx|en_pipe_tx|en_pipe3_tx
		parameter hssi_pipe_gen1_2_txswing = "dis_txswing", // dis_txswing|en_txswing
		
		// parameters for twentynm_hssi_pipe_gen3
		parameter hssi_pipe_gen3_bypass_rx_detection_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_rx_preset = 3'b0,
		parameter hssi_pipe_gen3_bypass_rx_preset_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_tx_coefficent = 18'b0,
		parameter hssi_pipe_gen3_bypass_tx_coefficent_enable = "false", // false|true
		parameter hssi_pipe_gen3_elecidle_delay_g3 = 3'b110,
		parameter hssi_pipe_gen3_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen3_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|disable_pcs
		parameter hssi_pipe_gen3_phy_status_delay_g12 = 3'b101,
		parameter hssi_pipe_gen3_phy_status_delay_g3 = 3'b101,
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g12 = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g3 = "dis_phystatus_rst_toggle_g3", // dis_phystatus_rst_toggle_g3|en_phystatus_rst_toggle_g3
		parameter hssi_pipe_gen3_rate_match_pad_insertion = "dis_rm_fifo_pad_ins", // dis_rm_fifo_pad_ins|en_rm_fifo_pad_ins
		parameter hssi_pipe_gen3_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen3_test_out_sel = "disable_test_out", // tx_test_out|rx_test_out|pipe_test_out1|pipe_test_out2|pipe_test_out3|pipe_ctrl_test_out|disable_test_out
		
		// parameters for twentynm_hssi_rx_pcs_pma_interface
		parameter hssi_rx_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|ten_g_pcs|direct_pld
		parameter hssi_rx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pcs_pma_interface_clkslip_sel = "pld", // pld|slip_eight_g_pcs
		parameter hssi_rx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pcs_pma_interface_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_rx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_rx_pcs_pma_interface_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_rx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_rx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_rx_pcs_pma_interface_prbs_ver = "prbs_off", // prbs_off|prbs_31|prbs_15|prbs_23|prbs_9|prbs_7
		parameter hssi_rx_pcs_pma_interface_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion = "rx_dyn_polinv_dis", // rx_dyn_polinv_dis|rx_dyn_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_lpbk_en = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok = "unforce_sig_ok", // unforce_sig_ok|force_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mask = "prbsmask128", // prbsmask128|prbsmask256|prbsmask512|prbsmask1024
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mode = "teng_mode", // teng_mode|eightg_mode
		parameter hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel = "sel_sig_det", // sel_sig_det|sel_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_static_polarity_inversion = "rx_stat_polinv_dis", // rx_stat_polinv_dis|rx_stat_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en = "uhsif_lpbk_dis", // uhsif_lpbk_dis|uhsif_lpbk_en
		parameter hssi_rx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_rx_pld_pcs_interface
		parameter hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx = "enable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx = "pma_64b_rx", // pma_32b_rx|pma_40b_rx|pma_64b_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_baser_mode_rx|interlaken_mode_rx|sfis_mode_rx|teng_sdi_mode_rx|basic_mode_rx|test_prp_mode_rx|test_prp_krfec_mode_rx|teng_1588_mode_rx|teng_baser_krfec_mode_rx|teng_1588_krfec_mode_rx|basic_krfec_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx = "disabled_prot_mode_rx", // pipe_g1_rx|pipe_g2_rx|pipe_g3_rx|cpri_rx|cpri_rx_tx_rx|gige_rx|gige_1588_rx|basic_rm_enable_rx|basic_rm_disable_rx|disabled_prot_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcie_g1_capable_rx|pcie_g2_capable_rx|pcie_g3_capable_rx|gige_rx|teng_baser_rx|teng_basekr_krfec_rx|fortyg_basekr_krfec_rx|cpri_8b10b_rx|interlaken_rx|sfis_rx|teng_sdi_rx|gige_1588_rx|teng_1588_baser_rx|teng_1588_basekr_krfec_rx|basic_8gpcs_rm_enable_rx|basic_8gpcs_rm_disable_rx|basic_10gpcs_rx|basic_10gpcs_krfec_rx|pcs_direct_rx|prp_rx|prp_krfec_rx|prbs_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx = "teng_mode_rx", // teng_mode_rx|non_teng_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_basekr_mode_rx|fortyg_basekr_mode_rx|teng_1588_basekr_mode_rx|basic_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|eightg_and_g3_pld_fifo_mode_rx|eightg_and_g3_reg_mode_rx|eightg_and_g3_reg_mode_hip_rx|teng_pld_fifo_mode_rx|teng_reg_mode_rx|teng_and_krfec_pld_fifo_mode_rx|teng_and_krfec_reg_mode_rx|pcs_direct_reg_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_block_sel = "pcs_direct", // eightg|teng|pcs_direct
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_rx_clk|pma_rx_clk_user
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_sel = "pld_rx_clk", // pld_rx_clk|pcs_rx_clk
		parameter hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en = "hip_rx_enable", // hip_rx_enable|hip_rx_disable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_rx_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_tx_pcs_pma_interface
		parameter hssi_tx_pcs_pma_interface_bypass_pma_txelecidle = "false", // false|true
		parameter hssi_tx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pcs_pma_interface_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx = "other_prot_mode", // pipe_g12|pipe_g3|other_prot_mode
		parameter hssi_tx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_tx_pcs_pma_interface_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_tx_pcs_pma_interface_pmagate_en = "pmagate_dis", // pmagate_dis|pmagate_en
		parameter hssi_tx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_tx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_tx_pcs_pma_interface_prbs_gen_pat = "prbs_gen_dis", // prbs_gen_dis|prbs_31|prbs_23|prbs_15|prbs_9|prbs_7
		parameter hssi_tx_pcs_pma_interface_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_tx_pcs_pma_interface_sq_wave_num = "sq_wave_4", // sq_wave_1|sq_wave_4|sq_wave_8|sq_wave_6|sq_wave_default
		parameter hssi_tx_pcs_pma_interface_sqwgen_clken = "sqwgen_clk_dis", // sqwgen_clk_dis|sqwgen_clk_en
		parameter hssi_tx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion = "tx_dyn_polinv_dis", // tx_dyn_polinv_dis|tx_dyn_polinv_en
		parameter hssi_tx_pcs_pma_interface_tx_pma_data_sel = "pld_dir", // pld_dir|pcie_gen3|eight_g_pcs|ten_g_pcs|prbs_pat|sq_wave_pat|block_sel_default|registered_uhsif_dat|directed_uhsif_dat
		parameter hssi_tx_pcs_pma_interface_tx_static_polarity_inversion = "tx_stat_polinv_dis", // tx_stat_polinv_dis|tx_stat_polinv_en
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock = "uhsif_filt_stepsz_b4lock_4", // uhsif_filt_stepsz_b4lock_2|uhsif_filt_stepsz_b4lock_4|uhsif_filt_stepsz_b4lock_6|uhsif_filt_stepsz_b4lock_8
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value = 4'b1011,
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock = "uhsif_filt_cntthr_b4lock_16", // uhsif_filt_cntthr_b4lock_8|uhsif_filt_cntthr_b4lock_16|uhsif_filt_cntthr_b4lock_24|uhsif_filt_cntthr_b4lock_32
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period = "uhsif_dcn_test_period_4", // uhsif_dcn_test_period_4|uhsif_dcn_test_period_8|uhsif_dcn_test_period_12|uhsif_dcn_test_period_16
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable = "uhsif_dcn_test_mode_disable", // uhsif_dcn_test_mode_enable|uhsif_dcn_test_mode_disable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh = "uhsif_dzt_cnt_thr_4", // uhsif_dzt_cnt_thr_2|uhsif_dzt_cnt_thr_4|uhsif_dzt_cnt_thr_6|uhsif_dzt_cnt_thr_8
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable = "uhsif_dzt_enable", // uhsif_dzt_disable|uhsif_dzt_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window = "uhsif_dzt_obr_win_32", // uhsif_dzt_obr_win_16|uhsif_dzt_obr_win_32|uhsif_dzt_obr_win_48|uhsif_dzt_obr_win_64
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size = "uhsif_dzt_skipsz_8", // uhsif_dzt_skipsz_4|uhsif_dzt_skipsz_8|uhsif_dzt_skipsz_12|uhsif_dzt_skipsz_16
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel = "uhsif_index_internal", // uhsif_index_internal|uhsif_index_cram
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin = "uhsif_dcn_margin_4", // uhsif_dcn_margin_2|uhsif_dcn_margin_3|uhsif_dcn_margin_4|uhsif_dcn_margin_5
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value = 8'b10000000,
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control = "uhsif_dft_dz_det_val_0", // uhsif_dft_dz_det_val_0|uhsif_dft_dz_det_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control = "uhsif_dft_up_val_0", // uhsif_dft_up_val_0|uhsif_dft_up_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_enable = "uhsif_disable", // uhsif_disable|uhsif_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock = "uhsif_lkd_segsz_aflock_2048", // uhsif_lkd_segsz_aflock_512|uhsif_lkd_segsz_aflock_1024|uhsif_lkd_segsz_aflock_2048|uhsif_lkd_segsz_aflock_4096
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock = "uhsif_lkd_segsz_b4lock_32", // uhsif_lkd_segsz_b4lock_16|uhsif_lkd_segsz_b4lock_32|uhsif_lkd_segsz_b4lock_64|uhsif_lkd_segsz_b4lock_128
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value = 4'b11,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value = 4'b11,
		
		// parameters for twentynm_hssi_tx_pld_pcs_interface
		parameter hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx = "enable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx = "pma_64b_tx", // pma_32b_tx|pma_40b_tx|pma_64b_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_baser_mode_tx|interlaken_mode_tx|sfis_mode_tx|teng_sdi_mode_tx|basic_mode_tx|test_prp_mode_tx|test_prp_krfec_mode_tx|teng_1588_mode_tx|teng_baser_krfec_mode_tx|teng_1588_krfec_mode_tx|basic_krfec_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx = "disabled_prot_mode_tx", // pipe_g1_tx|pipe_g2_tx|pipe_g3_tx|cpri_tx|cpri_rx_tx_tx|gige_tx|gige_1588_tx|basic_tx|disabled_prot_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcie_g1_capable_tx|pcie_g2_capable_tx|pcie_g3_capable_tx|gige_tx|teng_baser_tx|teng_basekr_krfec_tx|fortyg_basekr_krfec_tx|cpri_8b10b_tx|interlaken_tx|sfis_tx|teng_sdi_tx|gige_1588_tx|teng_1588_baser_tx|teng_1588_basekr_krfec_tx|basic_8gpcs_tx|basic_10gpcs_tx|basic_10gpcs_krfec_tx|pcs_direct_tx|uhsif_tx|prp_tx|prp_krfec_tx|prbs_tx|sqwave_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx = "teng_mode_tx", // teng_mode_tx|non_teng_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_basekr_mode_tx|fortyg_basekr_mode_tx|teng_1588_basekr_mode_tx|basic_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|eightg_and_g3_pld_fifo_mode_tx|eightg_and_g3_reg_mode_tx|eightg_and_g3_reg_mode_hip_tx|eightg_and_g3_fastreg_mode_tx|teng_pld_fifo_mode_tx|teng_reg_mode_tx|teng_fastreg_mode_tx|teng_and_krfec_pld_fifo_mode_tx|teng_and_krfec_reg_mode_tx|teng_and_krfec_fastreg_mode_tx|pcs_direct_fastreg_mode_tx|uhsif_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_tx_clk|pma_tx_clk_user
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_source = "teng", // eightg|teng|pma_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_data_source = "hip_disable", // hip_disable|hip_enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en = "delay1_clk_disable", // delay1_clk_enable|delay1_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel = "pld_tx_clk", // pld_tx_clk|pcs_tx_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl = "delay1_path0", // delay1_path0|delay1_path1|delay1_path2|delay1_path3|delay1_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel = "one_ff_delay", // one_ff_delay|two_ff_delay
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en = "delay2_clk_disable", // delay2_clk_enable|delay2_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl = "delay2_path0", // delay2_path0|delay2_path1|delay2_path2|delay2_path3|delay2_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_tx_pld_pcs_interface_reconfig_settings = "{}" // 
	//PARAM_LIST_END
	)
	(
	//PORT_LIST_START
		input wire	[8:0]	in_avmmaddress,
		input wire		in_avmmclk,
		input wire		in_avmmread,
		input wire		in_avmmrstn,
		input wire		in_avmmwrite,
		input wire	[7:0]	in_avmmwritedata,
		input wire	[4:0]	in_bond_pcs10g_in_bot,
		input wire	[4:0]	in_bond_pcs10g_in_top,
		input wire	[12:0]	in_bond_pcs8g_in_bot,
		input wire	[12:0]	in_bond_pcs8g_in_top,
		input wire	[11:0]	in_bond_pmaif_in_bot,
		input wire	[11:0]	in_bond_pmaif_in_top,
		input wire	[63:0]	in_hip_tx_data,
		input wire		in_iocsr_clk,
		input wire	[5:0]	in_iocsr_config,
		input wire		in_iocsr_rdy,
		input wire		in_iocsr_rdy_dly,
		input wire		in_pld_10g_krfec_rx_clr_errblk_cnt,
		input wire		in_pld_10g_krfec_rx_pld_rst_n,
		input wire		in_pld_10g_krfec_tx_pld_rst_n,
		input wire		in_pld_10g_rx_align_clr,
		input wire		in_pld_10g_rx_clr_ber_count,
		input wire		in_pld_10g_rx_rd_en,
		input wire	[6:0]	in_pld_10g_tx_bitslip,
		input wire		in_pld_10g_tx_burst_en,
		input wire		in_pld_10g_tx_data_valid,
		input wire	[1:0]	in_pld_10g_tx_diag_status,
		input wire		in_pld_10g_tx_wordslip,
		input wire		in_pld_8g_a1a2_size,
		input wire		in_pld_8g_bitloc_rev_en,
		input wire		in_pld_8g_byte_rev_en,
		input wire	[2:0]	in_pld_8g_eidleinfersel,
		input wire		in_pld_8g_encdt,
		input wire		in_pld_8g_g3_rx_pld_rst_n,
		input wire		in_pld_8g_g3_tx_pld_rst_n,
		input wire		in_pld_8g_rddisable_tx,
		input wire		in_pld_8g_rdenable_rx,
		input wire		in_pld_8g_refclk_dig2,
		input wire		in_pld_8g_rxpolarity,
		input wire	[4:0]	in_pld_8g_tx_boundary_sel,
		input wire		in_pld_8g_wrdisable_rx,
		input wire		in_pld_8g_wrenable_tx,
		input wire		in_pld_atpg_los_en_n,
		input wire		in_pld_bitslip,
		input wire	[17:0]	in_pld_g3_current_coeff,
		input wire	[2:0]	in_pld_g3_current_rxpreset,
		input wire		in_pld_ltr,
		input wire		in_pld_mem_krfec_atpg_rst_n,
		input wire		in_pld_partial_reconfig,
		input wire		in_pld_pcs_refclk_dig,
		input wire		in_pld_pma_adapt_start,
		input wire		in_pld_pma_csr_test_dis,
		input wire		in_pld_pma_early_eios,
		input wire	[5:0]	in_pld_pma_eye_monitor,
		input wire		in_pld_pma_ltd_b,
		input wire		in_pld_pma_nrpi_freeze,
		input wire	[1:0]	in_pld_pma_pcie_switch,
		input wire		in_pld_pma_ppm_lock,
		input wire	[4:0]	in_pld_pma_reserved_out,
		input wire		in_pld_pma_rs_lpbk_b,
		input wire		in_pld_pma_rx_qpi_pullup,
		input wire		in_pld_pma_rxpma_rstb,
		input wire		in_pld_pma_tx_bitslip,
		input wire		in_pld_pma_tx_bonding_rstb,
		input wire		in_pld_pma_tx_qpi_pulldn,
		input wire		in_pld_pma_tx_qpi_pullup,
		input wire		in_pld_pma_txdetectrx,
		input wire		in_pld_pma_txpma_rstb,
		input wire		in_pld_pmaif_rx_pld_rst_n,
		input wire		in_pld_pmaif_rxclkslip,
		input wire		in_pld_pmaif_tx_pld_rst_n,
		input wire		in_pld_polinv_rx,
		input wire		in_pld_polinv_tx,
		input wire	[1:0]	in_pld_rate,
		input wire	[9:0]	in_pld_reserved_in,
		input wire		in_pld_rx_clk,
		input wire		in_pld_rx_prbs_err_clr,
		input wire		in_pld_scan_mode_n,
		input wire		in_pld_scan_shift_n,
		input wire		in_pld_syncsm_en,
		input wire		in_pld_tx_clk,
		input wire	[17:0]	in_pld_tx_control,
		input wire	[127:0]	in_pld_tx_data,
		input wire		in_pld_txelecidle,
		input wire		in_pld_uhsif_tx_clk,
		input wire		in_pma_adapt_done,
		input wire		in_pma_clklow,
		input wire		in_pma_fref,
		input wire		in_pma_hclk,
		input wire	[1:0]	in_pma_pcie_sw_done,
		input wire		in_pma_pfdmode_lock,
		input wire	[4:0]	in_pma_reserved_in,
		input wire		in_pma_rx_clkdiv_user,
		input wire		in_pma_rx_detect_valid,
		input wire		in_pma_rx_found,
		input wire		in_pma_rx_pma_clk,
		input wire	[63:0]	in_pma_rx_pma_data,
		input wire		in_pma_rx_signal_ok,
		input wire		in_pma_rxpll_lock,
		input wire		in_pma_signal_det,
		input wire	[7:0]	in_pma_testbus,
		input wire		in_pma_tx_clkdiv_user,
		input wire		in_pma_tx_pma_clk,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen1_2,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen3,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pld_pcs_interface,
		output wire		out_blockselect_hssi_10g_rx_pcs,
		output wire		out_blockselect_hssi_10g_tx_pcs,
		output wire		out_blockselect_hssi_8g_rx_pcs,
		output wire		out_blockselect_hssi_8g_tx_pcs,
		output wire		out_blockselect_hssi_common_pcs_pma_interface,
		output wire		out_blockselect_hssi_common_pld_pcs_interface,
		output wire		out_blockselect_hssi_fifo_rx_pcs,
		output wire		out_blockselect_hssi_fifo_tx_pcs,
		output wire		out_blockselect_hssi_gen3_rx_pcs,
		output wire		out_blockselect_hssi_gen3_tx_pcs,
		output wire		out_blockselect_hssi_krfec_rx_pcs,
		output wire		out_blockselect_hssi_krfec_tx_pcs,
		output wire		out_blockselect_hssi_pipe_gen1_2,
		output wire		out_blockselect_hssi_pipe_gen3,
		output wire		out_blockselect_hssi_rx_pcs_pma_interface,
		output wire		out_blockselect_hssi_rx_pld_pcs_interface,
		output wire		out_blockselect_hssi_tx_pcs_pma_interface,
		output wire		out_blockselect_hssi_tx_pld_pcs_interface,
		output wire	[4:0]	out_bond_pcs10g_out_bot,
		output wire	[4:0]	out_bond_pcs10g_out_top,
		output wire	[12:0]	out_bond_pcs8g_out_bot,
		output wire	[12:0]	out_bond_pcs8g_out_top,
		output wire	[11:0]	out_bond_pmaif_out_bot,
		output wire	[11:0]	out_bond_pmaif_out_top,
		output wire	[2:0]	out_hip_clk_out,
		output wire	[7:0]	out_hip_ctrl_out,
		output wire		out_hip_iocsr_rdy,
		output wire		out_hip_iocsr_rdy_dly,
		output wire		out_hip_nfrzdrv,
		output wire		out_hip_npor,
		output wire	[50:0]	out_hip_rx_data,
		output wire		out_hip_usermode,
		output wire		out_pld_10g_krfec_rx_blk_lock,
		output wire	[1:0]	out_pld_10g_krfec_rx_diag_data_status,
		output wire		out_pld_10g_krfec_rx_frame,
		output wire		out_pld_10g_krfec_tx_frame,
		output wire		out_pld_10g_rx_align_val,
		output wire		out_pld_10g_rx_crc32_err,
		output wire		out_pld_10g_rx_data_valid,
		output wire		out_pld_10g_rx_empty,
		output wire		out_pld_10g_rx_fifo_del,
		output wire		out_pld_10g_rx_fifo_insert,
		output wire	[4:0]	out_pld_10g_rx_fifo_num,
		output wire		out_pld_10g_rx_frame_lock,
		output wire		out_pld_10g_rx_hi_ber,
		output wire		out_pld_10g_rx_oflw_err,
		output wire		out_pld_10g_rx_pempty,
		output wire		out_pld_10g_rx_pfull,
		output wire		out_pld_10g_tx_burst_en_exe,
		output wire		out_pld_10g_tx_empty,
		output wire	[3:0]	out_pld_10g_tx_fifo_num,
		output wire		out_pld_10g_tx_full,
		output wire		out_pld_10g_tx_pempty,
		output wire		out_pld_10g_tx_pfull,
		output wire		out_pld_10g_tx_wordslip_exe,
		output wire	[3:0]	out_pld_8g_a1a2_k1k2_flag,
		output wire		out_pld_8g_empty_rmf,
		output wire		out_pld_8g_empty_rx,
		output wire		out_pld_8g_empty_tx,
		output wire		out_pld_8g_full_rmf,
		output wire		out_pld_8g_full_rx,
		output wire		out_pld_8g_full_tx,
		output wire		out_pld_8g_rxelecidle,
		output wire		out_pld_8g_signal_detect_out,
		output wire	[4:0]	out_pld_8g_wa_boundary,
		output wire		out_pld_krfec_tx_alignment,
		output wire		out_pld_pcs_rx_clk_out,
		output wire		out_pld_pcs_tx_clk_out,
		output wire		out_pld_pma_adapt_done,
		output wire		out_pld_pma_clkdiv_rx_user,
		output wire		out_pld_pma_clkdiv_tx_user,
		output wire		out_pld_pma_clklow,
		output wire		out_pld_pma_fref,
		output wire		out_pld_pma_hclk,
		output wire	[1:0]	out_pld_pma_pcie_sw_done,
		output wire		out_pld_pma_pfdmode_lock,
		output wire	[4:0]	out_pld_pma_reserved_in,
		output wire		out_pld_pma_rx_clk_out,
		output wire		out_pld_pma_rx_detect_valid,
		output wire		out_pld_pma_rx_found,
		output wire		out_pld_pma_rxpll_lock,
		output wire		out_pld_pma_signal_ok,
		output wire	[7:0]	out_pld_pma_testbus,
		output wire		out_pld_pma_tx_clk_out,
		output wire		out_pld_pmaif_mask_tx_pll,
		output wire	[9:0]	out_pld_reserved_out,
		output wire	[19:0]	out_pld_rx_control,
		output wire	[127:0]	out_pld_rx_data,
		output wire		out_pld_rx_prbs_done,
		output wire		out_pld_rx_prbs_err,
		output wire	[19:0]	out_pld_test_data,
		output wire		out_pld_uhsif_lock,
		output wire		out_pld_uhsif_tx_clk_out,
		output wire		out_pma_adapt_start,
		output wire		out_pma_atpg_los_en_n,
		output wire		out_pma_csr_test_dis,
		output wire	[17:0]	out_pma_current_coeff,
		output wire	[2:0]	out_pma_current_rxpreset,
		output wire		out_pma_early_eios,
		output wire	[5:0]	out_pma_eye_monitor,
		output wire	[1:0]	out_pma_interface_select,
		output wire		out_pma_ltd_b,
		output wire		out_pma_ltr,
		output wire		out_pma_nfrzdrv,
		output wire		out_pma_nrpi_freeze,
		output wire	[1:0]	out_pma_pcie_switch,
		output wire		out_pma_ppm_lock,
		output wire	[4:0]	out_pma_reserved_out,
		output wire		out_pma_rs_lpbk_b,
		output wire		out_pma_rx_clkslip,
		output wire		out_pma_rx_qpi_pullup,
		output wire		out_pma_rxpma_rstb,
		output wire		out_pma_scan_mode_n,
		output wire		out_pma_scan_shift_n,
		output wire		out_pma_tx_bitslip,
		output wire		out_pma_tx_bonding_rstb,
		output wire		out_pma_tx_elec_idle,
		output wire	[63:0]	out_pma_tx_pma_data,
		output wire		out_pma_tx_qpi_pulldn,
		output wire		out_pma_tx_qpi_pullup,
		output wire		out_pma_tx_txdetectrx,
		output wire		out_pma_txpma_rstb
	//PORT_LIST_END
	);
	//wire declarations
	
	// wires for module twentynm_hssi_fifo_tx_pcs
	wire	[7:0]	w_hssi_fifo_tx_pcs_avmmreaddata;
	wire		w_hssi_fifo_tx_pcs_blockselect;
	wire	[72:0]	w_hssi_fifo_tx_pcs_data_out_10g;
	wire	[63:0]	w_hssi_fifo_tx_pcs_data_out_8g_phase_comp;
	
	// wires for module twentynm_hssi_gen3_rx_pcs
	wire	[7:0]	w_hssi_gen3_rx_pcs_avmmreaddata;
	wire		w_hssi_gen3_rx_pcs_blk_algnd_int;
	wire		w_hssi_gen3_rx_pcs_blk_start;
	wire		w_hssi_gen3_rx_pcs_blockselect;
	wire		w_hssi_gen3_rx_pcs_clkcomp_delete_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_insert_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_overfl_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_undfl_int;
	wire	[31:0]	w_hssi_gen3_rx_pcs_data_out;
	wire		w_hssi_gen3_rx_pcs_data_valid;
	wire		w_hssi_gen3_rx_pcs_ei_det_int;
	wire		w_hssi_gen3_rx_pcs_ei_partial_det_int;
	wire		w_hssi_gen3_rx_pcs_err_decode_int;
	wire		w_hssi_gen3_rx_pcs_i_det_int;
	wire		w_hssi_gen3_rx_pcs_lpbk_blk_start;
	wire	[33:0]	w_hssi_gen3_rx_pcs_lpbk_data;
	wire		w_hssi_gen3_rx_pcs_lpbk_data_valid;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk;
	wire	[39:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n;
	wire		w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int;
	wire	[19:0]	w_hssi_gen3_rx_pcs_rx_test_out;
	wire	[1:0]	w_hssi_gen3_rx_pcs_sync_hdr;
	
	// wires for module twentynm_hssi_krfec_tx_pcs
	wire	[7:0]	w_hssi_krfec_tx_pcs_avmmreaddata;
	wire		w_hssi_krfec_tx_pcs_blockselect;
	wire		w_hssi_krfec_tx_pcs_tx_alignment;
	wire	[63:0]	w_hssi_krfec_tx_pcs_tx_data_out;
	wire		w_hssi_krfec_tx_pcs_tx_frame;
	wire	[19:0]	w_hssi_krfec_tx_pcs_tx_test_data;
	
	// wires for module twentynm_hssi_krfec_rx_pcs
	wire	[7:0]	w_hssi_krfec_rx_pcs_avmmreaddata;
	wire		w_hssi_krfec_rx_pcs_blockselect;
	wire		w_hssi_krfec_rx_pcs_rx_block_lock;
	wire	[9:0]	w_hssi_krfec_rx_pcs_rx_control_out;
	wire	[63:0]	w_hssi_krfec_rx_pcs_rx_data_out;
	wire	[1:0]	w_hssi_krfec_rx_pcs_rx_data_status;
	wire		w_hssi_krfec_rx_pcs_rx_data_valid_out;
	wire		w_hssi_krfec_rx_pcs_rx_frame;
	wire		w_hssi_krfec_rx_pcs_rx_signal_ok_out;
	
	// wires for module twentynm_hssi_rx_pld_pcs_interface
	wire	[7:0]	w_hssi_rx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_rx_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_hip_rx_ctrl;
	wire	[50:0]	w_hssi_rx_pld_pcs_interface_hip_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
	wire	[3:0]	w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary;
	wire		w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_pld_rx_control;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_pld_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
	
	// wires for module twentynm_hssi_common_pld_pcs_interface
	wire	[7:0]	w_hssi_common_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_common_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_hip_cmn_clk;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_hip_cmn_ctrl;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
	wire		w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_hip_npor;
	wire		w_hssi_common_pld_pcs_interface_hip_usermode;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n;
	wire	[17:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel;
	wire		w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_clklow;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_fref;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_hclk;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_pld_pma_reserved_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
	wire	[7:0]	w_hssi_common_pld_pcs_interface_pld_pma_testbus;
	wire		w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
	wire	[9:0]	w_hssi_common_pld_pcs_interface_pld_reserved_out;
	wire	[19:0]	w_hssi_common_pld_pcs_interface_pld_test_data;
	wire		w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
	wire		w_hssi_common_pld_pcs_interface_scan_mode_n;
	
	// wires for module twentynm_hssi_10g_rx_pcs
	wire	[7:0]	w_hssi_10g_rx_pcs_avmmreaddata;
	wire		w_hssi_10g_rx_pcs_blockselect;
	wire		w_hssi_10g_rx_pcs_rx_align_val;
	wire		w_hssi_10g_rx_pcs_rx_blk_lock;
	wire		w_hssi_10g_rx_pcs_rx_clk_out;
	wire		w_hssi_10g_rx_pcs_rx_clk_out_pld_if;
	wire	[19:0]	w_hssi_10g_rx_pcs_rx_control;
	wire		w_hssi_10g_rx_pcs_rx_crc32_err;
	wire	[127:0]	w_hssi_10g_rx_pcs_rx_data;
	wire		w_hssi_10g_rx_pcs_rx_data_valid;
	wire		w_hssi_10g_rx_pcs_rx_dft_clk_out;
	wire	[1:0]	w_hssi_10g_rx_pcs_rx_diag_status;
	wire		w_hssi_10g_rx_pcs_rx_empty;
	wire		w_hssi_10g_rx_pcs_rx_fec_clk;
	wire		w_hssi_10g_rx_pcs_rx_fifo_del;
	wire		w_hssi_10g_rx_pcs_rx_fifo_insert;
	wire	[4:0]	w_hssi_10g_rx_pcs_rx_fifo_num;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_clk;
	wire	[73:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_data;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_en;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_ptr;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_frame_lock;
	wire		w_hssi_10g_rx_pcs_rx_hi_ber;
	wire		w_hssi_10g_rx_pcs_rx_master_clk;
	wire		w_hssi_10g_rx_pcs_rx_master_clk_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_oflw_err;
	wire		w_hssi_10g_rx_pcs_rx_pempty;
	wire		w_hssi_10g_rx_pcs_rx_pfull;
	wire		w_hssi_10g_rx_pcs_rx_random_err;
	wire		w_hssi_10g_rx_pcs_rx_rx_frame;
	
	// wires for module twentynm_hssi_tx_pld_pcs_interface
	wire	[7:0]	w_hssi_tx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_tx_pld_pcs_interface_blockselect;
	wire		w_hssi_tx_pld_pcs_interface_hip_tx_clk;
	wire	[6:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en;
	wire	[17:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control;
	wire	[8:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg;
	wire	[127:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start;
	wire	[4:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle;
	wire	[2:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
	wire		w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
	
	// wires for module twentynm_hssi_tx_pcs_pma_interface
	wire	[7:0]	w_hssi_tx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_tx_pcs_pma_interface_blockselect;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out;
	wire	[4:0]	w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk;
	wire		w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_pma_tx_pma_data;
	wire		w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_1;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_2;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_3;
	
	// wires for module twentynm_hssi_rx_pcs_pma_interface
	wire	[7:0]	w_hssi_rx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_rx_pcs_pma_interface_blockselect;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni;
	wire	[31:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok;
	wire		w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk;
	wire	[5:0]	w_hssi_rx_pcs_pma_interface_pma_eye_monitor;
	wire		w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
	wire		w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test;
	
	// wires for module twentynm_hssi_10g_tx_pcs
	wire	[7:0]	w_hssi_10g_tx_pcs_avmmreaddata;
	wire		w_hssi_10g_tx_pcs_blockselect;
	wire		w_hssi_10g_tx_pcs_distdwn_out_dv;
	wire		w_hssi_10g_tx_pcs_distdwn_out_rden;
	wire		w_hssi_10g_tx_pcs_distdwn_out_wren;
	wire		w_hssi_10g_tx_pcs_distup_out_dv;
	wire		w_hssi_10g_tx_pcs_distup_out_rden;
	wire		w_hssi_10g_tx_pcs_distup_out_wren;
	wire		w_hssi_10g_tx_pcs_tx_burst_en_exe;
	wire		w_hssi_10g_tx_pcs_tx_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pma_if;
	wire	[8:0]	w_hssi_10g_tx_pcs_tx_control_out_krfec;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_data_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_data_valid_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_dft_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_empty;
	wire		w_hssi_10g_tx_pcs_tx_fec_clk;
	wire	[3:0]	w_hssi_10g_tx_pcs_tx_fifo_num;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_rd_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_clk;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_en;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_frame;
	wire		w_hssi_10g_tx_pcs_tx_full;
	wire		w_hssi_10g_tx_pcs_tx_master_clk;
	wire		w_hssi_10g_tx_pcs_tx_master_clk_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_pempty;
	wire		w_hssi_10g_tx_pcs_tx_pfull;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_data;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_gating_val;
	wire	[19:0]	w_hssi_10g_tx_pcs_tx_test_data;
	wire		w_hssi_10g_tx_pcs_tx_wordslip_exe;
	
	// wires for module twentynm_hssi_8g_tx_pcs
	wire	[7:0]	w_hssi_8g_tx_pcs_avmmreaddata;
	wire		w_hssi_8g_tx_pcs_blockselect;
	wire		w_hssi_8g_tx_pcs_clk_out;
	wire		w_hssi_8g_tx_pcs_clk_out_gen3;
	wire	[19:0]	w_hssi_8g_tx_pcs_dataout;
	wire		w_hssi_8g_tx_pcs_dyn_clk_switch_n;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn;
	wire		w_hssi_8g_tx_pcs_g3_tx_pma_rstn;
	wire	[2:0]	w_hssi_8g_tx_pcs_non_gray_eidleinfersel;
	wire		w_hssi_8g_tx_pcs_ph_fifo_overflow;
	wire		w_hssi_8g_tx_pcs_ph_fifo_underflow;
	wire		w_hssi_8g_tx_pcs_phfifo_txdeemph;
	wire	[2:0]	w_hssi_8g_tx_pcs_phfifo_txmargin;
	wire		w_hssi_8g_tx_pcs_phfifo_txswing;
	wire		w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out;
	wire	[1:0]	w_hssi_8g_tx_pcs_pipe_power_down_out;
	wire		w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3;
	wire		w_hssi_8g_tx_pcs_pmaif_asn_rstn;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_refclk_b;
	wire		w_hssi_8g_tx_pcs_refclk_b_reset;
	wire		w_hssi_8g_tx_pcs_rxpolarity_int;
	wire		w_hssi_8g_tx_pcs_soft_reset_wclk1_n;
	wire		w_hssi_8g_tx_pcs_sw_fifo_wr_clk;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_blk_start_out;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_ctrlplane_testbus;
	wire	[31:0]	w_hssi_8g_tx_pcs_tx_data_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_data_valid_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_datak_out;
	wire		w_hssi_8g_tx_pcs_tx_detect_rxloopback_int;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_tx_pipe_clk;
	wire		w_hssi_8g_tx_pcs_tx_pipe_electidle;
	wire		w_hssi_8g_tx_pcs_tx_pipe_soft_reset;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_sync_hdr_out;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_testbus;
	wire		w_hssi_8g_tx_pcs_txcompliance_out;
	wire		w_hssi_8g_tx_pcs_txelecidle_out;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk;
	wire	[63:0]	w_hssi_8g_tx_pcs_wr_data_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_en_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo;
	
	// wires for module twentynm_hssi_pipe_gen3
	wire	[7:0]	w_hssi_pipe_gen3_avmmreaddata;
	wire		w_hssi_pipe_gen3_blockselect;
	wire		w_hssi_pipe_gen3_gen3_clk_sel;
	wire		w_hssi_pipe_gen3_pcs_rst;
	wire		w_hssi_pipe_gen3_phystatus;
	wire	[17:0]	w_hssi_pipe_gen3_pma_current_coeff;
	wire	[2:0]	w_hssi_pipe_gen3_pma_current_rxpreset;
	wire		w_hssi_pipe_gen3_pma_tx_elec_idle;
	wire		w_hssi_pipe_gen3_pma_txdetectrx;
	wire		w_hssi_pipe_gen3_rev_lpbk_8gpcs_out;
	wire		w_hssi_pipe_gen3_rev_lpbk_int;
	wire	[3:0]	w_hssi_pipe_gen3_rx_blk_start;
	wire	[1:0]	w_hssi_pipe_gen3_rx_sync_hdr;
	wire	[63:0]	w_hssi_pipe_gen3_rxd_8gpcs_out;
	wire	[3:0]	w_hssi_pipe_gen3_rxdataskip;
	wire		w_hssi_pipe_gen3_rxelecidle;
	wire		w_hssi_pipe_gen3_rxpolarity_8gpcs_out;
	wire		w_hssi_pipe_gen3_rxpolarity_int;
	wire	[2:0]	w_hssi_pipe_gen3_rxstatus;
	wire		w_hssi_pipe_gen3_rxvalid;
	wire		w_hssi_pipe_gen3_shutdown_clk;
	wire	[19:0]	w_hssi_pipe_gen3_test_out;
	wire		w_hssi_pipe_gen3_tx_blk_start_int;
	wire	[1:0]	w_hssi_pipe_gen3_tx_sync_hdr_int;
	wire	[31:0]	w_hssi_pipe_gen3_txdata_int;
	wire	[3:0]	w_hssi_pipe_gen3_txdatak_int;
	wire		w_hssi_pipe_gen3_txdataskip_int;
	
	// wires for module twentynm_hssi_pipe_gen1_2
	wire	[7:0]	w_hssi_pipe_gen1_2_avmmreaddata;
	wire		w_hssi_pipe_gen1_2_blockselect;
	wire	[17:0]	w_hssi_pipe_gen1_2_current_coeff;
	wire		w_hssi_pipe_gen1_2_phystatus;
	wire		w_hssi_pipe_gen1_2_polarity_inversion_rx;
	wire		w_hssi_pipe_gen1_2_rev_loopbk;
	wire		w_hssi_pipe_gen1_2_rxelecidle;
	wire		w_hssi_pipe_gen1_2_rxelectricalidle_out;
	wire	[2:0]	w_hssi_pipe_gen1_2_rxstatus;
	wire		w_hssi_pipe_gen1_2_rxvalid;
	wire		w_hssi_pipe_gen1_2_tx_elec_idle_out;
	wire		w_hssi_pipe_gen1_2_txdetectrx;
	
	// wires for module twentynm_hssi_gen3_tx_pcs
	wire	[7:0]	w_hssi_gen3_tx_pcs_avmmreaddata;
	wire		w_hssi_gen3_tx_pcs_blockselect;
	wire	[31:0]	w_hssi_gen3_tx_pcs_data_out;
	wire	[35:0]	w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out;
	wire	[31:0]	w_hssi_gen3_tx_pcs_par_lpbk_out;
	wire	[19:0]	w_hssi_gen3_tx_pcs_tx_test_out;
	
	// wires for module twentynm_hssi_8g_rx_pcs
	wire	[3:0]	w_hssi_8g_rx_pcs_a1a2k1k2flag;
	wire	[7:0]	w_hssi_8g_rx_pcs_avmmreaddata;
	wire		w_hssi_8g_rx_pcs_blockselect;
	wire	[19:0]	w_hssi_8g_rx_pcs_chnl_test_bus_out;
	wire		w_hssi_8g_rx_pcs_clock_to_pld;
	wire	[63:0]	w_hssi_8g_rx_pcs_dataout;
	wire		w_hssi_8g_rx_pcs_dis_pc_byte;
	wire		w_hssi_8g_rx_pcs_eidle_detected;
	wire	[2:0]	w_hssi_8g_rx_pcs_eios_det_cdr_ctrl;
	wire		w_hssi_8g_rx_pcs_g3_rx_pma_rstn;
	wire		w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn;
	wire		w_hssi_8g_rx_pcs_gen2ngen1;
	wire	[19:0]	w_hssi_8g_rx_pcs_parallel_rev_loopback;
	wire		w_hssi_8g_rx_pcs_pc_fifo_empty;
	wire		w_hssi_8g_rx_pcs_pcfifofull;
	wire		w_hssi_8g_rx_pcs_phystatus;
	wire	[63:0]	w_hssi_8g_rx_pcs_pipe_data;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_up;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo;
	wire	[7:0]	w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rm_fifo_empty;
	wire		w_hssi_8g_rx_pcs_rm_fifo_full;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_blk_start;
	wire		w_hssi_8g_rx_pcs_rx_clk_out_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clkslip;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_data_valid;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rx_pipe_clk;
	wire		w_hssi_8g_rx_pcs_rx_pipe_soft_reset;
	wire		w_hssi_8g_rx_pcs_rx_pma_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_sync_hdr;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_up;
	wire	[2:0]	w_hssi_8g_rx_pcs_rxstatus;
	wire		w_hssi_8g_rx_pcs_rxvalid;
	wire		w_hssi_8g_rx_pcs_signal_detect_out;
	wire	[4:0]	w_hssi_8g_rx_pcs_word_align_boundary;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk;
	wire	[79:0]	w_hssi_8g_rx_pcs_wr_data_rx_phfifo;
	wire	[31:0]	w_hssi_8g_rx_pcs_wr_data_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo;
	
	// wires for module twentynm_hssi_fifo_rx_pcs
	wire	[7:0]	w_hssi_fifo_rx_pcs_avmmreaddata;
	wire		w_hssi_fifo_rx_pcs_blockselect;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out2_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out_8g_clock_comp;
	wire	[79:0]	w_hssi_fifo_rx_pcs_data_out_8g_phase_comp;
	wire	[39:0]	w_hssi_fifo_rx_pcs_data_out_gen3;
	
	// wires for module twentynm_hssi_common_pcs_pma_interface
	wire	[7:0]	w_hssi_common_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_common_pcs_pma_interface_blockselect;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in;
	wire	[19:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out;
	wire	[7:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus;
	wire		w_hssi_common_pcs_pma_interface_pma_adapt_start;
	wire		w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
	wire		w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
	wire	[17:0]	w_hssi_common_pcs_pma_interface_pma_current_coeff;
	wire	[2:0]	w_hssi_common_pcs_pma_interface_pma_current_rxpreset;
	wire		w_hssi_common_pcs_pma_interface_pma_early_eios;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_interface_select;
	wire		w_hssi_common_pcs_pma_interface_pma_ltd_b;
	wire		w_hssi_common_pcs_pma_interface_pma_ltr;
	wire		w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
	wire		w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_pcie_switch;
	wire		w_hssi_common_pcs_pma_interface_pma_ppm_lock;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_pma_reserved_out;
	wire		w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
	wire		w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up;
	
	
	generate
		
		//module instantiations
		
		// instantiating twentynm_hssi_10g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_rx_pcs
			twentynm_hssi_10g_rx_pcs #(
				.advanced_user_mode(hssi_10g_rx_pcs_advanced_user_mode),
				.align_del(hssi_10g_rx_pcs_align_del),
				.ber_bit_err_total_cnt(hssi_10g_rx_pcs_ber_bit_err_total_cnt),
				.ber_clken(hssi_10g_rx_pcs_ber_clken),
				.ber_xus_timer_window(hssi_10g_rx_pcs_ber_xus_timer_window),
				.bitslip_mode(hssi_10g_rx_pcs_bitslip_mode),
				.blksync_bitslip_type(hssi_10g_rx_pcs_blksync_bitslip_type),
				.blksync_bitslip_wait_cnt(hssi_10g_rx_pcs_blksync_bitslip_wait_cnt),
				.blksync_bitslip_wait_type(hssi_10g_rx_pcs_blksync_bitslip_wait_type),
				.blksync_bypass(hssi_10g_rx_pcs_blksync_bypass),
				.blksync_clken(hssi_10g_rx_pcs_blksync_clken),
				.blksync_enum_invalid_sh_cnt(hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt),
				.blksync_knum_sh_cnt_postlock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock),
				.blksync_knum_sh_cnt_prelock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock),
				.blksync_pipeln(hssi_10g_rx_pcs_blksync_pipeln),
				.clr_errblk_cnt_en(hssi_10g_rx_pcs_clr_errblk_cnt_en),
				.control_del(hssi_10g_rx_pcs_control_del),
				.crcchk_bypass(hssi_10g_rx_pcs_crcchk_bypass),
				.crcchk_clken(hssi_10g_rx_pcs_crcchk_clken),
				.crcchk_inv(hssi_10g_rx_pcs_crcchk_inv),
				.crcchk_pipeln(hssi_10g_rx_pcs_crcchk_pipeln),
				.crcflag_pipeln(hssi_10g_rx_pcs_crcflag_pipeln),
				.ctrl_bit_reverse(hssi_10g_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_10g_rx_pcs_data_bit_reverse),
				.dec64b66b_clken(hssi_10g_rx_pcs_dec64b66b_clken),
				.dec_64b66b_rxsm_bypass(hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass),
				.descrm_bypass(hssi_10g_rx_pcs_descrm_bypass),
				.descrm_clken(hssi_10g_rx_pcs_descrm_clken),
				.descrm_mode(hssi_10g_rx_pcs_descrm_mode),
				.descrm_pipeln(hssi_10g_rx_pcs_descrm_pipeln),
				.dft_clk_out_sel(hssi_10g_rx_pcs_dft_clk_out_sel),
				.dis_signal_ok(hssi_10g_rx_pcs_dis_signal_ok),
				.dispchk_bypass(hssi_10g_rx_pcs_dispchk_bypass),
				.empty_flag_type(hssi_10g_rx_pcs_empty_flag_type),
				.fast_path(hssi_10g_rx_pcs_fast_path),
				.fec_clken(hssi_10g_rx_pcs_fec_clken),
				.fec_enable(hssi_10g_rx_pcs_fec_enable),
				.fifo_double_read(hssi_10g_rx_pcs_fifo_double_read),
				.fifo_stop_rd(hssi_10g_rx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_rx_pcs_fifo_stop_wr),
				.force_align(hssi_10g_rx_pcs_force_align),
				.frmsync_bypass(hssi_10g_rx_pcs_frmsync_bypass),
				.frmsync_clken(hssi_10g_rx_pcs_frmsync_clken),
				.frmsync_enum_scrm(hssi_10g_rx_pcs_frmsync_enum_scrm),
				.frmsync_enum_sync(hssi_10g_rx_pcs_frmsync_enum_sync),
				.frmsync_flag_type(hssi_10g_rx_pcs_frmsync_flag_type),
				.frmsync_knum_sync(hssi_10g_rx_pcs_frmsync_knum_sync),
				.frmsync_mfrm_length(hssi_10g_rx_pcs_frmsync_mfrm_length),
				.frmsync_pipeln(hssi_10g_rx_pcs_frmsync_pipeln),
				.full_flag_type(hssi_10g_rx_pcs_full_flag_type),
				.gb_rx_idwidth(hssi_10g_rx_pcs_gb_rx_idwidth),
				.gb_rx_odwidth(hssi_10g_rx_pcs_gb_rx_odwidth),
				.gbexp_clken(hssi_10g_rx_pcs_gbexp_clken),
				.low_latency_en(hssi_10g_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_10g_rx_pcs_lpbk_mode),
				.master_clk_sel(hssi_10g_rx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_rx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_rx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_rx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_rx_pcs_pld_if_type),
				.prot_mode(hssi_10g_rx_pcs_prot_mode),
				.rand_clken(hssi_10g_rx_pcs_rand_clken),
				.rd_clk_sel(hssi_10g_rx_pcs_rd_clk_sel),
				.rdfifo_clken(hssi_10g_rx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_rx_pcs_reconfig_settings),
				.rx_fifo_write_ctrl(hssi_10g_rx_pcs_rx_fifo_write_ctrl),
				.rx_scrm_width(hssi_10g_rx_pcs_rx_scrm_width),
				.rx_sh_location(hssi_10g_rx_pcs_rx_sh_location),
				.rx_signal_ok_sel(hssi_10g_rx_pcs_rx_signal_ok_sel),
				.rx_sm_bypass(hssi_10g_rx_pcs_rx_sm_bypass),
				.rx_sm_hiber(hssi_10g_rx_pcs_rx_sm_hiber),
				.rx_sm_pipeln(hssi_10g_rx_pcs_rx_sm_pipeln),
				.rx_testbus_sel(hssi_10g_rx_pcs_rx_testbus_sel),
				.rx_true_b2b(hssi_10g_rx_pcs_rx_true_b2b),
				.rxfifo_empty(hssi_10g_rx_pcs_rxfifo_empty),
				.rxfifo_full(hssi_10g_rx_pcs_rxfifo_full),
				.rxfifo_mode(hssi_10g_rx_pcs_rxfifo_mode),
				.rxfifo_pempty(hssi_10g_rx_pcs_rxfifo_pempty),
				.rxfifo_pfull(hssi_10g_rx_pcs_rxfifo_pfull),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.stretch_num_stages(hssi_10g_rx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_rx_pcs_sup_mode),
				.test_mode(hssi_10g_rx_pcs_test_mode),
				.wrfifo_clken(hssi_10g_rx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_rx_pcs_blockselect),
				.rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.rx_control(w_hssi_10g_rx_pcs_rx_control),
				.rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.rx_data(w_hssi_10g_rx_pcs_rx_data),
				.rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.rx_diag_status(w_hssi_10g_rx_pcs_rx_diag_status),
				.rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.rx_fec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.rx_fifo_num(w_hssi_10g_rx_pcs_rx_fifo_num),
				.rx_fifo_rd_ptr(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr),
				.rx_fifo_rd_ptr2(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2),
				.rx_fifo_wr_clk(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.rx_fifo_wr_data(w_hssi_10g_rx_pcs_rx_fifo_wr_data),
				.rx_fifo_wr_en(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.rx_fifo_wr_ptr(w_hssi_10g_rx_pcs_rx_fifo_wr_ptr),
				.rx_fifo_wr_rst_n(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.rx_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_rx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_rx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.rx_control_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0]}),
				.rx_control_in_krfec({w_hssi_krfec_rx_pcs_rx_control_out[9], w_hssi_krfec_rx_pcs_rx_control_out[8], w_hssi_krfec_rx_pcs_rx_control_out[7], w_hssi_krfec_rx_pcs_rx_control_out[6], w_hssi_krfec_rx_pcs_rx_control_out[5], w_hssi_krfec_rx_pcs_rx_control_out[4], w_hssi_krfec_rx_pcs_rx_control_out[3], w_hssi_krfec_rx_pcs_rx_control_out[2], w_hssi_krfec_rx_pcs_rx_control_out[1], w_hssi_krfec_rx_pcs_rx_control_out[0]}),
				.rx_data_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0]}),
				.rx_data_in_krfec({w_hssi_krfec_rx_pcs_rx_data_out[63], w_hssi_krfec_rx_pcs_rx_data_out[62], w_hssi_krfec_rx_pcs_rx_data_out[61], w_hssi_krfec_rx_pcs_rx_data_out[60], w_hssi_krfec_rx_pcs_rx_data_out[59], w_hssi_krfec_rx_pcs_rx_data_out[58], w_hssi_krfec_rx_pcs_rx_data_out[57], w_hssi_krfec_rx_pcs_rx_data_out[56], w_hssi_krfec_rx_pcs_rx_data_out[55], w_hssi_krfec_rx_pcs_rx_data_out[54], w_hssi_krfec_rx_pcs_rx_data_out[53], w_hssi_krfec_rx_pcs_rx_data_out[52], w_hssi_krfec_rx_pcs_rx_data_out[51], w_hssi_krfec_rx_pcs_rx_data_out[50], w_hssi_krfec_rx_pcs_rx_data_out[49], w_hssi_krfec_rx_pcs_rx_data_out[48], w_hssi_krfec_rx_pcs_rx_data_out[47], w_hssi_krfec_rx_pcs_rx_data_out[46], w_hssi_krfec_rx_pcs_rx_data_out[45], w_hssi_krfec_rx_pcs_rx_data_out[44], w_hssi_krfec_rx_pcs_rx_data_out[43], w_hssi_krfec_rx_pcs_rx_data_out[42], w_hssi_krfec_rx_pcs_rx_data_out[41], w_hssi_krfec_rx_pcs_rx_data_out[40], w_hssi_krfec_rx_pcs_rx_data_out[39], w_hssi_krfec_rx_pcs_rx_data_out[38], w_hssi_krfec_rx_pcs_rx_data_out[37], w_hssi_krfec_rx_pcs_rx_data_out[36], w_hssi_krfec_rx_pcs_rx_data_out[35], w_hssi_krfec_rx_pcs_rx_data_out[34], w_hssi_krfec_rx_pcs_rx_data_out[33], w_hssi_krfec_rx_pcs_rx_data_out[32], w_hssi_krfec_rx_pcs_rx_data_out[31], w_hssi_krfec_rx_pcs_rx_data_out[30], w_hssi_krfec_rx_pcs_rx_data_out[29], w_hssi_krfec_rx_pcs_rx_data_out[28], w_hssi_krfec_rx_pcs_rx_data_out[27], w_hssi_krfec_rx_pcs_rx_data_out[26], w_hssi_krfec_rx_pcs_rx_data_out[25], w_hssi_krfec_rx_pcs_rx_data_out[24], w_hssi_krfec_rx_pcs_rx_data_out[23], w_hssi_krfec_rx_pcs_rx_data_out[22], w_hssi_krfec_rx_pcs_rx_data_out[21], w_hssi_krfec_rx_pcs_rx_data_out[20], w_hssi_krfec_rx_pcs_rx_data_out[19], w_hssi_krfec_rx_pcs_rx_data_out[18], w_hssi_krfec_rx_pcs_rx_data_out[17], w_hssi_krfec_rx_pcs_rx_data_out[16], w_hssi_krfec_rx_pcs_rx_data_out[15], w_hssi_krfec_rx_pcs_rx_data_out[14], w_hssi_krfec_rx_pcs_rx_data_out[13], w_hssi_krfec_rx_pcs_rx_data_out[12], w_hssi_krfec_rx_pcs_rx_data_out[11], w_hssi_krfec_rx_pcs_rx_data_out[10], w_hssi_krfec_rx_pcs_rx_data_out[9], w_hssi_krfec_rx_pcs_rx_data_out[8], w_hssi_krfec_rx_pcs_rx_data_out[7], w_hssi_krfec_rx_pcs_rx_data_out[6], w_hssi_krfec_rx_pcs_rx_data_out[5], w_hssi_krfec_rx_pcs_rx_data_out[4], w_hssi_krfec_rx_pcs_rx_data_out[3], w_hssi_krfec_rx_pcs_rx_data_out[2], w_hssi_krfec_rx_pcs_rx_data_out[1], w_hssi_krfec_rx_pcs_rx_data_out[0]}),
				.rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.rx_data_valid_in_krfec(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_10g[73], w_hssi_fifo_rx_pcs_data_out_10g[72], w_hssi_fifo_rx_pcs_data_out_10g[71], w_hssi_fifo_rx_pcs_data_out_10g[70], w_hssi_fifo_rx_pcs_data_out_10g[69], w_hssi_fifo_rx_pcs_data_out_10g[68], w_hssi_fifo_rx_pcs_data_out_10g[67], w_hssi_fifo_rx_pcs_data_out_10g[66], w_hssi_fifo_rx_pcs_data_out_10g[65], w_hssi_fifo_rx_pcs_data_out_10g[64], w_hssi_fifo_rx_pcs_data_out_10g[63], w_hssi_fifo_rx_pcs_data_out_10g[62], w_hssi_fifo_rx_pcs_data_out_10g[61], w_hssi_fifo_rx_pcs_data_out_10g[60], w_hssi_fifo_rx_pcs_data_out_10g[59], w_hssi_fifo_rx_pcs_data_out_10g[58], w_hssi_fifo_rx_pcs_data_out_10g[57], w_hssi_fifo_rx_pcs_data_out_10g[56], w_hssi_fifo_rx_pcs_data_out_10g[55], w_hssi_fifo_rx_pcs_data_out_10g[54], w_hssi_fifo_rx_pcs_data_out_10g[53], w_hssi_fifo_rx_pcs_data_out_10g[52], w_hssi_fifo_rx_pcs_data_out_10g[51], w_hssi_fifo_rx_pcs_data_out_10g[50], w_hssi_fifo_rx_pcs_data_out_10g[49], w_hssi_fifo_rx_pcs_data_out_10g[48], w_hssi_fifo_rx_pcs_data_out_10g[47], w_hssi_fifo_rx_pcs_data_out_10g[46], w_hssi_fifo_rx_pcs_data_out_10g[45], w_hssi_fifo_rx_pcs_data_out_10g[44], w_hssi_fifo_rx_pcs_data_out_10g[43], w_hssi_fifo_rx_pcs_data_out_10g[42], w_hssi_fifo_rx_pcs_data_out_10g[41], w_hssi_fifo_rx_pcs_data_out_10g[40], w_hssi_fifo_rx_pcs_data_out_10g[39], w_hssi_fifo_rx_pcs_data_out_10g[38], w_hssi_fifo_rx_pcs_data_out_10g[37], w_hssi_fifo_rx_pcs_data_out_10g[36], w_hssi_fifo_rx_pcs_data_out_10g[35], w_hssi_fifo_rx_pcs_data_out_10g[34], w_hssi_fifo_rx_pcs_data_out_10g[33], w_hssi_fifo_rx_pcs_data_out_10g[32], w_hssi_fifo_rx_pcs_data_out_10g[31], w_hssi_fifo_rx_pcs_data_out_10g[30], w_hssi_fifo_rx_pcs_data_out_10g[29], w_hssi_fifo_rx_pcs_data_out_10g[28], w_hssi_fifo_rx_pcs_data_out_10g[27], w_hssi_fifo_rx_pcs_data_out_10g[26], w_hssi_fifo_rx_pcs_data_out_10g[25], w_hssi_fifo_rx_pcs_data_out_10g[24], w_hssi_fifo_rx_pcs_data_out_10g[23], w_hssi_fifo_rx_pcs_data_out_10g[22], w_hssi_fifo_rx_pcs_data_out_10g[21], w_hssi_fifo_rx_pcs_data_out_10g[20], w_hssi_fifo_rx_pcs_data_out_10g[19], w_hssi_fifo_rx_pcs_data_out_10g[18], w_hssi_fifo_rx_pcs_data_out_10g[17], w_hssi_fifo_rx_pcs_data_out_10g[16], w_hssi_fifo_rx_pcs_data_out_10g[15], w_hssi_fifo_rx_pcs_data_out_10g[14], w_hssi_fifo_rx_pcs_data_out_10g[13], w_hssi_fifo_rx_pcs_data_out_10g[12], w_hssi_fifo_rx_pcs_data_out_10g[11], w_hssi_fifo_rx_pcs_data_out_10g[10], w_hssi_fifo_rx_pcs_data_out_10g[9], w_hssi_fifo_rx_pcs_data_out_10g[8], w_hssi_fifo_rx_pcs_data_out_10g[7], w_hssi_fifo_rx_pcs_data_out_10g[6], w_hssi_fifo_rx_pcs_data_out_10g[5], w_hssi_fifo_rx_pcs_data_out_10g[4], w_hssi_fifo_rx_pcs_data_out_10g[3], w_hssi_fifo_rx_pcs_data_out_10g[2], w_hssi_fifo_rx_pcs_data_out_10g[1], w_hssi_fifo_rx_pcs_data_out_10g[0]}),
				.rx_fifo_rd_data_dw({w_hssi_fifo_rx_pcs_data_out2_10g[73], w_hssi_fifo_rx_pcs_data_out2_10g[72], w_hssi_fifo_rx_pcs_data_out2_10g[71], w_hssi_fifo_rx_pcs_data_out2_10g[70], w_hssi_fifo_rx_pcs_data_out2_10g[69], w_hssi_fifo_rx_pcs_data_out2_10g[68], w_hssi_fifo_rx_pcs_data_out2_10g[67], w_hssi_fifo_rx_pcs_data_out2_10g[66], w_hssi_fifo_rx_pcs_data_out2_10g[65], w_hssi_fifo_rx_pcs_data_out2_10g[64], w_hssi_fifo_rx_pcs_data_out2_10g[63], w_hssi_fifo_rx_pcs_data_out2_10g[62], w_hssi_fifo_rx_pcs_data_out2_10g[61], w_hssi_fifo_rx_pcs_data_out2_10g[60], w_hssi_fifo_rx_pcs_data_out2_10g[59], w_hssi_fifo_rx_pcs_data_out2_10g[58], w_hssi_fifo_rx_pcs_data_out2_10g[57], w_hssi_fifo_rx_pcs_data_out2_10g[56], w_hssi_fifo_rx_pcs_data_out2_10g[55], w_hssi_fifo_rx_pcs_data_out2_10g[54], w_hssi_fifo_rx_pcs_data_out2_10g[53], w_hssi_fifo_rx_pcs_data_out2_10g[52], w_hssi_fifo_rx_pcs_data_out2_10g[51], w_hssi_fifo_rx_pcs_data_out2_10g[50], w_hssi_fifo_rx_pcs_data_out2_10g[49], w_hssi_fifo_rx_pcs_data_out2_10g[48], w_hssi_fifo_rx_pcs_data_out2_10g[47], w_hssi_fifo_rx_pcs_data_out2_10g[46], w_hssi_fifo_rx_pcs_data_out2_10g[45], w_hssi_fifo_rx_pcs_data_out2_10g[44], w_hssi_fifo_rx_pcs_data_out2_10g[43], w_hssi_fifo_rx_pcs_data_out2_10g[42], w_hssi_fifo_rx_pcs_data_out2_10g[41], w_hssi_fifo_rx_pcs_data_out2_10g[40], w_hssi_fifo_rx_pcs_data_out2_10g[39], w_hssi_fifo_rx_pcs_data_out2_10g[38], w_hssi_fifo_rx_pcs_data_out2_10g[37], w_hssi_fifo_rx_pcs_data_out2_10g[36], w_hssi_fifo_rx_pcs_data_out2_10g[35], w_hssi_fifo_rx_pcs_data_out2_10g[34], w_hssi_fifo_rx_pcs_data_out2_10g[33], w_hssi_fifo_rx_pcs_data_out2_10g[32], w_hssi_fifo_rx_pcs_data_out2_10g[31], w_hssi_fifo_rx_pcs_data_out2_10g[30], w_hssi_fifo_rx_pcs_data_out2_10g[29], w_hssi_fifo_rx_pcs_data_out2_10g[28], w_hssi_fifo_rx_pcs_data_out2_10g[27], w_hssi_fifo_rx_pcs_data_out2_10g[26], w_hssi_fifo_rx_pcs_data_out2_10g[25], w_hssi_fifo_rx_pcs_data_out2_10g[24], w_hssi_fifo_rx_pcs_data_out2_10g[23], w_hssi_fifo_rx_pcs_data_out2_10g[22], w_hssi_fifo_rx_pcs_data_out2_10g[21], w_hssi_fifo_rx_pcs_data_out2_10g[20], w_hssi_fifo_rx_pcs_data_out2_10g[19], w_hssi_fifo_rx_pcs_data_out2_10g[18], w_hssi_fifo_rx_pcs_data_out2_10g[17], w_hssi_fifo_rx_pcs_data_out2_10g[16], w_hssi_fifo_rx_pcs_data_out2_10g[15], w_hssi_fifo_rx_pcs_data_out2_10g[14], w_hssi_fifo_rx_pcs_data_out2_10g[13], w_hssi_fifo_rx_pcs_data_out2_10g[12], w_hssi_fifo_rx_pcs_data_out2_10g[11], w_hssi_fifo_rx_pcs_data_out2_10g[10], w_hssi_fifo_rx_pcs_data_out2_10g[9], w_hssi_fifo_rx_pcs_data_out2_10g[8], w_hssi_fifo_rx_pcs_data_out2_10g[7], w_hssi_fifo_rx_pcs_data_out2_10g[6], w_hssi_fifo_rx_pcs_data_out2_10g[5], w_hssi_fifo_rx_pcs_data_out2_10g[4], w_hssi_fifo_rx_pcs_data_out2_10g[3], w_hssi_fifo_rx_pcs_data_out2_10g[2], w_hssi_fifo_rx_pcs_data_out2_10g[1], w_hssi_fifo_rx_pcs_data_out2_10g[0]}),
				.rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.rx_pma_data({w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0]}),
				.rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.signal_ok_krfec(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_10g_reg(),
				.pld_10g_krfec_rx_blk_lock_10g_txclk_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_txclk_reg(),
				.pld_10g_krfec_rx_frame_10g_reg(),
				.pld_10g_krfec_rx_frame_10g_txclk_reg(),
				.pld_10g_krfec_rx_pld_rst_n_fifo(),
				.pld_10g_krfec_rx_pld_rst_n_reg(),
				.pld_10g_krfec_rx_pld_rst_n_txclk_reg(),
				.pld_10g_rx_align_clr_fifo(),
				.pld_10g_rx_align_clr_reg(),
				.pld_10g_rx_align_clr_txclk_reg(),
				.pld_10g_rx_align_val_fifo(),
				.pld_10g_rx_align_val_reg(),
				.pld_10g_rx_align_val_txclk_reg(),
				.pld_10g_rx_clr_ber_count_reg(),
				.pld_10g_rx_clr_ber_count_txclk_reg(),
				.pld_10g_rx_crc32_err_reg(),
				.pld_10g_rx_crc32_err_txclk_reg(),
				.pld_10g_rx_data_valid_10g_reg(),
				.pld_10g_rx_data_valid_fifo(),
				.pld_10g_rx_data_valid_pcsdirect_reg(),
				.pld_10g_rx_data_valid_txclk_reg(),
				.pld_10g_rx_empty_fifo(),
				.pld_10g_rx_fifo_del_reg(),
				.pld_10g_rx_fifo_del_txclk_reg(),
				.pld_10g_rx_fifo_insert_fifo(),
				.pld_10g_rx_fifo_num_reg(),
				.pld_10g_rx_fifo_num_txclk_reg(),
				.pld_10g_rx_frame_lock_reg(),
				.pld_10g_rx_frame_lock_txclk_reg(),
				.pld_10g_rx_hi_ber_reg(),
				.pld_10g_rx_hi_ber_txclk_reg(),
				.pld_10g_rx_oflw_err_reg(),
				.pld_10g_rx_oflw_err_txclk_reg(),
				.pld_10g_rx_pempty_fifo(),
				.pld_10g_rx_pfull_reg(),
				.pld_10g_rx_pfull_txclk_reg(),
				.pld_10g_rx_rd_en_fifo(),
				.pld_pcs_rx_clk_out_10g_txclk_wire(),
				.pld_pcs_rx_clk_out_10g_wire(),
				.pld_rx_control_10g_reg(),
				.pld_rx_control_10g_txclk_reg(),
				.pld_rx_data_10g_reg(),
				.pld_rx_data_10g_txclk_reg(),
				.pld_rx_prbs_err_10g_txclk_reg(),
				.pld_rx_prbs_err_clr_10g_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_10g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_align_val = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_blk_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_control[19:0] = 20'b0;
				assign w_hssi_10g_rx_pcs_rx_crc32_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_data[127:0] = 128'b0;
				assign w_hssi_10g_rx_pcs_rx_data_valid = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_dft_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_diag_status[1:0] = 2'b0;
				assign w_hssi_10g_rx_pcs_rx_empty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fec_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_del = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_insert = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_data[73:0] = 74'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_frame_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_hi_ber = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_oflw_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pempty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pfull = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_random_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_rx_frame = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_10g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_tx_pcs
			twentynm_hssi_10g_tx_pcs #(
				.advanced_user_mode(hssi_10g_tx_pcs_advanced_user_mode),
				.bitslip_en(hssi_10g_tx_pcs_bitslip_en),
				.bonding_dft_en(hssi_10g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_10g_tx_pcs_bonding_dft_val),
				.comp_cnt(hssi_10g_tx_pcs_comp_cnt),
				.compin_sel(hssi_10g_tx_pcs_compin_sel),
				.crcgen_bypass(hssi_10g_tx_pcs_crcgen_bypass),
				.crcgen_clken(hssi_10g_tx_pcs_crcgen_clken),
				.crcgen_err(hssi_10g_tx_pcs_crcgen_err),
				.crcgen_inv(hssi_10g_tx_pcs_crcgen_inv),
				.ctrl_bit_reverse(hssi_10g_tx_pcs_ctrl_bit_reverse),
				.ctrl_plane_bonding(hssi_10g_tx_pcs_ctrl_plane_bonding),
				.data_bit_reverse(hssi_10g_tx_pcs_data_bit_reverse),
				.dft_clk_out_sel(hssi_10g_tx_pcs_dft_clk_out_sel),
				.dispgen_bypass(hssi_10g_tx_pcs_dispgen_bypass),
				.dispgen_clken(hssi_10g_tx_pcs_dispgen_clken),
				.dispgen_err(hssi_10g_tx_pcs_dispgen_err),
				.dispgen_pipeln(hssi_10g_tx_pcs_dispgen_pipeln),
				.distdwn_bypass_pipeln(hssi_10g_tx_pcs_distdwn_bypass_pipeln),
				.distdwn_master(hssi_10g_tx_pcs_distdwn_master),
				.distup_bypass_pipeln(hssi_10g_tx_pcs_distup_bypass_pipeln),
				.distup_master(hssi_10g_tx_pcs_distup_master),
				.dv_bond(hssi_10g_tx_pcs_dv_bond),
				.empty_flag_type(hssi_10g_tx_pcs_empty_flag_type),
				.enc64b66b_txsm_clken(hssi_10g_tx_pcs_enc64b66b_txsm_clken),
				.enc_64b66b_txsm_bypass(hssi_10g_tx_pcs_enc_64b66b_txsm_bypass),
				.fastpath(hssi_10g_tx_pcs_fastpath),
				.fec_clken(hssi_10g_tx_pcs_fec_clken),
				.fec_enable(hssi_10g_tx_pcs_fec_enable),
				.fifo_double_write(hssi_10g_tx_pcs_fifo_double_write),
				.fifo_reg_fast(hssi_10g_tx_pcs_fifo_reg_fast),
				.fifo_stop_rd(hssi_10g_tx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_tx_pcs_fifo_stop_wr),
				.frmgen_burst(hssi_10g_tx_pcs_frmgen_burst),
				.frmgen_bypass(hssi_10g_tx_pcs_frmgen_bypass),
				.frmgen_clken(hssi_10g_tx_pcs_frmgen_clken),
				.frmgen_mfrm_length(hssi_10g_tx_pcs_frmgen_mfrm_length),
				.frmgen_pipeln(hssi_10g_tx_pcs_frmgen_pipeln),
				.frmgen_pyld_ins(hssi_10g_tx_pcs_frmgen_pyld_ins),
				.frmgen_wordslip(hssi_10g_tx_pcs_frmgen_wordslip),
				.full_flag_type(hssi_10g_tx_pcs_full_flag_type),
				.gb_pipeln_bypass(hssi_10g_tx_pcs_gb_pipeln_bypass),
				.gb_tx_idwidth(hssi_10g_tx_pcs_gb_tx_idwidth),
				.gb_tx_odwidth(hssi_10g_tx_pcs_gb_tx_odwidth),
				.gbred_clken(hssi_10g_tx_pcs_gbred_clken),
				.indv(hssi_10g_tx_pcs_indv),
				.low_latency_en(hssi_10g_tx_pcs_low_latency_en),
				.master_clk_sel(hssi_10g_tx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_tx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_tx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_tx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_tx_pcs_pld_if_type),
				.prot_mode(hssi_10g_tx_pcs_prot_mode),
				.pseudo_random(hssi_10g_tx_pcs_pseudo_random),
				.pseudo_seed_a(hssi_10g_tx_pcs_pseudo_seed_a),
				.pseudo_seed_b(hssi_10g_tx_pcs_pseudo_seed_b),
				.random_disp(hssi_10g_tx_pcs_random_disp),
				.rdfifo_clken(hssi_10g_tx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_tx_pcs_reconfig_settings),
				.scrm_bypass(hssi_10g_tx_pcs_scrm_bypass),
				.scrm_clken(hssi_10g_tx_pcs_scrm_clken),
				.scrm_mode(hssi_10g_tx_pcs_scrm_mode),
				.scrm_pipeln(hssi_10g_tx_pcs_scrm_pipeln),
				.sh_err(hssi_10g_tx_pcs_sh_err),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sop_mark(hssi_10g_tx_pcs_sop_mark),
				.stretch_num_stages(hssi_10g_tx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_tx_pcs_sup_mode),
				.test_mode(hssi_10g_tx_pcs_test_mode),
				.tx_scrm_err(hssi_10g_tx_pcs_tx_scrm_err),
				.tx_scrm_width(hssi_10g_tx_pcs_tx_scrm_width),
				.tx_sh_location(hssi_10g_tx_pcs_tx_sh_location),
				.tx_sm_bypass(hssi_10g_tx_pcs_tx_sm_bypass),
				.tx_sm_pipeln(hssi_10g_tx_pcs_tx_sm_pipeln),
				.tx_testbus_sel(hssi_10g_tx_pcs_tx_testbus_sel),
				.txfifo_empty(hssi_10g_tx_pcs_txfifo_empty),
				.txfifo_full(hssi_10g_tx_pcs_txfifo_full),
				.txfifo_mode(hssi_10g_tx_pcs_txfifo_mode),
				.txfifo_pempty(hssi_10g_tx_pcs_txfifo_pempty),
				.txfifo_pfull(hssi_10g_tx_pcs_txfifo_pfull),
				.wr_clk_sel(hssi_10g_tx_pcs_wr_clk_sel),
				.wrfifo_clken(hssi_10g_tx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_tx_pcs_blockselect),
				.distdwn_out_dv(w_hssi_10g_tx_pcs_distdwn_out_dv),
				.distdwn_out_rden(w_hssi_10g_tx_pcs_distdwn_out_rden),
				.distdwn_out_wren(w_hssi_10g_tx_pcs_distdwn_out_wren),
				.distup_out_dv(w_hssi_10g_tx_pcs_distup_out_dv),
				.distup_out_rden(w_hssi_10g_tx_pcs_distup_out_rden),
				.distup_out_wren(w_hssi_10g_tx_pcs_distup_out_wren),
				.tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pma_if(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.tx_control_out_krfec(w_hssi_10g_tx_pcs_tx_control_out_krfec),
				.tx_data_out_krfec(w_hssi_10g_tx_pcs_tx_data_out_krfec),
				.tx_data_valid_out_krfec(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.tx_fec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_fifo_num(w_hssi_10g_tx_pcs_tx_fifo_num),
				.tx_fifo_rd_ptr(w_hssi_10g_tx_pcs_tx_fifo_rd_ptr),
				.tx_fifo_wr_clk(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.tx_fifo_wr_data(w_hssi_10g_tx_pcs_tx_fifo_wr_data),
				.tx_fifo_wr_data_dw(w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw),
				.tx_fifo_wr_en(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.tx_fifo_wr_ptr(w_hssi_10g_tx_pcs_tx_fifo_wr_ptr),
				.tx_fifo_wr_rst_n(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.tx_full(w_hssi_10g_tx_pcs_tx_full),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				.tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.tx_pma_data(w_hssi_10g_tx_pcs_tx_pma_data),
				.tx_pma_gating_val(w_hssi_10g_tx_pcs_tx_pma_gating_val),
				.tx_test_data(w_hssi_10g_tx_pcs_tx_test_data),
				.tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.distdwn_in_dv(in_bond_pcs10g_in_bot[2]),
				.distdwn_in_rden(in_bond_pcs10g_in_bot[4]),
				.distdwn_in_wren(in_bond_pcs10g_in_bot[3]),
				.distup_in_dv(in_bond_pcs10g_in_top[2]),
				.distup_in_rden(in_bond_pcs10g_in_top[4]),
				.distup_in_wren(in_bond_pcs10g_in_top[3]),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_tx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_tx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.tx_bitslip({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0]}),
				.tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.tx_control({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0]}),
				.tx_control_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0]}),
				.tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0]}),
				.tx_data_in_krfec({w_hssi_krfec_tx_pcs_tx_data_out[63], w_hssi_krfec_tx_pcs_tx_data_out[62], w_hssi_krfec_tx_pcs_tx_data_out[61], w_hssi_krfec_tx_pcs_tx_data_out[60], w_hssi_krfec_tx_pcs_tx_data_out[59], w_hssi_krfec_tx_pcs_tx_data_out[58], w_hssi_krfec_tx_pcs_tx_data_out[57], w_hssi_krfec_tx_pcs_tx_data_out[56], w_hssi_krfec_tx_pcs_tx_data_out[55], w_hssi_krfec_tx_pcs_tx_data_out[54], w_hssi_krfec_tx_pcs_tx_data_out[53], w_hssi_krfec_tx_pcs_tx_data_out[52], w_hssi_krfec_tx_pcs_tx_data_out[51], w_hssi_krfec_tx_pcs_tx_data_out[50], w_hssi_krfec_tx_pcs_tx_data_out[49], w_hssi_krfec_tx_pcs_tx_data_out[48], w_hssi_krfec_tx_pcs_tx_data_out[47], w_hssi_krfec_tx_pcs_tx_data_out[46], w_hssi_krfec_tx_pcs_tx_data_out[45], w_hssi_krfec_tx_pcs_tx_data_out[44], w_hssi_krfec_tx_pcs_tx_data_out[43], w_hssi_krfec_tx_pcs_tx_data_out[42], w_hssi_krfec_tx_pcs_tx_data_out[41], w_hssi_krfec_tx_pcs_tx_data_out[40], w_hssi_krfec_tx_pcs_tx_data_out[39], w_hssi_krfec_tx_pcs_tx_data_out[38], w_hssi_krfec_tx_pcs_tx_data_out[37], w_hssi_krfec_tx_pcs_tx_data_out[36], w_hssi_krfec_tx_pcs_tx_data_out[35], w_hssi_krfec_tx_pcs_tx_data_out[34], w_hssi_krfec_tx_pcs_tx_data_out[33], w_hssi_krfec_tx_pcs_tx_data_out[32], w_hssi_krfec_tx_pcs_tx_data_out[31], w_hssi_krfec_tx_pcs_tx_data_out[30], w_hssi_krfec_tx_pcs_tx_data_out[29], w_hssi_krfec_tx_pcs_tx_data_out[28], w_hssi_krfec_tx_pcs_tx_data_out[27], w_hssi_krfec_tx_pcs_tx_data_out[26], w_hssi_krfec_tx_pcs_tx_data_out[25], w_hssi_krfec_tx_pcs_tx_data_out[24], w_hssi_krfec_tx_pcs_tx_data_out[23], w_hssi_krfec_tx_pcs_tx_data_out[22], w_hssi_krfec_tx_pcs_tx_data_out[21], w_hssi_krfec_tx_pcs_tx_data_out[20], w_hssi_krfec_tx_pcs_tx_data_out[19], w_hssi_krfec_tx_pcs_tx_data_out[18], w_hssi_krfec_tx_pcs_tx_data_out[17], w_hssi_krfec_tx_pcs_tx_data_out[16], w_hssi_krfec_tx_pcs_tx_data_out[15], w_hssi_krfec_tx_pcs_tx_data_out[14], w_hssi_krfec_tx_pcs_tx_data_out[13], w_hssi_krfec_tx_pcs_tx_data_out[12], w_hssi_krfec_tx_pcs_tx_data_out[11], w_hssi_krfec_tx_pcs_tx_data_out[10], w_hssi_krfec_tx_pcs_tx_data_out[9], w_hssi_krfec_tx_pcs_tx_data_out[8], w_hssi_krfec_tx_pcs_tx_data_out[7], w_hssi_krfec_tx_pcs_tx_data_out[6], w_hssi_krfec_tx_pcs_tx_data_out[5], w_hssi_krfec_tx_pcs_tx_data_out[4], w_hssi_krfec_tx_pcs_tx_data_out[3], w_hssi_krfec_tx_pcs_tx_data_out[2], w_hssi_krfec_tx_pcs_tx_data_out[1], w_hssi_krfec_tx_pcs_tx_data_out[0]}),
				.tx_data_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0]}),
				.tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.tx_diag_status({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0]}),
				.tx_fifo_rd_data({w_hssi_fifo_tx_pcs_data_out_10g[72], w_hssi_fifo_tx_pcs_data_out_10g[71], w_hssi_fifo_tx_pcs_data_out_10g[70], w_hssi_fifo_tx_pcs_data_out_10g[69], w_hssi_fifo_tx_pcs_data_out_10g[68], w_hssi_fifo_tx_pcs_data_out_10g[67], w_hssi_fifo_tx_pcs_data_out_10g[66], w_hssi_fifo_tx_pcs_data_out_10g[65], w_hssi_fifo_tx_pcs_data_out_10g[64], w_hssi_fifo_tx_pcs_data_out_10g[63], w_hssi_fifo_tx_pcs_data_out_10g[62], w_hssi_fifo_tx_pcs_data_out_10g[61], w_hssi_fifo_tx_pcs_data_out_10g[60], w_hssi_fifo_tx_pcs_data_out_10g[59], w_hssi_fifo_tx_pcs_data_out_10g[58], w_hssi_fifo_tx_pcs_data_out_10g[57], w_hssi_fifo_tx_pcs_data_out_10g[56], w_hssi_fifo_tx_pcs_data_out_10g[55], w_hssi_fifo_tx_pcs_data_out_10g[54], w_hssi_fifo_tx_pcs_data_out_10g[53], w_hssi_fifo_tx_pcs_data_out_10g[52], w_hssi_fifo_tx_pcs_data_out_10g[51], w_hssi_fifo_tx_pcs_data_out_10g[50], w_hssi_fifo_tx_pcs_data_out_10g[49], w_hssi_fifo_tx_pcs_data_out_10g[48], w_hssi_fifo_tx_pcs_data_out_10g[47], w_hssi_fifo_tx_pcs_data_out_10g[46], w_hssi_fifo_tx_pcs_data_out_10g[45], w_hssi_fifo_tx_pcs_data_out_10g[44], w_hssi_fifo_tx_pcs_data_out_10g[43], w_hssi_fifo_tx_pcs_data_out_10g[42], w_hssi_fifo_tx_pcs_data_out_10g[41], w_hssi_fifo_tx_pcs_data_out_10g[40], w_hssi_fifo_tx_pcs_data_out_10g[39], w_hssi_fifo_tx_pcs_data_out_10g[38], w_hssi_fifo_tx_pcs_data_out_10g[37], w_hssi_fifo_tx_pcs_data_out_10g[36], w_hssi_fifo_tx_pcs_data_out_10g[35], w_hssi_fifo_tx_pcs_data_out_10g[34], w_hssi_fifo_tx_pcs_data_out_10g[33], w_hssi_fifo_tx_pcs_data_out_10g[32], w_hssi_fifo_tx_pcs_data_out_10g[31], w_hssi_fifo_tx_pcs_data_out_10g[30], w_hssi_fifo_tx_pcs_data_out_10g[29], w_hssi_fifo_tx_pcs_data_out_10g[28], w_hssi_fifo_tx_pcs_data_out_10g[27], w_hssi_fifo_tx_pcs_data_out_10g[26], w_hssi_fifo_tx_pcs_data_out_10g[25], w_hssi_fifo_tx_pcs_data_out_10g[24], w_hssi_fifo_tx_pcs_data_out_10g[23], w_hssi_fifo_tx_pcs_data_out_10g[22], w_hssi_fifo_tx_pcs_data_out_10g[21], w_hssi_fifo_tx_pcs_data_out_10g[20], w_hssi_fifo_tx_pcs_data_out_10g[19], w_hssi_fifo_tx_pcs_data_out_10g[18], w_hssi_fifo_tx_pcs_data_out_10g[17], w_hssi_fifo_tx_pcs_data_out_10g[16], w_hssi_fifo_tx_pcs_data_out_10g[15], w_hssi_fifo_tx_pcs_data_out_10g[14], w_hssi_fifo_tx_pcs_data_out_10g[13], w_hssi_fifo_tx_pcs_data_out_10g[12], w_hssi_fifo_tx_pcs_data_out_10g[11], w_hssi_fifo_tx_pcs_data_out_10g[10], w_hssi_fifo_tx_pcs_data_out_10g[9], w_hssi_fifo_tx_pcs_data_out_10g[8], w_hssi_fifo_tx_pcs_data_out_10g[7], w_hssi_fifo_tx_pcs_data_out_10g[6], w_hssi_fifo_tx_pcs_data_out_10g[5], w_hssi_fifo_tx_pcs_data_out_10g[4], w_hssi_fifo_tx_pcs_data_out_10g[3], w_hssi_fifo_tx_pcs_data_out_10g[2], w_hssi_fifo_tx_pcs_data_out_10g[1], w_hssi_fifo_tx_pcs_data_out_10g[0]}),
				.tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_10g_reg(),
				.pld_10g_krfec_tx_pld_rst_n_fifo(),
				.pld_10g_krfec_tx_pld_rst_n_reg(),
				.pld_10g_tx_bitslip_reg(),
				.pld_10g_tx_burst_en_exe_reg(),
				.pld_10g_tx_data_valid_10g_reg(),
				.pld_10g_tx_data_valid_fifo(),
				.pld_10g_tx_data_valid_reg(),
				.pld_10g_tx_diag_status_reg(),
				.pld_10g_tx_empty_reg(),
				.pld_10g_tx_fifo_num_reg(),
				.pld_10g_tx_full_fifo(),
				.pld_10g_tx_full_reg(),
				.pld_10g_tx_pempty_reg(),
				.pld_10g_tx_pfull_fifo(),
				.pld_10g_tx_wordslip_exe_reg(),
				.pld_10g_tx_wordslip_reg(),
				.pld_pcs_tx_clk_out_10g_wire(),
				.pld_tx_burst_en_reg(),
				.pld_tx_control_lo_10g_reg(),
				.pld_tx_data_10g_fifo(),
				.pld_tx_data_lo_10g_reg()
			);
		end // if generate
		else begin
				assign w_hssi_10g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_burst_en_exe = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pma_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_control_out_krfec[8:0] = 9'b0;
				assign w_hssi_10g_tx_pcs_tx_data_out_krfec[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_data_valid_out_krfec = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_dft_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_empty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fec_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_full = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_pempty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pfull = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_gating_val[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_test_data[19:0] = 20'b0;
				assign w_hssi_10g_tx_pcs_tx_wordslip_exe = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_rx_pcs
			twentynm_hssi_8g_rx_pcs #(
				.auto_error_replacement(hssi_8g_rx_pcs_auto_error_replacement),
				.auto_speed_nego(hssi_8g_rx_pcs_auto_speed_nego),
				.bit_reversal(hssi_8g_rx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_rx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_rx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_rx_pcs_bypass_pipeline_reg),
				.byte_deserializer(hssi_8g_rx_pcs_byte_deserializer),
				.cdr_ctrl_rxvalid_mask(hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask),
				.clkcmp_pattern_n(hssi_8g_rx_pcs_clkcmp_pattern_n),
				.clkcmp_pattern_p(hssi_8g_rx_pcs_clkcmp_pattern_p),
				.clock_gate_bds_dec_asn(hssi_8g_rx_pcs_clock_gate_bds_dec_asn),
				.clock_gate_cdr_eidle(hssi_8g_rx_pcs_clock_gate_cdr_eidle),
				.clock_gate_dw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk),
				.clock_gate_dw_rm_rd(hssi_8g_rx_pcs_clock_gate_dw_rm_rd),
				.clock_gate_dw_rm_wr(hssi_8g_rx_pcs_clock_gate_dw_rm_wr),
				.clock_gate_dw_wa(hssi_8g_rx_pcs_clock_gate_dw_wa),
				.clock_gate_pc_rdclk(hssi_8g_rx_pcs_clock_gate_pc_rdclk),
				.clock_gate_sw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk),
				.clock_gate_sw_rm_rd(hssi_8g_rx_pcs_clock_gate_sw_rm_rd),
				.clock_gate_sw_rm_wr(hssi_8g_rx_pcs_clock_gate_sw_rm_wr),
				.clock_gate_sw_wa(hssi_8g_rx_pcs_clock_gate_sw_wa),
				.clock_observation_in_pld_core(hssi_8g_rx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_rx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_rx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_rx_pcs_ctrl_plane_bonding_distribution),
				.eidle_entry_eios(hssi_8g_rx_pcs_eidle_entry_eios),
				.eidle_entry_iei(hssi_8g_rx_pcs_eidle_entry_iei),
				.eidle_entry_sd(hssi_8g_rx_pcs_eidle_entry_sd),
				.eightb_tenb_decoder(hssi_8g_rx_pcs_eightb_tenb_decoder),
				.err_flags_sel(hssi_8g_rx_pcs_err_flags_sel),
				.fixed_pat_det(hssi_8g_rx_pcs_fixed_pat_det),
				.fixed_pat_num(hssi_8g_rx_pcs_fixed_pat_num),
				.force_signal_detect(hssi_8g_rx_pcs_force_signal_detect),
				.gen3_clk_en(hssi_8g_rx_pcs_gen3_clk_en),
				.gen3_rx_clk_sel(hssi_8g_rx_pcs_gen3_rx_clk_sel),
				.gen3_tx_clk_sel(hssi_8g_rx_pcs_gen3_tx_clk_sel),
				.hip_mode(hssi_8g_rx_pcs_hip_mode),
				.ibm_invalid_code(hssi_8g_rx_pcs_ibm_invalid_code),
				.invalid_code_flag_only(hssi_8g_rx_pcs_invalid_code_flag_only),
				.pad_or_edb_error_replace(hssi_8g_rx_pcs_pad_or_edb_error_replace),
				.pcs_bypass(hssi_8g_rx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_rx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_rx_pcs_phase_compensation_fifo),
				.pipe_if_enable(hssi_8g_rx_pcs_pipe_if_enable),
				.pma_dw(hssi_8g_rx_pcs_pma_dw),
				.polinv_8b10b_dec(hssi_8g_rx_pcs_polinv_8b10b_dec),
				.prot_mode(hssi_8g_rx_pcs_prot_mode),
				.rate_match(hssi_8g_rx_pcs_rate_match),
				.rate_match_del_thres(hssi_8g_rx_pcs_rate_match_del_thres),
				.rate_match_empty_thres(hssi_8g_rx_pcs_rate_match_empty_thres),
				.rate_match_full_thres(hssi_8g_rx_pcs_rate_match_full_thres),
				.rate_match_ins_thres(hssi_8g_rx_pcs_rate_match_ins_thres),
				.rate_match_start_thres(hssi_8g_rx_pcs_rate_match_start_thres),
				.reconfig_settings(hssi_8g_rx_pcs_reconfig_settings),
				.rx_clk2(hssi_8g_rx_pcs_rx_clk2),
				.rx_clk_free_running(hssi_8g_rx_pcs_rx_clk_free_running),
				.rx_pcs_urst(hssi_8g_rx_pcs_rx_pcs_urst),
				.rx_rcvd_clk(hssi_8g_rx_pcs_rx_rcvd_clk),
				.rx_rd_clk(hssi_8g_rx_pcs_rx_rd_clk),
				.rx_refclk(hssi_8g_rx_pcs_rx_refclk),
				.rx_wr_clk(hssi_8g_rx_pcs_rx_wr_clk),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_rx_pcs_sup_mode),
				.symbol_swap(hssi_8g_rx_pcs_symbol_swap),
				.sync_sm_idle_eios(hssi_8g_rx_pcs_sync_sm_idle_eios),
				.test_bus_sel(hssi_8g_rx_pcs_test_bus_sel),
				.tx_rx_parallel_loopback(hssi_8g_rx_pcs_tx_rx_parallel_loopback),
				.wa_boundary_lock_ctrl(hssi_8g_rx_pcs_wa_boundary_lock_ctrl),
				.wa_clk_slip_spacing(hssi_8g_rx_pcs_wa_clk_slip_spacing),
				.wa_det_latency_sync_status_beh(hssi_8g_rx_pcs_wa_det_latency_sync_status_beh),
				.wa_disp_err_flag(hssi_8g_rx_pcs_wa_disp_err_flag),
				.wa_kchar(hssi_8g_rx_pcs_wa_kchar),
				.wa_pd(hssi_8g_rx_pcs_wa_pd),
				.wa_pd_data(hssi_8g_rx_pcs_wa_pd_data),
				.wa_pd_polarity(hssi_8g_rx_pcs_wa_pd_polarity),
				.wa_pld_controlled(hssi_8g_rx_pcs_wa_pld_controlled),
				.wa_renumber_data(hssi_8g_rx_pcs_wa_renumber_data),
				.wa_rgnumber_data(hssi_8g_rx_pcs_wa_rgnumber_data),
				.wa_rknumber_data(hssi_8g_rx_pcs_wa_rknumber_data),
				.wa_rosnumber_data(hssi_8g_rx_pcs_wa_rosnumber_data),
				.wa_rvnumber_data(hssi_8g_rx_pcs_wa_rvnumber_data),
				.wa_sync_sm_ctrl(hssi_8g_rx_pcs_wa_sync_sm_ctrl),
				.wait_cnt(hssi_8g_rx_pcs_wait_cnt)
			) inst_twentynm_hssi_8g_rx_pcs (
				// OUTPUTS
				.a1a2k1k2flag(w_hssi_8g_rx_pcs_a1a2k1k2flag),
				.avmmreaddata(w_hssi_8g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_rx_pcs_blockselect),
				.chnl_test_bus_out(w_hssi_8g_rx_pcs_chnl_test_bus_out),
				.clock_to_pld(w_hssi_8g_rx_pcs_clock_to_pld),
				.dataout(w_hssi_8g_rx_pcs_dataout),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidle_detected(w_hssi_8g_rx_pcs_eidle_detected),
				.eios_det_cdr_ctrl(w_hssi_8g_rx_pcs_eios_det_cdr_ctrl),
				.g3_rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.g3_rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.gen2ngen1(w_hssi_8g_rx_pcs_gen2ngen1),
				.parallel_rev_loopback(w_hssi_8g_rx_pcs_parallel_rev_loopback),
				.pc_fifo_empty(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.pcfifofull(w_hssi_8g_rx_pcs_pcfifofull),
				.phystatus(w_hssi_8g_rx_pcs_phystatus),
				.pipe_data(w_hssi_8g_rx_pcs_pipe_data),
				.rd_enable_out_chnl_down(w_hssi_8g_rx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_rx_pcs_rd_enable_out_chnl_up),
				.rd_ptr1_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo),
				.rd_ptr2_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo),
				.rd_ptr_rx_phfifo(w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.reset_pc_ptrs_out_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down),
				.reset_pc_ptrs_out_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up),
				.rm_fifo_empty(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.rm_fifo_full(w_hssi_8g_rx_pcs_rm_fifo_full),
				.rx_blk_start(w_hssi_8g_rx_pcs_rx_blk_start),
				.rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.rx_data_valid(w_hssi_8g_rx_pcs_rx_data_valid),
				.rx_div_sync_out_chnl_down(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down),
				.rx_div_sync_out_chnl_up(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up),
				.rx_pipe_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.rx_pipe_soft_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rx_pma_clk_gen3(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_rcvd_clk_gen3(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_rstn_sync2wrfifo_8g(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.rx_sync_hdr(w_hssi_8g_rx_pcs_rx_sync_hdr),
				.rx_we_out_chnl_down(w_hssi_8g_rx_pcs_rx_we_out_chnl_down),
				.rx_we_out_chnl_up(w_hssi_8g_rx_pcs_rx_we_out_chnl_up),
				.rxstatus(w_hssi_8g_rx_pcs_rxstatus),
				.rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.word_align_boundary(w_hssi_8g_rx_pcs_word_align_boundary),
				.wr_clk_rx_phfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_rx_phfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_rx_rmfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_rx_rmfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_data_rx_phfifo(w_hssi_8g_rx_pcs_wr_data_rx_phfifo),
				.wr_data_rx_rmfifo(w_hssi_8g_rx_pcs_wr_data_rx_rmfifo),
				.wr_en_rx_phfifo(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_rx_rmfifo(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_rx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_rx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_rx_phfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo),
				.wr_ptr_rx_rmfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo),
				.wr_rst_n_rx_phfifo(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_rx_rmfifo(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				// INPUTS
				.a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bit_reversal_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.datain({w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0]}),
				.disable_pc_fifo_byte_serdes(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4]),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.eidleinfersel({w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0]}),
				.eios_detected_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.enable_comma_detect(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.gen3_clk_sel(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.hrd_rst(1'b0),
				.inferred_rxvalid_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.pc_fifo_rd_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.pc_fifo_wrdisable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.phystatus_int(w_hssi_pipe_gen1_2_phystatus),
				.phystatus_pcs_gen3(w_hssi_pipe_gen3_phystatus),
				.pipe_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.polarity_inversion(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.rd_data1_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0]}),
				.rd_data2_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0]}),
				.rd_data_rx_phfifo({w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[3]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[3]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.reset_pc_ptrs_asn(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5]),
				.reset_pc_ptrs_in_chnl_down(in_bond_pcs8g_in_bot[12]),
				.reset_pc_ptrs_in_chnl_up(in_bond_pcs8g_in_top[12]),
				.reset_ppm_cntrs_pcs_pma(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7]),
				.rm_fifo_read_enable(1'b0),
				.rm_fifo_write_enable(1'b0),
				.rx_blk_start_pcs_gen3({w_hssi_pipe_gen3_rx_blk_start[3], w_hssi_pipe_gen3_rx_blk_start[2], w_hssi_pipe_gen3_rx_blk_start[1], w_hssi_pipe_gen3_rx_blk_start[0]}),
				.rx_data_pcs_gen3({w_hssi_pipe_gen3_rxd_8gpcs_out[63], w_hssi_pipe_gen3_rxd_8gpcs_out[62], w_hssi_pipe_gen3_rxd_8gpcs_out[61], w_hssi_pipe_gen3_rxd_8gpcs_out[60], w_hssi_pipe_gen3_rxd_8gpcs_out[59], w_hssi_pipe_gen3_rxd_8gpcs_out[58], w_hssi_pipe_gen3_rxd_8gpcs_out[57], w_hssi_pipe_gen3_rxd_8gpcs_out[56], w_hssi_pipe_gen3_rxd_8gpcs_out[55], w_hssi_pipe_gen3_rxd_8gpcs_out[54], w_hssi_pipe_gen3_rxd_8gpcs_out[53], w_hssi_pipe_gen3_rxd_8gpcs_out[52], w_hssi_pipe_gen3_rxd_8gpcs_out[51], w_hssi_pipe_gen3_rxd_8gpcs_out[50], w_hssi_pipe_gen3_rxd_8gpcs_out[49], w_hssi_pipe_gen3_rxd_8gpcs_out[48], w_hssi_pipe_gen3_rxd_8gpcs_out[47], w_hssi_pipe_gen3_rxd_8gpcs_out[46], w_hssi_pipe_gen3_rxd_8gpcs_out[45], w_hssi_pipe_gen3_rxd_8gpcs_out[44], w_hssi_pipe_gen3_rxd_8gpcs_out[43], w_hssi_pipe_gen3_rxd_8gpcs_out[42], w_hssi_pipe_gen3_rxd_8gpcs_out[41], w_hssi_pipe_gen3_rxd_8gpcs_out[40], w_hssi_pipe_gen3_rxd_8gpcs_out[39], w_hssi_pipe_gen3_rxd_8gpcs_out[38], w_hssi_pipe_gen3_rxd_8gpcs_out[37], w_hssi_pipe_gen3_rxd_8gpcs_out[36], w_hssi_pipe_gen3_rxd_8gpcs_out[35], w_hssi_pipe_gen3_rxd_8gpcs_out[34], w_hssi_pipe_gen3_rxd_8gpcs_out[33], w_hssi_pipe_gen3_rxd_8gpcs_out[32], w_hssi_pipe_gen3_rxd_8gpcs_out[31], w_hssi_pipe_gen3_rxd_8gpcs_out[30], w_hssi_pipe_gen3_rxd_8gpcs_out[29], w_hssi_pipe_gen3_rxd_8gpcs_out[28], w_hssi_pipe_gen3_rxd_8gpcs_out[27], w_hssi_pipe_gen3_rxd_8gpcs_out[26], w_hssi_pipe_gen3_rxd_8gpcs_out[25], w_hssi_pipe_gen3_rxd_8gpcs_out[24], w_hssi_pipe_gen3_rxd_8gpcs_out[23], w_hssi_pipe_gen3_rxd_8gpcs_out[22], w_hssi_pipe_gen3_rxd_8gpcs_out[21], w_hssi_pipe_gen3_rxd_8gpcs_out[20], w_hssi_pipe_gen3_rxd_8gpcs_out[19], w_hssi_pipe_gen3_rxd_8gpcs_out[18], w_hssi_pipe_gen3_rxd_8gpcs_out[17], w_hssi_pipe_gen3_rxd_8gpcs_out[16], w_hssi_pipe_gen3_rxd_8gpcs_out[15], w_hssi_pipe_gen3_rxd_8gpcs_out[14], w_hssi_pipe_gen3_rxd_8gpcs_out[13], w_hssi_pipe_gen3_rxd_8gpcs_out[12], w_hssi_pipe_gen3_rxd_8gpcs_out[11], w_hssi_pipe_gen3_rxd_8gpcs_out[10], w_hssi_pipe_gen3_rxd_8gpcs_out[9], w_hssi_pipe_gen3_rxd_8gpcs_out[8], w_hssi_pipe_gen3_rxd_8gpcs_out[7], w_hssi_pipe_gen3_rxd_8gpcs_out[6], w_hssi_pipe_gen3_rxd_8gpcs_out[5], w_hssi_pipe_gen3_rxd_8gpcs_out[4], w_hssi_pipe_gen3_rxd_8gpcs_out[3], w_hssi_pipe_gen3_rxd_8gpcs_out[2], w_hssi_pipe_gen3_rxd_8gpcs_out[1], w_hssi_pipe_gen3_rxd_8gpcs_out[0]}),
				.rx_data_valid_pcs_gen3({w_hssi_pipe_gen3_rxdataskip[3], w_hssi_pipe_gen3_rxdataskip[2], w_hssi_pipe_gen3_rxdataskip[1], w_hssi_pipe_gen3_rxdataskip[0]}),
				.rx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[1], in_bond_pcs8g_in_bot[0]}),
				.rx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[1], in_bond_pcs8g_in_top[0]}),
				.rx_pcs_rst(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.rx_sync_hdr_pcs_gen3({w_hssi_pipe_gen3_rx_sync_hdr[1], w_hssi_pipe_gen3_rx_sync_hdr[0]}),
				.rx_we_in_chnl_down({in_bond_pcs8g_in_bot[5], in_bond_pcs8g_in_bot[4]}),
				.rx_we_in_chnl_up({in_bond_pcs8g_in_top[5], in_bond_pcs8g_in_top[4]}),
				.rxstatus_int({w_hssi_pipe_gen1_2_rxstatus[2], w_hssi_pipe_gen1_2_rxstatus[1], w_hssi_pipe_gen1_2_rxstatus[0]}),
				.rxstatus_pcs_gen3({w_hssi_pipe_gen3_rxstatus[2], w_hssi_pipe_gen3_rxstatus[1], w_hssi_pipe_gen3_rxstatus[0]}),
				.rxvalid_int(w_hssi_pipe_gen1_2_rxvalid),
				.rxvalid_pcs_gen3(w_hssi_pipe_gen3_rxvalid),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.sig_det_from_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_ctrlplane_testbus({w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0]}),
				.tx_div_sync({w_hssi_8g_tx_pcs_tx_div_sync[1], w_hssi_8g_tx_pcs_tx_div_sync[0]}),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.tx_testbus({w_hssi_8g_tx_pcs_tx_testbus[19], w_hssi_8g_tx_pcs_tx_testbus[18], w_hssi_8g_tx_pcs_tx_testbus[17], w_hssi_8g_tx_pcs_tx_testbus[16], w_hssi_8g_tx_pcs_tx_testbus[15], w_hssi_8g_tx_pcs_tx_testbus[14], w_hssi_8g_tx_pcs_tx_testbus[13], w_hssi_8g_tx_pcs_tx_testbus[12], w_hssi_8g_tx_pcs_tx_testbus[11], w_hssi_8g_tx_pcs_tx_testbus[10], w_hssi_8g_tx_pcs_tx_testbus[9], w_hssi_8g_tx_pcs_tx_testbus[8], w_hssi_8g_tx_pcs_tx_testbus[7], w_hssi_8g_tx_pcs_tx_testbus[6], w_hssi_8g_tx_pcs_tx_testbus[5], w_hssi_8g_tx_pcs_tx_testbus[4], w_hssi_8g_tx_pcs_tx_testbus[3], w_hssi_8g_tx_pcs_tx_testbus[2], w_hssi_8g_tx_pcs_tx_testbus[1], w_hssi_8g_tx_pcs_tx_testbus[0]}),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[2]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[2]),
				
				// UNUSED
				.byte_deserializer_pcs_clk_div_by_2_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_wire(),
				.byte_deserializer_pcs_clk_div_by_2_wire(),
				.byte_deserializer_pcs_clk_div_by_4_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_2_reg(),
				.byte_deserializer_pld_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_4_txclk_reg(),
				.pld_8g_a1a2_k1k2_flag_reg(),
				.pld_8g_a1a2_k1k2_flag_txclk_reg(),
				.pld_8g_a1a2_size_reg(),
				.pld_8g_a1a2_size_txclk_reg(),
				.pld_8g_bitloc_rev_en_reg(),
				.pld_8g_bitloc_rev_en_txclk_reg(),
				.pld_8g_byte_rev_en_reg(),
				.pld_8g_byte_rev_en_txclk_reg(),
				.pld_8g_elecidle_reg(),
				.pld_8g_empty_rmf_lowlatency_reg(),
				.pld_8g_empty_rmf_lowlatency_txclk_reg(),
				.pld_8g_empty_rmf_reg(),
				.pld_8g_empty_rmf_txclk_reg(),
				.pld_8g_empty_rx_fifo(),
				.pld_8g_empty_rx_reg(),
				.pld_8g_empty_rx_txclk_reg(),
				.pld_8g_encdt_reg(),
				.pld_8g_encdt_txclk_reg(),
				.pld_8g_full_rmf_reg(),
				.pld_8g_full_rmf_txclk_reg(),
				.pld_8g_full_rx_fifo(),
				.pld_8g_full_rx_reg(),
				.pld_8g_full_rx_txclk_reg(),
				.pld_8g_g3_rx_pld_rst_n_reg(),
				.pld_8g_g3_rx_pld_rst_n_txclk_reg(),
				.pld_8g_rxelecidle_txclk_reg(),
				.pld_8g_rxpolarity_reg(),
				.pld_8g_rxpolarity_txclk_reg(),
				.pld_8g_wa_boundary_reg(),
				.pld_8g_wrdisable_rx_reg(),
				.pld_8g_wrdisable_rx_txclk_reg(),
				.pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_rx_clk_out_8g_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_wire(),
				.pld_rx_control_8g_reg(),
				.pld_rx_control_8g_txclk_reg(),
				.pld_rx_data_8g_reg(),
				.pld_rx_data_8g_txclk_reg(),
				.pld_syncsm_en_reg(),
				.pld_syncsm_en_txclk_reg(),
				.rm_fifo_partial_empty(),
				.rm_fifo_partial_full(),
				.sta_rx_clk2_by2_1(),
				.sta_rx_clk2_by2_1_out(),
				.sta_rx_clk2_by2_2(),
				.sta_rx_clk2_by2_2_out(),
				.sta_rx_clk2_by4_1(),
				.sta_rx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_rx_pcs_a1a2k1k2flag[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_rx_pcs_chnl_test_bus_out[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_clock_to_pld = 1'b0;
				assign w_hssi_8g_rx_pcs_dataout[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_dis_pc_byte = 1'b0;
				assign w_hssi_8g_rx_pcs_eidle_detected = 1'b0;
				assign w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_pma_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_gen2ngen1 = 1'b0;
				assign w_hssi_8g_rx_pcs_parallel_rev_loopback[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_pc_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_pcfifofull = 1'b0;
				assign w_hssi_8g_rx_pcs_phystatus = 1'b0;
				assign w_hssi_8g_rx_pcs_pipe_data[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_full = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clkslip = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_data_valid[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pma_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rxstatus[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_rxvalid = 1'b0;
				assign w_hssi_8g_rx_pcs_signal_detect_out = 1'b0;
				assign w_hssi_8g_rx_pcs_word_align_boundary[4:0] = 5'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79:0] = 80'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31:0] = 32'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_rmfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_tx_pcs
			twentynm_hssi_8g_tx_pcs #(
				.auto_speed_nego_gen2(hssi_8g_tx_pcs_auto_speed_nego_gen2),
				.bit_reversal(hssi_8g_tx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_tx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_tx_pcs_bypass_pipeline_reg),
				.byte_serializer(hssi_8g_tx_pcs_byte_serializer),
				.clock_gate_bs_enc(hssi_8g_tx_pcs_clock_gate_bs_enc),
				.clock_gate_dw_fifowr(hssi_8g_tx_pcs_clock_gate_dw_fifowr),
				.clock_gate_fiford(hssi_8g_tx_pcs_clock_gate_fiford),
				.clock_gate_sw_fifowr(hssi_8g_tx_pcs_clock_gate_sw_fifowr),
				.clock_observation_in_pld_core(hssi_8g_tx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_tx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_tx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_tx_pcs_ctrl_plane_bonding_distribution),
				.data_selection_8b10b_encoder_input(hssi_8g_tx_pcs_data_selection_8b10b_encoder_input),
				.dynamic_clk_switch(hssi_8g_tx_pcs_dynamic_clk_switch),
				.eightb_tenb_disp_ctrl(hssi_8g_tx_pcs_eightb_tenb_disp_ctrl),
				.eightb_tenb_encoder(hssi_8g_tx_pcs_eightb_tenb_encoder),
				.force_echar(hssi_8g_tx_pcs_force_echar),
				.force_kchar(hssi_8g_tx_pcs_force_kchar),
				.gen3_tx_clk_sel(hssi_8g_tx_pcs_gen3_tx_clk_sel),
				.gen3_tx_pipe_clk_sel(hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel),
				.hip_mode(hssi_8g_tx_pcs_hip_mode),
				.pcs_bypass(hssi_8g_tx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_tx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_tx_pcs_phase_compensation_fifo),
				.phfifo_write_clk_sel(hssi_8g_tx_pcs_phfifo_write_clk_sel),
				.pma_dw(hssi_8g_tx_pcs_pma_dw),
				.prot_mode(hssi_8g_tx_pcs_prot_mode),
				.reconfig_settings(hssi_8g_tx_pcs_reconfig_settings),
				.refclk_b_clk_sel(hssi_8g_tx_pcs_refclk_b_clk_sel),
				.revloop_back_rm(hssi_8g_tx_pcs_revloop_back_rm),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_tx_pcs_sup_mode),
				.symbol_swap(hssi_8g_tx_pcs_symbol_swap),
				.tx_bitslip(hssi_8g_tx_pcs_tx_bitslip),
				.tx_compliance_controlled_disparity(hssi_8g_tx_pcs_tx_compliance_controlled_disparity),
				.tx_fast_pld_reg(hssi_8g_tx_pcs_tx_fast_pld_reg),
				.txclk_freerun(hssi_8g_tx_pcs_txclk_freerun),
				.txpcs_urst(hssi_8g_tx_pcs_txpcs_urst)
			) inst_twentynm_hssi_8g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_8g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_tx_pcs_blockselect),
				.clk_out(w_hssi_8g_tx_pcs_clk_out),
				.clk_out_gen3(w_hssi_8g_tx_pcs_clk_out_gen3),
				.dataout(w_hssi_8g_tx_pcs_dataout),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.fifo_select_out_chnl_down(w_hssi_8g_tx_pcs_fifo_select_out_chnl_down),
				.fifo_select_out_chnl_up(w_hssi_8g_tx_pcs_fifo_select_out_chnl_up),
				.g3_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.g3_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
				.non_gray_eidleinfersel(w_hssi_8g_tx_pcs_non_gray_eidleinfersel),
				.ph_fifo_overflow(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.ph_fifo_underflow(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.phfifo_txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.phfifo_txmargin(w_hssi_8g_tx_pcs_phfifo_txmargin),
				.phfifo_txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				.pipe_en_rev_parallel_lpbk_out(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.pipe_power_down_out(w_hssi_8g_tx_pcs_pipe_power_down_out),
				.pipe_tx_clk_out_gen3(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pmaif_asn_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.rd_enable_out_chnl_down(w_hssi_8g_tx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_tx_pcs_rd_enable_out_chnl_up),
				.rd_ptr_tx_phfifo(w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rxpolarity_int(w_hssi_8g_tx_pcs_rxpolarity_int),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.tx_blk_start_out(w_hssi_8g_tx_pcs_tx_blk_start_out),
				.tx_clk_out_8g_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.tx_ctrlplane_testbus(w_hssi_8g_tx_pcs_tx_ctrlplane_testbus),
				.tx_data_out(w_hssi_8g_tx_pcs_tx_data_out),
				.tx_data_valid_out(w_hssi_8g_tx_pcs_tx_data_valid_out),
				.tx_datak_out(w_hssi_8g_tx_pcs_tx_datak_out),
				.tx_detect_rxloopback_int(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.tx_div_sync(w_hssi_8g_tx_pcs_tx_div_sync),
				.tx_div_sync_out_chnl_down(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down),
				.tx_div_sync_out_chnl_up(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up),
				.tx_pipe_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.tx_pipe_electidle(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_soft_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.tx_sync_hdr_out(w_hssi_8g_tx_pcs_tx_sync_hdr_out),
				.tx_testbus(w_hssi_8g_tx_pcs_tx_testbus),
				.txcompliance_out(w_hssi_8g_tx_pcs_txcompliance_out),
				.txelecidle_out(w_hssi_8g_tx_pcs_txelecidle_out),
				.wr_clk_tx_phfifo_dw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_tx_phfifo_sw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_data_tx_phfifo(w_hssi_8g_tx_pcs_wr_data_tx_phfifo),
				.wr_en_tx_phfifo(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_tx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_tx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_tx_phfifo(w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo),
				.wr_rst_n_tx_phfifo(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bitslip_boundary_select({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0]}),
				.clk_sel_gen3(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.coreclk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.datain({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.detectrxloopin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidleinfersel({w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0]}),
				.en_rev_parallel_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.fifo_select_in_chnl_down({in_bond_pcs8g_in_bot[11], in_bond_pcs8g_in_bot[10]}),
				.fifo_select_in_chnl_up({in_bond_pcs8g_in_top[11], in_bond_pcs8g_in_top[10]}),
				.hrdrst(1'b0),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.ph_fifo_rd_disable(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.pipe_en_rev_parallel_lpbk_in(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.pipe_tx_deemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.pipe_tx_margin({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0]}),
				.powerdn({w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0]}),
				.rate_switch(w_hssi_8g_rx_pcs_gen2ngen1),
				.rd_data_tx_phfifo({w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[9]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[9]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.rev_parallel_lpbk_data({w_hssi_8g_rx_pcs_parallel_rev_loopback[19], w_hssi_8g_rx_pcs_parallel_rev_loopback[18], w_hssi_8g_rx_pcs_parallel_rev_loopback[17], w_hssi_8g_rx_pcs_parallel_rev_loopback[16], w_hssi_8g_rx_pcs_parallel_rev_loopback[15], w_hssi_8g_rx_pcs_parallel_rev_loopback[14], w_hssi_8g_rx_pcs_parallel_rev_loopback[13], w_hssi_8g_rx_pcs_parallel_rev_loopback[12], w_hssi_8g_rx_pcs_parallel_rev_loopback[11], w_hssi_8g_rx_pcs_parallel_rev_loopback[10], w_hssi_8g_rx_pcs_parallel_rev_loopback[9], w_hssi_8g_rx_pcs_parallel_rev_loopback[8], w_hssi_8g_rx_pcs_parallel_rev_loopback[7], w_hssi_8g_rx_pcs_parallel_rev_loopback[6], w_hssi_8g_rx_pcs_parallel_rev_loopback[5], w_hssi_8g_rx_pcs_parallel_rev_loopback[4], w_hssi_8g_rx_pcs_parallel_rev_loopback[3], w_hssi_8g_rx_pcs_parallel_rev_loopback[2], w_hssi_8g_rx_pcs_parallel_rev_loopback[1], w_hssi_8g_rx_pcs_parallel_rev_loopback[0]}),
				.rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.tx_blk_start({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0]}),
				.tx_data_valid({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0]}),
				.tx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[7], in_bond_pcs8g_in_bot[6]}),
				.tx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[7], in_bond_pcs8g_in_top[6]}),
				.tx_pcs_reset(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.tx_sync_hdr({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0]}),
				.txd_fast_reg({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0]}),
				.txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[8]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[8]),
				.wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				
				// UNUSED
				.byte_serializer_pcs_clk_div_by_2_reg(),
				.byte_serializer_pcs_clk_div_by_2_wire(),
				.byte_serializer_pcs_clk_div_by_4_reg(),
				.byte_serializer_pld_clk_div_by_2_reg(),
				.byte_serializer_pld_clk_div_by_4_reg(),
				.pld_8g_empty_tx_fifo(),
				.pld_8g_empty_tx_reg(),
				.pld_8g_full_tx_fifo(),
				.pld_8g_full_tx_reg(),
				.pld_8g_g3_tx_pld_rst_n_reg(),
				.pld_8g_rddisable_tx_reg(),
				.pld_8g_tx_boundary_sel_reg(),
				.pld_pcs_tx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_tx_clk_out_8g_wire(),
				.pld_tx_data_8g_fifo(),
				.pld_tx_data_lo_8g_reg(),
				.sta_tx_clk2_by2_1(),
				.sta_tx_clk2_by2_1_out(),
				.sta_tx_clk2_by4_1(),
				.sta_tx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_dataout[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_dyn_clk_switch_n = 1'b1;		// Override default tieoff
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_g3_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_overflow = 1'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_underflow = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txdeemph = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txmargin[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txswing = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_power_down_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_pmaif_asn_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_refclk_b = 1'b0;
				assign w_hssi_8g_tx_pcs_refclk_b_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_rxpolarity_int = 1'b0;
				assign w_hssi_8g_tx_pcs_soft_reset_wclk1_n = 1'b0;
				assign w_hssi_8g_tx_pcs_sw_fifo_wr_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_blk_start_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_tx_data_out[31:0] = 32'b0;
				assign w_hssi_8g_tx_pcs_tx_data_valid_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_datak_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_detect_rxloopback_int = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_electidle = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_sync_hdr_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_txcompliance_out = 1'b0;
				assign w_hssi_8g_tx_pcs_txelecidle_out = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63:0] = 64'b0;
				assign w_hssi_8g_tx_pcs_wr_en_tx_phfifo = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pcs_pma_interface
			twentynm_hssi_common_pcs_pma_interface #(
				.asn_clk_enable(hssi_common_pcs_pma_interface_asn_clk_enable),
				.asn_enable(hssi_common_pcs_pma_interface_asn_enable),
				.block_sel(hssi_common_pcs_pma_interface_block_sel),
				.bypass_early_eios(hssi_common_pcs_pma_interface_bypass_early_eios),
				.bypass_pcie_switch(hssi_common_pcs_pma_interface_bypass_pcie_switch),
				.bypass_pma_ltr(hssi_common_pcs_pma_interface_bypass_pma_ltr),
				.bypass_pma_sw_done(hssi_common_pcs_pma_interface_bypass_pma_sw_done),
				.bypass_ppm_lock(hssi_common_pcs_pma_interface_bypass_ppm_lock),
				.bypass_send_syncp_fbkp(hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp),
				.bypass_txdetectrx(hssi_common_pcs_pma_interface_bypass_txdetectrx),
				.cdr_control(hssi_common_pcs_pma_interface_cdr_control),
				.cid_enable(hssi_common_pcs_pma_interface_cid_enable),
				.cp_cons_sel(hssi_common_pcs_pma_interface_cp_cons_sel),
				.cp_dwn_mstr(hssi_common_pcs_pma_interface_cp_dwn_mstr),
				.cp_up_mstr(hssi_common_pcs_pma_interface_cp_up_mstr),
				.ctrl_plane_bonding(hssi_common_pcs_pma_interface_ctrl_plane_bonding),
				.data_mask_count(hssi_common_pcs_pma_interface_data_mask_count),
				.data_mask_count_multi(hssi_common_pcs_pma_interface_data_mask_count_multi),
				.dft_observation_clock_selection(hssi_common_pcs_pma_interface_dft_observation_clock_selection),
				.early_eios_counter(hssi_common_pcs_pma_interface_early_eios_counter),
				.force_freqdet(hssi_common_pcs_pma_interface_force_freqdet),
				.free_run_clk_enable(hssi_common_pcs_pma_interface_free_run_clk_enable),
				.ignore_sigdet_g23(hssi_common_pcs_pma_interface_ignore_sigdet_g23),
				.pc_en_counter(hssi_common_pcs_pma_interface_pc_en_counter),
				.pc_rst_counter(hssi_common_pcs_pma_interface_pc_rst_counter),
				.pcie_hip_mode(hssi_common_pcs_pma_interface_pcie_hip_mode),
				.ph_fifo_reg_mode(hssi_common_pcs_pma_interface_ph_fifo_reg_mode),
				.phfifo_flush_wait(hssi_common_pcs_pma_interface_phfifo_flush_wait),
				.pipe_if_g3pcs(hssi_common_pcs_pma_interface_pipe_if_g3pcs),
				.pma_done_counter(hssi_common_pcs_pma_interface_pma_done_counter),
				.pma_if_dft_en(hssi_common_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_common_pcs_pma_interface_pma_if_dft_val),
				.ppm_cnt_rst(hssi_common_pcs_pma_interface_ppm_cnt_rst),
				.ppm_deassert_early(hssi_common_pcs_pma_interface_ppm_deassert_early),
				.ppm_det_buckets(hssi_common_pcs_pma_interface_ppm_det_buckets),
				.ppm_gen1_2_cnt(hssi_common_pcs_pma_interface_ppm_gen1_2_cnt),
				.ppm_post_eidle_delay(hssi_common_pcs_pma_interface_ppm_post_eidle_delay),
				.ppmsel(hssi_common_pcs_pma_interface_ppmsel),
				.prot_mode(hssi_common_pcs_pma_interface_prot_mode),
				.reconfig_settings(hssi_common_pcs_pma_interface_reconfig_settings),
				.rxvalid_mask(hssi_common_pcs_pma_interface_rxvalid_mask),
				.sigdet_wait_counter(hssi_common_pcs_pma_interface_sigdet_wait_counter),
				.sigdet_wait_counter_multi(hssi_common_pcs_pma_interface_sigdet_wait_counter_multi),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sim_mode(hssi_common_pcs_pma_interface_sim_mode),
				.spd_chg_rst_wait_cnt_en(hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en),
				.sup_mode(hssi_common_pcs_pma_interface_sup_mode),
				.testout_sel(hssi_common_pcs_pma_interface_testout_sel),
				.wait_clk_on_off_timer(hssi_common_pcs_pma_interface_wait_clk_on_off_timer),
				.wait_pipe_synchronizing(hssi_common_pcs_pma_interface_wait_pipe_synchronizing),
				.wait_send_syncp_fbkp(hssi_common_pcs_pma_interface_wait_send_syncp_fbkp)
			) inst_twentynm_hssi_common_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_common_pcs_pma_interface_blockselect),
				.int_pmaif_8g_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in),
				.int_pmaif_8g_eios_detected(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.int_pmaif_8g_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.int_pmaif_8g_power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.int_pmaif_g3_pcs_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in),
				.int_pmaif_pldif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pmaif_pldif_pcie_sw_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done),
				.int_pmaif_pldif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pmaif_pldif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pmaif_pldif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pmaif_pldif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pmaif_pldif_pma_reserved_in(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in),
				.int_pmaif_pldif_test_out(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out),
				.int_pmaif_pldif_testbus(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus),
				.pma_adapt_start(w_hssi_common_pcs_pma_interface_pma_adapt_start),
				.pma_atpg_los_en_n(w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n),
				.pma_csr_test_dis(w_hssi_common_pcs_pma_interface_pma_csr_test_dis),
				.pma_current_coeff(w_hssi_common_pcs_pma_interface_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_common_pcs_pma_interface_pma_current_rxpreset),
				.pma_early_eios(w_hssi_common_pcs_pma_interface_pma_early_eios),
				.pma_interface_select(w_hssi_common_pcs_pma_interface_pma_interface_select),
				.pma_ltd_b(w_hssi_common_pcs_pma_interface_pma_ltd_b),
				.pma_ltr(w_hssi_common_pcs_pma_interface_pma_ltr),
				.pma_nfrzdrv(w_hssi_common_pcs_pma_interface_pma_nfrzdrv),
				.pma_nrpi_freeze(w_hssi_common_pcs_pma_interface_pma_nrpi_freeze),
				.pma_pcie_switch(w_hssi_common_pcs_pma_interface_pma_pcie_switch),
				.pma_ppm_lock(w_hssi_common_pcs_pma_interface_pma_ppm_lock),
				.pma_reserved_out(w_hssi_common_pcs_pma_interface_pma_reserved_out),
				.pma_rs_lpbk_b(w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b),
				.pma_rx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup),
				.pma_scan_mode_n(w_hssi_common_pcs_pma_interface_pma_scan_mode_n),
				.pma_scan_shift_n(w_hssi_common_pcs_pma_interface_pma_scan_shift_n),
				.pma_tx_bitslip(w_hssi_common_pcs_pma_interface_pma_tx_bitslip),
				.pma_tx_bonding_rstb(w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb),
				.pma_tx_qpi_pulldn(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn),
				.pma_tx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup),
				.pma_tx_txdetectrx(w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx),
				.pmaif_bundling_out_down(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down),
				.pmaif_bundling_out_up(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_8g_current_coeff({w_hssi_pipe_gen1_2_current_coeff[17], w_hssi_pipe_gen1_2_current_coeff[16], w_hssi_pipe_gen1_2_current_coeff[15], w_hssi_pipe_gen1_2_current_coeff[14], w_hssi_pipe_gen1_2_current_coeff[13], w_hssi_pipe_gen1_2_current_coeff[12], w_hssi_pipe_gen1_2_current_coeff[11], w_hssi_pipe_gen1_2_current_coeff[10], w_hssi_pipe_gen1_2_current_coeff[9], w_hssi_pipe_gen1_2_current_coeff[8], w_hssi_pipe_gen1_2_current_coeff[7], w_hssi_pipe_gen1_2_current_coeff[6], w_hssi_pipe_gen1_2_current_coeff[5], w_hssi_pipe_gen1_2_current_coeff[4], w_hssi_pipe_gen1_2_current_coeff[3], w_hssi_pipe_gen1_2_current_coeff[2], w_hssi_pipe_gen1_2_current_coeff[1], w_hssi_pipe_gen1_2_current_coeff[0]}),
				.int_pmaif_8g_eios_det({w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0]}),
				.int_pmaif_8g_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.int_pmaif_8g_rev_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.int_pmaif_8g_tx_clk_out_gen3(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.int_pmaif_8g_txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				.int_pmaif_g3_eios_det({w_hssi_gen3_rx_pcs_ei_det_int, w_hssi_gen3_rx_pcs_ei_partial_det_int, w_hssi_gen3_rx_pcs_i_det_int}),
				.int_pmaif_g3_pma_current_coeff({w_hssi_pipe_gen3_pma_current_coeff[17], w_hssi_pipe_gen3_pma_current_coeff[16], w_hssi_pipe_gen3_pma_current_coeff[15], w_hssi_pipe_gen3_pma_current_coeff[14], w_hssi_pipe_gen3_pma_current_coeff[13], w_hssi_pipe_gen3_pma_current_coeff[12], w_hssi_pipe_gen3_pma_current_coeff[11], w_hssi_pipe_gen3_pma_current_coeff[10], w_hssi_pipe_gen3_pma_current_coeff[9], w_hssi_pipe_gen3_pma_current_coeff[8], w_hssi_pipe_gen3_pma_current_coeff[7], w_hssi_pipe_gen3_pma_current_coeff[6], w_hssi_pipe_gen3_pma_current_coeff[5], w_hssi_pipe_gen3_pma_current_coeff[4], w_hssi_pipe_gen3_pma_current_coeff[3], w_hssi_pipe_gen3_pma_current_coeff[2], w_hssi_pipe_gen3_pma_current_coeff[1], w_hssi_pipe_gen3_pma_current_coeff[0]}),
				.int_pmaif_g3_pma_current_rxpreset({w_hssi_pipe_gen3_pma_current_rxpreset[2], w_hssi_pipe_gen3_pma_current_rxpreset[1], w_hssi_pipe_gen3_pma_current_rxpreset[0]}),
				.int_pmaif_g3_pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.int_pmaif_g3_rev_lpbk(w_hssi_pipe_gen3_rev_lpbk_int),
				.int_pmaif_pldif_8g_tx_pld_rstn(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pmaif_pldif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pmaif_pldif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pmaif_pldif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pmaif_pldif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pmaif_pldif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pmaif_pldif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pmaif_pldif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pmaif_pldif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pmaif_pldif_pcie_switch({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0]}),
				.int_pmaif_pldif_pma_reserved_out({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0]}),
				.int_pmaif_pldif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pmaif_pldif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pmaif_pldif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pmaif_pldif_rate({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0]}),
				.int_pmaif_pldif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pmaif_pldif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pmaif_pldif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.int_pmaif_pldif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pmaif_pldif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pmaif_pldif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pmaif_pldif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pmaif_pldif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pmaif_pldif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.int_tx_dft_obsrv_clk({w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0]}),
				.iocsr_clk(in_iocsr_clk),
				.iocsr_config({in_iocsr_config[5], in_iocsr_config[4], in_iocsr_config[3], in_iocsr_config[2], in_iocsr_config[1], in_iocsr_config[0]}),
				.iocsr_rdy(in_iocsr_rdy),
				.iocsr_rdy_dly(in_iocsr_rdy_dly),
				.pma_adapt_done(in_pma_adapt_done),
				.pma_clklow(in_pma_clklow),
				.pma_fref(in_pma_fref),
				.pma_hclk(in_pma_hclk),
				.pma_pcie_sw_done({in_pma_pcie_sw_done[1], in_pma_pcie_sw_done[0]}),
				.pma_pfdmode_lock(in_pma_pfdmode_lock),
				.pma_reserved_in({in_pma_reserved_in[4], in_pma_reserved_in[3], in_pma_reserved_in[2], in_pma_reserved_in[1], in_pma_reserved_in[0]}),
				.pma_signal_det(in_pma_signal_det),
				.pma_testbus({in_pma_testbus[7], in_pma_testbus[6], in_pma_testbus[5], in_pma_testbus[4], in_pma_testbus[3], in_pma_testbus[2], in_pma_testbus[1], in_pma_testbus[0]}),
				.pmaif_bundling_in_down({in_bond_pmaif_in_bot[11], in_bond_pmaif_in_bot[10], in_bond_pmaif_in_bot[9], in_bond_pmaif_in_bot[8], in_bond_pmaif_in_bot[7], in_bond_pmaif_in_bot[6], in_bond_pmaif_in_bot[5], in_bond_pmaif_in_bot[4], in_bond_pmaif_in_bot[3], in_bond_pmaif_in_bot[2], in_bond_pmaif_in_bot[1], in_bond_pmaif_in_bot[0]}),
				.pmaif_bundling_in_up({in_bond_pmaif_in_top[11], in_bond_pmaif_in_top[10], in_bond_pmaif_in_top[9], in_bond_pmaif_in_top[8], in_bond_pmaif_in_top[7], in_bond_pmaif_in_top[6], in_bond_pmaif_in_top[5], in_bond_pmaif_in_top[4], in_bond_pmaif_in_top[3], in_bond_pmaif_in_top[2], in_bond_pmaif_in_top[1], in_bond_pmaif_in_top[0]}),
				.rx_pmaif_test_out({w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0]}),
				.rx_prbs_ver_test({w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0]}),
				.tx_prbs_gen_test({w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0]}),
				.uhsif_test_out_1({w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0]}),
				.uhsif_test_out_2({w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0]}),
				.uhsif_test_out_3({w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0]}),
				
				// UNUSED
				.int_pmaif_avmm_iocsr_clk(),
				.int_pmaif_avmm_iocsr_config(),
				.int_pmaif_avmm_iocsr_rdy(),
				.int_pmaif_avmm_iocsr_rdy_dly(),
				.int_pmaif_pldif_interface_select(),
				.pma_tx_pma_syncp(),
				.sta_pma_hclk_by2()
			);
		end // if generate
		else begin
				assign w_hssi_common_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19:0] = 20'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_pma_adapt_start = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_csr_test_dis = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pcs_pma_interface_pma_early_eios = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_interface_select[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltd_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltr = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nfrzdrv = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nrpi_freeze = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ppm_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_tx_bitslip = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx = in_pld_pma_txdetectrx;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11:0] = 12'b0;
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11:0] = 12'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pld_pcs_interface
			twentynm_hssi_common_pld_pcs_interface #(
				.dft_clk_out_en(hssi_common_pld_pcs_interface_dft_clk_out_en),
				.dft_clk_out_sel(hssi_common_pld_pcs_interface_dft_clk_out_sel),
				.hrdrstctrl_en(hssi_common_pld_pcs_interface_hrdrstctrl_en),
				.pcs_testbus_block_sel(hssi_common_pld_pcs_interface_pcs_testbus_block_sel),
				.reconfig_settings(hssi_common_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm2" )       //PARAM_HIDE
			) inst_twentynm_hssi_common_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_common_pld_pcs_interface_blockselect),
				.hip_cmn_clk(w_hssi_common_pld_pcs_interface_hip_cmn_clk),
				.hip_cmn_ctrl(w_hssi_common_pld_pcs_interface_hip_cmn_ctrl),
				.hip_iocsr_rdy(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy),
				.hip_iocsr_rdy_dly(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly),
				.hip_nfrzdrv(w_hssi_common_pld_pcs_interface_hip_nfrzdrv),
				.hip_npor(w_hssi_common_pld_pcs_interface_hip_npor),
				.hip_usermode(w_hssi_common_pld_pcs_interface_hip_usermode),
				.int_pldif_10g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.int_pldif_10g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.int_pldif_8g_eidleinfersel(w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel),
				.int_pldif_8g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.int_pldif_8g_refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.int_pldif_8g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.int_pldif_g3_current_coeff(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff),
				.int_pldif_g3_current_rxpreset(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset),
				.int_pldif_krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.int_pldif_krfec_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.int_pldif_krfec_scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				.int_pldif_mem_atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.int_pldif_mem_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.int_pldif_pmaif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pldif_pmaif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pldif_pmaif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pldif_pmaif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pldif_pmaif_eye_monitor(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor),
				.int_pldif_pmaif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pldif_pmaif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pldif_pmaif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pldif_pmaif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pldif_pmaif_pcie_switch(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch),
				.int_pldif_pmaif_pma_reserved_out(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out),
				.int_pldif_pmaif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pldif_pmaif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pldif_pmaif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pldif_pmaif_rate(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate),
				.int_pldif_pmaif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pldif_pmaif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pldif_pmaif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pldif_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_pldif_pmaif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pldif_pmaif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pldif_pmaif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pldif_pmaif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pldif_pmaif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pldif_pmaif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pldif_pmaif_uhsif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.pld_pma_adapt_done(w_hssi_common_pld_pcs_interface_pld_pma_adapt_done),
				.pld_pma_clklow(w_hssi_common_pld_pcs_interface_pld_pma_clklow),
				.pld_pma_fref(w_hssi_common_pld_pcs_interface_pld_pma_fref),
				.pld_pma_hclk(w_hssi_common_pld_pcs_interface_pld_pma_hclk),
				.pld_pma_pcie_sw_done(w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done),
				.pld_pma_pfdmode_lock(w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock),
				.pld_pma_reserved_in(w_hssi_common_pld_pcs_interface_pld_pma_reserved_in),
				.pld_pma_rx_detect_valid(w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid),
				.pld_pma_rx_found(w_hssi_common_pld_pcs_interface_pld_pma_rx_found),
				.pld_pma_rxpll_lock(w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock),
				.pld_pma_testbus(w_hssi_common_pld_pcs_interface_pld_pma_testbus),
				.pld_pmaif_mask_tx_pll(w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll),
				.pld_reserved_out(w_hssi_common_pld_pcs_interface_pld_reserved_out),
				.pld_test_data(w_hssi_common_pld_pcs_interface_pld_test_data),
				.pld_uhsif_lock(w_hssi_common_pld_pcs_interface_pld_uhsif_lock),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.int_pldif_10g_test_data({w_hssi_10g_tx_pcs_tx_test_data[19], w_hssi_10g_tx_pcs_tx_test_data[18], w_hssi_10g_tx_pcs_tx_test_data[17], w_hssi_10g_tx_pcs_tx_test_data[16], w_hssi_10g_tx_pcs_tx_test_data[15], w_hssi_10g_tx_pcs_tx_test_data[14], w_hssi_10g_tx_pcs_tx_test_data[13], w_hssi_10g_tx_pcs_tx_test_data[12], w_hssi_10g_tx_pcs_tx_test_data[11], w_hssi_10g_tx_pcs_tx_test_data[10], w_hssi_10g_tx_pcs_tx_test_data[9], w_hssi_10g_tx_pcs_tx_test_data[8], w_hssi_10g_tx_pcs_tx_test_data[7], w_hssi_10g_tx_pcs_tx_test_data[6], w_hssi_10g_tx_pcs_tx_test_data[5], w_hssi_10g_tx_pcs_tx_test_data[4], w_hssi_10g_tx_pcs_tx_test_data[3], w_hssi_10g_tx_pcs_tx_test_data[2], w_hssi_10g_tx_pcs_tx_test_data[1], w_hssi_10g_tx_pcs_tx_test_data[0]}),
				.int_pldif_10g_tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.int_pldif_8g_chnl_test_bus_out({w_hssi_8g_rx_pcs_chnl_test_bus_out[19], w_hssi_8g_rx_pcs_chnl_test_bus_out[18], w_hssi_8g_rx_pcs_chnl_test_bus_out[17], w_hssi_8g_rx_pcs_chnl_test_bus_out[16], w_hssi_8g_rx_pcs_chnl_test_bus_out[15], w_hssi_8g_rx_pcs_chnl_test_bus_out[14], w_hssi_8g_rx_pcs_chnl_test_bus_out[13], w_hssi_8g_rx_pcs_chnl_test_bus_out[12], w_hssi_8g_rx_pcs_chnl_test_bus_out[11], w_hssi_8g_rx_pcs_chnl_test_bus_out[10], w_hssi_8g_rx_pcs_chnl_test_bus_out[9], w_hssi_8g_rx_pcs_chnl_test_bus_out[8], w_hssi_8g_rx_pcs_chnl_test_bus_out[7], w_hssi_8g_rx_pcs_chnl_test_bus_out[6], w_hssi_8g_rx_pcs_chnl_test_bus_out[5], w_hssi_8g_rx_pcs_chnl_test_bus_out[4], w_hssi_8g_rx_pcs_chnl_test_bus_out[3], w_hssi_8g_rx_pcs_chnl_test_bus_out[2], w_hssi_8g_rx_pcs_chnl_test_bus_out[1], w_hssi_8g_rx_pcs_chnl_test_bus_out[0]}),
				.int_pldif_8g_rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.int_pldif_8g_tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.int_pldif_g3_test_out({w_hssi_pipe_gen3_test_out[19], w_hssi_pipe_gen3_test_out[18], w_hssi_pipe_gen3_test_out[17], w_hssi_pipe_gen3_test_out[16], w_hssi_pipe_gen3_test_out[15], w_hssi_pipe_gen3_test_out[14], w_hssi_pipe_gen3_test_out[13], w_hssi_pipe_gen3_test_out[12], w_hssi_pipe_gen3_test_out[11], w_hssi_pipe_gen3_test_out[10], w_hssi_pipe_gen3_test_out[9], w_hssi_pipe_gen3_test_out[8], w_hssi_pipe_gen3_test_out[7], w_hssi_pipe_gen3_test_out[6], w_hssi_pipe_gen3_test_out[5], w_hssi_pipe_gen3_test_out[4], w_hssi_pipe_gen3_test_out[3], w_hssi_pipe_gen3_test_out[2], w_hssi_pipe_gen3_test_out[1], w_hssi_pipe_gen3_test_out[0]}),
				.int_pldif_krfec_test_data({w_hssi_krfec_tx_pcs_tx_test_data[19], w_hssi_krfec_tx_pcs_tx_test_data[18], w_hssi_krfec_tx_pcs_tx_test_data[17], w_hssi_krfec_tx_pcs_tx_test_data[16], w_hssi_krfec_tx_pcs_tx_test_data[15], w_hssi_krfec_tx_pcs_tx_test_data[14], w_hssi_krfec_tx_pcs_tx_test_data[13], w_hssi_krfec_tx_pcs_tx_test_data[12], w_hssi_krfec_tx_pcs_tx_test_data[11], w_hssi_krfec_tx_pcs_tx_test_data[10], w_hssi_krfec_tx_pcs_tx_test_data[9], w_hssi_krfec_tx_pcs_tx_test_data[8], w_hssi_krfec_tx_pcs_tx_test_data[7], w_hssi_krfec_tx_pcs_tx_test_data[6], w_hssi_krfec_tx_pcs_tx_test_data[5], w_hssi_krfec_tx_pcs_tx_test_data[4], w_hssi_krfec_tx_pcs_tx_test_data[3], w_hssi_krfec_tx_pcs_tx_test_data[2], w_hssi_krfec_tx_pcs_tx_test_data[1], w_hssi_krfec_tx_pcs_tx_test_data[0]}),
				.int_pldif_pmaif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pldif_pmaif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pldif_pmaif_pcie_sw_done({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0]}),
				.int_pldif_pmaif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pldif_pmaif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pldif_pmaif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pldif_pmaif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pldif_pmaif_pma_reserved_in({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0]}),
				.int_pldif_pmaif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pldif_pmaif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_test_out({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0]}),
				.int_pldif_pmaif_testbus({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0]}),
				.int_pldif_pmaif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.pld_8g_eidleinfersel({in_pld_8g_eidleinfersel[2], in_pld_8g_eidleinfersel[1], in_pld_8g_eidleinfersel[0]}),
				.pld_8g_refclk_dig2(in_pld_8g_refclk_dig2),
				.pld_atpg_los_en_n(in_pld_atpg_los_en_n),
				.pld_g3_current_coeff({in_pld_g3_current_coeff[17], in_pld_g3_current_coeff[16], in_pld_g3_current_coeff[15], in_pld_g3_current_coeff[14], in_pld_g3_current_coeff[13], in_pld_g3_current_coeff[12], in_pld_g3_current_coeff[11], in_pld_g3_current_coeff[10], in_pld_g3_current_coeff[9], in_pld_g3_current_coeff[8], in_pld_g3_current_coeff[7], in_pld_g3_current_coeff[6], in_pld_g3_current_coeff[5], in_pld_g3_current_coeff[4], in_pld_g3_current_coeff[3], in_pld_g3_current_coeff[2], in_pld_g3_current_coeff[1], in_pld_g3_current_coeff[0]}),
				.pld_g3_current_rxpreset({in_pld_g3_current_rxpreset[2], in_pld_g3_current_rxpreset[1], in_pld_g3_current_rxpreset[0]}),
				.pld_ltr(in_pld_ltr),
				.pld_mem_krfec_atpg_rst_n(in_pld_mem_krfec_atpg_rst_n),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pcs_refclk_dig(in_pld_pcs_refclk_dig),
				.pld_pma_adapt_start(in_pld_pma_adapt_start),
				.pld_pma_csr_test_dis(in_pld_pma_csr_test_dis),
				.pld_pma_early_eios(in_pld_pma_early_eios),
				.pld_pma_eye_monitor({in_pld_pma_eye_monitor[5], in_pld_pma_eye_monitor[4], in_pld_pma_eye_monitor[3], in_pld_pma_eye_monitor[2], in_pld_pma_eye_monitor[1], in_pld_pma_eye_monitor[0]}),
				.pld_pma_ltd_b(in_pld_pma_ltd_b),
				.pld_pma_nrpi_freeze(in_pld_pma_nrpi_freeze),
				.pld_pma_pcie_switch({in_pld_pma_pcie_switch[1], in_pld_pma_pcie_switch[0]}),
				.pld_pma_ppm_lock(in_pld_pma_ppm_lock),
				.pld_pma_reserved_out({in_pld_pma_reserved_out[4], in_pld_pma_reserved_out[3], in_pld_pma_reserved_out[2], in_pld_pma_reserved_out[1], in_pld_pma_reserved_out[0]}),
				.pld_pma_rs_lpbk_b(in_pld_pma_rs_lpbk_b),
				.pld_pma_rx_qpi_pullup(in_pld_pma_rx_qpi_pullup),
				.pld_pma_tx_bitslip(in_pld_pma_tx_bitslip),
				.pld_pma_tx_bonding_rstb(in_pld_pma_tx_bonding_rstb),
				.pld_pma_tx_qpi_pulldn(in_pld_pma_tx_qpi_pulldn),
				.pld_pma_tx_qpi_pullup(in_pld_pma_tx_qpi_pullup),
				.pld_pma_txdetectrx(in_pld_pma_txdetectrx),
				.pld_rate({in_pld_rate[1], in_pld_rate[0]}),
				.pld_reserved_in({in_pld_reserved_in[9], in_pld_reserved_in[8], in_pld_reserved_in[7], in_pld_reserved_in[6], in_pld_reserved_in[5], in_pld_reserved_in[4], in_pld_reserved_in[3], in_pld_reserved_in[2], in_pld_reserved_in[1], in_pld_reserved_in[0]}),
				.pld_scan_mode_n(in_pld_scan_mode_n),
				.pld_scan_shift_n(in_pld_scan_shift_n),
				
				// UNUSED
				.int_pldif_8g_ltr(),
				.int_pldif_avmm_pld_avmm1_request(),
				.int_pldif_avmm_pld_avmm2_request(),
				.int_pldif_avmm_refclk_dig_en(),
				.int_pldif_g3_scan_mode_n(),
				.pld_8g_eidleinfersel_fifo(),
				.pld_8g_eidleinfersel_reg(),
				.pld_partial_reconfig_fifo(),
				.pld_partial_reconfig_rx_div_by_2_rxclk_wire(),
				.pld_partial_reconfig_rx_div_by_2_txclk_wire(),
				.pld_partial_reconfig_rxclk_reg(),
				.pld_partial_reconfig_tx_div_by_2_wire(),
				.pld_partial_reconfig_txclk_reg(),
				.pld_rate_reg(),
				.pld_test_data_reg()
			);
		end // if generate
		else begin
				assign w_hssi_common_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_clk[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_npor = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_usermode = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2 = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_adapt_done = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_clklow = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_fref = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_hclk = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_found = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_testbus[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_reserved_out[9:0] = 10'b0;
				assign w_hssi_common_pld_pcs_interface_pld_test_data[19:0] = 20'b0;
				assign w_hssi_common_pld_pcs_interface_pld_uhsif_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_scan_mode_n = 1'b1;		// Override default tieoff
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_rx_pcs
			twentynm_hssi_fifo_rx_pcs #(
				.double_read_mode(hssi_fifo_rx_pcs_double_read_mode),
				.prot_mode(hssi_fifo_rx_pcs_prot_mode),
				.silicon_rev( "20nm2" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_rx_pcs_blockselect),
				.data_out2_10g(w_hssi_fifo_rx_pcs_data_out2_10g),
				.data_out2_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp),
				.data_out_10g(w_hssi_fifo_rx_pcs_data_out_10g),
				.data_out_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out_8g_clock_comp),
				.data_out_8g_phase_comp(w_hssi_fifo_rx_pcs_data_out_8g_phase_comp),
				.data_out_gen3(w_hssi_fifo_rx_pcs_data_out_gen3),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_data[73], w_hssi_10g_rx_pcs_rx_fifo_wr_data[72], w_hssi_10g_rx_pcs_rx_fifo_wr_data[71], w_hssi_10g_rx_pcs_rx_fifo_wr_data[70], w_hssi_10g_rx_pcs_rx_fifo_wr_data[69], w_hssi_10g_rx_pcs_rx_fifo_wr_data[68], w_hssi_10g_rx_pcs_rx_fifo_wr_data[67], w_hssi_10g_rx_pcs_rx_fifo_wr_data[66], w_hssi_10g_rx_pcs_rx_fifo_wr_data[65], w_hssi_10g_rx_pcs_rx_fifo_wr_data[64], w_hssi_10g_rx_pcs_rx_fifo_wr_data[63], w_hssi_10g_rx_pcs_rx_fifo_wr_data[62], w_hssi_10g_rx_pcs_rx_fifo_wr_data[61], w_hssi_10g_rx_pcs_rx_fifo_wr_data[60], w_hssi_10g_rx_pcs_rx_fifo_wr_data[59], w_hssi_10g_rx_pcs_rx_fifo_wr_data[58], w_hssi_10g_rx_pcs_rx_fifo_wr_data[57], w_hssi_10g_rx_pcs_rx_fifo_wr_data[56], w_hssi_10g_rx_pcs_rx_fifo_wr_data[55], w_hssi_10g_rx_pcs_rx_fifo_wr_data[54], w_hssi_10g_rx_pcs_rx_fifo_wr_data[53], w_hssi_10g_rx_pcs_rx_fifo_wr_data[52], w_hssi_10g_rx_pcs_rx_fifo_wr_data[51], w_hssi_10g_rx_pcs_rx_fifo_wr_data[50], w_hssi_10g_rx_pcs_rx_fifo_wr_data[49], w_hssi_10g_rx_pcs_rx_fifo_wr_data[48], w_hssi_10g_rx_pcs_rx_fifo_wr_data[47], w_hssi_10g_rx_pcs_rx_fifo_wr_data[46], w_hssi_10g_rx_pcs_rx_fifo_wr_data[45], w_hssi_10g_rx_pcs_rx_fifo_wr_data[44], w_hssi_10g_rx_pcs_rx_fifo_wr_data[43], w_hssi_10g_rx_pcs_rx_fifo_wr_data[42], w_hssi_10g_rx_pcs_rx_fifo_wr_data[41], w_hssi_10g_rx_pcs_rx_fifo_wr_data[40], w_hssi_10g_rx_pcs_rx_fifo_wr_data[39], w_hssi_10g_rx_pcs_rx_fifo_wr_data[38], w_hssi_10g_rx_pcs_rx_fifo_wr_data[37], w_hssi_10g_rx_pcs_rx_fifo_wr_data[36], w_hssi_10g_rx_pcs_rx_fifo_wr_data[35], w_hssi_10g_rx_pcs_rx_fifo_wr_data[34], w_hssi_10g_rx_pcs_rx_fifo_wr_data[33], w_hssi_10g_rx_pcs_rx_fifo_wr_data[32], w_hssi_10g_rx_pcs_rx_fifo_wr_data[31], w_hssi_10g_rx_pcs_rx_fifo_wr_data[30], w_hssi_10g_rx_pcs_rx_fifo_wr_data[29], w_hssi_10g_rx_pcs_rx_fifo_wr_data[28], w_hssi_10g_rx_pcs_rx_fifo_wr_data[27], w_hssi_10g_rx_pcs_rx_fifo_wr_data[26], w_hssi_10g_rx_pcs_rx_fifo_wr_data[25], w_hssi_10g_rx_pcs_rx_fifo_wr_data[24], w_hssi_10g_rx_pcs_rx_fifo_wr_data[23], w_hssi_10g_rx_pcs_rx_fifo_wr_data[22], w_hssi_10g_rx_pcs_rx_fifo_wr_data[21], w_hssi_10g_rx_pcs_rx_fifo_wr_data[20], w_hssi_10g_rx_pcs_rx_fifo_wr_data[19], w_hssi_10g_rx_pcs_rx_fifo_wr_data[18], w_hssi_10g_rx_pcs_rx_fifo_wr_data[17], w_hssi_10g_rx_pcs_rx_fifo_wr_data[16], w_hssi_10g_rx_pcs_rx_fifo_wr_data[15], w_hssi_10g_rx_pcs_rx_fifo_wr_data[14], w_hssi_10g_rx_pcs_rx_fifo_wr_data[13], w_hssi_10g_rx_pcs_rx_fifo_wr_data[12], w_hssi_10g_rx_pcs_rx_fifo_wr_data[11], w_hssi_10g_rx_pcs_rx_fifo_wr_data[10], w_hssi_10g_rx_pcs_rx_fifo_wr_data[9], w_hssi_10g_rx_pcs_rx_fifo_wr_data[8], w_hssi_10g_rx_pcs_rx_fifo_wr_data[7], w_hssi_10g_rx_pcs_rx_fifo_wr_data[6], w_hssi_10g_rx_pcs_rx_fifo_wr_data[5], w_hssi_10g_rx_pcs_rx_fifo_wr_data[4], w_hssi_10g_rx_pcs_rx_fifo_wr_data[3], w_hssi_10g_rx_pcs_rx_fifo_wr_data[2], w_hssi_10g_rx_pcs_rx_fifo_wr_data[1], w_hssi_10g_rx_pcs_rx_fifo_wr_data[0]}),
				.data_in_8g_clock_comp({w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0]}),
				.data_in_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr2_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0]}),
				.rd_ptr2_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0]}),
				.rd_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0]}),
				.rd_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.wr_clk_8g_clock_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_8g_clock_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.wr_en_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.wr_en_8g_clock_comp(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_en_8g_phase_comp(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.wr_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0]}),
				.wr_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0]}),
				.wr_rst_n_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.wr_rst_n_8g_clock_comp(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_n_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_rx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79:0] = 80'b0;
				assign w_hssi_fifo_rx_pcs_data_out_gen3[39:0] = 40'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_tx_pcs
			twentynm_hssi_fifo_tx_pcs #(
				.double_write_mode(hssi_fifo_tx_pcs_double_write_mode),
				.prot_mode(hssi_fifo_tx_pcs_prot_mode),
				.silicon_rev( "20nm2" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_tx_pcs_blockselect),
				.data_out_10g(w_hssi_fifo_tx_pcs_data_out_10g),
				.data_out_8g_phase_comp(w_hssi_fifo_tx_pcs_data_out_8g_phase_comp),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in2_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0]}),
				.data_in_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_en_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.wr_en_8g_phase_comp(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0]}),
				.wr_rst_n_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_tx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_tx_pcs_data_out_10g[72:0] = 73'b0;
				assign w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63:0] = 64'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_rx_pcs
			twentynm_hssi_gen3_rx_pcs #(
				.block_sync(hssi_gen3_rx_pcs_block_sync),
				.block_sync_sm(hssi_gen3_rx_pcs_block_sync_sm),
				.cdr_ctrl_force_unalgn(hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn),
				.lpbk_force(hssi_gen3_rx_pcs_lpbk_force),
				.mode(hssi_gen3_rx_pcs_mode),
				.rate_match_fifo(hssi_gen3_rx_pcs_rate_match_fifo),
				.rate_match_fifo_latency(hssi_gen3_rx_pcs_rate_match_fifo_latency),
				.reconfig_settings(hssi_gen3_rx_pcs_reconfig_settings),
				.reverse_lpbk(hssi_gen3_rx_pcs_reverse_lpbk),
				.rx_b4gb_par_lpbk(hssi_gen3_rx_pcs_rx_b4gb_par_lpbk),
				.rx_force_balign(hssi_gen3_rx_pcs_rx_force_balign),
				.rx_ins_del_one_skip(hssi_gen3_rx_pcs_rx_ins_del_one_skip),
				.rx_num_fixed_pat(hssi_gen3_rx_pcs_rx_num_fixed_pat),
				.rx_test_out_sel(hssi_gen3_rx_pcs_rx_test_out_sel),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_rx_pcs_sup_mode)
			) inst_twentynm_hssi_gen3_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_rx_pcs_avmmreaddata),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.blk_start(w_hssi_gen3_rx_pcs_blk_start),
				.blockselect(w_hssi_gen3_rx_pcs_blockselect),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.data_out(w_hssi_gen3_rx_pcs_data_out),
				.data_valid(w_hssi_gen3_rx_pcs_data_valid),
				.ei_det_int(w_hssi_gen3_rx_pcs_ei_det_int),
				.ei_partial_det_int(w_hssi_gen3_rx_pcs_ei_partial_det_int),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.i_det_int(w_hssi_gen3_rx_pcs_i_det_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data(w_hssi_gen3_rx_pcs_lpbk_data),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.mem_rx_fifo_rd_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr),
				.mem_rx_fifo_wr_clk(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.mem_rx_fifo_wr_data(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data),
				.mem_rx_fifo_wr_en(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.mem_rx_fifo_wr_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr),
				.mem_rx_fifo_wr_rst_n(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_test_out(w_hssi_gen3_rx_pcs_rx_test_out),
				.sync_hdr(w_hssi_gen3_rx_pcs_sync_hdr),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0]}),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.mem_rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_gen3[39], w_hssi_fifo_rx_pcs_data_out_gen3[38], w_hssi_fifo_rx_pcs_data_out_gen3[37], w_hssi_fifo_rx_pcs_data_out_gen3[36], w_hssi_fifo_rx_pcs_data_out_gen3[35], w_hssi_fifo_rx_pcs_data_out_gen3[34], w_hssi_fifo_rx_pcs_data_out_gen3[33], w_hssi_fifo_rx_pcs_data_out_gen3[32], w_hssi_fifo_rx_pcs_data_out_gen3[31], w_hssi_fifo_rx_pcs_data_out_gen3[30], w_hssi_fifo_rx_pcs_data_out_gen3[29], w_hssi_fifo_rx_pcs_data_out_gen3[28], w_hssi_fifo_rx_pcs_data_out_gen3[27], w_hssi_fifo_rx_pcs_data_out_gen3[26], w_hssi_fifo_rx_pcs_data_out_gen3[25], w_hssi_fifo_rx_pcs_data_out_gen3[24], w_hssi_fifo_rx_pcs_data_out_gen3[23], w_hssi_fifo_rx_pcs_data_out_gen3[22], w_hssi_fifo_rx_pcs_data_out_gen3[21], w_hssi_fifo_rx_pcs_data_out_gen3[20], w_hssi_fifo_rx_pcs_data_out_gen3[19], w_hssi_fifo_rx_pcs_data_out_gen3[18], w_hssi_fifo_rx_pcs_data_out_gen3[17], w_hssi_fifo_rx_pcs_data_out_gen3[16], w_hssi_fifo_rx_pcs_data_out_gen3[15], w_hssi_fifo_rx_pcs_data_out_gen3[14], w_hssi_fifo_rx_pcs_data_out_gen3[13], w_hssi_fifo_rx_pcs_data_out_gen3[12], w_hssi_fifo_rx_pcs_data_out_gen3[11], w_hssi_fifo_rx_pcs_data_out_gen3[10], w_hssi_fifo_rx_pcs_data_out_gen3[9], w_hssi_fifo_rx_pcs_data_out_gen3[8], w_hssi_fifo_rx_pcs_data_out_gen3[7], w_hssi_fifo_rx_pcs_data_out_gen3[6], w_hssi_fifo_rx_pcs_data_out_gen3[5], w_hssi_fifo_rx_pcs_data_out_gen3[4], w_hssi_fifo_rx_pcs_data_out_gen3[3], w_hssi_fifo_rx_pcs_data_out_gen3[2], w_hssi_fifo_rx_pcs_data_out_gen3[1], w_hssi_fifo_rx_pcs_data_out_gen3[0]}),
				.par_lpbk_b4gb_in({w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0]}),
				.par_lpbk_in({w_hssi_gen3_tx_pcs_par_lpbk_out[31], w_hssi_gen3_tx_pcs_par_lpbk_out[30], w_hssi_gen3_tx_pcs_par_lpbk_out[29], w_hssi_gen3_tx_pcs_par_lpbk_out[28], w_hssi_gen3_tx_pcs_par_lpbk_out[27], w_hssi_gen3_tx_pcs_par_lpbk_out[26], w_hssi_gen3_tx_pcs_par_lpbk_out[25], w_hssi_gen3_tx_pcs_par_lpbk_out[24], w_hssi_gen3_tx_pcs_par_lpbk_out[23], w_hssi_gen3_tx_pcs_par_lpbk_out[22], w_hssi_gen3_tx_pcs_par_lpbk_out[21], w_hssi_gen3_tx_pcs_par_lpbk_out[20], w_hssi_gen3_tx_pcs_par_lpbk_out[19], w_hssi_gen3_tx_pcs_par_lpbk_out[18], w_hssi_gen3_tx_pcs_par_lpbk_out[17], w_hssi_gen3_tx_pcs_par_lpbk_out[16], w_hssi_gen3_tx_pcs_par_lpbk_out[15], w_hssi_gen3_tx_pcs_par_lpbk_out[14], w_hssi_gen3_tx_pcs_par_lpbk_out[13], w_hssi_gen3_tx_pcs_par_lpbk_out[12], w_hssi_gen3_tx_pcs_par_lpbk_out[11], w_hssi_gen3_tx_pcs_par_lpbk_out[10], w_hssi_gen3_tx_pcs_par_lpbk_out[9], w_hssi_gen3_tx_pcs_par_lpbk_out[8], w_hssi_gen3_tx_pcs_par_lpbk_out[7], w_hssi_gen3_tx_pcs_par_lpbk_out[6], w_hssi_gen3_tx_pcs_par_lpbk_out[5], w_hssi_gen3_tx_pcs_par_lpbk_out[4], w_hssi_gen3_tx_pcs_par_lpbk_out[3], w_hssi_gen3_tx_pcs_par_lpbk_out[2], w_hssi_gen3_tx_pcs_par_lpbk_out[1], w_hssi_gen3_tx_pcs_par_lpbk_out[0]}),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.rcvd_clk(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_pma_clk(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.rxpolarity(w_hssi_pipe_gen3_rxpolarity_int),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.sync_sm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.txdatak_in({w_hssi_pipe_gen3_txdatak_int[3], w_hssi_pipe_gen3_txdatak_int[2], w_hssi_pipe_gen3_txdatak_int[1], w_hssi_pipe_gen3_txdatak_int[0]}),
				
				// UNUSED
				.blk_lockd_int(),
				.skp_det_int()
			);
		end // if generate
		else begin
				assign w_hssi_gen3_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_rx_pcs_blk_algnd_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_delete_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_insert_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_overfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_undfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_rx_pcs_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_partial_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_err_decode_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_i_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data[33:0] = 34'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39:0] = 40'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_rx_test_out[19:0] = 20'b0;
				assign w_hssi_gen3_rx_pcs_sync_hdr[1:0] = 2'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_tx_pcs
			twentynm_hssi_gen3_tx_pcs #(
				.mode(hssi_gen3_tx_pcs_mode),
				.reverse_lpbk(hssi_gen3_tx_pcs_reverse_lpbk),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_tx_pcs_sup_mode),
				.tx_bitslip(hssi_gen3_tx_pcs_tx_bitslip),
				.tx_gbox_byp(hssi_gen3_tx_pcs_tx_gbox_byp)
			) inst_twentynm_hssi_gen3_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_gen3_tx_pcs_blockselect),
				.data_out(w_hssi_gen3_tx_pcs_data_out),
				.par_lpbk_b4gb_out(w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out),
				.par_lpbk_out(w_hssi_gen3_tx_pcs_par_lpbk_out),
				.tx_test_out(w_hssi_gen3_tx_pcs_tx_test_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_start_in(w_hssi_pipe_gen3_tx_blk_start_int),
				.data_in({w_hssi_pipe_gen3_txdata_int[31], w_hssi_pipe_gen3_txdata_int[30], w_hssi_pipe_gen3_txdata_int[29], w_hssi_pipe_gen3_txdata_int[28], w_hssi_pipe_gen3_txdata_int[27], w_hssi_pipe_gen3_txdata_int[26], w_hssi_pipe_gen3_txdata_int[25], w_hssi_pipe_gen3_txdata_int[24], w_hssi_pipe_gen3_txdata_int[23], w_hssi_pipe_gen3_txdata_int[22], w_hssi_pipe_gen3_txdata_int[21], w_hssi_pipe_gen3_txdata_int[20], w_hssi_pipe_gen3_txdata_int[19], w_hssi_pipe_gen3_txdata_int[18], w_hssi_pipe_gen3_txdata_int[17], w_hssi_pipe_gen3_txdata_int[16], w_hssi_pipe_gen3_txdata_int[15], w_hssi_pipe_gen3_txdata_int[14], w_hssi_pipe_gen3_txdata_int[13], w_hssi_pipe_gen3_txdata_int[12], w_hssi_pipe_gen3_txdata_int[11], w_hssi_pipe_gen3_txdata_int[10], w_hssi_pipe_gen3_txdata_int[9], w_hssi_pipe_gen3_txdata_int[8], w_hssi_pipe_gen3_txdata_int[7], w_hssi_pipe_gen3_txdata_int[6], w_hssi_pipe_gen3_txdata_int[5], w_hssi_pipe_gen3_txdata_int[4], w_hssi_pipe_gen3_txdata_int[3], w_hssi_pipe_gen3_txdata_int[2], w_hssi_pipe_gen3_txdata_int[1], w_hssi_pipe_gen3_txdata_int[0]}),
				.data_valid(w_hssi_pipe_gen3_txdataskip_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data_in({w_hssi_gen3_rx_pcs_lpbk_data[33], w_hssi_gen3_rx_pcs_lpbk_data[32], w_hssi_gen3_rx_pcs_lpbk_data[31], w_hssi_gen3_rx_pcs_lpbk_data[30], w_hssi_gen3_rx_pcs_lpbk_data[29], w_hssi_gen3_rx_pcs_lpbk_data[28], w_hssi_gen3_rx_pcs_lpbk_data[27], w_hssi_gen3_rx_pcs_lpbk_data[26], w_hssi_gen3_rx_pcs_lpbk_data[25], w_hssi_gen3_rx_pcs_lpbk_data[24], w_hssi_gen3_rx_pcs_lpbk_data[23], w_hssi_gen3_rx_pcs_lpbk_data[22], w_hssi_gen3_rx_pcs_lpbk_data[21], w_hssi_gen3_rx_pcs_lpbk_data[20], w_hssi_gen3_rx_pcs_lpbk_data[19], w_hssi_gen3_rx_pcs_lpbk_data[18], w_hssi_gen3_rx_pcs_lpbk_data[17], w_hssi_gen3_rx_pcs_lpbk_data[16], w_hssi_gen3_rx_pcs_lpbk_data[15], w_hssi_gen3_rx_pcs_lpbk_data[14], w_hssi_gen3_rx_pcs_lpbk_data[13], w_hssi_gen3_rx_pcs_lpbk_data[12], w_hssi_gen3_rx_pcs_lpbk_data[11], w_hssi_gen3_rx_pcs_lpbk_data[10], w_hssi_gen3_rx_pcs_lpbk_data[9], w_hssi_gen3_rx_pcs_lpbk_data[8], w_hssi_gen3_rx_pcs_lpbk_data[7], w_hssi_gen3_rx_pcs_lpbk_data[6], w_hssi_gen3_rx_pcs_lpbk_data[5], w_hssi_gen3_rx_pcs_lpbk_data[4], w_hssi_gen3_rx_pcs_lpbk_data[3], w_hssi_gen3_rx_pcs_lpbk_data[2], w_hssi_gen3_rx_pcs_lpbk_data[1], w_hssi_gen3_rx_pcs_lpbk_data[0]}),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.sync_in({w_hssi_pipe_gen3_tx_sync_hdr_int[1], w_hssi_pipe_gen3_tx_sync_hdr_int[0]}),
				.tx_pma_clk(w_hssi_8g_tx_pcs_clk_out_gen3),
				.tx_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn)
			);
		end // if generate
		else begin
				assign w_hssi_gen3_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_tx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_tx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35:0] = 36'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_tx_test_out[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_rx_pcs
			twentynm_hssi_krfec_rx_pcs #(
				.blksync_cor_en(hssi_krfec_rx_pcs_blksync_cor_en),
				.bypass_gb(hssi_krfec_rx_pcs_bypass_gb),
				.clr_ctrl(hssi_krfec_rx_pcs_clr_ctrl),
				.ctrl_bit_reverse(hssi_krfec_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_rx_pcs_data_bit_reverse),
				.dv_start(hssi_krfec_rx_pcs_dv_start),
				.err_mark_type(hssi_krfec_rx_pcs_err_mark_type),
				.error_marking_en(hssi_krfec_rx_pcs_error_marking_en),
				.low_latency_en(hssi_krfec_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_krfec_rx_pcs_lpbk_mode),
				.parity_invalid_enum(hssi_krfec_rx_pcs_parity_invalid_enum),
				.parity_valid_num(hssi_krfec_rx_pcs_parity_valid_num),
				.pipeln_blksync(hssi_krfec_rx_pcs_pipeln_blksync),
				.pipeln_descrm(hssi_krfec_rx_pcs_pipeln_descrm),
				.pipeln_errcorrect(hssi_krfec_rx_pcs_pipeln_errcorrect),
				.pipeln_errtrap_ind(hssi_krfec_rx_pcs_pipeln_errtrap_ind),
				.pipeln_errtrap_lfsr(hssi_krfec_rx_pcs_pipeln_errtrap_lfsr),
				.pipeln_errtrap_loc(hssi_krfec_rx_pcs_pipeln_errtrap_loc),
				.pipeln_errtrap_pat(hssi_krfec_rx_pcs_pipeln_errtrap_pat),
				.pipeln_gearbox(hssi_krfec_rx_pcs_pipeln_gearbox),
				.pipeln_syndrm(hssi_krfec_rx_pcs_pipeln_syndrm),
				.pipeln_trans_dec(hssi_krfec_rx_pcs_pipeln_trans_dec),
				.prot_mode(hssi_krfec_rx_pcs_prot_mode),
				.receive_order(hssi_krfec_rx_pcs_receive_order),
				.reconfig_settings(hssi_krfec_rx_pcs_reconfig_settings),
				.rx_testbus_sel(hssi_krfec_rx_pcs_rx_testbus_sel),
				.signal_ok_en(hssi_krfec_rx_pcs_signal_ok_en),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_rx_pcs_sup_mode)
			) inst_twentynm_hssi_krfec_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_rx_pcs_blockselect),
				.rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.rx_control_out(w_hssi_krfec_rx_pcs_rx_control_out),
				.rx_data_out(w_hssi_krfec_rx_pcs_rx_data_out),
				.rx_data_status(w_hssi_krfec_rx_pcs_rx_data_status),
				.rx_data_valid_out(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.rx_signal_ok_out(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.rx_data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0]}),
				.rx_krfec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_krfec_reg(),
				.pld_10g_krfec_rx_blk_lock_krfec_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg(),
				.pld_10g_krfec_rx_frame_krfec_reg(),
				.pld_10g_krfec_rx_frame_krfec_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_rx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_block_lock = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_control_out[9:0] = 10'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_status[1:0] = 2'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_valid_out = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_frame = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_signal_ok_out = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_tx_pcs
			twentynm_hssi_krfec_tx_pcs #(
				.burst_err(hssi_krfec_tx_pcs_burst_err),
				.burst_err_len(hssi_krfec_tx_pcs_burst_err_len),
				.ctrl_bit_reverse(hssi_krfec_tx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_tx_pcs_data_bit_reverse),
				.enc_frame_query(hssi_krfec_tx_pcs_enc_frame_query),
				.low_latency_en(hssi_krfec_tx_pcs_low_latency_en),
				.pipeln_encoder(hssi_krfec_tx_pcs_pipeln_encoder),
				.pipeln_scrambler(hssi_krfec_tx_pcs_pipeln_scrambler),
				.prot_mode(hssi_krfec_tx_pcs_prot_mode),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_tx_pcs_sup_mode),
				.transcode_err(hssi_krfec_tx_pcs_transcode_err),
				.transmit_order(hssi_krfec_tx_pcs_transmit_order),
				.tx_testbus_sel(hssi_krfec_tx_pcs_tx_testbus_sel)
			) inst_twentynm_hssi_krfec_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_tx_pcs_blockselect),
				.tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.tx_data_out(w_hssi_krfec_tx_pcs_tx_data_out),
				.tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.tx_test_data(w_hssi_krfec_tx_pcs_tx_test_data),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.tx_control_in({w_hssi_10g_tx_pcs_tx_control_out_krfec[8], w_hssi_10g_tx_pcs_tx_control_out_krfec[7], w_hssi_10g_tx_pcs_tx_control_out_krfec[6], w_hssi_10g_tx_pcs_tx_control_out_krfec[5], w_hssi_10g_tx_pcs_tx_control_out_krfec[4], w_hssi_10g_tx_pcs_tx_control_out_krfec[3], w_hssi_10g_tx_pcs_tx_control_out_krfec[2], w_hssi_10g_tx_pcs_tx_control_out_krfec[1], w_hssi_10g_tx_pcs_tx_control_out_krfec[0]}),
				.tx_data_in({w_hssi_10g_tx_pcs_tx_data_out_krfec[63], w_hssi_10g_tx_pcs_tx_data_out_krfec[62], w_hssi_10g_tx_pcs_tx_data_out_krfec[61], w_hssi_10g_tx_pcs_tx_data_out_krfec[60], w_hssi_10g_tx_pcs_tx_data_out_krfec[59], w_hssi_10g_tx_pcs_tx_data_out_krfec[58], w_hssi_10g_tx_pcs_tx_data_out_krfec[57], w_hssi_10g_tx_pcs_tx_data_out_krfec[56], w_hssi_10g_tx_pcs_tx_data_out_krfec[55], w_hssi_10g_tx_pcs_tx_data_out_krfec[54], w_hssi_10g_tx_pcs_tx_data_out_krfec[53], w_hssi_10g_tx_pcs_tx_data_out_krfec[52], w_hssi_10g_tx_pcs_tx_data_out_krfec[51], w_hssi_10g_tx_pcs_tx_data_out_krfec[50], w_hssi_10g_tx_pcs_tx_data_out_krfec[49], w_hssi_10g_tx_pcs_tx_data_out_krfec[48], w_hssi_10g_tx_pcs_tx_data_out_krfec[47], w_hssi_10g_tx_pcs_tx_data_out_krfec[46], w_hssi_10g_tx_pcs_tx_data_out_krfec[45], w_hssi_10g_tx_pcs_tx_data_out_krfec[44], w_hssi_10g_tx_pcs_tx_data_out_krfec[43], w_hssi_10g_tx_pcs_tx_data_out_krfec[42], w_hssi_10g_tx_pcs_tx_data_out_krfec[41], w_hssi_10g_tx_pcs_tx_data_out_krfec[40], w_hssi_10g_tx_pcs_tx_data_out_krfec[39], w_hssi_10g_tx_pcs_tx_data_out_krfec[38], w_hssi_10g_tx_pcs_tx_data_out_krfec[37], w_hssi_10g_tx_pcs_tx_data_out_krfec[36], w_hssi_10g_tx_pcs_tx_data_out_krfec[35], w_hssi_10g_tx_pcs_tx_data_out_krfec[34], w_hssi_10g_tx_pcs_tx_data_out_krfec[33], w_hssi_10g_tx_pcs_tx_data_out_krfec[32], w_hssi_10g_tx_pcs_tx_data_out_krfec[31], w_hssi_10g_tx_pcs_tx_data_out_krfec[30], w_hssi_10g_tx_pcs_tx_data_out_krfec[29], w_hssi_10g_tx_pcs_tx_data_out_krfec[28], w_hssi_10g_tx_pcs_tx_data_out_krfec[27], w_hssi_10g_tx_pcs_tx_data_out_krfec[26], w_hssi_10g_tx_pcs_tx_data_out_krfec[25], w_hssi_10g_tx_pcs_tx_data_out_krfec[24], w_hssi_10g_tx_pcs_tx_data_out_krfec[23], w_hssi_10g_tx_pcs_tx_data_out_krfec[22], w_hssi_10g_tx_pcs_tx_data_out_krfec[21], w_hssi_10g_tx_pcs_tx_data_out_krfec[20], w_hssi_10g_tx_pcs_tx_data_out_krfec[19], w_hssi_10g_tx_pcs_tx_data_out_krfec[18], w_hssi_10g_tx_pcs_tx_data_out_krfec[17], w_hssi_10g_tx_pcs_tx_data_out_krfec[16], w_hssi_10g_tx_pcs_tx_data_out_krfec[15], w_hssi_10g_tx_pcs_tx_data_out_krfec[14], w_hssi_10g_tx_pcs_tx_data_out_krfec[13], w_hssi_10g_tx_pcs_tx_data_out_krfec[12], w_hssi_10g_tx_pcs_tx_data_out_krfec[11], w_hssi_10g_tx_pcs_tx_data_out_krfec[10], w_hssi_10g_tx_pcs_tx_data_out_krfec[9], w_hssi_10g_tx_pcs_tx_data_out_krfec[8], w_hssi_10g_tx_pcs_tx_data_out_krfec[7], w_hssi_10g_tx_pcs_tx_data_out_krfec[6], w_hssi_10g_tx_pcs_tx_data_out_krfec[5], w_hssi_10g_tx_pcs_tx_data_out_krfec[4], w_hssi_10g_tx_pcs_tx_data_out_krfec[3], w_hssi_10g_tx_pcs_tx_data_out_krfec[2], w_hssi_10g_tx_pcs_tx_data_out_krfec[1], w_hssi_10g_tx_pcs_tx_data_out_krfec[0]}),
				.tx_data_valid_in(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_krfec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_krfec_reg(),
				.pld_krfec_tx_alignment_plddirect_reg(),
				.pld_krfec_tx_alignment_reg()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_tx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_alignment = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_test_data[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen1_2
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen1_2
			twentynm_hssi_pipe_gen1_2 #(
				.elec_idle_delay_val(hssi_pipe_gen1_2_elec_idle_delay_val),
				.error_replace_pad(hssi_pipe_gen1_2_error_replace_pad),
				.hip_mode(hssi_pipe_gen1_2_hip_mode),
				.ind_error_reporting(hssi_pipe_gen1_2_ind_error_reporting),
				.phystatus_delay_val(hssi_pipe_gen1_2_phystatus_delay_val),
				.phystatus_rst_toggle(hssi_pipe_gen1_2_phystatus_rst_toggle),
				.pipe_byte_de_serializer_en(hssi_pipe_gen1_2_pipe_byte_de_serializer_en),
				.prot_mode(hssi_pipe_gen1_2_prot_mode),
				.reconfig_settings(hssi_pipe_gen1_2_reconfig_settings),
				.rx_pipe_enable(hssi_pipe_gen1_2_rx_pipe_enable),
				.rxdetect_bypass(hssi_pipe_gen1_2_rxdetect_bypass),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen1_2_sup_mode),
				.tx_pipe_enable(hssi_pipe_gen1_2_tx_pipe_enable),
				.txswing(hssi_pipe_gen1_2_txswing)
			) inst_twentynm_hssi_pipe_gen1_2 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen1_2_avmmreaddata),
				.blockselect(w_hssi_pipe_gen1_2_blockselect),
				.current_coeff(w_hssi_pipe_gen1_2_current_coeff),
				.phystatus(w_hssi_pipe_gen1_2_phystatus),
				.polarity_inversion_rx(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rev_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.rxelectricalidle_out(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxstatus(w_hssi_pipe_gen1_2_rxstatus),
				.rxvalid(w_hssi_pipe_gen1_2_rxvalid),
				.tx_elec_idle_out(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pipe_rx_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.power_state_transition_done_ena(1'b0),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rev_loopbk_pcs_gen3(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.revloopback(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.rx_pipe_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rxd({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxelectricalidle(w_hssi_8g_rx_pcs_eidle_detected),
				.rxelectricalidle_pcs_gen3(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.rxpolarity_pcs_gen3(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.tx_elec_idle_comp(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.txd_ch({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswingport(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.pld_8g_rxpolarity_pipe3_reg(),
				.rxd_ch(),
				.txd()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen1_2_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen1_2_blockselect = 1'b0;
				assign w_hssi_pipe_gen1_2_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen1_2_phystatus = 1'b0;
				assign w_hssi_pipe_gen1_2_polarity_inversion_rx = 1'b0;
				assign w_hssi_pipe_gen1_2_rev_loopbk = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelectricalidle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen1_2_rxvalid = 1'b0;
				assign w_hssi_pipe_gen1_2_tx_elec_idle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_txdetectrx = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen3
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen3
			twentynm_hssi_pipe_gen3 #(
				.bypass_rx_detection_enable(hssi_pipe_gen3_bypass_rx_detection_enable),
				.bypass_rx_preset(hssi_pipe_gen3_bypass_rx_preset),
				.bypass_rx_preset_enable(hssi_pipe_gen3_bypass_rx_preset_enable),
				.bypass_tx_coefficent(hssi_pipe_gen3_bypass_tx_coefficent),
				.bypass_tx_coefficent_enable(hssi_pipe_gen3_bypass_tx_coefficent_enable),
				.elecidle_delay_g3(hssi_pipe_gen3_elecidle_delay_g3),
				.ind_error_reporting(hssi_pipe_gen3_ind_error_reporting),
				.mode(hssi_pipe_gen3_mode),
				.phy_status_delay_g12(hssi_pipe_gen3_phy_status_delay_g12),
				.phy_status_delay_g3(hssi_pipe_gen3_phy_status_delay_g3),
				.phystatus_rst_toggle_g12(hssi_pipe_gen3_phystatus_rst_toggle_g12),
				.phystatus_rst_toggle_g3(hssi_pipe_gen3_phystatus_rst_toggle_g3),
				.rate_match_pad_insertion(hssi_pipe_gen3_rate_match_pad_insertion),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen3_sup_mode),
				.test_out_sel(hssi_pipe_gen3_test_out_sel)
			) inst_twentynm_hssi_pipe_gen3 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen3_avmmreaddata),
				.blockselect(w_hssi_pipe_gen3_blockselect),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.phystatus(w_hssi_pipe_gen3_phystatus),
				.pma_current_coeff(w_hssi_pipe_gen3_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_pipe_gen3_pma_current_rxpreset),
				.pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.rev_lpbk_8gpcs_out(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.rev_lpbk_int(w_hssi_pipe_gen3_rev_lpbk_int),
				.rx_blk_start(w_hssi_pipe_gen3_rx_blk_start),
				.rx_sync_hdr(w_hssi_pipe_gen3_rx_sync_hdr),
				.rxd_8gpcs_out(w_hssi_pipe_gen3_rxd_8gpcs_out),
				.rxdataskip(w_hssi_pipe_gen3_rxdataskip),
				.rxelecidle(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity_8gpcs_out(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.rxpolarity_int(w_hssi_pipe_gen3_rxpolarity_int),
				.rxstatus(w_hssi_pipe_gen3_rxstatus),
				.rxvalid(w_hssi_pipe_gen3_rxvalid),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.test_out(w_hssi_pipe_gen3_test_out),
				.tx_blk_start_int(w_hssi_pipe_gen3_tx_blk_start_int),
				.tx_sync_hdr_int(w_hssi_pipe_gen3_tx_sync_hdr_int),
				.txdata_int(w_hssi_pipe_gen3_txdata_int),
				.txdatak_int(w_hssi_pipe_gen3_txdatak_int),
				.txdataskip_int(w_hssi_pipe_gen3_txdataskip_int),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.current_coeff({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0]}),
				.current_rxpreset({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0]}),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.pcs_asn_bundling_in({w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0]}),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pipe_tx_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_blk_start_int(w_hssi_gen3_rx_pcs_blk_start),
				.rx_sync_hdr_int({w_hssi_gen3_rx_pcs_sync_hdr[1], w_hssi_gen3_rx_pcs_sync_hdr[0]}),
				.rx_test_out({w_hssi_gen3_rx_pcs_rx_test_out[19], w_hssi_gen3_rx_pcs_rx_test_out[18], w_hssi_gen3_rx_pcs_rx_test_out[17], w_hssi_gen3_rx_pcs_rx_test_out[16], w_hssi_gen3_rx_pcs_rx_test_out[15], w_hssi_gen3_rx_pcs_rx_test_out[14], w_hssi_gen3_rx_pcs_rx_test_out[13], w_hssi_gen3_rx_pcs_rx_test_out[12], w_hssi_gen3_rx_pcs_rx_test_out[11], w_hssi_gen3_rx_pcs_rx_test_out[10], w_hssi_gen3_rx_pcs_rx_test_out[9], w_hssi_gen3_rx_pcs_rx_test_out[8], w_hssi_gen3_rx_pcs_rx_test_out[7], w_hssi_gen3_rx_pcs_rx_test_out[6], w_hssi_gen3_rx_pcs_rx_test_out[5], w_hssi_gen3_rx_pcs_rx_test_out[4], w_hssi_gen3_rx_pcs_rx_test_out[3], w_hssi_gen3_rx_pcs_rx_test_out[2], w_hssi_gen3_rx_pcs_rx_test_out[1], w_hssi_gen3_rx_pcs_rx_test_out[0]}),
				.rxd_8gpcs_in({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxdata_int({w_hssi_gen3_rx_pcs_data_out[31], w_hssi_gen3_rx_pcs_data_out[30], w_hssi_gen3_rx_pcs_data_out[29], w_hssi_gen3_rx_pcs_data_out[28], w_hssi_gen3_rx_pcs_data_out[27], w_hssi_gen3_rx_pcs_data_out[26], w_hssi_gen3_rx_pcs_data_out[25], w_hssi_gen3_rx_pcs_data_out[24], w_hssi_gen3_rx_pcs_data_out[23], w_hssi_gen3_rx_pcs_data_out[22], w_hssi_gen3_rx_pcs_data_out[21], w_hssi_gen3_rx_pcs_data_out[20], w_hssi_gen3_rx_pcs_data_out[19], w_hssi_gen3_rx_pcs_data_out[18], w_hssi_gen3_rx_pcs_data_out[17], w_hssi_gen3_rx_pcs_data_out[16], w_hssi_gen3_rx_pcs_data_out[15], w_hssi_gen3_rx_pcs_data_out[14], w_hssi_gen3_rx_pcs_data_out[13], w_hssi_gen3_rx_pcs_data_out[12], w_hssi_gen3_rx_pcs_data_out[11], w_hssi_gen3_rx_pcs_data_out[10], w_hssi_gen3_rx_pcs_data_out[9], w_hssi_gen3_rx_pcs_data_out[8], w_hssi_gen3_rx_pcs_data_out[7], w_hssi_gen3_rx_pcs_data_out[6], w_hssi_gen3_rx_pcs_data_out[5], w_hssi_gen3_rx_pcs_data_out[4], w_hssi_gen3_rx_pcs_data_out[3], w_hssi_gen3_rx_pcs_data_out[2], w_hssi_gen3_rx_pcs_data_out[1], w_hssi_gen3_rx_pcs_data_out[0]}),
				.rxdatak_int({1'b0, 1'b0, 1'b0, 1'b0}),
				.rxdataskip_int(w_hssi_gen3_rx_pcs_data_valid),
				.rxelecidle_8gpcs_in(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.tx_blk_start(w_hssi_8g_tx_pcs_tx_blk_start_out[0]),
				.tx_sync_hdr({w_hssi_8g_tx_pcs_tx_sync_hdr_out[1], w_hssi_8g_tx_pcs_tx_sync_hdr_out[0]}),
				.tx_test_out({w_hssi_gen3_tx_pcs_tx_test_out[19], w_hssi_gen3_tx_pcs_tx_test_out[18], w_hssi_gen3_tx_pcs_tx_test_out[17], w_hssi_gen3_tx_pcs_tx_test_out[16], w_hssi_gen3_tx_pcs_tx_test_out[15], w_hssi_gen3_tx_pcs_tx_test_out[14], w_hssi_gen3_tx_pcs_tx_test_out[13], w_hssi_gen3_tx_pcs_tx_test_out[12], w_hssi_gen3_tx_pcs_tx_test_out[11], w_hssi_gen3_tx_pcs_tx_test_out[10], w_hssi_gen3_tx_pcs_tx_test_out[9], w_hssi_gen3_tx_pcs_tx_test_out[8], w_hssi_gen3_tx_pcs_tx_test_out[7], w_hssi_gen3_tx_pcs_tx_test_out[6], w_hssi_gen3_tx_pcs_tx_test_out[5], w_hssi_gen3_tx_pcs_tx_test_out[4], w_hssi_gen3_tx_pcs_tx_test_out[3], w_hssi_gen3_tx_pcs_tx_test_out[2], w_hssi_gen3_tx_pcs_tx_test_out[1], w_hssi_gen3_tx_pcs_tx_test_out[0]}),
				.txcompliance(w_hssi_8g_tx_pcs_txcompliance_out),
				.txdata({w_hssi_8g_tx_pcs_tx_data_out[31], w_hssi_8g_tx_pcs_tx_data_out[30], w_hssi_8g_tx_pcs_tx_data_out[29], w_hssi_8g_tx_pcs_tx_data_out[28], w_hssi_8g_tx_pcs_tx_data_out[27], w_hssi_8g_tx_pcs_tx_data_out[26], w_hssi_8g_tx_pcs_tx_data_out[25], w_hssi_8g_tx_pcs_tx_data_out[24], w_hssi_8g_tx_pcs_tx_data_out[23], w_hssi_8g_tx_pcs_tx_data_out[22], w_hssi_8g_tx_pcs_tx_data_out[21], w_hssi_8g_tx_pcs_tx_data_out[20], w_hssi_8g_tx_pcs_tx_data_out[19], w_hssi_8g_tx_pcs_tx_data_out[18], w_hssi_8g_tx_pcs_tx_data_out[17], w_hssi_8g_tx_pcs_tx_data_out[16], w_hssi_8g_tx_pcs_tx_data_out[15], w_hssi_8g_tx_pcs_tx_data_out[14], w_hssi_8g_tx_pcs_tx_data_out[13], w_hssi_8g_tx_pcs_tx_data_out[12], w_hssi_8g_tx_pcs_tx_data_out[11], w_hssi_8g_tx_pcs_tx_data_out[10], w_hssi_8g_tx_pcs_tx_data_out[9], w_hssi_8g_tx_pcs_tx_data_out[8], w_hssi_8g_tx_pcs_tx_data_out[7], w_hssi_8g_tx_pcs_tx_data_out[6], w_hssi_8g_tx_pcs_tx_data_out[5], w_hssi_8g_tx_pcs_tx_data_out[4], w_hssi_8g_tx_pcs_tx_data_out[3], w_hssi_8g_tx_pcs_tx_data_out[2], w_hssi_8g_tx_pcs_tx_data_out[1], w_hssi_8g_tx_pcs_tx_data_out[0]}),
				.txdatak({w_hssi_8g_tx_pcs_tx_datak_out[3], w_hssi_8g_tx_pcs_tx_datak_out[2], w_hssi_8g_tx_pcs_tx_datak_out[1], w_hssi_8g_tx_pcs_tx_datak_out[0]}),
				.txdataskip(w_hssi_8g_tx_pcs_tx_data_valid_out[0]),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_8g_tx_pcs_txelecidle_out),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.dis_pc_byte(),
				.pma_rx_det_pd(),
				.pma_txdeemph(),
				.pma_txmargin(),
				.pma_txswing(),
				.reset_pc_prts()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen3_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen3_blockselect = 1'b0;
				assign w_hssi_pipe_gen3_gen3_clk_sel = 1'b0;
				assign w_hssi_pipe_gen3_pcs_rst = 1'b0;
				assign w_hssi_pipe_gen3_phystatus = 1'b0;
				assign w_hssi_pipe_gen3_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen3_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_pma_tx_elec_idle = 1'b0;
				assign w_hssi_pipe_gen3_pma_txdetectrx = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_int = 1'b0;
				assign w_hssi_pipe_gen3_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_rxd_8gpcs_out[63:0] = 64'b0;
				assign w_hssi_pipe_gen3_rxdataskip[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_int = 1'b0;
				assign w_hssi_pipe_gen3_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_rxvalid = 1'b0;
				assign w_hssi_pipe_gen3_shutdown_clk = 1'b0;
				assign w_hssi_pipe_gen3_test_out[19:0] = 20'b0;
				assign w_hssi_pipe_gen3_tx_blk_start_int = 1'b0;
				assign w_hssi_pipe_gen3_tx_sync_hdr_int[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_txdata_int[31:0] = 32'b0;
				assign w_hssi_pipe_gen3_txdatak_int[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_txdataskip_int = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pcs_pma_interface
			twentynm_hssi_rx_pcs_pma_interface #(
				.block_sel(hssi_rx_pcs_pma_interface_block_sel),
				.channel_operation_mode(hssi_rx_pcs_pma_interface_channel_operation_mode),
				.clkslip_sel(hssi_rx_pcs_pma_interface_clkslip_sel),
				.lpbk_en(hssi_rx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_rx_pcs_pma_interface_master_clk_sel),
				.pldif_datawidth_mode(hssi_rx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_rx(hssi_rx_pcs_pma_interface_pma_dw_rx),
				.pma_if_dft_en(hssi_rx_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_rx_pcs_pma_interface_pma_if_dft_val),
				.prbs9_dwidth(hssi_rx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_rx_pcs_pma_interface_prbs_clken),
				.prbs_ver(hssi_rx_pcs_pma_interface_prbs_ver),
				.prot_mode_rx(hssi_rx_pcs_pma_interface_prot_mode_rx),
				.reconfig_settings(hssi_rx_pcs_pma_interface_reconfig_settings),
				.rx_dyn_polarity_inversion(hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion),
				.rx_lpbk_en(hssi_rx_pcs_pma_interface_rx_lpbk_en),
				.rx_prbs_force_signal_ok(hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok),
				.rx_prbs_mask(hssi_rx_pcs_pma_interface_rx_prbs_mask),
				.rx_prbs_mode(hssi_rx_pcs_pma_interface_rx_prbs_mode),
				.rx_signalok_signaldet_sel(hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel),
				.rx_static_polarity_inversion(hssi_rx_pcs_pma_interface_rx_static_polarity_inversion),
				.rx_uhsif_lpbk_en(hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sup_mode(hssi_rx_pcs_pma_interface_sup_mode)
			) inst_twentynm_hssi_rx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.int_pmaif_10g_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data),
				.int_pmaif_10g_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.int_pmaif_8g_pudi(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi),
				.int_pmaif_8g_rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.int_pmaif_8g_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.int_pmaif_8g_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.int_pmaif_8g_sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.int_pmaif_g3_pma_data_in(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in),
				.int_pmaif_g3_pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.int_pmaif_g3_pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.int_pmaif_g3_pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.int_pmaif_krfec_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data),
				.int_pmaif_krfec_rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.int_pmaif_pldif_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pmaif_pldif_prbs_err_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pmaif_pldif_rx_clkdiv(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pmaif_pldif_rx_clkdiv_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pmaif_pldif_rx_data(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data),
				.int_pmaif_pldif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pmaif_pldif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pmaif_pldif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pmaif_pldif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.pma_eye_monitor(w_hssi_rx_pcs_pma_interface_pma_eye_monitor),
				.pma_rx_clkslip(w_hssi_rx_pcs_pma_interface_pma_rx_clkslip),
				.pma_rxpma_rstb(w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb),
				.rx_pmaif_test_out(w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out),
				.rx_prbs_ver_test(w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.int_pmaif_8g_rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.int_pmaif_pldif_eye_monitor({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0]}),
				.int_pmaif_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pmaif_pldif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pmaif_pldif_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pmaif_pldif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pma_rx_clkdiv_user(in_pma_rx_clkdiv_user),
				.pma_rx_detect_valid(in_pma_rx_detect_valid),
				.pma_rx_found(in_pma_rx_found),
				.pma_rx_pma_clk(in_pma_rx_pma_clk),
				.pma_rx_pma_data({in_pma_rx_pma_data[63], in_pma_rx_pma_data[62], in_pma_rx_pma_data[61], in_pma_rx_pma_data[60], in_pma_rx_pma_data[59], in_pma_rx_pma_data[58], in_pma_rx_pma_data[57], in_pma_rx_pma_data[56], in_pma_rx_pma_data[55], in_pma_rx_pma_data[54], in_pma_rx_pma_data[53], in_pma_rx_pma_data[52], in_pma_rx_pma_data[51], in_pma_rx_pma_data[50], in_pma_rx_pma_data[49], in_pma_rx_pma_data[48], in_pma_rx_pma_data[47], in_pma_rx_pma_data[46], in_pma_rx_pma_data[45], in_pma_rx_pma_data[44], in_pma_rx_pma_data[43], in_pma_rx_pma_data[42], in_pma_rx_pma_data[41], in_pma_rx_pma_data[40], in_pma_rx_pma_data[39], in_pma_rx_pma_data[38], in_pma_rx_pma_data[37], in_pma_rx_pma_data[36], in_pma_rx_pma_data[35], in_pma_rx_pma_data[34], in_pma_rx_pma_data[33], in_pma_rx_pma_data[32], in_pma_rx_pma_data[31], in_pma_rx_pma_data[30], in_pma_rx_pma_data[29], in_pma_rx_pma_data[28], in_pma_rx_pma_data[27], in_pma_rx_pma_data[26], in_pma_rx_pma_data[25], in_pma_rx_pma_data[24], in_pma_rx_pma_data[23], in_pma_rx_pma_data[22], in_pma_rx_pma_data[21], in_pma_rx_pma_data[20], in_pma_rx_pma_data[19], in_pma_rx_pma_data[18], in_pma_rx_pma_data[17], in_pma_rx_pma_data[16], in_pma_rx_pma_data[15], in_pma_rx_pma_data[14], in_pma_rx_pma_data[13], in_pma_rx_pma_data[12], in_pma_rx_pma_data[11], in_pma_rx_pma_data[10], in_pma_rx_pma_data[9], in_pma_rx_pma_data[8], in_pma_rx_pma_data[7], in_pma_rx_pma_data[6], in_pma_rx_pma_data[5], in_pma_rx_pma_data[4], in_pma_rx_pma_data[3], in_pma_rx_pma_data[2], in_pma_rx_pma_data[1], in_pma_rx_pma_data[0]}),
				.pma_rx_signal_ok(in_pma_rx_signal_ok),
				.pma_rxpll_lock(in_pma_rxpll_lock),
				.pma_signal_det(in_pma_signal_det),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.tx_pma_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0]}),
				.tx_pma_uhsif_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0]}),
				
				// UNUSED
				.int_pmaif_g3_rcvd_clk(),
				.prbs_err_lt()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31:0] = 32'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5:0] = 6'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rx_clkslip = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pld_pcs_interface
			twentynm_hssi_rx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx),
				.hd_10g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx),
				.hd_10g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx),
				.hd_10g_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx),
				.hd_10g_lpbk_en(hssi_rx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx),
				.hd_10g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx),
				.hd_10g_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx),
				.hd_10g_test_bus_mode(hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode),
				.hd_8g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx),
				.hd_8g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx),
				.hd_8g_hip_mode(hssi_rx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_rx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx),
				.hd_8g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx),
				.hd_chnl_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_clklow_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz),
				.hd_chnl_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx),
				.hd_chnl_fref_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz),
				.hd_chnl_frequency_rules_en(hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_rx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_rx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx),
				.hd_chnl_lpbk_en(hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx),
				.hd_chnl_pld_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz),
				.hd_chnl_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx),
				.hd_chnl_pma_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz),
				.hd_chnl_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx),
				.hd_chnl_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx),
				.hd_chnl_transparent_pcs_rx(hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx),
				.hd_fifo_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx),
				.hd_fifo_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx),
				.hd_g3_prot_mode(hssi_rx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx),
				.hd_krfec_lpbk_en(hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx),
				.hd_krfec_test_bus_mode(hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode),
				.hd_pldif_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx),
				.hd_pmaif_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_lpbk_en(hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx),
				.hd_pmaif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx),
				.hd_pmaif_sim_mode(hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_rx_block_sel(hssi_rx_pld_pcs_interface_pcs_rx_block_sel),
				.pcs_rx_clk_out_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel),
				.pcs_rx_clk_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_sel),
				.pcs_rx_hip_clk_en(hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en),
				.pcs_rx_output_sel(hssi_rx_pld_pcs_interface_pcs_rx_output_sel),
				.reconfig_settings(hssi_rx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm2" )       //PARAM_HIDE
			) inst_twentynm_hssi_rx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pld_pcs_interface_blockselect),
				.hip_rx_ctrl(w_hssi_rx_pld_pcs_interface_hip_rx_ctrl),
				.hip_rx_data(w_hssi_rx_pld_pcs_interface_hip_rx_data),
				.int_pldif_10g_rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.int_pldif_10g_rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.int_pldif_10g_rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.int_pldif_10g_rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.int_pldif_10g_rx_control_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb),
				.int_pldif_10g_rx_data_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb),
				.int_pldif_10g_rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.int_pldif_10g_rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.int_pldif_10g_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.int_pldif_10g_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.int_pldif_10g_rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.int_pldif_8g_a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.int_pldif_8g_bitloc_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.int_pldif_8g_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.int_pldif_8g_byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.int_pldif_8g_encdt(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.int_pldif_8g_pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.int_pldif_8g_rdenable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.int_pldif_8g_rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.int_pldif_8g_rxurstpcs_n(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.int_pldif_8g_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.int_pldif_8g_wrdisable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.int_pldif_g3_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.int_pldif_krfec_rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.int_pldif_pmaif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pldif_pmaif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pldif_pmaif_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pldif_pmaif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pld_10g_krfec_rx_blk_lock(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock),
				.pld_10g_krfec_rx_diag_data_status(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status),
				.pld_10g_krfec_rx_frame(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame),
				.pld_10g_rx_align_val(w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val),
				.pld_10g_rx_crc32_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err),
				.pld_10g_rx_data_valid(w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid),
				.pld_10g_rx_empty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty),
				.pld_10g_rx_fifo_del(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del),
				.pld_10g_rx_fifo_insert(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert),
				.pld_10g_rx_fifo_num(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num),
				.pld_10g_rx_frame_lock(w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock),
				.pld_10g_rx_hi_ber(w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber),
				.pld_10g_rx_oflw_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err),
				.pld_10g_rx_pempty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty),
				.pld_10g_rx_pfull(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull),
				.pld_8g_a1a2_k1k2_flag(w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag),
				.pld_8g_empty_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf),
				.pld_8g_empty_rx(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx),
				.pld_8g_full_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf),
				.pld_8g_full_rx(w_hssi_rx_pld_pcs_interface_pld_8g_full_rx),
				.pld_8g_rxelecidle(w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle),
				.pld_8g_signal_detect_out(w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out),
				.pld_8g_wa_boundary(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary),
				.pld_pcs_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out),
				.pld_pma_clkdiv_rx_user(w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user),
				.pld_pma_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out),
				.pld_pma_signal_ok(w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok),
				.pld_rx_control(w_hssi_rx_pld_pcs_interface_pld_rx_control),
				.pld_rx_data(w_hssi_rx_pld_pcs_interface_pld_rx_data),
				.pld_rx_prbs_done(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done),
				.pld_rx_prbs_err(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.int_pldif_10g_rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.int_pldif_10g_rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.int_pldif_10g_rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_10g_rx_control({w_hssi_10g_rx_pcs_rx_control[19], w_hssi_10g_rx_pcs_rx_control[18], w_hssi_10g_rx_pcs_rx_control[17], w_hssi_10g_rx_pcs_rx_control[16], w_hssi_10g_rx_pcs_rx_control[15], w_hssi_10g_rx_pcs_rx_control[14], w_hssi_10g_rx_pcs_rx_control[13], w_hssi_10g_rx_pcs_rx_control[12], w_hssi_10g_rx_pcs_rx_control[11], w_hssi_10g_rx_pcs_rx_control[10], w_hssi_10g_rx_pcs_rx_control[9], w_hssi_10g_rx_pcs_rx_control[8], w_hssi_10g_rx_pcs_rx_control[7], w_hssi_10g_rx_pcs_rx_control[6], w_hssi_10g_rx_pcs_rx_control[5], w_hssi_10g_rx_pcs_rx_control[4], w_hssi_10g_rx_pcs_rx_control[3], w_hssi_10g_rx_pcs_rx_control[2], w_hssi_10g_rx_pcs_rx_control[1], w_hssi_10g_rx_pcs_rx_control[0]}),
				.int_pldif_10g_rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.int_pldif_10g_rx_data({w_hssi_10g_rx_pcs_rx_data[127], w_hssi_10g_rx_pcs_rx_data[126], w_hssi_10g_rx_pcs_rx_data[125], w_hssi_10g_rx_pcs_rx_data[124], w_hssi_10g_rx_pcs_rx_data[123], w_hssi_10g_rx_pcs_rx_data[122], w_hssi_10g_rx_pcs_rx_data[121], w_hssi_10g_rx_pcs_rx_data[120], w_hssi_10g_rx_pcs_rx_data[119], w_hssi_10g_rx_pcs_rx_data[118], w_hssi_10g_rx_pcs_rx_data[117], w_hssi_10g_rx_pcs_rx_data[116], w_hssi_10g_rx_pcs_rx_data[115], w_hssi_10g_rx_pcs_rx_data[114], w_hssi_10g_rx_pcs_rx_data[113], w_hssi_10g_rx_pcs_rx_data[112], w_hssi_10g_rx_pcs_rx_data[111], w_hssi_10g_rx_pcs_rx_data[110], w_hssi_10g_rx_pcs_rx_data[109], w_hssi_10g_rx_pcs_rx_data[108], w_hssi_10g_rx_pcs_rx_data[107], w_hssi_10g_rx_pcs_rx_data[106], w_hssi_10g_rx_pcs_rx_data[105], w_hssi_10g_rx_pcs_rx_data[104], w_hssi_10g_rx_pcs_rx_data[103], w_hssi_10g_rx_pcs_rx_data[102], w_hssi_10g_rx_pcs_rx_data[101], w_hssi_10g_rx_pcs_rx_data[100], w_hssi_10g_rx_pcs_rx_data[99], w_hssi_10g_rx_pcs_rx_data[98], w_hssi_10g_rx_pcs_rx_data[97], w_hssi_10g_rx_pcs_rx_data[96], w_hssi_10g_rx_pcs_rx_data[95], w_hssi_10g_rx_pcs_rx_data[94], w_hssi_10g_rx_pcs_rx_data[93], w_hssi_10g_rx_pcs_rx_data[92], w_hssi_10g_rx_pcs_rx_data[91], w_hssi_10g_rx_pcs_rx_data[90], w_hssi_10g_rx_pcs_rx_data[89], w_hssi_10g_rx_pcs_rx_data[88], w_hssi_10g_rx_pcs_rx_data[87], w_hssi_10g_rx_pcs_rx_data[86], w_hssi_10g_rx_pcs_rx_data[85], w_hssi_10g_rx_pcs_rx_data[84], w_hssi_10g_rx_pcs_rx_data[83], w_hssi_10g_rx_pcs_rx_data[82], w_hssi_10g_rx_pcs_rx_data[81], w_hssi_10g_rx_pcs_rx_data[80], w_hssi_10g_rx_pcs_rx_data[79], w_hssi_10g_rx_pcs_rx_data[78], w_hssi_10g_rx_pcs_rx_data[77], w_hssi_10g_rx_pcs_rx_data[76], w_hssi_10g_rx_pcs_rx_data[75], w_hssi_10g_rx_pcs_rx_data[74], w_hssi_10g_rx_pcs_rx_data[73], w_hssi_10g_rx_pcs_rx_data[72], w_hssi_10g_rx_pcs_rx_data[71], w_hssi_10g_rx_pcs_rx_data[70], w_hssi_10g_rx_pcs_rx_data[69], w_hssi_10g_rx_pcs_rx_data[68], w_hssi_10g_rx_pcs_rx_data[67], w_hssi_10g_rx_pcs_rx_data[66], w_hssi_10g_rx_pcs_rx_data[65], w_hssi_10g_rx_pcs_rx_data[64], w_hssi_10g_rx_pcs_rx_data[63], w_hssi_10g_rx_pcs_rx_data[62], w_hssi_10g_rx_pcs_rx_data[61], w_hssi_10g_rx_pcs_rx_data[60], w_hssi_10g_rx_pcs_rx_data[59], w_hssi_10g_rx_pcs_rx_data[58], w_hssi_10g_rx_pcs_rx_data[57], w_hssi_10g_rx_pcs_rx_data[56], w_hssi_10g_rx_pcs_rx_data[55], w_hssi_10g_rx_pcs_rx_data[54], w_hssi_10g_rx_pcs_rx_data[53], w_hssi_10g_rx_pcs_rx_data[52], w_hssi_10g_rx_pcs_rx_data[51], w_hssi_10g_rx_pcs_rx_data[50], w_hssi_10g_rx_pcs_rx_data[49], w_hssi_10g_rx_pcs_rx_data[48], w_hssi_10g_rx_pcs_rx_data[47], w_hssi_10g_rx_pcs_rx_data[46], w_hssi_10g_rx_pcs_rx_data[45], w_hssi_10g_rx_pcs_rx_data[44], w_hssi_10g_rx_pcs_rx_data[43], w_hssi_10g_rx_pcs_rx_data[42], w_hssi_10g_rx_pcs_rx_data[41], w_hssi_10g_rx_pcs_rx_data[40], w_hssi_10g_rx_pcs_rx_data[39], w_hssi_10g_rx_pcs_rx_data[38], w_hssi_10g_rx_pcs_rx_data[37], w_hssi_10g_rx_pcs_rx_data[36], w_hssi_10g_rx_pcs_rx_data[35], w_hssi_10g_rx_pcs_rx_data[34], w_hssi_10g_rx_pcs_rx_data[33], w_hssi_10g_rx_pcs_rx_data[32], w_hssi_10g_rx_pcs_rx_data[31], w_hssi_10g_rx_pcs_rx_data[30], w_hssi_10g_rx_pcs_rx_data[29], w_hssi_10g_rx_pcs_rx_data[28], w_hssi_10g_rx_pcs_rx_data[27], w_hssi_10g_rx_pcs_rx_data[26], w_hssi_10g_rx_pcs_rx_data[25], w_hssi_10g_rx_pcs_rx_data[24], w_hssi_10g_rx_pcs_rx_data[23], w_hssi_10g_rx_pcs_rx_data[22], w_hssi_10g_rx_pcs_rx_data[21], w_hssi_10g_rx_pcs_rx_data[20], w_hssi_10g_rx_pcs_rx_data[19], w_hssi_10g_rx_pcs_rx_data[18], w_hssi_10g_rx_pcs_rx_data[17], w_hssi_10g_rx_pcs_rx_data[16], w_hssi_10g_rx_pcs_rx_data[15], w_hssi_10g_rx_pcs_rx_data[14], w_hssi_10g_rx_pcs_rx_data[13], w_hssi_10g_rx_pcs_rx_data[12], w_hssi_10g_rx_pcs_rx_data[11], w_hssi_10g_rx_pcs_rx_data[10], w_hssi_10g_rx_pcs_rx_data[9], w_hssi_10g_rx_pcs_rx_data[8], w_hssi_10g_rx_pcs_rx_data[7], w_hssi_10g_rx_pcs_rx_data[6], w_hssi_10g_rx_pcs_rx_data[5], w_hssi_10g_rx_pcs_rx_data[4], w_hssi_10g_rx_pcs_rx_data[3], w_hssi_10g_rx_pcs_rx_data[2], w_hssi_10g_rx_pcs_rx_data[1], w_hssi_10g_rx_pcs_rx_data[0]}),
				.int_pldif_10g_rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.int_pldif_10g_rx_diag_status({w_hssi_10g_rx_pcs_rx_diag_status[1], w_hssi_10g_rx_pcs_rx_diag_status[0]}),
				.int_pldif_10g_rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.int_pldif_10g_rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.int_pldif_10g_rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.int_pldif_10g_rx_fifo_num({w_hssi_10g_rx_pcs_rx_fifo_num[4], w_hssi_10g_rx_pcs_rx_fifo_num[3], w_hssi_10g_rx_pcs_rx_fifo_num[2], w_hssi_10g_rx_pcs_rx_fifo_num[1], w_hssi_10g_rx_pcs_rx_fifo_num[0]}),
				.int_pldif_10g_rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.int_pldif_10g_rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.int_pldif_10g_rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.int_pldif_10g_rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.int_pldif_10g_rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.int_pldif_10g_rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				.int_pldif_8g_a1a2_k1k2_flag({w_hssi_8g_rx_pcs_a1a2k1k2flag[3], w_hssi_8g_rx_pcs_a1a2k1k2flag[2], w_hssi_8g_rx_pcs_a1a2k1k2flag[1], w_hssi_8g_rx_pcs_a1a2k1k2flag[0]}),
				.int_pldif_8g_empty_rmf(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.int_pldif_8g_empty_rx(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.int_pldif_8g_full_rmf(w_hssi_8g_rx_pcs_rm_fifo_full),
				.int_pldif_8g_full_rx(w_hssi_8g_rx_pcs_pcfifofull),
				.int_pldif_8g_phystatus(w_hssi_8g_rx_pcs_phystatus),
				.int_pldif_8g_rx_blk_start({w_hssi_8g_rx_pcs_rx_blk_start[3], w_hssi_8g_rx_pcs_rx_blk_start[2], w_hssi_8g_rx_pcs_rx_blk_start[1], w_hssi_8g_rx_pcs_rx_blk_start[0]}),
				.int_pldif_8g_rx_clk(w_hssi_8g_rx_pcs_clock_to_pld),
				.int_pldif_8g_rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_8g_rx_data_valid({w_hssi_8g_rx_pcs_rx_data_valid[3], w_hssi_8g_rx_pcs_rx_data_valid[2], w_hssi_8g_rx_pcs_rx_data_valid[1], w_hssi_8g_rx_pcs_rx_data_valid[0]}),
				.int_pldif_8g_rx_rstn_sync2wrfifo(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.int_pldif_8g_rx_sync_hdr({w_hssi_8g_rx_pcs_rx_sync_hdr[1], w_hssi_8g_rx_pcs_rx_sync_hdr[0]}),
				.int_pldif_8g_rxd({w_hssi_8g_rx_pcs_dataout[63], w_hssi_8g_rx_pcs_dataout[62], w_hssi_8g_rx_pcs_dataout[61], w_hssi_8g_rx_pcs_dataout[60], w_hssi_8g_rx_pcs_dataout[59], w_hssi_8g_rx_pcs_dataout[58], w_hssi_8g_rx_pcs_dataout[57], w_hssi_8g_rx_pcs_dataout[56], w_hssi_8g_rx_pcs_dataout[55], w_hssi_8g_rx_pcs_dataout[54], w_hssi_8g_rx_pcs_dataout[53], w_hssi_8g_rx_pcs_dataout[52], w_hssi_8g_rx_pcs_dataout[51], w_hssi_8g_rx_pcs_dataout[50], w_hssi_8g_rx_pcs_dataout[49], w_hssi_8g_rx_pcs_dataout[48], w_hssi_8g_rx_pcs_dataout[47], w_hssi_8g_rx_pcs_dataout[46], w_hssi_8g_rx_pcs_dataout[45], w_hssi_8g_rx_pcs_dataout[44], w_hssi_8g_rx_pcs_dataout[43], w_hssi_8g_rx_pcs_dataout[42], w_hssi_8g_rx_pcs_dataout[41], w_hssi_8g_rx_pcs_dataout[40], w_hssi_8g_rx_pcs_dataout[39], w_hssi_8g_rx_pcs_dataout[38], w_hssi_8g_rx_pcs_dataout[37], w_hssi_8g_rx_pcs_dataout[36], w_hssi_8g_rx_pcs_dataout[35], w_hssi_8g_rx_pcs_dataout[34], w_hssi_8g_rx_pcs_dataout[33], w_hssi_8g_rx_pcs_dataout[32], w_hssi_8g_rx_pcs_dataout[31], w_hssi_8g_rx_pcs_dataout[30], w_hssi_8g_rx_pcs_dataout[29], w_hssi_8g_rx_pcs_dataout[28], w_hssi_8g_rx_pcs_dataout[27], w_hssi_8g_rx_pcs_dataout[26], w_hssi_8g_rx_pcs_dataout[25], w_hssi_8g_rx_pcs_dataout[24], w_hssi_8g_rx_pcs_dataout[23], w_hssi_8g_rx_pcs_dataout[22], w_hssi_8g_rx_pcs_dataout[21], w_hssi_8g_rx_pcs_dataout[20], w_hssi_8g_rx_pcs_dataout[19], w_hssi_8g_rx_pcs_dataout[18], w_hssi_8g_rx_pcs_dataout[17], w_hssi_8g_rx_pcs_dataout[16], w_hssi_8g_rx_pcs_dataout[15], w_hssi_8g_rx_pcs_dataout[14], w_hssi_8g_rx_pcs_dataout[13], w_hssi_8g_rx_pcs_dataout[12], w_hssi_8g_rx_pcs_dataout[11], w_hssi_8g_rx_pcs_dataout[10], w_hssi_8g_rx_pcs_dataout[9], w_hssi_8g_rx_pcs_dataout[8], w_hssi_8g_rx_pcs_dataout[7], w_hssi_8g_rx_pcs_dataout[6], w_hssi_8g_rx_pcs_dataout[5], w_hssi_8g_rx_pcs_dataout[4], w_hssi_8g_rx_pcs_dataout[3], w_hssi_8g_rx_pcs_dataout[2], w_hssi_8g_rx_pcs_dataout[1], w_hssi_8g_rx_pcs_dataout[0]}),
				.int_pldif_8g_rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.int_pldif_8g_rxstatus({w_hssi_8g_rx_pcs_rxstatus[2], w_hssi_8g_rx_pcs_rxstatus[1], w_hssi_8g_rx_pcs_rxstatus[0]}),
				.int_pldif_8g_rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.int_pldif_8g_signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.int_pldif_8g_wa_boundary({w_hssi_8g_rx_pcs_word_align_boundary[4], w_hssi_8g_rx_pcs_word_align_boundary[3], w_hssi_8g_rx_pcs_word_align_boundary[2], w_hssi_8g_rx_pcs_word_align_boundary[1], w_hssi_8g_rx_pcs_word_align_boundary[0]}),
				.int_pldif_krfec_rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.int_pldif_krfec_rx_data_status({w_hssi_krfec_rx_pcs_rx_data_status[1], w_hssi_krfec_rx_pcs_rx_data_status[0]}),
				.int_pldif_krfec_rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.int_pldif_pmaif_clkdiv_rx(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pldif_pmaif_clkdiv_rx_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pldif_pmaif_rx_data({w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0]}),
				.int_pldif_pmaif_rx_prbs_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pldif_pmaif_rx_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.pld_10g_krfec_rx_clr_errblk_cnt(in_pld_10g_krfec_rx_clr_errblk_cnt),
				.pld_10g_krfec_rx_pld_rst_n(in_pld_10g_krfec_rx_pld_rst_n),
				.pld_10g_rx_align_clr(in_pld_10g_rx_align_clr),
				.pld_10g_rx_clr_ber_count(in_pld_10g_rx_clr_ber_count),
				.pld_10g_rx_rd_en(in_pld_10g_rx_rd_en),
				.pld_8g_a1a2_size(in_pld_8g_a1a2_size),
				.pld_8g_bitloc_rev_en(in_pld_8g_bitloc_rev_en),
				.pld_8g_byte_rev_en(in_pld_8g_byte_rev_en),
				.pld_8g_encdt(in_pld_8g_encdt),
				.pld_8g_g3_rx_pld_rst_n(in_pld_8g_g3_rx_pld_rst_n),
				.pld_8g_rdenable_rx(in_pld_8g_rdenable_rx),
				.pld_8g_rxpolarity(in_pld_8g_rxpolarity),
				.pld_8g_wrdisable_rx(in_pld_8g_wrdisable_rx),
				.pld_bitslip(in_pld_bitslip),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_rxpma_rstb(in_pld_pma_rxpma_rstb),
				.pld_pmaif_rx_pld_rst_n(in_pld_pmaif_rx_pld_rst_n),
				.pld_pmaif_rxclkslip(in_pld_pmaif_rxclkslip),
				.pld_polinv_rx(in_pld_polinv_rx),
				.pld_rx_clk(in_pld_rx_clk),
				.pld_rx_prbs_err_clr(in_pld_rx_prbs_err_clr),
				.pld_syncsm_en(in_pld_syncsm_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.int_pldif_pmaif_rx_pld_clk(),
				.pld_8g_wa_boundary_txclk_fastreg(),
				.pld_8g_wa_boundary_txclk_reg(),
				.pld_bitslip_10g_txclk_reg(),
				.pld_bitslip_8g_txclk_reg(),
				.pld_bitslip_rxclk_parallel_loopback_reg(),
				.pld_bitslip_rxclk_reg(),
				.pld_pcs_rx_clk_out_pcsdirect_wire(),
				.pld_pma_rx_clk_out_10g_or_pcsdirect_wire(),
				.pld_pma_rx_clk_out_8g_wire(),
				.pld_pmaif_rx_pld_rst_n_reg(),
				.pld_pmaif_tx_pld_rst_n_txclk_reg(),
				.pld_polinv_rx_reg(),
				.pld_rx_clk_fifo(),
				.pld_rx_control_fifo(),
				.pld_rx_control_pcsdirect_reg(),
				.pld_rx_data_fifo(),
				.pld_rx_data_pcsdirect_reg(),
				.pld_rx_prbs_done_reg(),
				.pld_rx_prbs_done_txclk_reg(),
				.pld_rx_prbs_err_clr_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_clr_reg(),
				.pld_rx_prbs_err_disprbs_reg(),
				.pld_rx_prbs_err_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_reg(),
				.pma_rx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_data[50:0] = 51'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3:0] = 4'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_control[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_data[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pcs_pma_interface
			twentynm_hssi_tx_pcs_pma_interface #(
				.bypass_pma_txelecidle(hssi_tx_pcs_pma_interface_bypass_pma_txelecidle),
				.channel_operation_mode(hssi_tx_pcs_pma_interface_channel_operation_mode),
				.lpbk_en(hssi_tx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_tx_pcs_pma_interface_master_clk_sel),
				.pcie_sub_prot_mode_tx(hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx),
				.pldif_datawidth_mode(hssi_tx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_tx(hssi_tx_pcs_pma_interface_pma_dw_tx),
				.pma_if_dft_en(hssi_tx_pcs_pma_interface_pma_if_dft_en),
				.pmagate_en(hssi_tx_pcs_pma_interface_pmagate_en),
				.prbs9_dwidth(hssi_tx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_tx_pcs_pma_interface_prbs_clken),
				.prbs_gen_pat(hssi_tx_pcs_pma_interface_prbs_gen_pat),
				.prot_mode_tx(hssi_tx_pcs_pma_interface_prot_mode_tx),
				.reconfig_settings(hssi_tx_pcs_pma_interface_reconfig_settings),
				.silicon_rev( "20nm2" ),       //PARAM_HIDE
				.sq_wave_num(hssi_tx_pcs_pma_interface_sq_wave_num),
				.sqwgen_clken(hssi_tx_pcs_pma_interface_sqwgen_clken),
				.sup_mode(hssi_tx_pcs_pma_interface_sup_mode),
				.tx_dyn_polarity_inversion(hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion),
				.tx_pma_data_sel(hssi_tx_pcs_pma_interface_tx_pma_data_sel),
				.tx_static_polarity_inversion(hssi_tx_pcs_pma_interface_tx_static_polarity_inversion),
				.uhsif_cnt_step_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock),
				.uhsif_cnt_thresh_filt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value),
				.uhsif_cnt_thresh_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock),
				.uhsif_dcn_test_update_period(hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period),
				.uhsif_dcn_testmode_enable(hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable),
				.uhsif_dead_zone_count_thresh(hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh),
				.uhsif_dead_zone_detection_enable(hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable),
				.uhsif_dead_zone_obser_window(hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window),
				.uhsif_dead_zone_skip_size(hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size),
				.uhsif_delay_cell_index_sel(hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel),
				.uhsif_delay_cell_margin(hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin),
				.uhsif_delay_cell_static_index_value(hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value),
				.uhsif_dft_dead_zone_control(hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control),
				.uhsif_dft_up_filt_control(hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control),
				.uhsif_enable(hssi_tx_pcs_pma_interface_uhsif_enable),
				.uhsif_lock_det_segsz_after_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock),
				.uhsif_lock_det_segsz_before_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock),
				.uhsif_lock_det_thresh_cnt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value),
				.uhsif_lock_det_thresh_cnt_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value),
				.uhsif_lock_det_thresh_diff_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value),
				.uhsif_lock_det_thresh_diff_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value)
			) inst_twentynm_hssi_tx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.int_pmaif_8g_txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.int_pmaif_pldif_tx_clkdiv(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pmaif_pldif_tx_clkdiv_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pmaif_pldif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.int_pmaif_pldif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.int_tx_dft_obsrv_clk(w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk),
				.pma_tx_elec_idle(w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle),
				.pma_tx_pma_data(w_hssi_tx_pcs_pma_interface_pma_tx_pma_data),
				.pma_txpma_rstb(w_hssi_tx_pcs_pma_interface_pma_txpma_rstb),
				.tx_pma_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback),
				.tx_pma_uhsif_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback),
				.tx_prbs_gen_test(w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test),
				.uhsif_test_out_1(w_hssi_tx_pcs_pma_interface_uhsif_test_out_1),
				.uhsif_test_out_2(w_hssi_tx_pcs_pma_interface_uhsif_test_out_2),
				.uhsif_test_out_3(w_hssi_tx_pcs_pma_interface_uhsif_test_out_3),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.int_pmaif_10g_tx_pma_data({w_hssi_10g_tx_pcs_tx_pma_data[63], w_hssi_10g_tx_pcs_tx_pma_data[62], w_hssi_10g_tx_pcs_tx_pma_data[61], w_hssi_10g_tx_pcs_tx_pma_data[60], w_hssi_10g_tx_pcs_tx_pma_data[59], w_hssi_10g_tx_pcs_tx_pma_data[58], w_hssi_10g_tx_pcs_tx_pma_data[57], w_hssi_10g_tx_pcs_tx_pma_data[56], w_hssi_10g_tx_pcs_tx_pma_data[55], w_hssi_10g_tx_pcs_tx_pma_data[54], w_hssi_10g_tx_pcs_tx_pma_data[53], w_hssi_10g_tx_pcs_tx_pma_data[52], w_hssi_10g_tx_pcs_tx_pma_data[51], w_hssi_10g_tx_pcs_tx_pma_data[50], w_hssi_10g_tx_pcs_tx_pma_data[49], w_hssi_10g_tx_pcs_tx_pma_data[48], w_hssi_10g_tx_pcs_tx_pma_data[47], w_hssi_10g_tx_pcs_tx_pma_data[46], w_hssi_10g_tx_pcs_tx_pma_data[45], w_hssi_10g_tx_pcs_tx_pma_data[44], w_hssi_10g_tx_pcs_tx_pma_data[43], w_hssi_10g_tx_pcs_tx_pma_data[42], w_hssi_10g_tx_pcs_tx_pma_data[41], w_hssi_10g_tx_pcs_tx_pma_data[40], w_hssi_10g_tx_pcs_tx_pma_data[39], w_hssi_10g_tx_pcs_tx_pma_data[38], w_hssi_10g_tx_pcs_tx_pma_data[37], w_hssi_10g_tx_pcs_tx_pma_data[36], w_hssi_10g_tx_pcs_tx_pma_data[35], w_hssi_10g_tx_pcs_tx_pma_data[34], w_hssi_10g_tx_pcs_tx_pma_data[33], w_hssi_10g_tx_pcs_tx_pma_data[32], w_hssi_10g_tx_pcs_tx_pma_data[31], w_hssi_10g_tx_pcs_tx_pma_data[30], w_hssi_10g_tx_pcs_tx_pma_data[29], w_hssi_10g_tx_pcs_tx_pma_data[28], w_hssi_10g_tx_pcs_tx_pma_data[27], w_hssi_10g_tx_pcs_tx_pma_data[26], w_hssi_10g_tx_pcs_tx_pma_data[25], w_hssi_10g_tx_pcs_tx_pma_data[24], w_hssi_10g_tx_pcs_tx_pma_data[23], w_hssi_10g_tx_pcs_tx_pma_data[22], w_hssi_10g_tx_pcs_tx_pma_data[21], w_hssi_10g_tx_pcs_tx_pma_data[20], w_hssi_10g_tx_pcs_tx_pma_data[19], w_hssi_10g_tx_pcs_tx_pma_data[18], w_hssi_10g_tx_pcs_tx_pma_data[17], w_hssi_10g_tx_pcs_tx_pma_data[16], w_hssi_10g_tx_pcs_tx_pma_data[15], w_hssi_10g_tx_pcs_tx_pma_data[14], w_hssi_10g_tx_pcs_tx_pma_data[13], w_hssi_10g_tx_pcs_tx_pma_data[12], w_hssi_10g_tx_pcs_tx_pma_data[11], w_hssi_10g_tx_pcs_tx_pma_data[10], w_hssi_10g_tx_pcs_tx_pma_data[9], w_hssi_10g_tx_pcs_tx_pma_data[8], w_hssi_10g_tx_pcs_tx_pma_data[7], w_hssi_10g_tx_pcs_tx_pma_data[6], w_hssi_10g_tx_pcs_tx_pma_data[5], w_hssi_10g_tx_pcs_tx_pma_data[4], w_hssi_10g_tx_pcs_tx_pma_data[3], w_hssi_10g_tx_pcs_tx_pma_data[2], w_hssi_10g_tx_pcs_tx_pma_data[1], w_hssi_10g_tx_pcs_tx_pma_data[0]}),
				.int_pmaif_10g_tx_pma_data_gate_val({w_hssi_10g_tx_pcs_tx_pma_gating_val[63], w_hssi_10g_tx_pcs_tx_pma_gating_val[62], w_hssi_10g_tx_pcs_tx_pma_gating_val[61], w_hssi_10g_tx_pcs_tx_pma_gating_val[60], w_hssi_10g_tx_pcs_tx_pma_gating_val[59], w_hssi_10g_tx_pcs_tx_pma_gating_val[58], w_hssi_10g_tx_pcs_tx_pma_gating_val[57], w_hssi_10g_tx_pcs_tx_pma_gating_val[56], w_hssi_10g_tx_pcs_tx_pma_gating_val[55], w_hssi_10g_tx_pcs_tx_pma_gating_val[54], w_hssi_10g_tx_pcs_tx_pma_gating_val[53], w_hssi_10g_tx_pcs_tx_pma_gating_val[52], w_hssi_10g_tx_pcs_tx_pma_gating_val[51], w_hssi_10g_tx_pcs_tx_pma_gating_val[50], w_hssi_10g_tx_pcs_tx_pma_gating_val[49], w_hssi_10g_tx_pcs_tx_pma_gating_val[48], w_hssi_10g_tx_pcs_tx_pma_gating_val[47], w_hssi_10g_tx_pcs_tx_pma_gating_val[46], w_hssi_10g_tx_pcs_tx_pma_gating_val[45], w_hssi_10g_tx_pcs_tx_pma_gating_val[44], w_hssi_10g_tx_pcs_tx_pma_gating_val[43], w_hssi_10g_tx_pcs_tx_pma_gating_val[42], w_hssi_10g_tx_pcs_tx_pma_gating_val[41], w_hssi_10g_tx_pcs_tx_pma_gating_val[40], w_hssi_10g_tx_pcs_tx_pma_gating_val[39], w_hssi_10g_tx_pcs_tx_pma_gating_val[38], w_hssi_10g_tx_pcs_tx_pma_gating_val[37], w_hssi_10g_tx_pcs_tx_pma_gating_val[36], w_hssi_10g_tx_pcs_tx_pma_gating_val[35], w_hssi_10g_tx_pcs_tx_pma_gating_val[34], w_hssi_10g_tx_pcs_tx_pma_gating_val[33], w_hssi_10g_tx_pcs_tx_pma_gating_val[32], w_hssi_10g_tx_pcs_tx_pma_gating_val[31], w_hssi_10g_tx_pcs_tx_pma_gating_val[30], w_hssi_10g_tx_pcs_tx_pma_gating_val[29], w_hssi_10g_tx_pcs_tx_pma_gating_val[28], w_hssi_10g_tx_pcs_tx_pma_gating_val[27], w_hssi_10g_tx_pcs_tx_pma_gating_val[26], w_hssi_10g_tx_pcs_tx_pma_gating_val[25], w_hssi_10g_tx_pcs_tx_pma_gating_val[24], w_hssi_10g_tx_pcs_tx_pma_gating_val[23], w_hssi_10g_tx_pcs_tx_pma_gating_val[22], w_hssi_10g_tx_pcs_tx_pma_gating_val[21], w_hssi_10g_tx_pcs_tx_pma_gating_val[20], w_hssi_10g_tx_pcs_tx_pma_gating_val[19], w_hssi_10g_tx_pcs_tx_pma_gating_val[18], w_hssi_10g_tx_pcs_tx_pma_gating_val[17], w_hssi_10g_tx_pcs_tx_pma_gating_val[16], w_hssi_10g_tx_pcs_tx_pma_gating_val[15], w_hssi_10g_tx_pcs_tx_pma_gating_val[14], w_hssi_10g_tx_pcs_tx_pma_gating_val[13], w_hssi_10g_tx_pcs_tx_pma_gating_val[12], w_hssi_10g_tx_pcs_tx_pma_gating_val[11], w_hssi_10g_tx_pcs_tx_pma_gating_val[10], w_hssi_10g_tx_pcs_tx_pma_gating_val[9], w_hssi_10g_tx_pcs_tx_pma_gating_val[8], w_hssi_10g_tx_pcs_tx_pma_gating_val[7], w_hssi_10g_tx_pcs_tx_pma_gating_val[6], w_hssi_10g_tx_pcs_tx_pma_gating_val[5], w_hssi_10g_tx_pcs_tx_pma_gating_val[4], w_hssi_10g_tx_pcs_tx_pma_gating_val[3], w_hssi_10g_tx_pcs_tx_pma_gating_val[2], w_hssi_10g_tx_pcs_tx_pma_gating_val[1], w_hssi_10g_tx_pcs_tx_pma_gating_val[0]}),
				.int_pmaif_8g_pudr({w_hssi_8g_tx_pcs_dataout[19], w_hssi_8g_tx_pcs_dataout[18], w_hssi_8g_tx_pcs_dataout[17], w_hssi_8g_tx_pcs_dataout[16], w_hssi_8g_tx_pcs_dataout[15], w_hssi_8g_tx_pcs_dataout[14], w_hssi_8g_tx_pcs_dataout[13], w_hssi_8g_tx_pcs_dataout[12], w_hssi_8g_tx_pcs_dataout[11], w_hssi_8g_tx_pcs_dataout[10], w_hssi_8g_tx_pcs_dataout[9], w_hssi_8g_tx_pcs_dataout[8], w_hssi_8g_tx_pcs_dataout[7], w_hssi_8g_tx_pcs_dataout[6], w_hssi_8g_tx_pcs_dataout[5], w_hssi_8g_tx_pcs_dataout[4], w_hssi_8g_tx_pcs_dataout[3], w_hssi_8g_tx_pcs_dataout[2], w_hssi_8g_tx_pcs_dataout[1], w_hssi_8g_tx_pcs_dataout[0]}),
				.int_pmaif_8g_tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.int_pmaif_8g_tx_elec_idle(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_pma_data_out({w_hssi_gen3_tx_pcs_data_out[31], w_hssi_gen3_tx_pcs_data_out[30], w_hssi_gen3_tx_pcs_data_out[29], w_hssi_gen3_tx_pcs_data_out[28], w_hssi_gen3_tx_pcs_data_out[27], w_hssi_gen3_tx_pcs_data_out[26], w_hssi_gen3_tx_pcs_data_out[25], w_hssi_gen3_tx_pcs_data_out[24], w_hssi_gen3_tx_pcs_data_out[23], w_hssi_gen3_tx_pcs_data_out[22], w_hssi_gen3_tx_pcs_data_out[21], w_hssi_gen3_tx_pcs_data_out[20], w_hssi_gen3_tx_pcs_data_out[19], w_hssi_gen3_tx_pcs_data_out[18], w_hssi_gen3_tx_pcs_data_out[17], w_hssi_gen3_tx_pcs_data_out[16], w_hssi_gen3_tx_pcs_data_out[15], w_hssi_gen3_tx_pcs_data_out[14], w_hssi_gen3_tx_pcs_data_out[13], w_hssi_gen3_tx_pcs_data_out[12], w_hssi_gen3_tx_pcs_data_out[11], w_hssi_gen3_tx_pcs_data_out[10], w_hssi_gen3_tx_pcs_data_out[9], w_hssi_gen3_tx_pcs_data_out[8], w_hssi_gen3_tx_pcs_data_out[7], w_hssi_gen3_tx_pcs_data_out[6], w_hssi_gen3_tx_pcs_data_out[5], w_hssi_gen3_tx_pcs_data_out[4], w_hssi_gen3_tx_pcs_data_out[3], w_hssi_gen3_tx_pcs_data_out[2], w_hssi_gen3_tx_pcs_data_out[1], w_hssi_gen3_tx_pcs_data_out[0]}),
				.int_pmaif_g3_pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.int_pmaif_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pmaif_pldif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pmaif_pldif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0]}),
				.int_pmaif_pldif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pmaif_pldif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.int_pmaif_pldif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pmaif_pldif_uhsif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0]}),
				.pma_tx_clkdiv_user(in_pma_tx_clkdiv_user),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.refclk_dig_uhsif(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.uhsif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.uhsif_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				
				// UNUSED
				.avmm_user_dataout(),
				.write_en(),
				.write_en_ack()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4:0] = 5'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_txpma_rstb = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pld_pcs_interface
			twentynm_hssi_tx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx),
				.hd_10g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx),
				.hd_10g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx),
				.hd_10g_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx),
				.hd_10g_lpbk_en(hssi_tx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx),
				.hd_10g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx),
				.hd_10g_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx),
				.hd_8g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx),
				.hd_8g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx),
				.hd_8g_hip_mode(hssi_tx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_tx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx),
				.hd_8g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx),
				.hd_chnl_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx),
				.hd_chnl_frequency_rules_en(hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_tx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_tx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx),
				.hd_chnl_lpbk_en(hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx),
				.hd_chnl_pld_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz),
				.hd_chnl_pld_uhsif_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz),
				.hd_chnl_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx),
				.hd_chnl_pma_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz),
				.hd_chnl_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx),
				.hd_chnl_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx),
				.hd_fifo_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx),
				.hd_fifo_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx),
				.hd_g3_prot_mode(hssi_tx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx),
				.hd_krfec_lpbk_en(hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx),
				.hd_pldif_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx),
				.hd_pmaif_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_ctrl_plane_bonding(hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding),
				.hd_pmaif_lpbk_en(hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx),
				.hd_pmaif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx),
				.hd_pmaif_sim_mode(hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_tx_clk_out_sel(hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel),
				.pcs_tx_clk_source(hssi_tx_pld_pcs_interface_pcs_tx_clk_source),
				.pcs_tx_data_source(hssi_tx_pld_pcs_interface_pcs_tx_data_source),
				.pcs_tx_delay1_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en),
				.pcs_tx_delay1_clk_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel),
				.pcs_tx_delay1_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl),
				.pcs_tx_delay1_data_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel),
				.pcs_tx_delay2_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en),
				.pcs_tx_delay2_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl),
				.pcs_tx_output_sel(hssi_tx_pld_pcs_interface_pcs_tx_output_sel),
				.reconfig_settings(hssi_tx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm2" )       //PARAM_HIDE
			) inst_twentynm_hssi_tx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pld_pcs_interface_blockselect),
				.hip_tx_clk(w_hssi_tx_pld_pcs_interface_hip_tx_clk),
				.int_pldif_10g_tx_bitslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip),
				.int_pldif_10g_tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.int_pldif_10g_tx_control(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control),
				.int_pldif_10g_tx_control_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg),
				.int_pldif_10g_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data),
				.int_pldif_10g_tx_data_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg),
				.int_pldif_10g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.int_pldif_10g_tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.int_pldif_10g_tx_diag_status(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status),
				.int_pldif_10g_tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.int_pldif_10g_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.int_pldif_10g_tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				.int_pldif_8g_pld_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.int_pldif_8g_powerdown(w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown),
				.int_pldif_8g_rddisable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.int_pldif_8g_rev_loopbk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.int_pldif_8g_tx_blk_start(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start),
				.int_pldif_8g_tx_boundary_sel(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel),
				.int_pldif_8g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid),
				.int_pldif_8g_tx_sync_hdr(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr),
				.int_pldif_8g_txd(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd),
				.int_pldif_8g_txd_fast_reg(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg),
				.int_pldif_8g_txdeemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.int_pldif_8g_txdetectrxloopback(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.int_pldif_8g_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.int_pldif_8g_txmargin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin),
				.int_pldif_8g_txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.int_pldif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.int_pldif_8g_wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				.int_pldif_pmaif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pldif_pmaif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pldif_pmaif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data),
				.int_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pldif_pmaif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pldif_pmaif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pldif_pmaif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pldif_pmaif_uhsif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data),
				.pld_10g_krfec_tx_frame(w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame),
				.pld_10g_tx_burst_en_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe),
				.pld_10g_tx_empty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty),
				.pld_10g_tx_fifo_num(w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num),
				.pld_10g_tx_full(w_hssi_tx_pld_pcs_interface_pld_10g_tx_full),
				.pld_10g_tx_pempty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty),
				.pld_10g_tx_pfull(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull),
				.pld_10g_tx_wordslip_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe),
				.pld_8g_empty_tx(w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx),
				.pld_8g_full_tx(w_hssi_tx_pld_pcs_interface_pld_8g_full_tx),
				.pld_krfec_tx_alignment(w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment),
				.pld_pcs_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out),
				.pld_pma_clkdiv_tx_user(w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user),
				.pld_pma_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out),
				.pld_uhsif_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.hip_tx_data({in_hip_tx_data[63], in_hip_tx_data[62], in_hip_tx_data[61], in_hip_tx_data[60], in_hip_tx_data[59], in_hip_tx_data[58], in_hip_tx_data[57], in_hip_tx_data[56], in_hip_tx_data[55], in_hip_tx_data[54], in_hip_tx_data[53], in_hip_tx_data[52], in_hip_tx_data[51], in_hip_tx_data[50], in_hip_tx_data[49], in_hip_tx_data[48], in_hip_tx_data[47], in_hip_tx_data[46], in_hip_tx_data[45], in_hip_tx_data[44], in_hip_tx_data[43], in_hip_tx_data[42], in_hip_tx_data[41], in_hip_tx_data[40], in_hip_tx_data[39], in_hip_tx_data[38], in_hip_tx_data[37], in_hip_tx_data[36], in_hip_tx_data[35], in_hip_tx_data[34], in_hip_tx_data[33], in_hip_tx_data[32], in_hip_tx_data[31], in_hip_tx_data[30], in_hip_tx_data[29], in_hip_tx_data[28], in_hip_tx_data[27], in_hip_tx_data[26], in_hip_tx_data[25], in_hip_tx_data[24], in_hip_tx_data[23], in_hip_tx_data[22], in_hip_tx_data[21], in_hip_tx_data[20], in_hip_tx_data[19], in_hip_tx_data[18], in_hip_tx_data[17], in_hip_tx_data[16], in_hip_tx_data[15], in_hip_tx_data[14], in_hip_tx_data[13], in_hip_tx_data[12], in_hip_tx_data[11], in_hip_tx_data[10], in_hip_tx_data[9], in_hip_tx_data[8], in_hip_tx_data[7], in_hip_tx_data[6], in_hip_tx_data[5], in_hip_tx_data[4], in_hip_tx_data[3], in_hip_tx_data[2], in_hip_tx_data[1], in_hip_tx_data[0]}),
				.int_pldif_10g_tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.int_pldif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.int_pldif_10g_tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_10g_tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.int_pldif_10g_tx_fifo_num({w_hssi_10g_tx_pcs_tx_fifo_num[3], w_hssi_10g_tx_pcs_tx_fifo_num[2], w_hssi_10g_tx_pcs_tx_fifo_num[1], w_hssi_10g_tx_pcs_tx_fifo_num[0]}),
				.int_pldif_10g_tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.int_pldif_10g_tx_full(w_hssi_10g_tx_pcs_tx_full),
				.int_pldif_10g_tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.int_pldif_10g_tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.int_pldif_10g_tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				.int_pldif_8g_empty_tx(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.int_pldif_8g_full_tx(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.int_pldif_8g_tx_clk_out(w_hssi_8g_tx_pcs_clk_out),
				.int_pldif_8g_tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_krfec_tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.int_pldif_krfec_tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.int_pldif_pmaif_clkdiv_tx(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pldif_pmaif_clkdiv_tx_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pldif_pmaif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.pld_10g_krfec_tx_pld_rst_n(in_pld_10g_krfec_tx_pld_rst_n),
				.pld_10g_tx_bitslip({in_pld_10g_tx_bitslip[6], in_pld_10g_tx_bitslip[5], in_pld_10g_tx_bitslip[4], in_pld_10g_tx_bitslip[3], in_pld_10g_tx_bitslip[2], in_pld_10g_tx_bitslip[1], in_pld_10g_tx_bitslip[0]}),
				.pld_10g_tx_burst_en(in_pld_10g_tx_burst_en),
				.pld_10g_tx_data_valid(in_pld_10g_tx_data_valid),
				.pld_10g_tx_diag_status({in_pld_10g_tx_diag_status[1], in_pld_10g_tx_diag_status[0]}),
				.pld_10g_tx_wordslip(in_pld_10g_tx_wordslip),
				.pld_8g_g3_tx_pld_rst_n(in_pld_8g_g3_tx_pld_rst_n),
				.pld_8g_rddisable_tx(in_pld_8g_rddisable_tx),
				.pld_8g_tx_boundary_sel({in_pld_8g_tx_boundary_sel[4], in_pld_8g_tx_boundary_sel[3], in_pld_8g_tx_boundary_sel[2], in_pld_8g_tx_boundary_sel[1], in_pld_8g_tx_boundary_sel[0]}),
				.pld_8g_wrenable_tx(in_pld_8g_wrenable_tx),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_txpma_rstb(in_pld_pma_txpma_rstb),
				.pld_pmaif_tx_pld_rst_n(in_pld_pmaif_tx_pld_rst_n),
				.pld_polinv_tx(in_pld_polinv_tx),
				.pld_tx_clk(in_pld_tx_clk),
				.pld_tx_control({in_pld_tx_control[17], in_pld_tx_control[16], in_pld_tx_control[15], in_pld_tx_control[14], in_pld_tx_control[13], in_pld_tx_control[12], in_pld_tx_control[11], in_pld_tx_control[10], in_pld_tx_control[9], in_pld_tx_control[8], in_pld_tx_control[7], in_pld_tx_control[6], in_pld_tx_control[5], in_pld_tx_control[4], in_pld_tx_control[3], in_pld_tx_control[2], in_pld_tx_control[1], in_pld_tx_control[0]}),
				.pld_tx_data({in_pld_tx_data[127], in_pld_tx_data[126], in_pld_tx_data[125], in_pld_tx_data[124], in_pld_tx_data[123], in_pld_tx_data[122], in_pld_tx_data[121], in_pld_tx_data[120], in_pld_tx_data[119], in_pld_tx_data[118], in_pld_tx_data[117], in_pld_tx_data[116], in_pld_tx_data[115], in_pld_tx_data[114], in_pld_tx_data[113], in_pld_tx_data[112], in_pld_tx_data[111], in_pld_tx_data[110], in_pld_tx_data[109], in_pld_tx_data[108], in_pld_tx_data[107], in_pld_tx_data[106], in_pld_tx_data[105], in_pld_tx_data[104], in_pld_tx_data[103], in_pld_tx_data[102], in_pld_tx_data[101], in_pld_tx_data[100], in_pld_tx_data[99], in_pld_tx_data[98], in_pld_tx_data[97], in_pld_tx_data[96], in_pld_tx_data[95], in_pld_tx_data[94], in_pld_tx_data[93], in_pld_tx_data[92], in_pld_tx_data[91], in_pld_tx_data[90], in_pld_tx_data[89], in_pld_tx_data[88], in_pld_tx_data[87], in_pld_tx_data[86], in_pld_tx_data[85], in_pld_tx_data[84], in_pld_tx_data[83], in_pld_tx_data[82], in_pld_tx_data[81], in_pld_tx_data[80], in_pld_tx_data[79], in_pld_tx_data[78], in_pld_tx_data[77], in_pld_tx_data[76], in_pld_tx_data[75], in_pld_tx_data[74], in_pld_tx_data[73], in_pld_tx_data[72], in_pld_tx_data[71], in_pld_tx_data[70], in_pld_tx_data[69], in_pld_tx_data[68], in_pld_tx_data[67], in_pld_tx_data[66], in_pld_tx_data[65], in_pld_tx_data[64], in_pld_tx_data[63], in_pld_tx_data[62], in_pld_tx_data[61], in_pld_tx_data[60], in_pld_tx_data[59], in_pld_tx_data[58], in_pld_tx_data[57], in_pld_tx_data[56], in_pld_tx_data[55], in_pld_tx_data[54], in_pld_tx_data[53], in_pld_tx_data[52], in_pld_tx_data[51], in_pld_tx_data[50], in_pld_tx_data[49], in_pld_tx_data[48], in_pld_tx_data[47], in_pld_tx_data[46], in_pld_tx_data[45], in_pld_tx_data[44], in_pld_tx_data[43], in_pld_tx_data[42], in_pld_tx_data[41], in_pld_tx_data[40], in_pld_tx_data[39], in_pld_tx_data[38], in_pld_tx_data[37], in_pld_tx_data[36], in_pld_tx_data[35], in_pld_tx_data[34], in_pld_tx_data[33], in_pld_tx_data[32], in_pld_tx_data[31], in_pld_tx_data[30], in_pld_tx_data[29], in_pld_tx_data[28], in_pld_tx_data[27], in_pld_tx_data[26], in_pld_tx_data[25], in_pld_tx_data[24], in_pld_tx_data[23], in_pld_tx_data[22], in_pld_tx_data[21], in_pld_tx_data[20], in_pld_tx_data[19], in_pld_tx_data[18], in_pld_tx_data[17], in_pld_tx_data[16], in_pld_tx_data[15], in_pld_tx_data[14], in_pld_tx_data[13], in_pld_tx_data[12], in_pld_tx_data[11], in_pld_tx_data[10], in_pld_tx_data[9], in_pld_tx_data[8], in_pld_tx_data[7], in_pld_tx_data[6], in_pld_tx_data[5], in_pld_tx_data[4], in_pld_tx_data[3], in_pld_tx_data[2], in_pld_tx_data[1], in_pld_tx_data[0]}),
				.pld_txelecidle(in_pld_txelecidle),
				.pld_uhsif_tx_clk(in_pld_uhsif_tx_clk),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.hip_clk_out_div_by_2_wire(),
				.hip_clk_out_wire(),
				.int_pldif_pmaif_tx_pld_clk(),
				.pld_10g_tx_burst_en_exe_10g_fastreg(),
				.pld_10g_tx_burst_en_exe_plddirect_reg(),
				.pld_10g_tx_data_valid_2ff_delay1_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay3_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg(),
				.pld_10g_tx_data_valid_fastreg(),
				.pld_10g_tx_data_valid_plddirect_fastreg(),
				.pld_pcs_tx_clk_out_pma_wire(),
				.pld_pma_tx_clk_out_wire(),
				.pld_pmaif_tx_pld_rst_n_reg(),
				.pld_polinv_tx_10g_pcsdirect_reg(),
				.pld_polinv_tx_8g_reg(),
				.pld_polinv_tx_pat_reg(),
				.pld_tx_clk_fifo(),
				.pld_tx_control_fifo(),
				.pld_tx_control_hi_10g_reg(),
				.pld_tx_control_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_10g_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_8g_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_control_lo_plddirect_fastreg(),
				.pld_tx_control_lo_plddirect_reg(),
				.pld_tx_data_hi_reg(),
				.pld_tx_data_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_10g_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_8g_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_data_lo_plddirect_fastreg(),
				.pld_tx_data_lo_plddirect_reg(),
				.pld_uhsif_reg(),
				.pma_tx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_hip_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6:0] = 7'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17:0] = 18'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8:0] = 9'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127:0] = 128'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4:0] = 5'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2:0] = 3'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_full = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_full_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out = 1'b0;
		end // if not generate
		
		//output assignments
		assign out_avmmreaddata_hssi_10g_rx_pcs = {w_hssi_10g_rx_pcs_avmmreaddata[7], w_hssi_10g_rx_pcs_avmmreaddata[6], w_hssi_10g_rx_pcs_avmmreaddata[5], w_hssi_10g_rx_pcs_avmmreaddata[4], w_hssi_10g_rx_pcs_avmmreaddata[3], w_hssi_10g_rx_pcs_avmmreaddata[2], w_hssi_10g_rx_pcs_avmmreaddata[1], w_hssi_10g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_10g_tx_pcs = {w_hssi_10g_tx_pcs_avmmreaddata[7], w_hssi_10g_tx_pcs_avmmreaddata[6], w_hssi_10g_tx_pcs_avmmreaddata[5], w_hssi_10g_tx_pcs_avmmreaddata[4], w_hssi_10g_tx_pcs_avmmreaddata[3], w_hssi_10g_tx_pcs_avmmreaddata[2], w_hssi_10g_tx_pcs_avmmreaddata[1], w_hssi_10g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_rx_pcs = {w_hssi_8g_rx_pcs_avmmreaddata[7], w_hssi_8g_rx_pcs_avmmreaddata[6], w_hssi_8g_rx_pcs_avmmreaddata[5], w_hssi_8g_rx_pcs_avmmreaddata[4], w_hssi_8g_rx_pcs_avmmreaddata[3], w_hssi_8g_rx_pcs_avmmreaddata[2], w_hssi_8g_rx_pcs_avmmreaddata[1], w_hssi_8g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_tx_pcs = {w_hssi_8g_tx_pcs_avmmreaddata[7], w_hssi_8g_tx_pcs_avmmreaddata[6], w_hssi_8g_tx_pcs_avmmreaddata[5], w_hssi_8g_tx_pcs_avmmreaddata[4], w_hssi_8g_tx_pcs_avmmreaddata[3], w_hssi_8g_tx_pcs_avmmreaddata[2], w_hssi_8g_tx_pcs_avmmreaddata[1], w_hssi_8g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pcs_pma_interface = {w_hssi_common_pcs_pma_interface_avmmreaddata[7], w_hssi_common_pcs_pma_interface_avmmreaddata[6], w_hssi_common_pcs_pma_interface_avmmreaddata[5], w_hssi_common_pcs_pma_interface_avmmreaddata[4], w_hssi_common_pcs_pma_interface_avmmreaddata[3], w_hssi_common_pcs_pma_interface_avmmreaddata[2], w_hssi_common_pcs_pma_interface_avmmreaddata[1], w_hssi_common_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pld_pcs_interface = {w_hssi_common_pld_pcs_interface_avmmreaddata[7], w_hssi_common_pld_pcs_interface_avmmreaddata[6], w_hssi_common_pld_pcs_interface_avmmreaddata[5], w_hssi_common_pld_pcs_interface_avmmreaddata[4], w_hssi_common_pld_pcs_interface_avmmreaddata[3], w_hssi_common_pld_pcs_interface_avmmreaddata[2], w_hssi_common_pld_pcs_interface_avmmreaddata[1], w_hssi_common_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_rx_pcs = {w_hssi_fifo_rx_pcs_avmmreaddata[7], w_hssi_fifo_rx_pcs_avmmreaddata[6], w_hssi_fifo_rx_pcs_avmmreaddata[5], w_hssi_fifo_rx_pcs_avmmreaddata[4], w_hssi_fifo_rx_pcs_avmmreaddata[3], w_hssi_fifo_rx_pcs_avmmreaddata[2], w_hssi_fifo_rx_pcs_avmmreaddata[1], w_hssi_fifo_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_tx_pcs = {w_hssi_fifo_tx_pcs_avmmreaddata[7], w_hssi_fifo_tx_pcs_avmmreaddata[6], w_hssi_fifo_tx_pcs_avmmreaddata[5], w_hssi_fifo_tx_pcs_avmmreaddata[4], w_hssi_fifo_tx_pcs_avmmreaddata[3], w_hssi_fifo_tx_pcs_avmmreaddata[2], w_hssi_fifo_tx_pcs_avmmreaddata[1], w_hssi_fifo_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_rx_pcs = {w_hssi_gen3_rx_pcs_avmmreaddata[7], w_hssi_gen3_rx_pcs_avmmreaddata[6], w_hssi_gen3_rx_pcs_avmmreaddata[5], w_hssi_gen3_rx_pcs_avmmreaddata[4], w_hssi_gen3_rx_pcs_avmmreaddata[3], w_hssi_gen3_rx_pcs_avmmreaddata[2], w_hssi_gen3_rx_pcs_avmmreaddata[1], w_hssi_gen3_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_tx_pcs = {w_hssi_gen3_tx_pcs_avmmreaddata[7], w_hssi_gen3_tx_pcs_avmmreaddata[6], w_hssi_gen3_tx_pcs_avmmreaddata[5], w_hssi_gen3_tx_pcs_avmmreaddata[4], w_hssi_gen3_tx_pcs_avmmreaddata[3], w_hssi_gen3_tx_pcs_avmmreaddata[2], w_hssi_gen3_tx_pcs_avmmreaddata[1], w_hssi_gen3_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_rx_pcs = {w_hssi_krfec_rx_pcs_avmmreaddata[7], w_hssi_krfec_rx_pcs_avmmreaddata[6], w_hssi_krfec_rx_pcs_avmmreaddata[5], w_hssi_krfec_rx_pcs_avmmreaddata[4], w_hssi_krfec_rx_pcs_avmmreaddata[3], w_hssi_krfec_rx_pcs_avmmreaddata[2], w_hssi_krfec_rx_pcs_avmmreaddata[1], w_hssi_krfec_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_tx_pcs = {w_hssi_krfec_tx_pcs_avmmreaddata[7], w_hssi_krfec_tx_pcs_avmmreaddata[6], w_hssi_krfec_tx_pcs_avmmreaddata[5], w_hssi_krfec_tx_pcs_avmmreaddata[4], w_hssi_krfec_tx_pcs_avmmreaddata[3], w_hssi_krfec_tx_pcs_avmmreaddata[2], w_hssi_krfec_tx_pcs_avmmreaddata[1], w_hssi_krfec_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen1_2 = {w_hssi_pipe_gen1_2_avmmreaddata[7], w_hssi_pipe_gen1_2_avmmreaddata[6], w_hssi_pipe_gen1_2_avmmreaddata[5], w_hssi_pipe_gen1_2_avmmreaddata[4], w_hssi_pipe_gen1_2_avmmreaddata[3], w_hssi_pipe_gen1_2_avmmreaddata[2], w_hssi_pipe_gen1_2_avmmreaddata[1], w_hssi_pipe_gen1_2_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen3 = {w_hssi_pipe_gen3_avmmreaddata[7], w_hssi_pipe_gen3_avmmreaddata[6], w_hssi_pipe_gen3_avmmreaddata[5], w_hssi_pipe_gen3_avmmreaddata[4], w_hssi_pipe_gen3_avmmreaddata[3], w_hssi_pipe_gen3_avmmreaddata[2], w_hssi_pipe_gen3_avmmreaddata[1], w_hssi_pipe_gen3_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pcs_pma_interface = {w_hssi_rx_pcs_pma_interface_avmmreaddata[7], w_hssi_rx_pcs_pma_interface_avmmreaddata[6], w_hssi_rx_pcs_pma_interface_avmmreaddata[5], w_hssi_rx_pcs_pma_interface_avmmreaddata[4], w_hssi_rx_pcs_pma_interface_avmmreaddata[3], w_hssi_rx_pcs_pma_interface_avmmreaddata[2], w_hssi_rx_pcs_pma_interface_avmmreaddata[1], w_hssi_rx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pld_pcs_interface = {w_hssi_rx_pld_pcs_interface_avmmreaddata[7], w_hssi_rx_pld_pcs_interface_avmmreaddata[6], w_hssi_rx_pld_pcs_interface_avmmreaddata[5], w_hssi_rx_pld_pcs_interface_avmmreaddata[4], w_hssi_rx_pld_pcs_interface_avmmreaddata[3], w_hssi_rx_pld_pcs_interface_avmmreaddata[2], w_hssi_rx_pld_pcs_interface_avmmreaddata[1], w_hssi_rx_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pcs_pma_interface = {w_hssi_tx_pcs_pma_interface_avmmreaddata[7], w_hssi_tx_pcs_pma_interface_avmmreaddata[6], w_hssi_tx_pcs_pma_interface_avmmreaddata[5], w_hssi_tx_pcs_pma_interface_avmmreaddata[4], w_hssi_tx_pcs_pma_interface_avmmreaddata[3], w_hssi_tx_pcs_pma_interface_avmmreaddata[2], w_hssi_tx_pcs_pma_interface_avmmreaddata[1], w_hssi_tx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pld_pcs_interface = {w_hssi_tx_pld_pcs_interface_avmmreaddata[7], w_hssi_tx_pld_pcs_interface_avmmreaddata[6], w_hssi_tx_pld_pcs_interface_avmmreaddata[5], w_hssi_tx_pld_pcs_interface_avmmreaddata[4], w_hssi_tx_pld_pcs_interface_avmmreaddata[3], w_hssi_tx_pld_pcs_interface_avmmreaddata[2], w_hssi_tx_pld_pcs_interface_avmmreaddata[1], w_hssi_tx_pld_pcs_interface_avmmreaddata[0]};
		assign out_blockselect_hssi_10g_rx_pcs = w_hssi_10g_rx_pcs_blockselect;
		assign out_blockselect_hssi_10g_tx_pcs = w_hssi_10g_tx_pcs_blockselect;
		assign out_blockselect_hssi_8g_rx_pcs = w_hssi_8g_rx_pcs_blockselect;
		assign out_blockselect_hssi_8g_tx_pcs = w_hssi_8g_tx_pcs_blockselect;
		assign out_blockselect_hssi_common_pcs_pma_interface = w_hssi_common_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_common_pld_pcs_interface = w_hssi_common_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_fifo_rx_pcs = w_hssi_fifo_rx_pcs_blockselect;
		assign out_blockselect_hssi_fifo_tx_pcs = w_hssi_fifo_tx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_rx_pcs = w_hssi_gen3_rx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_tx_pcs = w_hssi_gen3_tx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_rx_pcs = w_hssi_krfec_rx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_tx_pcs = w_hssi_krfec_tx_pcs_blockselect;
		assign out_blockselect_hssi_pipe_gen1_2 = w_hssi_pipe_gen1_2_blockselect;
		assign out_blockselect_hssi_pipe_gen3 = w_hssi_pipe_gen3_blockselect;
		assign out_blockselect_hssi_rx_pcs_pma_interface = w_hssi_rx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_rx_pld_pcs_interface = w_hssi_rx_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_tx_pcs_pma_interface = w_hssi_tx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_tx_pld_pcs_interface = w_hssi_tx_pld_pcs_interface_blockselect;
		assign out_bond_pcs10g_out_bot = {w_hssi_10g_tx_pcs_distdwn_out_rden, w_hssi_10g_tx_pcs_distdwn_out_wren, w_hssi_10g_tx_pcs_distdwn_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs10g_out_top = {w_hssi_10g_tx_pcs_distup_out_rden, w_hssi_10g_tx_pcs_distup_out_wren, w_hssi_10g_tx_pcs_distup_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs8g_out_bot = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down, w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_down, w_hssi_8g_tx_pcs_wr_enable_out_chnl_down, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_down, w_hssi_8g_rx_pcs_wr_enable_out_chnl_down, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[0]};
		assign out_bond_pcs8g_out_top = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up, w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_up, w_hssi_8g_tx_pcs_wr_enable_out_chnl_up, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_up, w_hssi_8g_rx_pcs_wr_enable_out_chnl_up, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[0]};
		assign out_bond_pmaif_out_bot = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[0]};
		assign out_bond_pmaif_out_top = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[0]};
		assign out_hip_clk_out = {w_hssi_common_pld_pcs_interface_hip_cmn_clk[1], w_hssi_common_pld_pcs_interface_hip_cmn_clk[0], w_hssi_tx_pld_pcs_interface_hip_tx_clk};
		assign out_hip_ctrl_out = {w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[4], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[3], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[2], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[1], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[0], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[0]};
		assign out_hip_iocsr_rdy = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
		assign out_hip_iocsr_rdy_dly = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
		assign out_hip_nfrzdrv = w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
		assign out_hip_npor = w_hssi_common_pld_pcs_interface_hip_npor;
		assign out_hip_rx_data = {w_hssi_rx_pld_pcs_interface_hip_rx_data[50], w_hssi_rx_pld_pcs_interface_hip_rx_data[49], w_hssi_rx_pld_pcs_interface_hip_rx_data[48], w_hssi_rx_pld_pcs_interface_hip_rx_data[47], w_hssi_rx_pld_pcs_interface_hip_rx_data[46], w_hssi_rx_pld_pcs_interface_hip_rx_data[45], w_hssi_rx_pld_pcs_interface_hip_rx_data[44], w_hssi_rx_pld_pcs_interface_hip_rx_data[43], w_hssi_rx_pld_pcs_interface_hip_rx_data[42], w_hssi_rx_pld_pcs_interface_hip_rx_data[41], w_hssi_rx_pld_pcs_interface_hip_rx_data[40], w_hssi_rx_pld_pcs_interface_hip_rx_data[39], w_hssi_rx_pld_pcs_interface_hip_rx_data[38], w_hssi_rx_pld_pcs_interface_hip_rx_data[37], w_hssi_rx_pld_pcs_interface_hip_rx_data[36], w_hssi_rx_pld_pcs_interface_hip_rx_data[35], w_hssi_rx_pld_pcs_interface_hip_rx_data[34], w_hssi_rx_pld_pcs_interface_hip_rx_data[33], w_hssi_rx_pld_pcs_interface_hip_rx_data[32], w_hssi_rx_pld_pcs_interface_hip_rx_data[31], w_hssi_rx_pld_pcs_interface_hip_rx_data[30], w_hssi_rx_pld_pcs_interface_hip_rx_data[29], w_hssi_rx_pld_pcs_interface_hip_rx_data[28], w_hssi_rx_pld_pcs_interface_hip_rx_data[27], w_hssi_rx_pld_pcs_interface_hip_rx_data[26], w_hssi_rx_pld_pcs_interface_hip_rx_data[25], w_hssi_rx_pld_pcs_interface_hip_rx_data[24], w_hssi_rx_pld_pcs_interface_hip_rx_data[23], w_hssi_rx_pld_pcs_interface_hip_rx_data[22], w_hssi_rx_pld_pcs_interface_hip_rx_data[21], w_hssi_rx_pld_pcs_interface_hip_rx_data[20], w_hssi_rx_pld_pcs_interface_hip_rx_data[19], w_hssi_rx_pld_pcs_interface_hip_rx_data[18], w_hssi_rx_pld_pcs_interface_hip_rx_data[17], w_hssi_rx_pld_pcs_interface_hip_rx_data[16], w_hssi_rx_pld_pcs_interface_hip_rx_data[15], w_hssi_rx_pld_pcs_interface_hip_rx_data[14], w_hssi_rx_pld_pcs_interface_hip_rx_data[13], w_hssi_rx_pld_pcs_interface_hip_rx_data[12], w_hssi_rx_pld_pcs_interface_hip_rx_data[11], w_hssi_rx_pld_pcs_interface_hip_rx_data[10], w_hssi_rx_pld_pcs_interface_hip_rx_data[9], w_hssi_rx_pld_pcs_interface_hip_rx_data[8], w_hssi_rx_pld_pcs_interface_hip_rx_data[7], w_hssi_rx_pld_pcs_interface_hip_rx_data[6], w_hssi_rx_pld_pcs_interface_hip_rx_data[5], w_hssi_rx_pld_pcs_interface_hip_rx_data[4], w_hssi_rx_pld_pcs_interface_hip_rx_data[3], w_hssi_rx_pld_pcs_interface_hip_rx_data[2], w_hssi_rx_pld_pcs_interface_hip_rx_data[1], w_hssi_rx_pld_pcs_interface_hip_rx_data[0]};
		assign out_hip_usermode = w_hssi_common_pld_pcs_interface_hip_usermode;
		assign out_pld_10g_krfec_rx_blk_lock = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
		assign out_pld_10g_krfec_rx_diag_data_status = {w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1], w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[0]};
		assign out_pld_10g_krfec_rx_frame = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
		assign out_pld_10g_krfec_tx_frame = w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
		assign out_pld_10g_rx_align_val = w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
		assign out_pld_10g_rx_crc32_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
		assign out_pld_10g_rx_data_valid = w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
		assign out_pld_10g_rx_empty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
		assign out_pld_10g_rx_fifo_del = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
		assign out_pld_10g_rx_fifo_insert = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
		assign out_pld_10g_rx_fifo_num = {w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[3], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[2], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[1], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[0]};
		assign out_pld_10g_rx_frame_lock = w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
		assign out_pld_10g_rx_hi_ber = w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
		assign out_pld_10g_rx_oflw_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
		assign out_pld_10g_rx_pempty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
		assign out_pld_10g_rx_pfull = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
		assign out_pld_10g_tx_burst_en_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
		assign out_pld_10g_tx_empty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
		assign out_pld_10g_tx_fifo_num = {w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[2], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[1], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[0]};
		assign out_pld_10g_tx_full = w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
		assign out_pld_10g_tx_pempty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
		assign out_pld_10g_tx_pfull = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
		assign out_pld_10g_tx_wordslip_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
		assign out_pld_8g_a1a2_k1k2_flag = {w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[2], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[1], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[0]};
		assign out_pld_8g_empty_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
		assign out_pld_8g_empty_rx = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
		assign out_pld_8g_empty_tx = w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
		assign out_pld_8g_full_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
		assign out_pld_8g_full_rx = w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
		assign out_pld_8g_full_tx = w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
		assign out_pld_8g_rxelecidle = w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
		assign out_pld_8g_signal_detect_out = w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
		assign out_pld_8g_wa_boundary = {w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0]};
		assign out_pld_krfec_tx_alignment = w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
		assign out_pld_pcs_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
		assign out_pld_pcs_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
		assign out_pld_pma_adapt_done = w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
		assign out_pld_pma_clkdiv_rx_user = w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
		assign out_pld_pma_clkdiv_tx_user = w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
		assign out_pld_pma_clklow = w_hssi_common_pld_pcs_interface_pld_pma_clklow;
		assign out_pld_pma_fref = w_hssi_common_pld_pcs_interface_pld_pma_fref;
		assign out_pld_pma_hclk = w_hssi_common_pld_pcs_interface_pld_pma_hclk;
		assign out_pld_pma_pcie_sw_done = {w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1], w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[0]};
		assign out_pld_pma_pfdmode_lock = w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
		assign out_pld_pma_reserved_in = {w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[3], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[2], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[1], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[0]};
		assign out_pld_pma_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
		assign out_pld_pma_rx_detect_valid = w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
		assign out_pld_pma_rx_found = w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
		assign out_pld_pma_rxpll_lock = w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
		assign out_pld_pma_signal_ok = w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
		assign out_pld_pma_testbus = {w_hssi_common_pld_pcs_interface_pld_pma_testbus[7], w_hssi_common_pld_pcs_interface_pld_pma_testbus[6], w_hssi_common_pld_pcs_interface_pld_pma_testbus[5], w_hssi_common_pld_pcs_interface_pld_pma_testbus[4], w_hssi_common_pld_pcs_interface_pld_pma_testbus[3], w_hssi_common_pld_pcs_interface_pld_pma_testbus[2], w_hssi_common_pld_pcs_interface_pld_pma_testbus[1], w_hssi_common_pld_pcs_interface_pld_pma_testbus[0]};
		assign out_pld_pma_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
		assign out_pld_pmaif_mask_tx_pll = w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
		assign out_pld_reserved_out = {w_hssi_common_pld_pcs_interface_pld_reserved_out[9], w_hssi_common_pld_pcs_interface_pld_reserved_out[8], w_hssi_common_pld_pcs_interface_pld_reserved_out[7], w_hssi_common_pld_pcs_interface_pld_reserved_out[6], w_hssi_common_pld_pcs_interface_pld_reserved_out[5], w_hssi_common_pld_pcs_interface_pld_reserved_out[4], w_hssi_common_pld_pcs_interface_pld_reserved_out[3], w_hssi_common_pld_pcs_interface_pld_reserved_out[2], w_hssi_common_pld_pcs_interface_pld_reserved_out[1], w_hssi_common_pld_pcs_interface_pld_reserved_out[0]};
		assign out_pld_rx_control = {w_hssi_rx_pld_pcs_interface_pld_rx_control[19], w_hssi_rx_pld_pcs_interface_pld_rx_control[18], w_hssi_rx_pld_pcs_interface_pld_rx_control[17], w_hssi_rx_pld_pcs_interface_pld_rx_control[16], w_hssi_rx_pld_pcs_interface_pld_rx_control[15], w_hssi_rx_pld_pcs_interface_pld_rx_control[14], w_hssi_rx_pld_pcs_interface_pld_rx_control[13], w_hssi_rx_pld_pcs_interface_pld_rx_control[12], w_hssi_rx_pld_pcs_interface_pld_rx_control[11], w_hssi_rx_pld_pcs_interface_pld_rx_control[10], w_hssi_rx_pld_pcs_interface_pld_rx_control[9], w_hssi_rx_pld_pcs_interface_pld_rx_control[8], w_hssi_rx_pld_pcs_interface_pld_rx_control[7], w_hssi_rx_pld_pcs_interface_pld_rx_control[6], w_hssi_rx_pld_pcs_interface_pld_rx_control[5], w_hssi_rx_pld_pcs_interface_pld_rx_control[4], w_hssi_rx_pld_pcs_interface_pld_rx_control[3], w_hssi_rx_pld_pcs_interface_pld_rx_control[2], w_hssi_rx_pld_pcs_interface_pld_rx_control[1], w_hssi_rx_pld_pcs_interface_pld_rx_control[0]};
		assign out_pld_rx_data = {w_hssi_rx_pld_pcs_interface_pld_rx_data[127], w_hssi_rx_pld_pcs_interface_pld_rx_data[126], w_hssi_rx_pld_pcs_interface_pld_rx_data[125], w_hssi_rx_pld_pcs_interface_pld_rx_data[124], w_hssi_rx_pld_pcs_interface_pld_rx_data[123], w_hssi_rx_pld_pcs_interface_pld_rx_data[122], w_hssi_rx_pld_pcs_interface_pld_rx_data[121], w_hssi_rx_pld_pcs_interface_pld_rx_data[120], w_hssi_rx_pld_pcs_interface_pld_rx_data[119], w_hssi_rx_pld_pcs_interface_pld_rx_data[118], w_hssi_rx_pld_pcs_interface_pld_rx_data[117], w_hssi_rx_pld_pcs_interface_pld_rx_data[116], w_hssi_rx_pld_pcs_interface_pld_rx_data[115], w_hssi_rx_pld_pcs_interface_pld_rx_data[114], w_hssi_rx_pld_pcs_interface_pld_rx_data[113], w_hssi_rx_pld_pcs_interface_pld_rx_data[112], w_hssi_rx_pld_pcs_interface_pld_rx_data[111], w_hssi_rx_pld_pcs_interface_pld_rx_data[110], w_hssi_rx_pld_pcs_interface_pld_rx_data[109], w_hssi_rx_pld_pcs_interface_pld_rx_data[108], w_hssi_rx_pld_pcs_interface_pld_rx_data[107], w_hssi_rx_pld_pcs_interface_pld_rx_data[106], w_hssi_rx_pld_pcs_interface_pld_rx_data[105], w_hssi_rx_pld_pcs_interface_pld_rx_data[104], w_hssi_rx_pld_pcs_interface_pld_rx_data[103], w_hssi_rx_pld_pcs_interface_pld_rx_data[102], w_hssi_rx_pld_pcs_interface_pld_rx_data[101], w_hssi_rx_pld_pcs_interface_pld_rx_data[100], w_hssi_rx_pld_pcs_interface_pld_rx_data[99], w_hssi_rx_pld_pcs_interface_pld_rx_data[98], w_hssi_rx_pld_pcs_interface_pld_rx_data[97], w_hssi_rx_pld_pcs_interface_pld_rx_data[96], w_hssi_rx_pld_pcs_interface_pld_rx_data[95], w_hssi_rx_pld_pcs_interface_pld_rx_data[94], w_hssi_rx_pld_pcs_interface_pld_rx_data[93], w_hssi_rx_pld_pcs_interface_pld_rx_data[92], w_hssi_rx_pld_pcs_interface_pld_rx_data[91], w_hssi_rx_pld_pcs_interface_pld_rx_data[90], w_hssi_rx_pld_pcs_interface_pld_rx_data[89], w_hssi_rx_pld_pcs_interface_pld_rx_data[88], w_hssi_rx_pld_pcs_interface_pld_rx_data[87], w_hssi_rx_pld_pcs_interface_pld_rx_data[86], w_hssi_rx_pld_pcs_interface_pld_rx_data[85], w_hssi_rx_pld_pcs_interface_pld_rx_data[84], w_hssi_rx_pld_pcs_interface_pld_rx_data[83], w_hssi_rx_pld_pcs_interface_pld_rx_data[82], w_hssi_rx_pld_pcs_interface_pld_rx_data[81], w_hssi_rx_pld_pcs_interface_pld_rx_data[80], w_hssi_rx_pld_pcs_interface_pld_rx_data[79], w_hssi_rx_pld_pcs_interface_pld_rx_data[78], w_hssi_rx_pld_pcs_interface_pld_rx_data[77], w_hssi_rx_pld_pcs_interface_pld_rx_data[76], w_hssi_rx_pld_pcs_interface_pld_rx_data[75], w_hssi_rx_pld_pcs_interface_pld_rx_data[74], w_hssi_rx_pld_pcs_interface_pld_rx_data[73], w_hssi_rx_pld_pcs_interface_pld_rx_data[72], w_hssi_rx_pld_pcs_interface_pld_rx_data[71], w_hssi_rx_pld_pcs_interface_pld_rx_data[70], w_hssi_rx_pld_pcs_interface_pld_rx_data[69], w_hssi_rx_pld_pcs_interface_pld_rx_data[68], w_hssi_rx_pld_pcs_interface_pld_rx_data[67], w_hssi_rx_pld_pcs_interface_pld_rx_data[66], w_hssi_rx_pld_pcs_interface_pld_rx_data[65], w_hssi_rx_pld_pcs_interface_pld_rx_data[64], w_hssi_rx_pld_pcs_interface_pld_rx_data[63], w_hssi_rx_pld_pcs_interface_pld_rx_data[62], w_hssi_rx_pld_pcs_interface_pld_rx_data[61], w_hssi_rx_pld_pcs_interface_pld_rx_data[60], w_hssi_rx_pld_pcs_interface_pld_rx_data[59], w_hssi_rx_pld_pcs_interface_pld_rx_data[58], w_hssi_rx_pld_pcs_interface_pld_rx_data[57], w_hssi_rx_pld_pcs_interface_pld_rx_data[56], w_hssi_rx_pld_pcs_interface_pld_rx_data[55], w_hssi_rx_pld_pcs_interface_pld_rx_data[54], w_hssi_rx_pld_pcs_interface_pld_rx_data[53], w_hssi_rx_pld_pcs_interface_pld_rx_data[52], w_hssi_rx_pld_pcs_interface_pld_rx_data[51], w_hssi_rx_pld_pcs_interface_pld_rx_data[50], w_hssi_rx_pld_pcs_interface_pld_rx_data[49], w_hssi_rx_pld_pcs_interface_pld_rx_data[48], w_hssi_rx_pld_pcs_interface_pld_rx_data[47], w_hssi_rx_pld_pcs_interface_pld_rx_data[46], w_hssi_rx_pld_pcs_interface_pld_rx_data[45], w_hssi_rx_pld_pcs_interface_pld_rx_data[44], w_hssi_rx_pld_pcs_interface_pld_rx_data[43], w_hssi_rx_pld_pcs_interface_pld_rx_data[42], w_hssi_rx_pld_pcs_interface_pld_rx_data[41], w_hssi_rx_pld_pcs_interface_pld_rx_data[40], w_hssi_rx_pld_pcs_interface_pld_rx_data[39], w_hssi_rx_pld_pcs_interface_pld_rx_data[38], w_hssi_rx_pld_pcs_interface_pld_rx_data[37], w_hssi_rx_pld_pcs_interface_pld_rx_data[36], w_hssi_rx_pld_pcs_interface_pld_rx_data[35], w_hssi_rx_pld_pcs_interface_pld_rx_data[34], w_hssi_rx_pld_pcs_interface_pld_rx_data[33], w_hssi_rx_pld_pcs_interface_pld_rx_data[32], w_hssi_rx_pld_pcs_interface_pld_rx_data[31], w_hssi_rx_pld_pcs_interface_pld_rx_data[30], w_hssi_rx_pld_pcs_interface_pld_rx_data[29], w_hssi_rx_pld_pcs_interface_pld_rx_data[28], w_hssi_rx_pld_pcs_interface_pld_rx_data[27], w_hssi_rx_pld_pcs_interface_pld_rx_data[26], w_hssi_rx_pld_pcs_interface_pld_rx_data[25], w_hssi_rx_pld_pcs_interface_pld_rx_data[24], w_hssi_rx_pld_pcs_interface_pld_rx_data[23], w_hssi_rx_pld_pcs_interface_pld_rx_data[22], w_hssi_rx_pld_pcs_interface_pld_rx_data[21], w_hssi_rx_pld_pcs_interface_pld_rx_data[20], w_hssi_rx_pld_pcs_interface_pld_rx_data[19], w_hssi_rx_pld_pcs_interface_pld_rx_data[18], w_hssi_rx_pld_pcs_interface_pld_rx_data[17], w_hssi_rx_pld_pcs_interface_pld_rx_data[16], w_hssi_rx_pld_pcs_interface_pld_rx_data[15], w_hssi_rx_pld_pcs_interface_pld_rx_data[14], w_hssi_rx_pld_pcs_interface_pld_rx_data[13], w_hssi_rx_pld_pcs_interface_pld_rx_data[12], w_hssi_rx_pld_pcs_interface_pld_rx_data[11], w_hssi_rx_pld_pcs_interface_pld_rx_data[10], w_hssi_rx_pld_pcs_interface_pld_rx_data[9], w_hssi_rx_pld_pcs_interface_pld_rx_data[8], w_hssi_rx_pld_pcs_interface_pld_rx_data[7], w_hssi_rx_pld_pcs_interface_pld_rx_data[6], w_hssi_rx_pld_pcs_interface_pld_rx_data[5], w_hssi_rx_pld_pcs_interface_pld_rx_data[4], w_hssi_rx_pld_pcs_interface_pld_rx_data[3], w_hssi_rx_pld_pcs_interface_pld_rx_data[2], w_hssi_rx_pld_pcs_interface_pld_rx_data[1], w_hssi_rx_pld_pcs_interface_pld_rx_data[0]};
		assign out_pld_rx_prbs_done = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
		assign out_pld_rx_prbs_err = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
		assign out_pld_test_data = {w_hssi_common_pld_pcs_interface_pld_test_data[19], w_hssi_common_pld_pcs_interface_pld_test_data[18], w_hssi_common_pld_pcs_interface_pld_test_data[17], w_hssi_common_pld_pcs_interface_pld_test_data[16], w_hssi_common_pld_pcs_interface_pld_test_data[15], w_hssi_common_pld_pcs_interface_pld_test_data[14], w_hssi_common_pld_pcs_interface_pld_test_data[13], w_hssi_common_pld_pcs_interface_pld_test_data[12], w_hssi_common_pld_pcs_interface_pld_test_data[11], w_hssi_common_pld_pcs_interface_pld_test_data[10], w_hssi_common_pld_pcs_interface_pld_test_data[9], w_hssi_common_pld_pcs_interface_pld_test_data[8], w_hssi_common_pld_pcs_interface_pld_test_data[7], w_hssi_common_pld_pcs_interface_pld_test_data[6], w_hssi_common_pld_pcs_interface_pld_test_data[5], w_hssi_common_pld_pcs_interface_pld_test_data[4], w_hssi_common_pld_pcs_interface_pld_test_data[3], w_hssi_common_pld_pcs_interface_pld_test_data[2], w_hssi_common_pld_pcs_interface_pld_test_data[1], w_hssi_common_pld_pcs_interface_pld_test_data[0]};
		assign out_pld_uhsif_lock = w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
		assign out_pld_uhsif_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
		assign out_pma_adapt_start = w_hssi_common_pcs_pma_interface_pma_adapt_start;
		assign out_pma_atpg_los_en_n = w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
		assign out_pma_csr_test_dis = w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
		assign out_pma_current_coeff = {w_hssi_common_pcs_pma_interface_pma_current_coeff[17], w_hssi_common_pcs_pma_interface_pma_current_coeff[16], w_hssi_common_pcs_pma_interface_pma_current_coeff[15], w_hssi_common_pcs_pma_interface_pma_current_coeff[14], w_hssi_common_pcs_pma_interface_pma_current_coeff[13], w_hssi_common_pcs_pma_interface_pma_current_coeff[12], w_hssi_common_pcs_pma_interface_pma_current_coeff[11], w_hssi_common_pcs_pma_interface_pma_current_coeff[10], w_hssi_common_pcs_pma_interface_pma_current_coeff[9], w_hssi_common_pcs_pma_interface_pma_current_coeff[8], w_hssi_common_pcs_pma_interface_pma_current_coeff[7], w_hssi_common_pcs_pma_interface_pma_current_coeff[6], w_hssi_common_pcs_pma_interface_pma_current_coeff[5], w_hssi_common_pcs_pma_interface_pma_current_coeff[4], w_hssi_common_pcs_pma_interface_pma_current_coeff[3], w_hssi_common_pcs_pma_interface_pma_current_coeff[2], w_hssi_common_pcs_pma_interface_pma_current_coeff[1], w_hssi_common_pcs_pma_interface_pma_current_coeff[0]};
		assign out_pma_current_rxpreset = {w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[1], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[0]};
		assign out_pma_early_eios = w_hssi_common_pcs_pma_interface_pma_early_eios;
		assign out_pma_eye_monitor = {w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0]};
		assign out_pma_interface_select = {w_hssi_common_pcs_pma_interface_pma_interface_select[1], w_hssi_common_pcs_pma_interface_pma_interface_select[0]};
		assign out_pma_ltd_b = w_hssi_common_pcs_pma_interface_pma_ltd_b;
		assign out_pma_ltr = w_hssi_common_pcs_pma_interface_pma_ltr;
		assign out_pma_nfrzdrv = w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
		assign out_pma_nrpi_freeze = w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
		assign out_pma_pcie_switch = {w_hssi_common_pcs_pma_interface_pma_pcie_switch[1], w_hssi_common_pcs_pma_interface_pma_pcie_switch[0]};
		assign out_pma_ppm_lock = w_hssi_common_pcs_pma_interface_pma_ppm_lock;
		assign out_pma_reserved_out = {w_hssi_common_pcs_pma_interface_pma_reserved_out[4], w_hssi_common_pcs_pma_interface_pma_reserved_out[3], w_hssi_common_pcs_pma_interface_pma_reserved_out[2], w_hssi_common_pcs_pma_interface_pma_reserved_out[1], w_hssi_common_pcs_pma_interface_pma_reserved_out[0]};
		assign out_pma_rs_lpbk_b = w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
		assign out_pma_rx_clkslip = w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
		assign out_pma_rx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
		assign out_pma_rxpma_rstb = w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
		assign out_pma_scan_mode_n = w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
		assign out_pma_scan_shift_n = w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
		assign out_pma_tx_bitslip = w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
		assign out_pma_tx_bonding_rstb = w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
		assign out_pma_tx_elec_idle = w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
		assign out_pma_tx_pma_data = {w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0]};
		assign out_pma_tx_qpi_pulldn = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
		assign out_pma_tx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
		assign out_pma_tx_txdetectrx = w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
		assign out_pma_txpma_rstb = w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	endgenerate
endmodule
module twentynm_pcs_rev_20nm3
	#(
	//PARAM_LIST_START
		parameter xcvr_native_mode = "mode_duplex",  // mode_duplex, mode_rx_only, mode_tx_only
		
		// parameters for twentynm_hssi_10g_rx_pcs
		parameter hssi_10g_rx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_align_del = "align_del_en", // align_del_dis|align_del_en
		parameter hssi_10g_rx_pcs_ber_bit_err_total_cnt = "bit_err_total_cnt_10g", // bit_err_total_cnt_10g
		parameter hssi_10g_rx_pcs_ber_clken = "ber_clk_dis", // ber_clk_dis|ber_clk_en
		parameter hssi_10g_rx_pcs_ber_xus_timer_window = 21'b100110001001010,
		parameter hssi_10g_rx_pcs_bitslip_mode = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_rx_pcs_blksync_bitslip_type = "bitslip_comb", // bitslip_comb|bitslip_reg
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_cnt = 3'b1,
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_type = "bitslip_match", // bitslip_match|bitslip_cnt
		parameter hssi_10g_rx_pcs_blksync_bypass = "blksync_bypass_dis", // blksync_bypass_dis|blksync_bypass_en
		parameter hssi_10g_rx_pcs_blksync_clken = "blksync_clk_dis", // blksync_clk_dis|blksync_clk_en
		parameter hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt = "enum_invalid_sh_cnt_10g", // enum_invalid_sh_cnt_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock = "knum_sh_cnt_postlock_10g", // knum_sh_cnt_postlock_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock = "knum_sh_cnt_prelock_10g", // knum_sh_cnt_prelock_10g
		parameter hssi_10g_rx_pcs_blksync_pipeln = "blksync_pipeln_dis", // blksync_pipeln_dis|blksync_pipeln_en
		parameter hssi_10g_rx_pcs_clr_errblk_cnt_en = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_control_del = "control_del_all", // control_del_all|control_del_none
		parameter hssi_10g_rx_pcs_crcchk_bypass = "crcchk_bypass_dis", // crcchk_bypass_dis|crcchk_bypass_en
		parameter hssi_10g_rx_pcs_crcchk_clken = "crcchk_clk_dis", // crcchk_clk_dis|crcchk_clk_en
		parameter hssi_10g_rx_pcs_crcchk_inv = "crcchk_inv_dis", // crcchk_inv_dis|crcchk_inv_en
		parameter hssi_10g_rx_pcs_crcchk_pipeln = "crcchk_pipeln_dis", // crcchk_pipeln_dis|crcchk_pipeln_en
		parameter hssi_10g_rx_pcs_crcflag_pipeln = "crcflag_pipeln_dis", // crcflag_pipeln_dis|crcflag_pipeln_en
		parameter hssi_10g_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_rx_pcs_dec64b66b_clken = "dec64b66b_clk_dis", // dec64b66b_clk_dis|dec64b66b_clk_en
		parameter hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass = "dec_64b66b_rxsm_bypass_dis", // dec_64b66b_rxsm_bypass_dis|dec_64b66b_rxsm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_bypass = "descrm_bypass_en", // descrm_bypass_dis|descrm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_clken = "descrm_clk_dis", // descrm_clk_dis|descrm_clk_en
		parameter hssi_10g_rx_pcs_descrm_mode = "async", // async|sync
		parameter hssi_10g_rx_pcs_descrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_dft_clk_out_sel = "rx_master_clk", // rx_master_clk|rx_gbexp_clk|rx_blksync_clk|rx_descrm_clk|rx_frmsync_clk|rx_64b66bdec_clk|rx_ber_clk|rx_rand_clk|rx_crcchk_clk|rx_wrfifo_clk|rx_rdfifo_clk|rx_fec_clk
		parameter hssi_10g_rx_pcs_dis_signal_ok = "dis_signal_ok_dis", // dis_signal_ok_dis|dis_signal_ok_en
		parameter hssi_10g_rx_pcs_dispchk_bypass = "dispchk_bypass_dis", // dispchk_bypass_dis|dispchk_bypass_en
		parameter hssi_10g_rx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_rx_pcs_fast_path = "fast_path_dis", // fast_path_dis|fast_path_en
		parameter hssi_10g_rx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_rx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_rx_pcs_fifo_double_read = "fifo_double_read_dis", // fifo_double_read_dis|fifo_double_read_en
		parameter hssi_10g_rx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_rx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_rx_pcs_force_align = "force_align_dis", // force_align_dis|force_align_en
		parameter hssi_10g_rx_pcs_frmsync_bypass = "frmsync_bypass_dis", // frmsync_bypass_dis|frmsync_bypass_en
		parameter hssi_10g_rx_pcs_frmsync_clken = "frmsync_clk_dis", // frmsync_clk_dis|frmsync_clk_en
		parameter hssi_10g_rx_pcs_frmsync_enum_scrm = "enum_scrm_default", // enum_scrm_default
		parameter hssi_10g_rx_pcs_frmsync_enum_sync = "enum_sync_default", // enum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_flag_type = "all_framing_words", // all_framing_words|location_only
		parameter hssi_10g_rx_pcs_frmsync_knum_sync = "knum_sync_default", // knum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_mfrm_length = 16'b100000000000,
		parameter hssi_10g_rx_pcs_frmsync_pipeln = "frmsync_pipeln_dis", // frmsync_pipeln_dis|frmsync_pipeln_en
		parameter hssi_10g_rx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_rx_pcs_gb_rx_idwidth = "width_32", // width_40|width_32|width_64
		parameter hssi_10g_rx_pcs_gb_rx_odwidth = "width_66", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_rx_pcs_gbexp_clken = "gbexp_clk_dis", // gbexp_clk_dis|gbexp_clk_en
		parameter hssi_10g_rx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_10g_rx_pcs_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_rx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_rx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_rx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_rx_pcs_pld_if_type = "fifo", // fifo|reg
		parameter hssi_10g_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_rx_pcs_rand_clken = "rand_clk_dis", // rand_clk_dis|rand_clk_en
		parameter hssi_10g_rx_pcs_rd_clk_sel = "rd_rx_pma_clk", // rd_rx_pld_clk|rd_rx_pma_clk|rd_refclk_dig
		parameter hssi_10g_rx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_rx_pcs_rx_fifo_write_ctrl = "blklock_stops", // blklock_stops|blklock_ignore
		parameter hssi_10g_rx_pcs_rx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_rx_pcs_rx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_rx_pcs_rx_signal_ok_sel = "synchronized_ver", // synchronized_ver|nonsync_ver
		parameter hssi_10g_rx_pcs_rx_sm_bypass = "rx_sm_bypass_dis", // rx_sm_bypass_dis|rx_sm_bypass_en
		parameter hssi_10g_rx_pcs_rx_sm_hiber = "rx_sm_hiber_en", // rx_sm_hiber_en|rx_sm_hiber_dis
		parameter hssi_10g_rx_pcs_rx_sm_pipeln = "rx_sm_pipeln_dis", // rx_sm_pipeln_dis|rx_sm_pipeln_en
		parameter hssi_10g_rx_pcs_rx_testbus_sel = "crc32_chk_testbus1", // crc32_chk_testbus1|crc32_chk_testbus2|frame_sync_testbus1|frame_sync_testbus2|dec64b66b_testbus|rxsm_testbus|ber_testbus|blksync_testbus1|blksync_testbus2|gearbox_exp_testbus|random_ver_testbus|descramble_testbus|blank_testbus|rx_fifo_testbus1|rx_fifo_testbus2
		parameter hssi_10g_rx_pcs_rx_true_b2b = "b2b", // single|b2b
		parameter hssi_10g_rx_pcs_rxfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_rx_pcs_rxfifo_full = "full_default", // full_default
		parameter hssi_10g_rx_pcs_rxfifo_mode = "phase_comp", // register_mode|clk_comp_10g|generic_interlaken|generic_basic|phase_comp|phase_comp_dv
		parameter hssi_10g_rx_pcs_rxfifo_pempty = 5'b10,
		parameter hssi_10g_rx_pcs_rxfifo_pfull = 5'b10111,
		parameter hssi_10g_rx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_rx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_rx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_10g_tx_pcs
		parameter hssi_10g_tx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_bitslip_en = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_10g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_10g_tx_pcs_comp_cnt = 8'b0,
		parameter hssi_10g_tx_pcs_compin_sel = "compin_master", // compin_master|compin_slave_top|compin_slave_bot|compin_default
		parameter hssi_10g_tx_pcs_crcgen_bypass = "crcgen_bypass_dis", // crcgen_bypass_dis|crcgen_bypass_en
		parameter hssi_10g_tx_pcs_crcgen_clken = "crcgen_clk_dis", // crcgen_clk_dis|crcgen_clk_en
		parameter hssi_10g_tx_pcs_crcgen_err = "crcgen_err_dis", // crcgen_err_dis|crcgen_err_en
		parameter hssi_10g_tx_pcs_crcgen_inv = "crcgen_inv_dis", // crcgen_inv_dis|crcgen_inv_en
		parameter hssi_10g_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_tx_pcs_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_10g_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_tx_pcs_dft_clk_out_sel = "tx_master_clk", // tx_master_clk|tx_rdfifo_clk|tx_frmgen_clk|tx_crcgen_clk|tx_64b66benc_txsm_clk|tx_scrm_clk|tx_dispgen_clk|tx_gbred_clk|tx_wrfifo_clk|tx_fec_clk
		parameter hssi_10g_tx_pcs_dispgen_bypass = "dispgen_bypass_dis", // dispgen_bypass_dis|dispgen_bypass_en
		parameter hssi_10g_tx_pcs_dispgen_clken = "dispgen_clk_dis", // dispgen_clk_dis|dispgen_clk_en
		parameter hssi_10g_tx_pcs_dispgen_err = "dispgen_err_dis", // dispgen_err_dis|dispgen_err_en
		parameter hssi_10g_tx_pcs_dispgen_pipeln = "dispgen_pipeln_dis", // dispgen_pipeln_dis|dispgen_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_bypass_pipeln = "distdwn_bypass_pipeln_dis", // distdwn_bypass_pipeln_dis|distdwn_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_master = "distdwn_master_en", // distdwn_master_en|distdwn_master_dis
		parameter hssi_10g_tx_pcs_distup_bypass_pipeln = "distup_bypass_pipeln_dis", // distup_bypass_pipeln_dis|distup_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distup_master = "distup_master_en", // distup_master_en|distup_master_dis
		parameter hssi_10g_tx_pcs_dv_bond = "dv_bond_dis", // dv_bond_en|dv_bond_dis
		parameter hssi_10g_tx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_tx_pcs_enc64b66b_txsm_clken = "enc64b66b_txsm_clk_dis", // enc64b66b_txsm_clk_dis|enc64b66b_txsm_clk_en
		parameter hssi_10g_tx_pcs_enc_64b66b_txsm_bypass = "enc_64b66b_txsm_bypass_dis", // enc_64b66b_txsm_bypass_dis|enc_64b66b_txsm_bypass_en
		parameter hssi_10g_tx_pcs_fastpath = "fastpath_dis", // fastpath_dis|fastpath_en
		parameter hssi_10g_tx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_tx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_tx_pcs_fifo_double_write = "fifo_double_write_dis", // fifo_double_write_dis|fifo_double_write_en
		parameter hssi_10g_tx_pcs_fifo_reg_fast = "fifo_reg_fast_dis", // fifo_reg_fast_dis|fifo_reg_fast_en
		parameter hssi_10g_tx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_tx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_tx_pcs_frmgen_burst = "frmgen_burst_dis", // frmgen_burst_dis|frmgen_burst_en
		parameter hssi_10g_tx_pcs_frmgen_bypass = "frmgen_bypass_dis", // frmgen_bypass_dis|frmgen_bypass_en
		parameter hssi_10g_tx_pcs_frmgen_clken = "frmgen_clk_dis", // frmgen_clk_dis|frmgen_clk_en
		parameter hssi_10g_tx_pcs_frmgen_mfrm_length = 16'b100000000000,
		parameter hssi_10g_tx_pcs_frmgen_pipeln = "frmgen_pipeln_dis", // frmgen_pipeln_dis|frmgen_pipeln_en
		parameter hssi_10g_tx_pcs_frmgen_pyld_ins = "frmgen_pyld_ins_dis", // frmgen_pyld_ins_dis|frmgen_pyld_ins_en
		parameter hssi_10g_tx_pcs_frmgen_wordslip = "frmgen_wordslip_dis", // frmgen_wordslip_dis|frmgen_wordslip_en
		parameter hssi_10g_tx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_tx_pcs_gb_pipeln_bypass = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_gb_tx_idwidth = "width_50", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_tx_pcs_gb_tx_odwidth = "width_32", // width_32|width_40|width_64
		parameter hssi_10g_tx_pcs_gbred_clken = "gbred_clk_dis", // gbred_clk_dis|gbred_clk_en
		parameter hssi_10g_tx_pcs_indv = "indv_en", // indv_en|indv_dis
		parameter hssi_10g_tx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_tx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_tx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_tx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del6|phcomp_rd_del5|phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_tx_pcs_pld_if_type = "fifo", // fifo|reg|fastreg
		parameter hssi_10g_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_tx_pcs_pseudo_random = "all_0", // two_lf|all_0
		parameter hssi_10g_tx_pcs_pseudo_seed_a = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_pseudo_seed_b = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_random_disp = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_tx_pcs_scrm_bypass = "scrm_bypass_dis", // scrm_bypass_dis|scrm_bypass_en
		parameter hssi_10g_tx_pcs_scrm_clken = "scrm_clk_dis", // scrm_clk_dis|scrm_clk_en
		parameter hssi_10g_tx_pcs_scrm_mode = "async", // async|sync
		parameter hssi_10g_tx_pcs_scrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_sh_err = "sh_err_dis", // sh_err_dis|sh_err_en
		parameter hssi_10g_tx_pcs_sop_mark = "sop_mark_dis", // sop_mark_en|sop_mark_dis
		parameter hssi_10g_tx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_tx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_tx_pcs_tx_scrm_err = "scrm_err_dis", // scrm_err_dis|scrm_err_en
		parameter hssi_10g_tx_pcs_tx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_tx_pcs_tx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_tx_pcs_tx_sm_bypass = "tx_sm_bypass_dis", // tx_sm_bypass_dis|tx_sm_bypass_en
		parameter hssi_10g_tx_pcs_tx_sm_pipeln = "tx_sm_pipeln_dis", // tx_sm_pipeln_dis|tx_sm_pipeln_en
		parameter hssi_10g_tx_pcs_tx_testbus_sel = "crc32_gen_testbus1", // crc32_gen_testbus1|crc32_gen_testbus2|disp_gen_testbus1|disp_gen_testbus2|frame_gen_testbus1|frame_gen_testbus2|enc64b66b_testbus|txsm_testbus|tx_cp_bond_testbus|gearbox_red_testbus|scramble_testbus|blank_testbus|tx_fifo_testbus1|tx_fifo_testbus2
		parameter hssi_10g_tx_pcs_txfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_tx_pcs_txfifo_full = "full_default", // full_default
		parameter hssi_10g_tx_pcs_txfifo_mode = "phase_comp", // register_mode|interlaken_generic|basic_generic|phase_comp
		parameter hssi_10g_tx_pcs_txfifo_pempty = 4'b10,
		parameter hssi_10g_tx_pcs_txfifo_pfull = 4'b1011,
		parameter hssi_10g_tx_pcs_wr_clk_sel = "wr_tx_pma_clk", // wr_tx_pld_clk|wr_tx_pma_clk|wr_refclk_dig
		parameter hssi_10g_tx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_8g_rx_pcs
		parameter hssi_8g_rx_pcs_auto_error_replacement = "dis_err_replace", // dis_err_replace|en_err_replace
		parameter hssi_8g_rx_pcs_auto_speed_nego = "dis_asn", // dis_asn|en_asn_g2_freq_scal
		parameter hssi_8g_rx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_rx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_rx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_rx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_rx_pcs_byte_deserializer = "dis_bds", // dis_bds|en_bds_by_2|en_bds_by_4|en_bds_by_2_det
		parameter hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask = "dis_rxvalid_mask", // dis_rxvalid_mask|en_rxvalid_mask
		parameter hssi_8g_rx_pcs_clkcmp_pattern_n = 20'b0,
		parameter hssi_8g_rx_pcs_clkcmp_pattern_p = 20'b0,
		parameter hssi_8g_rx_pcs_clock_gate_bds_dec_asn = "dis_bds_dec_asn_clk_gating", // dis_bds_dec_asn_clk_gating|en_bds_dec_asn_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_cdr_eidle = "dis_cdr_eidle_clk_gating", // dis_cdr_eidle_clk_gating|en_cdr_eidle_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk = "dis_dw_pc_wrclk_gating", // dis_dw_pc_wrclk_gating|en_dw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_rd = "dis_dw_rm_rdclk_gating", // dis_dw_rm_rdclk_gating|en_dw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_wr = "dis_dw_rm_wrclk_gating", // dis_dw_rm_wrclk_gating|en_dw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_wa = "dis_dw_wa_clk_gating", // dis_dw_wa_clk_gating|en_dw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_pc_rdclk = "dis_pc_rdclk_gating", // dis_pc_rdclk_gating|en_pc_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk = "dis_sw_pc_wrclk_gating", // dis_sw_pc_wrclk_gating|en_sw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_rd = "dis_sw_rm_rdclk_gating", // dis_sw_rm_rdclk_gating|en_sw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_wr = "dis_sw_rm_wrclk_gating", // dis_sw_rm_wrclk_gating|en_sw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_wa = "dis_sw_wa_clk_gating", // dis_sw_wa_clk_gating|en_sw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_observation_in_pld_core = "internal_sw_wa_clk", // internal_sw_wa_clk|internal_dw_wa_clk|internal_cdr_eidle_clk|internal_sm_rm_wr_clk|internal_dw_rm_wr_clk|internal_clk_2_b|internal_sw_rm_rd_clk|internal_dw_rm_rd_clk|internal_sw_rx_wr_clk|internal_dw_rx_wr_clk|internal_rx_rd_clk|internal_rx_pma_clk_gen3|internal_rx_rcvd_clk_gen3
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_rx_pcs_eidle_entry_eios = "dis_eidle_eios", // dis_eidle_eios|en_eidle_eios
		parameter hssi_8g_rx_pcs_eidle_entry_iei = "dis_eidle_iei", // dis_eidle_iei|en_eidle_iei
		parameter hssi_8g_rx_pcs_eidle_entry_sd = "dis_eidle_sd", // dis_eidle_sd|en_eidle_sd
		parameter hssi_8g_rx_pcs_eightb_tenb_decoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_rx_pcs_err_flags_sel = "err_flags_wa", // err_flags_wa|err_flags_8b10b
		parameter hssi_8g_rx_pcs_fixed_pat_det = "dis_fixed_patdet", // dis_fixed_patdet|en_fixed_patdet
		parameter hssi_8g_rx_pcs_fixed_pat_num = 4'b1111,
		parameter hssi_8g_rx_pcs_force_signal_detect = "en_force_signal_detect", // en_force_signal_detect|dis_force_signal_detect
		parameter hssi_8g_rx_pcs_gen3_clk_en = "disable_clk", // disable_clk|enable_clk
		parameter hssi_8g_rx_pcs_gen3_rx_clk_sel = "rcvd_clk", // en_dig_clk1_8g|rcvd_clk
		parameter hssi_8g_rx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // en_dig_clk2_8g|tx_pma_clk
		parameter hssi_8g_rx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_rx_pcs_ibm_invalid_code = "dis_ibm_invalid_code", // dis_ibm_invalid_code|en_ibm_invalid_code
		parameter hssi_8g_rx_pcs_invalid_code_flag_only = "dis_invalid_code_only", // dis_invalid_code_only|en_invalid_code_only
		parameter hssi_8g_rx_pcs_pad_or_edb_error_replace = "replace_edb", // replace_edb|replace_edb_dynamic|replace_pad
		parameter hssi_8g_rx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_rx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_rx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_rx_pcs_pipe_if_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_8g_rx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_rx_pcs_polinv_8b10b_dec = "dis_polinv_8b10b_dec", // dis_polinv_8b10b_dec|en_polinv_8b10b_dec
		parameter hssi_8g_rx_pcs_prot_mode = "gige", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic_rm_enable|basic_rm_disable|disabled_prot_mode
		parameter hssi_8g_rx_pcs_rate_match = "dis_rm", // dis_rm|gige_rm|pipe_rm|pipe_rm_0ppm|sw_basic_rm|dw_basic_rm
		parameter hssi_8g_rx_pcs_rate_match_del_thres = "dis_rm_del_thres", // dis_rm_del_thres|gige_rm_del_thres|pipe_rm_del_thres|pipe_rm_0ppm_del_thres|sw_basic_rm_del_thres|dw_basic_rm_del_thres
		parameter hssi_8g_rx_pcs_rate_match_empty_thres = "dis_rm_empty_thres", // dis_rm_empty_thres|gige_rm_empty_thres|pipe_rm_empty_thres|pipe_rm_0ppm_empty_thres|sw_basic_rm_empty_thres|dw_basic_rm_empty_thres
		parameter hssi_8g_rx_pcs_rate_match_full_thres = "dis_rm_full_thres", // dis_rm_full_thres|gige_rm_full_thres|pipe_rm_full_thres|pipe_rm_0ppm_full_thres|sw_basic_rm_full_thres|dw_basic_rm_full_thres
		parameter hssi_8g_rx_pcs_rate_match_ins_thres = "dis_rm_ins_thres", // dis_rm_ins_thres|gige_rm_ins_thres|pipe_rm_ins_thres|pipe_rm_0ppm_ins_thres|sw_basic_rm_ins_thres|dw_basic_rm_ins_thres
		parameter hssi_8g_rx_pcs_rate_match_start_thres = "dis_rm_start_thres", // dis_rm_start_thres|gige_rm_start_thres|pipe_rm_start_thres|pipe_rm_0ppm_start_thres|sw_basic_rm_start_thres|dw_basic_rm_start_thres
		parameter hssi_8g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_rx_pcs_rx_clk2 = "rcvd_clk_clk2", // rcvd_clk_clk2|tx_pma_clock_clk2|refclk_dig2_clk2
		parameter hssi_8g_rx_pcs_rx_clk_free_running = "en_rx_clk_free_run", // dis_rx_clk_free_run|en_rx_clk_free_run
		parameter hssi_8g_rx_pcs_rx_pcs_urst = "en_rx_pcs_urst", // dis_rx_pcs_urst|en_rx_pcs_urst
		parameter hssi_8g_rx_pcs_rx_rcvd_clk = "rcvd_clk_rcvd_clk", // rcvd_clk_rcvd_clk|tx_pma_clock_rcvd_clk
		parameter hssi_8g_rx_pcs_rx_rd_clk = "pld_rx_clk", // pld_rx_clk|rx_clk
		parameter hssi_8g_rx_pcs_rx_refclk = "dis_refclk_sel", // dis_refclk_sel|en_refclk_sel
		parameter hssi_8g_rx_pcs_rx_wr_clk = "rx_clk2_div_1_2_4", // rx_clk2_div_1_2_4|txfifo_rd_clk
		parameter hssi_8g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_rx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_rx_pcs_sync_sm_idle_eios = "dis_syncsm_idle", // dis_syncsm_idle|en_syncsm_idle
		parameter hssi_8g_rx_pcs_test_bus_sel = "tx_testbus", // tx_testbus|tx_ctrl_plane_testbus|wa_testbus|rm_testbus|rx_ctrl_testbus|pcie_ctrl_testbus|rx_ctrl_plane_testbus
		parameter hssi_8g_rx_pcs_tx_rx_parallel_loopback = "dis_plpbk", // dis_plpbk|en_plpbk
		parameter hssi_8g_rx_pcs_wa_boundary_lock_ctrl = "bit_slip", // bit_slip|sync_sm|deterministic_latency|auto_align_pld_ctrl
		parameter hssi_8g_rx_pcs_wa_clk_slip_spacing = 10'b10000,
		parameter hssi_8g_rx_pcs_wa_det_latency_sync_status_beh = "assert_sync_status_non_imm", // assert_sync_status_imm|assert_sync_status_non_imm|dont_care_assert_sync
		parameter hssi_8g_rx_pcs_wa_disp_err_flag = "dis_disp_err_flag", // dis_disp_err_flag|en_disp_err_flag
		parameter hssi_8g_rx_pcs_wa_kchar = "dis_kchar", // dis_kchar|en_kchar
		parameter hssi_8g_rx_pcs_wa_pd = "wa_pd_10", // wa_pd_7|wa_pd_10|wa_pd_20|wa_pd_40|wa_pd_8_sw|wa_pd_8_dw|wa_pd_16_sw|wa_pd_16_dw|wa_pd_32
		parameter hssi_8g_rx_pcs_wa_pd_data = 40'b0,
		parameter hssi_8g_rx_pcs_wa_pd_polarity = "dis_pd_both_pol", // dis_pd_both_pol|en_pd_both_pol|dont_care_both_pol
		parameter hssi_8g_rx_pcs_wa_pld_controlled = "dis_pld_ctrl", // dis_pld_ctrl|pld_ctrl_sw|rising_edge_sensitive_dw|level_sensitive_dw
		parameter hssi_8g_rx_pcs_wa_renumber_data = 6'b0,
		parameter hssi_8g_rx_pcs_wa_rgnumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rknumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rosnumber_data = 2'b0,
		parameter hssi_8g_rx_pcs_wa_rvnumber_data = 13'b0,
		parameter hssi_8g_rx_pcs_wa_sync_sm_ctrl = "gige_sync_sm", // gige_sync_sm|pipe_sync_sm|sw_basic_sync_sm|dw_basic_sync_sm|fibre_channel_sync_sm
		parameter hssi_8g_rx_pcs_wait_cnt = 12'b0,
		
		// parameters for twentynm_hssi_8g_tx_pcs
		parameter hssi_8g_tx_pcs_auto_speed_nego_gen2 = "dis_asn_g2", // dis_asn_g2|en_asn_g2_freq_scal
		parameter hssi_8g_tx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_tx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_tx_pcs_byte_serializer = "dis_bs", // dis_bs|en_bs_by_2|en_bs_by_4
		parameter hssi_8g_tx_pcs_clock_gate_bs_enc = "dis_bs_enc_clk_gating", // dis_bs_enc_clk_gating|en_bs_enc_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_dw_fifowr = "dis_dw_fifowr_clk_gating", // dis_dw_fifowr_clk_gating|en_dw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_fiford = "dis_fiford_clk_gating", // dis_fiford_clk_gating|en_fiford_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_sw_fifowr = "dis_sw_fifowr_clk_gating", // dis_sw_fifowr_clk_gating|en_sw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_observation_in_pld_core = "internal_refclk_b", // internal_refclk_b|internal_fifo_rd_clk|internal_sw_fifo_wr_clk|internal_dw_fifo_wr_clk|internal_tx_clk_out_gen3|internal_pipe_tx_clk_out_gen3
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_tx_pcs_data_selection_8b10b_encoder_input = "normal_data_path", // normal_data_path|gige_idle_conversion
		parameter hssi_8g_tx_pcs_dynamic_clk_switch = "dis_dyn_clk_switch", // dis_dyn_clk_switch|en_dyn_clk_switch
		parameter hssi_8g_tx_pcs_eightb_tenb_disp_ctrl = "dis_disp_ctrl", // dis_disp_ctrl|en_disp_ctrl|en_ib_disp_ctrl
		parameter hssi_8g_tx_pcs_eightb_tenb_encoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_tx_pcs_force_echar = "dis_force_echar", // dis_force_echar|en_force_echar
		parameter hssi_8g_tx_pcs_force_kchar = "dis_force_kchar", // dis_force_kchar|en_force_kchar
		parameter hssi_8g_tx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // dis_tx_clk|tx_pma_clk
		parameter hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel = "func_clk", // dis_tx_pipe_clk|func_clk
		parameter hssi_8g_tx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_tx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_tx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_tx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_tx_pcs_phfifo_write_clk_sel = "pld_tx_clk", // pld_tx_clk|tx_clk
		parameter hssi_8g_tx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_tx_pcs_prot_mode = "basic", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic|disabled_prot_mode
		parameter hssi_8g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_tx_pcs_refclk_b_clk_sel = "tx_pma_clock", // tx_pma_clock|refclk_dig
		parameter hssi_8g_tx_pcs_revloop_back_rm = "dis_rev_loopback_rx_rm", // dis_rev_loopback_rx_rm|en_rev_loopback_rx_rm
		parameter hssi_8g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_tx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_tx_pcs_tx_bitslip = "dis_tx_bitslip", // dis_tx_bitslip|en_tx_bitslip
		parameter hssi_8g_tx_pcs_tx_compliance_controlled_disparity = "dis_txcompliance", // dis_txcompliance|en_txcompliance_pipe2p0|en_txcompliance_pipe3p0
		parameter hssi_8g_tx_pcs_tx_fast_pld_reg = "dis_tx_fast_pld_reg", // dis_tx_fast_pld_reg|en_tx_fast_pld_reg
		parameter hssi_8g_tx_pcs_txclk_freerun = "dis_freerun_tx", // dis_freerun_tx|en_freerun_tx
		parameter hssi_8g_tx_pcs_txpcs_urst = "en_txpcs_urst", // dis_txpcs_urst|en_txpcs_urst
		
		// parameters for twentynm_hssi_common_pcs_pma_interface
		parameter hssi_common_pcs_pma_interface_asn_clk_enable = "false", // false|true
		parameter hssi_common_pcs_pma_interface_asn_enable = "dis_asn", // dis_asn|en_asn
		parameter hssi_common_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|pcie_gen3
		parameter hssi_common_pcs_pma_interface_bypass_early_eios = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pcie_switch = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_ltr = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_sw_done = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_ppm_lock = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_txdetectrx = "false", // false|true
		parameter hssi_common_pcs_pma_interface_cdr_control = "en_cdr_ctrl", // dis_cdr_ctrl|en_cdr_ctrl
		parameter hssi_common_pcs_pma_interface_cid_enable = "en_cid_mode", // dis_cid_mode|en_cid_mode
		parameter hssi_common_pcs_pma_interface_cp_cons_sel = "cp_cons_default", // cp_cons_master|cp_cons_slave_abv|cp_cons_slave_blw|cp_cons_default
		parameter hssi_common_pcs_pma_interface_cp_dwn_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_cp_up_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_blw|ctrl_slave_abv
		parameter hssi_common_pcs_pma_interface_data_mask_count = 16'b100111000100,
		parameter hssi_common_pcs_pma_interface_data_mask_count_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_dft_observation_clock_selection = "dft_clk_obsrv_tx0", // dft_clk_obsrv_tx0|dft_clk_obsrv_tx1|dft_clk_obsrv_tx2|dft_clk_obsrv_tx3|dft_clk_obsrv_tx4|dft_clk_obsrv_rx|dft_clk_obsrv_hclk|dft_clk_obsrv_fref|dft_clk_obsrv_clklow|dft_clk_obsrv_asn0|dft_clk_obsrv_asn1
		parameter hssi_common_pcs_pma_interface_early_eios_counter = 8'b110010,
		parameter hssi_common_pcs_pma_interface_force_freqdet = "force_freqdet_dis", // force_freqdet_dis|force1_freqdet_en|force0_freqdet_en
		parameter hssi_common_pcs_pma_interface_free_run_clk_enable = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ignore_sigdet_g23 = "false", // false|true
		parameter hssi_common_pcs_pma_interface_pc_en_counter = 7'b110111,
		parameter hssi_common_pcs_pma_interface_pc_rst_counter = 5'b10111,
		parameter hssi_common_pcs_pma_interface_pcie_hip_mode = "hip_disable", // hip_enable|hip_disable
		parameter hssi_common_pcs_pma_interface_ph_fifo_reg_mode = "phfifo_reg_mode_dis", // phfifo_reg_mode_dis|phfifo_reg_mode_en
		parameter hssi_common_pcs_pma_interface_phfifo_flush_wait = 6'b100100,
		parameter hssi_common_pcs_pma_interface_pipe_if_g3pcs = "pipe_if_8gpcs", // pipe_if_g3pcs|pipe_if_8gpcs
		parameter hssi_common_pcs_pma_interface_pma_done_counter = 18'b101010101110011000,
		parameter hssi_common_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_common_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_common_pcs_pma_interface_ppm_cnt_rst = "ppm_cnt_rst_dis", // ppm_cnt_rst_dis|ppm_cnt_rst_en
		parameter hssi_common_pcs_pma_interface_ppm_deassert_early = "deassert_early_dis", // deassert_early_dis|deassert_early_en
		parameter hssi_common_pcs_pma_interface_ppm_det_buckets = "ppm_100_bucket", // disable_prot|ppm_300_bucket|ppm_100_bucket|ppm_300_100_bucket
		parameter hssi_common_pcs_pma_interface_ppm_gen1_2_cnt = "cnt_32k", // cnt_32k|cnt_64k
		parameter hssi_common_pcs_pma_interface_ppm_post_eidle_delay = "cnt_200_cycles", // cnt_200_cycles|cnt_400_cycles
		parameter hssi_common_pcs_pma_interface_ppmsel = "ppmsel_300", // ppmsel_disable|ppmsel_5000|ppmsel_2500|ppmsel_1000|ppmsel_500|ppmsel_300|ppmsel_250|ppmsel_200|ppmsel_125|ppmsel_100|ppmsel_62p5|ppm_other
		parameter hssi_common_pcs_pma_interface_prot_mode = "disable_prot_mode", // disable_prot_mode|pipe_g12|pipe_g3|other_protocols
		parameter hssi_common_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_common_pcs_pma_interface_rxvalid_mask = "rxvalid_mask_en", // rxvalid_mask_dis|rxvalid_mask_en
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter = 12'b100111000100,
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_sim_mode = "disable", // disable|enable
		parameter hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en = "true", // false|true
		parameter hssi_common_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_common_pcs_pma_interface_testout_sel = "ppm_det_test", // ppm_det_test|asn_test|pma_pll_test|rxpmaif_test|prbs_gen_test|prbs_ver_test|uhsif_1_test|uhsif_2_test|uhsif_3_test
		parameter hssi_common_pcs_pma_interface_wait_clk_on_off_timer = 4'b100,
		parameter hssi_common_pcs_pma_interface_wait_pipe_synchronizing = 5'b10111,
		parameter hssi_common_pcs_pma_interface_wait_send_syncp_fbkp = 11'b11111010,
		
		// parameters for twentynm_hssi_common_pld_pcs_interface
		parameter hssi_common_pld_pcs_interface_dft_clk_out_en = "dft_clk_out_disable", // dft_clk_out_disable|dft_clk_out_enable
		parameter hssi_common_pld_pcs_interface_dft_clk_out_sel = "teng_rx_dft_clk", // teng_rx_dft_clk|teng_tx_dft_clk|eightg_rx_dft_clk|eightg_tx_dft_clk|pmaif_dft_clk
		parameter hssi_common_pld_pcs_interface_hrdrstctrl_en = "hrst_dis", // hrst_dis|hrst_en
		parameter hssi_common_pld_pcs_interface_pcs_testbus_block_sel = "eightg", // eightg|g3pcs|teng|krfec|pma_if
		parameter hssi_common_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_fifo_rx_pcs
		parameter hssi_fifo_rx_pcs_double_read_mode = "double_read_dis", // double_read_en|double_read_dis
		parameter hssi_fifo_rx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_fifo_tx_pcs
		parameter hssi_fifo_tx_pcs_double_write_mode = "double_write_dis", // double_write_en|double_write_dis
		parameter hssi_fifo_tx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_gen3_rx_pcs
		parameter hssi_gen3_rx_pcs_block_sync = "enable_block_sync", // bypass_block_sync|enable_block_sync
		parameter hssi_gen3_rx_pcs_block_sync_sm = "enable_blk_sync_sm", // disable_blk_sync_sm|enable_blk_sync_sm
		parameter hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn = "enable", // disable|enable
		parameter hssi_gen3_rx_pcs_lpbk_force = "lpbk_frce_dis", // lpbk_frce_dis|lpbk_frce_en
		parameter hssi_gen3_rx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_rx_pcs_rate_match_fifo = "enable_rm_fifo_600ppm", // bypass_rm_fifo|enable_rm_fifo_600ppm|enable_rm_fifo_0ppm
		parameter hssi_gen3_rx_pcs_rate_match_fifo_latency = "regular_latency", // regular_latency|low_latency
		parameter hssi_gen3_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_gen3_rx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_b4gb_par_lpbk = "b4gb_par_lpbk_dis", // b4gb_par_lpbk_dis|b4gb_par_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_force_balign = "en_force_balign", // en_force_balign|dis_force_balign
		parameter hssi_gen3_rx_pcs_rx_ins_del_one_skip = "ins_del_one_skip_en", // ins_del_one_skip_dis|ins_del_one_skip_en
		parameter hssi_gen3_rx_pcs_rx_num_fixed_pat = 4'b1000,
		parameter hssi_gen3_rx_pcs_rx_test_out_sel = "rx_test_out0", // rx_test_out0|rx_test_out1
		parameter hssi_gen3_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_gen3_tx_pcs
		parameter hssi_gen3_tx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_tx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_gen3_tx_pcs_tx_bitslip = 5'b0,
		parameter hssi_gen3_tx_pcs_tx_gbox_byp = "bypass_gbox", // bypass_gbox|enable_gbox
		
		// parameters for twentynm_hssi_krfec_rx_pcs
		parameter hssi_krfec_rx_pcs_blksync_cor_en = "detect", // detect|correct
		parameter hssi_krfec_rx_pcs_bypass_gb = "bypass_dis", // bypass_dis|bypass_en
		parameter hssi_krfec_rx_pcs_clr_ctrl = "both_enabled", // both_enabled|corr_cnt_only|uncorr_cnt_only
		parameter hssi_krfec_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_rx_pcs_dv_start = "with_blklock", // with_blksync|with_blklock
		parameter hssi_krfec_rx_pcs_err_mark_type = "err_mark_10g", // err_mark_10g|err_mark_40g
		parameter hssi_krfec_rx_pcs_error_marking_en = "err_mark_dis", // err_mark_dis|err_mark_en
		parameter hssi_krfec_rx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_krfec_rx_pcs_parity_invalid_enum = 8'b1000,
		parameter hssi_krfec_rx_pcs_parity_valid_num = 4'b100,
		parameter hssi_krfec_rx_pcs_pipeln_blksync = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_descrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errcorrect = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_ind = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_lfsr = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_loc = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_pat = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_gearbox = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_syndrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_trans_dec = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_rx_pcs_receive_order = "receive_lsb", // receive_lsb|receive_msb
		parameter hssi_krfec_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_krfec_rx_pcs_rx_testbus_sel = "overall", // overall|fast_search|fast_search_cntrs|blksync|blksync_cntrs|decoder_master_sm|decoder_master_sm_cntrs|syndrm_sm|syndrm1|syndrm2|errtrap_sm|errtrap_ind1|errtrap_ind2|errtrap_ind3|errtrap_ind4|errtrap_ind5|errtrap_loc|errtrap_pat1|errtrap_pat2|errtrap_pat3|errtrap_pat4|decoder_rd_sm|gb_and_trans
		parameter hssi_krfec_rx_pcs_signal_ok_en = "sig_ok_dis", // sig_ok_dis|sig_ok_en
		parameter hssi_krfec_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_krfec_tx_pcs
		parameter hssi_krfec_tx_pcs_burst_err = "burst_err_dis", // burst_err_dis|burst_err_en
		parameter hssi_krfec_tx_pcs_burst_err_len = "burst_err_len1", // burst_err_len1|burst_err_len2|burst_err_len3|burst_err_len4|burst_err_len5|burst_err_len6|burst_err_len7|burst_err_len8|burst_err_len9|burst_err_len10|burst_err_len11|burst_err_len12|burst_err_len13|burst_err_len14|burst_err_len15|burst_err_len16
		parameter hssi_krfec_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_tx_pcs_enc_frame_query = "enc_query_dis", // enc_query_dis|enc_query_en
		parameter hssi_krfec_tx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_encoder = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_scrambler = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_krfec_tx_pcs_transcode_err = "trans_err_dis", // trans_err_dis|trans_err_en
		parameter hssi_krfec_tx_pcs_transmit_order = "transmit_lsb", // transmit_lsb|transmit_msb
		parameter hssi_krfec_tx_pcs_tx_testbus_sel = "overall", // overall|encoder1|encoder2|scramble1|scramble2|scramble3|gearbox
		
		// parameters for twentynm_hssi_pipe_gen1_2
		parameter hssi_pipe_gen1_2_elec_idle_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_error_replace_pad = "replace_edb", // replace_edb|replace_pad
		parameter hssi_pipe_gen1_2_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_pipe_gen1_2_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen1_2_phystatus_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_phystatus_rst_toggle = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen1_2_pipe_byte_de_serializer_en = "dont_care_bds", // dis_bds|en_bds_by_2|dont_care_bds
		parameter hssi_pipe_gen1_2_prot_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|basic|disabled_prot_mode
		parameter hssi_pipe_gen1_2_reconfig_settings = "{}", // 
		parameter hssi_pipe_gen1_2_rx_pipe_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_pipe_gen1_2_rxdetect_bypass = "dis_rxdetect_bypass", // dis_rxdetect_bypass|en_rxdetect_bypass
		parameter hssi_pipe_gen1_2_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen1_2_tx_pipe_enable = "dis_pipe_tx", // dis_pipe_tx|en_pipe_tx|en_pipe3_tx
		parameter hssi_pipe_gen1_2_txswing = "dis_txswing", // dis_txswing|en_txswing
		
		// parameters for twentynm_hssi_pipe_gen3
		parameter hssi_pipe_gen3_bypass_rx_detection_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_rx_preset = 3'b0,
		parameter hssi_pipe_gen3_bypass_rx_preset_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_tx_coefficent = 18'b0,
		parameter hssi_pipe_gen3_bypass_tx_coefficent_enable = "false", // false|true
		parameter hssi_pipe_gen3_elecidle_delay_g3 = 3'b110,
		parameter hssi_pipe_gen3_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen3_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|disable_pcs
		parameter hssi_pipe_gen3_phy_status_delay_g12 = 3'b101,
		parameter hssi_pipe_gen3_phy_status_delay_g3 = 3'b101,
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g12 = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g3 = "dis_phystatus_rst_toggle_g3", // dis_phystatus_rst_toggle_g3|en_phystatus_rst_toggle_g3
		parameter hssi_pipe_gen3_rate_match_pad_insertion = "dis_rm_fifo_pad_ins", // dis_rm_fifo_pad_ins|en_rm_fifo_pad_ins
		parameter hssi_pipe_gen3_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen3_test_out_sel = "disable_test_out", // tx_test_out|rx_test_out|pipe_test_out1|pipe_test_out2|pipe_test_out3|pipe_ctrl_test_out|disable_test_out
		
		// parameters for twentynm_hssi_rx_pcs_pma_interface
		parameter hssi_rx_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|ten_g_pcs|direct_pld
		parameter hssi_rx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pcs_pma_interface_clkslip_sel = "pld", // pld|slip_eight_g_pcs
		parameter hssi_rx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pcs_pma_interface_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_rx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_rx_pcs_pma_interface_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_rx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_rx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_rx_pcs_pma_interface_prbs_ver = "prbs_off", // prbs_off|prbs_31|prbs_15|prbs_23|prbs_9|prbs_7
		parameter hssi_rx_pcs_pma_interface_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion = "rx_dyn_polinv_dis", // rx_dyn_polinv_dis|rx_dyn_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_lpbk_en = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok = "unforce_sig_ok", // unforce_sig_ok|force_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mask = "prbsmask128", // prbsmask128|prbsmask256|prbsmask512|prbsmask1024
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mode = "teng_mode", // teng_mode|eightg_mode
		parameter hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel = "sel_sig_det", // sel_sig_det|sel_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_static_polarity_inversion = "rx_stat_polinv_dis", // rx_stat_polinv_dis|rx_stat_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en = "uhsif_lpbk_dis", // uhsif_lpbk_dis|uhsif_lpbk_en
		parameter hssi_rx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_rx_pld_pcs_interface
		parameter hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx = "enable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx = "pma_64b_rx", // pma_32b_rx|pma_40b_rx|pma_64b_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_baser_mode_rx|interlaken_mode_rx|sfis_mode_rx|teng_sdi_mode_rx|basic_mode_rx|test_prp_mode_rx|test_prp_krfec_mode_rx|teng_1588_mode_rx|teng_baser_krfec_mode_rx|teng_1588_krfec_mode_rx|basic_krfec_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx = "disabled_prot_mode_rx", // pipe_g1_rx|pipe_g2_rx|pipe_g3_rx|cpri_rx|cpri_rx_tx_rx|gige_rx|gige_1588_rx|basic_rm_enable_rx|basic_rm_disable_rx|disabled_prot_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcie_g1_capable_rx|pcie_g2_capable_rx|pcie_g3_capable_rx|gige_rx|teng_baser_rx|teng_basekr_krfec_rx|fortyg_basekr_krfec_rx|cpri_8b10b_rx|interlaken_rx|sfis_rx|teng_sdi_rx|gige_1588_rx|teng_1588_baser_rx|teng_1588_basekr_krfec_rx|basic_8gpcs_rm_enable_rx|basic_8gpcs_rm_disable_rx|basic_10gpcs_rx|basic_10gpcs_krfec_rx|pcs_direct_rx|prp_rx|prp_krfec_rx|prbs_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx = "teng_mode_rx", // teng_mode_rx|non_teng_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_basekr_mode_rx|fortyg_basekr_mode_rx|teng_1588_basekr_mode_rx|basic_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|eightg_and_g3_pld_fifo_mode_rx|eightg_and_g3_reg_mode_rx|eightg_and_g3_reg_mode_hip_rx|teng_pld_fifo_mode_rx|teng_reg_mode_rx|teng_and_krfec_pld_fifo_mode_rx|teng_and_krfec_reg_mode_rx|pcs_direct_reg_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_block_sel = "pcs_direct", // eightg|teng|pcs_direct
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_rx_clk|pma_rx_clk_user
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_sel = "pld_rx_clk", // pld_rx_clk|pcs_rx_clk
		parameter hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en = "hip_rx_enable", // hip_rx_enable|hip_rx_disable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_rx_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_tx_pcs_pma_interface
		parameter hssi_tx_pcs_pma_interface_bypass_pma_txelecidle = "false", // false|true
		parameter hssi_tx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pcs_pma_interface_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx = "other_prot_mode", // pipe_g12|pipe_g3|other_prot_mode
		parameter hssi_tx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_tx_pcs_pma_interface_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_tx_pcs_pma_interface_pmagate_en = "pmagate_dis", // pmagate_dis|pmagate_en
		parameter hssi_tx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_tx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_tx_pcs_pma_interface_prbs_gen_pat = "prbs_gen_dis", // prbs_gen_dis|prbs_31|prbs_23|prbs_15|prbs_9|prbs_7
		parameter hssi_tx_pcs_pma_interface_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_tx_pcs_pma_interface_sq_wave_num = "sq_wave_4", // sq_wave_1|sq_wave_4|sq_wave_8|sq_wave_6|sq_wave_default
		parameter hssi_tx_pcs_pma_interface_sqwgen_clken = "sqwgen_clk_dis", // sqwgen_clk_dis|sqwgen_clk_en
		parameter hssi_tx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion = "tx_dyn_polinv_dis", // tx_dyn_polinv_dis|tx_dyn_polinv_en
		parameter hssi_tx_pcs_pma_interface_tx_pma_data_sel = "pld_dir", // pld_dir|pcie_gen3|eight_g_pcs|ten_g_pcs|prbs_pat|sq_wave_pat|block_sel_default|registered_uhsif_dat|directed_uhsif_dat
		parameter hssi_tx_pcs_pma_interface_tx_static_polarity_inversion = "tx_stat_polinv_dis", // tx_stat_polinv_dis|tx_stat_polinv_en
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock = "uhsif_filt_stepsz_b4lock_4", // uhsif_filt_stepsz_b4lock_2|uhsif_filt_stepsz_b4lock_4|uhsif_filt_stepsz_b4lock_6|uhsif_filt_stepsz_b4lock_8
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value = 4'b1011,
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock = "uhsif_filt_cntthr_b4lock_16", // uhsif_filt_cntthr_b4lock_8|uhsif_filt_cntthr_b4lock_16|uhsif_filt_cntthr_b4lock_24|uhsif_filt_cntthr_b4lock_32
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period = "uhsif_dcn_test_period_4", // uhsif_dcn_test_period_4|uhsif_dcn_test_period_8|uhsif_dcn_test_period_12|uhsif_dcn_test_period_16
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable = "uhsif_dcn_test_mode_disable", // uhsif_dcn_test_mode_enable|uhsif_dcn_test_mode_disable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh = "uhsif_dzt_cnt_thr_4", // uhsif_dzt_cnt_thr_2|uhsif_dzt_cnt_thr_4|uhsif_dzt_cnt_thr_6|uhsif_dzt_cnt_thr_8
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable = "uhsif_dzt_enable", // uhsif_dzt_disable|uhsif_dzt_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window = "uhsif_dzt_obr_win_32", // uhsif_dzt_obr_win_16|uhsif_dzt_obr_win_32|uhsif_dzt_obr_win_48|uhsif_dzt_obr_win_64
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size = "uhsif_dzt_skipsz_8", // uhsif_dzt_skipsz_4|uhsif_dzt_skipsz_8|uhsif_dzt_skipsz_12|uhsif_dzt_skipsz_16
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel = "uhsif_index_internal", // uhsif_index_internal|uhsif_index_cram
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin = "uhsif_dcn_margin_4", // uhsif_dcn_margin_2|uhsif_dcn_margin_3|uhsif_dcn_margin_4|uhsif_dcn_margin_5
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value = 8'b10000000,
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control = "uhsif_dft_dz_det_val_0", // uhsif_dft_dz_det_val_0|uhsif_dft_dz_det_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control = "uhsif_dft_up_val_0", // uhsif_dft_up_val_0|uhsif_dft_up_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_enable = "uhsif_disable", // uhsif_disable|uhsif_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock = "uhsif_lkd_segsz_aflock_2048", // uhsif_lkd_segsz_aflock_512|uhsif_lkd_segsz_aflock_1024|uhsif_lkd_segsz_aflock_2048|uhsif_lkd_segsz_aflock_4096
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock = "uhsif_lkd_segsz_b4lock_32", // uhsif_lkd_segsz_b4lock_16|uhsif_lkd_segsz_b4lock_32|uhsif_lkd_segsz_b4lock_64|uhsif_lkd_segsz_b4lock_128
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value = 4'b11,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value = 4'b11,
		
		// parameters for twentynm_hssi_tx_pld_pcs_interface
		parameter hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx = "enable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx = "pma_64b_tx", // pma_32b_tx|pma_40b_tx|pma_64b_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_baser_mode_tx|interlaken_mode_tx|sfis_mode_tx|teng_sdi_mode_tx|basic_mode_tx|test_prp_mode_tx|test_prp_krfec_mode_tx|teng_1588_mode_tx|teng_baser_krfec_mode_tx|teng_1588_krfec_mode_tx|basic_krfec_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx = "disabled_prot_mode_tx", // pipe_g1_tx|pipe_g2_tx|pipe_g3_tx|cpri_tx|cpri_rx_tx_tx|gige_tx|gige_1588_tx|basic_tx|disabled_prot_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcie_g1_capable_tx|pcie_g2_capable_tx|pcie_g3_capable_tx|gige_tx|teng_baser_tx|teng_basekr_krfec_tx|fortyg_basekr_krfec_tx|cpri_8b10b_tx|interlaken_tx|sfis_tx|teng_sdi_tx|gige_1588_tx|teng_1588_baser_tx|teng_1588_basekr_krfec_tx|basic_8gpcs_tx|basic_10gpcs_tx|basic_10gpcs_krfec_tx|pcs_direct_tx|uhsif_tx|prp_tx|prp_krfec_tx|prbs_tx|sqwave_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx = "teng_mode_tx", // teng_mode_tx|non_teng_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_basekr_mode_tx|fortyg_basekr_mode_tx|teng_1588_basekr_mode_tx|basic_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|eightg_and_g3_pld_fifo_mode_tx|eightg_and_g3_reg_mode_tx|eightg_and_g3_reg_mode_hip_tx|eightg_and_g3_fastreg_mode_tx|teng_pld_fifo_mode_tx|teng_reg_mode_tx|teng_fastreg_mode_tx|teng_and_krfec_pld_fifo_mode_tx|teng_and_krfec_reg_mode_tx|teng_and_krfec_fastreg_mode_tx|pcs_direct_fastreg_mode_tx|uhsif_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_tx_clk|pma_tx_clk_user
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_source = "teng", // eightg|teng|pma_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_data_source = "hip_disable", // hip_disable|hip_enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en = "delay1_clk_disable", // delay1_clk_enable|delay1_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel = "pld_tx_clk", // pld_tx_clk|pcs_tx_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl = "delay1_path0", // delay1_path0|delay1_path1|delay1_path2|delay1_path3|delay1_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel = "one_ff_delay", // one_ff_delay|two_ff_delay
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en = "delay2_clk_disable", // delay2_clk_enable|delay2_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl = "delay2_path0", // delay2_path0|delay2_path1|delay2_path2|delay2_path3|delay2_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_tx_pld_pcs_interface_reconfig_settings = "{}" // 
	//PARAM_LIST_END
	)
	(
	//PORT_LIST_START
		input wire	[8:0]	in_avmmaddress,
		input wire		in_avmmclk,
		input wire		in_avmmread,
		input wire		in_avmmrstn,
		input wire		in_avmmwrite,
		input wire	[7:0]	in_avmmwritedata,
		input wire	[4:0]	in_bond_pcs10g_in_bot,
		input wire	[4:0]	in_bond_pcs10g_in_top,
		input wire	[12:0]	in_bond_pcs8g_in_bot,
		input wire	[12:0]	in_bond_pcs8g_in_top,
		input wire	[11:0]	in_bond_pmaif_in_bot,
		input wire	[11:0]	in_bond_pmaif_in_top,
		input wire	[63:0]	in_hip_tx_data,
		input wire		in_iocsr_clk,
		input wire	[5:0]	in_iocsr_config,
		input wire		in_iocsr_rdy,
		input wire		in_iocsr_rdy_dly,
		input wire		in_pld_10g_krfec_rx_clr_errblk_cnt,
		input wire		in_pld_10g_krfec_rx_pld_rst_n,
		input wire		in_pld_10g_krfec_tx_pld_rst_n,
		input wire		in_pld_10g_rx_align_clr,
		input wire		in_pld_10g_rx_clr_ber_count,
		input wire		in_pld_10g_rx_rd_en,
		input wire	[6:0]	in_pld_10g_tx_bitslip,
		input wire		in_pld_10g_tx_burst_en,
		input wire		in_pld_10g_tx_data_valid,
		input wire	[1:0]	in_pld_10g_tx_diag_status,
		input wire		in_pld_10g_tx_wordslip,
		input wire		in_pld_8g_a1a2_size,
		input wire		in_pld_8g_bitloc_rev_en,
		input wire		in_pld_8g_byte_rev_en,
		input wire	[2:0]	in_pld_8g_eidleinfersel,
		input wire		in_pld_8g_encdt,
		input wire		in_pld_8g_g3_rx_pld_rst_n,
		input wire		in_pld_8g_g3_tx_pld_rst_n,
		input wire		in_pld_8g_rddisable_tx,
		input wire		in_pld_8g_rdenable_rx,
		input wire		in_pld_8g_refclk_dig2,
		input wire		in_pld_8g_rxpolarity,
		input wire	[4:0]	in_pld_8g_tx_boundary_sel,
		input wire		in_pld_8g_wrdisable_rx,
		input wire		in_pld_8g_wrenable_tx,
		input wire		in_pld_atpg_los_en_n,
		input wire		in_pld_bitslip,
		input wire	[17:0]	in_pld_g3_current_coeff,
		input wire	[2:0]	in_pld_g3_current_rxpreset,
		input wire		in_pld_ltr,
		input wire		in_pld_mem_krfec_atpg_rst_n,
		input wire		in_pld_partial_reconfig,
		input wire		in_pld_pcs_refclk_dig,
		input wire		in_pld_pma_adapt_start,
		input wire		in_pld_pma_csr_test_dis,
		input wire		in_pld_pma_early_eios,
		input wire	[5:0]	in_pld_pma_eye_monitor,
		input wire		in_pld_pma_ltd_b,
		input wire		in_pld_pma_nrpi_freeze,
		input wire	[1:0]	in_pld_pma_pcie_switch,
		input wire		in_pld_pma_ppm_lock,
		input wire	[4:0]	in_pld_pma_reserved_out,
		input wire		in_pld_pma_rs_lpbk_b,
		input wire		in_pld_pma_rx_qpi_pullup,
		input wire		in_pld_pma_rxpma_rstb,
		input wire		in_pld_pma_tx_bitslip,
		input wire		in_pld_pma_tx_bonding_rstb,
		input wire		in_pld_pma_tx_qpi_pulldn,
		input wire		in_pld_pma_tx_qpi_pullup,
		input wire		in_pld_pma_txdetectrx,
		input wire		in_pld_pma_txpma_rstb,
		input wire		in_pld_pmaif_rx_pld_rst_n,
		input wire		in_pld_pmaif_rxclkslip,
		input wire		in_pld_pmaif_tx_pld_rst_n,
		input wire		in_pld_polinv_rx,
		input wire		in_pld_polinv_tx,
		input wire	[1:0]	in_pld_rate,
		input wire	[9:0]	in_pld_reserved_in,
		input wire		in_pld_rx_clk,
		input wire		in_pld_rx_prbs_err_clr,
		input wire		in_pld_scan_mode_n,
		input wire		in_pld_scan_shift_n,
		input wire		in_pld_syncsm_en,
		input wire		in_pld_tx_clk,
		input wire	[17:0]	in_pld_tx_control,
		input wire	[127:0]	in_pld_tx_data,
		input wire		in_pld_txelecidle,
		input wire		in_pld_uhsif_tx_clk,
		input wire		in_pma_adapt_done,
		input wire		in_pma_clklow,
		input wire		in_pma_fref,
		input wire		in_pma_hclk,
		input wire	[1:0]	in_pma_pcie_sw_done,
		input wire		in_pma_pfdmode_lock,
		input wire	[4:0]	in_pma_reserved_in,
		input wire		in_pma_rx_clkdiv_user,
		input wire		in_pma_rx_detect_valid,
		input wire		in_pma_rx_found,
		input wire		in_pma_rx_pma_clk,
		input wire	[63:0]	in_pma_rx_pma_data,
		input wire		in_pma_rx_signal_ok,
		input wire		in_pma_rxpll_lock,
		input wire		in_pma_signal_det,
		input wire	[7:0]	in_pma_testbus,
		input wire		in_pma_tx_clkdiv_user,
		input wire		in_pma_tx_pma_clk,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen1_2,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen3,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pld_pcs_interface,
		output wire		out_blockselect_hssi_10g_rx_pcs,
		output wire		out_blockselect_hssi_10g_tx_pcs,
		output wire		out_blockselect_hssi_8g_rx_pcs,
		output wire		out_blockselect_hssi_8g_tx_pcs,
		output wire		out_blockselect_hssi_common_pcs_pma_interface,
		output wire		out_blockselect_hssi_common_pld_pcs_interface,
		output wire		out_blockselect_hssi_fifo_rx_pcs,
		output wire		out_blockselect_hssi_fifo_tx_pcs,
		output wire		out_blockselect_hssi_gen3_rx_pcs,
		output wire		out_blockselect_hssi_gen3_tx_pcs,
		output wire		out_blockselect_hssi_krfec_rx_pcs,
		output wire		out_blockselect_hssi_krfec_tx_pcs,
		output wire		out_blockselect_hssi_pipe_gen1_2,
		output wire		out_blockselect_hssi_pipe_gen3,
		output wire		out_blockselect_hssi_rx_pcs_pma_interface,
		output wire		out_blockselect_hssi_rx_pld_pcs_interface,
		output wire		out_blockselect_hssi_tx_pcs_pma_interface,
		output wire		out_blockselect_hssi_tx_pld_pcs_interface,
		output wire	[4:0]	out_bond_pcs10g_out_bot,
		output wire	[4:0]	out_bond_pcs10g_out_top,
		output wire	[12:0]	out_bond_pcs8g_out_bot,
		output wire	[12:0]	out_bond_pcs8g_out_top,
		output wire	[11:0]	out_bond_pmaif_out_bot,
		output wire	[11:0]	out_bond_pmaif_out_top,
		output wire	[2:0]	out_hip_clk_out,
		output wire	[7:0]	out_hip_ctrl_out,
		output wire		out_hip_iocsr_rdy,
		output wire		out_hip_iocsr_rdy_dly,
		output wire		out_hip_nfrzdrv,
		output wire		out_hip_npor,
		output wire	[50:0]	out_hip_rx_data,
		output wire		out_hip_usermode,
		output wire		out_pld_10g_krfec_rx_blk_lock,
		output wire	[1:0]	out_pld_10g_krfec_rx_diag_data_status,
		output wire		out_pld_10g_krfec_rx_frame,
		output wire		out_pld_10g_krfec_tx_frame,
		output wire		out_pld_10g_rx_align_val,
		output wire		out_pld_10g_rx_crc32_err,
		output wire		out_pld_10g_rx_data_valid,
		output wire		out_pld_10g_rx_empty,
		output wire		out_pld_10g_rx_fifo_del,
		output wire		out_pld_10g_rx_fifo_insert,
		output wire	[4:0]	out_pld_10g_rx_fifo_num,
		output wire		out_pld_10g_rx_frame_lock,
		output wire		out_pld_10g_rx_hi_ber,
		output wire		out_pld_10g_rx_oflw_err,
		output wire		out_pld_10g_rx_pempty,
		output wire		out_pld_10g_rx_pfull,
		output wire		out_pld_10g_tx_burst_en_exe,
		output wire		out_pld_10g_tx_empty,
		output wire	[3:0]	out_pld_10g_tx_fifo_num,
		output wire		out_pld_10g_tx_full,
		output wire		out_pld_10g_tx_pempty,
		output wire		out_pld_10g_tx_pfull,
		output wire		out_pld_10g_tx_wordslip_exe,
		output wire	[3:0]	out_pld_8g_a1a2_k1k2_flag,
		output wire		out_pld_8g_empty_rmf,
		output wire		out_pld_8g_empty_rx,
		output wire		out_pld_8g_empty_tx,
		output wire		out_pld_8g_full_rmf,
		output wire		out_pld_8g_full_rx,
		output wire		out_pld_8g_full_tx,
		output wire		out_pld_8g_rxelecidle,
		output wire		out_pld_8g_signal_detect_out,
		output wire	[4:0]	out_pld_8g_wa_boundary,
		output wire		out_pld_krfec_tx_alignment,
		output wire		out_pld_pcs_rx_clk_out,
		output wire		out_pld_pcs_tx_clk_out,
		output wire		out_pld_pma_adapt_done,
		output wire		out_pld_pma_clkdiv_rx_user,
		output wire		out_pld_pma_clkdiv_tx_user,
		output wire		out_pld_pma_clklow,
		output wire		out_pld_pma_fref,
		output wire		out_pld_pma_hclk,
		output wire	[1:0]	out_pld_pma_pcie_sw_done,
		output wire		out_pld_pma_pfdmode_lock,
		output wire	[4:0]	out_pld_pma_reserved_in,
		output wire		out_pld_pma_rx_clk_out,
		output wire		out_pld_pma_rx_detect_valid,
		output wire		out_pld_pma_rx_found,
		output wire		out_pld_pma_rxpll_lock,
		output wire		out_pld_pma_signal_ok,
		output wire	[7:0]	out_pld_pma_testbus,
		output wire		out_pld_pma_tx_clk_out,
		output wire		out_pld_pmaif_mask_tx_pll,
		output wire	[9:0]	out_pld_reserved_out,
		output wire	[19:0]	out_pld_rx_control,
		output wire	[127:0]	out_pld_rx_data,
		output wire		out_pld_rx_prbs_done,
		output wire		out_pld_rx_prbs_err,
		output wire	[19:0]	out_pld_test_data,
		output wire		out_pld_uhsif_lock,
		output wire		out_pld_uhsif_tx_clk_out,
		output wire		out_pma_adapt_start,
		output wire		out_pma_atpg_los_en_n,
		output wire		out_pma_csr_test_dis,
		output wire	[17:0]	out_pma_current_coeff,
		output wire	[2:0]	out_pma_current_rxpreset,
		output wire		out_pma_early_eios,
		output wire	[5:0]	out_pma_eye_monitor,
		output wire	[1:0]	out_pma_interface_select,
		output wire		out_pma_ltd_b,
		output wire		out_pma_ltr,
		output wire		out_pma_nfrzdrv,
		output wire		out_pma_nrpi_freeze,
		output wire	[1:0]	out_pma_pcie_switch,
		output wire		out_pma_ppm_lock,
		output wire	[4:0]	out_pma_reserved_out,
		output wire		out_pma_rs_lpbk_b,
		output wire		out_pma_rx_clkslip,
		output wire		out_pma_rx_qpi_pullup,
		output wire		out_pma_rxpma_rstb,
		output wire		out_pma_scan_mode_n,
		output wire		out_pma_scan_shift_n,
		output wire		out_pma_tx_bitslip,
		output wire		out_pma_tx_bonding_rstb,
		output wire		out_pma_tx_elec_idle,
		output wire	[63:0]	out_pma_tx_pma_data,
		output wire		out_pma_tx_qpi_pulldn,
		output wire		out_pma_tx_qpi_pullup,
		output wire		out_pma_tx_txdetectrx,
		output wire		out_pma_txpma_rstb
	//PORT_LIST_END
	);
	//wire declarations
	
	// wires for module twentynm_hssi_fifo_tx_pcs
	wire	[7:0]	w_hssi_fifo_tx_pcs_avmmreaddata;
	wire		w_hssi_fifo_tx_pcs_blockselect;
	wire	[72:0]	w_hssi_fifo_tx_pcs_data_out_10g;
	wire	[63:0]	w_hssi_fifo_tx_pcs_data_out_8g_phase_comp;
	
	// wires for module twentynm_hssi_gen3_rx_pcs
	wire	[7:0]	w_hssi_gen3_rx_pcs_avmmreaddata;
	wire		w_hssi_gen3_rx_pcs_blk_algnd_int;
	wire		w_hssi_gen3_rx_pcs_blk_start;
	wire		w_hssi_gen3_rx_pcs_blockselect;
	wire		w_hssi_gen3_rx_pcs_clkcomp_delete_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_insert_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_overfl_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_undfl_int;
	wire	[31:0]	w_hssi_gen3_rx_pcs_data_out;
	wire		w_hssi_gen3_rx_pcs_data_valid;
	wire		w_hssi_gen3_rx_pcs_ei_det_int;
	wire		w_hssi_gen3_rx_pcs_ei_partial_det_int;
	wire		w_hssi_gen3_rx_pcs_err_decode_int;
	wire		w_hssi_gen3_rx_pcs_i_det_int;
	wire		w_hssi_gen3_rx_pcs_lpbk_blk_start;
	wire	[33:0]	w_hssi_gen3_rx_pcs_lpbk_data;
	wire		w_hssi_gen3_rx_pcs_lpbk_data_valid;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk;
	wire	[39:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n;
	wire		w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int;
	wire	[19:0]	w_hssi_gen3_rx_pcs_rx_test_out;
	wire	[1:0]	w_hssi_gen3_rx_pcs_sync_hdr;
	
	// wires for module twentynm_hssi_krfec_tx_pcs
	wire	[7:0]	w_hssi_krfec_tx_pcs_avmmreaddata;
	wire		w_hssi_krfec_tx_pcs_blockselect;
	wire		w_hssi_krfec_tx_pcs_tx_alignment;
	wire	[63:0]	w_hssi_krfec_tx_pcs_tx_data_out;
	wire		w_hssi_krfec_tx_pcs_tx_frame;
	wire	[19:0]	w_hssi_krfec_tx_pcs_tx_test_data;
	
	// wires for module twentynm_hssi_krfec_rx_pcs
	wire	[7:0]	w_hssi_krfec_rx_pcs_avmmreaddata;
	wire		w_hssi_krfec_rx_pcs_blockselect;
	wire		w_hssi_krfec_rx_pcs_rx_block_lock;
	wire	[9:0]	w_hssi_krfec_rx_pcs_rx_control_out;
	wire	[63:0]	w_hssi_krfec_rx_pcs_rx_data_out;
	wire	[1:0]	w_hssi_krfec_rx_pcs_rx_data_status;
	wire		w_hssi_krfec_rx_pcs_rx_data_valid_out;
	wire		w_hssi_krfec_rx_pcs_rx_frame;
	wire		w_hssi_krfec_rx_pcs_rx_signal_ok_out;
	
	// wires for module twentynm_hssi_rx_pld_pcs_interface
	wire	[7:0]	w_hssi_rx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_rx_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_hip_rx_ctrl;
	wire	[50:0]	w_hssi_rx_pld_pcs_interface_hip_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
	wire	[3:0]	w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary;
	wire		w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_pld_rx_control;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_pld_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
	
	// wires for module twentynm_hssi_common_pld_pcs_interface
	wire	[7:0]	w_hssi_common_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_common_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_hip_cmn_clk;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_hip_cmn_ctrl;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
	wire		w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_hip_npor;
	wire		w_hssi_common_pld_pcs_interface_hip_usermode;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n;
	wire	[17:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel;
	wire		w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_clklow;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_fref;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_hclk;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_pld_pma_reserved_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
	wire	[7:0]	w_hssi_common_pld_pcs_interface_pld_pma_testbus;
	wire		w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
	wire	[9:0]	w_hssi_common_pld_pcs_interface_pld_reserved_out;
	wire	[19:0]	w_hssi_common_pld_pcs_interface_pld_test_data;
	wire		w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
	wire		w_hssi_common_pld_pcs_interface_scan_mode_n;
	
	// wires for module twentynm_hssi_10g_rx_pcs
	wire	[7:0]	w_hssi_10g_rx_pcs_avmmreaddata;
	wire		w_hssi_10g_rx_pcs_blockselect;
	wire		w_hssi_10g_rx_pcs_rx_align_val;
	wire		w_hssi_10g_rx_pcs_rx_blk_lock;
	wire		w_hssi_10g_rx_pcs_rx_clk_out;
	wire		w_hssi_10g_rx_pcs_rx_clk_out_pld_if;
	wire	[19:0]	w_hssi_10g_rx_pcs_rx_control;
	wire		w_hssi_10g_rx_pcs_rx_crc32_err;
	wire	[127:0]	w_hssi_10g_rx_pcs_rx_data;
	wire		w_hssi_10g_rx_pcs_rx_data_valid;
	wire		w_hssi_10g_rx_pcs_rx_dft_clk_out;
	wire	[1:0]	w_hssi_10g_rx_pcs_rx_diag_status;
	wire		w_hssi_10g_rx_pcs_rx_empty;
	wire		w_hssi_10g_rx_pcs_rx_fec_clk;
	wire		w_hssi_10g_rx_pcs_rx_fifo_del;
	wire		w_hssi_10g_rx_pcs_rx_fifo_insert;
	wire	[4:0]	w_hssi_10g_rx_pcs_rx_fifo_num;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_clk;
	wire	[73:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_data;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_en;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_ptr;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_frame_lock;
	wire		w_hssi_10g_rx_pcs_rx_hi_ber;
	wire		w_hssi_10g_rx_pcs_rx_master_clk;
	wire		w_hssi_10g_rx_pcs_rx_master_clk_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_oflw_err;
	wire		w_hssi_10g_rx_pcs_rx_pempty;
	wire		w_hssi_10g_rx_pcs_rx_pfull;
	wire		w_hssi_10g_rx_pcs_rx_random_err;
	wire		w_hssi_10g_rx_pcs_rx_rx_frame;
	
	// wires for module twentynm_hssi_tx_pld_pcs_interface
	wire	[7:0]	w_hssi_tx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_tx_pld_pcs_interface_blockselect;
	wire		w_hssi_tx_pld_pcs_interface_hip_tx_clk;
	wire	[6:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en;
	wire	[17:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control;
	wire	[8:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg;
	wire	[127:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start;
	wire	[4:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle;
	wire	[2:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
	wire		w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
	
	// wires for module twentynm_hssi_tx_pcs_pma_interface
	wire	[7:0]	w_hssi_tx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_tx_pcs_pma_interface_blockselect;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out;
	wire	[4:0]	w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk;
	wire		w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_pma_tx_pma_data;
	wire		w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_1;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_2;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_3;
	
	// wires for module twentynm_hssi_rx_pcs_pma_interface
	wire	[7:0]	w_hssi_rx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_rx_pcs_pma_interface_blockselect;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni;
	wire	[31:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok;
	wire		w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk;
	wire	[5:0]	w_hssi_rx_pcs_pma_interface_pma_eye_monitor;
	wire		w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
	wire		w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test;
	
	// wires for module twentynm_hssi_10g_tx_pcs
	wire	[7:0]	w_hssi_10g_tx_pcs_avmmreaddata;
	wire		w_hssi_10g_tx_pcs_blockselect;
	wire		w_hssi_10g_tx_pcs_distdwn_out_dv;
	wire		w_hssi_10g_tx_pcs_distdwn_out_rden;
	wire		w_hssi_10g_tx_pcs_distdwn_out_wren;
	wire		w_hssi_10g_tx_pcs_distup_out_dv;
	wire		w_hssi_10g_tx_pcs_distup_out_rden;
	wire		w_hssi_10g_tx_pcs_distup_out_wren;
	wire		w_hssi_10g_tx_pcs_tx_burst_en_exe;
	wire		w_hssi_10g_tx_pcs_tx_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pma_if;
	wire	[8:0]	w_hssi_10g_tx_pcs_tx_control_out_krfec;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_data_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_data_valid_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_dft_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_empty;
	wire		w_hssi_10g_tx_pcs_tx_fec_clk;
	wire	[3:0]	w_hssi_10g_tx_pcs_tx_fifo_num;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_rd_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_clk;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_en;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_frame;
	wire		w_hssi_10g_tx_pcs_tx_full;
	wire		w_hssi_10g_tx_pcs_tx_master_clk;
	wire		w_hssi_10g_tx_pcs_tx_master_clk_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_pempty;
	wire		w_hssi_10g_tx_pcs_tx_pfull;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_data;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_gating_val;
	wire	[19:0]	w_hssi_10g_tx_pcs_tx_test_data;
	wire		w_hssi_10g_tx_pcs_tx_wordslip_exe;
	
	// wires for module twentynm_hssi_8g_tx_pcs
	wire	[7:0]	w_hssi_8g_tx_pcs_avmmreaddata;
	wire		w_hssi_8g_tx_pcs_blockselect;
	wire		w_hssi_8g_tx_pcs_clk_out;
	wire		w_hssi_8g_tx_pcs_clk_out_gen3;
	wire	[19:0]	w_hssi_8g_tx_pcs_dataout;
	wire		w_hssi_8g_tx_pcs_dyn_clk_switch_n;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn;
	wire		w_hssi_8g_tx_pcs_g3_tx_pma_rstn;
	wire	[2:0]	w_hssi_8g_tx_pcs_non_gray_eidleinfersel;
	wire		w_hssi_8g_tx_pcs_ph_fifo_overflow;
	wire		w_hssi_8g_tx_pcs_ph_fifo_underflow;
	wire		w_hssi_8g_tx_pcs_phfifo_txdeemph;
	wire	[2:0]	w_hssi_8g_tx_pcs_phfifo_txmargin;
	wire		w_hssi_8g_tx_pcs_phfifo_txswing;
	wire		w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out;
	wire	[1:0]	w_hssi_8g_tx_pcs_pipe_power_down_out;
	wire		w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3;
	wire		w_hssi_8g_tx_pcs_pmaif_asn_rstn;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_refclk_b;
	wire		w_hssi_8g_tx_pcs_refclk_b_reset;
	wire		w_hssi_8g_tx_pcs_rxpolarity_int;
	wire		w_hssi_8g_tx_pcs_soft_reset_wclk1_n;
	wire		w_hssi_8g_tx_pcs_sw_fifo_wr_clk;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_blk_start_out;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_ctrlplane_testbus;
	wire	[31:0]	w_hssi_8g_tx_pcs_tx_data_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_data_valid_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_datak_out;
	wire		w_hssi_8g_tx_pcs_tx_detect_rxloopback_int;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_tx_pipe_clk;
	wire		w_hssi_8g_tx_pcs_tx_pipe_electidle;
	wire		w_hssi_8g_tx_pcs_tx_pipe_soft_reset;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_sync_hdr_out;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_testbus;
	wire		w_hssi_8g_tx_pcs_txcompliance_out;
	wire		w_hssi_8g_tx_pcs_txelecidle_out;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk;
	wire	[63:0]	w_hssi_8g_tx_pcs_wr_data_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_en_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo;
	
	// wires for module twentynm_hssi_pipe_gen3
	wire	[7:0]	w_hssi_pipe_gen3_avmmreaddata;
	wire		w_hssi_pipe_gen3_blockselect;
	wire		w_hssi_pipe_gen3_gen3_clk_sel;
	wire		w_hssi_pipe_gen3_pcs_rst;
	wire		w_hssi_pipe_gen3_phystatus;
	wire	[17:0]	w_hssi_pipe_gen3_pma_current_coeff;
	wire	[2:0]	w_hssi_pipe_gen3_pma_current_rxpreset;
	wire		w_hssi_pipe_gen3_pma_tx_elec_idle;
	wire		w_hssi_pipe_gen3_pma_txdetectrx;
	wire		w_hssi_pipe_gen3_rev_lpbk_8gpcs_out;
	wire		w_hssi_pipe_gen3_rev_lpbk_int;
	wire	[3:0]	w_hssi_pipe_gen3_rx_blk_start;
	wire	[1:0]	w_hssi_pipe_gen3_rx_sync_hdr;
	wire	[63:0]	w_hssi_pipe_gen3_rxd_8gpcs_out;
	wire	[3:0]	w_hssi_pipe_gen3_rxdataskip;
	wire		w_hssi_pipe_gen3_rxelecidle;
	wire		w_hssi_pipe_gen3_rxpolarity_8gpcs_out;
	wire		w_hssi_pipe_gen3_rxpolarity_int;
	wire	[2:0]	w_hssi_pipe_gen3_rxstatus;
	wire		w_hssi_pipe_gen3_rxvalid;
	wire		w_hssi_pipe_gen3_shutdown_clk;
	wire	[19:0]	w_hssi_pipe_gen3_test_out;
	wire		w_hssi_pipe_gen3_tx_blk_start_int;
	wire	[1:0]	w_hssi_pipe_gen3_tx_sync_hdr_int;
	wire	[31:0]	w_hssi_pipe_gen3_txdata_int;
	wire	[3:0]	w_hssi_pipe_gen3_txdatak_int;
	wire		w_hssi_pipe_gen3_txdataskip_int;
	
	// wires for module twentynm_hssi_pipe_gen1_2
	wire	[7:0]	w_hssi_pipe_gen1_2_avmmreaddata;
	wire		w_hssi_pipe_gen1_2_blockselect;
	wire	[17:0]	w_hssi_pipe_gen1_2_current_coeff;
	wire		w_hssi_pipe_gen1_2_phystatus;
	wire		w_hssi_pipe_gen1_2_polarity_inversion_rx;
	wire		w_hssi_pipe_gen1_2_rev_loopbk;
	wire		w_hssi_pipe_gen1_2_rxelecidle;
	wire		w_hssi_pipe_gen1_2_rxelectricalidle_out;
	wire	[2:0]	w_hssi_pipe_gen1_2_rxstatus;
	wire		w_hssi_pipe_gen1_2_rxvalid;
	wire		w_hssi_pipe_gen1_2_tx_elec_idle_out;
	wire		w_hssi_pipe_gen1_2_txdetectrx;
	
	// wires for module twentynm_hssi_gen3_tx_pcs
	wire	[7:0]	w_hssi_gen3_tx_pcs_avmmreaddata;
	wire		w_hssi_gen3_tx_pcs_blockselect;
	wire	[31:0]	w_hssi_gen3_tx_pcs_data_out;
	wire	[35:0]	w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out;
	wire	[31:0]	w_hssi_gen3_tx_pcs_par_lpbk_out;
	wire	[19:0]	w_hssi_gen3_tx_pcs_tx_test_out;
	
	// wires for module twentynm_hssi_8g_rx_pcs
	wire	[3:0]	w_hssi_8g_rx_pcs_a1a2k1k2flag;
	wire	[7:0]	w_hssi_8g_rx_pcs_avmmreaddata;
	wire		w_hssi_8g_rx_pcs_blockselect;
	wire	[19:0]	w_hssi_8g_rx_pcs_chnl_test_bus_out;
	wire		w_hssi_8g_rx_pcs_clock_to_pld;
	wire	[63:0]	w_hssi_8g_rx_pcs_dataout;
	wire		w_hssi_8g_rx_pcs_dis_pc_byte;
	wire		w_hssi_8g_rx_pcs_eidle_detected;
	wire	[2:0]	w_hssi_8g_rx_pcs_eios_det_cdr_ctrl;
	wire		w_hssi_8g_rx_pcs_g3_rx_pma_rstn;
	wire		w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn;
	wire		w_hssi_8g_rx_pcs_gen2ngen1;
	wire	[19:0]	w_hssi_8g_rx_pcs_parallel_rev_loopback;
	wire		w_hssi_8g_rx_pcs_pc_fifo_empty;
	wire		w_hssi_8g_rx_pcs_pcfifofull;
	wire		w_hssi_8g_rx_pcs_phystatus;
	wire	[63:0]	w_hssi_8g_rx_pcs_pipe_data;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_up;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo;
	wire	[7:0]	w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rm_fifo_empty;
	wire		w_hssi_8g_rx_pcs_rm_fifo_full;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_blk_start;
	wire		w_hssi_8g_rx_pcs_rx_clk_out_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clkslip;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_data_valid;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rx_pipe_clk;
	wire		w_hssi_8g_rx_pcs_rx_pipe_soft_reset;
	wire		w_hssi_8g_rx_pcs_rx_pma_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_sync_hdr;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_up;
	wire	[2:0]	w_hssi_8g_rx_pcs_rxstatus;
	wire		w_hssi_8g_rx_pcs_rxvalid;
	wire		w_hssi_8g_rx_pcs_signal_detect_out;
	wire	[4:0]	w_hssi_8g_rx_pcs_word_align_boundary;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk;
	wire	[79:0]	w_hssi_8g_rx_pcs_wr_data_rx_phfifo;
	wire	[31:0]	w_hssi_8g_rx_pcs_wr_data_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo;
	
	// wires for module twentynm_hssi_fifo_rx_pcs
	wire	[7:0]	w_hssi_fifo_rx_pcs_avmmreaddata;
	wire		w_hssi_fifo_rx_pcs_blockselect;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out2_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out_8g_clock_comp;
	wire	[79:0]	w_hssi_fifo_rx_pcs_data_out_8g_phase_comp;
	wire	[39:0]	w_hssi_fifo_rx_pcs_data_out_gen3;
	
	// wires for module twentynm_hssi_common_pcs_pma_interface
	wire	[7:0]	w_hssi_common_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_common_pcs_pma_interface_blockselect;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in;
	wire	[19:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out;
	wire	[7:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus;
	wire		w_hssi_common_pcs_pma_interface_pma_adapt_start;
	wire		w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
	wire		w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
	wire	[17:0]	w_hssi_common_pcs_pma_interface_pma_current_coeff;
	wire	[2:0]	w_hssi_common_pcs_pma_interface_pma_current_rxpreset;
	wire		w_hssi_common_pcs_pma_interface_pma_early_eios;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_interface_select;
	wire		w_hssi_common_pcs_pma_interface_pma_ltd_b;
	wire		w_hssi_common_pcs_pma_interface_pma_ltr;
	wire		w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
	wire		w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_pcie_switch;
	wire		w_hssi_common_pcs_pma_interface_pma_ppm_lock;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_pma_reserved_out;
	wire		w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
	wire		w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up;
	
	
	generate
		
		//module instantiations
		
		// instantiating twentynm_hssi_10g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_rx_pcs
			twentynm_hssi_10g_rx_pcs #(
				.advanced_user_mode(hssi_10g_rx_pcs_advanced_user_mode),
				.align_del(hssi_10g_rx_pcs_align_del),
				.ber_bit_err_total_cnt(hssi_10g_rx_pcs_ber_bit_err_total_cnt),
				.ber_clken(hssi_10g_rx_pcs_ber_clken),
				.ber_xus_timer_window(hssi_10g_rx_pcs_ber_xus_timer_window),
				.bitslip_mode(hssi_10g_rx_pcs_bitslip_mode),
				.blksync_bitslip_type(hssi_10g_rx_pcs_blksync_bitslip_type),
				.blksync_bitslip_wait_cnt(hssi_10g_rx_pcs_blksync_bitslip_wait_cnt),
				.blksync_bitslip_wait_type(hssi_10g_rx_pcs_blksync_bitslip_wait_type),
				.blksync_bypass(hssi_10g_rx_pcs_blksync_bypass),
				.blksync_clken(hssi_10g_rx_pcs_blksync_clken),
				.blksync_enum_invalid_sh_cnt(hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt),
				.blksync_knum_sh_cnt_postlock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock),
				.blksync_knum_sh_cnt_prelock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock),
				.blksync_pipeln(hssi_10g_rx_pcs_blksync_pipeln),
				.clr_errblk_cnt_en(hssi_10g_rx_pcs_clr_errblk_cnt_en),
				.control_del(hssi_10g_rx_pcs_control_del),
				.crcchk_bypass(hssi_10g_rx_pcs_crcchk_bypass),
				.crcchk_clken(hssi_10g_rx_pcs_crcchk_clken),
				.crcchk_inv(hssi_10g_rx_pcs_crcchk_inv),
				.crcchk_pipeln(hssi_10g_rx_pcs_crcchk_pipeln),
				.crcflag_pipeln(hssi_10g_rx_pcs_crcflag_pipeln),
				.ctrl_bit_reverse(hssi_10g_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_10g_rx_pcs_data_bit_reverse),
				.dec64b66b_clken(hssi_10g_rx_pcs_dec64b66b_clken),
				.dec_64b66b_rxsm_bypass(hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass),
				.descrm_bypass(hssi_10g_rx_pcs_descrm_bypass),
				.descrm_clken(hssi_10g_rx_pcs_descrm_clken),
				.descrm_mode(hssi_10g_rx_pcs_descrm_mode),
				.descrm_pipeln(hssi_10g_rx_pcs_descrm_pipeln),
				.dft_clk_out_sel(hssi_10g_rx_pcs_dft_clk_out_sel),
				.dis_signal_ok(hssi_10g_rx_pcs_dis_signal_ok),
				.dispchk_bypass(hssi_10g_rx_pcs_dispchk_bypass),
				.empty_flag_type(hssi_10g_rx_pcs_empty_flag_type),
				.fast_path(hssi_10g_rx_pcs_fast_path),
				.fec_clken(hssi_10g_rx_pcs_fec_clken),
				.fec_enable(hssi_10g_rx_pcs_fec_enable),
				.fifo_double_read(hssi_10g_rx_pcs_fifo_double_read),
				.fifo_stop_rd(hssi_10g_rx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_rx_pcs_fifo_stop_wr),
				.force_align(hssi_10g_rx_pcs_force_align),
				.frmsync_bypass(hssi_10g_rx_pcs_frmsync_bypass),
				.frmsync_clken(hssi_10g_rx_pcs_frmsync_clken),
				.frmsync_enum_scrm(hssi_10g_rx_pcs_frmsync_enum_scrm),
				.frmsync_enum_sync(hssi_10g_rx_pcs_frmsync_enum_sync),
				.frmsync_flag_type(hssi_10g_rx_pcs_frmsync_flag_type),
				.frmsync_knum_sync(hssi_10g_rx_pcs_frmsync_knum_sync),
				.frmsync_mfrm_length(hssi_10g_rx_pcs_frmsync_mfrm_length),
				.frmsync_pipeln(hssi_10g_rx_pcs_frmsync_pipeln),
				.full_flag_type(hssi_10g_rx_pcs_full_flag_type),
				.gb_rx_idwidth(hssi_10g_rx_pcs_gb_rx_idwidth),
				.gb_rx_odwidth(hssi_10g_rx_pcs_gb_rx_odwidth),
				.gbexp_clken(hssi_10g_rx_pcs_gbexp_clken),
				.low_latency_en(hssi_10g_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_10g_rx_pcs_lpbk_mode),
				.master_clk_sel(hssi_10g_rx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_rx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_rx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_rx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_rx_pcs_pld_if_type),
				.prot_mode(hssi_10g_rx_pcs_prot_mode),
				.rand_clken(hssi_10g_rx_pcs_rand_clken),
				.rd_clk_sel(hssi_10g_rx_pcs_rd_clk_sel),
				.rdfifo_clken(hssi_10g_rx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_rx_pcs_reconfig_settings),
				.rx_fifo_write_ctrl(hssi_10g_rx_pcs_rx_fifo_write_ctrl),
				.rx_scrm_width(hssi_10g_rx_pcs_rx_scrm_width),
				.rx_sh_location(hssi_10g_rx_pcs_rx_sh_location),
				.rx_signal_ok_sel(hssi_10g_rx_pcs_rx_signal_ok_sel),
				.rx_sm_bypass(hssi_10g_rx_pcs_rx_sm_bypass),
				.rx_sm_hiber(hssi_10g_rx_pcs_rx_sm_hiber),
				.rx_sm_pipeln(hssi_10g_rx_pcs_rx_sm_pipeln),
				.rx_testbus_sel(hssi_10g_rx_pcs_rx_testbus_sel),
				.rx_true_b2b(hssi_10g_rx_pcs_rx_true_b2b),
				.rxfifo_empty(hssi_10g_rx_pcs_rxfifo_empty),
				.rxfifo_full(hssi_10g_rx_pcs_rxfifo_full),
				.rxfifo_mode(hssi_10g_rx_pcs_rxfifo_mode),
				.rxfifo_pempty(hssi_10g_rx_pcs_rxfifo_pempty),
				.rxfifo_pfull(hssi_10g_rx_pcs_rxfifo_pfull),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.stretch_num_stages(hssi_10g_rx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_rx_pcs_sup_mode),
				.test_mode(hssi_10g_rx_pcs_test_mode),
				.wrfifo_clken(hssi_10g_rx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_rx_pcs_blockselect),
				.rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.rx_control(w_hssi_10g_rx_pcs_rx_control),
				.rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.rx_data(w_hssi_10g_rx_pcs_rx_data),
				.rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.rx_diag_status(w_hssi_10g_rx_pcs_rx_diag_status),
				.rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.rx_fec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.rx_fifo_num(w_hssi_10g_rx_pcs_rx_fifo_num),
				.rx_fifo_rd_ptr(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr),
				.rx_fifo_rd_ptr2(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2),
				.rx_fifo_wr_clk(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.rx_fifo_wr_data(w_hssi_10g_rx_pcs_rx_fifo_wr_data),
				.rx_fifo_wr_en(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.rx_fifo_wr_ptr(w_hssi_10g_rx_pcs_rx_fifo_wr_ptr),
				.rx_fifo_wr_rst_n(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.rx_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_rx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_rx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.rx_control_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0]}),
				.rx_control_in_krfec({w_hssi_krfec_rx_pcs_rx_control_out[9], w_hssi_krfec_rx_pcs_rx_control_out[8], w_hssi_krfec_rx_pcs_rx_control_out[7], w_hssi_krfec_rx_pcs_rx_control_out[6], w_hssi_krfec_rx_pcs_rx_control_out[5], w_hssi_krfec_rx_pcs_rx_control_out[4], w_hssi_krfec_rx_pcs_rx_control_out[3], w_hssi_krfec_rx_pcs_rx_control_out[2], w_hssi_krfec_rx_pcs_rx_control_out[1], w_hssi_krfec_rx_pcs_rx_control_out[0]}),
				.rx_data_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0]}),
				.rx_data_in_krfec({w_hssi_krfec_rx_pcs_rx_data_out[63], w_hssi_krfec_rx_pcs_rx_data_out[62], w_hssi_krfec_rx_pcs_rx_data_out[61], w_hssi_krfec_rx_pcs_rx_data_out[60], w_hssi_krfec_rx_pcs_rx_data_out[59], w_hssi_krfec_rx_pcs_rx_data_out[58], w_hssi_krfec_rx_pcs_rx_data_out[57], w_hssi_krfec_rx_pcs_rx_data_out[56], w_hssi_krfec_rx_pcs_rx_data_out[55], w_hssi_krfec_rx_pcs_rx_data_out[54], w_hssi_krfec_rx_pcs_rx_data_out[53], w_hssi_krfec_rx_pcs_rx_data_out[52], w_hssi_krfec_rx_pcs_rx_data_out[51], w_hssi_krfec_rx_pcs_rx_data_out[50], w_hssi_krfec_rx_pcs_rx_data_out[49], w_hssi_krfec_rx_pcs_rx_data_out[48], w_hssi_krfec_rx_pcs_rx_data_out[47], w_hssi_krfec_rx_pcs_rx_data_out[46], w_hssi_krfec_rx_pcs_rx_data_out[45], w_hssi_krfec_rx_pcs_rx_data_out[44], w_hssi_krfec_rx_pcs_rx_data_out[43], w_hssi_krfec_rx_pcs_rx_data_out[42], w_hssi_krfec_rx_pcs_rx_data_out[41], w_hssi_krfec_rx_pcs_rx_data_out[40], w_hssi_krfec_rx_pcs_rx_data_out[39], w_hssi_krfec_rx_pcs_rx_data_out[38], w_hssi_krfec_rx_pcs_rx_data_out[37], w_hssi_krfec_rx_pcs_rx_data_out[36], w_hssi_krfec_rx_pcs_rx_data_out[35], w_hssi_krfec_rx_pcs_rx_data_out[34], w_hssi_krfec_rx_pcs_rx_data_out[33], w_hssi_krfec_rx_pcs_rx_data_out[32], w_hssi_krfec_rx_pcs_rx_data_out[31], w_hssi_krfec_rx_pcs_rx_data_out[30], w_hssi_krfec_rx_pcs_rx_data_out[29], w_hssi_krfec_rx_pcs_rx_data_out[28], w_hssi_krfec_rx_pcs_rx_data_out[27], w_hssi_krfec_rx_pcs_rx_data_out[26], w_hssi_krfec_rx_pcs_rx_data_out[25], w_hssi_krfec_rx_pcs_rx_data_out[24], w_hssi_krfec_rx_pcs_rx_data_out[23], w_hssi_krfec_rx_pcs_rx_data_out[22], w_hssi_krfec_rx_pcs_rx_data_out[21], w_hssi_krfec_rx_pcs_rx_data_out[20], w_hssi_krfec_rx_pcs_rx_data_out[19], w_hssi_krfec_rx_pcs_rx_data_out[18], w_hssi_krfec_rx_pcs_rx_data_out[17], w_hssi_krfec_rx_pcs_rx_data_out[16], w_hssi_krfec_rx_pcs_rx_data_out[15], w_hssi_krfec_rx_pcs_rx_data_out[14], w_hssi_krfec_rx_pcs_rx_data_out[13], w_hssi_krfec_rx_pcs_rx_data_out[12], w_hssi_krfec_rx_pcs_rx_data_out[11], w_hssi_krfec_rx_pcs_rx_data_out[10], w_hssi_krfec_rx_pcs_rx_data_out[9], w_hssi_krfec_rx_pcs_rx_data_out[8], w_hssi_krfec_rx_pcs_rx_data_out[7], w_hssi_krfec_rx_pcs_rx_data_out[6], w_hssi_krfec_rx_pcs_rx_data_out[5], w_hssi_krfec_rx_pcs_rx_data_out[4], w_hssi_krfec_rx_pcs_rx_data_out[3], w_hssi_krfec_rx_pcs_rx_data_out[2], w_hssi_krfec_rx_pcs_rx_data_out[1], w_hssi_krfec_rx_pcs_rx_data_out[0]}),
				.rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.rx_data_valid_in_krfec(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_10g[73], w_hssi_fifo_rx_pcs_data_out_10g[72], w_hssi_fifo_rx_pcs_data_out_10g[71], w_hssi_fifo_rx_pcs_data_out_10g[70], w_hssi_fifo_rx_pcs_data_out_10g[69], w_hssi_fifo_rx_pcs_data_out_10g[68], w_hssi_fifo_rx_pcs_data_out_10g[67], w_hssi_fifo_rx_pcs_data_out_10g[66], w_hssi_fifo_rx_pcs_data_out_10g[65], w_hssi_fifo_rx_pcs_data_out_10g[64], w_hssi_fifo_rx_pcs_data_out_10g[63], w_hssi_fifo_rx_pcs_data_out_10g[62], w_hssi_fifo_rx_pcs_data_out_10g[61], w_hssi_fifo_rx_pcs_data_out_10g[60], w_hssi_fifo_rx_pcs_data_out_10g[59], w_hssi_fifo_rx_pcs_data_out_10g[58], w_hssi_fifo_rx_pcs_data_out_10g[57], w_hssi_fifo_rx_pcs_data_out_10g[56], w_hssi_fifo_rx_pcs_data_out_10g[55], w_hssi_fifo_rx_pcs_data_out_10g[54], w_hssi_fifo_rx_pcs_data_out_10g[53], w_hssi_fifo_rx_pcs_data_out_10g[52], w_hssi_fifo_rx_pcs_data_out_10g[51], w_hssi_fifo_rx_pcs_data_out_10g[50], w_hssi_fifo_rx_pcs_data_out_10g[49], w_hssi_fifo_rx_pcs_data_out_10g[48], w_hssi_fifo_rx_pcs_data_out_10g[47], w_hssi_fifo_rx_pcs_data_out_10g[46], w_hssi_fifo_rx_pcs_data_out_10g[45], w_hssi_fifo_rx_pcs_data_out_10g[44], w_hssi_fifo_rx_pcs_data_out_10g[43], w_hssi_fifo_rx_pcs_data_out_10g[42], w_hssi_fifo_rx_pcs_data_out_10g[41], w_hssi_fifo_rx_pcs_data_out_10g[40], w_hssi_fifo_rx_pcs_data_out_10g[39], w_hssi_fifo_rx_pcs_data_out_10g[38], w_hssi_fifo_rx_pcs_data_out_10g[37], w_hssi_fifo_rx_pcs_data_out_10g[36], w_hssi_fifo_rx_pcs_data_out_10g[35], w_hssi_fifo_rx_pcs_data_out_10g[34], w_hssi_fifo_rx_pcs_data_out_10g[33], w_hssi_fifo_rx_pcs_data_out_10g[32], w_hssi_fifo_rx_pcs_data_out_10g[31], w_hssi_fifo_rx_pcs_data_out_10g[30], w_hssi_fifo_rx_pcs_data_out_10g[29], w_hssi_fifo_rx_pcs_data_out_10g[28], w_hssi_fifo_rx_pcs_data_out_10g[27], w_hssi_fifo_rx_pcs_data_out_10g[26], w_hssi_fifo_rx_pcs_data_out_10g[25], w_hssi_fifo_rx_pcs_data_out_10g[24], w_hssi_fifo_rx_pcs_data_out_10g[23], w_hssi_fifo_rx_pcs_data_out_10g[22], w_hssi_fifo_rx_pcs_data_out_10g[21], w_hssi_fifo_rx_pcs_data_out_10g[20], w_hssi_fifo_rx_pcs_data_out_10g[19], w_hssi_fifo_rx_pcs_data_out_10g[18], w_hssi_fifo_rx_pcs_data_out_10g[17], w_hssi_fifo_rx_pcs_data_out_10g[16], w_hssi_fifo_rx_pcs_data_out_10g[15], w_hssi_fifo_rx_pcs_data_out_10g[14], w_hssi_fifo_rx_pcs_data_out_10g[13], w_hssi_fifo_rx_pcs_data_out_10g[12], w_hssi_fifo_rx_pcs_data_out_10g[11], w_hssi_fifo_rx_pcs_data_out_10g[10], w_hssi_fifo_rx_pcs_data_out_10g[9], w_hssi_fifo_rx_pcs_data_out_10g[8], w_hssi_fifo_rx_pcs_data_out_10g[7], w_hssi_fifo_rx_pcs_data_out_10g[6], w_hssi_fifo_rx_pcs_data_out_10g[5], w_hssi_fifo_rx_pcs_data_out_10g[4], w_hssi_fifo_rx_pcs_data_out_10g[3], w_hssi_fifo_rx_pcs_data_out_10g[2], w_hssi_fifo_rx_pcs_data_out_10g[1], w_hssi_fifo_rx_pcs_data_out_10g[0]}),
				.rx_fifo_rd_data_dw({w_hssi_fifo_rx_pcs_data_out2_10g[73], w_hssi_fifo_rx_pcs_data_out2_10g[72], w_hssi_fifo_rx_pcs_data_out2_10g[71], w_hssi_fifo_rx_pcs_data_out2_10g[70], w_hssi_fifo_rx_pcs_data_out2_10g[69], w_hssi_fifo_rx_pcs_data_out2_10g[68], w_hssi_fifo_rx_pcs_data_out2_10g[67], w_hssi_fifo_rx_pcs_data_out2_10g[66], w_hssi_fifo_rx_pcs_data_out2_10g[65], w_hssi_fifo_rx_pcs_data_out2_10g[64], w_hssi_fifo_rx_pcs_data_out2_10g[63], w_hssi_fifo_rx_pcs_data_out2_10g[62], w_hssi_fifo_rx_pcs_data_out2_10g[61], w_hssi_fifo_rx_pcs_data_out2_10g[60], w_hssi_fifo_rx_pcs_data_out2_10g[59], w_hssi_fifo_rx_pcs_data_out2_10g[58], w_hssi_fifo_rx_pcs_data_out2_10g[57], w_hssi_fifo_rx_pcs_data_out2_10g[56], w_hssi_fifo_rx_pcs_data_out2_10g[55], w_hssi_fifo_rx_pcs_data_out2_10g[54], w_hssi_fifo_rx_pcs_data_out2_10g[53], w_hssi_fifo_rx_pcs_data_out2_10g[52], w_hssi_fifo_rx_pcs_data_out2_10g[51], w_hssi_fifo_rx_pcs_data_out2_10g[50], w_hssi_fifo_rx_pcs_data_out2_10g[49], w_hssi_fifo_rx_pcs_data_out2_10g[48], w_hssi_fifo_rx_pcs_data_out2_10g[47], w_hssi_fifo_rx_pcs_data_out2_10g[46], w_hssi_fifo_rx_pcs_data_out2_10g[45], w_hssi_fifo_rx_pcs_data_out2_10g[44], w_hssi_fifo_rx_pcs_data_out2_10g[43], w_hssi_fifo_rx_pcs_data_out2_10g[42], w_hssi_fifo_rx_pcs_data_out2_10g[41], w_hssi_fifo_rx_pcs_data_out2_10g[40], w_hssi_fifo_rx_pcs_data_out2_10g[39], w_hssi_fifo_rx_pcs_data_out2_10g[38], w_hssi_fifo_rx_pcs_data_out2_10g[37], w_hssi_fifo_rx_pcs_data_out2_10g[36], w_hssi_fifo_rx_pcs_data_out2_10g[35], w_hssi_fifo_rx_pcs_data_out2_10g[34], w_hssi_fifo_rx_pcs_data_out2_10g[33], w_hssi_fifo_rx_pcs_data_out2_10g[32], w_hssi_fifo_rx_pcs_data_out2_10g[31], w_hssi_fifo_rx_pcs_data_out2_10g[30], w_hssi_fifo_rx_pcs_data_out2_10g[29], w_hssi_fifo_rx_pcs_data_out2_10g[28], w_hssi_fifo_rx_pcs_data_out2_10g[27], w_hssi_fifo_rx_pcs_data_out2_10g[26], w_hssi_fifo_rx_pcs_data_out2_10g[25], w_hssi_fifo_rx_pcs_data_out2_10g[24], w_hssi_fifo_rx_pcs_data_out2_10g[23], w_hssi_fifo_rx_pcs_data_out2_10g[22], w_hssi_fifo_rx_pcs_data_out2_10g[21], w_hssi_fifo_rx_pcs_data_out2_10g[20], w_hssi_fifo_rx_pcs_data_out2_10g[19], w_hssi_fifo_rx_pcs_data_out2_10g[18], w_hssi_fifo_rx_pcs_data_out2_10g[17], w_hssi_fifo_rx_pcs_data_out2_10g[16], w_hssi_fifo_rx_pcs_data_out2_10g[15], w_hssi_fifo_rx_pcs_data_out2_10g[14], w_hssi_fifo_rx_pcs_data_out2_10g[13], w_hssi_fifo_rx_pcs_data_out2_10g[12], w_hssi_fifo_rx_pcs_data_out2_10g[11], w_hssi_fifo_rx_pcs_data_out2_10g[10], w_hssi_fifo_rx_pcs_data_out2_10g[9], w_hssi_fifo_rx_pcs_data_out2_10g[8], w_hssi_fifo_rx_pcs_data_out2_10g[7], w_hssi_fifo_rx_pcs_data_out2_10g[6], w_hssi_fifo_rx_pcs_data_out2_10g[5], w_hssi_fifo_rx_pcs_data_out2_10g[4], w_hssi_fifo_rx_pcs_data_out2_10g[3], w_hssi_fifo_rx_pcs_data_out2_10g[2], w_hssi_fifo_rx_pcs_data_out2_10g[1], w_hssi_fifo_rx_pcs_data_out2_10g[0]}),
				.rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.rx_pma_data({w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0]}),
				.rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.signal_ok_krfec(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_10g_reg(),
				.pld_10g_krfec_rx_blk_lock_10g_txclk_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_txclk_reg(),
				.pld_10g_krfec_rx_frame_10g_reg(),
				.pld_10g_krfec_rx_frame_10g_txclk_reg(),
				.pld_10g_krfec_rx_pld_rst_n_fifo(),
				.pld_10g_krfec_rx_pld_rst_n_reg(),
				.pld_10g_krfec_rx_pld_rst_n_txclk_reg(),
				.pld_10g_rx_align_clr_fifo(),
				.pld_10g_rx_align_clr_reg(),
				.pld_10g_rx_align_clr_txclk_reg(),
				.pld_10g_rx_align_val_fifo(),
				.pld_10g_rx_align_val_reg(),
				.pld_10g_rx_align_val_txclk_reg(),
				.pld_10g_rx_clr_ber_count_reg(),
				.pld_10g_rx_clr_ber_count_txclk_reg(),
				.pld_10g_rx_crc32_err_reg(),
				.pld_10g_rx_crc32_err_txclk_reg(),
				.pld_10g_rx_data_valid_10g_reg(),
				.pld_10g_rx_data_valid_fifo(),
				.pld_10g_rx_data_valid_pcsdirect_reg(),
				.pld_10g_rx_data_valid_txclk_reg(),
				.pld_10g_rx_empty_fifo(),
				.pld_10g_rx_fifo_del_reg(),
				.pld_10g_rx_fifo_del_txclk_reg(),
				.pld_10g_rx_fifo_insert_fifo(),
				.pld_10g_rx_fifo_num_reg(),
				.pld_10g_rx_fifo_num_txclk_reg(),
				.pld_10g_rx_frame_lock_reg(),
				.pld_10g_rx_frame_lock_txclk_reg(),
				.pld_10g_rx_hi_ber_reg(),
				.pld_10g_rx_hi_ber_txclk_reg(),
				.pld_10g_rx_oflw_err_reg(),
				.pld_10g_rx_oflw_err_txclk_reg(),
				.pld_10g_rx_pempty_fifo(),
				.pld_10g_rx_pfull_reg(),
				.pld_10g_rx_pfull_txclk_reg(),
				.pld_10g_rx_rd_en_fifo(),
				.pld_pcs_rx_clk_out_10g_txclk_wire(),
				.pld_pcs_rx_clk_out_10g_wire(),
				.pld_rx_control_10g_reg(),
				.pld_rx_control_10g_txclk_reg(),
				.pld_rx_data_10g_reg(),
				.pld_rx_data_10g_txclk_reg(),
				.pld_rx_prbs_err_10g_txclk_reg(),
				.pld_rx_prbs_err_clr_10g_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_10g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_align_val = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_blk_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_control[19:0] = 20'b0;
				assign w_hssi_10g_rx_pcs_rx_crc32_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_data[127:0] = 128'b0;
				assign w_hssi_10g_rx_pcs_rx_data_valid = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_dft_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_diag_status[1:0] = 2'b0;
				assign w_hssi_10g_rx_pcs_rx_empty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fec_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_del = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_insert = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_data[73:0] = 74'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_frame_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_hi_ber = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_oflw_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pempty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pfull = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_random_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_rx_frame = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_10g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_tx_pcs
			twentynm_hssi_10g_tx_pcs #(
				.advanced_user_mode(hssi_10g_tx_pcs_advanced_user_mode),
				.bitslip_en(hssi_10g_tx_pcs_bitslip_en),
				.bonding_dft_en(hssi_10g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_10g_tx_pcs_bonding_dft_val),
				.comp_cnt(hssi_10g_tx_pcs_comp_cnt),
				.compin_sel(hssi_10g_tx_pcs_compin_sel),
				.crcgen_bypass(hssi_10g_tx_pcs_crcgen_bypass),
				.crcgen_clken(hssi_10g_tx_pcs_crcgen_clken),
				.crcgen_err(hssi_10g_tx_pcs_crcgen_err),
				.crcgen_inv(hssi_10g_tx_pcs_crcgen_inv),
				.ctrl_bit_reverse(hssi_10g_tx_pcs_ctrl_bit_reverse),
				.ctrl_plane_bonding(hssi_10g_tx_pcs_ctrl_plane_bonding),
				.data_bit_reverse(hssi_10g_tx_pcs_data_bit_reverse),
				.dft_clk_out_sel(hssi_10g_tx_pcs_dft_clk_out_sel),
				.dispgen_bypass(hssi_10g_tx_pcs_dispgen_bypass),
				.dispgen_clken(hssi_10g_tx_pcs_dispgen_clken),
				.dispgen_err(hssi_10g_tx_pcs_dispgen_err),
				.dispgen_pipeln(hssi_10g_tx_pcs_dispgen_pipeln),
				.distdwn_bypass_pipeln(hssi_10g_tx_pcs_distdwn_bypass_pipeln),
				.distdwn_master(hssi_10g_tx_pcs_distdwn_master),
				.distup_bypass_pipeln(hssi_10g_tx_pcs_distup_bypass_pipeln),
				.distup_master(hssi_10g_tx_pcs_distup_master),
				.dv_bond(hssi_10g_tx_pcs_dv_bond),
				.empty_flag_type(hssi_10g_tx_pcs_empty_flag_type),
				.enc64b66b_txsm_clken(hssi_10g_tx_pcs_enc64b66b_txsm_clken),
				.enc_64b66b_txsm_bypass(hssi_10g_tx_pcs_enc_64b66b_txsm_bypass),
				.fastpath(hssi_10g_tx_pcs_fastpath),
				.fec_clken(hssi_10g_tx_pcs_fec_clken),
				.fec_enable(hssi_10g_tx_pcs_fec_enable),
				.fifo_double_write(hssi_10g_tx_pcs_fifo_double_write),
				.fifo_reg_fast(hssi_10g_tx_pcs_fifo_reg_fast),
				.fifo_stop_rd(hssi_10g_tx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_tx_pcs_fifo_stop_wr),
				.frmgen_burst(hssi_10g_tx_pcs_frmgen_burst),
				.frmgen_bypass(hssi_10g_tx_pcs_frmgen_bypass),
				.frmgen_clken(hssi_10g_tx_pcs_frmgen_clken),
				.frmgen_mfrm_length(hssi_10g_tx_pcs_frmgen_mfrm_length),
				.frmgen_pipeln(hssi_10g_tx_pcs_frmgen_pipeln),
				.frmgen_pyld_ins(hssi_10g_tx_pcs_frmgen_pyld_ins),
				.frmgen_wordslip(hssi_10g_tx_pcs_frmgen_wordslip),
				.full_flag_type(hssi_10g_tx_pcs_full_flag_type),
				.gb_pipeln_bypass(hssi_10g_tx_pcs_gb_pipeln_bypass),
				.gb_tx_idwidth(hssi_10g_tx_pcs_gb_tx_idwidth),
				.gb_tx_odwidth(hssi_10g_tx_pcs_gb_tx_odwidth),
				.gbred_clken(hssi_10g_tx_pcs_gbred_clken),
				.indv(hssi_10g_tx_pcs_indv),
				.low_latency_en(hssi_10g_tx_pcs_low_latency_en),
				.master_clk_sel(hssi_10g_tx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_tx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_tx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_tx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_tx_pcs_pld_if_type),
				.prot_mode(hssi_10g_tx_pcs_prot_mode),
				.pseudo_random(hssi_10g_tx_pcs_pseudo_random),
				.pseudo_seed_a(hssi_10g_tx_pcs_pseudo_seed_a),
				.pseudo_seed_b(hssi_10g_tx_pcs_pseudo_seed_b),
				.random_disp(hssi_10g_tx_pcs_random_disp),
				.rdfifo_clken(hssi_10g_tx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_tx_pcs_reconfig_settings),
				.scrm_bypass(hssi_10g_tx_pcs_scrm_bypass),
				.scrm_clken(hssi_10g_tx_pcs_scrm_clken),
				.scrm_mode(hssi_10g_tx_pcs_scrm_mode),
				.scrm_pipeln(hssi_10g_tx_pcs_scrm_pipeln),
				.sh_err(hssi_10g_tx_pcs_sh_err),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sop_mark(hssi_10g_tx_pcs_sop_mark),
				.stretch_num_stages(hssi_10g_tx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_tx_pcs_sup_mode),
				.test_mode(hssi_10g_tx_pcs_test_mode),
				.tx_scrm_err(hssi_10g_tx_pcs_tx_scrm_err),
				.tx_scrm_width(hssi_10g_tx_pcs_tx_scrm_width),
				.tx_sh_location(hssi_10g_tx_pcs_tx_sh_location),
				.tx_sm_bypass(hssi_10g_tx_pcs_tx_sm_bypass),
				.tx_sm_pipeln(hssi_10g_tx_pcs_tx_sm_pipeln),
				.tx_testbus_sel(hssi_10g_tx_pcs_tx_testbus_sel),
				.txfifo_empty(hssi_10g_tx_pcs_txfifo_empty),
				.txfifo_full(hssi_10g_tx_pcs_txfifo_full),
				.txfifo_mode(hssi_10g_tx_pcs_txfifo_mode),
				.txfifo_pempty(hssi_10g_tx_pcs_txfifo_pempty),
				.txfifo_pfull(hssi_10g_tx_pcs_txfifo_pfull),
				.wr_clk_sel(hssi_10g_tx_pcs_wr_clk_sel),
				.wrfifo_clken(hssi_10g_tx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_tx_pcs_blockselect),
				.distdwn_out_dv(w_hssi_10g_tx_pcs_distdwn_out_dv),
				.distdwn_out_rden(w_hssi_10g_tx_pcs_distdwn_out_rden),
				.distdwn_out_wren(w_hssi_10g_tx_pcs_distdwn_out_wren),
				.distup_out_dv(w_hssi_10g_tx_pcs_distup_out_dv),
				.distup_out_rden(w_hssi_10g_tx_pcs_distup_out_rden),
				.distup_out_wren(w_hssi_10g_tx_pcs_distup_out_wren),
				.tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pma_if(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.tx_control_out_krfec(w_hssi_10g_tx_pcs_tx_control_out_krfec),
				.tx_data_out_krfec(w_hssi_10g_tx_pcs_tx_data_out_krfec),
				.tx_data_valid_out_krfec(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.tx_fec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_fifo_num(w_hssi_10g_tx_pcs_tx_fifo_num),
				.tx_fifo_rd_ptr(w_hssi_10g_tx_pcs_tx_fifo_rd_ptr),
				.tx_fifo_wr_clk(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.tx_fifo_wr_data(w_hssi_10g_tx_pcs_tx_fifo_wr_data),
				.tx_fifo_wr_data_dw(w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw),
				.tx_fifo_wr_en(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.tx_fifo_wr_ptr(w_hssi_10g_tx_pcs_tx_fifo_wr_ptr),
				.tx_fifo_wr_rst_n(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.tx_full(w_hssi_10g_tx_pcs_tx_full),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				.tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.tx_pma_data(w_hssi_10g_tx_pcs_tx_pma_data),
				.tx_pma_gating_val(w_hssi_10g_tx_pcs_tx_pma_gating_val),
				.tx_test_data(w_hssi_10g_tx_pcs_tx_test_data),
				.tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.distdwn_in_dv(in_bond_pcs10g_in_bot[2]),
				.distdwn_in_rden(in_bond_pcs10g_in_bot[4]),
				.distdwn_in_wren(in_bond_pcs10g_in_bot[3]),
				.distup_in_dv(in_bond_pcs10g_in_top[2]),
				.distup_in_rden(in_bond_pcs10g_in_top[4]),
				.distup_in_wren(in_bond_pcs10g_in_top[3]),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_tx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_tx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.tx_bitslip({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0]}),
				.tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.tx_control({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0]}),
				.tx_control_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0]}),
				.tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0]}),
				.tx_data_in_krfec({w_hssi_krfec_tx_pcs_tx_data_out[63], w_hssi_krfec_tx_pcs_tx_data_out[62], w_hssi_krfec_tx_pcs_tx_data_out[61], w_hssi_krfec_tx_pcs_tx_data_out[60], w_hssi_krfec_tx_pcs_tx_data_out[59], w_hssi_krfec_tx_pcs_tx_data_out[58], w_hssi_krfec_tx_pcs_tx_data_out[57], w_hssi_krfec_tx_pcs_tx_data_out[56], w_hssi_krfec_tx_pcs_tx_data_out[55], w_hssi_krfec_tx_pcs_tx_data_out[54], w_hssi_krfec_tx_pcs_tx_data_out[53], w_hssi_krfec_tx_pcs_tx_data_out[52], w_hssi_krfec_tx_pcs_tx_data_out[51], w_hssi_krfec_tx_pcs_tx_data_out[50], w_hssi_krfec_tx_pcs_tx_data_out[49], w_hssi_krfec_tx_pcs_tx_data_out[48], w_hssi_krfec_tx_pcs_tx_data_out[47], w_hssi_krfec_tx_pcs_tx_data_out[46], w_hssi_krfec_tx_pcs_tx_data_out[45], w_hssi_krfec_tx_pcs_tx_data_out[44], w_hssi_krfec_tx_pcs_tx_data_out[43], w_hssi_krfec_tx_pcs_tx_data_out[42], w_hssi_krfec_tx_pcs_tx_data_out[41], w_hssi_krfec_tx_pcs_tx_data_out[40], w_hssi_krfec_tx_pcs_tx_data_out[39], w_hssi_krfec_tx_pcs_tx_data_out[38], w_hssi_krfec_tx_pcs_tx_data_out[37], w_hssi_krfec_tx_pcs_tx_data_out[36], w_hssi_krfec_tx_pcs_tx_data_out[35], w_hssi_krfec_tx_pcs_tx_data_out[34], w_hssi_krfec_tx_pcs_tx_data_out[33], w_hssi_krfec_tx_pcs_tx_data_out[32], w_hssi_krfec_tx_pcs_tx_data_out[31], w_hssi_krfec_tx_pcs_tx_data_out[30], w_hssi_krfec_tx_pcs_tx_data_out[29], w_hssi_krfec_tx_pcs_tx_data_out[28], w_hssi_krfec_tx_pcs_tx_data_out[27], w_hssi_krfec_tx_pcs_tx_data_out[26], w_hssi_krfec_tx_pcs_tx_data_out[25], w_hssi_krfec_tx_pcs_tx_data_out[24], w_hssi_krfec_tx_pcs_tx_data_out[23], w_hssi_krfec_tx_pcs_tx_data_out[22], w_hssi_krfec_tx_pcs_tx_data_out[21], w_hssi_krfec_tx_pcs_tx_data_out[20], w_hssi_krfec_tx_pcs_tx_data_out[19], w_hssi_krfec_tx_pcs_tx_data_out[18], w_hssi_krfec_tx_pcs_tx_data_out[17], w_hssi_krfec_tx_pcs_tx_data_out[16], w_hssi_krfec_tx_pcs_tx_data_out[15], w_hssi_krfec_tx_pcs_tx_data_out[14], w_hssi_krfec_tx_pcs_tx_data_out[13], w_hssi_krfec_tx_pcs_tx_data_out[12], w_hssi_krfec_tx_pcs_tx_data_out[11], w_hssi_krfec_tx_pcs_tx_data_out[10], w_hssi_krfec_tx_pcs_tx_data_out[9], w_hssi_krfec_tx_pcs_tx_data_out[8], w_hssi_krfec_tx_pcs_tx_data_out[7], w_hssi_krfec_tx_pcs_tx_data_out[6], w_hssi_krfec_tx_pcs_tx_data_out[5], w_hssi_krfec_tx_pcs_tx_data_out[4], w_hssi_krfec_tx_pcs_tx_data_out[3], w_hssi_krfec_tx_pcs_tx_data_out[2], w_hssi_krfec_tx_pcs_tx_data_out[1], w_hssi_krfec_tx_pcs_tx_data_out[0]}),
				.tx_data_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0]}),
				.tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.tx_diag_status({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0]}),
				.tx_fifo_rd_data({w_hssi_fifo_tx_pcs_data_out_10g[72], w_hssi_fifo_tx_pcs_data_out_10g[71], w_hssi_fifo_tx_pcs_data_out_10g[70], w_hssi_fifo_tx_pcs_data_out_10g[69], w_hssi_fifo_tx_pcs_data_out_10g[68], w_hssi_fifo_tx_pcs_data_out_10g[67], w_hssi_fifo_tx_pcs_data_out_10g[66], w_hssi_fifo_tx_pcs_data_out_10g[65], w_hssi_fifo_tx_pcs_data_out_10g[64], w_hssi_fifo_tx_pcs_data_out_10g[63], w_hssi_fifo_tx_pcs_data_out_10g[62], w_hssi_fifo_tx_pcs_data_out_10g[61], w_hssi_fifo_tx_pcs_data_out_10g[60], w_hssi_fifo_tx_pcs_data_out_10g[59], w_hssi_fifo_tx_pcs_data_out_10g[58], w_hssi_fifo_tx_pcs_data_out_10g[57], w_hssi_fifo_tx_pcs_data_out_10g[56], w_hssi_fifo_tx_pcs_data_out_10g[55], w_hssi_fifo_tx_pcs_data_out_10g[54], w_hssi_fifo_tx_pcs_data_out_10g[53], w_hssi_fifo_tx_pcs_data_out_10g[52], w_hssi_fifo_tx_pcs_data_out_10g[51], w_hssi_fifo_tx_pcs_data_out_10g[50], w_hssi_fifo_tx_pcs_data_out_10g[49], w_hssi_fifo_tx_pcs_data_out_10g[48], w_hssi_fifo_tx_pcs_data_out_10g[47], w_hssi_fifo_tx_pcs_data_out_10g[46], w_hssi_fifo_tx_pcs_data_out_10g[45], w_hssi_fifo_tx_pcs_data_out_10g[44], w_hssi_fifo_tx_pcs_data_out_10g[43], w_hssi_fifo_tx_pcs_data_out_10g[42], w_hssi_fifo_tx_pcs_data_out_10g[41], w_hssi_fifo_tx_pcs_data_out_10g[40], w_hssi_fifo_tx_pcs_data_out_10g[39], w_hssi_fifo_tx_pcs_data_out_10g[38], w_hssi_fifo_tx_pcs_data_out_10g[37], w_hssi_fifo_tx_pcs_data_out_10g[36], w_hssi_fifo_tx_pcs_data_out_10g[35], w_hssi_fifo_tx_pcs_data_out_10g[34], w_hssi_fifo_tx_pcs_data_out_10g[33], w_hssi_fifo_tx_pcs_data_out_10g[32], w_hssi_fifo_tx_pcs_data_out_10g[31], w_hssi_fifo_tx_pcs_data_out_10g[30], w_hssi_fifo_tx_pcs_data_out_10g[29], w_hssi_fifo_tx_pcs_data_out_10g[28], w_hssi_fifo_tx_pcs_data_out_10g[27], w_hssi_fifo_tx_pcs_data_out_10g[26], w_hssi_fifo_tx_pcs_data_out_10g[25], w_hssi_fifo_tx_pcs_data_out_10g[24], w_hssi_fifo_tx_pcs_data_out_10g[23], w_hssi_fifo_tx_pcs_data_out_10g[22], w_hssi_fifo_tx_pcs_data_out_10g[21], w_hssi_fifo_tx_pcs_data_out_10g[20], w_hssi_fifo_tx_pcs_data_out_10g[19], w_hssi_fifo_tx_pcs_data_out_10g[18], w_hssi_fifo_tx_pcs_data_out_10g[17], w_hssi_fifo_tx_pcs_data_out_10g[16], w_hssi_fifo_tx_pcs_data_out_10g[15], w_hssi_fifo_tx_pcs_data_out_10g[14], w_hssi_fifo_tx_pcs_data_out_10g[13], w_hssi_fifo_tx_pcs_data_out_10g[12], w_hssi_fifo_tx_pcs_data_out_10g[11], w_hssi_fifo_tx_pcs_data_out_10g[10], w_hssi_fifo_tx_pcs_data_out_10g[9], w_hssi_fifo_tx_pcs_data_out_10g[8], w_hssi_fifo_tx_pcs_data_out_10g[7], w_hssi_fifo_tx_pcs_data_out_10g[6], w_hssi_fifo_tx_pcs_data_out_10g[5], w_hssi_fifo_tx_pcs_data_out_10g[4], w_hssi_fifo_tx_pcs_data_out_10g[3], w_hssi_fifo_tx_pcs_data_out_10g[2], w_hssi_fifo_tx_pcs_data_out_10g[1], w_hssi_fifo_tx_pcs_data_out_10g[0]}),
				.tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_10g_reg(),
				.pld_10g_krfec_tx_pld_rst_n_fifo(),
				.pld_10g_krfec_tx_pld_rst_n_reg(),
				.pld_10g_tx_bitslip_reg(),
				.pld_10g_tx_burst_en_exe_reg(),
				.pld_10g_tx_data_valid_10g_reg(),
				.pld_10g_tx_data_valid_fifo(),
				.pld_10g_tx_data_valid_reg(),
				.pld_10g_tx_diag_status_reg(),
				.pld_10g_tx_empty_reg(),
				.pld_10g_tx_fifo_num_reg(),
				.pld_10g_tx_full_fifo(),
				.pld_10g_tx_full_reg(),
				.pld_10g_tx_pempty_reg(),
				.pld_10g_tx_pfull_fifo(),
				.pld_10g_tx_wordslip_exe_reg(),
				.pld_10g_tx_wordslip_reg(),
				.pld_pcs_tx_clk_out_10g_wire(),
				.pld_tx_burst_en_reg(),
				.pld_tx_control_lo_10g_reg(),
				.pld_tx_data_10g_fifo(),
				.pld_tx_data_lo_10g_reg()
			);
		end // if generate
		else begin
				assign w_hssi_10g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_burst_en_exe = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pma_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_control_out_krfec[8:0] = 9'b0;
				assign w_hssi_10g_tx_pcs_tx_data_out_krfec[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_data_valid_out_krfec = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_dft_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_empty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fec_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_full = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_pempty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pfull = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_gating_val[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_test_data[19:0] = 20'b0;
				assign w_hssi_10g_tx_pcs_tx_wordslip_exe = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_rx_pcs
			twentynm_hssi_8g_rx_pcs #(
				.auto_error_replacement(hssi_8g_rx_pcs_auto_error_replacement),
				.auto_speed_nego(hssi_8g_rx_pcs_auto_speed_nego),
				.bit_reversal(hssi_8g_rx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_rx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_rx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_rx_pcs_bypass_pipeline_reg),
				.byte_deserializer(hssi_8g_rx_pcs_byte_deserializer),
				.cdr_ctrl_rxvalid_mask(hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask),
				.clkcmp_pattern_n(hssi_8g_rx_pcs_clkcmp_pattern_n),
				.clkcmp_pattern_p(hssi_8g_rx_pcs_clkcmp_pattern_p),
				.clock_gate_bds_dec_asn(hssi_8g_rx_pcs_clock_gate_bds_dec_asn),
				.clock_gate_cdr_eidle(hssi_8g_rx_pcs_clock_gate_cdr_eidle),
				.clock_gate_dw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk),
				.clock_gate_dw_rm_rd(hssi_8g_rx_pcs_clock_gate_dw_rm_rd),
				.clock_gate_dw_rm_wr(hssi_8g_rx_pcs_clock_gate_dw_rm_wr),
				.clock_gate_dw_wa(hssi_8g_rx_pcs_clock_gate_dw_wa),
				.clock_gate_pc_rdclk(hssi_8g_rx_pcs_clock_gate_pc_rdclk),
				.clock_gate_sw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk),
				.clock_gate_sw_rm_rd(hssi_8g_rx_pcs_clock_gate_sw_rm_rd),
				.clock_gate_sw_rm_wr(hssi_8g_rx_pcs_clock_gate_sw_rm_wr),
				.clock_gate_sw_wa(hssi_8g_rx_pcs_clock_gate_sw_wa),
				.clock_observation_in_pld_core(hssi_8g_rx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_rx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_rx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_rx_pcs_ctrl_plane_bonding_distribution),
				.eidle_entry_eios(hssi_8g_rx_pcs_eidle_entry_eios),
				.eidle_entry_iei(hssi_8g_rx_pcs_eidle_entry_iei),
				.eidle_entry_sd(hssi_8g_rx_pcs_eidle_entry_sd),
				.eightb_tenb_decoder(hssi_8g_rx_pcs_eightb_tenb_decoder),
				.err_flags_sel(hssi_8g_rx_pcs_err_flags_sel),
				.fixed_pat_det(hssi_8g_rx_pcs_fixed_pat_det),
				.fixed_pat_num(hssi_8g_rx_pcs_fixed_pat_num),
				.force_signal_detect(hssi_8g_rx_pcs_force_signal_detect),
				.gen3_clk_en(hssi_8g_rx_pcs_gen3_clk_en),
				.gen3_rx_clk_sel(hssi_8g_rx_pcs_gen3_rx_clk_sel),
				.gen3_tx_clk_sel(hssi_8g_rx_pcs_gen3_tx_clk_sel),
				.hip_mode(hssi_8g_rx_pcs_hip_mode),
				.ibm_invalid_code(hssi_8g_rx_pcs_ibm_invalid_code),
				.invalid_code_flag_only(hssi_8g_rx_pcs_invalid_code_flag_only),
				.pad_or_edb_error_replace(hssi_8g_rx_pcs_pad_or_edb_error_replace),
				.pcs_bypass(hssi_8g_rx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_rx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_rx_pcs_phase_compensation_fifo),
				.pipe_if_enable(hssi_8g_rx_pcs_pipe_if_enable),
				.pma_dw(hssi_8g_rx_pcs_pma_dw),
				.polinv_8b10b_dec(hssi_8g_rx_pcs_polinv_8b10b_dec),
				.prot_mode(hssi_8g_rx_pcs_prot_mode),
				.rate_match(hssi_8g_rx_pcs_rate_match),
				.rate_match_del_thres(hssi_8g_rx_pcs_rate_match_del_thres),
				.rate_match_empty_thres(hssi_8g_rx_pcs_rate_match_empty_thres),
				.rate_match_full_thres(hssi_8g_rx_pcs_rate_match_full_thres),
				.rate_match_ins_thres(hssi_8g_rx_pcs_rate_match_ins_thres),
				.rate_match_start_thres(hssi_8g_rx_pcs_rate_match_start_thres),
				.reconfig_settings(hssi_8g_rx_pcs_reconfig_settings),
				.rx_clk2(hssi_8g_rx_pcs_rx_clk2),
				.rx_clk_free_running(hssi_8g_rx_pcs_rx_clk_free_running),
				.rx_pcs_urst(hssi_8g_rx_pcs_rx_pcs_urst),
				.rx_rcvd_clk(hssi_8g_rx_pcs_rx_rcvd_clk),
				.rx_rd_clk(hssi_8g_rx_pcs_rx_rd_clk),
				.rx_refclk(hssi_8g_rx_pcs_rx_refclk),
				.rx_wr_clk(hssi_8g_rx_pcs_rx_wr_clk),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_rx_pcs_sup_mode),
				.symbol_swap(hssi_8g_rx_pcs_symbol_swap),
				.sync_sm_idle_eios(hssi_8g_rx_pcs_sync_sm_idle_eios),
				.test_bus_sel(hssi_8g_rx_pcs_test_bus_sel),
				.tx_rx_parallel_loopback(hssi_8g_rx_pcs_tx_rx_parallel_loopback),
				.wa_boundary_lock_ctrl(hssi_8g_rx_pcs_wa_boundary_lock_ctrl),
				.wa_clk_slip_spacing(hssi_8g_rx_pcs_wa_clk_slip_spacing),
				.wa_det_latency_sync_status_beh(hssi_8g_rx_pcs_wa_det_latency_sync_status_beh),
				.wa_disp_err_flag(hssi_8g_rx_pcs_wa_disp_err_flag),
				.wa_kchar(hssi_8g_rx_pcs_wa_kchar),
				.wa_pd(hssi_8g_rx_pcs_wa_pd),
				.wa_pd_data(hssi_8g_rx_pcs_wa_pd_data),
				.wa_pd_polarity(hssi_8g_rx_pcs_wa_pd_polarity),
				.wa_pld_controlled(hssi_8g_rx_pcs_wa_pld_controlled),
				.wa_renumber_data(hssi_8g_rx_pcs_wa_renumber_data),
				.wa_rgnumber_data(hssi_8g_rx_pcs_wa_rgnumber_data),
				.wa_rknumber_data(hssi_8g_rx_pcs_wa_rknumber_data),
				.wa_rosnumber_data(hssi_8g_rx_pcs_wa_rosnumber_data),
				.wa_rvnumber_data(hssi_8g_rx_pcs_wa_rvnumber_data),
				.wa_sync_sm_ctrl(hssi_8g_rx_pcs_wa_sync_sm_ctrl),
				.wait_cnt(hssi_8g_rx_pcs_wait_cnt)
			) inst_twentynm_hssi_8g_rx_pcs (
				// OUTPUTS
				.a1a2k1k2flag(w_hssi_8g_rx_pcs_a1a2k1k2flag),
				.avmmreaddata(w_hssi_8g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_rx_pcs_blockselect),
				.chnl_test_bus_out(w_hssi_8g_rx_pcs_chnl_test_bus_out),
				.clock_to_pld(w_hssi_8g_rx_pcs_clock_to_pld),
				.dataout(w_hssi_8g_rx_pcs_dataout),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidle_detected(w_hssi_8g_rx_pcs_eidle_detected),
				.eios_det_cdr_ctrl(w_hssi_8g_rx_pcs_eios_det_cdr_ctrl),
				.g3_rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.g3_rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.gen2ngen1(w_hssi_8g_rx_pcs_gen2ngen1),
				.parallel_rev_loopback(w_hssi_8g_rx_pcs_parallel_rev_loopback),
				.pc_fifo_empty(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.pcfifofull(w_hssi_8g_rx_pcs_pcfifofull),
				.phystatus(w_hssi_8g_rx_pcs_phystatus),
				.pipe_data(w_hssi_8g_rx_pcs_pipe_data),
				.rd_enable_out_chnl_down(w_hssi_8g_rx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_rx_pcs_rd_enable_out_chnl_up),
				.rd_ptr1_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo),
				.rd_ptr2_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo),
				.rd_ptr_rx_phfifo(w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.reset_pc_ptrs_out_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down),
				.reset_pc_ptrs_out_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up),
				.rm_fifo_empty(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.rm_fifo_full(w_hssi_8g_rx_pcs_rm_fifo_full),
				.rx_blk_start(w_hssi_8g_rx_pcs_rx_blk_start),
				.rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.rx_data_valid(w_hssi_8g_rx_pcs_rx_data_valid),
				.rx_div_sync_out_chnl_down(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down),
				.rx_div_sync_out_chnl_up(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up),
				.rx_pipe_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.rx_pipe_soft_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rx_pma_clk_gen3(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_rcvd_clk_gen3(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_rstn_sync2wrfifo_8g(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.rx_sync_hdr(w_hssi_8g_rx_pcs_rx_sync_hdr),
				.rx_we_out_chnl_down(w_hssi_8g_rx_pcs_rx_we_out_chnl_down),
				.rx_we_out_chnl_up(w_hssi_8g_rx_pcs_rx_we_out_chnl_up),
				.rxstatus(w_hssi_8g_rx_pcs_rxstatus),
				.rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.word_align_boundary(w_hssi_8g_rx_pcs_word_align_boundary),
				.wr_clk_rx_phfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_rx_phfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_rx_rmfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_rx_rmfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_data_rx_phfifo(w_hssi_8g_rx_pcs_wr_data_rx_phfifo),
				.wr_data_rx_rmfifo(w_hssi_8g_rx_pcs_wr_data_rx_rmfifo),
				.wr_en_rx_phfifo(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_rx_rmfifo(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_rx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_rx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_rx_phfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo),
				.wr_ptr_rx_rmfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo),
				.wr_rst_n_rx_phfifo(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_rx_rmfifo(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				// INPUTS
				.a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bit_reversal_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.datain({w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0]}),
				.disable_pc_fifo_byte_serdes(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4]),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.eidleinfersel({w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0]}),
				.eios_detected_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.enable_comma_detect(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.gen3_clk_sel(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.hrd_rst(1'b0),
				.inferred_rxvalid_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.pc_fifo_rd_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.pc_fifo_wrdisable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.phystatus_int(w_hssi_pipe_gen1_2_phystatus),
				.phystatus_pcs_gen3(w_hssi_pipe_gen3_phystatus),
				.pipe_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.polarity_inversion(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.rd_data1_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0]}),
				.rd_data2_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0]}),
				.rd_data_rx_phfifo({w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[3]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[3]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.reset_pc_ptrs_asn(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5]),
				.reset_pc_ptrs_in_chnl_down(in_bond_pcs8g_in_bot[12]),
				.reset_pc_ptrs_in_chnl_up(in_bond_pcs8g_in_top[12]),
				.reset_ppm_cntrs_pcs_pma(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7]),
				.rm_fifo_read_enable(1'b0),
				.rm_fifo_write_enable(1'b0),
				.rx_blk_start_pcs_gen3({w_hssi_pipe_gen3_rx_blk_start[3], w_hssi_pipe_gen3_rx_blk_start[2], w_hssi_pipe_gen3_rx_blk_start[1], w_hssi_pipe_gen3_rx_blk_start[0]}),
				.rx_data_pcs_gen3({w_hssi_pipe_gen3_rxd_8gpcs_out[63], w_hssi_pipe_gen3_rxd_8gpcs_out[62], w_hssi_pipe_gen3_rxd_8gpcs_out[61], w_hssi_pipe_gen3_rxd_8gpcs_out[60], w_hssi_pipe_gen3_rxd_8gpcs_out[59], w_hssi_pipe_gen3_rxd_8gpcs_out[58], w_hssi_pipe_gen3_rxd_8gpcs_out[57], w_hssi_pipe_gen3_rxd_8gpcs_out[56], w_hssi_pipe_gen3_rxd_8gpcs_out[55], w_hssi_pipe_gen3_rxd_8gpcs_out[54], w_hssi_pipe_gen3_rxd_8gpcs_out[53], w_hssi_pipe_gen3_rxd_8gpcs_out[52], w_hssi_pipe_gen3_rxd_8gpcs_out[51], w_hssi_pipe_gen3_rxd_8gpcs_out[50], w_hssi_pipe_gen3_rxd_8gpcs_out[49], w_hssi_pipe_gen3_rxd_8gpcs_out[48], w_hssi_pipe_gen3_rxd_8gpcs_out[47], w_hssi_pipe_gen3_rxd_8gpcs_out[46], w_hssi_pipe_gen3_rxd_8gpcs_out[45], w_hssi_pipe_gen3_rxd_8gpcs_out[44], w_hssi_pipe_gen3_rxd_8gpcs_out[43], w_hssi_pipe_gen3_rxd_8gpcs_out[42], w_hssi_pipe_gen3_rxd_8gpcs_out[41], w_hssi_pipe_gen3_rxd_8gpcs_out[40], w_hssi_pipe_gen3_rxd_8gpcs_out[39], w_hssi_pipe_gen3_rxd_8gpcs_out[38], w_hssi_pipe_gen3_rxd_8gpcs_out[37], w_hssi_pipe_gen3_rxd_8gpcs_out[36], w_hssi_pipe_gen3_rxd_8gpcs_out[35], w_hssi_pipe_gen3_rxd_8gpcs_out[34], w_hssi_pipe_gen3_rxd_8gpcs_out[33], w_hssi_pipe_gen3_rxd_8gpcs_out[32], w_hssi_pipe_gen3_rxd_8gpcs_out[31], w_hssi_pipe_gen3_rxd_8gpcs_out[30], w_hssi_pipe_gen3_rxd_8gpcs_out[29], w_hssi_pipe_gen3_rxd_8gpcs_out[28], w_hssi_pipe_gen3_rxd_8gpcs_out[27], w_hssi_pipe_gen3_rxd_8gpcs_out[26], w_hssi_pipe_gen3_rxd_8gpcs_out[25], w_hssi_pipe_gen3_rxd_8gpcs_out[24], w_hssi_pipe_gen3_rxd_8gpcs_out[23], w_hssi_pipe_gen3_rxd_8gpcs_out[22], w_hssi_pipe_gen3_rxd_8gpcs_out[21], w_hssi_pipe_gen3_rxd_8gpcs_out[20], w_hssi_pipe_gen3_rxd_8gpcs_out[19], w_hssi_pipe_gen3_rxd_8gpcs_out[18], w_hssi_pipe_gen3_rxd_8gpcs_out[17], w_hssi_pipe_gen3_rxd_8gpcs_out[16], w_hssi_pipe_gen3_rxd_8gpcs_out[15], w_hssi_pipe_gen3_rxd_8gpcs_out[14], w_hssi_pipe_gen3_rxd_8gpcs_out[13], w_hssi_pipe_gen3_rxd_8gpcs_out[12], w_hssi_pipe_gen3_rxd_8gpcs_out[11], w_hssi_pipe_gen3_rxd_8gpcs_out[10], w_hssi_pipe_gen3_rxd_8gpcs_out[9], w_hssi_pipe_gen3_rxd_8gpcs_out[8], w_hssi_pipe_gen3_rxd_8gpcs_out[7], w_hssi_pipe_gen3_rxd_8gpcs_out[6], w_hssi_pipe_gen3_rxd_8gpcs_out[5], w_hssi_pipe_gen3_rxd_8gpcs_out[4], w_hssi_pipe_gen3_rxd_8gpcs_out[3], w_hssi_pipe_gen3_rxd_8gpcs_out[2], w_hssi_pipe_gen3_rxd_8gpcs_out[1], w_hssi_pipe_gen3_rxd_8gpcs_out[0]}),
				.rx_data_valid_pcs_gen3({w_hssi_pipe_gen3_rxdataskip[3], w_hssi_pipe_gen3_rxdataskip[2], w_hssi_pipe_gen3_rxdataskip[1], w_hssi_pipe_gen3_rxdataskip[0]}),
				.rx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[1], in_bond_pcs8g_in_bot[0]}),
				.rx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[1], in_bond_pcs8g_in_top[0]}),
				.rx_pcs_rst(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.rx_sync_hdr_pcs_gen3({w_hssi_pipe_gen3_rx_sync_hdr[1], w_hssi_pipe_gen3_rx_sync_hdr[0]}),
				.rx_we_in_chnl_down({in_bond_pcs8g_in_bot[5], in_bond_pcs8g_in_bot[4]}),
				.rx_we_in_chnl_up({in_bond_pcs8g_in_top[5], in_bond_pcs8g_in_top[4]}),
				.rxstatus_int({w_hssi_pipe_gen1_2_rxstatus[2], w_hssi_pipe_gen1_2_rxstatus[1], w_hssi_pipe_gen1_2_rxstatus[0]}),
				.rxstatus_pcs_gen3({w_hssi_pipe_gen3_rxstatus[2], w_hssi_pipe_gen3_rxstatus[1], w_hssi_pipe_gen3_rxstatus[0]}),
				.rxvalid_int(w_hssi_pipe_gen1_2_rxvalid),
				.rxvalid_pcs_gen3(w_hssi_pipe_gen3_rxvalid),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.sig_det_from_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_ctrlplane_testbus({w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0]}),
				.tx_div_sync({w_hssi_8g_tx_pcs_tx_div_sync[1], w_hssi_8g_tx_pcs_tx_div_sync[0]}),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.tx_testbus({w_hssi_8g_tx_pcs_tx_testbus[19], w_hssi_8g_tx_pcs_tx_testbus[18], w_hssi_8g_tx_pcs_tx_testbus[17], w_hssi_8g_tx_pcs_tx_testbus[16], w_hssi_8g_tx_pcs_tx_testbus[15], w_hssi_8g_tx_pcs_tx_testbus[14], w_hssi_8g_tx_pcs_tx_testbus[13], w_hssi_8g_tx_pcs_tx_testbus[12], w_hssi_8g_tx_pcs_tx_testbus[11], w_hssi_8g_tx_pcs_tx_testbus[10], w_hssi_8g_tx_pcs_tx_testbus[9], w_hssi_8g_tx_pcs_tx_testbus[8], w_hssi_8g_tx_pcs_tx_testbus[7], w_hssi_8g_tx_pcs_tx_testbus[6], w_hssi_8g_tx_pcs_tx_testbus[5], w_hssi_8g_tx_pcs_tx_testbus[4], w_hssi_8g_tx_pcs_tx_testbus[3], w_hssi_8g_tx_pcs_tx_testbus[2], w_hssi_8g_tx_pcs_tx_testbus[1], w_hssi_8g_tx_pcs_tx_testbus[0]}),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[2]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[2]),
				
				// UNUSED
				.byte_deserializer_pcs_clk_div_by_2_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_wire(),
				.byte_deserializer_pcs_clk_div_by_2_wire(),
				.byte_deserializer_pcs_clk_div_by_4_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_2_reg(),
				.byte_deserializer_pld_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_4_txclk_reg(),
				.pld_8g_a1a2_k1k2_flag_reg(),
				.pld_8g_a1a2_k1k2_flag_txclk_reg(),
				.pld_8g_a1a2_size_reg(),
				.pld_8g_a1a2_size_txclk_reg(),
				.pld_8g_bitloc_rev_en_reg(),
				.pld_8g_bitloc_rev_en_txclk_reg(),
				.pld_8g_byte_rev_en_reg(),
				.pld_8g_byte_rev_en_txclk_reg(),
				.pld_8g_elecidle_reg(),
				.pld_8g_empty_rmf_lowlatency_reg(),
				.pld_8g_empty_rmf_lowlatency_txclk_reg(),
				.pld_8g_empty_rmf_reg(),
				.pld_8g_empty_rmf_txclk_reg(),
				.pld_8g_empty_rx_fifo(),
				.pld_8g_empty_rx_reg(),
				.pld_8g_empty_rx_txclk_reg(),
				.pld_8g_encdt_reg(),
				.pld_8g_encdt_txclk_reg(),
				.pld_8g_full_rmf_reg(),
				.pld_8g_full_rmf_txclk_reg(),
				.pld_8g_full_rx_fifo(),
				.pld_8g_full_rx_reg(),
				.pld_8g_full_rx_txclk_reg(),
				.pld_8g_g3_rx_pld_rst_n_reg(),
				.pld_8g_g3_rx_pld_rst_n_txclk_reg(),
				.pld_8g_rxelecidle_txclk_reg(),
				.pld_8g_rxpolarity_reg(),
				.pld_8g_rxpolarity_txclk_reg(),
				.pld_8g_wa_boundary_reg(),
				.pld_8g_wrdisable_rx_reg(),
				.pld_8g_wrdisable_rx_txclk_reg(),
				.pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_rx_clk_out_8g_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_wire(),
				.pld_rx_control_8g_reg(),
				.pld_rx_control_8g_txclk_reg(),
				.pld_rx_data_8g_reg(),
				.pld_rx_data_8g_txclk_reg(),
				.pld_syncsm_en_reg(),
				.pld_syncsm_en_txclk_reg(),
				.rm_fifo_partial_empty(),
				.rm_fifo_partial_full(),
				.sta_rx_clk2_by2_1(),
				.sta_rx_clk2_by2_1_out(),
				.sta_rx_clk2_by2_2(),
				.sta_rx_clk2_by2_2_out(),
				.sta_rx_clk2_by4_1(),
				.sta_rx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_rx_pcs_a1a2k1k2flag[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_rx_pcs_chnl_test_bus_out[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_clock_to_pld = 1'b0;
				assign w_hssi_8g_rx_pcs_dataout[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_dis_pc_byte = 1'b0;
				assign w_hssi_8g_rx_pcs_eidle_detected = 1'b0;
				assign w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_pma_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_gen2ngen1 = 1'b0;
				assign w_hssi_8g_rx_pcs_parallel_rev_loopback[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_pc_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_pcfifofull = 1'b0;
				assign w_hssi_8g_rx_pcs_phystatus = 1'b0;
				assign w_hssi_8g_rx_pcs_pipe_data[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_full = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clkslip = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_data_valid[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pma_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rxstatus[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_rxvalid = 1'b0;
				assign w_hssi_8g_rx_pcs_signal_detect_out = 1'b0;
				assign w_hssi_8g_rx_pcs_word_align_boundary[4:0] = 5'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79:0] = 80'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31:0] = 32'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_rmfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_tx_pcs
			twentynm_hssi_8g_tx_pcs #(
				.auto_speed_nego_gen2(hssi_8g_tx_pcs_auto_speed_nego_gen2),
				.bit_reversal(hssi_8g_tx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_tx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_tx_pcs_bypass_pipeline_reg),
				.byte_serializer(hssi_8g_tx_pcs_byte_serializer),
				.clock_gate_bs_enc(hssi_8g_tx_pcs_clock_gate_bs_enc),
				.clock_gate_dw_fifowr(hssi_8g_tx_pcs_clock_gate_dw_fifowr),
				.clock_gate_fiford(hssi_8g_tx_pcs_clock_gate_fiford),
				.clock_gate_sw_fifowr(hssi_8g_tx_pcs_clock_gate_sw_fifowr),
				.clock_observation_in_pld_core(hssi_8g_tx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_tx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_tx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_tx_pcs_ctrl_plane_bonding_distribution),
				.data_selection_8b10b_encoder_input(hssi_8g_tx_pcs_data_selection_8b10b_encoder_input),
				.dynamic_clk_switch(hssi_8g_tx_pcs_dynamic_clk_switch),
				.eightb_tenb_disp_ctrl(hssi_8g_tx_pcs_eightb_tenb_disp_ctrl),
				.eightb_tenb_encoder(hssi_8g_tx_pcs_eightb_tenb_encoder),
				.force_echar(hssi_8g_tx_pcs_force_echar),
				.force_kchar(hssi_8g_tx_pcs_force_kchar),
				.gen3_tx_clk_sel(hssi_8g_tx_pcs_gen3_tx_clk_sel),
				.gen3_tx_pipe_clk_sel(hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel),
				.hip_mode(hssi_8g_tx_pcs_hip_mode),
				.pcs_bypass(hssi_8g_tx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_tx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_tx_pcs_phase_compensation_fifo),
				.phfifo_write_clk_sel(hssi_8g_tx_pcs_phfifo_write_clk_sel),
				.pma_dw(hssi_8g_tx_pcs_pma_dw),
				.prot_mode(hssi_8g_tx_pcs_prot_mode),
				.reconfig_settings(hssi_8g_tx_pcs_reconfig_settings),
				.refclk_b_clk_sel(hssi_8g_tx_pcs_refclk_b_clk_sel),
				.revloop_back_rm(hssi_8g_tx_pcs_revloop_back_rm),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_tx_pcs_sup_mode),
				.symbol_swap(hssi_8g_tx_pcs_symbol_swap),
				.tx_bitslip(hssi_8g_tx_pcs_tx_bitslip),
				.tx_compliance_controlled_disparity(hssi_8g_tx_pcs_tx_compliance_controlled_disparity),
				.tx_fast_pld_reg(hssi_8g_tx_pcs_tx_fast_pld_reg),
				.txclk_freerun(hssi_8g_tx_pcs_txclk_freerun),
				.txpcs_urst(hssi_8g_tx_pcs_txpcs_urst)
			) inst_twentynm_hssi_8g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_8g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_tx_pcs_blockselect),
				.clk_out(w_hssi_8g_tx_pcs_clk_out),
				.clk_out_gen3(w_hssi_8g_tx_pcs_clk_out_gen3),
				.dataout(w_hssi_8g_tx_pcs_dataout),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.fifo_select_out_chnl_down(w_hssi_8g_tx_pcs_fifo_select_out_chnl_down),
				.fifo_select_out_chnl_up(w_hssi_8g_tx_pcs_fifo_select_out_chnl_up),
				.g3_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.g3_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
				.non_gray_eidleinfersel(w_hssi_8g_tx_pcs_non_gray_eidleinfersel),
				.ph_fifo_overflow(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.ph_fifo_underflow(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.phfifo_txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.phfifo_txmargin(w_hssi_8g_tx_pcs_phfifo_txmargin),
				.phfifo_txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				.pipe_en_rev_parallel_lpbk_out(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.pipe_power_down_out(w_hssi_8g_tx_pcs_pipe_power_down_out),
				.pipe_tx_clk_out_gen3(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pmaif_asn_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.rd_enable_out_chnl_down(w_hssi_8g_tx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_tx_pcs_rd_enable_out_chnl_up),
				.rd_ptr_tx_phfifo(w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rxpolarity_int(w_hssi_8g_tx_pcs_rxpolarity_int),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.tx_blk_start_out(w_hssi_8g_tx_pcs_tx_blk_start_out),
				.tx_clk_out_8g_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.tx_ctrlplane_testbus(w_hssi_8g_tx_pcs_tx_ctrlplane_testbus),
				.tx_data_out(w_hssi_8g_tx_pcs_tx_data_out),
				.tx_data_valid_out(w_hssi_8g_tx_pcs_tx_data_valid_out),
				.tx_datak_out(w_hssi_8g_tx_pcs_tx_datak_out),
				.tx_detect_rxloopback_int(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.tx_div_sync(w_hssi_8g_tx_pcs_tx_div_sync),
				.tx_div_sync_out_chnl_down(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down),
				.tx_div_sync_out_chnl_up(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up),
				.tx_pipe_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.tx_pipe_electidle(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_soft_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.tx_sync_hdr_out(w_hssi_8g_tx_pcs_tx_sync_hdr_out),
				.tx_testbus(w_hssi_8g_tx_pcs_tx_testbus),
				.txcompliance_out(w_hssi_8g_tx_pcs_txcompliance_out),
				.txelecidle_out(w_hssi_8g_tx_pcs_txelecidle_out),
				.wr_clk_tx_phfifo_dw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_tx_phfifo_sw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_data_tx_phfifo(w_hssi_8g_tx_pcs_wr_data_tx_phfifo),
				.wr_en_tx_phfifo(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_tx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_tx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_tx_phfifo(w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo),
				.wr_rst_n_tx_phfifo(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bitslip_boundary_select({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0]}),
				.clk_sel_gen3(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.coreclk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.datain({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.detectrxloopin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidleinfersel({w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0]}),
				.en_rev_parallel_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.fifo_select_in_chnl_down({in_bond_pcs8g_in_bot[11], in_bond_pcs8g_in_bot[10]}),
				.fifo_select_in_chnl_up({in_bond_pcs8g_in_top[11], in_bond_pcs8g_in_top[10]}),
				.hrdrst(1'b0),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.ph_fifo_rd_disable(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.pipe_en_rev_parallel_lpbk_in(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.pipe_tx_deemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.pipe_tx_margin({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0]}),
				.powerdn({w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0]}),
				.rate_switch(w_hssi_8g_rx_pcs_gen2ngen1),
				.rd_data_tx_phfifo({w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[9]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[9]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.rev_parallel_lpbk_data({w_hssi_8g_rx_pcs_parallel_rev_loopback[19], w_hssi_8g_rx_pcs_parallel_rev_loopback[18], w_hssi_8g_rx_pcs_parallel_rev_loopback[17], w_hssi_8g_rx_pcs_parallel_rev_loopback[16], w_hssi_8g_rx_pcs_parallel_rev_loopback[15], w_hssi_8g_rx_pcs_parallel_rev_loopback[14], w_hssi_8g_rx_pcs_parallel_rev_loopback[13], w_hssi_8g_rx_pcs_parallel_rev_loopback[12], w_hssi_8g_rx_pcs_parallel_rev_loopback[11], w_hssi_8g_rx_pcs_parallel_rev_loopback[10], w_hssi_8g_rx_pcs_parallel_rev_loopback[9], w_hssi_8g_rx_pcs_parallel_rev_loopback[8], w_hssi_8g_rx_pcs_parallel_rev_loopback[7], w_hssi_8g_rx_pcs_parallel_rev_loopback[6], w_hssi_8g_rx_pcs_parallel_rev_loopback[5], w_hssi_8g_rx_pcs_parallel_rev_loopback[4], w_hssi_8g_rx_pcs_parallel_rev_loopback[3], w_hssi_8g_rx_pcs_parallel_rev_loopback[2], w_hssi_8g_rx_pcs_parallel_rev_loopback[1], w_hssi_8g_rx_pcs_parallel_rev_loopback[0]}),
				.rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.tx_blk_start({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0]}),
				.tx_data_valid({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0]}),
				.tx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[7], in_bond_pcs8g_in_bot[6]}),
				.tx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[7], in_bond_pcs8g_in_top[6]}),
				.tx_pcs_reset(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.tx_sync_hdr({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0]}),
				.txd_fast_reg({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0]}),
				.txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[8]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[8]),
				.wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				
				// UNUSED
				.byte_serializer_pcs_clk_div_by_2_reg(),
				.byte_serializer_pcs_clk_div_by_2_wire(),
				.byte_serializer_pcs_clk_div_by_4_reg(),
				.byte_serializer_pld_clk_div_by_2_reg(),
				.byte_serializer_pld_clk_div_by_4_reg(),
				.pld_8g_empty_tx_fifo(),
				.pld_8g_empty_tx_reg(),
				.pld_8g_full_tx_fifo(),
				.pld_8g_full_tx_reg(),
				.pld_8g_g3_tx_pld_rst_n_reg(),
				.pld_8g_rddisable_tx_reg(),
				.pld_8g_tx_boundary_sel_reg(),
				.pld_pcs_tx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_tx_clk_out_8g_wire(),
				.pld_tx_data_8g_fifo(),
				.pld_tx_data_lo_8g_reg(),
				.sta_tx_clk2_by2_1(),
				.sta_tx_clk2_by2_1_out(),
				.sta_tx_clk2_by4_1(),
				.sta_tx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_dataout[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_dyn_clk_switch_n = 1'b1;		// Override default tieoff
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_g3_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_overflow = 1'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_underflow = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txdeemph = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txmargin[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txswing = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_power_down_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_pmaif_asn_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_refclk_b = 1'b0;
				assign w_hssi_8g_tx_pcs_refclk_b_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_rxpolarity_int = 1'b0;
				assign w_hssi_8g_tx_pcs_soft_reset_wclk1_n = 1'b0;
				assign w_hssi_8g_tx_pcs_sw_fifo_wr_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_blk_start_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_tx_data_out[31:0] = 32'b0;
				assign w_hssi_8g_tx_pcs_tx_data_valid_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_datak_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_detect_rxloopback_int = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_electidle = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_sync_hdr_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_txcompliance_out = 1'b0;
				assign w_hssi_8g_tx_pcs_txelecidle_out = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63:0] = 64'b0;
				assign w_hssi_8g_tx_pcs_wr_en_tx_phfifo = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pcs_pma_interface
			twentynm_hssi_common_pcs_pma_interface #(
				.asn_clk_enable(hssi_common_pcs_pma_interface_asn_clk_enable),
				.asn_enable(hssi_common_pcs_pma_interface_asn_enable),
				.block_sel(hssi_common_pcs_pma_interface_block_sel),
				.bypass_early_eios(hssi_common_pcs_pma_interface_bypass_early_eios),
				.bypass_pcie_switch(hssi_common_pcs_pma_interface_bypass_pcie_switch),
				.bypass_pma_ltr(hssi_common_pcs_pma_interface_bypass_pma_ltr),
				.bypass_pma_sw_done(hssi_common_pcs_pma_interface_bypass_pma_sw_done),
				.bypass_ppm_lock(hssi_common_pcs_pma_interface_bypass_ppm_lock),
				.bypass_send_syncp_fbkp(hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp),
				.bypass_txdetectrx(hssi_common_pcs_pma_interface_bypass_txdetectrx),
				.cdr_control(hssi_common_pcs_pma_interface_cdr_control),
				.cid_enable(hssi_common_pcs_pma_interface_cid_enable),
				.cp_cons_sel(hssi_common_pcs_pma_interface_cp_cons_sel),
				.cp_dwn_mstr(hssi_common_pcs_pma_interface_cp_dwn_mstr),
				.cp_up_mstr(hssi_common_pcs_pma_interface_cp_up_mstr),
				.ctrl_plane_bonding(hssi_common_pcs_pma_interface_ctrl_plane_bonding),
				.data_mask_count(hssi_common_pcs_pma_interface_data_mask_count),
				.data_mask_count_multi(hssi_common_pcs_pma_interface_data_mask_count_multi),
				.dft_observation_clock_selection(hssi_common_pcs_pma_interface_dft_observation_clock_selection),
				.early_eios_counter(hssi_common_pcs_pma_interface_early_eios_counter),
				.force_freqdet(hssi_common_pcs_pma_interface_force_freqdet),
				.free_run_clk_enable(hssi_common_pcs_pma_interface_free_run_clk_enable),
				.ignore_sigdet_g23(hssi_common_pcs_pma_interface_ignore_sigdet_g23),
				.pc_en_counter(hssi_common_pcs_pma_interface_pc_en_counter),
				.pc_rst_counter(hssi_common_pcs_pma_interface_pc_rst_counter),
				.pcie_hip_mode(hssi_common_pcs_pma_interface_pcie_hip_mode),
				.ph_fifo_reg_mode(hssi_common_pcs_pma_interface_ph_fifo_reg_mode),
				.phfifo_flush_wait(hssi_common_pcs_pma_interface_phfifo_flush_wait),
				.pipe_if_g3pcs(hssi_common_pcs_pma_interface_pipe_if_g3pcs),
				.pma_done_counter(hssi_common_pcs_pma_interface_pma_done_counter),
				.pma_if_dft_en(hssi_common_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_common_pcs_pma_interface_pma_if_dft_val),
				.ppm_cnt_rst(hssi_common_pcs_pma_interface_ppm_cnt_rst),
				.ppm_deassert_early(hssi_common_pcs_pma_interface_ppm_deassert_early),
				.ppm_det_buckets(hssi_common_pcs_pma_interface_ppm_det_buckets),
				.ppm_gen1_2_cnt(hssi_common_pcs_pma_interface_ppm_gen1_2_cnt),
				.ppm_post_eidle_delay(hssi_common_pcs_pma_interface_ppm_post_eidle_delay),
				.ppmsel(hssi_common_pcs_pma_interface_ppmsel),
				.prot_mode(hssi_common_pcs_pma_interface_prot_mode),
				.reconfig_settings(hssi_common_pcs_pma_interface_reconfig_settings),
				.rxvalid_mask(hssi_common_pcs_pma_interface_rxvalid_mask),
				.sigdet_wait_counter(hssi_common_pcs_pma_interface_sigdet_wait_counter),
				.sigdet_wait_counter_multi(hssi_common_pcs_pma_interface_sigdet_wait_counter_multi),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sim_mode(hssi_common_pcs_pma_interface_sim_mode),
				.spd_chg_rst_wait_cnt_en(hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en),
				.sup_mode(hssi_common_pcs_pma_interface_sup_mode),
				.testout_sel(hssi_common_pcs_pma_interface_testout_sel),
				.wait_clk_on_off_timer(hssi_common_pcs_pma_interface_wait_clk_on_off_timer),
				.wait_pipe_synchronizing(hssi_common_pcs_pma_interface_wait_pipe_synchronizing),
				.wait_send_syncp_fbkp(hssi_common_pcs_pma_interface_wait_send_syncp_fbkp)
			) inst_twentynm_hssi_common_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_common_pcs_pma_interface_blockselect),
				.int_pmaif_8g_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in),
				.int_pmaif_8g_eios_detected(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.int_pmaif_8g_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.int_pmaif_8g_power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.int_pmaif_g3_pcs_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in),
				.int_pmaif_pldif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pmaif_pldif_pcie_sw_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done),
				.int_pmaif_pldif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pmaif_pldif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pmaif_pldif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pmaif_pldif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pmaif_pldif_pma_reserved_in(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in),
				.int_pmaif_pldif_test_out(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out),
				.int_pmaif_pldif_testbus(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus),
				.pma_adapt_start(w_hssi_common_pcs_pma_interface_pma_adapt_start),
				.pma_atpg_los_en_n(w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n),
				.pma_csr_test_dis(w_hssi_common_pcs_pma_interface_pma_csr_test_dis),
				.pma_current_coeff(w_hssi_common_pcs_pma_interface_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_common_pcs_pma_interface_pma_current_rxpreset),
				.pma_early_eios(w_hssi_common_pcs_pma_interface_pma_early_eios),
				.pma_interface_select(w_hssi_common_pcs_pma_interface_pma_interface_select),
				.pma_ltd_b(w_hssi_common_pcs_pma_interface_pma_ltd_b),
				.pma_ltr(w_hssi_common_pcs_pma_interface_pma_ltr),
				.pma_nfrzdrv(w_hssi_common_pcs_pma_interface_pma_nfrzdrv),
				.pma_nrpi_freeze(w_hssi_common_pcs_pma_interface_pma_nrpi_freeze),
				.pma_pcie_switch(w_hssi_common_pcs_pma_interface_pma_pcie_switch),
				.pma_ppm_lock(w_hssi_common_pcs_pma_interface_pma_ppm_lock),
				.pma_reserved_out(w_hssi_common_pcs_pma_interface_pma_reserved_out),
				.pma_rs_lpbk_b(w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b),
				.pma_rx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup),
				.pma_scan_mode_n(w_hssi_common_pcs_pma_interface_pma_scan_mode_n),
				.pma_scan_shift_n(w_hssi_common_pcs_pma_interface_pma_scan_shift_n),
				.pma_tx_bitslip(w_hssi_common_pcs_pma_interface_pma_tx_bitslip),
				.pma_tx_bonding_rstb(w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb),
				.pma_tx_qpi_pulldn(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn),
				.pma_tx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup),
				.pma_tx_txdetectrx(w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx),
				.pmaif_bundling_out_down(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down),
				.pmaif_bundling_out_up(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_8g_current_coeff({w_hssi_pipe_gen1_2_current_coeff[17], w_hssi_pipe_gen1_2_current_coeff[16], w_hssi_pipe_gen1_2_current_coeff[15], w_hssi_pipe_gen1_2_current_coeff[14], w_hssi_pipe_gen1_2_current_coeff[13], w_hssi_pipe_gen1_2_current_coeff[12], w_hssi_pipe_gen1_2_current_coeff[11], w_hssi_pipe_gen1_2_current_coeff[10], w_hssi_pipe_gen1_2_current_coeff[9], w_hssi_pipe_gen1_2_current_coeff[8], w_hssi_pipe_gen1_2_current_coeff[7], w_hssi_pipe_gen1_2_current_coeff[6], w_hssi_pipe_gen1_2_current_coeff[5], w_hssi_pipe_gen1_2_current_coeff[4], w_hssi_pipe_gen1_2_current_coeff[3], w_hssi_pipe_gen1_2_current_coeff[2], w_hssi_pipe_gen1_2_current_coeff[1], w_hssi_pipe_gen1_2_current_coeff[0]}),
				.int_pmaif_8g_eios_det({w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0]}),
				.int_pmaif_8g_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.int_pmaif_8g_rev_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.int_pmaif_8g_tx_clk_out_gen3(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.int_pmaif_8g_txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				.int_pmaif_g3_eios_det({w_hssi_gen3_rx_pcs_ei_det_int, w_hssi_gen3_rx_pcs_ei_partial_det_int, w_hssi_gen3_rx_pcs_i_det_int}),
				.int_pmaif_g3_pma_current_coeff({w_hssi_pipe_gen3_pma_current_coeff[17], w_hssi_pipe_gen3_pma_current_coeff[16], w_hssi_pipe_gen3_pma_current_coeff[15], w_hssi_pipe_gen3_pma_current_coeff[14], w_hssi_pipe_gen3_pma_current_coeff[13], w_hssi_pipe_gen3_pma_current_coeff[12], w_hssi_pipe_gen3_pma_current_coeff[11], w_hssi_pipe_gen3_pma_current_coeff[10], w_hssi_pipe_gen3_pma_current_coeff[9], w_hssi_pipe_gen3_pma_current_coeff[8], w_hssi_pipe_gen3_pma_current_coeff[7], w_hssi_pipe_gen3_pma_current_coeff[6], w_hssi_pipe_gen3_pma_current_coeff[5], w_hssi_pipe_gen3_pma_current_coeff[4], w_hssi_pipe_gen3_pma_current_coeff[3], w_hssi_pipe_gen3_pma_current_coeff[2], w_hssi_pipe_gen3_pma_current_coeff[1], w_hssi_pipe_gen3_pma_current_coeff[0]}),
				.int_pmaif_g3_pma_current_rxpreset({w_hssi_pipe_gen3_pma_current_rxpreset[2], w_hssi_pipe_gen3_pma_current_rxpreset[1], w_hssi_pipe_gen3_pma_current_rxpreset[0]}),
				.int_pmaif_g3_pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.int_pmaif_g3_rev_lpbk(w_hssi_pipe_gen3_rev_lpbk_int),
				.int_pmaif_pldif_8g_tx_pld_rstn(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pmaif_pldif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pmaif_pldif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pmaif_pldif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pmaif_pldif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pmaif_pldif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pmaif_pldif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pmaif_pldif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pmaif_pldif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pmaif_pldif_pcie_switch({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0]}),
				.int_pmaif_pldif_pma_reserved_out({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0]}),
				.int_pmaif_pldif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pmaif_pldif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pmaif_pldif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pmaif_pldif_rate({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0]}),
				.int_pmaif_pldif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pmaif_pldif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pmaif_pldif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.int_pmaif_pldif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pmaif_pldif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pmaif_pldif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pmaif_pldif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pmaif_pldif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pmaif_pldif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.int_tx_dft_obsrv_clk({w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0]}),
				.iocsr_clk(in_iocsr_clk),
				.iocsr_config({in_iocsr_config[5], in_iocsr_config[4], in_iocsr_config[3], in_iocsr_config[2], in_iocsr_config[1], in_iocsr_config[0]}),
				.iocsr_rdy(in_iocsr_rdy),
				.iocsr_rdy_dly(in_iocsr_rdy_dly),
				.pma_adapt_done(in_pma_adapt_done),
				.pma_clklow(in_pma_clklow),
				.pma_fref(in_pma_fref),
				.pma_hclk(in_pma_hclk),
				.pma_pcie_sw_done({in_pma_pcie_sw_done[1], in_pma_pcie_sw_done[0]}),
				.pma_pfdmode_lock(in_pma_pfdmode_lock),
				.pma_reserved_in({in_pma_reserved_in[4], in_pma_reserved_in[3], in_pma_reserved_in[2], in_pma_reserved_in[1], in_pma_reserved_in[0]}),
				.pma_signal_det(in_pma_signal_det),
				.pma_testbus({in_pma_testbus[7], in_pma_testbus[6], in_pma_testbus[5], in_pma_testbus[4], in_pma_testbus[3], in_pma_testbus[2], in_pma_testbus[1], in_pma_testbus[0]}),
				.pmaif_bundling_in_down({in_bond_pmaif_in_bot[11], in_bond_pmaif_in_bot[10], in_bond_pmaif_in_bot[9], in_bond_pmaif_in_bot[8], in_bond_pmaif_in_bot[7], in_bond_pmaif_in_bot[6], in_bond_pmaif_in_bot[5], in_bond_pmaif_in_bot[4], in_bond_pmaif_in_bot[3], in_bond_pmaif_in_bot[2], in_bond_pmaif_in_bot[1], in_bond_pmaif_in_bot[0]}),
				.pmaif_bundling_in_up({in_bond_pmaif_in_top[11], in_bond_pmaif_in_top[10], in_bond_pmaif_in_top[9], in_bond_pmaif_in_top[8], in_bond_pmaif_in_top[7], in_bond_pmaif_in_top[6], in_bond_pmaif_in_top[5], in_bond_pmaif_in_top[4], in_bond_pmaif_in_top[3], in_bond_pmaif_in_top[2], in_bond_pmaif_in_top[1], in_bond_pmaif_in_top[0]}),
				.rx_pmaif_test_out({w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0]}),
				.rx_prbs_ver_test({w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0]}),
				.tx_prbs_gen_test({w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0]}),
				.uhsif_test_out_1({w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0]}),
				.uhsif_test_out_2({w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0]}),
				.uhsif_test_out_3({w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0]}),
				
				// UNUSED
				.int_pmaif_avmm_iocsr_clk(),
				.int_pmaif_avmm_iocsr_config(),
				.int_pmaif_avmm_iocsr_rdy(),
				.int_pmaif_avmm_iocsr_rdy_dly(),
				.int_pmaif_pldif_interface_select(),
				.pma_tx_pma_syncp(),
				.sta_pma_hclk_by2()
			);
		end // if generate
		else begin
				assign w_hssi_common_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19:0] = 20'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_pma_adapt_start = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_csr_test_dis = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pcs_pma_interface_pma_early_eios = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_interface_select[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltd_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltr = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nfrzdrv = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nrpi_freeze = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ppm_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_tx_bitslip = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx = in_pld_pma_txdetectrx;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11:0] = 12'b0;
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11:0] = 12'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pld_pcs_interface
			twentynm_hssi_common_pld_pcs_interface #(
				.dft_clk_out_en(hssi_common_pld_pcs_interface_dft_clk_out_en),
				.dft_clk_out_sel(hssi_common_pld_pcs_interface_dft_clk_out_sel),
				.hrdrstctrl_en(hssi_common_pld_pcs_interface_hrdrstctrl_en),
				.pcs_testbus_block_sel(hssi_common_pld_pcs_interface_pcs_testbus_block_sel),
				.reconfig_settings(hssi_common_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm3" )       //PARAM_HIDE
			) inst_twentynm_hssi_common_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_common_pld_pcs_interface_blockselect),
				.hip_cmn_clk(w_hssi_common_pld_pcs_interface_hip_cmn_clk),
				.hip_cmn_ctrl(w_hssi_common_pld_pcs_interface_hip_cmn_ctrl),
				.hip_iocsr_rdy(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy),
				.hip_iocsr_rdy_dly(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly),
				.hip_nfrzdrv(w_hssi_common_pld_pcs_interface_hip_nfrzdrv),
				.hip_npor(w_hssi_common_pld_pcs_interface_hip_npor),
				.hip_usermode(w_hssi_common_pld_pcs_interface_hip_usermode),
				.int_pldif_10g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.int_pldif_10g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.int_pldif_8g_eidleinfersel(w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel),
				.int_pldif_8g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.int_pldif_8g_refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.int_pldif_8g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.int_pldif_g3_current_coeff(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff),
				.int_pldif_g3_current_rxpreset(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset),
				.int_pldif_krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.int_pldif_krfec_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.int_pldif_krfec_scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				.int_pldif_mem_atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.int_pldif_mem_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.int_pldif_pmaif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pldif_pmaif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pldif_pmaif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pldif_pmaif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pldif_pmaif_eye_monitor(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor),
				.int_pldif_pmaif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pldif_pmaif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pldif_pmaif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pldif_pmaif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pldif_pmaif_pcie_switch(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch),
				.int_pldif_pmaif_pma_reserved_out(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out),
				.int_pldif_pmaif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pldif_pmaif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pldif_pmaif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pldif_pmaif_rate(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate),
				.int_pldif_pmaif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pldif_pmaif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pldif_pmaif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pldif_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_pldif_pmaif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pldif_pmaif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pldif_pmaif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pldif_pmaif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pldif_pmaif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pldif_pmaif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pldif_pmaif_uhsif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.pld_pma_adapt_done(w_hssi_common_pld_pcs_interface_pld_pma_adapt_done),
				.pld_pma_clklow(w_hssi_common_pld_pcs_interface_pld_pma_clklow),
				.pld_pma_fref(w_hssi_common_pld_pcs_interface_pld_pma_fref),
				.pld_pma_hclk(w_hssi_common_pld_pcs_interface_pld_pma_hclk),
				.pld_pma_pcie_sw_done(w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done),
				.pld_pma_pfdmode_lock(w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock),
				.pld_pma_reserved_in(w_hssi_common_pld_pcs_interface_pld_pma_reserved_in),
				.pld_pma_rx_detect_valid(w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid),
				.pld_pma_rx_found(w_hssi_common_pld_pcs_interface_pld_pma_rx_found),
				.pld_pma_rxpll_lock(w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock),
				.pld_pma_testbus(w_hssi_common_pld_pcs_interface_pld_pma_testbus),
				.pld_pmaif_mask_tx_pll(w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll),
				.pld_reserved_out(w_hssi_common_pld_pcs_interface_pld_reserved_out),
				.pld_test_data(w_hssi_common_pld_pcs_interface_pld_test_data),
				.pld_uhsif_lock(w_hssi_common_pld_pcs_interface_pld_uhsif_lock),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.int_pldif_10g_test_data({w_hssi_10g_tx_pcs_tx_test_data[19], w_hssi_10g_tx_pcs_tx_test_data[18], w_hssi_10g_tx_pcs_tx_test_data[17], w_hssi_10g_tx_pcs_tx_test_data[16], w_hssi_10g_tx_pcs_tx_test_data[15], w_hssi_10g_tx_pcs_tx_test_data[14], w_hssi_10g_tx_pcs_tx_test_data[13], w_hssi_10g_tx_pcs_tx_test_data[12], w_hssi_10g_tx_pcs_tx_test_data[11], w_hssi_10g_tx_pcs_tx_test_data[10], w_hssi_10g_tx_pcs_tx_test_data[9], w_hssi_10g_tx_pcs_tx_test_data[8], w_hssi_10g_tx_pcs_tx_test_data[7], w_hssi_10g_tx_pcs_tx_test_data[6], w_hssi_10g_tx_pcs_tx_test_data[5], w_hssi_10g_tx_pcs_tx_test_data[4], w_hssi_10g_tx_pcs_tx_test_data[3], w_hssi_10g_tx_pcs_tx_test_data[2], w_hssi_10g_tx_pcs_tx_test_data[1], w_hssi_10g_tx_pcs_tx_test_data[0]}),
				.int_pldif_10g_tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.int_pldif_8g_chnl_test_bus_out({w_hssi_8g_rx_pcs_chnl_test_bus_out[19], w_hssi_8g_rx_pcs_chnl_test_bus_out[18], w_hssi_8g_rx_pcs_chnl_test_bus_out[17], w_hssi_8g_rx_pcs_chnl_test_bus_out[16], w_hssi_8g_rx_pcs_chnl_test_bus_out[15], w_hssi_8g_rx_pcs_chnl_test_bus_out[14], w_hssi_8g_rx_pcs_chnl_test_bus_out[13], w_hssi_8g_rx_pcs_chnl_test_bus_out[12], w_hssi_8g_rx_pcs_chnl_test_bus_out[11], w_hssi_8g_rx_pcs_chnl_test_bus_out[10], w_hssi_8g_rx_pcs_chnl_test_bus_out[9], w_hssi_8g_rx_pcs_chnl_test_bus_out[8], w_hssi_8g_rx_pcs_chnl_test_bus_out[7], w_hssi_8g_rx_pcs_chnl_test_bus_out[6], w_hssi_8g_rx_pcs_chnl_test_bus_out[5], w_hssi_8g_rx_pcs_chnl_test_bus_out[4], w_hssi_8g_rx_pcs_chnl_test_bus_out[3], w_hssi_8g_rx_pcs_chnl_test_bus_out[2], w_hssi_8g_rx_pcs_chnl_test_bus_out[1], w_hssi_8g_rx_pcs_chnl_test_bus_out[0]}),
				.int_pldif_8g_rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.int_pldif_8g_tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.int_pldif_g3_test_out({w_hssi_pipe_gen3_test_out[19], w_hssi_pipe_gen3_test_out[18], w_hssi_pipe_gen3_test_out[17], w_hssi_pipe_gen3_test_out[16], w_hssi_pipe_gen3_test_out[15], w_hssi_pipe_gen3_test_out[14], w_hssi_pipe_gen3_test_out[13], w_hssi_pipe_gen3_test_out[12], w_hssi_pipe_gen3_test_out[11], w_hssi_pipe_gen3_test_out[10], w_hssi_pipe_gen3_test_out[9], w_hssi_pipe_gen3_test_out[8], w_hssi_pipe_gen3_test_out[7], w_hssi_pipe_gen3_test_out[6], w_hssi_pipe_gen3_test_out[5], w_hssi_pipe_gen3_test_out[4], w_hssi_pipe_gen3_test_out[3], w_hssi_pipe_gen3_test_out[2], w_hssi_pipe_gen3_test_out[1], w_hssi_pipe_gen3_test_out[0]}),
				.int_pldif_krfec_test_data({w_hssi_krfec_tx_pcs_tx_test_data[19], w_hssi_krfec_tx_pcs_tx_test_data[18], w_hssi_krfec_tx_pcs_tx_test_data[17], w_hssi_krfec_tx_pcs_tx_test_data[16], w_hssi_krfec_tx_pcs_tx_test_data[15], w_hssi_krfec_tx_pcs_tx_test_data[14], w_hssi_krfec_tx_pcs_tx_test_data[13], w_hssi_krfec_tx_pcs_tx_test_data[12], w_hssi_krfec_tx_pcs_tx_test_data[11], w_hssi_krfec_tx_pcs_tx_test_data[10], w_hssi_krfec_tx_pcs_tx_test_data[9], w_hssi_krfec_tx_pcs_tx_test_data[8], w_hssi_krfec_tx_pcs_tx_test_data[7], w_hssi_krfec_tx_pcs_tx_test_data[6], w_hssi_krfec_tx_pcs_tx_test_data[5], w_hssi_krfec_tx_pcs_tx_test_data[4], w_hssi_krfec_tx_pcs_tx_test_data[3], w_hssi_krfec_tx_pcs_tx_test_data[2], w_hssi_krfec_tx_pcs_tx_test_data[1], w_hssi_krfec_tx_pcs_tx_test_data[0]}),
				.int_pldif_pmaif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pldif_pmaif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pldif_pmaif_pcie_sw_done({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0]}),
				.int_pldif_pmaif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pldif_pmaif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pldif_pmaif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pldif_pmaif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pldif_pmaif_pma_reserved_in({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0]}),
				.int_pldif_pmaif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pldif_pmaif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_test_out({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0]}),
				.int_pldif_pmaif_testbus({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0]}),
				.int_pldif_pmaif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.pld_8g_eidleinfersel({in_pld_8g_eidleinfersel[2], in_pld_8g_eidleinfersel[1], in_pld_8g_eidleinfersel[0]}),
				.pld_8g_refclk_dig2(in_pld_8g_refclk_dig2),
				.pld_atpg_los_en_n(in_pld_atpg_los_en_n),
				.pld_g3_current_coeff({in_pld_g3_current_coeff[17], in_pld_g3_current_coeff[16], in_pld_g3_current_coeff[15], in_pld_g3_current_coeff[14], in_pld_g3_current_coeff[13], in_pld_g3_current_coeff[12], in_pld_g3_current_coeff[11], in_pld_g3_current_coeff[10], in_pld_g3_current_coeff[9], in_pld_g3_current_coeff[8], in_pld_g3_current_coeff[7], in_pld_g3_current_coeff[6], in_pld_g3_current_coeff[5], in_pld_g3_current_coeff[4], in_pld_g3_current_coeff[3], in_pld_g3_current_coeff[2], in_pld_g3_current_coeff[1], in_pld_g3_current_coeff[0]}),
				.pld_g3_current_rxpreset({in_pld_g3_current_rxpreset[2], in_pld_g3_current_rxpreset[1], in_pld_g3_current_rxpreset[0]}),
				.pld_ltr(in_pld_ltr),
				.pld_mem_krfec_atpg_rst_n(in_pld_mem_krfec_atpg_rst_n),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pcs_refclk_dig(in_pld_pcs_refclk_dig),
				.pld_pma_adapt_start(in_pld_pma_adapt_start),
				.pld_pma_csr_test_dis(in_pld_pma_csr_test_dis),
				.pld_pma_early_eios(in_pld_pma_early_eios),
				.pld_pma_eye_monitor({in_pld_pma_eye_monitor[5], in_pld_pma_eye_monitor[4], in_pld_pma_eye_monitor[3], in_pld_pma_eye_monitor[2], in_pld_pma_eye_monitor[1], in_pld_pma_eye_monitor[0]}),
				.pld_pma_ltd_b(in_pld_pma_ltd_b),
				.pld_pma_nrpi_freeze(in_pld_pma_nrpi_freeze),
				.pld_pma_pcie_switch({in_pld_pma_pcie_switch[1], in_pld_pma_pcie_switch[0]}),
				.pld_pma_ppm_lock(in_pld_pma_ppm_lock),
				.pld_pma_reserved_out({in_pld_pma_reserved_out[4], in_pld_pma_reserved_out[3], in_pld_pma_reserved_out[2], in_pld_pma_reserved_out[1], in_pld_pma_reserved_out[0]}),
				.pld_pma_rs_lpbk_b(in_pld_pma_rs_lpbk_b),
				.pld_pma_rx_qpi_pullup(in_pld_pma_rx_qpi_pullup),
				.pld_pma_tx_bitslip(in_pld_pma_tx_bitslip),
				.pld_pma_tx_bonding_rstb(in_pld_pma_tx_bonding_rstb),
				.pld_pma_tx_qpi_pulldn(in_pld_pma_tx_qpi_pulldn),
				.pld_pma_tx_qpi_pullup(in_pld_pma_tx_qpi_pullup),
				.pld_pma_txdetectrx(in_pld_pma_txdetectrx),
				.pld_rate({in_pld_rate[1], in_pld_rate[0]}),
				.pld_reserved_in({in_pld_reserved_in[9], in_pld_reserved_in[8], in_pld_reserved_in[7], in_pld_reserved_in[6], in_pld_reserved_in[5], in_pld_reserved_in[4], in_pld_reserved_in[3], in_pld_reserved_in[2], in_pld_reserved_in[1], in_pld_reserved_in[0]}),
				.pld_scan_mode_n(in_pld_scan_mode_n),
				.pld_scan_shift_n(in_pld_scan_shift_n),
				
				// UNUSED
				.int_pldif_8g_ltr(),
				.int_pldif_avmm_pld_avmm1_request(),
				.int_pldif_avmm_pld_avmm2_request(),
				.int_pldif_avmm_refclk_dig_en(),
				.int_pldif_g3_scan_mode_n(),
				.pld_8g_eidleinfersel_fifo(),
				.pld_8g_eidleinfersel_reg(),
				.pld_partial_reconfig_fifo(),
				.pld_partial_reconfig_rx_div_by_2_rxclk_wire(),
				.pld_partial_reconfig_rx_div_by_2_txclk_wire(),
				.pld_partial_reconfig_rxclk_reg(),
				.pld_partial_reconfig_tx_div_by_2_wire(),
				.pld_partial_reconfig_txclk_reg(),
				.pld_rate_reg(),
				.pld_test_data_reg()
			);
		end // if generate
		else begin
				assign w_hssi_common_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_clk[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_npor = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_usermode = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2 = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_adapt_done = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_clklow = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_fref = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_hclk = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_found = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_testbus[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_reserved_out[9:0] = 10'b0;
				assign w_hssi_common_pld_pcs_interface_pld_test_data[19:0] = 20'b0;
				assign w_hssi_common_pld_pcs_interface_pld_uhsif_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_scan_mode_n = 1'b1;		// Override default tieoff
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_rx_pcs
			twentynm_hssi_fifo_rx_pcs #(
				.double_read_mode(hssi_fifo_rx_pcs_double_read_mode),
				.prot_mode(hssi_fifo_rx_pcs_prot_mode),
				.silicon_rev( "20nm3" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_rx_pcs_blockselect),
				.data_out2_10g(w_hssi_fifo_rx_pcs_data_out2_10g),
				.data_out2_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp),
				.data_out_10g(w_hssi_fifo_rx_pcs_data_out_10g),
				.data_out_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out_8g_clock_comp),
				.data_out_8g_phase_comp(w_hssi_fifo_rx_pcs_data_out_8g_phase_comp),
				.data_out_gen3(w_hssi_fifo_rx_pcs_data_out_gen3),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_data[73], w_hssi_10g_rx_pcs_rx_fifo_wr_data[72], w_hssi_10g_rx_pcs_rx_fifo_wr_data[71], w_hssi_10g_rx_pcs_rx_fifo_wr_data[70], w_hssi_10g_rx_pcs_rx_fifo_wr_data[69], w_hssi_10g_rx_pcs_rx_fifo_wr_data[68], w_hssi_10g_rx_pcs_rx_fifo_wr_data[67], w_hssi_10g_rx_pcs_rx_fifo_wr_data[66], w_hssi_10g_rx_pcs_rx_fifo_wr_data[65], w_hssi_10g_rx_pcs_rx_fifo_wr_data[64], w_hssi_10g_rx_pcs_rx_fifo_wr_data[63], w_hssi_10g_rx_pcs_rx_fifo_wr_data[62], w_hssi_10g_rx_pcs_rx_fifo_wr_data[61], w_hssi_10g_rx_pcs_rx_fifo_wr_data[60], w_hssi_10g_rx_pcs_rx_fifo_wr_data[59], w_hssi_10g_rx_pcs_rx_fifo_wr_data[58], w_hssi_10g_rx_pcs_rx_fifo_wr_data[57], w_hssi_10g_rx_pcs_rx_fifo_wr_data[56], w_hssi_10g_rx_pcs_rx_fifo_wr_data[55], w_hssi_10g_rx_pcs_rx_fifo_wr_data[54], w_hssi_10g_rx_pcs_rx_fifo_wr_data[53], w_hssi_10g_rx_pcs_rx_fifo_wr_data[52], w_hssi_10g_rx_pcs_rx_fifo_wr_data[51], w_hssi_10g_rx_pcs_rx_fifo_wr_data[50], w_hssi_10g_rx_pcs_rx_fifo_wr_data[49], w_hssi_10g_rx_pcs_rx_fifo_wr_data[48], w_hssi_10g_rx_pcs_rx_fifo_wr_data[47], w_hssi_10g_rx_pcs_rx_fifo_wr_data[46], w_hssi_10g_rx_pcs_rx_fifo_wr_data[45], w_hssi_10g_rx_pcs_rx_fifo_wr_data[44], w_hssi_10g_rx_pcs_rx_fifo_wr_data[43], w_hssi_10g_rx_pcs_rx_fifo_wr_data[42], w_hssi_10g_rx_pcs_rx_fifo_wr_data[41], w_hssi_10g_rx_pcs_rx_fifo_wr_data[40], w_hssi_10g_rx_pcs_rx_fifo_wr_data[39], w_hssi_10g_rx_pcs_rx_fifo_wr_data[38], w_hssi_10g_rx_pcs_rx_fifo_wr_data[37], w_hssi_10g_rx_pcs_rx_fifo_wr_data[36], w_hssi_10g_rx_pcs_rx_fifo_wr_data[35], w_hssi_10g_rx_pcs_rx_fifo_wr_data[34], w_hssi_10g_rx_pcs_rx_fifo_wr_data[33], w_hssi_10g_rx_pcs_rx_fifo_wr_data[32], w_hssi_10g_rx_pcs_rx_fifo_wr_data[31], w_hssi_10g_rx_pcs_rx_fifo_wr_data[30], w_hssi_10g_rx_pcs_rx_fifo_wr_data[29], w_hssi_10g_rx_pcs_rx_fifo_wr_data[28], w_hssi_10g_rx_pcs_rx_fifo_wr_data[27], w_hssi_10g_rx_pcs_rx_fifo_wr_data[26], w_hssi_10g_rx_pcs_rx_fifo_wr_data[25], w_hssi_10g_rx_pcs_rx_fifo_wr_data[24], w_hssi_10g_rx_pcs_rx_fifo_wr_data[23], w_hssi_10g_rx_pcs_rx_fifo_wr_data[22], w_hssi_10g_rx_pcs_rx_fifo_wr_data[21], w_hssi_10g_rx_pcs_rx_fifo_wr_data[20], w_hssi_10g_rx_pcs_rx_fifo_wr_data[19], w_hssi_10g_rx_pcs_rx_fifo_wr_data[18], w_hssi_10g_rx_pcs_rx_fifo_wr_data[17], w_hssi_10g_rx_pcs_rx_fifo_wr_data[16], w_hssi_10g_rx_pcs_rx_fifo_wr_data[15], w_hssi_10g_rx_pcs_rx_fifo_wr_data[14], w_hssi_10g_rx_pcs_rx_fifo_wr_data[13], w_hssi_10g_rx_pcs_rx_fifo_wr_data[12], w_hssi_10g_rx_pcs_rx_fifo_wr_data[11], w_hssi_10g_rx_pcs_rx_fifo_wr_data[10], w_hssi_10g_rx_pcs_rx_fifo_wr_data[9], w_hssi_10g_rx_pcs_rx_fifo_wr_data[8], w_hssi_10g_rx_pcs_rx_fifo_wr_data[7], w_hssi_10g_rx_pcs_rx_fifo_wr_data[6], w_hssi_10g_rx_pcs_rx_fifo_wr_data[5], w_hssi_10g_rx_pcs_rx_fifo_wr_data[4], w_hssi_10g_rx_pcs_rx_fifo_wr_data[3], w_hssi_10g_rx_pcs_rx_fifo_wr_data[2], w_hssi_10g_rx_pcs_rx_fifo_wr_data[1], w_hssi_10g_rx_pcs_rx_fifo_wr_data[0]}),
				.data_in_8g_clock_comp({w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0]}),
				.data_in_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr2_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0]}),
				.rd_ptr2_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0]}),
				.rd_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0]}),
				.rd_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.wr_clk_8g_clock_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_8g_clock_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.wr_en_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.wr_en_8g_clock_comp(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_en_8g_phase_comp(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.wr_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0]}),
				.wr_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0]}),
				.wr_rst_n_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.wr_rst_n_8g_clock_comp(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_n_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_rx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79:0] = 80'b0;
				assign w_hssi_fifo_rx_pcs_data_out_gen3[39:0] = 40'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_tx_pcs
			twentynm_hssi_fifo_tx_pcs #(
				.double_write_mode(hssi_fifo_tx_pcs_double_write_mode),
				.prot_mode(hssi_fifo_tx_pcs_prot_mode),
				.silicon_rev( "20nm3" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_tx_pcs_blockselect),
				.data_out_10g(w_hssi_fifo_tx_pcs_data_out_10g),
				.data_out_8g_phase_comp(w_hssi_fifo_tx_pcs_data_out_8g_phase_comp),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in2_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0]}),
				.data_in_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_en_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.wr_en_8g_phase_comp(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0]}),
				.wr_rst_n_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_tx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_tx_pcs_data_out_10g[72:0] = 73'b0;
				assign w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63:0] = 64'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_rx_pcs
			twentynm_hssi_gen3_rx_pcs #(
				.block_sync(hssi_gen3_rx_pcs_block_sync),
				.block_sync_sm(hssi_gen3_rx_pcs_block_sync_sm),
				.cdr_ctrl_force_unalgn(hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn),
				.lpbk_force(hssi_gen3_rx_pcs_lpbk_force),
				.mode(hssi_gen3_rx_pcs_mode),
				.rate_match_fifo(hssi_gen3_rx_pcs_rate_match_fifo),
				.rate_match_fifo_latency(hssi_gen3_rx_pcs_rate_match_fifo_latency),
				.reconfig_settings(hssi_gen3_rx_pcs_reconfig_settings),
				.reverse_lpbk(hssi_gen3_rx_pcs_reverse_lpbk),
				.rx_b4gb_par_lpbk(hssi_gen3_rx_pcs_rx_b4gb_par_lpbk),
				.rx_force_balign(hssi_gen3_rx_pcs_rx_force_balign),
				.rx_ins_del_one_skip(hssi_gen3_rx_pcs_rx_ins_del_one_skip),
				.rx_num_fixed_pat(hssi_gen3_rx_pcs_rx_num_fixed_pat),
				.rx_test_out_sel(hssi_gen3_rx_pcs_rx_test_out_sel),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_rx_pcs_sup_mode)
			) inst_twentynm_hssi_gen3_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_rx_pcs_avmmreaddata),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.blk_start(w_hssi_gen3_rx_pcs_blk_start),
				.blockselect(w_hssi_gen3_rx_pcs_blockselect),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.data_out(w_hssi_gen3_rx_pcs_data_out),
				.data_valid(w_hssi_gen3_rx_pcs_data_valid),
				.ei_det_int(w_hssi_gen3_rx_pcs_ei_det_int),
				.ei_partial_det_int(w_hssi_gen3_rx_pcs_ei_partial_det_int),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.i_det_int(w_hssi_gen3_rx_pcs_i_det_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data(w_hssi_gen3_rx_pcs_lpbk_data),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.mem_rx_fifo_rd_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr),
				.mem_rx_fifo_wr_clk(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.mem_rx_fifo_wr_data(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data),
				.mem_rx_fifo_wr_en(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.mem_rx_fifo_wr_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr),
				.mem_rx_fifo_wr_rst_n(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_test_out(w_hssi_gen3_rx_pcs_rx_test_out),
				.sync_hdr(w_hssi_gen3_rx_pcs_sync_hdr),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0]}),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.mem_rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_gen3[39], w_hssi_fifo_rx_pcs_data_out_gen3[38], w_hssi_fifo_rx_pcs_data_out_gen3[37], w_hssi_fifo_rx_pcs_data_out_gen3[36], w_hssi_fifo_rx_pcs_data_out_gen3[35], w_hssi_fifo_rx_pcs_data_out_gen3[34], w_hssi_fifo_rx_pcs_data_out_gen3[33], w_hssi_fifo_rx_pcs_data_out_gen3[32], w_hssi_fifo_rx_pcs_data_out_gen3[31], w_hssi_fifo_rx_pcs_data_out_gen3[30], w_hssi_fifo_rx_pcs_data_out_gen3[29], w_hssi_fifo_rx_pcs_data_out_gen3[28], w_hssi_fifo_rx_pcs_data_out_gen3[27], w_hssi_fifo_rx_pcs_data_out_gen3[26], w_hssi_fifo_rx_pcs_data_out_gen3[25], w_hssi_fifo_rx_pcs_data_out_gen3[24], w_hssi_fifo_rx_pcs_data_out_gen3[23], w_hssi_fifo_rx_pcs_data_out_gen3[22], w_hssi_fifo_rx_pcs_data_out_gen3[21], w_hssi_fifo_rx_pcs_data_out_gen3[20], w_hssi_fifo_rx_pcs_data_out_gen3[19], w_hssi_fifo_rx_pcs_data_out_gen3[18], w_hssi_fifo_rx_pcs_data_out_gen3[17], w_hssi_fifo_rx_pcs_data_out_gen3[16], w_hssi_fifo_rx_pcs_data_out_gen3[15], w_hssi_fifo_rx_pcs_data_out_gen3[14], w_hssi_fifo_rx_pcs_data_out_gen3[13], w_hssi_fifo_rx_pcs_data_out_gen3[12], w_hssi_fifo_rx_pcs_data_out_gen3[11], w_hssi_fifo_rx_pcs_data_out_gen3[10], w_hssi_fifo_rx_pcs_data_out_gen3[9], w_hssi_fifo_rx_pcs_data_out_gen3[8], w_hssi_fifo_rx_pcs_data_out_gen3[7], w_hssi_fifo_rx_pcs_data_out_gen3[6], w_hssi_fifo_rx_pcs_data_out_gen3[5], w_hssi_fifo_rx_pcs_data_out_gen3[4], w_hssi_fifo_rx_pcs_data_out_gen3[3], w_hssi_fifo_rx_pcs_data_out_gen3[2], w_hssi_fifo_rx_pcs_data_out_gen3[1], w_hssi_fifo_rx_pcs_data_out_gen3[0]}),
				.par_lpbk_b4gb_in({w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0]}),
				.par_lpbk_in({w_hssi_gen3_tx_pcs_par_lpbk_out[31], w_hssi_gen3_tx_pcs_par_lpbk_out[30], w_hssi_gen3_tx_pcs_par_lpbk_out[29], w_hssi_gen3_tx_pcs_par_lpbk_out[28], w_hssi_gen3_tx_pcs_par_lpbk_out[27], w_hssi_gen3_tx_pcs_par_lpbk_out[26], w_hssi_gen3_tx_pcs_par_lpbk_out[25], w_hssi_gen3_tx_pcs_par_lpbk_out[24], w_hssi_gen3_tx_pcs_par_lpbk_out[23], w_hssi_gen3_tx_pcs_par_lpbk_out[22], w_hssi_gen3_tx_pcs_par_lpbk_out[21], w_hssi_gen3_tx_pcs_par_lpbk_out[20], w_hssi_gen3_tx_pcs_par_lpbk_out[19], w_hssi_gen3_tx_pcs_par_lpbk_out[18], w_hssi_gen3_tx_pcs_par_lpbk_out[17], w_hssi_gen3_tx_pcs_par_lpbk_out[16], w_hssi_gen3_tx_pcs_par_lpbk_out[15], w_hssi_gen3_tx_pcs_par_lpbk_out[14], w_hssi_gen3_tx_pcs_par_lpbk_out[13], w_hssi_gen3_tx_pcs_par_lpbk_out[12], w_hssi_gen3_tx_pcs_par_lpbk_out[11], w_hssi_gen3_tx_pcs_par_lpbk_out[10], w_hssi_gen3_tx_pcs_par_lpbk_out[9], w_hssi_gen3_tx_pcs_par_lpbk_out[8], w_hssi_gen3_tx_pcs_par_lpbk_out[7], w_hssi_gen3_tx_pcs_par_lpbk_out[6], w_hssi_gen3_tx_pcs_par_lpbk_out[5], w_hssi_gen3_tx_pcs_par_lpbk_out[4], w_hssi_gen3_tx_pcs_par_lpbk_out[3], w_hssi_gen3_tx_pcs_par_lpbk_out[2], w_hssi_gen3_tx_pcs_par_lpbk_out[1], w_hssi_gen3_tx_pcs_par_lpbk_out[0]}),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.rcvd_clk(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_pma_clk(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.rxpolarity(w_hssi_pipe_gen3_rxpolarity_int),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.sync_sm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.txdatak_in({w_hssi_pipe_gen3_txdatak_int[3], w_hssi_pipe_gen3_txdatak_int[2], w_hssi_pipe_gen3_txdatak_int[1], w_hssi_pipe_gen3_txdatak_int[0]}),
				
				// UNUSED
				.blk_lockd_int(),
				.skp_det_int()
			);
		end // if generate
		else begin
				assign w_hssi_gen3_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_rx_pcs_blk_algnd_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_delete_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_insert_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_overfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_undfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_rx_pcs_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_partial_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_err_decode_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_i_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data[33:0] = 34'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39:0] = 40'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_rx_test_out[19:0] = 20'b0;
				assign w_hssi_gen3_rx_pcs_sync_hdr[1:0] = 2'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_tx_pcs
			twentynm_hssi_gen3_tx_pcs #(
				.mode(hssi_gen3_tx_pcs_mode),
				.reverse_lpbk(hssi_gen3_tx_pcs_reverse_lpbk),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_tx_pcs_sup_mode),
				.tx_bitslip(hssi_gen3_tx_pcs_tx_bitslip),
				.tx_gbox_byp(hssi_gen3_tx_pcs_tx_gbox_byp)
			) inst_twentynm_hssi_gen3_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_gen3_tx_pcs_blockselect),
				.data_out(w_hssi_gen3_tx_pcs_data_out),
				.par_lpbk_b4gb_out(w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out),
				.par_lpbk_out(w_hssi_gen3_tx_pcs_par_lpbk_out),
				.tx_test_out(w_hssi_gen3_tx_pcs_tx_test_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_start_in(w_hssi_pipe_gen3_tx_blk_start_int),
				.data_in({w_hssi_pipe_gen3_txdata_int[31], w_hssi_pipe_gen3_txdata_int[30], w_hssi_pipe_gen3_txdata_int[29], w_hssi_pipe_gen3_txdata_int[28], w_hssi_pipe_gen3_txdata_int[27], w_hssi_pipe_gen3_txdata_int[26], w_hssi_pipe_gen3_txdata_int[25], w_hssi_pipe_gen3_txdata_int[24], w_hssi_pipe_gen3_txdata_int[23], w_hssi_pipe_gen3_txdata_int[22], w_hssi_pipe_gen3_txdata_int[21], w_hssi_pipe_gen3_txdata_int[20], w_hssi_pipe_gen3_txdata_int[19], w_hssi_pipe_gen3_txdata_int[18], w_hssi_pipe_gen3_txdata_int[17], w_hssi_pipe_gen3_txdata_int[16], w_hssi_pipe_gen3_txdata_int[15], w_hssi_pipe_gen3_txdata_int[14], w_hssi_pipe_gen3_txdata_int[13], w_hssi_pipe_gen3_txdata_int[12], w_hssi_pipe_gen3_txdata_int[11], w_hssi_pipe_gen3_txdata_int[10], w_hssi_pipe_gen3_txdata_int[9], w_hssi_pipe_gen3_txdata_int[8], w_hssi_pipe_gen3_txdata_int[7], w_hssi_pipe_gen3_txdata_int[6], w_hssi_pipe_gen3_txdata_int[5], w_hssi_pipe_gen3_txdata_int[4], w_hssi_pipe_gen3_txdata_int[3], w_hssi_pipe_gen3_txdata_int[2], w_hssi_pipe_gen3_txdata_int[1], w_hssi_pipe_gen3_txdata_int[0]}),
				.data_valid(w_hssi_pipe_gen3_txdataskip_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data_in({w_hssi_gen3_rx_pcs_lpbk_data[33], w_hssi_gen3_rx_pcs_lpbk_data[32], w_hssi_gen3_rx_pcs_lpbk_data[31], w_hssi_gen3_rx_pcs_lpbk_data[30], w_hssi_gen3_rx_pcs_lpbk_data[29], w_hssi_gen3_rx_pcs_lpbk_data[28], w_hssi_gen3_rx_pcs_lpbk_data[27], w_hssi_gen3_rx_pcs_lpbk_data[26], w_hssi_gen3_rx_pcs_lpbk_data[25], w_hssi_gen3_rx_pcs_lpbk_data[24], w_hssi_gen3_rx_pcs_lpbk_data[23], w_hssi_gen3_rx_pcs_lpbk_data[22], w_hssi_gen3_rx_pcs_lpbk_data[21], w_hssi_gen3_rx_pcs_lpbk_data[20], w_hssi_gen3_rx_pcs_lpbk_data[19], w_hssi_gen3_rx_pcs_lpbk_data[18], w_hssi_gen3_rx_pcs_lpbk_data[17], w_hssi_gen3_rx_pcs_lpbk_data[16], w_hssi_gen3_rx_pcs_lpbk_data[15], w_hssi_gen3_rx_pcs_lpbk_data[14], w_hssi_gen3_rx_pcs_lpbk_data[13], w_hssi_gen3_rx_pcs_lpbk_data[12], w_hssi_gen3_rx_pcs_lpbk_data[11], w_hssi_gen3_rx_pcs_lpbk_data[10], w_hssi_gen3_rx_pcs_lpbk_data[9], w_hssi_gen3_rx_pcs_lpbk_data[8], w_hssi_gen3_rx_pcs_lpbk_data[7], w_hssi_gen3_rx_pcs_lpbk_data[6], w_hssi_gen3_rx_pcs_lpbk_data[5], w_hssi_gen3_rx_pcs_lpbk_data[4], w_hssi_gen3_rx_pcs_lpbk_data[3], w_hssi_gen3_rx_pcs_lpbk_data[2], w_hssi_gen3_rx_pcs_lpbk_data[1], w_hssi_gen3_rx_pcs_lpbk_data[0]}),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.sync_in({w_hssi_pipe_gen3_tx_sync_hdr_int[1], w_hssi_pipe_gen3_tx_sync_hdr_int[0]}),
				.tx_pma_clk(w_hssi_8g_tx_pcs_clk_out_gen3),
				.tx_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn)
			);
		end // if generate
		else begin
				assign w_hssi_gen3_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_tx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_tx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35:0] = 36'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_tx_test_out[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_rx_pcs
			twentynm_hssi_krfec_rx_pcs #(
				.blksync_cor_en(hssi_krfec_rx_pcs_blksync_cor_en),
				.bypass_gb(hssi_krfec_rx_pcs_bypass_gb),
				.clr_ctrl(hssi_krfec_rx_pcs_clr_ctrl),
				.ctrl_bit_reverse(hssi_krfec_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_rx_pcs_data_bit_reverse),
				.dv_start(hssi_krfec_rx_pcs_dv_start),
				.err_mark_type(hssi_krfec_rx_pcs_err_mark_type),
				.error_marking_en(hssi_krfec_rx_pcs_error_marking_en),
				.low_latency_en(hssi_krfec_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_krfec_rx_pcs_lpbk_mode),
				.parity_invalid_enum(hssi_krfec_rx_pcs_parity_invalid_enum),
				.parity_valid_num(hssi_krfec_rx_pcs_parity_valid_num),
				.pipeln_blksync(hssi_krfec_rx_pcs_pipeln_blksync),
				.pipeln_descrm(hssi_krfec_rx_pcs_pipeln_descrm),
				.pipeln_errcorrect(hssi_krfec_rx_pcs_pipeln_errcorrect),
				.pipeln_errtrap_ind(hssi_krfec_rx_pcs_pipeln_errtrap_ind),
				.pipeln_errtrap_lfsr(hssi_krfec_rx_pcs_pipeln_errtrap_lfsr),
				.pipeln_errtrap_loc(hssi_krfec_rx_pcs_pipeln_errtrap_loc),
				.pipeln_errtrap_pat(hssi_krfec_rx_pcs_pipeln_errtrap_pat),
				.pipeln_gearbox(hssi_krfec_rx_pcs_pipeln_gearbox),
				.pipeln_syndrm(hssi_krfec_rx_pcs_pipeln_syndrm),
				.pipeln_trans_dec(hssi_krfec_rx_pcs_pipeln_trans_dec),
				.prot_mode(hssi_krfec_rx_pcs_prot_mode),
				.receive_order(hssi_krfec_rx_pcs_receive_order),
				.reconfig_settings(hssi_krfec_rx_pcs_reconfig_settings),
				.rx_testbus_sel(hssi_krfec_rx_pcs_rx_testbus_sel),
				.signal_ok_en(hssi_krfec_rx_pcs_signal_ok_en),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_rx_pcs_sup_mode)
			) inst_twentynm_hssi_krfec_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_rx_pcs_blockselect),
				.rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.rx_control_out(w_hssi_krfec_rx_pcs_rx_control_out),
				.rx_data_out(w_hssi_krfec_rx_pcs_rx_data_out),
				.rx_data_status(w_hssi_krfec_rx_pcs_rx_data_status),
				.rx_data_valid_out(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.rx_signal_ok_out(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.rx_data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0]}),
				.rx_krfec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_krfec_reg(),
				.pld_10g_krfec_rx_blk_lock_krfec_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg(),
				.pld_10g_krfec_rx_frame_krfec_reg(),
				.pld_10g_krfec_rx_frame_krfec_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_rx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_block_lock = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_control_out[9:0] = 10'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_status[1:0] = 2'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_valid_out = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_frame = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_signal_ok_out = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_tx_pcs
			twentynm_hssi_krfec_tx_pcs #(
				.burst_err(hssi_krfec_tx_pcs_burst_err),
				.burst_err_len(hssi_krfec_tx_pcs_burst_err_len),
				.ctrl_bit_reverse(hssi_krfec_tx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_tx_pcs_data_bit_reverse),
				.enc_frame_query(hssi_krfec_tx_pcs_enc_frame_query),
				.low_latency_en(hssi_krfec_tx_pcs_low_latency_en),
				.pipeln_encoder(hssi_krfec_tx_pcs_pipeln_encoder),
				.pipeln_scrambler(hssi_krfec_tx_pcs_pipeln_scrambler),
				.prot_mode(hssi_krfec_tx_pcs_prot_mode),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_tx_pcs_sup_mode),
				.transcode_err(hssi_krfec_tx_pcs_transcode_err),
				.transmit_order(hssi_krfec_tx_pcs_transmit_order),
				.tx_testbus_sel(hssi_krfec_tx_pcs_tx_testbus_sel)
			) inst_twentynm_hssi_krfec_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_tx_pcs_blockselect),
				.tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.tx_data_out(w_hssi_krfec_tx_pcs_tx_data_out),
				.tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.tx_test_data(w_hssi_krfec_tx_pcs_tx_test_data),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.tx_control_in({w_hssi_10g_tx_pcs_tx_control_out_krfec[8], w_hssi_10g_tx_pcs_tx_control_out_krfec[7], w_hssi_10g_tx_pcs_tx_control_out_krfec[6], w_hssi_10g_tx_pcs_tx_control_out_krfec[5], w_hssi_10g_tx_pcs_tx_control_out_krfec[4], w_hssi_10g_tx_pcs_tx_control_out_krfec[3], w_hssi_10g_tx_pcs_tx_control_out_krfec[2], w_hssi_10g_tx_pcs_tx_control_out_krfec[1], w_hssi_10g_tx_pcs_tx_control_out_krfec[0]}),
				.tx_data_in({w_hssi_10g_tx_pcs_tx_data_out_krfec[63], w_hssi_10g_tx_pcs_tx_data_out_krfec[62], w_hssi_10g_tx_pcs_tx_data_out_krfec[61], w_hssi_10g_tx_pcs_tx_data_out_krfec[60], w_hssi_10g_tx_pcs_tx_data_out_krfec[59], w_hssi_10g_tx_pcs_tx_data_out_krfec[58], w_hssi_10g_tx_pcs_tx_data_out_krfec[57], w_hssi_10g_tx_pcs_tx_data_out_krfec[56], w_hssi_10g_tx_pcs_tx_data_out_krfec[55], w_hssi_10g_tx_pcs_tx_data_out_krfec[54], w_hssi_10g_tx_pcs_tx_data_out_krfec[53], w_hssi_10g_tx_pcs_tx_data_out_krfec[52], w_hssi_10g_tx_pcs_tx_data_out_krfec[51], w_hssi_10g_tx_pcs_tx_data_out_krfec[50], w_hssi_10g_tx_pcs_tx_data_out_krfec[49], w_hssi_10g_tx_pcs_tx_data_out_krfec[48], w_hssi_10g_tx_pcs_tx_data_out_krfec[47], w_hssi_10g_tx_pcs_tx_data_out_krfec[46], w_hssi_10g_tx_pcs_tx_data_out_krfec[45], w_hssi_10g_tx_pcs_tx_data_out_krfec[44], w_hssi_10g_tx_pcs_tx_data_out_krfec[43], w_hssi_10g_tx_pcs_tx_data_out_krfec[42], w_hssi_10g_tx_pcs_tx_data_out_krfec[41], w_hssi_10g_tx_pcs_tx_data_out_krfec[40], w_hssi_10g_tx_pcs_tx_data_out_krfec[39], w_hssi_10g_tx_pcs_tx_data_out_krfec[38], w_hssi_10g_tx_pcs_tx_data_out_krfec[37], w_hssi_10g_tx_pcs_tx_data_out_krfec[36], w_hssi_10g_tx_pcs_tx_data_out_krfec[35], w_hssi_10g_tx_pcs_tx_data_out_krfec[34], w_hssi_10g_tx_pcs_tx_data_out_krfec[33], w_hssi_10g_tx_pcs_tx_data_out_krfec[32], w_hssi_10g_tx_pcs_tx_data_out_krfec[31], w_hssi_10g_tx_pcs_tx_data_out_krfec[30], w_hssi_10g_tx_pcs_tx_data_out_krfec[29], w_hssi_10g_tx_pcs_tx_data_out_krfec[28], w_hssi_10g_tx_pcs_tx_data_out_krfec[27], w_hssi_10g_tx_pcs_tx_data_out_krfec[26], w_hssi_10g_tx_pcs_tx_data_out_krfec[25], w_hssi_10g_tx_pcs_tx_data_out_krfec[24], w_hssi_10g_tx_pcs_tx_data_out_krfec[23], w_hssi_10g_tx_pcs_tx_data_out_krfec[22], w_hssi_10g_tx_pcs_tx_data_out_krfec[21], w_hssi_10g_tx_pcs_tx_data_out_krfec[20], w_hssi_10g_tx_pcs_tx_data_out_krfec[19], w_hssi_10g_tx_pcs_tx_data_out_krfec[18], w_hssi_10g_tx_pcs_tx_data_out_krfec[17], w_hssi_10g_tx_pcs_tx_data_out_krfec[16], w_hssi_10g_tx_pcs_tx_data_out_krfec[15], w_hssi_10g_tx_pcs_tx_data_out_krfec[14], w_hssi_10g_tx_pcs_tx_data_out_krfec[13], w_hssi_10g_tx_pcs_tx_data_out_krfec[12], w_hssi_10g_tx_pcs_tx_data_out_krfec[11], w_hssi_10g_tx_pcs_tx_data_out_krfec[10], w_hssi_10g_tx_pcs_tx_data_out_krfec[9], w_hssi_10g_tx_pcs_tx_data_out_krfec[8], w_hssi_10g_tx_pcs_tx_data_out_krfec[7], w_hssi_10g_tx_pcs_tx_data_out_krfec[6], w_hssi_10g_tx_pcs_tx_data_out_krfec[5], w_hssi_10g_tx_pcs_tx_data_out_krfec[4], w_hssi_10g_tx_pcs_tx_data_out_krfec[3], w_hssi_10g_tx_pcs_tx_data_out_krfec[2], w_hssi_10g_tx_pcs_tx_data_out_krfec[1], w_hssi_10g_tx_pcs_tx_data_out_krfec[0]}),
				.tx_data_valid_in(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_krfec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_krfec_reg(),
				.pld_krfec_tx_alignment_plddirect_reg(),
				.pld_krfec_tx_alignment_reg()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_tx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_alignment = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_test_data[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen1_2
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen1_2
			twentynm_hssi_pipe_gen1_2 #(
				.elec_idle_delay_val(hssi_pipe_gen1_2_elec_idle_delay_val),
				.error_replace_pad(hssi_pipe_gen1_2_error_replace_pad),
				.hip_mode(hssi_pipe_gen1_2_hip_mode),
				.ind_error_reporting(hssi_pipe_gen1_2_ind_error_reporting),
				.phystatus_delay_val(hssi_pipe_gen1_2_phystatus_delay_val),
				.phystatus_rst_toggle(hssi_pipe_gen1_2_phystatus_rst_toggle),
				.pipe_byte_de_serializer_en(hssi_pipe_gen1_2_pipe_byte_de_serializer_en),
				.prot_mode(hssi_pipe_gen1_2_prot_mode),
				.reconfig_settings(hssi_pipe_gen1_2_reconfig_settings),
				.rx_pipe_enable(hssi_pipe_gen1_2_rx_pipe_enable),
				.rxdetect_bypass(hssi_pipe_gen1_2_rxdetect_bypass),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen1_2_sup_mode),
				.tx_pipe_enable(hssi_pipe_gen1_2_tx_pipe_enable),
				.txswing(hssi_pipe_gen1_2_txswing)
			) inst_twentynm_hssi_pipe_gen1_2 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen1_2_avmmreaddata),
				.blockselect(w_hssi_pipe_gen1_2_blockselect),
				.current_coeff(w_hssi_pipe_gen1_2_current_coeff),
				.phystatus(w_hssi_pipe_gen1_2_phystatus),
				.polarity_inversion_rx(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rev_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.rxelectricalidle_out(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxstatus(w_hssi_pipe_gen1_2_rxstatus),
				.rxvalid(w_hssi_pipe_gen1_2_rxvalid),
				.tx_elec_idle_out(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pipe_rx_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.power_state_transition_done_ena(1'b0),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rev_loopbk_pcs_gen3(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.revloopback(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.rx_pipe_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rxd({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxelectricalidle(w_hssi_8g_rx_pcs_eidle_detected),
				.rxelectricalidle_pcs_gen3(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.rxpolarity_pcs_gen3(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.tx_elec_idle_comp(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.txd_ch({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswingport(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.pld_8g_rxpolarity_pipe3_reg(),
				.rxd_ch(),
				.txd()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen1_2_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen1_2_blockselect = 1'b0;
				assign w_hssi_pipe_gen1_2_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen1_2_phystatus = 1'b0;
				assign w_hssi_pipe_gen1_2_polarity_inversion_rx = 1'b0;
				assign w_hssi_pipe_gen1_2_rev_loopbk = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelectricalidle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen1_2_rxvalid = 1'b0;
				assign w_hssi_pipe_gen1_2_tx_elec_idle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_txdetectrx = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen3
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen3
			twentynm_hssi_pipe_gen3 #(
				.bypass_rx_detection_enable(hssi_pipe_gen3_bypass_rx_detection_enable),
				.bypass_rx_preset(hssi_pipe_gen3_bypass_rx_preset),
				.bypass_rx_preset_enable(hssi_pipe_gen3_bypass_rx_preset_enable),
				.bypass_tx_coefficent(hssi_pipe_gen3_bypass_tx_coefficent),
				.bypass_tx_coefficent_enable(hssi_pipe_gen3_bypass_tx_coefficent_enable),
				.elecidle_delay_g3(hssi_pipe_gen3_elecidle_delay_g3),
				.ind_error_reporting(hssi_pipe_gen3_ind_error_reporting),
				.mode(hssi_pipe_gen3_mode),
				.phy_status_delay_g12(hssi_pipe_gen3_phy_status_delay_g12),
				.phy_status_delay_g3(hssi_pipe_gen3_phy_status_delay_g3),
				.phystatus_rst_toggle_g12(hssi_pipe_gen3_phystatus_rst_toggle_g12),
				.phystatus_rst_toggle_g3(hssi_pipe_gen3_phystatus_rst_toggle_g3),
				.rate_match_pad_insertion(hssi_pipe_gen3_rate_match_pad_insertion),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen3_sup_mode),
				.test_out_sel(hssi_pipe_gen3_test_out_sel)
			) inst_twentynm_hssi_pipe_gen3 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen3_avmmreaddata),
				.blockselect(w_hssi_pipe_gen3_blockselect),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.phystatus(w_hssi_pipe_gen3_phystatus),
				.pma_current_coeff(w_hssi_pipe_gen3_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_pipe_gen3_pma_current_rxpreset),
				.pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.rev_lpbk_8gpcs_out(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.rev_lpbk_int(w_hssi_pipe_gen3_rev_lpbk_int),
				.rx_blk_start(w_hssi_pipe_gen3_rx_blk_start),
				.rx_sync_hdr(w_hssi_pipe_gen3_rx_sync_hdr),
				.rxd_8gpcs_out(w_hssi_pipe_gen3_rxd_8gpcs_out),
				.rxdataskip(w_hssi_pipe_gen3_rxdataskip),
				.rxelecidle(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity_8gpcs_out(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.rxpolarity_int(w_hssi_pipe_gen3_rxpolarity_int),
				.rxstatus(w_hssi_pipe_gen3_rxstatus),
				.rxvalid(w_hssi_pipe_gen3_rxvalid),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.test_out(w_hssi_pipe_gen3_test_out),
				.tx_blk_start_int(w_hssi_pipe_gen3_tx_blk_start_int),
				.tx_sync_hdr_int(w_hssi_pipe_gen3_tx_sync_hdr_int),
				.txdata_int(w_hssi_pipe_gen3_txdata_int),
				.txdatak_int(w_hssi_pipe_gen3_txdatak_int),
				.txdataskip_int(w_hssi_pipe_gen3_txdataskip_int),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.current_coeff({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0]}),
				.current_rxpreset({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0]}),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.pcs_asn_bundling_in({w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0]}),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pipe_tx_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_blk_start_int(w_hssi_gen3_rx_pcs_blk_start),
				.rx_sync_hdr_int({w_hssi_gen3_rx_pcs_sync_hdr[1], w_hssi_gen3_rx_pcs_sync_hdr[0]}),
				.rx_test_out({w_hssi_gen3_rx_pcs_rx_test_out[19], w_hssi_gen3_rx_pcs_rx_test_out[18], w_hssi_gen3_rx_pcs_rx_test_out[17], w_hssi_gen3_rx_pcs_rx_test_out[16], w_hssi_gen3_rx_pcs_rx_test_out[15], w_hssi_gen3_rx_pcs_rx_test_out[14], w_hssi_gen3_rx_pcs_rx_test_out[13], w_hssi_gen3_rx_pcs_rx_test_out[12], w_hssi_gen3_rx_pcs_rx_test_out[11], w_hssi_gen3_rx_pcs_rx_test_out[10], w_hssi_gen3_rx_pcs_rx_test_out[9], w_hssi_gen3_rx_pcs_rx_test_out[8], w_hssi_gen3_rx_pcs_rx_test_out[7], w_hssi_gen3_rx_pcs_rx_test_out[6], w_hssi_gen3_rx_pcs_rx_test_out[5], w_hssi_gen3_rx_pcs_rx_test_out[4], w_hssi_gen3_rx_pcs_rx_test_out[3], w_hssi_gen3_rx_pcs_rx_test_out[2], w_hssi_gen3_rx_pcs_rx_test_out[1], w_hssi_gen3_rx_pcs_rx_test_out[0]}),
				.rxd_8gpcs_in({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxdata_int({w_hssi_gen3_rx_pcs_data_out[31], w_hssi_gen3_rx_pcs_data_out[30], w_hssi_gen3_rx_pcs_data_out[29], w_hssi_gen3_rx_pcs_data_out[28], w_hssi_gen3_rx_pcs_data_out[27], w_hssi_gen3_rx_pcs_data_out[26], w_hssi_gen3_rx_pcs_data_out[25], w_hssi_gen3_rx_pcs_data_out[24], w_hssi_gen3_rx_pcs_data_out[23], w_hssi_gen3_rx_pcs_data_out[22], w_hssi_gen3_rx_pcs_data_out[21], w_hssi_gen3_rx_pcs_data_out[20], w_hssi_gen3_rx_pcs_data_out[19], w_hssi_gen3_rx_pcs_data_out[18], w_hssi_gen3_rx_pcs_data_out[17], w_hssi_gen3_rx_pcs_data_out[16], w_hssi_gen3_rx_pcs_data_out[15], w_hssi_gen3_rx_pcs_data_out[14], w_hssi_gen3_rx_pcs_data_out[13], w_hssi_gen3_rx_pcs_data_out[12], w_hssi_gen3_rx_pcs_data_out[11], w_hssi_gen3_rx_pcs_data_out[10], w_hssi_gen3_rx_pcs_data_out[9], w_hssi_gen3_rx_pcs_data_out[8], w_hssi_gen3_rx_pcs_data_out[7], w_hssi_gen3_rx_pcs_data_out[6], w_hssi_gen3_rx_pcs_data_out[5], w_hssi_gen3_rx_pcs_data_out[4], w_hssi_gen3_rx_pcs_data_out[3], w_hssi_gen3_rx_pcs_data_out[2], w_hssi_gen3_rx_pcs_data_out[1], w_hssi_gen3_rx_pcs_data_out[0]}),
				.rxdatak_int({1'b0, 1'b0, 1'b0, 1'b0}),
				.rxdataskip_int(w_hssi_gen3_rx_pcs_data_valid),
				.rxelecidle_8gpcs_in(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.tx_blk_start(w_hssi_8g_tx_pcs_tx_blk_start_out[0]),
				.tx_sync_hdr({w_hssi_8g_tx_pcs_tx_sync_hdr_out[1], w_hssi_8g_tx_pcs_tx_sync_hdr_out[0]}),
				.tx_test_out({w_hssi_gen3_tx_pcs_tx_test_out[19], w_hssi_gen3_tx_pcs_tx_test_out[18], w_hssi_gen3_tx_pcs_tx_test_out[17], w_hssi_gen3_tx_pcs_tx_test_out[16], w_hssi_gen3_tx_pcs_tx_test_out[15], w_hssi_gen3_tx_pcs_tx_test_out[14], w_hssi_gen3_tx_pcs_tx_test_out[13], w_hssi_gen3_tx_pcs_tx_test_out[12], w_hssi_gen3_tx_pcs_tx_test_out[11], w_hssi_gen3_tx_pcs_tx_test_out[10], w_hssi_gen3_tx_pcs_tx_test_out[9], w_hssi_gen3_tx_pcs_tx_test_out[8], w_hssi_gen3_tx_pcs_tx_test_out[7], w_hssi_gen3_tx_pcs_tx_test_out[6], w_hssi_gen3_tx_pcs_tx_test_out[5], w_hssi_gen3_tx_pcs_tx_test_out[4], w_hssi_gen3_tx_pcs_tx_test_out[3], w_hssi_gen3_tx_pcs_tx_test_out[2], w_hssi_gen3_tx_pcs_tx_test_out[1], w_hssi_gen3_tx_pcs_tx_test_out[0]}),
				.txcompliance(w_hssi_8g_tx_pcs_txcompliance_out),
				.txdata({w_hssi_8g_tx_pcs_tx_data_out[31], w_hssi_8g_tx_pcs_tx_data_out[30], w_hssi_8g_tx_pcs_tx_data_out[29], w_hssi_8g_tx_pcs_tx_data_out[28], w_hssi_8g_tx_pcs_tx_data_out[27], w_hssi_8g_tx_pcs_tx_data_out[26], w_hssi_8g_tx_pcs_tx_data_out[25], w_hssi_8g_tx_pcs_tx_data_out[24], w_hssi_8g_tx_pcs_tx_data_out[23], w_hssi_8g_tx_pcs_tx_data_out[22], w_hssi_8g_tx_pcs_tx_data_out[21], w_hssi_8g_tx_pcs_tx_data_out[20], w_hssi_8g_tx_pcs_tx_data_out[19], w_hssi_8g_tx_pcs_tx_data_out[18], w_hssi_8g_tx_pcs_tx_data_out[17], w_hssi_8g_tx_pcs_tx_data_out[16], w_hssi_8g_tx_pcs_tx_data_out[15], w_hssi_8g_tx_pcs_tx_data_out[14], w_hssi_8g_tx_pcs_tx_data_out[13], w_hssi_8g_tx_pcs_tx_data_out[12], w_hssi_8g_tx_pcs_tx_data_out[11], w_hssi_8g_tx_pcs_tx_data_out[10], w_hssi_8g_tx_pcs_tx_data_out[9], w_hssi_8g_tx_pcs_tx_data_out[8], w_hssi_8g_tx_pcs_tx_data_out[7], w_hssi_8g_tx_pcs_tx_data_out[6], w_hssi_8g_tx_pcs_tx_data_out[5], w_hssi_8g_tx_pcs_tx_data_out[4], w_hssi_8g_tx_pcs_tx_data_out[3], w_hssi_8g_tx_pcs_tx_data_out[2], w_hssi_8g_tx_pcs_tx_data_out[1], w_hssi_8g_tx_pcs_tx_data_out[0]}),
				.txdatak({w_hssi_8g_tx_pcs_tx_datak_out[3], w_hssi_8g_tx_pcs_tx_datak_out[2], w_hssi_8g_tx_pcs_tx_datak_out[1], w_hssi_8g_tx_pcs_tx_datak_out[0]}),
				.txdataskip(w_hssi_8g_tx_pcs_tx_data_valid_out[0]),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_8g_tx_pcs_txelecidle_out),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.dis_pc_byte(),
				.pma_rx_det_pd(),
				.pma_txdeemph(),
				.pma_txmargin(),
				.pma_txswing(),
				.reset_pc_prts()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen3_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen3_blockselect = 1'b0;
				assign w_hssi_pipe_gen3_gen3_clk_sel = 1'b0;
				assign w_hssi_pipe_gen3_pcs_rst = 1'b0;
				assign w_hssi_pipe_gen3_phystatus = 1'b0;
				assign w_hssi_pipe_gen3_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen3_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_pma_tx_elec_idle = 1'b0;
				assign w_hssi_pipe_gen3_pma_txdetectrx = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_int = 1'b0;
				assign w_hssi_pipe_gen3_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_rxd_8gpcs_out[63:0] = 64'b0;
				assign w_hssi_pipe_gen3_rxdataskip[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_int = 1'b0;
				assign w_hssi_pipe_gen3_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_rxvalid = 1'b0;
				assign w_hssi_pipe_gen3_shutdown_clk = 1'b0;
				assign w_hssi_pipe_gen3_test_out[19:0] = 20'b0;
				assign w_hssi_pipe_gen3_tx_blk_start_int = 1'b0;
				assign w_hssi_pipe_gen3_tx_sync_hdr_int[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_txdata_int[31:0] = 32'b0;
				assign w_hssi_pipe_gen3_txdatak_int[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_txdataskip_int = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pcs_pma_interface
			twentynm_hssi_rx_pcs_pma_interface #(
				.block_sel(hssi_rx_pcs_pma_interface_block_sel),
				.channel_operation_mode(hssi_rx_pcs_pma_interface_channel_operation_mode),
				.clkslip_sel(hssi_rx_pcs_pma_interface_clkslip_sel),
				.lpbk_en(hssi_rx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_rx_pcs_pma_interface_master_clk_sel),
				.pldif_datawidth_mode(hssi_rx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_rx(hssi_rx_pcs_pma_interface_pma_dw_rx),
				.pma_if_dft_en(hssi_rx_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_rx_pcs_pma_interface_pma_if_dft_val),
				.prbs9_dwidth(hssi_rx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_rx_pcs_pma_interface_prbs_clken),
				.prbs_ver(hssi_rx_pcs_pma_interface_prbs_ver),
				.prot_mode_rx(hssi_rx_pcs_pma_interface_prot_mode_rx),
				.reconfig_settings(hssi_rx_pcs_pma_interface_reconfig_settings),
				.rx_dyn_polarity_inversion(hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion),
				.rx_lpbk_en(hssi_rx_pcs_pma_interface_rx_lpbk_en),
				.rx_prbs_force_signal_ok(hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok),
				.rx_prbs_mask(hssi_rx_pcs_pma_interface_rx_prbs_mask),
				.rx_prbs_mode(hssi_rx_pcs_pma_interface_rx_prbs_mode),
				.rx_signalok_signaldet_sel(hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel),
				.rx_static_polarity_inversion(hssi_rx_pcs_pma_interface_rx_static_polarity_inversion),
				.rx_uhsif_lpbk_en(hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sup_mode(hssi_rx_pcs_pma_interface_sup_mode)
			) inst_twentynm_hssi_rx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.int_pmaif_10g_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data),
				.int_pmaif_10g_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.int_pmaif_8g_pudi(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi),
				.int_pmaif_8g_rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.int_pmaif_8g_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.int_pmaif_8g_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.int_pmaif_8g_sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.int_pmaif_g3_pma_data_in(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in),
				.int_pmaif_g3_pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.int_pmaif_g3_pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.int_pmaif_g3_pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.int_pmaif_krfec_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data),
				.int_pmaif_krfec_rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.int_pmaif_pldif_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pmaif_pldif_prbs_err_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pmaif_pldif_rx_clkdiv(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pmaif_pldif_rx_clkdiv_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pmaif_pldif_rx_data(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data),
				.int_pmaif_pldif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pmaif_pldif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pmaif_pldif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pmaif_pldif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.pma_eye_monitor(w_hssi_rx_pcs_pma_interface_pma_eye_monitor),
				.pma_rx_clkslip(w_hssi_rx_pcs_pma_interface_pma_rx_clkslip),
				.pma_rxpma_rstb(w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb),
				.rx_pmaif_test_out(w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out),
				.rx_prbs_ver_test(w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.int_pmaif_8g_rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.int_pmaif_pldif_eye_monitor({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0]}),
				.int_pmaif_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pmaif_pldif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pmaif_pldif_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pmaif_pldif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pma_rx_clkdiv_user(in_pma_rx_clkdiv_user),
				.pma_rx_detect_valid(in_pma_rx_detect_valid),
				.pma_rx_found(in_pma_rx_found),
				.pma_rx_pma_clk(in_pma_rx_pma_clk),
				.pma_rx_pma_data({in_pma_rx_pma_data[63], in_pma_rx_pma_data[62], in_pma_rx_pma_data[61], in_pma_rx_pma_data[60], in_pma_rx_pma_data[59], in_pma_rx_pma_data[58], in_pma_rx_pma_data[57], in_pma_rx_pma_data[56], in_pma_rx_pma_data[55], in_pma_rx_pma_data[54], in_pma_rx_pma_data[53], in_pma_rx_pma_data[52], in_pma_rx_pma_data[51], in_pma_rx_pma_data[50], in_pma_rx_pma_data[49], in_pma_rx_pma_data[48], in_pma_rx_pma_data[47], in_pma_rx_pma_data[46], in_pma_rx_pma_data[45], in_pma_rx_pma_data[44], in_pma_rx_pma_data[43], in_pma_rx_pma_data[42], in_pma_rx_pma_data[41], in_pma_rx_pma_data[40], in_pma_rx_pma_data[39], in_pma_rx_pma_data[38], in_pma_rx_pma_data[37], in_pma_rx_pma_data[36], in_pma_rx_pma_data[35], in_pma_rx_pma_data[34], in_pma_rx_pma_data[33], in_pma_rx_pma_data[32], in_pma_rx_pma_data[31], in_pma_rx_pma_data[30], in_pma_rx_pma_data[29], in_pma_rx_pma_data[28], in_pma_rx_pma_data[27], in_pma_rx_pma_data[26], in_pma_rx_pma_data[25], in_pma_rx_pma_data[24], in_pma_rx_pma_data[23], in_pma_rx_pma_data[22], in_pma_rx_pma_data[21], in_pma_rx_pma_data[20], in_pma_rx_pma_data[19], in_pma_rx_pma_data[18], in_pma_rx_pma_data[17], in_pma_rx_pma_data[16], in_pma_rx_pma_data[15], in_pma_rx_pma_data[14], in_pma_rx_pma_data[13], in_pma_rx_pma_data[12], in_pma_rx_pma_data[11], in_pma_rx_pma_data[10], in_pma_rx_pma_data[9], in_pma_rx_pma_data[8], in_pma_rx_pma_data[7], in_pma_rx_pma_data[6], in_pma_rx_pma_data[5], in_pma_rx_pma_data[4], in_pma_rx_pma_data[3], in_pma_rx_pma_data[2], in_pma_rx_pma_data[1], in_pma_rx_pma_data[0]}),
				.pma_rx_signal_ok(in_pma_rx_signal_ok),
				.pma_rxpll_lock(in_pma_rxpll_lock),
				.pma_signal_det(in_pma_signal_det),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.tx_pma_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0]}),
				.tx_pma_uhsif_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0]}),
				
				// UNUSED
				.int_pmaif_g3_rcvd_clk(),
				.prbs_err_lt()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31:0] = 32'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5:0] = 6'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rx_clkslip = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pld_pcs_interface
			twentynm_hssi_rx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx),
				.hd_10g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx),
				.hd_10g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx),
				.hd_10g_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx),
				.hd_10g_lpbk_en(hssi_rx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx),
				.hd_10g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx),
				.hd_10g_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx),
				.hd_10g_test_bus_mode(hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode),
				.hd_8g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx),
				.hd_8g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx),
				.hd_8g_hip_mode(hssi_rx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_rx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx),
				.hd_8g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx),
				.hd_chnl_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_clklow_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz),
				.hd_chnl_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx),
				.hd_chnl_fref_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz),
				.hd_chnl_frequency_rules_en(hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_rx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_rx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx),
				.hd_chnl_lpbk_en(hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx),
				.hd_chnl_pld_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz),
				.hd_chnl_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx),
				.hd_chnl_pma_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz),
				.hd_chnl_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx),
				.hd_chnl_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx),
				.hd_chnl_transparent_pcs_rx(hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx),
				.hd_fifo_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx),
				.hd_fifo_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx),
				.hd_g3_prot_mode(hssi_rx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx),
				.hd_krfec_lpbk_en(hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx),
				.hd_krfec_test_bus_mode(hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode),
				.hd_pldif_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx),
				.hd_pmaif_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_lpbk_en(hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx),
				.hd_pmaif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx),
				.hd_pmaif_sim_mode(hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_rx_block_sel(hssi_rx_pld_pcs_interface_pcs_rx_block_sel),
				.pcs_rx_clk_out_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel),
				.pcs_rx_clk_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_sel),
				.pcs_rx_hip_clk_en(hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en),
				.pcs_rx_output_sel(hssi_rx_pld_pcs_interface_pcs_rx_output_sel),
				.reconfig_settings(hssi_rx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm3" )       //PARAM_HIDE
			) inst_twentynm_hssi_rx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pld_pcs_interface_blockselect),
				.hip_rx_ctrl(w_hssi_rx_pld_pcs_interface_hip_rx_ctrl),
				.hip_rx_data(w_hssi_rx_pld_pcs_interface_hip_rx_data),
				.int_pldif_10g_rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.int_pldif_10g_rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.int_pldif_10g_rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.int_pldif_10g_rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.int_pldif_10g_rx_control_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb),
				.int_pldif_10g_rx_data_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb),
				.int_pldif_10g_rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.int_pldif_10g_rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.int_pldif_10g_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.int_pldif_10g_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.int_pldif_10g_rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.int_pldif_8g_a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.int_pldif_8g_bitloc_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.int_pldif_8g_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.int_pldif_8g_byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.int_pldif_8g_encdt(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.int_pldif_8g_pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.int_pldif_8g_rdenable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.int_pldif_8g_rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.int_pldif_8g_rxurstpcs_n(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.int_pldif_8g_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.int_pldif_8g_wrdisable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.int_pldif_g3_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.int_pldif_krfec_rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.int_pldif_pmaif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pldif_pmaif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pldif_pmaif_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pldif_pmaif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pld_10g_krfec_rx_blk_lock(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock),
				.pld_10g_krfec_rx_diag_data_status(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status),
				.pld_10g_krfec_rx_frame(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame),
				.pld_10g_rx_align_val(w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val),
				.pld_10g_rx_crc32_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err),
				.pld_10g_rx_data_valid(w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid),
				.pld_10g_rx_empty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty),
				.pld_10g_rx_fifo_del(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del),
				.pld_10g_rx_fifo_insert(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert),
				.pld_10g_rx_fifo_num(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num),
				.pld_10g_rx_frame_lock(w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock),
				.pld_10g_rx_hi_ber(w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber),
				.pld_10g_rx_oflw_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err),
				.pld_10g_rx_pempty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty),
				.pld_10g_rx_pfull(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull),
				.pld_8g_a1a2_k1k2_flag(w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag),
				.pld_8g_empty_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf),
				.pld_8g_empty_rx(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx),
				.pld_8g_full_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf),
				.pld_8g_full_rx(w_hssi_rx_pld_pcs_interface_pld_8g_full_rx),
				.pld_8g_rxelecidle(w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle),
				.pld_8g_signal_detect_out(w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out),
				.pld_8g_wa_boundary(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary),
				.pld_pcs_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out),
				.pld_pma_clkdiv_rx_user(w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user),
				.pld_pma_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out),
				.pld_pma_signal_ok(w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok),
				.pld_rx_control(w_hssi_rx_pld_pcs_interface_pld_rx_control),
				.pld_rx_data(w_hssi_rx_pld_pcs_interface_pld_rx_data),
				.pld_rx_prbs_done(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done),
				.pld_rx_prbs_err(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.int_pldif_10g_rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.int_pldif_10g_rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.int_pldif_10g_rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_10g_rx_control({w_hssi_10g_rx_pcs_rx_control[19], w_hssi_10g_rx_pcs_rx_control[18], w_hssi_10g_rx_pcs_rx_control[17], w_hssi_10g_rx_pcs_rx_control[16], w_hssi_10g_rx_pcs_rx_control[15], w_hssi_10g_rx_pcs_rx_control[14], w_hssi_10g_rx_pcs_rx_control[13], w_hssi_10g_rx_pcs_rx_control[12], w_hssi_10g_rx_pcs_rx_control[11], w_hssi_10g_rx_pcs_rx_control[10], w_hssi_10g_rx_pcs_rx_control[9], w_hssi_10g_rx_pcs_rx_control[8], w_hssi_10g_rx_pcs_rx_control[7], w_hssi_10g_rx_pcs_rx_control[6], w_hssi_10g_rx_pcs_rx_control[5], w_hssi_10g_rx_pcs_rx_control[4], w_hssi_10g_rx_pcs_rx_control[3], w_hssi_10g_rx_pcs_rx_control[2], w_hssi_10g_rx_pcs_rx_control[1], w_hssi_10g_rx_pcs_rx_control[0]}),
				.int_pldif_10g_rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.int_pldif_10g_rx_data({w_hssi_10g_rx_pcs_rx_data[127], w_hssi_10g_rx_pcs_rx_data[126], w_hssi_10g_rx_pcs_rx_data[125], w_hssi_10g_rx_pcs_rx_data[124], w_hssi_10g_rx_pcs_rx_data[123], w_hssi_10g_rx_pcs_rx_data[122], w_hssi_10g_rx_pcs_rx_data[121], w_hssi_10g_rx_pcs_rx_data[120], w_hssi_10g_rx_pcs_rx_data[119], w_hssi_10g_rx_pcs_rx_data[118], w_hssi_10g_rx_pcs_rx_data[117], w_hssi_10g_rx_pcs_rx_data[116], w_hssi_10g_rx_pcs_rx_data[115], w_hssi_10g_rx_pcs_rx_data[114], w_hssi_10g_rx_pcs_rx_data[113], w_hssi_10g_rx_pcs_rx_data[112], w_hssi_10g_rx_pcs_rx_data[111], w_hssi_10g_rx_pcs_rx_data[110], w_hssi_10g_rx_pcs_rx_data[109], w_hssi_10g_rx_pcs_rx_data[108], w_hssi_10g_rx_pcs_rx_data[107], w_hssi_10g_rx_pcs_rx_data[106], w_hssi_10g_rx_pcs_rx_data[105], w_hssi_10g_rx_pcs_rx_data[104], w_hssi_10g_rx_pcs_rx_data[103], w_hssi_10g_rx_pcs_rx_data[102], w_hssi_10g_rx_pcs_rx_data[101], w_hssi_10g_rx_pcs_rx_data[100], w_hssi_10g_rx_pcs_rx_data[99], w_hssi_10g_rx_pcs_rx_data[98], w_hssi_10g_rx_pcs_rx_data[97], w_hssi_10g_rx_pcs_rx_data[96], w_hssi_10g_rx_pcs_rx_data[95], w_hssi_10g_rx_pcs_rx_data[94], w_hssi_10g_rx_pcs_rx_data[93], w_hssi_10g_rx_pcs_rx_data[92], w_hssi_10g_rx_pcs_rx_data[91], w_hssi_10g_rx_pcs_rx_data[90], w_hssi_10g_rx_pcs_rx_data[89], w_hssi_10g_rx_pcs_rx_data[88], w_hssi_10g_rx_pcs_rx_data[87], w_hssi_10g_rx_pcs_rx_data[86], w_hssi_10g_rx_pcs_rx_data[85], w_hssi_10g_rx_pcs_rx_data[84], w_hssi_10g_rx_pcs_rx_data[83], w_hssi_10g_rx_pcs_rx_data[82], w_hssi_10g_rx_pcs_rx_data[81], w_hssi_10g_rx_pcs_rx_data[80], w_hssi_10g_rx_pcs_rx_data[79], w_hssi_10g_rx_pcs_rx_data[78], w_hssi_10g_rx_pcs_rx_data[77], w_hssi_10g_rx_pcs_rx_data[76], w_hssi_10g_rx_pcs_rx_data[75], w_hssi_10g_rx_pcs_rx_data[74], w_hssi_10g_rx_pcs_rx_data[73], w_hssi_10g_rx_pcs_rx_data[72], w_hssi_10g_rx_pcs_rx_data[71], w_hssi_10g_rx_pcs_rx_data[70], w_hssi_10g_rx_pcs_rx_data[69], w_hssi_10g_rx_pcs_rx_data[68], w_hssi_10g_rx_pcs_rx_data[67], w_hssi_10g_rx_pcs_rx_data[66], w_hssi_10g_rx_pcs_rx_data[65], w_hssi_10g_rx_pcs_rx_data[64], w_hssi_10g_rx_pcs_rx_data[63], w_hssi_10g_rx_pcs_rx_data[62], w_hssi_10g_rx_pcs_rx_data[61], w_hssi_10g_rx_pcs_rx_data[60], w_hssi_10g_rx_pcs_rx_data[59], w_hssi_10g_rx_pcs_rx_data[58], w_hssi_10g_rx_pcs_rx_data[57], w_hssi_10g_rx_pcs_rx_data[56], w_hssi_10g_rx_pcs_rx_data[55], w_hssi_10g_rx_pcs_rx_data[54], w_hssi_10g_rx_pcs_rx_data[53], w_hssi_10g_rx_pcs_rx_data[52], w_hssi_10g_rx_pcs_rx_data[51], w_hssi_10g_rx_pcs_rx_data[50], w_hssi_10g_rx_pcs_rx_data[49], w_hssi_10g_rx_pcs_rx_data[48], w_hssi_10g_rx_pcs_rx_data[47], w_hssi_10g_rx_pcs_rx_data[46], w_hssi_10g_rx_pcs_rx_data[45], w_hssi_10g_rx_pcs_rx_data[44], w_hssi_10g_rx_pcs_rx_data[43], w_hssi_10g_rx_pcs_rx_data[42], w_hssi_10g_rx_pcs_rx_data[41], w_hssi_10g_rx_pcs_rx_data[40], w_hssi_10g_rx_pcs_rx_data[39], w_hssi_10g_rx_pcs_rx_data[38], w_hssi_10g_rx_pcs_rx_data[37], w_hssi_10g_rx_pcs_rx_data[36], w_hssi_10g_rx_pcs_rx_data[35], w_hssi_10g_rx_pcs_rx_data[34], w_hssi_10g_rx_pcs_rx_data[33], w_hssi_10g_rx_pcs_rx_data[32], w_hssi_10g_rx_pcs_rx_data[31], w_hssi_10g_rx_pcs_rx_data[30], w_hssi_10g_rx_pcs_rx_data[29], w_hssi_10g_rx_pcs_rx_data[28], w_hssi_10g_rx_pcs_rx_data[27], w_hssi_10g_rx_pcs_rx_data[26], w_hssi_10g_rx_pcs_rx_data[25], w_hssi_10g_rx_pcs_rx_data[24], w_hssi_10g_rx_pcs_rx_data[23], w_hssi_10g_rx_pcs_rx_data[22], w_hssi_10g_rx_pcs_rx_data[21], w_hssi_10g_rx_pcs_rx_data[20], w_hssi_10g_rx_pcs_rx_data[19], w_hssi_10g_rx_pcs_rx_data[18], w_hssi_10g_rx_pcs_rx_data[17], w_hssi_10g_rx_pcs_rx_data[16], w_hssi_10g_rx_pcs_rx_data[15], w_hssi_10g_rx_pcs_rx_data[14], w_hssi_10g_rx_pcs_rx_data[13], w_hssi_10g_rx_pcs_rx_data[12], w_hssi_10g_rx_pcs_rx_data[11], w_hssi_10g_rx_pcs_rx_data[10], w_hssi_10g_rx_pcs_rx_data[9], w_hssi_10g_rx_pcs_rx_data[8], w_hssi_10g_rx_pcs_rx_data[7], w_hssi_10g_rx_pcs_rx_data[6], w_hssi_10g_rx_pcs_rx_data[5], w_hssi_10g_rx_pcs_rx_data[4], w_hssi_10g_rx_pcs_rx_data[3], w_hssi_10g_rx_pcs_rx_data[2], w_hssi_10g_rx_pcs_rx_data[1], w_hssi_10g_rx_pcs_rx_data[0]}),
				.int_pldif_10g_rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.int_pldif_10g_rx_diag_status({w_hssi_10g_rx_pcs_rx_diag_status[1], w_hssi_10g_rx_pcs_rx_diag_status[0]}),
				.int_pldif_10g_rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.int_pldif_10g_rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.int_pldif_10g_rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.int_pldif_10g_rx_fifo_num({w_hssi_10g_rx_pcs_rx_fifo_num[4], w_hssi_10g_rx_pcs_rx_fifo_num[3], w_hssi_10g_rx_pcs_rx_fifo_num[2], w_hssi_10g_rx_pcs_rx_fifo_num[1], w_hssi_10g_rx_pcs_rx_fifo_num[0]}),
				.int_pldif_10g_rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.int_pldif_10g_rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.int_pldif_10g_rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.int_pldif_10g_rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.int_pldif_10g_rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.int_pldif_10g_rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				.int_pldif_8g_a1a2_k1k2_flag({w_hssi_8g_rx_pcs_a1a2k1k2flag[3], w_hssi_8g_rx_pcs_a1a2k1k2flag[2], w_hssi_8g_rx_pcs_a1a2k1k2flag[1], w_hssi_8g_rx_pcs_a1a2k1k2flag[0]}),
				.int_pldif_8g_empty_rmf(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.int_pldif_8g_empty_rx(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.int_pldif_8g_full_rmf(w_hssi_8g_rx_pcs_rm_fifo_full),
				.int_pldif_8g_full_rx(w_hssi_8g_rx_pcs_pcfifofull),
				.int_pldif_8g_phystatus(w_hssi_8g_rx_pcs_phystatus),
				.int_pldif_8g_rx_blk_start({w_hssi_8g_rx_pcs_rx_blk_start[3], w_hssi_8g_rx_pcs_rx_blk_start[2], w_hssi_8g_rx_pcs_rx_blk_start[1], w_hssi_8g_rx_pcs_rx_blk_start[0]}),
				.int_pldif_8g_rx_clk(w_hssi_8g_rx_pcs_clock_to_pld),
				.int_pldif_8g_rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_8g_rx_data_valid({w_hssi_8g_rx_pcs_rx_data_valid[3], w_hssi_8g_rx_pcs_rx_data_valid[2], w_hssi_8g_rx_pcs_rx_data_valid[1], w_hssi_8g_rx_pcs_rx_data_valid[0]}),
				.int_pldif_8g_rx_rstn_sync2wrfifo(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.int_pldif_8g_rx_sync_hdr({w_hssi_8g_rx_pcs_rx_sync_hdr[1], w_hssi_8g_rx_pcs_rx_sync_hdr[0]}),
				.int_pldif_8g_rxd({w_hssi_8g_rx_pcs_dataout[63], w_hssi_8g_rx_pcs_dataout[62], w_hssi_8g_rx_pcs_dataout[61], w_hssi_8g_rx_pcs_dataout[60], w_hssi_8g_rx_pcs_dataout[59], w_hssi_8g_rx_pcs_dataout[58], w_hssi_8g_rx_pcs_dataout[57], w_hssi_8g_rx_pcs_dataout[56], w_hssi_8g_rx_pcs_dataout[55], w_hssi_8g_rx_pcs_dataout[54], w_hssi_8g_rx_pcs_dataout[53], w_hssi_8g_rx_pcs_dataout[52], w_hssi_8g_rx_pcs_dataout[51], w_hssi_8g_rx_pcs_dataout[50], w_hssi_8g_rx_pcs_dataout[49], w_hssi_8g_rx_pcs_dataout[48], w_hssi_8g_rx_pcs_dataout[47], w_hssi_8g_rx_pcs_dataout[46], w_hssi_8g_rx_pcs_dataout[45], w_hssi_8g_rx_pcs_dataout[44], w_hssi_8g_rx_pcs_dataout[43], w_hssi_8g_rx_pcs_dataout[42], w_hssi_8g_rx_pcs_dataout[41], w_hssi_8g_rx_pcs_dataout[40], w_hssi_8g_rx_pcs_dataout[39], w_hssi_8g_rx_pcs_dataout[38], w_hssi_8g_rx_pcs_dataout[37], w_hssi_8g_rx_pcs_dataout[36], w_hssi_8g_rx_pcs_dataout[35], w_hssi_8g_rx_pcs_dataout[34], w_hssi_8g_rx_pcs_dataout[33], w_hssi_8g_rx_pcs_dataout[32], w_hssi_8g_rx_pcs_dataout[31], w_hssi_8g_rx_pcs_dataout[30], w_hssi_8g_rx_pcs_dataout[29], w_hssi_8g_rx_pcs_dataout[28], w_hssi_8g_rx_pcs_dataout[27], w_hssi_8g_rx_pcs_dataout[26], w_hssi_8g_rx_pcs_dataout[25], w_hssi_8g_rx_pcs_dataout[24], w_hssi_8g_rx_pcs_dataout[23], w_hssi_8g_rx_pcs_dataout[22], w_hssi_8g_rx_pcs_dataout[21], w_hssi_8g_rx_pcs_dataout[20], w_hssi_8g_rx_pcs_dataout[19], w_hssi_8g_rx_pcs_dataout[18], w_hssi_8g_rx_pcs_dataout[17], w_hssi_8g_rx_pcs_dataout[16], w_hssi_8g_rx_pcs_dataout[15], w_hssi_8g_rx_pcs_dataout[14], w_hssi_8g_rx_pcs_dataout[13], w_hssi_8g_rx_pcs_dataout[12], w_hssi_8g_rx_pcs_dataout[11], w_hssi_8g_rx_pcs_dataout[10], w_hssi_8g_rx_pcs_dataout[9], w_hssi_8g_rx_pcs_dataout[8], w_hssi_8g_rx_pcs_dataout[7], w_hssi_8g_rx_pcs_dataout[6], w_hssi_8g_rx_pcs_dataout[5], w_hssi_8g_rx_pcs_dataout[4], w_hssi_8g_rx_pcs_dataout[3], w_hssi_8g_rx_pcs_dataout[2], w_hssi_8g_rx_pcs_dataout[1], w_hssi_8g_rx_pcs_dataout[0]}),
				.int_pldif_8g_rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.int_pldif_8g_rxstatus({w_hssi_8g_rx_pcs_rxstatus[2], w_hssi_8g_rx_pcs_rxstatus[1], w_hssi_8g_rx_pcs_rxstatus[0]}),
				.int_pldif_8g_rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.int_pldif_8g_signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.int_pldif_8g_wa_boundary({w_hssi_8g_rx_pcs_word_align_boundary[4], w_hssi_8g_rx_pcs_word_align_boundary[3], w_hssi_8g_rx_pcs_word_align_boundary[2], w_hssi_8g_rx_pcs_word_align_boundary[1], w_hssi_8g_rx_pcs_word_align_boundary[0]}),
				.int_pldif_krfec_rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.int_pldif_krfec_rx_data_status({w_hssi_krfec_rx_pcs_rx_data_status[1], w_hssi_krfec_rx_pcs_rx_data_status[0]}),
				.int_pldif_krfec_rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.int_pldif_pmaif_clkdiv_rx(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pldif_pmaif_clkdiv_rx_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pldif_pmaif_rx_data({w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0]}),
				.int_pldif_pmaif_rx_prbs_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pldif_pmaif_rx_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.pld_10g_krfec_rx_clr_errblk_cnt(in_pld_10g_krfec_rx_clr_errblk_cnt),
				.pld_10g_krfec_rx_pld_rst_n(in_pld_10g_krfec_rx_pld_rst_n),
				.pld_10g_rx_align_clr(in_pld_10g_rx_align_clr),
				.pld_10g_rx_clr_ber_count(in_pld_10g_rx_clr_ber_count),
				.pld_10g_rx_rd_en(in_pld_10g_rx_rd_en),
				.pld_8g_a1a2_size(in_pld_8g_a1a2_size),
				.pld_8g_bitloc_rev_en(in_pld_8g_bitloc_rev_en),
				.pld_8g_byte_rev_en(in_pld_8g_byte_rev_en),
				.pld_8g_encdt(in_pld_8g_encdt),
				.pld_8g_g3_rx_pld_rst_n(in_pld_8g_g3_rx_pld_rst_n),
				.pld_8g_rdenable_rx(in_pld_8g_rdenable_rx),
				.pld_8g_rxpolarity(in_pld_8g_rxpolarity),
				.pld_8g_wrdisable_rx(in_pld_8g_wrdisable_rx),
				.pld_bitslip(in_pld_bitslip),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_rxpma_rstb(in_pld_pma_rxpma_rstb),
				.pld_pmaif_rx_pld_rst_n(in_pld_pmaif_rx_pld_rst_n),
				.pld_pmaif_rxclkslip(in_pld_pmaif_rxclkslip),
				.pld_polinv_rx(in_pld_polinv_rx),
				.pld_rx_clk(in_pld_rx_clk),
				.pld_rx_prbs_err_clr(in_pld_rx_prbs_err_clr),
				.pld_syncsm_en(in_pld_syncsm_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.int_pldif_pmaif_rx_pld_clk(),
				.pld_8g_wa_boundary_txclk_fastreg(),
				.pld_8g_wa_boundary_txclk_reg(),
				.pld_bitslip_10g_txclk_reg(),
				.pld_bitslip_8g_txclk_reg(),
				.pld_bitslip_rxclk_parallel_loopback_reg(),
				.pld_bitslip_rxclk_reg(),
				.pld_pcs_rx_clk_out_pcsdirect_wire(),
				.pld_pma_rx_clk_out_10g_or_pcsdirect_wire(),
				.pld_pma_rx_clk_out_8g_wire(),
				.pld_pmaif_rx_pld_rst_n_reg(),
				.pld_pmaif_tx_pld_rst_n_txclk_reg(),
				.pld_polinv_rx_reg(),
				.pld_rx_clk_fifo(),
				.pld_rx_control_fifo(),
				.pld_rx_control_pcsdirect_reg(),
				.pld_rx_data_fifo(),
				.pld_rx_data_pcsdirect_reg(),
				.pld_rx_prbs_done_reg(),
				.pld_rx_prbs_done_txclk_reg(),
				.pld_rx_prbs_err_clr_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_clr_reg(),
				.pld_rx_prbs_err_disprbs_reg(),
				.pld_rx_prbs_err_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_reg(),
				.pma_rx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_data[50:0] = 51'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3:0] = 4'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_control[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_data[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pcs_pma_interface
			twentynm_hssi_tx_pcs_pma_interface #(
				.bypass_pma_txelecidle(hssi_tx_pcs_pma_interface_bypass_pma_txelecidle),
				.channel_operation_mode(hssi_tx_pcs_pma_interface_channel_operation_mode),
				.lpbk_en(hssi_tx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_tx_pcs_pma_interface_master_clk_sel),
				.pcie_sub_prot_mode_tx(hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx),
				.pldif_datawidth_mode(hssi_tx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_tx(hssi_tx_pcs_pma_interface_pma_dw_tx),
				.pma_if_dft_en(hssi_tx_pcs_pma_interface_pma_if_dft_en),
				.pmagate_en(hssi_tx_pcs_pma_interface_pmagate_en),
				.prbs9_dwidth(hssi_tx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_tx_pcs_pma_interface_prbs_clken),
				.prbs_gen_pat(hssi_tx_pcs_pma_interface_prbs_gen_pat),
				.prot_mode_tx(hssi_tx_pcs_pma_interface_prot_mode_tx),
				.reconfig_settings(hssi_tx_pcs_pma_interface_reconfig_settings),
				.silicon_rev( "20nm3" ),       //PARAM_HIDE
				.sq_wave_num(hssi_tx_pcs_pma_interface_sq_wave_num),
				.sqwgen_clken(hssi_tx_pcs_pma_interface_sqwgen_clken),
				.sup_mode(hssi_tx_pcs_pma_interface_sup_mode),
				.tx_dyn_polarity_inversion(hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion),
				.tx_pma_data_sel(hssi_tx_pcs_pma_interface_tx_pma_data_sel),
				.tx_static_polarity_inversion(hssi_tx_pcs_pma_interface_tx_static_polarity_inversion),
				.uhsif_cnt_step_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock),
				.uhsif_cnt_thresh_filt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value),
				.uhsif_cnt_thresh_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock),
				.uhsif_dcn_test_update_period(hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period),
				.uhsif_dcn_testmode_enable(hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable),
				.uhsif_dead_zone_count_thresh(hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh),
				.uhsif_dead_zone_detection_enable(hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable),
				.uhsif_dead_zone_obser_window(hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window),
				.uhsif_dead_zone_skip_size(hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size),
				.uhsif_delay_cell_index_sel(hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel),
				.uhsif_delay_cell_margin(hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin),
				.uhsif_delay_cell_static_index_value(hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value),
				.uhsif_dft_dead_zone_control(hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control),
				.uhsif_dft_up_filt_control(hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control),
				.uhsif_enable(hssi_tx_pcs_pma_interface_uhsif_enable),
				.uhsif_lock_det_segsz_after_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock),
				.uhsif_lock_det_segsz_before_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock),
				.uhsif_lock_det_thresh_cnt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value),
				.uhsif_lock_det_thresh_cnt_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value),
				.uhsif_lock_det_thresh_diff_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value),
				.uhsif_lock_det_thresh_diff_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value)
			) inst_twentynm_hssi_tx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.int_pmaif_8g_txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.int_pmaif_pldif_tx_clkdiv(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pmaif_pldif_tx_clkdiv_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pmaif_pldif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.int_pmaif_pldif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.int_tx_dft_obsrv_clk(w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk),
				.pma_tx_elec_idle(w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle),
				.pma_tx_pma_data(w_hssi_tx_pcs_pma_interface_pma_tx_pma_data),
				.pma_txpma_rstb(w_hssi_tx_pcs_pma_interface_pma_txpma_rstb),
				.tx_pma_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback),
				.tx_pma_uhsif_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback),
				.tx_prbs_gen_test(w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test),
				.uhsif_test_out_1(w_hssi_tx_pcs_pma_interface_uhsif_test_out_1),
				.uhsif_test_out_2(w_hssi_tx_pcs_pma_interface_uhsif_test_out_2),
				.uhsif_test_out_3(w_hssi_tx_pcs_pma_interface_uhsif_test_out_3),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.int_pmaif_10g_tx_pma_data({w_hssi_10g_tx_pcs_tx_pma_data[63], w_hssi_10g_tx_pcs_tx_pma_data[62], w_hssi_10g_tx_pcs_tx_pma_data[61], w_hssi_10g_tx_pcs_tx_pma_data[60], w_hssi_10g_tx_pcs_tx_pma_data[59], w_hssi_10g_tx_pcs_tx_pma_data[58], w_hssi_10g_tx_pcs_tx_pma_data[57], w_hssi_10g_tx_pcs_tx_pma_data[56], w_hssi_10g_tx_pcs_tx_pma_data[55], w_hssi_10g_tx_pcs_tx_pma_data[54], w_hssi_10g_tx_pcs_tx_pma_data[53], w_hssi_10g_tx_pcs_tx_pma_data[52], w_hssi_10g_tx_pcs_tx_pma_data[51], w_hssi_10g_tx_pcs_tx_pma_data[50], w_hssi_10g_tx_pcs_tx_pma_data[49], w_hssi_10g_tx_pcs_tx_pma_data[48], w_hssi_10g_tx_pcs_tx_pma_data[47], w_hssi_10g_tx_pcs_tx_pma_data[46], w_hssi_10g_tx_pcs_tx_pma_data[45], w_hssi_10g_tx_pcs_tx_pma_data[44], w_hssi_10g_tx_pcs_tx_pma_data[43], w_hssi_10g_tx_pcs_tx_pma_data[42], w_hssi_10g_tx_pcs_tx_pma_data[41], w_hssi_10g_tx_pcs_tx_pma_data[40], w_hssi_10g_tx_pcs_tx_pma_data[39], w_hssi_10g_tx_pcs_tx_pma_data[38], w_hssi_10g_tx_pcs_tx_pma_data[37], w_hssi_10g_tx_pcs_tx_pma_data[36], w_hssi_10g_tx_pcs_tx_pma_data[35], w_hssi_10g_tx_pcs_tx_pma_data[34], w_hssi_10g_tx_pcs_tx_pma_data[33], w_hssi_10g_tx_pcs_tx_pma_data[32], w_hssi_10g_tx_pcs_tx_pma_data[31], w_hssi_10g_tx_pcs_tx_pma_data[30], w_hssi_10g_tx_pcs_tx_pma_data[29], w_hssi_10g_tx_pcs_tx_pma_data[28], w_hssi_10g_tx_pcs_tx_pma_data[27], w_hssi_10g_tx_pcs_tx_pma_data[26], w_hssi_10g_tx_pcs_tx_pma_data[25], w_hssi_10g_tx_pcs_tx_pma_data[24], w_hssi_10g_tx_pcs_tx_pma_data[23], w_hssi_10g_tx_pcs_tx_pma_data[22], w_hssi_10g_tx_pcs_tx_pma_data[21], w_hssi_10g_tx_pcs_tx_pma_data[20], w_hssi_10g_tx_pcs_tx_pma_data[19], w_hssi_10g_tx_pcs_tx_pma_data[18], w_hssi_10g_tx_pcs_tx_pma_data[17], w_hssi_10g_tx_pcs_tx_pma_data[16], w_hssi_10g_tx_pcs_tx_pma_data[15], w_hssi_10g_tx_pcs_tx_pma_data[14], w_hssi_10g_tx_pcs_tx_pma_data[13], w_hssi_10g_tx_pcs_tx_pma_data[12], w_hssi_10g_tx_pcs_tx_pma_data[11], w_hssi_10g_tx_pcs_tx_pma_data[10], w_hssi_10g_tx_pcs_tx_pma_data[9], w_hssi_10g_tx_pcs_tx_pma_data[8], w_hssi_10g_tx_pcs_tx_pma_data[7], w_hssi_10g_tx_pcs_tx_pma_data[6], w_hssi_10g_tx_pcs_tx_pma_data[5], w_hssi_10g_tx_pcs_tx_pma_data[4], w_hssi_10g_tx_pcs_tx_pma_data[3], w_hssi_10g_tx_pcs_tx_pma_data[2], w_hssi_10g_tx_pcs_tx_pma_data[1], w_hssi_10g_tx_pcs_tx_pma_data[0]}),
				.int_pmaif_10g_tx_pma_data_gate_val({w_hssi_10g_tx_pcs_tx_pma_gating_val[63], w_hssi_10g_tx_pcs_tx_pma_gating_val[62], w_hssi_10g_tx_pcs_tx_pma_gating_val[61], w_hssi_10g_tx_pcs_tx_pma_gating_val[60], w_hssi_10g_tx_pcs_tx_pma_gating_val[59], w_hssi_10g_tx_pcs_tx_pma_gating_val[58], w_hssi_10g_tx_pcs_tx_pma_gating_val[57], w_hssi_10g_tx_pcs_tx_pma_gating_val[56], w_hssi_10g_tx_pcs_tx_pma_gating_val[55], w_hssi_10g_tx_pcs_tx_pma_gating_val[54], w_hssi_10g_tx_pcs_tx_pma_gating_val[53], w_hssi_10g_tx_pcs_tx_pma_gating_val[52], w_hssi_10g_tx_pcs_tx_pma_gating_val[51], w_hssi_10g_tx_pcs_tx_pma_gating_val[50], w_hssi_10g_tx_pcs_tx_pma_gating_val[49], w_hssi_10g_tx_pcs_tx_pma_gating_val[48], w_hssi_10g_tx_pcs_tx_pma_gating_val[47], w_hssi_10g_tx_pcs_tx_pma_gating_val[46], w_hssi_10g_tx_pcs_tx_pma_gating_val[45], w_hssi_10g_tx_pcs_tx_pma_gating_val[44], w_hssi_10g_tx_pcs_tx_pma_gating_val[43], w_hssi_10g_tx_pcs_tx_pma_gating_val[42], w_hssi_10g_tx_pcs_tx_pma_gating_val[41], w_hssi_10g_tx_pcs_tx_pma_gating_val[40], w_hssi_10g_tx_pcs_tx_pma_gating_val[39], w_hssi_10g_tx_pcs_tx_pma_gating_val[38], w_hssi_10g_tx_pcs_tx_pma_gating_val[37], w_hssi_10g_tx_pcs_tx_pma_gating_val[36], w_hssi_10g_tx_pcs_tx_pma_gating_val[35], w_hssi_10g_tx_pcs_tx_pma_gating_val[34], w_hssi_10g_tx_pcs_tx_pma_gating_val[33], w_hssi_10g_tx_pcs_tx_pma_gating_val[32], w_hssi_10g_tx_pcs_tx_pma_gating_val[31], w_hssi_10g_tx_pcs_tx_pma_gating_val[30], w_hssi_10g_tx_pcs_tx_pma_gating_val[29], w_hssi_10g_tx_pcs_tx_pma_gating_val[28], w_hssi_10g_tx_pcs_tx_pma_gating_val[27], w_hssi_10g_tx_pcs_tx_pma_gating_val[26], w_hssi_10g_tx_pcs_tx_pma_gating_val[25], w_hssi_10g_tx_pcs_tx_pma_gating_val[24], w_hssi_10g_tx_pcs_tx_pma_gating_val[23], w_hssi_10g_tx_pcs_tx_pma_gating_val[22], w_hssi_10g_tx_pcs_tx_pma_gating_val[21], w_hssi_10g_tx_pcs_tx_pma_gating_val[20], w_hssi_10g_tx_pcs_tx_pma_gating_val[19], w_hssi_10g_tx_pcs_tx_pma_gating_val[18], w_hssi_10g_tx_pcs_tx_pma_gating_val[17], w_hssi_10g_tx_pcs_tx_pma_gating_val[16], w_hssi_10g_tx_pcs_tx_pma_gating_val[15], w_hssi_10g_tx_pcs_tx_pma_gating_val[14], w_hssi_10g_tx_pcs_tx_pma_gating_val[13], w_hssi_10g_tx_pcs_tx_pma_gating_val[12], w_hssi_10g_tx_pcs_tx_pma_gating_val[11], w_hssi_10g_tx_pcs_tx_pma_gating_val[10], w_hssi_10g_tx_pcs_tx_pma_gating_val[9], w_hssi_10g_tx_pcs_tx_pma_gating_val[8], w_hssi_10g_tx_pcs_tx_pma_gating_val[7], w_hssi_10g_tx_pcs_tx_pma_gating_val[6], w_hssi_10g_tx_pcs_tx_pma_gating_val[5], w_hssi_10g_tx_pcs_tx_pma_gating_val[4], w_hssi_10g_tx_pcs_tx_pma_gating_val[3], w_hssi_10g_tx_pcs_tx_pma_gating_val[2], w_hssi_10g_tx_pcs_tx_pma_gating_val[1], w_hssi_10g_tx_pcs_tx_pma_gating_val[0]}),
				.int_pmaif_8g_pudr({w_hssi_8g_tx_pcs_dataout[19], w_hssi_8g_tx_pcs_dataout[18], w_hssi_8g_tx_pcs_dataout[17], w_hssi_8g_tx_pcs_dataout[16], w_hssi_8g_tx_pcs_dataout[15], w_hssi_8g_tx_pcs_dataout[14], w_hssi_8g_tx_pcs_dataout[13], w_hssi_8g_tx_pcs_dataout[12], w_hssi_8g_tx_pcs_dataout[11], w_hssi_8g_tx_pcs_dataout[10], w_hssi_8g_tx_pcs_dataout[9], w_hssi_8g_tx_pcs_dataout[8], w_hssi_8g_tx_pcs_dataout[7], w_hssi_8g_tx_pcs_dataout[6], w_hssi_8g_tx_pcs_dataout[5], w_hssi_8g_tx_pcs_dataout[4], w_hssi_8g_tx_pcs_dataout[3], w_hssi_8g_tx_pcs_dataout[2], w_hssi_8g_tx_pcs_dataout[1], w_hssi_8g_tx_pcs_dataout[0]}),
				.int_pmaif_8g_tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.int_pmaif_8g_tx_elec_idle(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_pma_data_out({w_hssi_gen3_tx_pcs_data_out[31], w_hssi_gen3_tx_pcs_data_out[30], w_hssi_gen3_tx_pcs_data_out[29], w_hssi_gen3_tx_pcs_data_out[28], w_hssi_gen3_tx_pcs_data_out[27], w_hssi_gen3_tx_pcs_data_out[26], w_hssi_gen3_tx_pcs_data_out[25], w_hssi_gen3_tx_pcs_data_out[24], w_hssi_gen3_tx_pcs_data_out[23], w_hssi_gen3_tx_pcs_data_out[22], w_hssi_gen3_tx_pcs_data_out[21], w_hssi_gen3_tx_pcs_data_out[20], w_hssi_gen3_tx_pcs_data_out[19], w_hssi_gen3_tx_pcs_data_out[18], w_hssi_gen3_tx_pcs_data_out[17], w_hssi_gen3_tx_pcs_data_out[16], w_hssi_gen3_tx_pcs_data_out[15], w_hssi_gen3_tx_pcs_data_out[14], w_hssi_gen3_tx_pcs_data_out[13], w_hssi_gen3_tx_pcs_data_out[12], w_hssi_gen3_tx_pcs_data_out[11], w_hssi_gen3_tx_pcs_data_out[10], w_hssi_gen3_tx_pcs_data_out[9], w_hssi_gen3_tx_pcs_data_out[8], w_hssi_gen3_tx_pcs_data_out[7], w_hssi_gen3_tx_pcs_data_out[6], w_hssi_gen3_tx_pcs_data_out[5], w_hssi_gen3_tx_pcs_data_out[4], w_hssi_gen3_tx_pcs_data_out[3], w_hssi_gen3_tx_pcs_data_out[2], w_hssi_gen3_tx_pcs_data_out[1], w_hssi_gen3_tx_pcs_data_out[0]}),
				.int_pmaif_g3_pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.int_pmaif_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pmaif_pldif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pmaif_pldif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0]}),
				.int_pmaif_pldif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pmaif_pldif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.int_pmaif_pldif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pmaif_pldif_uhsif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0]}),
				.pma_tx_clkdiv_user(in_pma_tx_clkdiv_user),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.refclk_dig_uhsif(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.uhsif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.uhsif_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				
				// UNUSED
				.avmm_user_dataout(),
				.write_en(),
				.write_en_ack()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4:0] = 5'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_txpma_rstb = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pld_pcs_interface
			twentynm_hssi_tx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx),
				.hd_10g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx),
				.hd_10g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx),
				.hd_10g_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx),
				.hd_10g_lpbk_en(hssi_tx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx),
				.hd_10g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx),
				.hd_10g_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx),
				.hd_8g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx),
				.hd_8g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx),
				.hd_8g_hip_mode(hssi_tx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_tx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx),
				.hd_8g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx),
				.hd_chnl_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx),
				.hd_chnl_frequency_rules_en(hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_tx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_tx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx),
				.hd_chnl_lpbk_en(hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx),
				.hd_chnl_pld_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz),
				.hd_chnl_pld_uhsif_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz),
				.hd_chnl_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx),
				.hd_chnl_pma_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz),
				.hd_chnl_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx),
				.hd_chnl_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx),
				.hd_fifo_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx),
				.hd_fifo_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx),
				.hd_g3_prot_mode(hssi_tx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx),
				.hd_krfec_lpbk_en(hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx),
				.hd_pldif_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx),
				.hd_pmaif_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_ctrl_plane_bonding(hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding),
				.hd_pmaif_lpbk_en(hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx),
				.hd_pmaif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx),
				.hd_pmaif_sim_mode(hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_tx_clk_out_sel(hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel),
				.pcs_tx_clk_source(hssi_tx_pld_pcs_interface_pcs_tx_clk_source),
				.pcs_tx_data_source(hssi_tx_pld_pcs_interface_pcs_tx_data_source),
				.pcs_tx_delay1_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en),
				.pcs_tx_delay1_clk_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel),
				.pcs_tx_delay1_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl),
				.pcs_tx_delay1_data_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel),
				.pcs_tx_delay2_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en),
				.pcs_tx_delay2_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl),
				.pcs_tx_output_sel(hssi_tx_pld_pcs_interface_pcs_tx_output_sel),
				.reconfig_settings(hssi_tx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm3" )       //PARAM_HIDE
			) inst_twentynm_hssi_tx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pld_pcs_interface_blockselect),
				.hip_tx_clk(w_hssi_tx_pld_pcs_interface_hip_tx_clk),
				.int_pldif_10g_tx_bitslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip),
				.int_pldif_10g_tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.int_pldif_10g_tx_control(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control),
				.int_pldif_10g_tx_control_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg),
				.int_pldif_10g_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data),
				.int_pldif_10g_tx_data_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg),
				.int_pldif_10g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.int_pldif_10g_tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.int_pldif_10g_tx_diag_status(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status),
				.int_pldif_10g_tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.int_pldif_10g_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.int_pldif_10g_tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				.int_pldif_8g_pld_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.int_pldif_8g_powerdown(w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown),
				.int_pldif_8g_rddisable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.int_pldif_8g_rev_loopbk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.int_pldif_8g_tx_blk_start(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start),
				.int_pldif_8g_tx_boundary_sel(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel),
				.int_pldif_8g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid),
				.int_pldif_8g_tx_sync_hdr(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr),
				.int_pldif_8g_txd(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd),
				.int_pldif_8g_txd_fast_reg(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg),
				.int_pldif_8g_txdeemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.int_pldif_8g_txdetectrxloopback(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.int_pldif_8g_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.int_pldif_8g_txmargin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin),
				.int_pldif_8g_txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.int_pldif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.int_pldif_8g_wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				.int_pldif_pmaif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pldif_pmaif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pldif_pmaif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data),
				.int_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pldif_pmaif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pldif_pmaif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pldif_pmaif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pldif_pmaif_uhsif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data),
				.pld_10g_krfec_tx_frame(w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame),
				.pld_10g_tx_burst_en_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe),
				.pld_10g_tx_empty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty),
				.pld_10g_tx_fifo_num(w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num),
				.pld_10g_tx_full(w_hssi_tx_pld_pcs_interface_pld_10g_tx_full),
				.pld_10g_tx_pempty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty),
				.pld_10g_tx_pfull(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull),
				.pld_10g_tx_wordslip_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe),
				.pld_8g_empty_tx(w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx),
				.pld_8g_full_tx(w_hssi_tx_pld_pcs_interface_pld_8g_full_tx),
				.pld_krfec_tx_alignment(w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment),
				.pld_pcs_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out),
				.pld_pma_clkdiv_tx_user(w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user),
				.pld_pma_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out),
				.pld_uhsif_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.hip_tx_data({in_hip_tx_data[63], in_hip_tx_data[62], in_hip_tx_data[61], in_hip_tx_data[60], in_hip_tx_data[59], in_hip_tx_data[58], in_hip_tx_data[57], in_hip_tx_data[56], in_hip_tx_data[55], in_hip_tx_data[54], in_hip_tx_data[53], in_hip_tx_data[52], in_hip_tx_data[51], in_hip_tx_data[50], in_hip_tx_data[49], in_hip_tx_data[48], in_hip_tx_data[47], in_hip_tx_data[46], in_hip_tx_data[45], in_hip_tx_data[44], in_hip_tx_data[43], in_hip_tx_data[42], in_hip_tx_data[41], in_hip_tx_data[40], in_hip_tx_data[39], in_hip_tx_data[38], in_hip_tx_data[37], in_hip_tx_data[36], in_hip_tx_data[35], in_hip_tx_data[34], in_hip_tx_data[33], in_hip_tx_data[32], in_hip_tx_data[31], in_hip_tx_data[30], in_hip_tx_data[29], in_hip_tx_data[28], in_hip_tx_data[27], in_hip_tx_data[26], in_hip_tx_data[25], in_hip_tx_data[24], in_hip_tx_data[23], in_hip_tx_data[22], in_hip_tx_data[21], in_hip_tx_data[20], in_hip_tx_data[19], in_hip_tx_data[18], in_hip_tx_data[17], in_hip_tx_data[16], in_hip_tx_data[15], in_hip_tx_data[14], in_hip_tx_data[13], in_hip_tx_data[12], in_hip_tx_data[11], in_hip_tx_data[10], in_hip_tx_data[9], in_hip_tx_data[8], in_hip_tx_data[7], in_hip_tx_data[6], in_hip_tx_data[5], in_hip_tx_data[4], in_hip_tx_data[3], in_hip_tx_data[2], in_hip_tx_data[1], in_hip_tx_data[0]}),
				.int_pldif_10g_tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.int_pldif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.int_pldif_10g_tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_10g_tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.int_pldif_10g_tx_fifo_num({w_hssi_10g_tx_pcs_tx_fifo_num[3], w_hssi_10g_tx_pcs_tx_fifo_num[2], w_hssi_10g_tx_pcs_tx_fifo_num[1], w_hssi_10g_tx_pcs_tx_fifo_num[0]}),
				.int_pldif_10g_tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.int_pldif_10g_tx_full(w_hssi_10g_tx_pcs_tx_full),
				.int_pldif_10g_tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.int_pldif_10g_tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.int_pldif_10g_tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				.int_pldif_8g_empty_tx(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.int_pldif_8g_full_tx(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.int_pldif_8g_tx_clk_out(w_hssi_8g_tx_pcs_clk_out),
				.int_pldif_8g_tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_krfec_tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.int_pldif_krfec_tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.int_pldif_pmaif_clkdiv_tx(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pldif_pmaif_clkdiv_tx_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pldif_pmaif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.pld_10g_krfec_tx_pld_rst_n(in_pld_10g_krfec_tx_pld_rst_n),
				.pld_10g_tx_bitslip({in_pld_10g_tx_bitslip[6], in_pld_10g_tx_bitslip[5], in_pld_10g_tx_bitslip[4], in_pld_10g_tx_bitslip[3], in_pld_10g_tx_bitslip[2], in_pld_10g_tx_bitslip[1], in_pld_10g_tx_bitslip[0]}),
				.pld_10g_tx_burst_en(in_pld_10g_tx_burst_en),
				.pld_10g_tx_data_valid(in_pld_10g_tx_data_valid),
				.pld_10g_tx_diag_status({in_pld_10g_tx_diag_status[1], in_pld_10g_tx_diag_status[0]}),
				.pld_10g_tx_wordslip(in_pld_10g_tx_wordslip),
				.pld_8g_g3_tx_pld_rst_n(in_pld_8g_g3_tx_pld_rst_n),
				.pld_8g_rddisable_tx(in_pld_8g_rddisable_tx),
				.pld_8g_tx_boundary_sel({in_pld_8g_tx_boundary_sel[4], in_pld_8g_tx_boundary_sel[3], in_pld_8g_tx_boundary_sel[2], in_pld_8g_tx_boundary_sel[1], in_pld_8g_tx_boundary_sel[0]}),
				.pld_8g_wrenable_tx(in_pld_8g_wrenable_tx),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_txpma_rstb(in_pld_pma_txpma_rstb),
				.pld_pmaif_tx_pld_rst_n(in_pld_pmaif_tx_pld_rst_n),
				.pld_polinv_tx(in_pld_polinv_tx),
				.pld_tx_clk(in_pld_tx_clk),
				.pld_tx_control({in_pld_tx_control[17], in_pld_tx_control[16], in_pld_tx_control[15], in_pld_tx_control[14], in_pld_tx_control[13], in_pld_tx_control[12], in_pld_tx_control[11], in_pld_tx_control[10], in_pld_tx_control[9], in_pld_tx_control[8], in_pld_tx_control[7], in_pld_tx_control[6], in_pld_tx_control[5], in_pld_tx_control[4], in_pld_tx_control[3], in_pld_tx_control[2], in_pld_tx_control[1], in_pld_tx_control[0]}),
				.pld_tx_data({in_pld_tx_data[127], in_pld_tx_data[126], in_pld_tx_data[125], in_pld_tx_data[124], in_pld_tx_data[123], in_pld_tx_data[122], in_pld_tx_data[121], in_pld_tx_data[120], in_pld_tx_data[119], in_pld_tx_data[118], in_pld_tx_data[117], in_pld_tx_data[116], in_pld_tx_data[115], in_pld_tx_data[114], in_pld_tx_data[113], in_pld_tx_data[112], in_pld_tx_data[111], in_pld_tx_data[110], in_pld_tx_data[109], in_pld_tx_data[108], in_pld_tx_data[107], in_pld_tx_data[106], in_pld_tx_data[105], in_pld_tx_data[104], in_pld_tx_data[103], in_pld_tx_data[102], in_pld_tx_data[101], in_pld_tx_data[100], in_pld_tx_data[99], in_pld_tx_data[98], in_pld_tx_data[97], in_pld_tx_data[96], in_pld_tx_data[95], in_pld_tx_data[94], in_pld_tx_data[93], in_pld_tx_data[92], in_pld_tx_data[91], in_pld_tx_data[90], in_pld_tx_data[89], in_pld_tx_data[88], in_pld_tx_data[87], in_pld_tx_data[86], in_pld_tx_data[85], in_pld_tx_data[84], in_pld_tx_data[83], in_pld_tx_data[82], in_pld_tx_data[81], in_pld_tx_data[80], in_pld_tx_data[79], in_pld_tx_data[78], in_pld_tx_data[77], in_pld_tx_data[76], in_pld_tx_data[75], in_pld_tx_data[74], in_pld_tx_data[73], in_pld_tx_data[72], in_pld_tx_data[71], in_pld_tx_data[70], in_pld_tx_data[69], in_pld_tx_data[68], in_pld_tx_data[67], in_pld_tx_data[66], in_pld_tx_data[65], in_pld_tx_data[64], in_pld_tx_data[63], in_pld_tx_data[62], in_pld_tx_data[61], in_pld_tx_data[60], in_pld_tx_data[59], in_pld_tx_data[58], in_pld_tx_data[57], in_pld_tx_data[56], in_pld_tx_data[55], in_pld_tx_data[54], in_pld_tx_data[53], in_pld_tx_data[52], in_pld_tx_data[51], in_pld_tx_data[50], in_pld_tx_data[49], in_pld_tx_data[48], in_pld_tx_data[47], in_pld_tx_data[46], in_pld_tx_data[45], in_pld_tx_data[44], in_pld_tx_data[43], in_pld_tx_data[42], in_pld_tx_data[41], in_pld_tx_data[40], in_pld_tx_data[39], in_pld_tx_data[38], in_pld_tx_data[37], in_pld_tx_data[36], in_pld_tx_data[35], in_pld_tx_data[34], in_pld_tx_data[33], in_pld_tx_data[32], in_pld_tx_data[31], in_pld_tx_data[30], in_pld_tx_data[29], in_pld_tx_data[28], in_pld_tx_data[27], in_pld_tx_data[26], in_pld_tx_data[25], in_pld_tx_data[24], in_pld_tx_data[23], in_pld_tx_data[22], in_pld_tx_data[21], in_pld_tx_data[20], in_pld_tx_data[19], in_pld_tx_data[18], in_pld_tx_data[17], in_pld_tx_data[16], in_pld_tx_data[15], in_pld_tx_data[14], in_pld_tx_data[13], in_pld_tx_data[12], in_pld_tx_data[11], in_pld_tx_data[10], in_pld_tx_data[9], in_pld_tx_data[8], in_pld_tx_data[7], in_pld_tx_data[6], in_pld_tx_data[5], in_pld_tx_data[4], in_pld_tx_data[3], in_pld_tx_data[2], in_pld_tx_data[1], in_pld_tx_data[0]}),
				.pld_txelecidle(in_pld_txelecidle),
				.pld_uhsif_tx_clk(in_pld_uhsif_tx_clk),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.hip_clk_out_div_by_2_wire(),
				.hip_clk_out_wire(),
				.int_pldif_pmaif_tx_pld_clk(),
				.pld_10g_tx_burst_en_exe_10g_fastreg(),
				.pld_10g_tx_burst_en_exe_plddirect_reg(),
				.pld_10g_tx_data_valid_2ff_delay1_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay3_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg(),
				.pld_10g_tx_data_valid_fastreg(),
				.pld_10g_tx_data_valid_plddirect_fastreg(),
				.pld_pcs_tx_clk_out_pma_wire(),
				.pld_pma_tx_clk_out_wire(),
				.pld_pmaif_tx_pld_rst_n_reg(),
				.pld_polinv_tx_10g_pcsdirect_reg(),
				.pld_polinv_tx_8g_reg(),
				.pld_polinv_tx_pat_reg(),
				.pld_tx_clk_fifo(),
				.pld_tx_control_fifo(),
				.pld_tx_control_hi_10g_reg(),
				.pld_tx_control_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_10g_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_8g_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_control_lo_plddirect_fastreg(),
				.pld_tx_control_lo_plddirect_reg(),
				.pld_tx_data_hi_reg(),
				.pld_tx_data_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_10g_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_8g_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_data_lo_plddirect_fastreg(),
				.pld_tx_data_lo_plddirect_reg(),
				.pld_uhsif_reg(),
				.pma_tx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_hip_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6:0] = 7'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17:0] = 18'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8:0] = 9'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127:0] = 128'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4:0] = 5'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2:0] = 3'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_full = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_full_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out = 1'b0;
		end // if not generate
		
		//output assignments
		assign out_avmmreaddata_hssi_10g_rx_pcs = {w_hssi_10g_rx_pcs_avmmreaddata[7], w_hssi_10g_rx_pcs_avmmreaddata[6], w_hssi_10g_rx_pcs_avmmreaddata[5], w_hssi_10g_rx_pcs_avmmreaddata[4], w_hssi_10g_rx_pcs_avmmreaddata[3], w_hssi_10g_rx_pcs_avmmreaddata[2], w_hssi_10g_rx_pcs_avmmreaddata[1], w_hssi_10g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_10g_tx_pcs = {w_hssi_10g_tx_pcs_avmmreaddata[7], w_hssi_10g_tx_pcs_avmmreaddata[6], w_hssi_10g_tx_pcs_avmmreaddata[5], w_hssi_10g_tx_pcs_avmmreaddata[4], w_hssi_10g_tx_pcs_avmmreaddata[3], w_hssi_10g_tx_pcs_avmmreaddata[2], w_hssi_10g_tx_pcs_avmmreaddata[1], w_hssi_10g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_rx_pcs = {w_hssi_8g_rx_pcs_avmmreaddata[7], w_hssi_8g_rx_pcs_avmmreaddata[6], w_hssi_8g_rx_pcs_avmmreaddata[5], w_hssi_8g_rx_pcs_avmmreaddata[4], w_hssi_8g_rx_pcs_avmmreaddata[3], w_hssi_8g_rx_pcs_avmmreaddata[2], w_hssi_8g_rx_pcs_avmmreaddata[1], w_hssi_8g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_tx_pcs = {w_hssi_8g_tx_pcs_avmmreaddata[7], w_hssi_8g_tx_pcs_avmmreaddata[6], w_hssi_8g_tx_pcs_avmmreaddata[5], w_hssi_8g_tx_pcs_avmmreaddata[4], w_hssi_8g_tx_pcs_avmmreaddata[3], w_hssi_8g_tx_pcs_avmmreaddata[2], w_hssi_8g_tx_pcs_avmmreaddata[1], w_hssi_8g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pcs_pma_interface = {w_hssi_common_pcs_pma_interface_avmmreaddata[7], w_hssi_common_pcs_pma_interface_avmmreaddata[6], w_hssi_common_pcs_pma_interface_avmmreaddata[5], w_hssi_common_pcs_pma_interface_avmmreaddata[4], w_hssi_common_pcs_pma_interface_avmmreaddata[3], w_hssi_common_pcs_pma_interface_avmmreaddata[2], w_hssi_common_pcs_pma_interface_avmmreaddata[1], w_hssi_common_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pld_pcs_interface = {w_hssi_common_pld_pcs_interface_avmmreaddata[7], w_hssi_common_pld_pcs_interface_avmmreaddata[6], w_hssi_common_pld_pcs_interface_avmmreaddata[5], w_hssi_common_pld_pcs_interface_avmmreaddata[4], w_hssi_common_pld_pcs_interface_avmmreaddata[3], w_hssi_common_pld_pcs_interface_avmmreaddata[2], w_hssi_common_pld_pcs_interface_avmmreaddata[1], w_hssi_common_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_rx_pcs = {w_hssi_fifo_rx_pcs_avmmreaddata[7], w_hssi_fifo_rx_pcs_avmmreaddata[6], w_hssi_fifo_rx_pcs_avmmreaddata[5], w_hssi_fifo_rx_pcs_avmmreaddata[4], w_hssi_fifo_rx_pcs_avmmreaddata[3], w_hssi_fifo_rx_pcs_avmmreaddata[2], w_hssi_fifo_rx_pcs_avmmreaddata[1], w_hssi_fifo_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_tx_pcs = {w_hssi_fifo_tx_pcs_avmmreaddata[7], w_hssi_fifo_tx_pcs_avmmreaddata[6], w_hssi_fifo_tx_pcs_avmmreaddata[5], w_hssi_fifo_tx_pcs_avmmreaddata[4], w_hssi_fifo_tx_pcs_avmmreaddata[3], w_hssi_fifo_tx_pcs_avmmreaddata[2], w_hssi_fifo_tx_pcs_avmmreaddata[1], w_hssi_fifo_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_rx_pcs = {w_hssi_gen3_rx_pcs_avmmreaddata[7], w_hssi_gen3_rx_pcs_avmmreaddata[6], w_hssi_gen3_rx_pcs_avmmreaddata[5], w_hssi_gen3_rx_pcs_avmmreaddata[4], w_hssi_gen3_rx_pcs_avmmreaddata[3], w_hssi_gen3_rx_pcs_avmmreaddata[2], w_hssi_gen3_rx_pcs_avmmreaddata[1], w_hssi_gen3_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_tx_pcs = {w_hssi_gen3_tx_pcs_avmmreaddata[7], w_hssi_gen3_tx_pcs_avmmreaddata[6], w_hssi_gen3_tx_pcs_avmmreaddata[5], w_hssi_gen3_tx_pcs_avmmreaddata[4], w_hssi_gen3_tx_pcs_avmmreaddata[3], w_hssi_gen3_tx_pcs_avmmreaddata[2], w_hssi_gen3_tx_pcs_avmmreaddata[1], w_hssi_gen3_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_rx_pcs = {w_hssi_krfec_rx_pcs_avmmreaddata[7], w_hssi_krfec_rx_pcs_avmmreaddata[6], w_hssi_krfec_rx_pcs_avmmreaddata[5], w_hssi_krfec_rx_pcs_avmmreaddata[4], w_hssi_krfec_rx_pcs_avmmreaddata[3], w_hssi_krfec_rx_pcs_avmmreaddata[2], w_hssi_krfec_rx_pcs_avmmreaddata[1], w_hssi_krfec_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_tx_pcs = {w_hssi_krfec_tx_pcs_avmmreaddata[7], w_hssi_krfec_tx_pcs_avmmreaddata[6], w_hssi_krfec_tx_pcs_avmmreaddata[5], w_hssi_krfec_tx_pcs_avmmreaddata[4], w_hssi_krfec_tx_pcs_avmmreaddata[3], w_hssi_krfec_tx_pcs_avmmreaddata[2], w_hssi_krfec_tx_pcs_avmmreaddata[1], w_hssi_krfec_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen1_2 = {w_hssi_pipe_gen1_2_avmmreaddata[7], w_hssi_pipe_gen1_2_avmmreaddata[6], w_hssi_pipe_gen1_2_avmmreaddata[5], w_hssi_pipe_gen1_2_avmmreaddata[4], w_hssi_pipe_gen1_2_avmmreaddata[3], w_hssi_pipe_gen1_2_avmmreaddata[2], w_hssi_pipe_gen1_2_avmmreaddata[1], w_hssi_pipe_gen1_2_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen3 = {w_hssi_pipe_gen3_avmmreaddata[7], w_hssi_pipe_gen3_avmmreaddata[6], w_hssi_pipe_gen3_avmmreaddata[5], w_hssi_pipe_gen3_avmmreaddata[4], w_hssi_pipe_gen3_avmmreaddata[3], w_hssi_pipe_gen3_avmmreaddata[2], w_hssi_pipe_gen3_avmmreaddata[1], w_hssi_pipe_gen3_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pcs_pma_interface = {w_hssi_rx_pcs_pma_interface_avmmreaddata[7], w_hssi_rx_pcs_pma_interface_avmmreaddata[6], w_hssi_rx_pcs_pma_interface_avmmreaddata[5], w_hssi_rx_pcs_pma_interface_avmmreaddata[4], w_hssi_rx_pcs_pma_interface_avmmreaddata[3], w_hssi_rx_pcs_pma_interface_avmmreaddata[2], w_hssi_rx_pcs_pma_interface_avmmreaddata[1], w_hssi_rx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pld_pcs_interface = {w_hssi_rx_pld_pcs_interface_avmmreaddata[7], w_hssi_rx_pld_pcs_interface_avmmreaddata[6], w_hssi_rx_pld_pcs_interface_avmmreaddata[5], w_hssi_rx_pld_pcs_interface_avmmreaddata[4], w_hssi_rx_pld_pcs_interface_avmmreaddata[3], w_hssi_rx_pld_pcs_interface_avmmreaddata[2], w_hssi_rx_pld_pcs_interface_avmmreaddata[1], w_hssi_rx_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pcs_pma_interface = {w_hssi_tx_pcs_pma_interface_avmmreaddata[7], w_hssi_tx_pcs_pma_interface_avmmreaddata[6], w_hssi_tx_pcs_pma_interface_avmmreaddata[5], w_hssi_tx_pcs_pma_interface_avmmreaddata[4], w_hssi_tx_pcs_pma_interface_avmmreaddata[3], w_hssi_tx_pcs_pma_interface_avmmreaddata[2], w_hssi_tx_pcs_pma_interface_avmmreaddata[1], w_hssi_tx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pld_pcs_interface = {w_hssi_tx_pld_pcs_interface_avmmreaddata[7], w_hssi_tx_pld_pcs_interface_avmmreaddata[6], w_hssi_tx_pld_pcs_interface_avmmreaddata[5], w_hssi_tx_pld_pcs_interface_avmmreaddata[4], w_hssi_tx_pld_pcs_interface_avmmreaddata[3], w_hssi_tx_pld_pcs_interface_avmmreaddata[2], w_hssi_tx_pld_pcs_interface_avmmreaddata[1], w_hssi_tx_pld_pcs_interface_avmmreaddata[0]};
		assign out_blockselect_hssi_10g_rx_pcs = w_hssi_10g_rx_pcs_blockselect;
		assign out_blockselect_hssi_10g_tx_pcs = w_hssi_10g_tx_pcs_blockselect;
		assign out_blockselect_hssi_8g_rx_pcs = w_hssi_8g_rx_pcs_blockselect;
		assign out_blockselect_hssi_8g_tx_pcs = w_hssi_8g_tx_pcs_blockselect;
		assign out_blockselect_hssi_common_pcs_pma_interface = w_hssi_common_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_common_pld_pcs_interface = w_hssi_common_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_fifo_rx_pcs = w_hssi_fifo_rx_pcs_blockselect;
		assign out_blockselect_hssi_fifo_tx_pcs = w_hssi_fifo_tx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_rx_pcs = w_hssi_gen3_rx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_tx_pcs = w_hssi_gen3_tx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_rx_pcs = w_hssi_krfec_rx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_tx_pcs = w_hssi_krfec_tx_pcs_blockselect;
		assign out_blockselect_hssi_pipe_gen1_2 = w_hssi_pipe_gen1_2_blockselect;
		assign out_blockselect_hssi_pipe_gen3 = w_hssi_pipe_gen3_blockselect;
		assign out_blockselect_hssi_rx_pcs_pma_interface = w_hssi_rx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_rx_pld_pcs_interface = w_hssi_rx_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_tx_pcs_pma_interface = w_hssi_tx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_tx_pld_pcs_interface = w_hssi_tx_pld_pcs_interface_blockselect;
		assign out_bond_pcs10g_out_bot = {w_hssi_10g_tx_pcs_distdwn_out_rden, w_hssi_10g_tx_pcs_distdwn_out_wren, w_hssi_10g_tx_pcs_distdwn_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs10g_out_top = {w_hssi_10g_tx_pcs_distup_out_rden, w_hssi_10g_tx_pcs_distup_out_wren, w_hssi_10g_tx_pcs_distup_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs8g_out_bot = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down, w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_down, w_hssi_8g_tx_pcs_wr_enable_out_chnl_down, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_down, w_hssi_8g_rx_pcs_wr_enable_out_chnl_down, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[0]};
		assign out_bond_pcs8g_out_top = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up, w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_up, w_hssi_8g_tx_pcs_wr_enable_out_chnl_up, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_up, w_hssi_8g_rx_pcs_wr_enable_out_chnl_up, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[0]};
		assign out_bond_pmaif_out_bot = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[0]};
		assign out_bond_pmaif_out_top = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[0]};
		assign out_hip_clk_out = {w_hssi_common_pld_pcs_interface_hip_cmn_clk[1], w_hssi_common_pld_pcs_interface_hip_cmn_clk[0], w_hssi_tx_pld_pcs_interface_hip_tx_clk};
		assign out_hip_ctrl_out = {w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[4], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[3], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[2], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[1], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[0], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[0]};
		assign out_hip_iocsr_rdy = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
		assign out_hip_iocsr_rdy_dly = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
		assign out_hip_nfrzdrv = w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
		assign out_hip_npor = w_hssi_common_pld_pcs_interface_hip_npor;
		assign out_hip_rx_data = {w_hssi_rx_pld_pcs_interface_hip_rx_data[50], w_hssi_rx_pld_pcs_interface_hip_rx_data[49], w_hssi_rx_pld_pcs_interface_hip_rx_data[48], w_hssi_rx_pld_pcs_interface_hip_rx_data[47], w_hssi_rx_pld_pcs_interface_hip_rx_data[46], w_hssi_rx_pld_pcs_interface_hip_rx_data[45], w_hssi_rx_pld_pcs_interface_hip_rx_data[44], w_hssi_rx_pld_pcs_interface_hip_rx_data[43], w_hssi_rx_pld_pcs_interface_hip_rx_data[42], w_hssi_rx_pld_pcs_interface_hip_rx_data[41], w_hssi_rx_pld_pcs_interface_hip_rx_data[40], w_hssi_rx_pld_pcs_interface_hip_rx_data[39], w_hssi_rx_pld_pcs_interface_hip_rx_data[38], w_hssi_rx_pld_pcs_interface_hip_rx_data[37], w_hssi_rx_pld_pcs_interface_hip_rx_data[36], w_hssi_rx_pld_pcs_interface_hip_rx_data[35], w_hssi_rx_pld_pcs_interface_hip_rx_data[34], w_hssi_rx_pld_pcs_interface_hip_rx_data[33], w_hssi_rx_pld_pcs_interface_hip_rx_data[32], w_hssi_rx_pld_pcs_interface_hip_rx_data[31], w_hssi_rx_pld_pcs_interface_hip_rx_data[30], w_hssi_rx_pld_pcs_interface_hip_rx_data[29], w_hssi_rx_pld_pcs_interface_hip_rx_data[28], w_hssi_rx_pld_pcs_interface_hip_rx_data[27], w_hssi_rx_pld_pcs_interface_hip_rx_data[26], w_hssi_rx_pld_pcs_interface_hip_rx_data[25], w_hssi_rx_pld_pcs_interface_hip_rx_data[24], w_hssi_rx_pld_pcs_interface_hip_rx_data[23], w_hssi_rx_pld_pcs_interface_hip_rx_data[22], w_hssi_rx_pld_pcs_interface_hip_rx_data[21], w_hssi_rx_pld_pcs_interface_hip_rx_data[20], w_hssi_rx_pld_pcs_interface_hip_rx_data[19], w_hssi_rx_pld_pcs_interface_hip_rx_data[18], w_hssi_rx_pld_pcs_interface_hip_rx_data[17], w_hssi_rx_pld_pcs_interface_hip_rx_data[16], w_hssi_rx_pld_pcs_interface_hip_rx_data[15], w_hssi_rx_pld_pcs_interface_hip_rx_data[14], w_hssi_rx_pld_pcs_interface_hip_rx_data[13], w_hssi_rx_pld_pcs_interface_hip_rx_data[12], w_hssi_rx_pld_pcs_interface_hip_rx_data[11], w_hssi_rx_pld_pcs_interface_hip_rx_data[10], w_hssi_rx_pld_pcs_interface_hip_rx_data[9], w_hssi_rx_pld_pcs_interface_hip_rx_data[8], w_hssi_rx_pld_pcs_interface_hip_rx_data[7], w_hssi_rx_pld_pcs_interface_hip_rx_data[6], w_hssi_rx_pld_pcs_interface_hip_rx_data[5], w_hssi_rx_pld_pcs_interface_hip_rx_data[4], w_hssi_rx_pld_pcs_interface_hip_rx_data[3], w_hssi_rx_pld_pcs_interface_hip_rx_data[2], w_hssi_rx_pld_pcs_interface_hip_rx_data[1], w_hssi_rx_pld_pcs_interface_hip_rx_data[0]};
		assign out_hip_usermode = w_hssi_common_pld_pcs_interface_hip_usermode;
		assign out_pld_10g_krfec_rx_blk_lock = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
		assign out_pld_10g_krfec_rx_diag_data_status = {w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1], w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[0]};
		assign out_pld_10g_krfec_rx_frame = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
		assign out_pld_10g_krfec_tx_frame = w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
		assign out_pld_10g_rx_align_val = w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
		assign out_pld_10g_rx_crc32_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
		assign out_pld_10g_rx_data_valid = w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
		assign out_pld_10g_rx_empty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
		assign out_pld_10g_rx_fifo_del = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
		assign out_pld_10g_rx_fifo_insert = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
		assign out_pld_10g_rx_fifo_num = {w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[3], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[2], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[1], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[0]};
		assign out_pld_10g_rx_frame_lock = w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
		assign out_pld_10g_rx_hi_ber = w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
		assign out_pld_10g_rx_oflw_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
		assign out_pld_10g_rx_pempty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
		assign out_pld_10g_rx_pfull = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
		assign out_pld_10g_tx_burst_en_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
		assign out_pld_10g_tx_empty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
		assign out_pld_10g_tx_fifo_num = {w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[2], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[1], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[0]};
		assign out_pld_10g_tx_full = w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
		assign out_pld_10g_tx_pempty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
		assign out_pld_10g_tx_pfull = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
		assign out_pld_10g_tx_wordslip_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
		assign out_pld_8g_a1a2_k1k2_flag = {w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[2], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[1], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[0]};
		assign out_pld_8g_empty_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
		assign out_pld_8g_empty_rx = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
		assign out_pld_8g_empty_tx = w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
		assign out_pld_8g_full_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
		assign out_pld_8g_full_rx = w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
		assign out_pld_8g_full_tx = w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
		assign out_pld_8g_rxelecidle = w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
		assign out_pld_8g_signal_detect_out = w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
		assign out_pld_8g_wa_boundary = {w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0]};
		assign out_pld_krfec_tx_alignment = w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
		assign out_pld_pcs_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
		assign out_pld_pcs_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
		assign out_pld_pma_adapt_done = w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
		assign out_pld_pma_clkdiv_rx_user = w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
		assign out_pld_pma_clkdiv_tx_user = w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
		assign out_pld_pma_clklow = w_hssi_common_pld_pcs_interface_pld_pma_clklow;
		assign out_pld_pma_fref = w_hssi_common_pld_pcs_interface_pld_pma_fref;
		assign out_pld_pma_hclk = w_hssi_common_pld_pcs_interface_pld_pma_hclk;
		assign out_pld_pma_pcie_sw_done = {w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1], w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[0]};
		assign out_pld_pma_pfdmode_lock = w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
		assign out_pld_pma_reserved_in = {w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[3], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[2], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[1], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[0]};
		assign out_pld_pma_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
		assign out_pld_pma_rx_detect_valid = w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
		assign out_pld_pma_rx_found = w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
		assign out_pld_pma_rxpll_lock = w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
		assign out_pld_pma_signal_ok = w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
		assign out_pld_pma_testbus = {w_hssi_common_pld_pcs_interface_pld_pma_testbus[7], w_hssi_common_pld_pcs_interface_pld_pma_testbus[6], w_hssi_common_pld_pcs_interface_pld_pma_testbus[5], w_hssi_common_pld_pcs_interface_pld_pma_testbus[4], w_hssi_common_pld_pcs_interface_pld_pma_testbus[3], w_hssi_common_pld_pcs_interface_pld_pma_testbus[2], w_hssi_common_pld_pcs_interface_pld_pma_testbus[1], w_hssi_common_pld_pcs_interface_pld_pma_testbus[0]};
		assign out_pld_pma_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
		assign out_pld_pmaif_mask_tx_pll = w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
		assign out_pld_reserved_out = {w_hssi_common_pld_pcs_interface_pld_reserved_out[9], w_hssi_common_pld_pcs_interface_pld_reserved_out[8], w_hssi_common_pld_pcs_interface_pld_reserved_out[7], w_hssi_common_pld_pcs_interface_pld_reserved_out[6], w_hssi_common_pld_pcs_interface_pld_reserved_out[5], w_hssi_common_pld_pcs_interface_pld_reserved_out[4], w_hssi_common_pld_pcs_interface_pld_reserved_out[3], w_hssi_common_pld_pcs_interface_pld_reserved_out[2], w_hssi_common_pld_pcs_interface_pld_reserved_out[1], w_hssi_common_pld_pcs_interface_pld_reserved_out[0]};
		assign out_pld_rx_control = {w_hssi_rx_pld_pcs_interface_pld_rx_control[19], w_hssi_rx_pld_pcs_interface_pld_rx_control[18], w_hssi_rx_pld_pcs_interface_pld_rx_control[17], w_hssi_rx_pld_pcs_interface_pld_rx_control[16], w_hssi_rx_pld_pcs_interface_pld_rx_control[15], w_hssi_rx_pld_pcs_interface_pld_rx_control[14], w_hssi_rx_pld_pcs_interface_pld_rx_control[13], w_hssi_rx_pld_pcs_interface_pld_rx_control[12], w_hssi_rx_pld_pcs_interface_pld_rx_control[11], w_hssi_rx_pld_pcs_interface_pld_rx_control[10], w_hssi_rx_pld_pcs_interface_pld_rx_control[9], w_hssi_rx_pld_pcs_interface_pld_rx_control[8], w_hssi_rx_pld_pcs_interface_pld_rx_control[7], w_hssi_rx_pld_pcs_interface_pld_rx_control[6], w_hssi_rx_pld_pcs_interface_pld_rx_control[5], w_hssi_rx_pld_pcs_interface_pld_rx_control[4], w_hssi_rx_pld_pcs_interface_pld_rx_control[3], w_hssi_rx_pld_pcs_interface_pld_rx_control[2], w_hssi_rx_pld_pcs_interface_pld_rx_control[1], w_hssi_rx_pld_pcs_interface_pld_rx_control[0]};
		assign out_pld_rx_data = {w_hssi_rx_pld_pcs_interface_pld_rx_data[127], w_hssi_rx_pld_pcs_interface_pld_rx_data[126], w_hssi_rx_pld_pcs_interface_pld_rx_data[125], w_hssi_rx_pld_pcs_interface_pld_rx_data[124], w_hssi_rx_pld_pcs_interface_pld_rx_data[123], w_hssi_rx_pld_pcs_interface_pld_rx_data[122], w_hssi_rx_pld_pcs_interface_pld_rx_data[121], w_hssi_rx_pld_pcs_interface_pld_rx_data[120], w_hssi_rx_pld_pcs_interface_pld_rx_data[119], w_hssi_rx_pld_pcs_interface_pld_rx_data[118], w_hssi_rx_pld_pcs_interface_pld_rx_data[117], w_hssi_rx_pld_pcs_interface_pld_rx_data[116], w_hssi_rx_pld_pcs_interface_pld_rx_data[115], w_hssi_rx_pld_pcs_interface_pld_rx_data[114], w_hssi_rx_pld_pcs_interface_pld_rx_data[113], w_hssi_rx_pld_pcs_interface_pld_rx_data[112], w_hssi_rx_pld_pcs_interface_pld_rx_data[111], w_hssi_rx_pld_pcs_interface_pld_rx_data[110], w_hssi_rx_pld_pcs_interface_pld_rx_data[109], w_hssi_rx_pld_pcs_interface_pld_rx_data[108], w_hssi_rx_pld_pcs_interface_pld_rx_data[107], w_hssi_rx_pld_pcs_interface_pld_rx_data[106], w_hssi_rx_pld_pcs_interface_pld_rx_data[105], w_hssi_rx_pld_pcs_interface_pld_rx_data[104], w_hssi_rx_pld_pcs_interface_pld_rx_data[103], w_hssi_rx_pld_pcs_interface_pld_rx_data[102], w_hssi_rx_pld_pcs_interface_pld_rx_data[101], w_hssi_rx_pld_pcs_interface_pld_rx_data[100], w_hssi_rx_pld_pcs_interface_pld_rx_data[99], w_hssi_rx_pld_pcs_interface_pld_rx_data[98], w_hssi_rx_pld_pcs_interface_pld_rx_data[97], w_hssi_rx_pld_pcs_interface_pld_rx_data[96], w_hssi_rx_pld_pcs_interface_pld_rx_data[95], w_hssi_rx_pld_pcs_interface_pld_rx_data[94], w_hssi_rx_pld_pcs_interface_pld_rx_data[93], w_hssi_rx_pld_pcs_interface_pld_rx_data[92], w_hssi_rx_pld_pcs_interface_pld_rx_data[91], w_hssi_rx_pld_pcs_interface_pld_rx_data[90], w_hssi_rx_pld_pcs_interface_pld_rx_data[89], w_hssi_rx_pld_pcs_interface_pld_rx_data[88], w_hssi_rx_pld_pcs_interface_pld_rx_data[87], w_hssi_rx_pld_pcs_interface_pld_rx_data[86], w_hssi_rx_pld_pcs_interface_pld_rx_data[85], w_hssi_rx_pld_pcs_interface_pld_rx_data[84], w_hssi_rx_pld_pcs_interface_pld_rx_data[83], w_hssi_rx_pld_pcs_interface_pld_rx_data[82], w_hssi_rx_pld_pcs_interface_pld_rx_data[81], w_hssi_rx_pld_pcs_interface_pld_rx_data[80], w_hssi_rx_pld_pcs_interface_pld_rx_data[79], w_hssi_rx_pld_pcs_interface_pld_rx_data[78], w_hssi_rx_pld_pcs_interface_pld_rx_data[77], w_hssi_rx_pld_pcs_interface_pld_rx_data[76], w_hssi_rx_pld_pcs_interface_pld_rx_data[75], w_hssi_rx_pld_pcs_interface_pld_rx_data[74], w_hssi_rx_pld_pcs_interface_pld_rx_data[73], w_hssi_rx_pld_pcs_interface_pld_rx_data[72], w_hssi_rx_pld_pcs_interface_pld_rx_data[71], w_hssi_rx_pld_pcs_interface_pld_rx_data[70], w_hssi_rx_pld_pcs_interface_pld_rx_data[69], w_hssi_rx_pld_pcs_interface_pld_rx_data[68], w_hssi_rx_pld_pcs_interface_pld_rx_data[67], w_hssi_rx_pld_pcs_interface_pld_rx_data[66], w_hssi_rx_pld_pcs_interface_pld_rx_data[65], w_hssi_rx_pld_pcs_interface_pld_rx_data[64], w_hssi_rx_pld_pcs_interface_pld_rx_data[63], w_hssi_rx_pld_pcs_interface_pld_rx_data[62], w_hssi_rx_pld_pcs_interface_pld_rx_data[61], w_hssi_rx_pld_pcs_interface_pld_rx_data[60], w_hssi_rx_pld_pcs_interface_pld_rx_data[59], w_hssi_rx_pld_pcs_interface_pld_rx_data[58], w_hssi_rx_pld_pcs_interface_pld_rx_data[57], w_hssi_rx_pld_pcs_interface_pld_rx_data[56], w_hssi_rx_pld_pcs_interface_pld_rx_data[55], w_hssi_rx_pld_pcs_interface_pld_rx_data[54], w_hssi_rx_pld_pcs_interface_pld_rx_data[53], w_hssi_rx_pld_pcs_interface_pld_rx_data[52], w_hssi_rx_pld_pcs_interface_pld_rx_data[51], w_hssi_rx_pld_pcs_interface_pld_rx_data[50], w_hssi_rx_pld_pcs_interface_pld_rx_data[49], w_hssi_rx_pld_pcs_interface_pld_rx_data[48], w_hssi_rx_pld_pcs_interface_pld_rx_data[47], w_hssi_rx_pld_pcs_interface_pld_rx_data[46], w_hssi_rx_pld_pcs_interface_pld_rx_data[45], w_hssi_rx_pld_pcs_interface_pld_rx_data[44], w_hssi_rx_pld_pcs_interface_pld_rx_data[43], w_hssi_rx_pld_pcs_interface_pld_rx_data[42], w_hssi_rx_pld_pcs_interface_pld_rx_data[41], w_hssi_rx_pld_pcs_interface_pld_rx_data[40], w_hssi_rx_pld_pcs_interface_pld_rx_data[39], w_hssi_rx_pld_pcs_interface_pld_rx_data[38], w_hssi_rx_pld_pcs_interface_pld_rx_data[37], w_hssi_rx_pld_pcs_interface_pld_rx_data[36], w_hssi_rx_pld_pcs_interface_pld_rx_data[35], w_hssi_rx_pld_pcs_interface_pld_rx_data[34], w_hssi_rx_pld_pcs_interface_pld_rx_data[33], w_hssi_rx_pld_pcs_interface_pld_rx_data[32], w_hssi_rx_pld_pcs_interface_pld_rx_data[31], w_hssi_rx_pld_pcs_interface_pld_rx_data[30], w_hssi_rx_pld_pcs_interface_pld_rx_data[29], w_hssi_rx_pld_pcs_interface_pld_rx_data[28], w_hssi_rx_pld_pcs_interface_pld_rx_data[27], w_hssi_rx_pld_pcs_interface_pld_rx_data[26], w_hssi_rx_pld_pcs_interface_pld_rx_data[25], w_hssi_rx_pld_pcs_interface_pld_rx_data[24], w_hssi_rx_pld_pcs_interface_pld_rx_data[23], w_hssi_rx_pld_pcs_interface_pld_rx_data[22], w_hssi_rx_pld_pcs_interface_pld_rx_data[21], w_hssi_rx_pld_pcs_interface_pld_rx_data[20], w_hssi_rx_pld_pcs_interface_pld_rx_data[19], w_hssi_rx_pld_pcs_interface_pld_rx_data[18], w_hssi_rx_pld_pcs_interface_pld_rx_data[17], w_hssi_rx_pld_pcs_interface_pld_rx_data[16], w_hssi_rx_pld_pcs_interface_pld_rx_data[15], w_hssi_rx_pld_pcs_interface_pld_rx_data[14], w_hssi_rx_pld_pcs_interface_pld_rx_data[13], w_hssi_rx_pld_pcs_interface_pld_rx_data[12], w_hssi_rx_pld_pcs_interface_pld_rx_data[11], w_hssi_rx_pld_pcs_interface_pld_rx_data[10], w_hssi_rx_pld_pcs_interface_pld_rx_data[9], w_hssi_rx_pld_pcs_interface_pld_rx_data[8], w_hssi_rx_pld_pcs_interface_pld_rx_data[7], w_hssi_rx_pld_pcs_interface_pld_rx_data[6], w_hssi_rx_pld_pcs_interface_pld_rx_data[5], w_hssi_rx_pld_pcs_interface_pld_rx_data[4], w_hssi_rx_pld_pcs_interface_pld_rx_data[3], w_hssi_rx_pld_pcs_interface_pld_rx_data[2], w_hssi_rx_pld_pcs_interface_pld_rx_data[1], w_hssi_rx_pld_pcs_interface_pld_rx_data[0]};
		assign out_pld_rx_prbs_done = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
		assign out_pld_rx_prbs_err = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
		assign out_pld_test_data = {w_hssi_common_pld_pcs_interface_pld_test_data[19], w_hssi_common_pld_pcs_interface_pld_test_data[18], w_hssi_common_pld_pcs_interface_pld_test_data[17], w_hssi_common_pld_pcs_interface_pld_test_data[16], w_hssi_common_pld_pcs_interface_pld_test_data[15], w_hssi_common_pld_pcs_interface_pld_test_data[14], w_hssi_common_pld_pcs_interface_pld_test_data[13], w_hssi_common_pld_pcs_interface_pld_test_data[12], w_hssi_common_pld_pcs_interface_pld_test_data[11], w_hssi_common_pld_pcs_interface_pld_test_data[10], w_hssi_common_pld_pcs_interface_pld_test_data[9], w_hssi_common_pld_pcs_interface_pld_test_data[8], w_hssi_common_pld_pcs_interface_pld_test_data[7], w_hssi_common_pld_pcs_interface_pld_test_data[6], w_hssi_common_pld_pcs_interface_pld_test_data[5], w_hssi_common_pld_pcs_interface_pld_test_data[4], w_hssi_common_pld_pcs_interface_pld_test_data[3], w_hssi_common_pld_pcs_interface_pld_test_data[2], w_hssi_common_pld_pcs_interface_pld_test_data[1], w_hssi_common_pld_pcs_interface_pld_test_data[0]};
		assign out_pld_uhsif_lock = w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
		assign out_pld_uhsif_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
		assign out_pma_adapt_start = w_hssi_common_pcs_pma_interface_pma_adapt_start;
		assign out_pma_atpg_los_en_n = w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
		assign out_pma_csr_test_dis = w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
		assign out_pma_current_coeff = {w_hssi_common_pcs_pma_interface_pma_current_coeff[17], w_hssi_common_pcs_pma_interface_pma_current_coeff[16], w_hssi_common_pcs_pma_interface_pma_current_coeff[15], w_hssi_common_pcs_pma_interface_pma_current_coeff[14], w_hssi_common_pcs_pma_interface_pma_current_coeff[13], w_hssi_common_pcs_pma_interface_pma_current_coeff[12], w_hssi_common_pcs_pma_interface_pma_current_coeff[11], w_hssi_common_pcs_pma_interface_pma_current_coeff[10], w_hssi_common_pcs_pma_interface_pma_current_coeff[9], w_hssi_common_pcs_pma_interface_pma_current_coeff[8], w_hssi_common_pcs_pma_interface_pma_current_coeff[7], w_hssi_common_pcs_pma_interface_pma_current_coeff[6], w_hssi_common_pcs_pma_interface_pma_current_coeff[5], w_hssi_common_pcs_pma_interface_pma_current_coeff[4], w_hssi_common_pcs_pma_interface_pma_current_coeff[3], w_hssi_common_pcs_pma_interface_pma_current_coeff[2], w_hssi_common_pcs_pma_interface_pma_current_coeff[1], w_hssi_common_pcs_pma_interface_pma_current_coeff[0]};
		assign out_pma_current_rxpreset = {w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[1], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[0]};
		assign out_pma_early_eios = w_hssi_common_pcs_pma_interface_pma_early_eios;
		assign out_pma_eye_monitor = {w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0]};
		assign out_pma_interface_select = {w_hssi_common_pcs_pma_interface_pma_interface_select[1], w_hssi_common_pcs_pma_interface_pma_interface_select[0]};
		assign out_pma_ltd_b = w_hssi_common_pcs_pma_interface_pma_ltd_b;
		assign out_pma_ltr = w_hssi_common_pcs_pma_interface_pma_ltr;
		assign out_pma_nfrzdrv = w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
		assign out_pma_nrpi_freeze = w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
		assign out_pma_pcie_switch = {w_hssi_common_pcs_pma_interface_pma_pcie_switch[1], w_hssi_common_pcs_pma_interface_pma_pcie_switch[0]};
		assign out_pma_ppm_lock = w_hssi_common_pcs_pma_interface_pma_ppm_lock;
		assign out_pma_reserved_out = {w_hssi_common_pcs_pma_interface_pma_reserved_out[4], w_hssi_common_pcs_pma_interface_pma_reserved_out[3], w_hssi_common_pcs_pma_interface_pma_reserved_out[2], w_hssi_common_pcs_pma_interface_pma_reserved_out[1], w_hssi_common_pcs_pma_interface_pma_reserved_out[0]};
		assign out_pma_rs_lpbk_b = w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
		assign out_pma_rx_clkslip = w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
		assign out_pma_rx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
		assign out_pma_rxpma_rstb = w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
		assign out_pma_scan_mode_n = w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
		assign out_pma_scan_shift_n = w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
		assign out_pma_tx_bitslip = w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
		assign out_pma_tx_bonding_rstb = w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
		assign out_pma_tx_elec_idle = w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
		assign out_pma_tx_pma_data = {w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0]};
		assign out_pma_tx_qpi_pulldn = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
		assign out_pma_tx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
		assign out_pma_tx_txdetectrx = w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
		assign out_pma_txpma_rstb = w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	endgenerate
endmodule
module twentynm_pcs_rev_20nm4
	#(
	//PARAM_LIST_START
		parameter xcvr_native_mode = "mode_duplex",  // mode_duplex, mode_rx_only, mode_tx_only
		
		// parameters for twentynm_hssi_10g_rx_pcs
		parameter hssi_10g_rx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_align_del = "align_del_en", // align_del_dis|align_del_en
		parameter hssi_10g_rx_pcs_ber_bit_err_total_cnt = "bit_err_total_cnt_10g", // bit_err_total_cnt_10g
		parameter hssi_10g_rx_pcs_ber_clken = "ber_clk_dis", // ber_clk_dis|ber_clk_en
		parameter hssi_10g_rx_pcs_ber_xus_timer_window = 21'b100110001001010,
		parameter hssi_10g_rx_pcs_bitslip_mode = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_rx_pcs_blksync_bitslip_type = "bitslip_comb", // bitslip_comb|bitslip_reg
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_cnt = 3'b1,
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_type = "bitslip_match", // bitslip_match|bitslip_cnt
		parameter hssi_10g_rx_pcs_blksync_bypass = "blksync_bypass_dis", // blksync_bypass_dis|blksync_bypass_en
		parameter hssi_10g_rx_pcs_blksync_clken = "blksync_clk_dis", // blksync_clk_dis|blksync_clk_en
		parameter hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt = "enum_invalid_sh_cnt_10g", // enum_invalid_sh_cnt_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock = "knum_sh_cnt_postlock_10g", // knum_sh_cnt_postlock_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock = "knum_sh_cnt_prelock_10g", // knum_sh_cnt_prelock_10g
		parameter hssi_10g_rx_pcs_blksync_pipeln = "blksync_pipeln_dis", // blksync_pipeln_dis|blksync_pipeln_en
		parameter hssi_10g_rx_pcs_clr_errblk_cnt_en = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_control_del = "control_del_all", // control_del_all|control_del_none
		parameter hssi_10g_rx_pcs_crcchk_bypass = "crcchk_bypass_dis", // crcchk_bypass_dis|crcchk_bypass_en
		parameter hssi_10g_rx_pcs_crcchk_clken = "crcchk_clk_dis", // crcchk_clk_dis|crcchk_clk_en
		parameter hssi_10g_rx_pcs_crcchk_inv = "crcchk_inv_dis", // crcchk_inv_dis|crcchk_inv_en
		parameter hssi_10g_rx_pcs_crcchk_pipeln = "crcchk_pipeln_dis", // crcchk_pipeln_dis|crcchk_pipeln_en
		parameter hssi_10g_rx_pcs_crcflag_pipeln = "crcflag_pipeln_dis", // crcflag_pipeln_dis|crcflag_pipeln_en
		parameter hssi_10g_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_rx_pcs_dec64b66b_clken = "dec64b66b_clk_dis", // dec64b66b_clk_dis|dec64b66b_clk_en
		parameter hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass = "dec_64b66b_rxsm_bypass_dis", // dec_64b66b_rxsm_bypass_dis|dec_64b66b_rxsm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_bypass = "descrm_bypass_en", // descrm_bypass_dis|descrm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_clken = "descrm_clk_dis", // descrm_clk_dis|descrm_clk_en
		parameter hssi_10g_rx_pcs_descrm_mode = "async", // async|sync
		parameter hssi_10g_rx_pcs_descrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_dft_clk_out_sel = "rx_master_clk", // rx_master_clk|rx_gbexp_clk|rx_blksync_clk|rx_descrm_clk|rx_frmsync_clk|rx_64b66bdec_clk|rx_ber_clk|rx_rand_clk|rx_crcchk_clk|rx_wrfifo_clk|rx_rdfifo_clk|rx_fec_clk
		parameter hssi_10g_rx_pcs_dis_signal_ok = "dis_signal_ok_dis", // dis_signal_ok_dis|dis_signal_ok_en
		parameter hssi_10g_rx_pcs_dispchk_bypass = "dispchk_bypass_dis", // dispchk_bypass_dis|dispchk_bypass_en
		parameter hssi_10g_rx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_rx_pcs_fast_path = "fast_path_dis", // fast_path_dis|fast_path_en
		parameter hssi_10g_rx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_rx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_rx_pcs_fifo_double_read = "fifo_double_read_dis", // fifo_double_read_dis|fifo_double_read_en
		parameter hssi_10g_rx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_rx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_rx_pcs_force_align = "force_align_dis", // force_align_dis|force_align_en
		parameter hssi_10g_rx_pcs_frmsync_bypass = "frmsync_bypass_dis", // frmsync_bypass_dis|frmsync_bypass_en
		parameter hssi_10g_rx_pcs_frmsync_clken = "frmsync_clk_dis", // frmsync_clk_dis|frmsync_clk_en
		parameter hssi_10g_rx_pcs_frmsync_enum_scrm = "enum_scrm_default", // enum_scrm_default
		parameter hssi_10g_rx_pcs_frmsync_enum_sync = "enum_sync_default", // enum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_flag_type = "all_framing_words", // all_framing_words|location_only
		parameter hssi_10g_rx_pcs_frmsync_knum_sync = "knum_sync_default", // knum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_mfrm_length = 16'b100000000000,
		parameter hssi_10g_rx_pcs_frmsync_pipeln = "frmsync_pipeln_dis", // frmsync_pipeln_dis|frmsync_pipeln_en
		parameter hssi_10g_rx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_rx_pcs_gb_rx_idwidth = "width_32", // width_40|width_32|width_64
		parameter hssi_10g_rx_pcs_gb_rx_odwidth = "width_66", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_rx_pcs_gbexp_clken = "gbexp_clk_dis", // gbexp_clk_dis|gbexp_clk_en
		parameter hssi_10g_rx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_10g_rx_pcs_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_rx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_rx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_rx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_rx_pcs_pld_if_type = "fifo", // fifo|reg
		parameter hssi_10g_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_rx_pcs_rand_clken = "rand_clk_dis", // rand_clk_dis|rand_clk_en
		parameter hssi_10g_rx_pcs_rd_clk_sel = "rd_rx_pma_clk", // rd_rx_pld_clk|rd_rx_pma_clk|rd_refclk_dig
		parameter hssi_10g_rx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_rx_pcs_rx_fifo_write_ctrl = "blklock_stops", // blklock_stops|blklock_ignore
		parameter hssi_10g_rx_pcs_rx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_rx_pcs_rx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_rx_pcs_rx_signal_ok_sel = "synchronized_ver", // synchronized_ver|nonsync_ver
		parameter hssi_10g_rx_pcs_rx_sm_bypass = "rx_sm_bypass_dis", // rx_sm_bypass_dis|rx_sm_bypass_en
		parameter hssi_10g_rx_pcs_rx_sm_hiber = "rx_sm_hiber_en", // rx_sm_hiber_en|rx_sm_hiber_dis
		parameter hssi_10g_rx_pcs_rx_sm_pipeln = "rx_sm_pipeln_dis", // rx_sm_pipeln_dis|rx_sm_pipeln_en
		parameter hssi_10g_rx_pcs_rx_testbus_sel = "crc32_chk_testbus1", // crc32_chk_testbus1|crc32_chk_testbus2|frame_sync_testbus1|frame_sync_testbus2|dec64b66b_testbus|rxsm_testbus|ber_testbus|blksync_testbus1|blksync_testbus2|gearbox_exp_testbus|random_ver_testbus|descramble_testbus|blank_testbus|rx_fifo_testbus1|rx_fifo_testbus2
		parameter hssi_10g_rx_pcs_rx_true_b2b = "b2b", // single|b2b
		parameter hssi_10g_rx_pcs_rxfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_rx_pcs_rxfifo_full = "full_default", // full_default
		parameter hssi_10g_rx_pcs_rxfifo_mode = "phase_comp", // register_mode|clk_comp_10g|generic_interlaken|generic_basic|phase_comp|phase_comp_dv
		parameter hssi_10g_rx_pcs_rxfifo_pempty = 5'b10,
		parameter hssi_10g_rx_pcs_rxfifo_pfull = 5'b10111,
		parameter hssi_10g_rx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_rx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_rx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_10g_tx_pcs
		parameter hssi_10g_tx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_bitslip_en = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_10g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_10g_tx_pcs_comp_cnt = 8'b0,
		parameter hssi_10g_tx_pcs_compin_sel = "compin_master", // compin_master|compin_slave_top|compin_slave_bot|compin_default
		parameter hssi_10g_tx_pcs_crcgen_bypass = "crcgen_bypass_dis", // crcgen_bypass_dis|crcgen_bypass_en
		parameter hssi_10g_tx_pcs_crcgen_clken = "crcgen_clk_dis", // crcgen_clk_dis|crcgen_clk_en
		parameter hssi_10g_tx_pcs_crcgen_err = "crcgen_err_dis", // crcgen_err_dis|crcgen_err_en
		parameter hssi_10g_tx_pcs_crcgen_inv = "crcgen_inv_dis", // crcgen_inv_dis|crcgen_inv_en
		parameter hssi_10g_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_tx_pcs_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_10g_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_tx_pcs_dft_clk_out_sel = "tx_master_clk", // tx_master_clk|tx_rdfifo_clk|tx_frmgen_clk|tx_crcgen_clk|tx_64b66benc_txsm_clk|tx_scrm_clk|tx_dispgen_clk|tx_gbred_clk|tx_wrfifo_clk|tx_fec_clk
		parameter hssi_10g_tx_pcs_dispgen_bypass = "dispgen_bypass_dis", // dispgen_bypass_dis|dispgen_bypass_en
		parameter hssi_10g_tx_pcs_dispgen_clken = "dispgen_clk_dis", // dispgen_clk_dis|dispgen_clk_en
		parameter hssi_10g_tx_pcs_dispgen_err = "dispgen_err_dis", // dispgen_err_dis|dispgen_err_en
		parameter hssi_10g_tx_pcs_dispgen_pipeln = "dispgen_pipeln_dis", // dispgen_pipeln_dis|dispgen_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_bypass_pipeln = "distdwn_bypass_pipeln_dis", // distdwn_bypass_pipeln_dis|distdwn_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_master = "distdwn_master_en", // distdwn_master_en|distdwn_master_dis
		parameter hssi_10g_tx_pcs_distup_bypass_pipeln = "distup_bypass_pipeln_dis", // distup_bypass_pipeln_dis|distup_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distup_master = "distup_master_en", // distup_master_en|distup_master_dis
		parameter hssi_10g_tx_pcs_dv_bond = "dv_bond_dis", // dv_bond_en|dv_bond_dis
		parameter hssi_10g_tx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_tx_pcs_enc64b66b_txsm_clken = "enc64b66b_txsm_clk_dis", // enc64b66b_txsm_clk_dis|enc64b66b_txsm_clk_en
		parameter hssi_10g_tx_pcs_enc_64b66b_txsm_bypass = "enc_64b66b_txsm_bypass_dis", // enc_64b66b_txsm_bypass_dis|enc_64b66b_txsm_bypass_en
		parameter hssi_10g_tx_pcs_fastpath = "fastpath_dis", // fastpath_dis|fastpath_en
		parameter hssi_10g_tx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_tx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_tx_pcs_fifo_double_write = "fifo_double_write_dis", // fifo_double_write_dis|fifo_double_write_en
		parameter hssi_10g_tx_pcs_fifo_reg_fast = "fifo_reg_fast_dis", // fifo_reg_fast_dis|fifo_reg_fast_en
		parameter hssi_10g_tx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_tx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_tx_pcs_frmgen_burst = "frmgen_burst_dis", // frmgen_burst_dis|frmgen_burst_en
		parameter hssi_10g_tx_pcs_frmgen_bypass = "frmgen_bypass_dis", // frmgen_bypass_dis|frmgen_bypass_en
		parameter hssi_10g_tx_pcs_frmgen_clken = "frmgen_clk_dis", // frmgen_clk_dis|frmgen_clk_en
		parameter hssi_10g_tx_pcs_frmgen_mfrm_length = 16'b100000000000,
		parameter hssi_10g_tx_pcs_frmgen_pipeln = "frmgen_pipeln_dis", // frmgen_pipeln_dis|frmgen_pipeln_en
		parameter hssi_10g_tx_pcs_frmgen_pyld_ins = "frmgen_pyld_ins_dis", // frmgen_pyld_ins_dis|frmgen_pyld_ins_en
		parameter hssi_10g_tx_pcs_frmgen_wordslip = "frmgen_wordslip_dis", // frmgen_wordslip_dis|frmgen_wordslip_en
		parameter hssi_10g_tx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_tx_pcs_gb_pipeln_bypass = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_gb_tx_idwidth = "width_50", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_tx_pcs_gb_tx_odwidth = "width_32", // width_32|width_40|width_64
		parameter hssi_10g_tx_pcs_gbred_clken = "gbred_clk_dis", // gbred_clk_dis|gbred_clk_en
		parameter hssi_10g_tx_pcs_indv = "indv_en", // indv_en|indv_dis
		parameter hssi_10g_tx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_tx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_tx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_tx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del6|phcomp_rd_del5|phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_tx_pcs_pld_if_type = "fifo", // fifo|reg|fastreg
		parameter hssi_10g_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_tx_pcs_pseudo_random = "all_0", // two_lf|all_0
		parameter hssi_10g_tx_pcs_pseudo_seed_a = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_pseudo_seed_b = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_random_disp = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_tx_pcs_scrm_bypass = "scrm_bypass_dis", // scrm_bypass_dis|scrm_bypass_en
		parameter hssi_10g_tx_pcs_scrm_clken = "scrm_clk_dis", // scrm_clk_dis|scrm_clk_en
		parameter hssi_10g_tx_pcs_scrm_mode = "async", // async|sync
		parameter hssi_10g_tx_pcs_scrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_sh_err = "sh_err_dis", // sh_err_dis|sh_err_en
		parameter hssi_10g_tx_pcs_sop_mark = "sop_mark_dis", // sop_mark_en|sop_mark_dis
		parameter hssi_10g_tx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_tx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_tx_pcs_tx_scrm_err = "scrm_err_dis", // scrm_err_dis|scrm_err_en
		parameter hssi_10g_tx_pcs_tx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_tx_pcs_tx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_tx_pcs_tx_sm_bypass = "tx_sm_bypass_dis", // tx_sm_bypass_dis|tx_sm_bypass_en
		parameter hssi_10g_tx_pcs_tx_sm_pipeln = "tx_sm_pipeln_dis", // tx_sm_pipeln_dis|tx_sm_pipeln_en
		parameter hssi_10g_tx_pcs_tx_testbus_sel = "crc32_gen_testbus1", // crc32_gen_testbus1|crc32_gen_testbus2|disp_gen_testbus1|disp_gen_testbus2|frame_gen_testbus1|frame_gen_testbus2|enc64b66b_testbus|txsm_testbus|tx_cp_bond_testbus|gearbox_red_testbus|scramble_testbus|blank_testbus|tx_fifo_testbus1|tx_fifo_testbus2
		parameter hssi_10g_tx_pcs_txfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_tx_pcs_txfifo_full = "full_default", // full_default
		parameter hssi_10g_tx_pcs_txfifo_mode = "phase_comp", // register_mode|interlaken_generic|basic_generic|phase_comp
		parameter hssi_10g_tx_pcs_txfifo_pempty = 4'b10,
		parameter hssi_10g_tx_pcs_txfifo_pfull = 4'b1011,
		parameter hssi_10g_tx_pcs_wr_clk_sel = "wr_tx_pma_clk", // wr_tx_pld_clk|wr_tx_pma_clk|wr_refclk_dig
		parameter hssi_10g_tx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_8g_rx_pcs
		parameter hssi_8g_rx_pcs_auto_error_replacement = "dis_err_replace", // dis_err_replace|en_err_replace
		parameter hssi_8g_rx_pcs_auto_speed_nego = "dis_asn", // dis_asn|en_asn_g2_freq_scal
		parameter hssi_8g_rx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_rx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_rx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_rx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_rx_pcs_byte_deserializer = "dis_bds", // dis_bds|en_bds_by_2|en_bds_by_4|en_bds_by_2_det
		parameter hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask = "dis_rxvalid_mask", // dis_rxvalid_mask|en_rxvalid_mask
		parameter hssi_8g_rx_pcs_clkcmp_pattern_n = 20'b0,
		parameter hssi_8g_rx_pcs_clkcmp_pattern_p = 20'b0,
		parameter hssi_8g_rx_pcs_clock_gate_bds_dec_asn = "dis_bds_dec_asn_clk_gating", // dis_bds_dec_asn_clk_gating|en_bds_dec_asn_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_cdr_eidle = "dis_cdr_eidle_clk_gating", // dis_cdr_eidle_clk_gating|en_cdr_eidle_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk = "dis_dw_pc_wrclk_gating", // dis_dw_pc_wrclk_gating|en_dw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_rd = "dis_dw_rm_rdclk_gating", // dis_dw_rm_rdclk_gating|en_dw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_wr = "dis_dw_rm_wrclk_gating", // dis_dw_rm_wrclk_gating|en_dw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_wa = "dis_dw_wa_clk_gating", // dis_dw_wa_clk_gating|en_dw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_pc_rdclk = "dis_pc_rdclk_gating", // dis_pc_rdclk_gating|en_pc_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk = "dis_sw_pc_wrclk_gating", // dis_sw_pc_wrclk_gating|en_sw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_rd = "dis_sw_rm_rdclk_gating", // dis_sw_rm_rdclk_gating|en_sw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_wr = "dis_sw_rm_wrclk_gating", // dis_sw_rm_wrclk_gating|en_sw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_wa = "dis_sw_wa_clk_gating", // dis_sw_wa_clk_gating|en_sw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_observation_in_pld_core = "internal_sw_wa_clk", // internal_sw_wa_clk|internal_dw_wa_clk|internal_cdr_eidle_clk|internal_sm_rm_wr_clk|internal_dw_rm_wr_clk|internal_clk_2_b|internal_sw_rm_rd_clk|internal_dw_rm_rd_clk|internal_sw_rx_wr_clk|internal_dw_rx_wr_clk|internal_rx_rd_clk|internal_rx_pma_clk_gen3|internal_rx_rcvd_clk_gen3
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_rx_pcs_eidle_entry_eios = "dis_eidle_eios", // dis_eidle_eios|en_eidle_eios
		parameter hssi_8g_rx_pcs_eidle_entry_iei = "dis_eidle_iei", // dis_eidle_iei|en_eidle_iei
		parameter hssi_8g_rx_pcs_eidle_entry_sd = "dis_eidle_sd", // dis_eidle_sd|en_eidle_sd
		parameter hssi_8g_rx_pcs_eightb_tenb_decoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_rx_pcs_err_flags_sel = "err_flags_wa", // err_flags_wa|err_flags_8b10b
		parameter hssi_8g_rx_pcs_fixed_pat_det = "dis_fixed_patdet", // dis_fixed_patdet|en_fixed_patdet
		parameter hssi_8g_rx_pcs_fixed_pat_num = 4'b1111,
		parameter hssi_8g_rx_pcs_force_signal_detect = "en_force_signal_detect", // en_force_signal_detect|dis_force_signal_detect
		parameter hssi_8g_rx_pcs_gen3_clk_en = "disable_clk", // disable_clk|enable_clk
		parameter hssi_8g_rx_pcs_gen3_rx_clk_sel = "rcvd_clk", // en_dig_clk1_8g|rcvd_clk
		parameter hssi_8g_rx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // en_dig_clk2_8g|tx_pma_clk
		parameter hssi_8g_rx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_rx_pcs_ibm_invalid_code = "dis_ibm_invalid_code", // dis_ibm_invalid_code|en_ibm_invalid_code
		parameter hssi_8g_rx_pcs_invalid_code_flag_only = "dis_invalid_code_only", // dis_invalid_code_only|en_invalid_code_only
		parameter hssi_8g_rx_pcs_pad_or_edb_error_replace = "replace_edb", // replace_edb|replace_edb_dynamic|replace_pad
		parameter hssi_8g_rx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_rx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_rx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_rx_pcs_pipe_if_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_8g_rx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_rx_pcs_polinv_8b10b_dec = "dis_polinv_8b10b_dec", // dis_polinv_8b10b_dec|en_polinv_8b10b_dec
		parameter hssi_8g_rx_pcs_prot_mode = "gige", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic_rm_enable|basic_rm_disable|disabled_prot_mode
		parameter hssi_8g_rx_pcs_rate_match = "dis_rm", // dis_rm|gige_rm|pipe_rm|pipe_rm_0ppm|sw_basic_rm|dw_basic_rm
		parameter hssi_8g_rx_pcs_rate_match_del_thres = "dis_rm_del_thres", // dis_rm_del_thres|gige_rm_del_thres|pipe_rm_del_thres|pipe_rm_0ppm_del_thres|sw_basic_rm_del_thres|dw_basic_rm_del_thres
		parameter hssi_8g_rx_pcs_rate_match_empty_thres = "dis_rm_empty_thres", // dis_rm_empty_thres|gige_rm_empty_thres|pipe_rm_empty_thres|pipe_rm_0ppm_empty_thres|sw_basic_rm_empty_thres|dw_basic_rm_empty_thres
		parameter hssi_8g_rx_pcs_rate_match_full_thres = "dis_rm_full_thres", // dis_rm_full_thres|gige_rm_full_thres|pipe_rm_full_thres|pipe_rm_0ppm_full_thres|sw_basic_rm_full_thres|dw_basic_rm_full_thres
		parameter hssi_8g_rx_pcs_rate_match_ins_thres = "dis_rm_ins_thres", // dis_rm_ins_thres|gige_rm_ins_thres|pipe_rm_ins_thres|pipe_rm_0ppm_ins_thres|sw_basic_rm_ins_thres|dw_basic_rm_ins_thres
		parameter hssi_8g_rx_pcs_rate_match_start_thres = "dis_rm_start_thres", // dis_rm_start_thres|gige_rm_start_thres|pipe_rm_start_thres|pipe_rm_0ppm_start_thres|sw_basic_rm_start_thres|dw_basic_rm_start_thres
		parameter hssi_8g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_rx_pcs_rx_clk2 = "rcvd_clk_clk2", // rcvd_clk_clk2|tx_pma_clock_clk2|refclk_dig2_clk2
		parameter hssi_8g_rx_pcs_rx_clk_free_running = "en_rx_clk_free_run", // dis_rx_clk_free_run|en_rx_clk_free_run
		parameter hssi_8g_rx_pcs_rx_pcs_urst = "en_rx_pcs_urst", // dis_rx_pcs_urst|en_rx_pcs_urst
		parameter hssi_8g_rx_pcs_rx_rcvd_clk = "rcvd_clk_rcvd_clk", // rcvd_clk_rcvd_clk|tx_pma_clock_rcvd_clk
		parameter hssi_8g_rx_pcs_rx_rd_clk = "pld_rx_clk", // pld_rx_clk|rx_clk
		parameter hssi_8g_rx_pcs_rx_refclk = "dis_refclk_sel", // dis_refclk_sel|en_refclk_sel
		parameter hssi_8g_rx_pcs_rx_wr_clk = "rx_clk2_div_1_2_4", // rx_clk2_div_1_2_4|txfifo_rd_clk
		parameter hssi_8g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_rx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_rx_pcs_sync_sm_idle_eios = "dis_syncsm_idle", // dis_syncsm_idle|en_syncsm_idle
		parameter hssi_8g_rx_pcs_test_bus_sel = "tx_testbus", // tx_testbus|tx_ctrl_plane_testbus|wa_testbus|rm_testbus|rx_ctrl_testbus|pcie_ctrl_testbus|rx_ctrl_plane_testbus
		parameter hssi_8g_rx_pcs_tx_rx_parallel_loopback = "dis_plpbk", // dis_plpbk|en_plpbk
		parameter hssi_8g_rx_pcs_wa_boundary_lock_ctrl = "bit_slip", // bit_slip|sync_sm|deterministic_latency|auto_align_pld_ctrl
		parameter hssi_8g_rx_pcs_wa_clk_slip_spacing = 10'b10000,
		parameter hssi_8g_rx_pcs_wa_det_latency_sync_status_beh = "assert_sync_status_non_imm", // assert_sync_status_imm|assert_sync_status_non_imm|dont_care_assert_sync
		parameter hssi_8g_rx_pcs_wa_disp_err_flag = "dis_disp_err_flag", // dis_disp_err_flag|en_disp_err_flag
		parameter hssi_8g_rx_pcs_wa_kchar = "dis_kchar", // dis_kchar|en_kchar
		parameter hssi_8g_rx_pcs_wa_pd = "wa_pd_10", // wa_pd_7|wa_pd_10|wa_pd_20|wa_pd_40|wa_pd_8_sw|wa_pd_8_dw|wa_pd_16_sw|wa_pd_16_dw|wa_pd_32
		parameter hssi_8g_rx_pcs_wa_pd_data = 40'b0,
		parameter hssi_8g_rx_pcs_wa_pd_polarity = "dis_pd_both_pol", // dis_pd_both_pol|en_pd_both_pol|dont_care_both_pol
		parameter hssi_8g_rx_pcs_wa_pld_controlled = "dis_pld_ctrl", // dis_pld_ctrl|pld_ctrl_sw|rising_edge_sensitive_dw|level_sensitive_dw
		parameter hssi_8g_rx_pcs_wa_renumber_data = 6'b0,
		parameter hssi_8g_rx_pcs_wa_rgnumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rknumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rosnumber_data = 2'b0,
		parameter hssi_8g_rx_pcs_wa_rvnumber_data = 13'b0,
		parameter hssi_8g_rx_pcs_wa_sync_sm_ctrl = "gige_sync_sm", // gige_sync_sm|pipe_sync_sm|sw_basic_sync_sm|dw_basic_sync_sm|fibre_channel_sync_sm
		parameter hssi_8g_rx_pcs_wait_cnt = 12'b0,
		
		// parameters for twentynm_hssi_8g_tx_pcs
		parameter hssi_8g_tx_pcs_auto_speed_nego_gen2 = "dis_asn_g2", // dis_asn_g2|en_asn_g2_freq_scal
		parameter hssi_8g_tx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_tx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_tx_pcs_byte_serializer = "dis_bs", // dis_bs|en_bs_by_2|en_bs_by_4
		parameter hssi_8g_tx_pcs_clock_gate_bs_enc = "dis_bs_enc_clk_gating", // dis_bs_enc_clk_gating|en_bs_enc_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_dw_fifowr = "dis_dw_fifowr_clk_gating", // dis_dw_fifowr_clk_gating|en_dw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_fiford = "dis_fiford_clk_gating", // dis_fiford_clk_gating|en_fiford_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_sw_fifowr = "dis_sw_fifowr_clk_gating", // dis_sw_fifowr_clk_gating|en_sw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_observation_in_pld_core = "internal_refclk_b", // internal_refclk_b|internal_fifo_rd_clk|internal_sw_fifo_wr_clk|internal_dw_fifo_wr_clk|internal_tx_clk_out_gen3|internal_pipe_tx_clk_out_gen3
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_tx_pcs_data_selection_8b10b_encoder_input = "normal_data_path", // normal_data_path|gige_idle_conversion
		parameter hssi_8g_tx_pcs_dynamic_clk_switch = "dis_dyn_clk_switch", // dis_dyn_clk_switch|en_dyn_clk_switch
		parameter hssi_8g_tx_pcs_eightb_tenb_disp_ctrl = "dis_disp_ctrl", // dis_disp_ctrl|en_disp_ctrl|en_ib_disp_ctrl
		parameter hssi_8g_tx_pcs_eightb_tenb_encoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_tx_pcs_force_echar = "dis_force_echar", // dis_force_echar|en_force_echar
		parameter hssi_8g_tx_pcs_force_kchar = "dis_force_kchar", // dis_force_kchar|en_force_kchar
		parameter hssi_8g_tx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // dis_tx_clk|tx_pma_clk
		parameter hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel = "func_clk", // dis_tx_pipe_clk|func_clk
		parameter hssi_8g_tx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_tx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_tx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_tx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_tx_pcs_phfifo_write_clk_sel = "pld_tx_clk", // pld_tx_clk|tx_clk
		parameter hssi_8g_tx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_tx_pcs_prot_mode = "basic", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic|disabled_prot_mode
		parameter hssi_8g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_tx_pcs_refclk_b_clk_sel = "tx_pma_clock", // tx_pma_clock|refclk_dig
		parameter hssi_8g_tx_pcs_revloop_back_rm = "dis_rev_loopback_rx_rm", // dis_rev_loopback_rx_rm|en_rev_loopback_rx_rm
		parameter hssi_8g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_tx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_tx_pcs_tx_bitslip = "dis_tx_bitslip", // dis_tx_bitslip|en_tx_bitslip
		parameter hssi_8g_tx_pcs_tx_compliance_controlled_disparity = "dis_txcompliance", // dis_txcompliance|en_txcompliance_pipe2p0|en_txcompliance_pipe3p0
		parameter hssi_8g_tx_pcs_tx_fast_pld_reg = "dis_tx_fast_pld_reg", // dis_tx_fast_pld_reg|en_tx_fast_pld_reg
		parameter hssi_8g_tx_pcs_txclk_freerun = "dis_freerun_tx", // dis_freerun_tx|en_freerun_tx
		parameter hssi_8g_tx_pcs_txpcs_urst = "en_txpcs_urst", // dis_txpcs_urst|en_txpcs_urst
		
		// parameters for twentynm_hssi_common_pcs_pma_interface
		parameter hssi_common_pcs_pma_interface_asn_clk_enable = "false", // false|true
		parameter hssi_common_pcs_pma_interface_asn_enable = "dis_asn", // dis_asn|en_asn
		parameter hssi_common_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|pcie_gen3
		parameter hssi_common_pcs_pma_interface_bypass_early_eios = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pcie_switch = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_ltr = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_sw_done = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_ppm_lock = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_txdetectrx = "false", // false|true
		parameter hssi_common_pcs_pma_interface_cdr_control = "en_cdr_ctrl", // dis_cdr_ctrl|en_cdr_ctrl
		parameter hssi_common_pcs_pma_interface_cid_enable = "en_cid_mode", // dis_cid_mode|en_cid_mode
		parameter hssi_common_pcs_pma_interface_cp_cons_sel = "cp_cons_default", // cp_cons_master|cp_cons_slave_abv|cp_cons_slave_blw|cp_cons_default
		parameter hssi_common_pcs_pma_interface_cp_dwn_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_cp_up_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_blw|ctrl_slave_abv
		parameter hssi_common_pcs_pma_interface_data_mask_count = 16'b100111000100,
		parameter hssi_common_pcs_pma_interface_data_mask_count_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_dft_observation_clock_selection = "dft_clk_obsrv_tx0", // dft_clk_obsrv_tx0|dft_clk_obsrv_tx1|dft_clk_obsrv_tx2|dft_clk_obsrv_tx3|dft_clk_obsrv_tx4|dft_clk_obsrv_rx|dft_clk_obsrv_hclk|dft_clk_obsrv_fref|dft_clk_obsrv_clklow|dft_clk_obsrv_asn0|dft_clk_obsrv_asn1
		parameter hssi_common_pcs_pma_interface_early_eios_counter = 8'b110010,
		parameter hssi_common_pcs_pma_interface_force_freqdet = "force_freqdet_dis", // force_freqdet_dis|force1_freqdet_en|force0_freqdet_en
		parameter hssi_common_pcs_pma_interface_free_run_clk_enable = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ignore_sigdet_g23 = "false", // false|true
		parameter hssi_common_pcs_pma_interface_pc_en_counter = 7'b110111,
		parameter hssi_common_pcs_pma_interface_pc_rst_counter = 5'b10111,
		parameter hssi_common_pcs_pma_interface_pcie_hip_mode = "hip_disable", // hip_enable|hip_disable
		parameter hssi_common_pcs_pma_interface_ph_fifo_reg_mode = "phfifo_reg_mode_dis", // phfifo_reg_mode_dis|phfifo_reg_mode_en
		parameter hssi_common_pcs_pma_interface_phfifo_flush_wait = 6'b100100,
		parameter hssi_common_pcs_pma_interface_pipe_if_g3pcs = "pipe_if_8gpcs", // pipe_if_g3pcs|pipe_if_8gpcs
		parameter hssi_common_pcs_pma_interface_pma_done_counter = 18'b101010101110011000,
		parameter hssi_common_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_common_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_common_pcs_pma_interface_ppm_cnt_rst = "ppm_cnt_rst_dis", // ppm_cnt_rst_dis|ppm_cnt_rst_en
		parameter hssi_common_pcs_pma_interface_ppm_deassert_early = "deassert_early_dis", // deassert_early_dis|deassert_early_en
		parameter hssi_common_pcs_pma_interface_ppm_det_buckets = "ppm_100_bucket", // disable_prot|ppm_300_bucket|ppm_100_bucket|ppm_300_100_bucket
		parameter hssi_common_pcs_pma_interface_ppm_gen1_2_cnt = "cnt_32k", // cnt_32k|cnt_64k
		parameter hssi_common_pcs_pma_interface_ppm_post_eidle_delay = "cnt_200_cycles", // cnt_200_cycles|cnt_400_cycles
		parameter hssi_common_pcs_pma_interface_ppmsel = "ppmsel_300", // ppmsel_disable|ppmsel_5000|ppmsel_2500|ppmsel_1000|ppmsel_500|ppmsel_300|ppmsel_250|ppmsel_200|ppmsel_125|ppmsel_100|ppmsel_62p5|ppm_other
		parameter hssi_common_pcs_pma_interface_prot_mode = "disable_prot_mode", // disable_prot_mode|pipe_g12|pipe_g3|other_protocols
		parameter hssi_common_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_common_pcs_pma_interface_rxvalid_mask = "rxvalid_mask_en", // rxvalid_mask_dis|rxvalid_mask_en
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter = 12'b100111000100,
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_sim_mode = "disable", // disable|enable
		parameter hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en = "true", // false|true
		parameter hssi_common_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_common_pcs_pma_interface_testout_sel = "ppm_det_test", // ppm_det_test|asn_test|pma_pll_test|rxpmaif_test|prbs_gen_test|prbs_ver_test|uhsif_1_test|uhsif_2_test|uhsif_3_test
		parameter hssi_common_pcs_pma_interface_wait_clk_on_off_timer = 4'b100,
		parameter hssi_common_pcs_pma_interface_wait_pipe_synchronizing = 5'b10111,
		parameter hssi_common_pcs_pma_interface_wait_send_syncp_fbkp = 11'b11111010,
		
		// parameters for twentynm_hssi_common_pld_pcs_interface
		parameter hssi_common_pld_pcs_interface_dft_clk_out_en = "dft_clk_out_disable", // dft_clk_out_disable|dft_clk_out_enable
		parameter hssi_common_pld_pcs_interface_dft_clk_out_sel = "teng_rx_dft_clk", // teng_rx_dft_clk|teng_tx_dft_clk|eightg_rx_dft_clk|eightg_tx_dft_clk|pmaif_dft_clk
		parameter hssi_common_pld_pcs_interface_hrdrstctrl_en = "hrst_dis", // hrst_dis|hrst_en
		parameter hssi_common_pld_pcs_interface_pcs_testbus_block_sel = "eightg", // eightg|g3pcs|teng|krfec|pma_if
		parameter hssi_common_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_fifo_rx_pcs
		parameter hssi_fifo_rx_pcs_double_read_mode = "double_read_dis", // double_read_en|double_read_dis
		parameter hssi_fifo_rx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_fifo_tx_pcs
		parameter hssi_fifo_tx_pcs_double_write_mode = "double_write_dis", // double_write_en|double_write_dis
		parameter hssi_fifo_tx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_gen3_rx_pcs
		parameter hssi_gen3_rx_pcs_block_sync = "enable_block_sync", // bypass_block_sync|enable_block_sync
		parameter hssi_gen3_rx_pcs_block_sync_sm = "enable_blk_sync_sm", // disable_blk_sync_sm|enable_blk_sync_sm
		parameter hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn = "enable", // disable|enable
		parameter hssi_gen3_rx_pcs_lpbk_force = "lpbk_frce_dis", // lpbk_frce_dis|lpbk_frce_en
		parameter hssi_gen3_rx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_rx_pcs_rate_match_fifo = "enable_rm_fifo_600ppm", // bypass_rm_fifo|enable_rm_fifo_600ppm|enable_rm_fifo_0ppm
		parameter hssi_gen3_rx_pcs_rate_match_fifo_latency = "regular_latency", // regular_latency|low_latency
		parameter hssi_gen3_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_gen3_rx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_b4gb_par_lpbk = "b4gb_par_lpbk_dis", // b4gb_par_lpbk_dis|b4gb_par_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_force_balign = "en_force_balign", // en_force_balign|dis_force_balign
		parameter hssi_gen3_rx_pcs_rx_ins_del_one_skip = "ins_del_one_skip_en", // ins_del_one_skip_dis|ins_del_one_skip_en
		parameter hssi_gen3_rx_pcs_rx_num_fixed_pat = 4'b1000,
		parameter hssi_gen3_rx_pcs_rx_test_out_sel = "rx_test_out0", // rx_test_out0|rx_test_out1
		parameter hssi_gen3_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_gen3_tx_pcs
		parameter hssi_gen3_tx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_tx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_gen3_tx_pcs_tx_bitslip = 5'b0,
		parameter hssi_gen3_tx_pcs_tx_gbox_byp = "bypass_gbox", // bypass_gbox|enable_gbox
		
		// parameters for twentynm_hssi_krfec_rx_pcs
		parameter hssi_krfec_rx_pcs_blksync_cor_en = "detect", // detect|correct
		parameter hssi_krfec_rx_pcs_bypass_gb = "bypass_dis", // bypass_dis|bypass_en
		parameter hssi_krfec_rx_pcs_clr_ctrl = "both_enabled", // both_enabled|corr_cnt_only|uncorr_cnt_only
		parameter hssi_krfec_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_rx_pcs_dv_start = "with_blklock", // with_blksync|with_blklock
		parameter hssi_krfec_rx_pcs_err_mark_type = "err_mark_10g", // err_mark_10g|err_mark_40g
		parameter hssi_krfec_rx_pcs_error_marking_en = "err_mark_dis", // err_mark_dis|err_mark_en
		parameter hssi_krfec_rx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_krfec_rx_pcs_parity_invalid_enum = 8'b1000,
		parameter hssi_krfec_rx_pcs_parity_valid_num = 4'b100,
		parameter hssi_krfec_rx_pcs_pipeln_blksync = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_descrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errcorrect = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_ind = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_lfsr = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_loc = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_pat = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_gearbox = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_syndrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_trans_dec = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_rx_pcs_receive_order = "receive_lsb", // receive_lsb|receive_msb
		parameter hssi_krfec_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_krfec_rx_pcs_rx_testbus_sel = "overall", // overall|fast_search|fast_search_cntrs|blksync|blksync_cntrs|decoder_master_sm|decoder_master_sm_cntrs|syndrm_sm|syndrm1|syndrm2|errtrap_sm|errtrap_ind1|errtrap_ind2|errtrap_ind3|errtrap_ind4|errtrap_ind5|errtrap_loc|errtrap_pat1|errtrap_pat2|errtrap_pat3|errtrap_pat4|decoder_rd_sm|gb_and_trans
		parameter hssi_krfec_rx_pcs_signal_ok_en = "sig_ok_dis", // sig_ok_dis|sig_ok_en
		parameter hssi_krfec_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_krfec_tx_pcs
		parameter hssi_krfec_tx_pcs_burst_err = "burst_err_dis", // burst_err_dis|burst_err_en
		parameter hssi_krfec_tx_pcs_burst_err_len = "burst_err_len1", // burst_err_len1|burst_err_len2|burst_err_len3|burst_err_len4|burst_err_len5|burst_err_len6|burst_err_len7|burst_err_len8|burst_err_len9|burst_err_len10|burst_err_len11|burst_err_len12|burst_err_len13|burst_err_len14|burst_err_len15|burst_err_len16
		parameter hssi_krfec_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_tx_pcs_enc_frame_query = "enc_query_dis", // enc_query_dis|enc_query_en
		parameter hssi_krfec_tx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_encoder = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_scrambler = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_krfec_tx_pcs_transcode_err = "trans_err_dis", // trans_err_dis|trans_err_en
		parameter hssi_krfec_tx_pcs_transmit_order = "transmit_lsb", // transmit_lsb|transmit_msb
		parameter hssi_krfec_tx_pcs_tx_testbus_sel = "overall", // overall|encoder1|encoder2|scramble1|scramble2|scramble3|gearbox
		
		// parameters for twentynm_hssi_pipe_gen1_2
		parameter hssi_pipe_gen1_2_elec_idle_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_error_replace_pad = "replace_edb", // replace_edb|replace_pad
		parameter hssi_pipe_gen1_2_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_pipe_gen1_2_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen1_2_phystatus_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_phystatus_rst_toggle = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen1_2_pipe_byte_de_serializer_en = "dont_care_bds", // dis_bds|en_bds_by_2|dont_care_bds
		parameter hssi_pipe_gen1_2_prot_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|basic|disabled_prot_mode
		parameter hssi_pipe_gen1_2_reconfig_settings = "{}", // 
		parameter hssi_pipe_gen1_2_rx_pipe_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_pipe_gen1_2_rxdetect_bypass = "dis_rxdetect_bypass", // dis_rxdetect_bypass|en_rxdetect_bypass
		parameter hssi_pipe_gen1_2_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen1_2_tx_pipe_enable = "dis_pipe_tx", // dis_pipe_tx|en_pipe_tx|en_pipe3_tx
		parameter hssi_pipe_gen1_2_txswing = "dis_txswing", // dis_txswing|en_txswing
		
		// parameters for twentynm_hssi_pipe_gen3
		parameter hssi_pipe_gen3_bypass_rx_detection_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_rx_preset = 3'b0,
		parameter hssi_pipe_gen3_bypass_rx_preset_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_tx_coefficent = 18'b0,
		parameter hssi_pipe_gen3_bypass_tx_coefficent_enable = "false", // false|true
		parameter hssi_pipe_gen3_elecidle_delay_g3 = 3'b110,
		parameter hssi_pipe_gen3_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen3_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|disable_pcs
		parameter hssi_pipe_gen3_phy_status_delay_g12 = 3'b101,
		parameter hssi_pipe_gen3_phy_status_delay_g3 = 3'b101,
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g12 = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g3 = "dis_phystatus_rst_toggle_g3", // dis_phystatus_rst_toggle_g3|en_phystatus_rst_toggle_g3
		parameter hssi_pipe_gen3_rate_match_pad_insertion = "dis_rm_fifo_pad_ins", // dis_rm_fifo_pad_ins|en_rm_fifo_pad_ins
		parameter hssi_pipe_gen3_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen3_test_out_sel = "disable_test_out", // tx_test_out|rx_test_out|pipe_test_out1|pipe_test_out2|pipe_test_out3|pipe_ctrl_test_out|disable_test_out
		
		// parameters for twentynm_hssi_rx_pcs_pma_interface
		parameter hssi_rx_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|ten_g_pcs|direct_pld
		parameter hssi_rx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pcs_pma_interface_clkslip_sel = "pld", // pld|slip_eight_g_pcs
		parameter hssi_rx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pcs_pma_interface_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_rx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_rx_pcs_pma_interface_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_rx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_rx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_rx_pcs_pma_interface_prbs_ver = "prbs_off", // prbs_off|prbs_31|prbs_15|prbs_23|prbs_9|prbs_7
		parameter hssi_rx_pcs_pma_interface_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion = "rx_dyn_polinv_dis", // rx_dyn_polinv_dis|rx_dyn_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_lpbk_en = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok = "unforce_sig_ok", // unforce_sig_ok|force_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mask = "prbsmask128", // prbsmask128|prbsmask256|prbsmask512|prbsmask1024
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mode = "teng_mode", // teng_mode|eightg_mode
		parameter hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel = "sel_sig_det", // sel_sig_det|sel_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_static_polarity_inversion = "rx_stat_polinv_dis", // rx_stat_polinv_dis|rx_stat_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en = "uhsif_lpbk_dis", // uhsif_lpbk_dis|uhsif_lpbk_en
		parameter hssi_rx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_rx_pld_pcs_interface
		parameter hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx = "enable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx = "pma_64b_rx", // pma_32b_rx|pma_40b_rx|pma_64b_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_baser_mode_rx|interlaken_mode_rx|sfis_mode_rx|teng_sdi_mode_rx|basic_mode_rx|test_prp_mode_rx|test_prp_krfec_mode_rx|teng_1588_mode_rx|teng_baser_krfec_mode_rx|teng_1588_krfec_mode_rx|basic_krfec_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx = "disabled_prot_mode_rx", // pipe_g1_rx|pipe_g2_rx|pipe_g3_rx|cpri_rx|cpri_rx_tx_rx|gige_rx|gige_1588_rx|basic_rm_enable_rx|basic_rm_disable_rx|disabled_prot_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcie_g1_capable_rx|pcie_g2_capable_rx|pcie_g3_capable_rx|gige_rx|teng_baser_rx|teng_basekr_krfec_rx|fortyg_basekr_krfec_rx|cpri_8b10b_rx|interlaken_rx|sfis_rx|teng_sdi_rx|gige_1588_rx|teng_1588_baser_rx|teng_1588_basekr_krfec_rx|basic_8gpcs_rm_enable_rx|basic_8gpcs_rm_disable_rx|basic_10gpcs_rx|basic_10gpcs_krfec_rx|pcs_direct_rx|prp_rx|prp_krfec_rx|prbs_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx = "teng_mode_rx", // teng_mode_rx|non_teng_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_basekr_mode_rx|fortyg_basekr_mode_rx|teng_1588_basekr_mode_rx|basic_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|eightg_and_g3_pld_fifo_mode_rx|eightg_and_g3_reg_mode_rx|eightg_and_g3_reg_mode_hip_rx|teng_pld_fifo_mode_rx|teng_reg_mode_rx|teng_and_krfec_pld_fifo_mode_rx|teng_and_krfec_reg_mode_rx|pcs_direct_reg_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_block_sel = "pcs_direct", // eightg|teng|pcs_direct
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_rx_clk|pma_rx_clk_user
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_sel = "pld_rx_clk", // pld_rx_clk|pcs_rx_clk
		parameter hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en = "hip_rx_enable", // hip_rx_enable|hip_rx_disable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_rx_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_tx_pcs_pma_interface
		parameter hssi_tx_pcs_pma_interface_bypass_pma_txelecidle = "false", // false|true
		parameter hssi_tx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pcs_pma_interface_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx = "other_prot_mode", // pipe_g12|pipe_g3|other_prot_mode
		parameter hssi_tx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_tx_pcs_pma_interface_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_tx_pcs_pma_interface_pmagate_en = "pmagate_dis", // pmagate_dis|pmagate_en
		parameter hssi_tx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_tx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_tx_pcs_pma_interface_prbs_gen_pat = "prbs_gen_dis", // prbs_gen_dis|prbs_31|prbs_23|prbs_15|prbs_9|prbs_7
		parameter hssi_tx_pcs_pma_interface_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_tx_pcs_pma_interface_sq_wave_num = "sq_wave_4", // sq_wave_1|sq_wave_4|sq_wave_8|sq_wave_6|sq_wave_default
		parameter hssi_tx_pcs_pma_interface_sqwgen_clken = "sqwgen_clk_dis", // sqwgen_clk_dis|sqwgen_clk_en
		parameter hssi_tx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion = "tx_dyn_polinv_dis", // tx_dyn_polinv_dis|tx_dyn_polinv_en
		parameter hssi_tx_pcs_pma_interface_tx_pma_data_sel = "pld_dir", // pld_dir|pcie_gen3|eight_g_pcs|ten_g_pcs|prbs_pat|sq_wave_pat|block_sel_default|registered_uhsif_dat|directed_uhsif_dat
		parameter hssi_tx_pcs_pma_interface_tx_static_polarity_inversion = "tx_stat_polinv_dis", // tx_stat_polinv_dis|tx_stat_polinv_en
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock = "uhsif_filt_stepsz_b4lock_4", // uhsif_filt_stepsz_b4lock_2|uhsif_filt_stepsz_b4lock_4|uhsif_filt_stepsz_b4lock_6|uhsif_filt_stepsz_b4lock_8
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value = 4'b1011,
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock = "uhsif_filt_cntthr_b4lock_16", // uhsif_filt_cntthr_b4lock_8|uhsif_filt_cntthr_b4lock_16|uhsif_filt_cntthr_b4lock_24|uhsif_filt_cntthr_b4lock_32
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period = "uhsif_dcn_test_period_4", // uhsif_dcn_test_period_4|uhsif_dcn_test_period_8|uhsif_dcn_test_period_12|uhsif_dcn_test_period_16
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable = "uhsif_dcn_test_mode_disable", // uhsif_dcn_test_mode_enable|uhsif_dcn_test_mode_disable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh = "uhsif_dzt_cnt_thr_4", // uhsif_dzt_cnt_thr_2|uhsif_dzt_cnt_thr_4|uhsif_dzt_cnt_thr_6|uhsif_dzt_cnt_thr_8
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable = "uhsif_dzt_enable", // uhsif_dzt_disable|uhsif_dzt_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window = "uhsif_dzt_obr_win_32", // uhsif_dzt_obr_win_16|uhsif_dzt_obr_win_32|uhsif_dzt_obr_win_48|uhsif_dzt_obr_win_64
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size = "uhsif_dzt_skipsz_8", // uhsif_dzt_skipsz_4|uhsif_dzt_skipsz_8|uhsif_dzt_skipsz_12|uhsif_dzt_skipsz_16
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel = "uhsif_index_internal", // uhsif_index_internal|uhsif_index_cram
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin = "uhsif_dcn_margin_4", // uhsif_dcn_margin_2|uhsif_dcn_margin_3|uhsif_dcn_margin_4|uhsif_dcn_margin_5
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value = 8'b10000000,
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control = "uhsif_dft_dz_det_val_0", // uhsif_dft_dz_det_val_0|uhsif_dft_dz_det_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control = "uhsif_dft_up_val_0", // uhsif_dft_up_val_0|uhsif_dft_up_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_enable = "uhsif_disable", // uhsif_disable|uhsif_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock = "uhsif_lkd_segsz_aflock_2048", // uhsif_lkd_segsz_aflock_512|uhsif_lkd_segsz_aflock_1024|uhsif_lkd_segsz_aflock_2048|uhsif_lkd_segsz_aflock_4096
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock = "uhsif_lkd_segsz_b4lock_32", // uhsif_lkd_segsz_b4lock_16|uhsif_lkd_segsz_b4lock_32|uhsif_lkd_segsz_b4lock_64|uhsif_lkd_segsz_b4lock_128
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value = 4'b11,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value = 4'b11,
		
		// parameters for twentynm_hssi_tx_pld_pcs_interface
		parameter hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx = "enable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx = "pma_64b_tx", // pma_32b_tx|pma_40b_tx|pma_64b_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_baser_mode_tx|interlaken_mode_tx|sfis_mode_tx|teng_sdi_mode_tx|basic_mode_tx|test_prp_mode_tx|test_prp_krfec_mode_tx|teng_1588_mode_tx|teng_baser_krfec_mode_tx|teng_1588_krfec_mode_tx|basic_krfec_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx = "disabled_prot_mode_tx", // pipe_g1_tx|pipe_g2_tx|pipe_g3_tx|cpri_tx|cpri_rx_tx_tx|gige_tx|gige_1588_tx|basic_tx|disabled_prot_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcie_g1_capable_tx|pcie_g2_capable_tx|pcie_g3_capable_tx|gige_tx|teng_baser_tx|teng_basekr_krfec_tx|fortyg_basekr_krfec_tx|cpri_8b10b_tx|interlaken_tx|sfis_tx|teng_sdi_tx|gige_1588_tx|teng_1588_baser_tx|teng_1588_basekr_krfec_tx|basic_8gpcs_tx|basic_10gpcs_tx|basic_10gpcs_krfec_tx|pcs_direct_tx|uhsif_tx|prp_tx|prp_krfec_tx|prbs_tx|sqwave_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx = "teng_mode_tx", // teng_mode_tx|non_teng_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_basekr_mode_tx|fortyg_basekr_mode_tx|teng_1588_basekr_mode_tx|basic_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|eightg_and_g3_pld_fifo_mode_tx|eightg_and_g3_reg_mode_tx|eightg_and_g3_reg_mode_hip_tx|eightg_and_g3_fastreg_mode_tx|teng_pld_fifo_mode_tx|teng_reg_mode_tx|teng_fastreg_mode_tx|teng_and_krfec_pld_fifo_mode_tx|teng_and_krfec_reg_mode_tx|teng_and_krfec_fastreg_mode_tx|pcs_direct_fastreg_mode_tx|uhsif_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_tx_clk|pma_tx_clk_user
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_source = "teng", // eightg|teng|pma_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_data_source = "hip_disable", // hip_disable|hip_enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en = "delay1_clk_disable", // delay1_clk_enable|delay1_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel = "pld_tx_clk", // pld_tx_clk|pcs_tx_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl = "delay1_path0", // delay1_path0|delay1_path1|delay1_path2|delay1_path3|delay1_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel = "one_ff_delay", // one_ff_delay|two_ff_delay
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en = "delay2_clk_disable", // delay2_clk_enable|delay2_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl = "delay2_path0", // delay2_path0|delay2_path1|delay2_path2|delay2_path3|delay2_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_tx_pld_pcs_interface_reconfig_settings = "{}" // 
	//PARAM_LIST_END
	)
	(
	//PORT_LIST_START
		input wire	[8:0]	in_avmmaddress,
		input wire		in_avmmclk,
		input wire		in_avmmread,
		input wire		in_avmmrstn,
		input wire		in_avmmwrite,
		input wire	[7:0]	in_avmmwritedata,
		input wire	[4:0]	in_bond_pcs10g_in_bot,
		input wire	[4:0]	in_bond_pcs10g_in_top,
		input wire	[12:0]	in_bond_pcs8g_in_bot,
		input wire	[12:0]	in_bond_pcs8g_in_top,
		input wire	[11:0]	in_bond_pmaif_in_bot,
		input wire	[11:0]	in_bond_pmaif_in_top,
		input wire	[63:0]	in_hip_tx_data,
		input wire		in_iocsr_clk,
		input wire	[5:0]	in_iocsr_config,
		input wire		in_iocsr_rdy,
		input wire		in_iocsr_rdy_dly,
		input wire		in_pld_10g_krfec_rx_clr_errblk_cnt,
		input wire		in_pld_10g_krfec_rx_pld_rst_n,
		input wire		in_pld_10g_krfec_tx_pld_rst_n,
		input wire		in_pld_10g_rx_align_clr,
		input wire		in_pld_10g_rx_clr_ber_count,
		input wire		in_pld_10g_rx_rd_en,
		input wire	[6:0]	in_pld_10g_tx_bitslip,
		input wire		in_pld_10g_tx_burst_en,
		input wire		in_pld_10g_tx_data_valid,
		input wire	[1:0]	in_pld_10g_tx_diag_status,
		input wire		in_pld_10g_tx_wordslip,
		input wire		in_pld_8g_a1a2_size,
		input wire		in_pld_8g_bitloc_rev_en,
		input wire		in_pld_8g_byte_rev_en,
		input wire	[2:0]	in_pld_8g_eidleinfersel,
		input wire		in_pld_8g_encdt,
		input wire		in_pld_8g_g3_rx_pld_rst_n,
		input wire		in_pld_8g_g3_tx_pld_rst_n,
		input wire		in_pld_8g_rddisable_tx,
		input wire		in_pld_8g_rdenable_rx,
		input wire		in_pld_8g_refclk_dig2,
		input wire		in_pld_8g_rxpolarity,
		input wire	[4:0]	in_pld_8g_tx_boundary_sel,
		input wire		in_pld_8g_wrdisable_rx,
		input wire		in_pld_8g_wrenable_tx,
		input wire		in_pld_atpg_los_en_n,
		input wire		in_pld_bitslip,
		input wire	[17:0]	in_pld_g3_current_coeff,
		input wire	[2:0]	in_pld_g3_current_rxpreset,
		input wire		in_pld_ltr,
		input wire		in_pld_mem_krfec_atpg_rst_n,
		input wire		in_pld_partial_reconfig,
		input wire		in_pld_pcs_refclk_dig,
		input wire		in_pld_pma_adapt_start,
		input wire		in_pld_pma_csr_test_dis,
		input wire		in_pld_pma_early_eios,
		input wire	[5:0]	in_pld_pma_eye_monitor,
		input wire		in_pld_pma_ltd_b,
		input wire		in_pld_pma_nrpi_freeze,
		input wire	[1:0]	in_pld_pma_pcie_switch,
		input wire		in_pld_pma_ppm_lock,
		input wire	[4:0]	in_pld_pma_reserved_out,
		input wire		in_pld_pma_rs_lpbk_b,
		input wire		in_pld_pma_rx_qpi_pullup,
		input wire		in_pld_pma_rxpma_rstb,
		input wire		in_pld_pma_tx_bitslip,
		input wire		in_pld_pma_tx_bonding_rstb,
		input wire		in_pld_pma_tx_qpi_pulldn,
		input wire		in_pld_pma_tx_qpi_pullup,
		input wire		in_pld_pma_txdetectrx,
		input wire		in_pld_pma_txpma_rstb,
		input wire		in_pld_pmaif_rx_pld_rst_n,
		input wire		in_pld_pmaif_rxclkslip,
		input wire		in_pld_pmaif_tx_pld_rst_n,
		input wire		in_pld_polinv_rx,
		input wire		in_pld_polinv_tx,
		input wire	[1:0]	in_pld_rate,
		input wire	[9:0]	in_pld_reserved_in,
		input wire		in_pld_rx_clk,
		input wire		in_pld_rx_prbs_err_clr,
		input wire		in_pld_scan_mode_n,
		input wire		in_pld_scan_shift_n,
		input wire		in_pld_syncsm_en,
		input wire		in_pld_tx_clk,
		input wire	[17:0]	in_pld_tx_control,
		input wire	[127:0]	in_pld_tx_data,
		input wire		in_pld_txelecidle,
		input wire		in_pld_uhsif_tx_clk,
		input wire		in_pma_adapt_done,
		input wire		in_pma_clklow,
		input wire		in_pma_fref,
		input wire		in_pma_hclk,
		input wire	[1:0]	in_pma_pcie_sw_done,
		input wire		in_pma_pfdmode_lock,
		input wire	[4:0]	in_pma_reserved_in,
		input wire		in_pma_rx_clkdiv_user,
		input wire		in_pma_rx_detect_valid,
		input wire		in_pma_rx_found,
		input wire		in_pma_rx_pma_clk,
		input wire	[63:0]	in_pma_rx_pma_data,
		input wire		in_pma_rx_signal_ok,
		input wire		in_pma_rxpll_lock,
		input wire		in_pma_signal_det,
		input wire	[7:0]	in_pma_testbus,
		input wire		in_pma_tx_clkdiv_user,
		input wire		in_pma_tx_pma_clk,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen1_2,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen3,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pld_pcs_interface,
		output wire		out_blockselect_hssi_10g_rx_pcs,
		output wire		out_blockselect_hssi_10g_tx_pcs,
		output wire		out_blockselect_hssi_8g_rx_pcs,
		output wire		out_blockselect_hssi_8g_tx_pcs,
		output wire		out_blockselect_hssi_common_pcs_pma_interface,
		output wire		out_blockselect_hssi_common_pld_pcs_interface,
		output wire		out_blockselect_hssi_fifo_rx_pcs,
		output wire		out_blockselect_hssi_fifo_tx_pcs,
		output wire		out_blockselect_hssi_gen3_rx_pcs,
		output wire		out_blockselect_hssi_gen3_tx_pcs,
		output wire		out_blockselect_hssi_krfec_rx_pcs,
		output wire		out_blockselect_hssi_krfec_tx_pcs,
		output wire		out_blockselect_hssi_pipe_gen1_2,
		output wire		out_blockselect_hssi_pipe_gen3,
		output wire		out_blockselect_hssi_rx_pcs_pma_interface,
		output wire		out_blockselect_hssi_rx_pld_pcs_interface,
		output wire		out_blockselect_hssi_tx_pcs_pma_interface,
		output wire		out_blockselect_hssi_tx_pld_pcs_interface,
		output wire	[4:0]	out_bond_pcs10g_out_bot,
		output wire	[4:0]	out_bond_pcs10g_out_top,
		output wire	[12:0]	out_bond_pcs8g_out_bot,
		output wire	[12:0]	out_bond_pcs8g_out_top,
		output wire	[11:0]	out_bond_pmaif_out_bot,
		output wire	[11:0]	out_bond_pmaif_out_top,
		output wire	[2:0]	out_hip_clk_out,
		output wire	[7:0]	out_hip_ctrl_out,
		output wire		out_hip_iocsr_rdy,
		output wire		out_hip_iocsr_rdy_dly,
		output wire		out_hip_nfrzdrv,
		output wire		out_hip_npor,
		output wire	[50:0]	out_hip_rx_data,
		output wire		out_hip_usermode,
		output wire		out_pld_10g_krfec_rx_blk_lock,
		output wire	[1:0]	out_pld_10g_krfec_rx_diag_data_status,
		output wire		out_pld_10g_krfec_rx_frame,
		output wire		out_pld_10g_krfec_tx_frame,
		output wire		out_pld_10g_rx_align_val,
		output wire		out_pld_10g_rx_crc32_err,
		output wire		out_pld_10g_rx_data_valid,
		output wire		out_pld_10g_rx_empty,
		output wire		out_pld_10g_rx_fifo_del,
		output wire		out_pld_10g_rx_fifo_insert,
		output wire	[4:0]	out_pld_10g_rx_fifo_num,
		output wire		out_pld_10g_rx_frame_lock,
		output wire		out_pld_10g_rx_hi_ber,
		output wire		out_pld_10g_rx_oflw_err,
		output wire		out_pld_10g_rx_pempty,
		output wire		out_pld_10g_rx_pfull,
		output wire		out_pld_10g_tx_burst_en_exe,
		output wire		out_pld_10g_tx_empty,
		output wire	[3:0]	out_pld_10g_tx_fifo_num,
		output wire		out_pld_10g_tx_full,
		output wire		out_pld_10g_tx_pempty,
		output wire		out_pld_10g_tx_pfull,
		output wire		out_pld_10g_tx_wordslip_exe,
		output wire	[3:0]	out_pld_8g_a1a2_k1k2_flag,
		output wire		out_pld_8g_empty_rmf,
		output wire		out_pld_8g_empty_rx,
		output wire		out_pld_8g_empty_tx,
		output wire		out_pld_8g_full_rmf,
		output wire		out_pld_8g_full_rx,
		output wire		out_pld_8g_full_tx,
		output wire		out_pld_8g_rxelecidle,
		output wire		out_pld_8g_signal_detect_out,
		output wire	[4:0]	out_pld_8g_wa_boundary,
		output wire		out_pld_krfec_tx_alignment,
		output wire		out_pld_pcs_rx_clk_out,
		output wire		out_pld_pcs_tx_clk_out,
		output wire		out_pld_pma_adapt_done,
		output wire		out_pld_pma_clkdiv_rx_user,
		output wire		out_pld_pma_clkdiv_tx_user,
		output wire		out_pld_pma_clklow,
		output wire		out_pld_pma_fref,
		output wire		out_pld_pma_hclk,
		output wire	[1:0]	out_pld_pma_pcie_sw_done,
		output wire		out_pld_pma_pfdmode_lock,
		output wire	[4:0]	out_pld_pma_reserved_in,
		output wire		out_pld_pma_rx_clk_out,
		output wire		out_pld_pma_rx_detect_valid,
		output wire		out_pld_pma_rx_found,
		output wire		out_pld_pma_rxpll_lock,
		output wire		out_pld_pma_signal_ok,
		output wire	[7:0]	out_pld_pma_testbus,
		output wire		out_pld_pma_tx_clk_out,
		output wire		out_pld_pmaif_mask_tx_pll,
		output wire	[9:0]	out_pld_reserved_out,
		output wire	[19:0]	out_pld_rx_control,
		output wire	[127:0]	out_pld_rx_data,
		output wire		out_pld_rx_prbs_done,
		output wire		out_pld_rx_prbs_err,
		output wire	[19:0]	out_pld_test_data,
		output wire		out_pld_uhsif_lock,
		output wire		out_pld_uhsif_tx_clk_out,
		output wire		out_pma_adapt_start,
		output wire		out_pma_atpg_los_en_n,
		output wire		out_pma_csr_test_dis,
		output wire	[17:0]	out_pma_current_coeff,
		output wire	[2:0]	out_pma_current_rxpreset,
		output wire		out_pma_early_eios,
		output wire	[5:0]	out_pma_eye_monitor,
		output wire	[1:0]	out_pma_interface_select,
		output wire		out_pma_ltd_b,
		output wire		out_pma_ltr,
		output wire		out_pma_nfrzdrv,
		output wire		out_pma_nrpi_freeze,
		output wire	[1:0]	out_pma_pcie_switch,
		output wire		out_pma_ppm_lock,
		output wire	[4:0]	out_pma_reserved_out,
		output wire		out_pma_rs_lpbk_b,
		output wire		out_pma_rx_clkslip,
		output wire		out_pma_rx_qpi_pullup,
		output wire		out_pma_rxpma_rstb,
		output wire		out_pma_scan_mode_n,
		output wire		out_pma_scan_shift_n,
		output wire		out_pma_tx_bitslip,
		output wire		out_pma_tx_bonding_rstb,
		output wire		out_pma_tx_elec_idle,
		output wire	[63:0]	out_pma_tx_pma_data,
		output wire		out_pma_tx_qpi_pulldn,
		output wire		out_pma_tx_qpi_pullup,
		output wire		out_pma_tx_txdetectrx,
		output wire		out_pma_txpma_rstb
	//PORT_LIST_END
	);
	//wire declarations
	
	// wires for module twentynm_hssi_fifo_tx_pcs
	wire	[7:0]	w_hssi_fifo_tx_pcs_avmmreaddata;
	wire		w_hssi_fifo_tx_pcs_blockselect;
	wire	[72:0]	w_hssi_fifo_tx_pcs_data_out_10g;
	wire	[63:0]	w_hssi_fifo_tx_pcs_data_out_8g_phase_comp;
	
	// wires for module twentynm_hssi_gen3_rx_pcs
	wire	[7:0]	w_hssi_gen3_rx_pcs_avmmreaddata;
	wire		w_hssi_gen3_rx_pcs_blk_algnd_int;
	wire		w_hssi_gen3_rx_pcs_blk_start;
	wire		w_hssi_gen3_rx_pcs_blockselect;
	wire		w_hssi_gen3_rx_pcs_clkcomp_delete_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_insert_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_overfl_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_undfl_int;
	wire	[31:0]	w_hssi_gen3_rx_pcs_data_out;
	wire		w_hssi_gen3_rx_pcs_data_valid;
	wire		w_hssi_gen3_rx_pcs_ei_det_int;
	wire		w_hssi_gen3_rx_pcs_ei_partial_det_int;
	wire		w_hssi_gen3_rx_pcs_err_decode_int;
	wire		w_hssi_gen3_rx_pcs_i_det_int;
	wire		w_hssi_gen3_rx_pcs_lpbk_blk_start;
	wire	[33:0]	w_hssi_gen3_rx_pcs_lpbk_data;
	wire		w_hssi_gen3_rx_pcs_lpbk_data_valid;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk;
	wire	[39:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n;
	wire		w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int;
	wire	[19:0]	w_hssi_gen3_rx_pcs_rx_test_out;
	wire	[1:0]	w_hssi_gen3_rx_pcs_sync_hdr;
	
	// wires for module twentynm_hssi_krfec_tx_pcs
	wire	[7:0]	w_hssi_krfec_tx_pcs_avmmreaddata;
	wire		w_hssi_krfec_tx_pcs_blockselect;
	wire		w_hssi_krfec_tx_pcs_tx_alignment;
	wire	[63:0]	w_hssi_krfec_tx_pcs_tx_data_out;
	wire		w_hssi_krfec_tx_pcs_tx_frame;
	wire	[19:0]	w_hssi_krfec_tx_pcs_tx_test_data;
	
	// wires for module twentynm_hssi_krfec_rx_pcs
	wire	[7:0]	w_hssi_krfec_rx_pcs_avmmreaddata;
	wire		w_hssi_krfec_rx_pcs_blockselect;
	wire		w_hssi_krfec_rx_pcs_rx_block_lock;
	wire	[9:0]	w_hssi_krfec_rx_pcs_rx_control_out;
	wire	[63:0]	w_hssi_krfec_rx_pcs_rx_data_out;
	wire	[1:0]	w_hssi_krfec_rx_pcs_rx_data_status;
	wire		w_hssi_krfec_rx_pcs_rx_data_valid_out;
	wire		w_hssi_krfec_rx_pcs_rx_frame;
	wire		w_hssi_krfec_rx_pcs_rx_signal_ok_out;
	
	// wires for module twentynm_hssi_rx_pld_pcs_interface
	wire	[7:0]	w_hssi_rx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_rx_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_hip_rx_ctrl;
	wire	[50:0]	w_hssi_rx_pld_pcs_interface_hip_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
	wire	[3:0]	w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary;
	wire		w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_pld_rx_control;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_pld_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
	
	// wires for module twentynm_hssi_common_pld_pcs_interface
	wire	[7:0]	w_hssi_common_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_common_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_hip_cmn_clk;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_hip_cmn_ctrl;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
	wire		w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_hip_npor;
	wire		w_hssi_common_pld_pcs_interface_hip_usermode;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n;
	wire	[17:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel;
	wire		w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_clklow;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_fref;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_hclk;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_pld_pma_reserved_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
	wire	[7:0]	w_hssi_common_pld_pcs_interface_pld_pma_testbus;
	wire		w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
	wire	[9:0]	w_hssi_common_pld_pcs_interface_pld_reserved_out;
	wire	[19:0]	w_hssi_common_pld_pcs_interface_pld_test_data;
	wire		w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
	wire		w_hssi_common_pld_pcs_interface_scan_mode_n;
	
	// wires for module twentynm_hssi_10g_rx_pcs
	wire	[7:0]	w_hssi_10g_rx_pcs_avmmreaddata;
	wire		w_hssi_10g_rx_pcs_blockselect;
	wire		w_hssi_10g_rx_pcs_rx_align_val;
	wire		w_hssi_10g_rx_pcs_rx_blk_lock;
	wire		w_hssi_10g_rx_pcs_rx_clk_out;
	wire		w_hssi_10g_rx_pcs_rx_clk_out_pld_if;
	wire	[19:0]	w_hssi_10g_rx_pcs_rx_control;
	wire		w_hssi_10g_rx_pcs_rx_crc32_err;
	wire	[127:0]	w_hssi_10g_rx_pcs_rx_data;
	wire		w_hssi_10g_rx_pcs_rx_data_valid;
	wire		w_hssi_10g_rx_pcs_rx_dft_clk_out;
	wire	[1:0]	w_hssi_10g_rx_pcs_rx_diag_status;
	wire		w_hssi_10g_rx_pcs_rx_empty;
	wire		w_hssi_10g_rx_pcs_rx_fec_clk;
	wire		w_hssi_10g_rx_pcs_rx_fifo_del;
	wire		w_hssi_10g_rx_pcs_rx_fifo_insert;
	wire	[4:0]	w_hssi_10g_rx_pcs_rx_fifo_num;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_clk;
	wire	[73:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_data;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_en;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_ptr;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_frame_lock;
	wire		w_hssi_10g_rx_pcs_rx_hi_ber;
	wire		w_hssi_10g_rx_pcs_rx_master_clk;
	wire		w_hssi_10g_rx_pcs_rx_master_clk_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_oflw_err;
	wire		w_hssi_10g_rx_pcs_rx_pempty;
	wire		w_hssi_10g_rx_pcs_rx_pfull;
	wire		w_hssi_10g_rx_pcs_rx_random_err;
	wire		w_hssi_10g_rx_pcs_rx_rx_frame;
	
	// wires for module twentynm_hssi_tx_pld_pcs_interface
	wire	[7:0]	w_hssi_tx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_tx_pld_pcs_interface_blockselect;
	wire		w_hssi_tx_pld_pcs_interface_hip_tx_clk;
	wire	[6:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en;
	wire	[17:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control;
	wire	[8:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg;
	wire	[127:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start;
	wire	[4:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle;
	wire	[2:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
	wire		w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
	
	// wires for module twentynm_hssi_tx_pcs_pma_interface
	wire	[7:0]	w_hssi_tx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_tx_pcs_pma_interface_blockselect;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out;
	wire	[4:0]	w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk;
	wire		w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_pma_tx_pma_data;
	wire		w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_1;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_2;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_3;
	
	// wires for module twentynm_hssi_rx_pcs_pma_interface
	wire	[7:0]	w_hssi_rx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_rx_pcs_pma_interface_blockselect;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni;
	wire	[31:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok;
	wire		w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk;
	wire	[5:0]	w_hssi_rx_pcs_pma_interface_pma_eye_monitor;
	wire		w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
	wire		w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test;
	
	// wires for module twentynm_hssi_10g_tx_pcs
	wire	[7:0]	w_hssi_10g_tx_pcs_avmmreaddata;
	wire		w_hssi_10g_tx_pcs_blockselect;
	wire		w_hssi_10g_tx_pcs_distdwn_out_dv;
	wire		w_hssi_10g_tx_pcs_distdwn_out_rden;
	wire		w_hssi_10g_tx_pcs_distdwn_out_wren;
	wire		w_hssi_10g_tx_pcs_distup_out_dv;
	wire		w_hssi_10g_tx_pcs_distup_out_rden;
	wire		w_hssi_10g_tx_pcs_distup_out_wren;
	wire		w_hssi_10g_tx_pcs_tx_burst_en_exe;
	wire		w_hssi_10g_tx_pcs_tx_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pma_if;
	wire	[8:0]	w_hssi_10g_tx_pcs_tx_control_out_krfec;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_data_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_data_valid_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_dft_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_empty;
	wire		w_hssi_10g_tx_pcs_tx_fec_clk;
	wire	[3:0]	w_hssi_10g_tx_pcs_tx_fifo_num;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_rd_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_clk;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_en;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_frame;
	wire		w_hssi_10g_tx_pcs_tx_full;
	wire		w_hssi_10g_tx_pcs_tx_master_clk;
	wire		w_hssi_10g_tx_pcs_tx_master_clk_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_pempty;
	wire		w_hssi_10g_tx_pcs_tx_pfull;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_data;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_gating_val;
	wire	[19:0]	w_hssi_10g_tx_pcs_tx_test_data;
	wire		w_hssi_10g_tx_pcs_tx_wordslip_exe;
	
	// wires for module twentynm_hssi_8g_tx_pcs
	wire	[7:0]	w_hssi_8g_tx_pcs_avmmreaddata;
	wire		w_hssi_8g_tx_pcs_blockselect;
	wire		w_hssi_8g_tx_pcs_clk_out;
	wire		w_hssi_8g_tx_pcs_clk_out_gen3;
	wire	[19:0]	w_hssi_8g_tx_pcs_dataout;
	wire		w_hssi_8g_tx_pcs_dyn_clk_switch_n;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn;
	wire		w_hssi_8g_tx_pcs_g3_tx_pma_rstn;
	wire	[2:0]	w_hssi_8g_tx_pcs_non_gray_eidleinfersel;
	wire		w_hssi_8g_tx_pcs_ph_fifo_overflow;
	wire		w_hssi_8g_tx_pcs_ph_fifo_underflow;
	wire		w_hssi_8g_tx_pcs_phfifo_txdeemph;
	wire	[2:0]	w_hssi_8g_tx_pcs_phfifo_txmargin;
	wire		w_hssi_8g_tx_pcs_phfifo_txswing;
	wire		w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out;
	wire	[1:0]	w_hssi_8g_tx_pcs_pipe_power_down_out;
	wire		w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3;
	wire		w_hssi_8g_tx_pcs_pmaif_asn_rstn;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_refclk_b;
	wire		w_hssi_8g_tx_pcs_refclk_b_reset;
	wire		w_hssi_8g_tx_pcs_rxpolarity_int;
	wire		w_hssi_8g_tx_pcs_soft_reset_wclk1_n;
	wire		w_hssi_8g_tx_pcs_sw_fifo_wr_clk;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_blk_start_out;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_ctrlplane_testbus;
	wire	[31:0]	w_hssi_8g_tx_pcs_tx_data_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_data_valid_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_datak_out;
	wire		w_hssi_8g_tx_pcs_tx_detect_rxloopback_int;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_tx_pipe_clk;
	wire		w_hssi_8g_tx_pcs_tx_pipe_electidle;
	wire		w_hssi_8g_tx_pcs_tx_pipe_soft_reset;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_sync_hdr_out;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_testbus;
	wire		w_hssi_8g_tx_pcs_txcompliance_out;
	wire		w_hssi_8g_tx_pcs_txelecidle_out;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk;
	wire	[63:0]	w_hssi_8g_tx_pcs_wr_data_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_en_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo;
	
	// wires for module twentynm_hssi_pipe_gen3
	wire	[7:0]	w_hssi_pipe_gen3_avmmreaddata;
	wire		w_hssi_pipe_gen3_blockselect;
	wire		w_hssi_pipe_gen3_gen3_clk_sel;
	wire		w_hssi_pipe_gen3_pcs_rst;
	wire		w_hssi_pipe_gen3_phystatus;
	wire	[17:0]	w_hssi_pipe_gen3_pma_current_coeff;
	wire	[2:0]	w_hssi_pipe_gen3_pma_current_rxpreset;
	wire		w_hssi_pipe_gen3_pma_tx_elec_idle;
	wire		w_hssi_pipe_gen3_pma_txdetectrx;
	wire		w_hssi_pipe_gen3_rev_lpbk_8gpcs_out;
	wire		w_hssi_pipe_gen3_rev_lpbk_int;
	wire	[3:0]	w_hssi_pipe_gen3_rx_blk_start;
	wire	[1:0]	w_hssi_pipe_gen3_rx_sync_hdr;
	wire	[63:0]	w_hssi_pipe_gen3_rxd_8gpcs_out;
	wire	[3:0]	w_hssi_pipe_gen3_rxdataskip;
	wire		w_hssi_pipe_gen3_rxelecidle;
	wire		w_hssi_pipe_gen3_rxpolarity_8gpcs_out;
	wire		w_hssi_pipe_gen3_rxpolarity_int;
	wire	[2:0]	w_hssi_pipe_gen3_rxstatus;
	wire		w_hssi_pipe_gen3_rxvalid;
	wire		w_hssi_pipe_gen3_shutdown_clk;
	wire	[19:0]	w_hssi_pipe_gen3_test_out;
	wire		w_hssi_pipe_gen3_tx_blk_start_int;
	wire	[1:0]	w_hssi_pipe_gen3_tx_sync_hdr_int;
	wire	[31:0]	w_hssi_pipe_gen3_txdata_int;
	wire	[3:0]	w_hssi_pipe_gen3_txdatak_int;
	wire		w_hssi_pipe_gen3_txdataskip_int;
	
	// wires for module twentynm_hssi_pipe_gen1_2
	wire	[7:0]	w_hssi_pipe_gen1_2_avmmreaddata;
	wire		w_hssi_pipe_gen1_2_blockselect;
	wire	[17:0]	w_hssi_pipe_gen1_2_current_coeff;
	wire		w_hssi_pipe_gen1_2_phystatus;
	wire		w_hssi_pipe_gen1_2_polarity_inversion_rx;
	wire		w_hssi_pipe_gen1_2_rev_loopbk;
	wire		w_hssi_pipe_gen1_2_rxelecidle;
	wire		w_hssi_pipe_gen1_2_rxelectricalidle_out;
	wire	[2:0]	w_hssi_pipe_gen1_2_rxstatus;
	wire		w_hssi_pipe_gen1_2_rxvalid;
	wire		w_hssi_pipe_gen1_2_tx_elec_idle_out;
	wire		w_hssi_pipe_gen1_2_txdetectrx;
	
	// wires for module twentynm_hssi_gen3_tx_pcs
	wire	[7:0]	w_hssi_gen3_tx_pcs_avmmreaddata;
	wire		w_hssi_gen3_tx_pcs_blockselect;
	wire	[31:0]	w_hssi_gen3_tx_pcs_data_out;
	wire	[35:0]	w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out;
	wire	[31:0]	w_hssi_gen3_tx_pcs_par_lpbk_out;
	wire	[19:0]	w_hssi_gen3_tx_pcs_tx_test_out;
	
	// wires for module twentynm_hssi_8g_rx_pcs
	wire	[3:0]	w_hssi_8g_rx_pcs_a1a2k1k2flag;
	wire	[7:0]	w_hssi_8g_rx_pcs_avmmreaddata;
	wire		w_hssi_8g_rx_pcs_blockselect;
	wire	[19:0]	w_hssi_8g_rx_pcs_chnl_test_bus_out;
	wire		w_hssi_8g_rx_pcs_clock_to_pld;
	wire	[63:0]	w_hssi_8g_rx_pcs_dataout;
	wire		w_hssi_8g_rx_pcs_dis_pc_byte;
	wire		w_hssi_8g_rx_pcs_eidle_detected;
	wire	[2:0]	w_hssi_8g_rx_pcs_eios_det_cdr_ctrl;
	wire		w_hssi_8g_rx_pcs_g3_rx_pma_rstn;
	wire		w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn;
	wire		w_hssi_8g_rx_pcs_gen2ngen1;
	wire	[19:0]	w_hssi_8g_rx_pcs_parallel_rev_loopback;
	wire		w_hssi_8g_rx_pcs_pc_fifo_empty;
	wire		w_hssi_8g_rx_pcs_pcfifofull;
	wire		w_hssi_8g_rx_pcs_phystatus;
	wire	[63:0]	w_hssi_8g_rx_pcs_pipe_data;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_up;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo;
	wire	[7:0]	w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rm_fifo_empty;
	wire		w_hssi_8g_rx_pcs_rm_fifo_full;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_blk_start;
	wire		w_hssi_8g_rx_pcs_rx_clk_out_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clkslip;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_data_valid;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rx_pipe_clk;
	wire		w_hssi_8g_rx_pcs_rx_pipe_soft_reset;
	wire		w_hssi_8g_rx_pcs_rx_pma_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_sync_hdr;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_up;
	wire	[2:0]	w_hssi_8g_rx_pcs_rxstatus;
	wire		w_hssi_8g_rx_pcs_rxvalid;
	wire		w_hssi_8g_rx_pcs_signal_detect_out;
	wire	[4:0]	w_hssi_8g_rx_pcs_word_align_boundary;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk;
	wire	[79:0]	w_hssi_8g_rx_pcs_wr_data_rx_phfifo;
	wire	[31:0]	w_hssi_8g_rx_pcs_wr_data_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo;
	
	// wires for module twentynm_hssi_fifo_rx_pcs
	wire	[7:0]	w_hssi_fifo_rx_pcs_avmmreaddata;
	wire		w_hssi_fifo_rx_pcs_blockselect;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out2_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out_8g_clock_comp;
	wire	[79:0]	w_hssi_fifo_rx_pcs_data_out_8g_phase_comp;
	wire	[39:0]	w_hssi_fifo_rx_pcs_data_out_gen3;
	
	// wires for module twentynm_hssi_common_pcs_pma_interface
	wire	[7:0]	w_hssi_common_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_common_pcs_pma_interface_blockselect;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in;
	wire	[19:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out;
	wire	[7:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus;
	wire		w_hssi_common_pcs_pma_interface_pma_adapt_start;
	wire		w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
	wire		w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
	wire	[17:0]	w_hssi_common_pcs_pma_interface_pma_current_coeff;
	wire	[2:0]	w_hssi_common_pcs_pma_interface_pma_current_rxpreset;
	wire		w_hssi_common_pcs_pma_interface_pma_early_eios;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_interface_select;
	wire		w_hssi_common_pcs_pma_interface_pma_ltd_b;
	wire		w_hssi_common_pcs_pma_interface_pma_ltr;
	wire		w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
	wire		w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_pcie_switch;
	wire		w_hssi_common_pcs_pma_interface_pma_ppm_lock;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_pma_reserved_out;
	wire		w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
	wire		w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up;
	
	
	generate
		
		//module instantiations
		
		// instantiating twentynm_hssi_10g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_rx_pcs
			twentynm_hssi_10g_rx_pcs #(
				.advanced_user_mode(hssi_10g_rx_pcs_advanced_user_mode),
				.align_del(hssi_10g_rx_pcs_align_del),
				.ber_bit_err_total_cnt(hssi_10g_rx_pcs_ber_bit_err_total_cnt),
				.ber_clken(hssi_10g_rx_pcs_ber_clken),
				.ber_xus_timer_window(hssi_10g_rx_pcs_ber_xus_timer_window),
				.bitslip_mode(hssi_10g_rx_pcs_bitslip_mode),
				.blksync_bitslip_type(hssi_10g_rx_pcs_blksync_bitslip_type),
				.blksync_bitslip_wait_cnt(hssi_10g_rx_pcs_blksync_bitslip_wait_cnt),
				.blksync_bitslip_wait_type(hssi_10g_rx_pcs_blksync_bitslip_wait_type),
				.blksync_bypass(hssi_10g_rx_pcs_blksync_bypass),
				.blksync_clken(hssi_10g_rx_pcs_blksync_clken),
				.blksync_enum_invalid_sh_cnt(hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt),
				.blksync_knum_sh_cnt_postlock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock),
				.blksync_knum_sh_cnt_prelock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock),
				.blksync_pipeln(hssi_10g_rx_pcs_blksync_pipeln),
				.clr_errblk_cnt_en(hssi_10g_rx_pcs_clr_errblk_cnt_en),
				.control_del(hssi_10g_rx_pcs_control_del),
				.crcchk_bypass(hssi_10g_rx_pcs_crcchk_bypass),
				.crcchk_clken(hssi_10g_rx_pcs_crcchk_clken),
				.crcchk_inv(hssi_10g_rx_pcs_crcchk_inv),
				.crcchk_pipeln(hssi_10g_rx_pcs_crcchk_pipeln),
				.crcflag_pipeln(hssi_10g_rx_pcs_crcflag_pipeln),
				.ctrl_bit_reverse(hssi_10g_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_10g_rx_pcs_data_bit_reverse),
				.dec64b66b_clken(hssi_10g_rx_pcs_dec64b66b_clken),
				.dec_64b66b_rxsm_bypass(hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass),
				.descrm_bypass(hssi_10g_rx_pcs_descrm_bypass),
				.descrm_clken(hssi_10g_rx_pcs_descrm_clken),
				.descrm_mode(hssi_10g_rx_pcs_descrm_mode),
				.descrm_pipeln(hssi_10g_rx_pcs_descrm_pipeln),
				.dft_clk_out_sel(hssi_10g_rx_pcs_dft_clk_out_sel),
				.dis_signal_ok(hssi_10g_rx_pcs_dis_signal_ok),
				.dispchk_bypass(hssi_10g_rx_pcs_dispchk_bypass),
				.empty_flag_type(hssi_10g_rx_pcs_empty_flag_type),
				.fast_path(hssi_10g_rx_pcs_fast_path),
				.fec_clken(hssi_10g_rx_pcs_fec_clken),
				.fec_enable(hssi_10g_rx_pcs_fec_enable),
				.fifo_double_read(hssi_10g_rx_pcs_fifo_double_read),
				.fifo_stop_rd(hssi_10g_rx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_rx_pcs_fifo_stop_wr),
				.force_align(hssi_10g_rx_pcs_force_align),
				.frmsync_bypass(hssi_10g_rx_pcs_frmsync_bypass),
				.frmsync_clken(hssi_10g_rx_pcs_frmsync_clken),
				.frmsync_enum_scrm(hssi_10g_rx_pcs_frmsync_enum_scrm),
				.frmsync_enum_sync(hssi_10g_rx_pcs_frmsync_enum_sync),
				.frmsync_flag_type(hssi_10g_rx_pcs_frmsync_flag_type),
				.frmsync_knum_sync(hssi_10g_rx_pcs_frmsync_knum_sync),
				.frmsync_mfrm_length(hssi_10g_rx_pcs_frmsync_mfrm_length),
				.frmsync_pipeln(hssi_10g_rx_pcs_frmsync_pipeln),
				.full_flag_type(hssi_10g_rx_pcs_full_flag_type),
				.gb_rx_idwidth(hssi_10g_rx_pcs_gb_rx_idwidth),
				.gb_rx_odwidth(hssi_10g_rx_pcs_gb_rx_odwidth),
				.gbexp_clken(hssi_10g_rx_pcs_gbexp_clken),
				.low_latency_en(hssi_10g_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_10g_rx_pcs_lpbk_mode),
				.master_clk_sel(hssi_10g_rx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_rx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_rx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_rx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_rx_pcs_pld_if_type),
				.prot_mode(hssi_10g_rx_pcs_prot_mode),
				.rand_clken(hssi_10g_rx_pcs_rand_clken),
				.rd_clk_sel(hssi_10g_rx_pcs_rd_clk_sel),
				.rdfifo_clken(hssi_10g_rx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_rx_pcs_reconfig_settings),
				.rx_fifo_write_ctrl(hssi_10g_rx_pcs_rx_fifo_write_ctrl),
				.rx_scrm_width(hssi_10g_rx_pcs_rx_scrm_width),
				.rx_sh_location(hssi_10g_rx_pcs_rx_sh_location),
				.rx_signal_ok_sel(hssi_10g_rx_pcs_rx_signal_ok_sel),
				.rx_sm_bypass(hssi_10g_rx_pcs_rx_sm_bypass),
				.rx_sm_hiber(hssi_10g_rx_pcs_rx_sm_hiber),
				.rx_sm_pipeln(hssi_10g_rx_pcs_rx_sm_pipeln),
				.rx_testbus_sel(hssi_10g_rx_pcs_rx_testbus_sel),
				.rx_true_b2b(hssi_10g_rx_pcs_rx_true_b2b),
				.rxfifo_empty(hssi_10g_rx_pcs_rxfifo_empty),
				.rxfifo_full(hssi_10g_rx_pcs_rxfifo_full),
				.rxfifo_mode(hssi_10g_rx_pcs_rxfifo_mode),
				.rxfifo_pempty(hssi_10g_rx_pcs_rxfifo_pempty),
				.rxfifo_pfull(hssi_10g_rx_pcs_rxfifo_pfull),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.stretch_num_stages(hssi_10g_rx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_rx_pcs_sup_mode),
				.test_mode(hssi_10g_rx_pcs_test_mode),
				.wrfifo_clken(hssi_10g_rx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_rx_pcs_blockselect),
				.rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.rx_control(w_hssi_10g_rx_pcs_rx_control),
				.rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.rx_data(w_hssi_10g_rx_pcs_rx_data),
				.rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.rx_diag_status(w_hssi_10g_rx_pcs_rx_diag_status),
				.rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.rx_fec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.rx_fifo_num(w_hssi_10g_rx_pcs_rx_fifo_num),
				.rx_fifo_rd_ptr(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr),
				.rx_fifo_rd_ptr2(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2),
				.rx_fifo_wr_clk(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.rx_fifo_wr_data(w_hssi_10g_rx_pcs_rx_fifo_wr_data),
				.rx_fifo_wr_en(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.rx_fifo_wr_ptr(w_hssi_10g_rx_pcs_rx_fifo_wr_ptr),
				.rx_fifo_wr_rst_n(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.rx_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_rx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_rx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.rx_control_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0]}),
				.rx_control_in_krfec({w_hssi_krfec_rx_pcs_rx_control_out[9], w_hssi_krfec_rx_pcs_rx_control_out[8], w_hssi_krfec_rx_pcs_rx_control_out[7], w_hssi_krfec_rx_pcs_rx_control_out[6], w_hssi_krfec_rx_pcs_rx_control_out[5], w_hssi_krfec_rx_pcs_rx_control_out[4], w_hssi_krfec_rx_pcs_rx_control_out[3], w_hssi_krfec_rx_pcs_rx_control_out[2], w_hssi_krfec_rx_pcs_rx_control_out[1], w_hssi_krfec_rx_pcs_rx_control_out[0]}),
				.rx_data_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0]}),
				.rx_data_in_krfec({w_hssi_krfec_rx_pcs_rx_data_out[63], w_hssi_krfec_rx_pcs_rx_data_out[62], w_hssi_krfec_rx_pcs_rx_data_out[61], w_hssi_krfec_rx_pcs_rx_data_out[60], w_hssi_krfec_rx_pcs_rx_data_out[59], w_hssi_krfec_rx_pcs_rx_data_out[58], w_hssi_krfec_rx_pcs_rx_data_out[57], w_hssi_krfec_rx_pcs_rx_data_out[56], w_hssi_krfec_rx_pcs_rx_data_out[55], w_hssi_krfec_rx_pcs_rx_data_out[54], w_hssi_krfec_rx_pcs_rx_data_out[53], w_hssi_krfec_rx_pcs_rx_data_out[52], w_hssi_krfec_rx_pcs_rx_data_out[51], w_hssi_krfec_rx_pcs_rx_data_out[50], w_hssi_krfec_rx_pcs_rx_data_out[49], w_hssi_krfec_rx_pcs_rx_data_out[48], w_hssi_krfec_rx_pcs_rx_data_out[47], w_hssi_krfec_rx_pcs_rx_data_out[46], w_hssi_krfec_rx_pcs_rx_data_out[45], w_hssi_krfec_rx_pcs_rx_data_out[44], w_hssi_krfec_rx_pcs_rx_data_out[43], w_hssi_krfec_rx_pcs_rx_data_out[42], w_hssi_krfec_rx_pcs_rx_data_out[41], w_hssi_krfec_rx_pcs_rx_data_out[40], w_hssi_krfec_rx_pcs_rx_data_out[39], w_hssi_krfec_rx_pcs_rx_data_out[38], w_hssi_krfec_rx_pcs_rx_data_out[37], w_hssi_krfec_rx_pcs_rx_data_out[36], w_hssi_krfec_rx_pcs_rx_data_out[35], w_hssi_krfec_rx_pcs_rx_data_out[34], w_hssi_krfec_rx_pcs_rx_data_out[33], w_hssi_krfec_rx_pcs_rx_data_out[32], w_hssi_krfec_rx_pcs_rx_data_out[31], w_hssi_krfec_rx_pcs_rx_data_out[30], w_hssi_krfec_rx_pcs_rx_data_out[29], w_hssi_krfec_rx_pcs_rx_data_out[28], w_hssi_krfec_rx_pcs_rx_data_out[27], w_hssi_krfec_rx_pcs_rx_data_out[26], w_hssi_krfec_rx_pcs_rx_data_out[25], w_hssi_krfec_rx_pcs_rx_data_out[24], w_hssi_krfec_rx_pcs_rx_data_out[23], w_hssi_krfec_rx_pcs_rx_data_out[22], w_hssi_krfec_rx_pcs_rx_data_out[21], w_hssi_krfec_rx_pcs_rx_data_out[20], w_hssi_krfec_rx_pcs_rx_data_out[19], w_hssi_krfec_rx_pcs_rx_data_out[18], w_hssi_krfec_rx_pcs_rx_data_out[17], w_hssi_krfec_rx_pcs_rx_data_out[16], w_hssi_krfec_rx_pcs_rx_data_out[15], w_hssi_krfec_rx_pcs_rx_data_out[14], w_hssi_krfec_rx_pcs_rx_data_out[13], w_hssi_krfec_rx_pcs_rx_data_out[12], w_hssi_krfec_rx_pcs_rx_data_out[11], w_hssi_krfec_rx_pcs_rx_data_out[10], w_hssi_krfec_rx_pcs_rx_data_out[9], w_hssi_krfec_rx_pcs_rx_data_out[8], w_hssi_krfec_rx_pcs_rx_data_out[7], w_hssi_krfec_rx_pcs_rx_data_out[6], w_hssi_krfec_rx_pcs_rx_data_out[5], w_hssi_krfec_rx_pcs_rx_data_out[4], w_hssi_krfec_rx_pcs_rx_data_out[3], w_hssi_krfec_rx_pcs_rx_data_out[2], w_hssi_krfec_rx_pcs_rx_data_out[1], w_hssi_krfec_rx_pcs_rx_data_out[0]}),
				.rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.rx_data_valid_in_krfec(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_10g[73], w_hssi_fifo_rx_pcs_data_out_10g[72], w_hssi_fifo_rx_pcs_data_out_10g[71], w_hssi_fifo_rx_pcs_data_out_10g[70], w_hssi_fifo_rx_pcs_data_out_10g[69], w_hssi_fifo_rx_pcs_data_out_10g[68], w_hssi_fifo_rx_pcs_data_out_10g[67], w_hssi_fifo_rx_pcs_data_out_10g[66], w_hssi_fifo_rx_pcs_data_out_10g[65], w_hssi_fifo_rx_pcs_data_out_10g[64], w_hssi_fifo_rx_pcs_data_out_10g[63], w_hssi_fifo_rx_pcs_data_out_10g[62], w_hssi_fifo_rx_pcs_data_out_10g[61], w_hssi_fifo_rx_pcs_data_out_10g[60], w_hssi_fifo_rx_pcs_data_out_10g[59], w_hssi_fifo_rx_pcs_data_out_10g[58], w_hssi_fifo_rx_pcs_data_out_10g[57], w_hssi_fifo_rx_pcs_data_out_10g[56], w_hssi_fifo_rx_pcs_data_out_10g[55], w_hssi_fifo_rx_pcs_data_out_10g[54], w_hssi_fifo_rx_pcs_data_out_10g[53], w_hssi_fifo_rx_pcs_data_out_10g[52], w_hssi_fifo_rx_pcs_data_out_10g[51], w_hssi_fifo_rx_pcs_data_out_10g[50], w_hssi_fifo_rx_pcs_data_out_10g[49], w_hssi_fifo_rx_pcs_data_out_10g[48], w_hssi_fifo_rx_pcs_data_out_10g[47], w_hssi_fifo_rx_pcs_data_out_10g[46], w_hssi_fifo_rx_pcs_data_out_10g[45], w_hssi_fifo_rx_pcs_data_out_10g[44], w_hssi_fifo_rx_pcs_data_out_10g[43], w_hssi_fifo_rx_pcs_data_out_10g[42], w_hssi_fifo_rx_pcs_data_out_10g[41], w_hssi_fifo_rx_pcs_data_out_10g[40], w_hssi_fifo_rx_pcs_data_out_10g[39], w_hssi_fifo_rx_pcs_data_out_10g[38], w_hssi_fifo_rx_pcs_data_out_10g[37], w_hssi_fifo_rx_pcs_data_out_10g[36], w_hssi_fifo_rx_pcs_data_out_10g[35], w_hssi_fifo_rx_pcs_data_out_10g[34], w_hssi_fifo_rx_pcs_data_out_10g[33], w_hssi_fifo_rx_pcs_data_out_10g[32], w_hssi_fifo_rx_pcs_data_out_10g[31], w_hssi_fifo_rx_pcs_data_out_10g[30], w_hssi_fifo_rx_pcs_data_out_10g[29], w_hssi_fifo_rx_pcs_data_out_10g[28], w_hssi_fifo_rx_pcs_data_out_10g[27], w_hssi_fifo_rx_pcs_data_out_10g[26], w_hssi_fifo_rx_pcs_data_out_10g[25], w_hssi_fifo_rx_pcs_data_out_10g[24], w_hssi_fifo_rx_pcs_data_out_10g[23], w_hssi_fifo_rx_pcs_data_out_10g[22], w_hssi_fifo_rx_pcs_data_out_10g[21], w_hssi_fifo_rx_pcs_data_out_10g[20], w_hssi_fifo_rx_pcs_data_out_10g[19], w_hssi_fifo_rx_pcs_data_out_10g[18], w_hssi_fifo_rx_pcs_data_out_10g[17], w_hssi_fifo_rx_pcs_data_out_10g[16], w_hssi_fifo_rx_pcs_data_out_10g[15], w_hssi_fifo_rx_pcs_data_out_10g[14], w_hssi_fifo_rx_pcs_data_out_10g[13], w_hssi_fifo_rx_pcs_data_out_10g[12], w_hssi_fifo_rx_pcs_data_out_10g[11], w_hssi_fifo_rx_pcs_data_out_10g[10], w_hssi_fifo_rx_pcs_data_out_10g[9], w_hssi_fifo_rx_pcs_data_out_10g[8], w_hssi_fifo_rx_pcs_data_out_10g[7], w_hssi_fifo_rx_pcs_data_out_10g[6], w_hssi_fifo_rx_pcs_data_out_10g[5], w_hssi_fifo_rx_pcs_data_out_10g[4], w_hssi_fifo_rx_pcs_data_out_10g[3], w_hssi_fifo_rx_pcs_data_out_10g[2], w_hssi_fifo_rx_pcs_data_out_10g[1], w_hssi_fifo_rx_pcs_data_out_10g[0]}),
				.rx_fifo_rd_data_dw({w_hssi_fifo_rx_pcs_data_out2_10g[73], w_hssi_fifo_rx_pcs_data_out2_10g[72], w_hssi_fifo_rx_pcs_data_out2_10g[71], w_hssi_fifo_rx_pcs_data_out2_10g[70], w_hssi_fifo_rx_pcs_data_out2_10g[69], w_hssi_fifo_rx_pcs_data_out2_10g[68], w_hssi_fifo_rx_pcs_data_out2_10g[67], w_hssi_fifo_rx_pcs_data_out2_10g[66], w_hssi_fifo_rx_pcs_data_out2_10g[65], w_hssi_fifo_rx_pcs_data_out2_10g[64], w_hssi_fifo_rx_pcs_data_out2_10g[63], w_hssi_fifo_rx_pcs_data_out2_10g[62], w_hssi_fifo_rx_pcs_data_out2_10g[61], w_hssi_fifo_rx_pcs_data_out2_10g[60], w_hssi_fifo_rx_pcs_data_out2_10g[59], w_hssi_fifo_rx_pcs_data_out2_10g[58], w_hssi_fifo_rx_pcs_data_out2_10g[57], w_hssi_fifo_rx_pcs_data_out2_10g[56], w_hssi_fifo_rx_pcs_data_out2_10g[55], w_hssi_fifo_rx_pcs_data_out2_10g[54], w_hssi_fifo_rx_pcs_data_out2_10g[53], w_hssi_fifo_rx_pcs_data_out2_10g[52], w_hssi_fifo_rx_pcs_data_out2_10g[51], w_hssi_fifo_rx_pcs_data_out2_10g[50], w_hssi_fifo_rx_pcs_data_out2_10g[49], w_hssi_fifo_rx_pcs_data_out2_10g[48], w_hssi_fifo_rx_pcs_data_out2_10g[47], w_hssi_fifo_rx_pcs_data_out2_10g[46], w_hssi_fifo_rx_pcs_data_out2_10g[45], w_hssi_fifo_rx_pcs_data_out2_10g[44], w_hssi_fifo_rx_pcs_data_out2_10g[43], w_hssi_fifo_rx_pcs_data_out2_10g[42], w_hssi_fifo_rx_pcs_data_out2_10g[41], w_hssi_fifo_rx_pcs_data_out2_10g[40], w_hssi_fifo_rx_pcs_data_out2_10g[39], w_hssi_fifo_rx_pcs_data_out2_10g[38], w_hssi_fifo_rx_pcs_data_out2_10g[37], w_hssi_fifo_rx_pcs_data_out2_10g[36], w_hssi_fifo_rx_pcs_data_out2_10g[35], w_hssi_fifo_rx_pcs_data_out2_10g[34], w_hssi_fifo_rx_pcs_data_out2_10g[33], w_hssi_fifo_rx_pcs_data_out2_10g[32], w_hssi_fifo_rx_pcs_data_out2_10g[31], w_hssi_fifo_rx_pcs_data_out2_10g[30], w_hssi_fifo_rx_pcs_data_out2_10g[29], w_hssi_fifo_rx_pcs_data_out2_10g[28], w_hssi_fifo_rx_pcs_data_out2_10g[27], w_hssi_fifo_rx_pcs_data_out2_10g[26], w_hssi_fifo_rx_pcs_data_out2_10g[25], w_hssi_fifo_rx_pcs_data_out2_10g[24], w_hssi_fifo_rx_pcs_data_out2_10g[23], w_hssi_fifo_rx_pcs_data_out2_10g[22], w_hssi_fifo_rx_pcs_data_out2_10g[21], w_hssi_fifo_rx_pcs_data_out2_10g[20], w_hssi_fifo_rx_pcs_data_out2_10g[19], w_hssi_fifo_rx_pcs_data_out2_10g[18], w_hssi_fifo_rx_pcs_data_out2_10g[17], w_hssi_fifo_rx_pcs_data_out2_10g[16], w_hssi_fifo_rx_pcs_data_out2_10g[15], w_hssi_fifo_rx_pcs_data_out2_10g[14], w_hssi_fifo_rx_pcs_data_out2_10g[13], w_hssi_fifo_rx_pcs_data_out2_10g[12], w_hssi_fifo_rx_pcs_data_out2_10g[11], w_hssi_fifo_rx_pcs_data_out2_10g[10], w_hssi_fifo_rx_pcs_data_out2_10g[9], w_hssi_fifo_rx_pcs_data_out2_10g[8], w_hssi_fifo_rx_pcs_data_out2_10g[7], w_hssi_fifo_rx_pcs_data_out2_10g[6], w_hssi_fifo_rx_pcs_data_out2_10g[5], w_hssi_fifo_rx_pcs_data_out2_10g[4], w_hssi_fifo_rx_pcs_data_out2_10g[3], w_hssi_fifo_rx_pcs_data_out2_10g[2], w_hssi_fifo_rx_pcs_data_out2_10g[1], w_hssi_fifo_rx_pcs_data_out2_10g[0]}),
				.rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.rx_pma_data({w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0]}),
				.rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.signal_ok_krfec(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_10g_reg(),
				.pld_10g_krfec_rx_blk_lock_10g_txclk_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_txclk_reg(),
				.pld_10g_krfec_rx_frame_10g_reg(),
				.pld_10g_krfec_rx_frame_10g_txclk_reg(),
				.pld_10g_krfec_rx_pld_rst_n_fifo(),
				.pld_10g_krfec_rx_pld_rst_n_reg(),
				.pld_10g_krfec_rx_pld_rst_n_txclk_reg(),
				.pld_10g_rx_align_clr_fifo(),
				.pld_10g_rx_align_clr_reg(),
				.pld_10g_rx_align_clr_txclk_reg(),
				.pld_10g_rx_align_val_fifo(),
				.pld_10g_rx_align_val_reg(),
				.pld_10g_rx_align_val_txclk_reg(),
				.pld_10g_rx_clr_ber_count_reg(),
				.pld_10g_rx_clr_ber_count_txclk_reg(),
				.pld_10g_rx_crc32_err_reg(),
				.pld_10g_rx_crc32_err_txclk_reg(),
				.pld_10g_rx_data_valid_10g_reg(),
				.pld_10g_rx_data_valid_fifo(),
				.pld_10g_rx_data_valid_pcsdirect_reg(),
				.pld_10g_rx_data_valid_txclk_reg(),
				.pld_10g_rx_empty_fifo(),
				.pld_10g_rx_fifo_del_reg(),
				.pld_10g_rx_fifo_del_txclk_reg(),
				.pld_10g_rx_fifo_insert_fifo(),
				.pld_10g_rx_fifo_num_reg(),
				.pld_10g_rx_fifo_num_txclk_reg(),
				.pld_10g_rx_frame_lock_reg(),
				.pld_10g_rx_frame_lock_txclk_reg(),
				.pld_10g_rx_hi_ber_reg(),
				.pld_10g_rx_hi_ber_txclk_reg(),
				.pld_10g_rx_oflw_err_reg(),
				.pld_10g_rx_oflw_err_txclk_reg(),
				.pld_10g_rx_pempty_fifo(),
				.pld_10g_rx_pfull_reg(),
				.pld_10g_rx_pfull_txclk_reg(),
				.pld_10g_rx_rd_en_fifo(),
				.pld_pcs_rx_clk_out_10g_txclk_wire(),
				.pld_pcs_rx_clk_out_10g_wire(),
				.pld_rx_control_10g_reg(),
				.pld_rx_control_10g_txclk_reg(),
				.pld_rx_data_10g_reg(),
				.pld_rx_data_10g_txclk_reg(),
				.pld_rx_prbs_err_10g_txclk_reg(),
				.pld_rx_prbs_err_clr_10g_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_10g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_align_val = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_blk_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_control[19:0] = 20'b0;
				assign w_hssi_10g_rx_pcs_rx_crc32_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_data[127:0] = 128'b0;
				assign w_hssi_10g_rx_pcs_rx_data_valid = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_dft_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_diag_status[1:0] = 2'b0;
				assign w_hssi_10g_rx_pcs_rx_empty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fec_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_del = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_insert = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_data[73:0] = 74'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_frame_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_hi_ber = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_oflw_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pempty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pfull = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_random_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_rx_frame = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_10g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_tx_pcs
			twentynm_hssi_10g_tx_pcs #(
				.advanced_user_mode(hssi_10g_tx_pcs_advanced_user_mode),
				.bitslip_en(hssi_10g_tx_pcs_bitslip_en),
				.bonding_dft_en(hssi_10g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_10g_tx_pcs_bonding_dft_val),
				.comp_cnt(hssi_10g_tx_pcs_comp_cnt),
				.compin_sel(hssi_10g_tx_pcs_compin_sel),
				.crcgen_bypass(hssi_10g_tx_pcs_crcgen_bypass),
				.crcgen_clken(hssi_10g_tx_pcs_crcgen_clken),
				.crcgen_err(hssi_10g_tx_pcs_crcgen_err),
				.crcgen_inv(hssi_10g_tx_pcs_crcgen_inv),
				.ctrl_bit_reverse(hssi_10g_tx_pcs_ctrl_bit_reverse),
				.ctrl_plane_bonding(hssi_10g_tx_pcs_ctrl_plane_bonding),
				.data_bit_reverse(hssi_10g_tx_pcs_data_bit_reverse),
				.dft_clk_out_sel(hssi_10g_tx_pcs_dft_clk_out_sel),
				.dispgen_bypass(hssi_10g_tx_pcs_dispgen_bypass),
				.dispgen_clken(hssi_10g_tx_pcs_dispgen_clken),
				.dispgen_err(hssi_10g_tx_pcs_dispgen_err),
				.dispgen_pipeln(hssi_10g_tx_pcs_dispgen_pipeln),
				.distdwn_bypass_pipeln(hssi_10g_tx_pcs_distdwn_bypass_pipeln),
				.distdwn_master(hssi_10g_tx_pcs_distdwn_master),
				.distup_bypass_pipeln(hssi_10g_tx_pcs_distup_bypass_pipeln),
				.distup_master(hssi_10g_tx_pcs_distup_master),
				.dv_bond(hssi_10g_tx_pcs_dv_bond),
				.empty_flag_type(hssi_10g_tx_pcs_empty_flag_type),
				.enc64b66b_txsm_clken(hssi_10g_tx_pcs_enc64b66b_txsm_clken),
				.enc_64b66b_txsm_bypass(hssi_10g_tx_pcs_enc_64b66b_txsm_bypass),
				.fastpath(hssi_10g_tx_pcs_fastpath),
				.fec_clken(hssi_10g_tx_pcs_fec_clken),
				.fec_enable(hssi_10g_tx_pcs_fec_enable),
				.fifo_double_write(hssi_10g_tx_pcs_fifo_double_write),
				.fifo_reg_fast(hssi_10g_tx_pcs_fifo_reg_fast),
				.fifo_stop_rd(hssi_10g_tx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_tx_pcs_fifo_stop_wr),
				.frmgen_burst(hssi_10g_tx_pcs_frmgen_burst),
				.frmgen_bypass(hssi_10g_tx_pcs_frmgen_bypass),
				.frmgen_clken(hssi_10g_tx_pcs_frmgen_clken),
				.frmgen_mfrm_length(hssi_10g_tx_pcs_frmgen_mfrm_length),
				.frmgen_pipeln(hssi_10g_tx_pcs_frmgen_pipeln),
				.frmgen_pyld_ins(hssi_10g_tx_pcs_frmgen_pyld_ins),
				.frmgen_wordslip(hssi_10g_tx_pcs_frmgen_wordslip),
				.full_flag_type(hssi_10g_tx_pcs_full_flag_type),
				.gb_pipeln_bypass(hssi_10g_tx_pcs_gb_pipeln_bypass),
				.gb_tx_idwidth(hssi_10g_tx_pcs_gb_tx_idwidth),
				.gb_tx_odwidth(hssi_10g_tx_pcs_gb_tx_odwidth),
				.gbred_clken(hssi_10g_tx_pcs_gbred_clken),
				.indv(hssi_10g_tx_pcs_indv),
				.low_latency_en(hssi_10g_tx_pcs_low_latency_en),
				.master_clk_sel(hssi_10g_tx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_tx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_tx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_tx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_tx_pcs_pld_if_type),
				.prot_mode(hssi_10g_tx_pcs_prot_mode),
				.pseudo_random(hssi_10g_tx_pcs_pseudo_random),
				.pseudo_seed_a(hssi_10g_tx_pcs_pseudo_seed_a),
				.pseudo_seed_b(hssi_10g_tx_pcs_pseudo_seed_b),
				.random_disp(hssi_10g_tx_pcs_random_disp),
				.rdfifo_clken(hssi_10g_tx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_tx_pcs_reconfig_settings),
				.scrm_bypass(hssi_10g_tx_pcs_scrm_bypass),
				.scrm_clken(hssi_10g_tx_pcs_scrm_clken),
				.scrm_mode(hssi_10g_tx_pcs_scrm_mode),
				.scrm_pipeln(hssi_10g_tx_pcs_scrm_pipeln),
				.sh_err(hssi_10g_tx_pcs_sh_err),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sop_mark(hssi_10g_tx_pcs_sop_mark),
				.stretch_num_stages(hssi_10g_tx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_tx_pcs_sup_mode),
				.test_mode(hssi_10g_tx_pcs_test_mode),
				.tx_scrm_err(hssi_10g_tx_pcs_tx_scrm_err),
				.tx_scrm_width(hssi_10g_tx_pcs_tx_scrm_width),
				.tx_sh_location(hssi_10g_tx_pcs_tx_sh_location),
				.tx_sm_bypass(hssi_10g_tx_pcs_tx_sm_bypass),
				.tx_sm_pipeln(hssi_10g_tx_pcs_tx_sm_pipeln),
				.tx_testbus_sel(hssi_10g_tx_pcs_tx_testbus_sel),
				.txfifo_empty(hssi_10g_tx_pcs_txfifo_empty),
				.txfifo_full(hssi_10g_tx_pcs_txfifo_full),
				.txfifo_mode(hssi_10g_tx_pcs_txfifo_mode),
				.txfifo_pempty(hssi_10g_tx_pcs_txfifo_pempty),
				.txfifo_pfull(hssi_10g_tx_pcs_txfifo_pfull),
				.wr_clk_sel(hssi_10g_tx_pcs_wr_clk_sel),
				.wrfifo_clken(hssi_10g_tx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_tx_pcs_blockselect),
				.distdwn_out_dv(w_hssi_10g_tx_pcs_distdwn_out_dv),
				.distdwn_out_rden(w_hssi_10g_tx_pcs_distdwn_out_rden),
				.distdwn_out_wren(w_hssi_10g_tx_pcs_distdwn_out_wren),
				.distup_out_dv(w_hssi_10g_tx_pcs_distup_out_dv),
				.distup_out_rden(w_hssi_10g_tx_pcs_distup_out_rden),
				.distup_out_wren(w_hssi_10g_tx_pcs_distup_out_wren),
				.tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pma_if(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.tx_control_out_krfec(w_hssi_10g_tx_pcs_tx_control_out_krfec),
				.tx_data_out_krfec(w_hssi_10g_tx_pcs_tx_data_out_krfec),
				.tx_data_valid_out_krfec(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.tx_fec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_fifo_num(w_hssi_10g_tx_pcs_tx_fifo_num),
				.tx_fifo_rd_ptr(w_hssi_10g_tx_pcs_tx_fifo_rd_ptr),
				.tx_fifo_wr_clk(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.tx_fifo_wr_data(w_hssi_10g_tx_pcs_tx_fifo_wr_data),
				.tx_fifo_wr_data_dw(w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw),
				.tx_fifo_wr_en(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.tx_fifo_wr_ptr(w_hssi_10g_tx_pcs_tx_fifo_wr_ptr),
				.tx_fifo_wr_rst_n(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.tx_full(w_hssi_10g_tx_pcs_tx_full),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				.tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.tx_pma_data(w_hssi_10g_tx_pcs_tx_pma_data),
				.tx_pma_gating_val(w_hssi_10g_tx_pcs_tx_pma_gating_val),
				.tx_test_data(w_hssi_10g_tx_pcs_tx_test_data),
				.tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.distdwn_in_dv(in_bond_pcs10g_in_bot[2]),
				.distdwn_in_rden(in_bond_pcs10g_in_bot[4]),
				.distdwn_in_wren(in_bond_pcs10g_in_bot[3]),
				.distup_in_dv(in_bond_pcs10g_in_top[2]),
				.distup_in_rden(in_bond_pcs10g_in_top[4]),
				.distup_in_wren(in_bond_pcs10g_in_top[3]),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_tx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_tx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.tx_bitslip({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0]}),
				.tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.tx_control({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0]}),
				.tx_control_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0]}),
				.tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0]}),
				.tx_data_in_krfec({w_hssi_krfec_tx_pcs_tx_data_out[63], w_hssi_krfec_tx_pcs_tx_data_out[62], w_hssi_krfec_tx_pcs_tx_data_out[61], w_hssi_krfec_tx_pcs_tx_data_out[60], w_hssi_krfec_tx_pcs_tx_data_out[59], w_hssi_krfec_tx_pcs_tx_data_out[58], w_hssi_krfec_tx_pcs_tx_data_out[57], w_hssi_krfec_tx_pcs_tx_data_out[56], w_hssi_krfec_tx_pcs_tx_data_out[55], w_hssi_krfec_tx_pcs_tx_data_out[54], w_hssi_krfec_tx_pcs_tx_data_out[53], w_hssi_krfec_tx_pcs_tx_data_out[52], w_hssi_krfec_tx_pcs_tx_data_out[51], w_hssi_krfec_tx_pcs_tx_data_out[50], w_hssi_krfec_tx_pcs_tx_data_out[49], w_hssi_krfec_tx_pcs_tx_data_out[48], w_hssi_krfec_tx_pcs_tx_data_out[47], w_hssi_krfec_tx_pcs_tx_data_out[46], w_hssi_krfec_tx_pcs_tx_data_out[45], w_hssi_krfec_tx_pcs_tx_data_out[44], w_hssi_krfec_tx_pcs_tx_data_out[43], w_hssi_krfec_tx_pcs_tx_data_out[42], w_hssi_krfec_tx_pcs_tx_data_out[41], w_hssi_krfec_tx_pcs_tx_data_out[40], w_hssi_krfec_tx_pcs_tx_data_out[39], w_hssi_krfec_tx_pcs_tx_data_out[38], w_hssi_krfec_tx_pcs_tx_data_out[37], w_hssi_krfec_tx_pcs_tx_data_out[36], w_hssi_krfec_tx_pcs_tx_data_out[35], w_hssi_krfec_tx_pcs_tx_data_out[34], w_hssi_krfec_tx_pcs_tx_data_out[33], w_hssi_krfec_tx_pcs_tx_data_out[32], w_hssi_krfec_tx_pcs_tx_data_out[31], w_hssi_krfec_tx_pcs_tx_data_out[30], w_hssi_krfec_tx_pcs_tx_data_out[29], w_hssi_krfec_tx_pcs_tx_data_out[28], w_hssi_krfec_tx_pcs_tx_data_out[27], w_hssi_krfec_tx_pcs_tx_data_out[26], w_hssi_krfec_tx_pcs_tx_data_out[25], w_hssi_krfec_tx_pcs_tx_data_out[24], w_hssi_krfec_tx_pcs_tx_data_out[23], w_hssi_krfec_tx_pcs_tx_data_out[22], w_hssi_krfec_tx_pcs_tx_data_out[21], w_hssi_krfec_tx_pcs_tx_data_out[20], w_hssi_krfec_tx_pcs_tx_data_out[19], w_hssi_krfec_tx_pcs_tx_data_out[18], w_hssi_krfec_tx_pcs_tx_data_out[17], w_hssi_krfec_tx_pcs_tx_data_out[16], w_hssi_krfec_tx_pcs_tx_data_out[15], w_hssi_krfec_tx_pcs_tx_data_out[14], w_hssi_krfec_tx_pcs_tx_data_out[13], w_hssi_krfec_tx_pcs_tx_data_out[12], w_hssi_krfec_tx_pcs_tx_data_out[11], w_hssi_krfec_tx_pcs_tx_data_out[10], w_hssi_krfec_tx_pcs_tx_data_out[9], w_hssi_krfec_tx_pcs_tx_data_out[8], w_hssi_krfec_tx_pcs_tx_data_out[7], w_hssi_krfec_tx_pcs_tx_data_out[6], w_hssi_krfec_tx_pcs_tx_data_out[5], w_hssi_krfec_tx_pcs_tx_data_out[4], w_hssi_krfec_tx_pcs_tx_data_out[3], w_hssi_krfec_tx_pcs_tx_data_out[2], w_hssi_krfec_tx_pcs_tx_data_out[1], w_hssi_krfec_tx_pcs_tx_data_out[0]}),
				.tx_data_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0]}),
				.tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.tx_diag_status({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0]}),
				.tx_fifo_rd_data({w_hssi_fifo_tx_pcs_data_out_10g[72], w_hssi_fifo_tx_pcs_data_out_10g[71], w_hssi_fifo_tx_pcs_data_out_10g[70], w_hssi_fifo_tx_pcs_data_out_10g[69], w_hssi_fifo_tx_pcs_data_out_10g[68], w_hssi_fifo_tx_pcs_data_out_10g[67], w_hssi_fifo_tx_pcs_data_out_10g[66], w_hssi_fifo_tx_pcs_data_out_10g[65], w_hssi_fifo_tx_pcs_data_out_10g[64], w_hssi_fifo_tx_pcs_data_out_10g[63], w_hssi_fifo_tx_pcs_data_out_10g[62], w_hssi_fifo_tx_pcs_data_out_10g[61], w_hssi_fifo_tx_pcs_data_out_10g[60], w_hssi_fifo_tx_pcs_data_out_10g[59], w_hssi_fifo_tx_pcs_data_out_10g[58], w_hssi_fifo_tx_pcs_data_out_10g[57], w_hssi_fifo_tx_pcs_data_out_10g[56], w_hssi_fifo_tx_pcs_data_out_10g[55], w_hssi_fifo_tx_pcs_data_out_10g[54], w_hssi_fifo_tx_pcs_data_out_10g[53], w_hssi_fifo_tx_pcs_data_out_10g[52], w_hssi_fifo_tx_pcs_data_out_10g[51], w_hssi_fifo_tx_pcs_data_out_10g[50], w_hssi_fifo_tx_pcs_data_out_10g[49], w_hssi_fifo_tx_pcs_data_out_10g[48], w_hssi_fifo_tx_pcs_data_out_10g[47], w_hssi_fifo_tx_pcs_data_out_10g[46], w_hssi_fifo_tx_pcs_data_out_10g[45], w_hssi_fifo_tx_pcs_data_out_10g[44], w_hssi_fifo_tx_pcs_data_out_10g[43], w_hssi_fifo_tx_pcs_data_out_10g[42], w_hssi_fifo_tx_pcs_data_out_10g[41], w_hssi_fifo_tx_pcs_data_out_10g[40], w_hssi_fifo_tx_pcs_data_out_10g[39], w_hssi_fifo_tx_pcs_data_out_10g[38], w_hssi_fifo_tx_pcs_data_out_10g[37], w_hssi_fifo_tx_pcs_data_out_10g[36], w_hssi_fifo_tx_pcs_data_out_10g[35], w_hssi_fifo_tx_pcs_data_out_10g[34], w_hssi_fifo_tx_pcs_data_out_10g[33], w_hssi_fifo_tx_pcs_data_out_10g[32], w_hssi_fifo_tx_pcs_data_out_10g[31], w_hssi_fifo_tx_pcs_data_out_10g[30], w_hssi_fifo_tx_pcs_data_out_10g[29], w_hssi_fifo_tx_pcs_data_out_10g[28], w_hssi_fifo_tx_pcs_data_out_10g[27], w_hssi_fifo_tx_pcs_data_out_10g[26], w_hssi_fifo_tx_pcs_data_out_10g[25], w_hssi_fifo_tx_pcs_data_out_10g[24], w_hssi_fifo_tx_pcs_data_out_10g[23], w_hssi_fifo_tx_pcs_data_out_10g[22], w_hssi_fifo_tx_pcs_data_out_10g[21], w_hssi_fifo_tx_pcs_data_out_10g[20], w_hssi_fifo_tx_pcs_data_out_10g[19], w_hssi_fifo_tx_pcs_data_out_10g[18], w_hssi_fifo_tx_pcs_data_out_10g[17], w_hssi_fifo_tx_pcs_data_out_10g[16], w_hssi_fifo_tx_pcs_data_out_10g[15], w_hssi_fifo_tx_pcs_data_out_10g[14], w_hssi_fifo_tx_pcs_data_out_10g[13], w_hssi_fifo_tx_pcs_data_out_10g[12], w_hssi_fifo_tx_pcs_data_out_10g[11], w_hssi_fifo_tx_pcs_data_out_10g[10], w_hssi_fifo_tx_pcs_data_out_10g[9], w_hssi_fifo_tx_pcs_data_out_10g[8], w_hssi_fifo_tx_pcs_data_out_10g[7], w_hssi_fifo_tx_pcs_data_out_10g[6], w_hssi_fifo_tx_pcs_data_out_10g[5], w_hssi_fifo_tx_pcs_data_out_10g[4], w_hssi_fifo_tx_pcs_data_out_10g[3], w_hssi_fifo_tx_pcs_data_out_10g[2], w_hssi_fifo_tx_pcs_data_out_10g[1], w_hssi_fifo_tx_pcs_data_out_10g[0]}),
				.tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_10g_reg(),
				.pld_10g_krfec_tx_pld_rst_n_fifo(),
				.pld_10g_krfec_tx_pld_rst_n_reg(),
				.pld_10g_tx_bitslip_reg(),
				.pld_10g_tx_burst_en_exe_reg(),
				.pld_10g_tx_data_valid_10g_reg(),
				.pld_10g_tx_data_valid_fifo(),
				.pld_10g_tx_data_valid_reg(),
				.pld_10g_tx_diag_status_reg(),
				.pld_10g_tx_empty_reg(),
				.pld_10g_tx_fifo_num_reg(),
				.pld_10g_tx_full_fifo(),
				.pld_10g_tx_full_reg(),
				.pld_10g_tx_pempty_reg(),
				.pld_10g_tx_pfull_fifo(),
				.pld_10g_tx_wordslip_exe_reg(),
				.pld_10g_tx_wordslip_reg(),
				.pld_pcs_tx_clk_out_10g_wire(),
				.pld_tx_burst_en_reg(),
				.pld_tx_control_lo_10g_reg(),
				.pld_tx_data_10g_fifo(),
				.pld_tx_data_lo_10g_reg()
			);
		end // if generate
		else begin
				assign w_hssi_10g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_burst_en_exe = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pma_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_control_out_krfec[8:0] = 9'b0;
				assign w_hssi_10g_tx_pcs_tx_data_out_krfec[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_data_valid_out_krfec = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_dft_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_empty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fec_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_full = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_pempty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pfull = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_gating_val[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_test_data[19:0] = 20'b0;
				assign w_hssi_10g_tx_pcs_tx_wordslip_exe = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_rx_pcs
			twentynm_hssi_8g_rx_pcs #(
				.auto_error_replacement(hssi_8g_rx_pcs_auto_error_replacement),
				.auto_speed_nego(hssi_8g_rx_pcs_auto_speed_nego),
				.bit_reversal(hssi_8g_rx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_rx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_rx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_rx_pcs_bypass_pipeline_reg),
				.byte_deserializer(hssi_8g_rx_pcs_byte_deserializer),
				.cdr_ctrl_rxvalid_mask(hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask),
				.clkcmp_pattern_n(hssi_8g_rx_pcs_clkcmp_pattern_n),
				.clkcmp_pattern_p(hssi_8g_rx_pcs_clkcmp_pattern_p),
				.clock_gate_bds_dec_asn(hssi_8g_rx_pcs_clock_gate_bds_dec_asn),
				.clock_gate_cdr_eidle(hssi_8g_rx_pcs_clock_gate_cdr_eidle),
				.clock_gate_dw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk),
				.clock_gate_dw_rm_rd(hssi_8g_rx_pcs_clock_gate_dw_rm_rd),
				.clock_gate_dw_rm_wr(hssi_8g_rx_pcs_clock_gate_dw_rm_wr),
				.clock_gate_dw_wa(hssi_8g_rx_pcs_clock_gate_dw_wa),
				.clock_gate_pc_rdclk(hssi_8g_rx_pcs_clock_gate_pc_rdclk),
				.clock_gate_sw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk),
				.clock_gate_sw_rm_rd(hssi_8g_rx_pcs_clock_gate_sw_rm_rd),
				.clock_gate_sw_rm_wr(hssi_8g_rx_pcs_clock_gate_sw_rm_wr),
				.clock_gate_sw_wa(hssi_8g_rx_pcs_clock_gate_sw_wa),
				.clock_observation_in_pld_core(hssi_8g_rx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_rx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_rx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_rx_pcs_ctrl_plane_bonding_distribution),
				.eidle_entry_eios(hssi_8g_rx_pcs_eidle_entry_eios),
				.eidle_entry_iei(hssi_8g_rx_pcs_eidle_entry_iei),
				.eidle_entry_sd(hssi_8g_rx_pcs_eidle_entry_sd),
				.eightb_tenb_decoder(hssi_8g_rx_pcs_eightb_tenb_decoder),
				.err_flags_sel(hssi_8g_rx_pcs_err_flags_sel),
				.fixed_pat_det(hssi_8g_rx_pcs_fixed_pat_det),
				.fixed_pat_num(hssi_8g_rx_pcs_fixed_pat_num),
				.force_signal_detect(hssi_8g_rx_pcs_force_signal_detect),
				.gen3_clk_en(hssi_8g_rx_pcs_gen3_clk_en),
				.gen3_rx_clk_sel(hssi_8g_rx_pcs_gen3_rx_clk_sel),
				.gen3_tx_clk_sel(hssi_8g_rx_pcs_gen3_tx_clk_sel),
				.hip_mode(hssi_8g_rx_pcs_hip_mode),
				.ibm_invalid_code(hssi_8g_rx_pcs_ibm_invalid_code),
				.invalid_code_flag_only(hssi_8g_rx_pcs_invalid_code_flag_only),
				.pad_or_edb_error_replace(hssi_8g_rx_pcs_pad_or_edb_error_replace),
				.pcs_bypass(hssi_8g_rx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_rx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_rx_pcs_phase_compensation_fifo),
				.pipe_if_enable(hssi_8g_rx_pcs_pipe_if_enable),
				.pma_dw(hssi_8g_rx_pcs_pma_dw),
				.polinv_8b10b_dec(hssi_8g_rx_pcs_polinv_8b10b_dec),
				.prot_mode(hssi_8g_rx_pcs_prot_mode),
				.rate_match(hssi_8g_rx_pcs_rate_match),
				.rate_match_del_thres(hssi_8g_rx_pcs_rate_match_del_thres),
				.rate_match_empty_thres(hssi_8g_rx_pcs_rate_match_empty_thres),
				.rate_match_full_thres(hssi_8g_rx_pcs_rate_match_full_thres),
				.rate_match_ins_thres(hssi_8g_rx_pcs_rate_match_ins_thres),
				.rate_match_start_thres(hssi_8g_rx_pcs_rate_match_start_thres),
				.reconfig_settings(hssi_8g_rx_pcs_reconfig_settings),
				.rx_clk2(hssi_8g_rx_pcs_rx_clk2),
				.rx_clk_free_running(hssi_8g_rx_pcs_rx_clk_free_running),
				.rx_pcs_urst(hssi_8g_rx_pcs_rx_pcs_urst),
				.rx_rcvd_clk(hssi_8g_rx_pcs_rx_rcvd_clk),
				.rx_rd_clk(hssi_8g_rx_pcs_rx_rd_clk),
				.rx_refclk(hssi_8g_rx_pcs_rx_refclk),
				.rx_wr_clk(hssi_8g_rx_pcs_rx_wr_clk),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_rx_pcs_sup_mode),
				.symbol_swap(hssi_8g_rx_pcs_symbol_swap),
				.sync_sm_idle_eios(hssi_8g_rx_pcs_sync_sm_idle_eios),
				.test_bus_sel(hssi_8g_rx_pcs_test_bus_sel),
				.tx_rx_parallel_loopback(hssi_8g_rx_pcs_tx_rx_parallel_loopback),
				.wa_boundary_lock_ctrl(hssi_8g_rx_pcs_wa_boundary_lock_ctrl),
				.wa_clk_slip_spacing(hssi_8g_rx_pcs_wa_clk_slip_spacing),
				.wa_det_latency_sync_status_beh(hssi_8g_rx_pcs_wa_det_latency_sync_status_beh),
				.wa_disp_err_flag(hssi_8g_rx_pcs_wa_disp_err_flag),
				.wa_kchar(hssi_8g_rx_pcs_wa_kchar),
				.wa_pd(hssi_8g_rx_pcs_wa_pd),
				.wa_pd_data(hssi_8g_rx_pcs_wa_pd_data),
				.wa_pd_polarity(hssi_8g_rx_pcs_wa_pd_polarity),
				.wa_pld_controlled(hssi_8g_rx_pcs_wa_pld_controlled),
				.wa_renumber_data(hssi_8g_rx_pcs_wa_renumber_data),
				.wa_rgnumber_data(hssi_8g_rx_pcs_wa_rgnumber_data),
				.wa_rknumber_data(hssi_8g_rx_pcs_wa_rknumber_data),
				.wa_rosnumber_data(hssi_8g_rx_pcs_wa_rosnumber_data),
				.wa_rvnumber_data(hssi_8g_rx_pcs_wa_rvnumber_data),
				.wa_sync_sm_ctrl(hssi_8g_rx_pcs_wa_sync_sm_ctrl),
				.wait_cnt(hssi_8g_rx_pcs_wait_cnt)
			) inst_twentynm_hssi_8g_rx_pcs (
				// OUTPUTS
				.a1a2k1k2flag(w_hssi_8g_rx_pcs_a1a2k1k2flag),
				.avmmreaddata(w_hssi_8g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_rx_pcs_blockselect),
				.chnl_test_bus_out(w_hssi_8g_rx_pcs_chnl_test_bus_out),
				.clock_to_pld(w_hssi_8g_rx_pcs_clock_to_pld),
				.dataout(w_hssi_8g_rx_pcs_dataout),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidle_detected(w_hssi_8g_rx_pcs_eidle_detected),
				.eios_det_cdr_ctrl(w_hssi_8g_rx_pcs_eios_det_cdr_ctrl),
				.g3_rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.g3_rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.gen2ngen1(w_hssi_8g_rx_pcs_gen2ngen1),
				.parallel_rev_loopback(w_hssi_8g_rx_pcs_parallel_rev_loopback),
				.pc_fifo_empty(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.pcfifofull(w_hssi_8g_rx_pcs_pcfifofull),
				.phystatus(w_hssi_8g_rx_pcs_phystatus),
				.pipe_data(w_hssi_8g_rx_pcs_pipe_data),
				.rd_enable_out_chnl_down(w_hssi_8g_rx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_rx_pcs_rd_enable_out_chnl_up),
				.rd_ptr1_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo),
				.rd_ptr2_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo),
				.rd_ptr_rx_phfifo(w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.reset_pc_ptrs_out_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down),
				.reset_pc_ptrs_out_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up),
				.rm_fifo_empty(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.rm_fifo_full(w_hssi_8g_rx_pcs_rm_fifo_full),
				.rx_blk_start(w_hssi_8g_rx_pcs_rx_blk_start),
				.rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.rx_data_valid(w_hssi_8g_rx_pcs_rx_data_valid),
				.rx_div_sync_out_chnl_down(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down),
				.rx_div_sync_out_chnl_up(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up),
				.rx_pipe_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.rx_pipe_soft_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rx_pma_clk_gen3(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_rcvd_clk_gen3(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_rstn_sync2wrfifo_8g(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.rx_sync_hdr(w_hssi_8g_rx_pcs_rx_sync_hdr),
				.rx_we_out_chnl_down(w_hssi_8g_rx_pcs_rx_we_out_chnl_down),
				.rx_we_out_chnl_up(w_hssi_8g_rx_pcs_rx_we_out_chnl_up),
				.rxstatus(w_hssi_8g_rx_pcs_rxstatus),
				.rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.word_align_boundary(w_hssi_8g_rx_pcs_word_align_boundary),
				.wr_clk_rx_phfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_rx_phfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_rx_rmfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_rx_rmfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_data_rx_phfifo(w_hssi_8g_rx_pcs_wr_data_rx_phfifo),
				.wr_data_rx_rmfifo(w_hssi_8g_rx_pcs_wr_data_rx_rmfifo),
				.wr_en_rx_phfifo(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_rx_rmfifo(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_rx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_rx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_rx_phfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo),
				.wr_ptr_rx_rmfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo),
				.wr_rst_n_rx_phfifo(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_rx_rmfifo(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				// INPUTS
				.a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bit_reversal_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.datain({w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0]}),
				.disable_pc_fifo_byte_serdes(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4]),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.eidleinfersel({w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0]}),
				.eios_detected_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.enable_comma_detect(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.gen3_clk_sel(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.hrd_rst(1'b0),
				.inferred_rxvalid_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.pc_fifo_rd_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.pc_fifo_wrdisable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.phystatus_int(w_hssi_pipe_gen1_2_phystatus),
				.phystatus_pcs_gen3(w_hssi_pipe_gen3_phystatus),
				.pipe_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.polarity_inversion(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.rd_data1_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0]}),
				.rd_data2_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0]}),
				.rd_data_rx_phfifo({w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[3]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[3]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.reset_pc_ptrs_asn(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5]),
				.reset_pc_ptrs_in_chnl_down(in_bond_pcs8g_in_bot[12]),
				.reset_pc_ptrs_in_chnl_up(in_bond_pcs8g_in_top[12]),
				.reset_ppm_cntrs_pcs_pma(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7]),
				.rm_fifo_read_enable(1'b0),
				.rm_fifo_write_enable(1'b0),
				.rx_blk_start_pcs_gen3({w_hssi_pipe_gen3_rx_blk_start[3], w_hssi_pipe_gen3_rx_blk_start[2], w_hssi_pipe_gen3_rx_blk_start[1], w_hssi_pipe_gen3_rx_blk_start[0]}),
				.rx_data_pcs_gen3({w_hssi_pipe_gen3_rxd_8gpcs_out[63], w_hssi_pipe_gen3_rxd_8gpcs_out[62], w_hssi_pipe_gen3_rxd_8gpcs_out[61], w_hssi_pipe_gen3_rxd_8gpcs_out[60], w_hssi_pipe_gen3_rxd_8gpcs_out[59], w_hssi_pipe_gen3_rxd_8gpcs_out[58], w_hssi_pipe_gen3_rxd_8gpcs_out[57], w_hssi_pipe_gen3_rxd_8gpcs_out[56], w_hssi_pipe_gen3_rxd_8gpcs_out[55], w_hssi_pipe_gen3_rxd_8gpcs_out[54], w_hssi_pipe_gen3_rxd_8gpcs_out[53], w_hssi_pipe_gen3_rxd_8gpcs_out[52], w_hssi_pipe_gen3_rxd_8gpcs_out[51], w_hssi_pipe_gen3_rxd_8gpcs_out[50], w_hssi_pipe_gen3_rxd_8gpcs_out[49], w_hssi_pipe_gen3_rxd_8gpcs_out[48], w_hssi_pipe_gen3_rxd_8gpcs_out[47], w_hssi_pipe_gen3_rxd_8gpcs_out[46], w_hssi_pipe_gen3_rxd_8gpcs_out[45], w_hssi_pipe_gen3_rxd_8gpcs_out[44], w_hssi_pipe_gen3_rxd_8gpcs_out[43], w_hssi_pipe_gen3_rxd_8gpcs_out[42], w_hssi_pipe_gen3_rxd_8gpcs_out[41], w_hssi_pipe_gen3_rxd_8gpcs_out[40], w_hssi_pipe_gen3_rxd_8gpcs_out[39], w_hssi_pipe_gen3_rxd_8gpcs_out[38], w_hssi_pipe_gen3_rxd_8gpcs_out[37], w_hssi_pipe_gen3_rxd_8gpcs_out[36], w_hssi_pipe_gen3_rxd_8gpcs_out[35], w_hssi_pipe_gen3_rxd_8gpcs_out[34], w_hssi_pipe_gen3_rxd_8gpcs_out[33], w_hssi_pipe_gen3_rxd_8gpcs_out[32], w_hssi_pipe_gen3_rxd_8gpcs_out[31], w_hssi_pipe_gen3_rxd_8gpcs_out[30], w_hssi_pipe_gen3_rxd_8gpcs_out[29], w_hssi_pipe_gen3_rxd_8gpcs_out[28], w_hssi_pipe_gen3_rxd_8gpcs_out[27], w_hssi_pipe_gen3_rxd_8gpcs_out[26], w_hssi_pipe_gen3_rxd_8gpcs_out[25], w_hssi_pipe_gen3_rxd_8gpcs_out[24], w_hssi_pipe_gen3_rxd_8gpcs_out[23], w_hssi_pipe_gen3_rxd_8gpcs_out[22], w_hssi_pipe_gen3_rxd_8gpcs_out[21], w_hssi_pipe_gen3_rxd_8gpcs_out[20], w_hssi_pipe_gen3_rxd_8gpcs_out[19], w_hssi_pipe_gen3_rxd_8gpcs_out[18], w_hssi_pipe_gen3_rxd_8gpcs_out[17], w_hssi_pipe_gen3_rxd_8gpcs_out[16], w_hssi_pipe_gen3_rxd_8gpcs_out[15], w_hssi_pipe_gen3_rxd_8gpcs_out[14], w_hssi_pipe_gen3_rxd_8gpcs_out[13], w_hssi_pipe_gen3_rxd_8gpcs_out[12], w_hssi_pipe_gen3_rxd_8gpcs_out[11], w_hssi_pipe_gen3_rxd_8gpcs_out[10], w_hssi_pipe_gen3_rxd_8gpcs_out[9], w_hssi_pipe_gen3_rxd_8gpcs_out[8], w_hssi_pipe_gen3_rxd_8gpcs_out[7], w_hssi_pipe_gen3_rxd_8gpcs_out[6], w_hssi_pipe_gen3_rxd_8gpcs_out[5], w_hssi_pipe_gen3_rxd_8gpcs_out[4], w_hssi_pipe_gen3_rxd_8gpcs_out[3], w_hssi_pipe_gen3_rxd_8gpcs_out[2], w_hssi_pipe_gen3_rxd_8gpcs_out[1], w_hssi_pipe_gen3_rxd_8gpcs_out[0]}),
				.rx_data_valid_pcs_gen3({w_hssi_pipe_gen3_rxdataskip[3], w_hssi_pipe_gen3_rxdataskip[2], w_hssi_pipe_gen3_rxdataskip[1], w_hssi_pipe_gen3_rxdataskip[0]}),
				.rx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[1], in_bond_pcs8g_in_bot[0]}),
				.rx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[1], in_bond_pcs8g_in_top[0]}),
				.rx_pcs_rst(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.rx_sync_hdr_pcs_gen3({w_hssi_pipe_gen3_rx_sync_hdr[1], w_hssi_pipe_gen3_rx_sync_hdr[0]}),
				.rx_we_in_chnl_down({in_bond_pcs8g_in_bot[5], in_bond_pcs8g_in_bot[4]}),
				.rx_we_in_chnl_up({in_bond_pcs8g_in_top[5], in_bond_pcs8g_in_top[4]}),
				.rxstatus_int({w_hssi_pipe_gen1_2_rxstatus[2], w_hssi_pipe_gen1_2_rxstatus[1], w_hssi_pipe_gen1_2_rxstatus[0]}),
				.rxstatus_pcs_gen3({w_hssi_pipe_gen3_rxstatus[2], w_hssi_pipe_gen3_rxstatus[1], w_hssi_pipe_gen3_rxstatus[0]}),
				.rxvalid_int(w_hssi_pipe_gen1_2_rxvalid),
				.rxvalid_pcs_gen3(w_hssi_pipe_gen3_rxvalid),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.sig_det_from_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_ctrlplane_testbus({w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0]}),
				.tx_div_sync({w_hssi_8g_tx_pcs_tx_div_sync[1], w_hssi_8g_tx_pcs_tx_div_sync[0]}),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.tx_testbus({w_hssi_8g_tx_pcs_tx_testbus[19], w_hssi_8g_tx_pcs_tx_testbus[18], w_hssi_8g_tx_pcs_tx_testbus[17], w_hssi_8g_tx_pcs_tx_testbus[16], w_hssi_8g_tx_pcs_tx_testbus[15], w_hssi_8g_tx_pcs_tx_testbus[14], w_hssi_8g_tx_pcs_tx_testbus[13], w_hssi_8g_tx_pcs_tx_testbus[12], w_hssi_8g_tx_pcs_tx_testbus[11], w_hssi_8g_tx_pcs_tx_testbus[10], w_hssi_8g_tx_pcs_tx_testbus[9], w_hssi_8g_tx_pcs_tx_testbus[8], w_hssi_8g_tx_pcs_tx_testbus[7], w_hssi_8g_tx_pcs_tx_testbus[6], w_hssi_8g_tx_pcs_tx_testbus[5], w_hssi_8g_tx_pcs_tx_testbus[4], w_hssi_8g_tx_pcs_tx_testbus[3], w_hssi_8g_tx_pcs_tx_testbus[2], w_hssi_8g_tx_pcs_tx_testbus[1], w_hssi_8g_tx_pcs_tx_testbus[0]}),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[2]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[2]),
				
				// UNUSED
				.byte_deserializer_pcs_clk_div_by_2_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_wire(),
				.byte_deserializer_pcs_clk_div_by_2_wire(),
				.byte_deserializer_pcs_clk_div_by_4_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_2_reg(),
				.byte_deserializer_pld_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_4_txclk_reg(),
				.pld_8g_a1a2_k1k2_flag_reg(),
				.pld_8g_a1a2_k1k2_flag_txclk_reg(),
				.pld_8g_a1a2_size_reg(),
				.pld_8g_a1a2_size_txclk_reg(),
				.pld_8g_bitloc_rev_en_reg(),
				.pld_8g_bitloc_rev_en_txclk_reg(),
				.pld_8g_byte_rev_en_reg(),
				.pld_8g_byte_rev_en_txclk_reg(),
				.pld_8g_elecidle_reg(),
				.pld_8g_empty_rmf_lowlatency_reg(),
				.pld_8g_empty_rmf_lowlatency_txclk_reg(),
				.pld_8g_empty_rmf_reg(),
				.pld_8g_empty_rmf_txclk_reg(),
				.pld_8g_empty_rx_fifo(),
				.pld_8g_empty_rx_reg(),
				.pld_8g_empty_rx_txclk_reg(),
				.pld_8g_encdt_reg(),
				.pld_8g_encdt_txclk_reg(),
				.pld_8g_full_rmf_reg(),
				.pld_8g_full_rmf_txclk_reg(),
				.pld_8g_full_rx_fifo(),
				.pld_8g_full_rx_reg(),
				.pld_8g_full_rx_txclk_reg(),
				.pld_8g_g3_rx_pld_rst_n_reg(),
				.pld_8g_g3_rx_pld_rst_n_txclk_reg(),
				.pld_8g_rxelecidle_txclk_reg(),
				.pld_8g_rxpolarity_reg(),
				.pld_8g_rxpolarity_txclk_reg(),
				.pld_8g_wa_boundary_reg(),
				.pld_8g_wrdisable_rx_reg(),
				.pld_8g_wrdisable_rx_txclk_reg(),
				.pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_rx_clk_out_8g_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_wire(),
				.pld_rx_control_8g_reg(),
				.pld_rx_control_8g_txclk_reg(),
				.pld_rx_data_8g_reg(),
				.pld_rx_data_8g_txclk_reg(),
				.pld_syncsm_en_reg(),
				.pld_syncsm_en_txclk_reg(),
				.rm_fifo_partial_empty(),
				.rm_fifo_partial_full(),
				.sta_rx_clk2_by2_1(),
				.sta_rx_clk2_by2_1_out(),
				.sta_rx_clk2_by2_2(),
				.sta_rx_clk2_by2_2_out(),
				.sta_rx_clk2_by4_1(),
				.sta_rx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_rx_pcs_a1a2k1k2flag[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_rx_pcs_chnl_test_bus_out[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_clock_to_pld = 1'b0;
				assign w_hssi_8g_rx_pcs_dataout[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_dis_pc_byte = 1'b0;
				assign w_hssi_8g_rx_pcs_eidle_detected = 1'b0;
				assign w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_pma_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_gen2ngen1 = 1'b0;
				assign w_hssi_8g_rx_pcs_parallel_rev_loopback[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_pc_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_pcfifofull = 1'b0;
				assign w_hssi_8g_rx_pcs_phystatus = 1'b0;
				assign w_hssi_8g_rx_pcs_pipe_data[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_full = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clkslip = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_data_valid[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pma_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rxstatus[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_rxvalid = 1'b0;
				assign w_hssi_8g_rx_pcs_signal_detect_out = 1'b0;
				assign w_hssi_8g_rx_pcs_word_align_boundary[4:0] = 5'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79:0] = 80'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31:0] = 32'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_rmfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_tx_pcs
			twentynm_hssi_8g_tx_pcs #(
				.auto_speed_nego_gen2(hssi_8g_tx_pcs_auto_speed_nego_gen2),
				.bit_reversal(hssi_8g_tx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_tx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_tx_pcs_bypass_pipeline_reg),
				.byte_serializer(hssi_8g_tx_pcs_byte_serializer),
				.clock_gate_bs_enc(hssi_8g_tx_pcs_clock_gate_bs_enc),
				.clock_gate_dw_fifowr(hssi_8g_tx_pcs_clock_gate_dw_fifowr),
				.clock_gate_fiford(hssi_8g_tx_pcs_clock_gate_fiford),
				.clock_gate_sw_fifowr(hssi_8g_tx_pcs_clock_gate_sw_fifowr),
				.clock_observation_in_pld_core(hssi_8g_tx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_tx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_tx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_tx_pcs_ctrl_plane_bonding_distribution),
				.data_selection_8b10b_encoder_input(hssi_8g_tx_pcs_data_selection_8b10b_encoder_input),
				.dynamic_clk_switch(hssi_8g_tx_pcs_dynamic_clk_switch),
				.eightb_tenb_disp_ctrl(hssi_8g_tx_pcs_eightb_tenb_disp_ctrl),
				.eightb_tenb_encoder(hssi_8g_tx_pcs_eightb_tenb_encoder),
				.force_echar(hssi_8g_tx_pcs_force_echar),
				.force_kchar(hssi_8g_tx_pcs_force_kchar),
				.gen3_tx_clk_sel(hssi_8g_tx_pcs_gen3_tx_clk_sel),
				.gen3_tx_pipe_clk_sel(hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel),
				.hip_mode(hssi_8g_tx_pcs_hip_mode),
				.pcs_bypass(hssi_8g_tx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_tx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_tx_pcs_phase_compensation_fifo),
				.phfifo_write_clk_sel(hssi_8g_tx_pcs_phfifo_write_clk_sel),
				.pma_dw(hssi_8g_tx_pcs_pma_dw),
				.prot_mode(hssi_8g_tx_pcs_prot_mode),
				.reconfig_settings(hssi_8g_tx_pcs_reconfig_settings),
				.refclk_b_clk_sel(hssi_8g_tx_pcs_refclk_b_clk_sel),
				.revloop_back_rm(hssi_8g_tx_pcs_revloop_back_rm),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_tx_pcs_sup_mode),
				.symbol_swap(hssi_8g_tx_pcs_symbol_swap),
				.tx_bitslip(hssi_8g_tx_pcs_tx_bitslip),
				.tx_compliance_controlled_disparity(hssi_8g_tx_pcs_tx_compliance_controlled_disparity),
				.tx_fast_pld_reg(hssi_8g_tx_pcs_tx_fast_pld_reg),
				.txclk_freerun(hssi_8g_tx_pcs_txclk_freerun),
				.txpcs_urst(hssi_8g_tx_pcs_txpcs_urst)
			) inst_twentynm_hssi_8g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_8g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_tx_pcs_blockselect),
				.clk_out(w_hssi_8g_tx_pcs_clk_out),
				.clk_out_gen3(w_hssi_8g_tx_pcs_clk_out_gen3),
				.dataout(w_hssi_8g_tx_pcs_dataout),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.fifo_select_out_chnl_down(w_hssi_8g_tx_pcs_fifo_select_out_chnl_down),
				.fifo_select_out_chnl_up(w_hssi_8g_tx_pcs_fifo_select_out_chnl_up),
				.g3_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.g3_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
				.non_gray_eidleinfersel(w_hssi_8g_tx_pcs_non_gray_eidleinfersel),
				.ph_fifo_overflow(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.ph_fifo_underflow(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.phfifo_txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.phfifo_txmargin(w_hssi_8g_tx_pcs_phfifo_txmargin),
				.phfifo_txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				.pipe_en_rev_parallel_lpbk_out(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.pipe_power_down_out(w_hssi_8g_tx_pcs_pipe_power_down_out),
				.pipe_tx_clk_out_gen3(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pmaif_asn_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.rd_enable_out_chnl_down(w_hssi_8g_tx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_tx_pcs_rd_enable_out_chnl_up),
				.rd_ptr_tx_phfifo(w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rxpolarity_int(w_hssi_8g_tx_pcs_rxpolarity_int),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.tx_blk_start_out(w_hssi_8g_tx_pcs_tx_blk_start_out),
				.tx_clk_out_8g_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.tx_ctrlplane_testbus(w_hssi_8g_tx_pcs_tx_ctrlplane_testbus),
				.tx_data_out(w_hssi_8g_tx_pcs_tx_data_out),
				.tx_data_valid_out(w_hssi_8g_tx_pcs_tx_data_valid_out),
				.tx_datak_out(w_hssi_8g_tx_pcs_tx_datak_out),
				.tx_detect_rxloopback_int(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.tx_div_sync(w_hssi_8g_tx_pcs_tx_div_sync),
				.tx_div_sync_out_chnl_down(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down),
				.tx_div_sync_out_chnl_up(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up),
				.tx_pipe_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.tx_pipe_electidle(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_soft_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.tx_sync_hdr_out(w_hssi_8g_tx_pcs_tx_sync_hdr_out),
				.tx_testbus(w_hssi_8g_tx_pcs_tx_testbus),
				.txcompliance_out(w_hssi_8g_tx_pcs_txcompliance_out),
				.txelecidle_out(w_hssi_8g_tx_pcs_txelecidle_out),
				.wr_clk_tx_phfifo_dw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_tx_phfifo_sw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_data_tx_phfifo(w_hssi_8g_tx_pcs_wr_data_tx_phfifo),
				.wr_en_tx_phfifo(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_tx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_tx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_tx_phfifo(w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo),
				.wr_rst_n_tx_phfifo(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bitslip_boundary_select({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0]}),
				.clk_sel_gen3(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.coreclk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.datain({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.detectrxloopin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidleinfersel({w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0]}),
				.en_rev_parallel_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.fifo_select_in_chnl_down({in_bond_pcs8g_in_bot[11], in_bond_pcs8g_in_bot[10]}),
				.fifo_select_in_chnl_up({in_bond_pcs8g_in_top[11], in_bond_pcs8g_in_top[10]}),
				.hrdrst(1'b0),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.ph_fifo_rd_disable(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.pipe_en_rev_parallel_lpbk_in(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.pipe_tx_deemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.pipe_tx_margin({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0]}),
				.powerdn({w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0]}),
				.rate_switch(w_hssi_8g_rx_pcs_gen2ngen1),
				.rd_data_tx_phfifo({w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[9]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[9]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.rev_parallel_lpbk_data({w_hssi_8g_rx_pcs_parallel_rev_loopback[19], w_hssi_8g_rx_pcs_parallel_rev_loopback[18], w_hssi_8g_rx_pcs_parallel_rev_loopback[17], w_hssi_8g_rx_pcs_parallel_rev_loopback[16], w_hssi_8g_rx_pcs_parallel_rev_loopback[15], w_hssi_8g_rx_pcs_parallel_rev_loopback[14], w_hssi_8g_rx_pcs_parallel_rev_loopback[13], w_hssi_8g_rx_pcs_parallel_rev_loopback[12], w_hssi_8g_rx_pcs_parallel_rev_loopback[11], w_hssi_8g_rx_pcs_parallel_rev_loopback[10], w_hssi_8g_rx_pcs_parallel_rev_loopback[9], w_hssi_8g_rx_pcs_parallel_rev_loopback[8], w_hssi_8g_rx_pcs_parallel_rev_loopback[7], w_hssi_8g_rx_pcs_parallel_rev_loopback[6], w_hssi_8g_rx_pcs_parallel_rev_loopback[5], w_hssi_8g_rx_pcs_parallel_rev_loopback[4], w_hssi_8g_rx_pcs_parallel_rev_loopback[3], w_hssi_8g_rx_pcs_parallel_rev_loopback[2], w_hssi_8g_rx_pcs_parallel_rev_loopback[1], w_hssi_8g_rx_pcs_parallel_rev_loopback[0]}),
				.rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.tx_blk_start({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0]}),
				.tx_data_valid({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0]}),
				.tx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[7], in_bond_pcs8g_in_bot[6]}),
				.tx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[7], in_bond_pcs8g_in_top[6]}),
				.tx_pcs_reset(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.tx_sync_hdr({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0]}),
				.txd_fast_reg({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0]}),
				.txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[8]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[8]),
				.wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				
				// UNUSED
				.byte_serializer_pcs_clk_div_by_2_reg(),
				.byte_serializer_pcs_clk_div_by_2_wire(),
				.byte_serializer_pcs_clk_div_by_4_reg(),
				.byte_serializer_pld_clk_div_by_2_reg(),
				.byte_serializer_pld_clk_div_by_4_reg(),
				.pld_8g_empty_tx_fifo(),
				.pld_8g_empty_tx_reg(),
				.pld_8g_full_tx_fifo(),
				.pld_8g_full_tx_reg(),
				.pld_8g_g3_tx_pld_rst_n_reg(),
				.pld_8g_rddisable_tx_reg(),
				.pld_8g_tx_boundary_sel_reg(),
				.pld_pcs_tx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_tx_clk_out_8g_wire(),
				.pld_tx_data_8g_fifo(),
				.pld_tx_data_lo_8g_reg(),
				.sta_tx_clk2_by2_1(),
				.sta_tx_clk2_by2_1_out(),
				.sta_tx_clk2_by4_1(),
				.sta_tx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_dataout[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_dyn_clk_switch_n = 1'b1;		// Override default tieoff
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_g3_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_overflow = 1'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_underflow = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txdeemph = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txmargin[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txswing = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_power_down_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_pmaif_asn_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_refclk_b = 1'b0;
				assign w_hssi_8g_tx_pcs_refclk_b_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_rxpolarity_int = 1'b0;
				assign w_hssi_8g_tx_pcs_soft_reset_wclk1_n = 1'b0;
				assign w_hssi_8g_tx_pcs_sw_fifo_wr_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_blk_start_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_tx_data_out[31:0] = 32'b0;
				assign w_hssi_8g_tx_pcs_tx_data_valid_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_datak_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_detect_rxloopback_int = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_electidle = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_sync_hdr_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_txcompliance_out = 1'b0;
				assign w_hssi_8g_tx_pcs_txelecidle_out = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63:0] = 64'b0;
				assign w_hssi_8g_tx_pcs_wr_en_tx_phfifo = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pcs_pma_interface
			twentynm_hssi_common_pcs_pma_interface #(
				.asn_clk_enable(hssi_common_pcs_pma_interface_asn_clk_enable),
				.asn_enable(hssi_common_pcs_pma_interface_asn_enable),
				.block_sel(hssi_common_pcs_pma_interface_block_sel),
				.bypass_early_eios(hssi_common_pcs_pma_interface_bypass_early_eios),
				.bypass_pcie_switch(hssi_common_pcs_pma_interface_bypass_pcie_switch),
				.bypass_pma_ltr(hssi_common_pcs_pma_interface_bypass_pma_ltr),
				.bypass_pma_sw_done(hssi_common_pcs_pma_interface_bypass_pma_sw_done),
				.bypass_ppm_lock(hssi_common_pcs_pma_interface_bypass_ppm_lock),
				.bypass_send_syncp_fbkp(hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp),
				.bypass_txdetectrx(hssi_common_pcs_pma_interface_bypass_txdetectrx),
				.cdr_control(hssi_common_pcs_pma_interface_cdr_control),
				.cid_enable(hssi_common_pcs_pma_interface_cid_enable),
				.cp_cons_sel(hssi_common_pcs_pma_interface_cp_cons_sel),
				.cp_dwn_mstr(hssi_common_pcs_pma_interface_cp_dwn_mstr),
				.cp_up_mstr(hssi_common_pcs_pma_interface_cp_up_mstr),
				.ctrl_plane_bonding(hssi_common_pcs_pma_interface_ctrl_plane_bonding),
				.data_mask_count(hssi_common_pcs_pma_interface_data_mask_count),
				.data_mask_count_multi(hssi_common_pcs_pma_interface_data_mask_count_multi),
				.dft_observation_clock_selection(hssi_common_pcs_pma_interface_dft_observation_clock_selection),
				.early_eios_counter(hssi_common_pcs_pma_interface_early_eios_counter),
				.force_freqdet(hssi_common_pcs_pma_interface_force_freqdet),
				.free_run_clk_enable(hssi_common_pcs_pma_interface_free_run_clk_enable),
				.ignore_sigdet_g23(hssi_common_pcs_pma_interface_ignore_sigdet_g23),
				.pc_en_counter(hssi_common_pcs_pma_interface_pc_en_counter),
				.pc_rst_counter(hssi_common_pcs_pma_interface_pc_rst_counter),
				.pcie_hip_mode(hssi_common_pcs_pma_interface_pcie_hip_mode),
				.ph_fifo_reg_mode(hssi_common_pcs_pma_interface_ph_fifo_reg_mode),
				.phfifo_flush_wait(hssi_common_pcs_pma_interface_phfifo_flush_wait),
				.pipe_if_g3pcs(hssi_common_pcs_pma_interface_pipe_if_g3pcs),
				.pma_done_counter(hssi_common_pcs_pma_interface_pma_done_counter),
				.pma_if_dft_en(hssi_common_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_common_pcs_pma_interface_pma_if_dft_val),
				.ppm_cnt_rst(hssi_common_pcs_pma_interface_ppm_cnt_rst),
				.ppm_deassert_early(hssi_common_pcs_pma_interface_ppm_deassert_early),
				.ppm_det_buckets(hssi_common_pcs_pma_interface_ppm_det_buckets),
				.ppm_gen1_2_cnt(hssi_common_pcs_pma_interface_ppm_gen1_2_cnt),
				.ppm_post_eidle_delay(hssi_common_pcs_pma_interface_ppm_post_eidle_delay),
				.ppmsel(hssi_common_pcs_pma_interface_ppmsel),
				.prot_mode(hssi_common_pcs_pma_interface_prot_mode),
				.reconfig_settings(hssi_common_pcs_pma_interface_reconfig_settings),
				.rxvalid_mask(hssi_common_pcs_pma_interface_rxvalid_mask),
				.sigdet_wait_counter(hssi_common_pcs_pma_interface_sigdet_wait_counter),
				.sigdet_wait_counter_multi(hssi_common_pcs_pma_interface_sigdet_wait_counter_multi),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sim_mode(hssi_common_pcs_pma_interface_sim_mode),
				.spd_chg_rst_wait_cnt_en(hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en),
				.sup_mode(hssi_common_pcs_pma_interface_sup_mode),
				.testout_sel(hssi_common_pcs_pma_interface_testout_sel),
				.wait_clk_on_off_timer(hssi_common_pcs_pma_interface_wait_clk_on_off_timer),
				.wait_pipe_synchronizing(hssi_common_pcs_pma_interface_wait_pipe_synchronizing),
				.wait_send_syncp_fbkp(hssi_common_pcs_pma_interface_wait_send_syncp_fbkp)
			) inst_twentynm_hssi_common_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_common_pcs_pma_interface_blockselect),
				.int_pmaif_8g_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in),
				.int_pmaif_8g_eios_detected(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.int_pmaif_8g_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.int_pmaif_8g_power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.int_pmaif_g3_pcs_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in),
				.int_pmaif_pldif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pmaif_pldif_pcie_sw_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done),
				.int_pmaif_pldif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pmaif_pldif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pmaif_pldif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pmaif_pldif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pmaif_pldif_pma_reserved_in(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in),
				.int_pmaif_pldif_test_out(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out),
				.int_pmaif_pldif_testbus(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus),
				.pma_adapt_start(w_hssi_common_pcs_pma_interface_pma_adapt_start),
				.pma_atpg_los_en_n(w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n),
				.pma_csr_test_dis(w_hssi_common_pcs_pma_interface_pma_csr_test_dis),
				.pma_current_coeff(w_hssi_common_pcs_pma_interface_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_common_pcs_pma_interface_pma_current_rxpreset),
				.pma_early_eios(w_hssi_common_pcs_pma_interface_pma_early_eios),
				.pma_interface_select(w_hssi_common_pcs_pma_interface_pma_interface_select),
				.pma_ltd_b(w_hssi_common_pcs_pma_interface_pma_ltd_b),
				.pma_ltr(w_hssi_common_pcs_pma_interface_pma_ltr),
				.pma_nfrzdrv(w_hssi_common_pcs_pma_interface_pma_nfrzdrv),
				.pma_nrpi_freeze(w_hssi_common_pcs_pma_interface_pma_nrpi_freeze),
				.pma_pcie_switch(w_hssi_common_pcs_pma_interface_pma_pcie_switch),
				.pma_ppm_lock(w_hssi_common_pcs_pma_interface_pma_ppm_lock),
				.pma_reserved_out(w_hssi_common_pcs_pma_interface_pma_reserved_out),
				.pma_rs_lpbk_b(w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b),
				.pma_rx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup),
				.pma_scan_mode_n(w_hssi_common_pcs_pma_interface_pma_scan_mode_n),
				.pma_scan_shift_n(w_hssi_common_pcs_pma_interface_pma_scan_shift_n),
				.pma_tx_bitslip(w_hssi_common_pcs_pma_interface_pma_tx_bitslip),
				.pma_tx_bonding_rstb(w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb),
				.pma_tx_qpi_pulldn(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn),
				.pma_tx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup),
				.pma_tx_txdetectrx(w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx),
				.pmaif_bundling_out_down(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down),
				.pmaif_bundling_out_up(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_8g_current_coeff({w_hssi_pipe_gen1_2_current_coeff[17], w_hssi_pipe_gen1_2_current_coeff[16], w_hssi_pipe_gen1_2_current_coeff[15], w_hssi_pipe_gen1_2_current_coeff[14], w_hssi_pipe_gen1_2_current_coeff[13], w_hssi_pipe_gen1_2_current_coeff[12], w_hssi_pipe_gen1_2_current_coeff[11], w_hssi_pipe_gen1_2_current_coeff[10], w_hssi_pipe_gen1_2_current_coeff[9], w_hssi_pipe_gen1_2_current_coeff[8], w_hssi_pipe_gen1_2_current_coeff[7], w_hssi_pipe_gen1_2_current_coeff[6], w_hssi_pipe_gen1_2_current_coeff[5], w_hssi_pipe_gen1_2_current_coeff[4], w_hssi_pipe_gen1_2_current_coeff[3], w_hssi_pipe_gen1_2_current_coeff[2], w_hssi_pipe_gen1_2_current_coeff[1], w_hssi_pipe_gen1_2_current_coeff[0]}),
				.int_pmaif_8g_eios_det({w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0]}),
				.int_pmaif_8g_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.int_pmaif_8g_rev_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.int_pmaif_8g_tx_clk_out_gen3(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.int_pmaif_8g_txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				.int_pmaif_g3_eios_det({w_hssi_gen3_rx_pcs_ei_det_int, w_hssi_gen3_rx_pcs_ei_partial_det_int, w_hssi_gen3_rx_pcs_i_det_int}),
				.int_pmaif_g3_pma_current_coeff({w_hssi_pipe_gen3_pma_current_coeff[17], w_hssi_pipe_gen3_pma_current_coeff[16], w_hssi_pipe_gen3_pma_current_coeff[15], w_hssi_pipe_gen3_pma_current_coeff[14], w_hssi_pipe_gen3_pma_current_coeff[13], w_hssi_pipe_gen3_pma_current_coeff[12], w_hssi_pipe_gen3_pma_current_coeff[11], w_hssi_pipe_gen3_pma_current_coeff[10], w_hssi_pipe_gen3_pma_current_coeff[9], w_hssi_pipe_gen3_pma_current_coeff[8], w_hssi_pipe_gen3_pma_current_coeff[7], w_hssi_pipe_gen3_pma_current_coeff[6], w_hssi_pipe_gen3_pma_current_coeff[5], w_hssi_pipe_gen3_pma_current_coeff[4], w_hssi_pipe_gen3_pma_current_coeff[3], w_hssi_pipe_gen3_pma_current_coeff[2], w_hssi_pipe_gen3_pma_current_coeff[1], w_hssi_pipe_gen3_pma_current_coeff[0]}),
				.int_pmaif_g3_pma_current_rxpreset({w_hssi_pipe_gen3_pma_current_rxpreset[2], w_hssi_pipe_gen3_pma_current_rxpreset[1], w_hssi_pipe_gen3_pma_current_rxpreset[0]}),
				.int_pmaif_g3_pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.int_pmaif_g3_rev_lpbk(w_hssi_pipe_gen3_rev_lpbk_int),
				.int_pmaif_pldif_8g_tx_pld_rstn(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pmaif_pldif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pmaif_pldif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pmaif_pldif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pmaif_pldif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pmaif_pldif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pmaif_pldif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pmaif_pldif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pmaif_pldif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pmaif_pldif_pcie_switch({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0]}),
				.int_pmaif_pldif_pma_reserved_out({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0]}),
				.int_pmaif_pldif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pmaif_pldif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pmaif_pldif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pmaif_pldif_rate({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0]}),
				.int_pmaif_pldif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pmaif_pldif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pmaif_pldif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.int_pmaif_pldif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pmaif_pldif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pmaif_pldif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pmaif_pldif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pmaif_pldif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pmaif_pldif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.int_tx_dft_obsrv_clk({w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0]}),
				.iocsr_clk(in_iocsr_clk),
				.iocsr_config({in_iocsr_config[5], in_iocsr_config[4], in_iocsr_config[3], in_iocsr_config[2], in_iocsr_config[1], in_iocsr_config[0]}),
				.iocsr_rdy(in_iocsr_rdy),
				.iocsr_rdy_dly(in_iocsr_rdy_dly),
				.pma_adapt_done(in_pma_adapt_done),
				.pma_clklow(in_pma_clklow),
				.pma_fref(in_pma_fref),
				.pma_hclk(in_pma_hclk),
				.pma_pcie_sw_done({in_pma_pcie_sw_done[1], in_pma_pcie_sw_done[0]}),
				.pma_pfdmode_lock(in_pma_pfdmode_lock),
				.pma_reserved_in({in_pma_reserved_in[4], in_pma_reserved_in[3], in_pma_reserved_in[2], in_pma_reserved_in[1], in_pma_reserved_in[0]}),
				.pma_signal_det(in_pma_signal_det),
				.pma_testbus({in_pma_testbus[7], in_pma_testbus[6], in_pma_testbus[5], in_pma_testbus[4], in_pma_testbus[3], in_pma_testbus[2], in_pma_testbus[1], in_pma_testbus[0]}),
				.pmaif_bundling_in_down({in_bond_pmaif_in_bot[11], in_bond_pmaif_in_bot[10], in_bond_pmaif_in_bot[9], in_bond_pmaif_in_bot[8], in_bond_pmaif_in_bot[7], in_bond_pmaif_in_bot[6], in_bond_pmaif_in_bot[5], in_bond_pmaif_in_bot[4], in_bond_pmaif_in_bot[3], in_bond_pmaif_in_bot[2], in_bond_pmaif_in_bot[1], in_bond_pmaif_in_bot[0]}),
				.pmaif_bundling_in_up({in_bond_pmaif_in_top[11], in_bond_pmaif_in_top[10], in_bond_pmaif_in_top[9], in_bond_pmaif_in_top[8], in_bond_pmaif_in_top[7], in_bond_pmaif_in_top[6], in_bond_pmaif_in_top[5], in_bond_pmaif_in_top[4], in_bond_pmaif_in_top[3], in_bond_pmaif_in_top[2], in_bond_pmaif_in_top[1], in_bond_pmaif_in_top[0]}),
				.rx_pmaif_test_out({w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0]}),
				.rx_prbs_ver_test({w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0]}),
				.tx_prbs_gen_test({w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0]}),
				.uhsif_test_out_1({w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0]}),
				.uhsif_test_out_2({w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0]}),
				.uhsif_test_out_3({w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0]}),
				
				// UNUSED
				.int_pmaif_avmm_iocsr_clk(),
				.int_pmaif_avmm_iocsr_config(),
				.int_pmaif_avmm_iocsr_rdy(),
				.int_pmaif_avmm_iocsr_rdy_dly(),
				.int_pmaif_pldif_interface_select(),
				.pma_tx_pma_syncp(),
				.sta_pma_hclk_by2()
			);
		end // if generate
		else begin
				assign w_hssi_common_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19:0] = 20'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_pma_adapt_start = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_csr_test_dis = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pcs_pma_interface_pma_early_eios = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_interface_select[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltd_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltr = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nfrzdrv = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nrpi_freeze = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ppm_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_tx_bitslip = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx = in_pld_pma_txdetectrx;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11:0] = 12'b0;
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11:0] = 12'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pld_pcs_interface
			twentynm_hssi_common_pld_pcs_interface #(
				.dft_clk_out_en(hssi_common_pld_pcs_interface_dft_clk_out_en),
				.dft_clk_out_sel(hssi_common_pld_pcs_interface_dft_clk_out_sel),
				.hrdrstctrl_en(hssi_common_pld_pcs_interface_hrdrstctrl_en),
				.pcs_testbus_block_sel(hssi_common_pld_pcs_interface_pcs_testbus_block_sel),
				.reconfig_settings(hssi_common_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm4" )       //PARAM_HIDE
			) inst_twentynm_hssi_common_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_common_pld_pcs_interface_blockselect),
				.hip_cmn_clk(w_hssi_common_pld_pcs_interface_hip_cmn_clk),
				.hip_cmn_ctrl(w_hssi_common_pld_pcs_interface_hip_cmn_ctrl),
				.hip_iocsr_rdy(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy),
				.hip_iocsr_rdy_dly(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly),
				.hip_nfrzdrv(w_hssi_common_pld_pcs_interface_hip_nfrzdrv),
				.hip_npor(w_hssi_common_pld_pcs_interface_hip_npor),
				.hip_usermode(w_hssi_common_pld_pcs_interface_hip_usermode),
				.int_pldif_10g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.int_pldif_10g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.int_pldif_8g_eidleinfersel(w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel),
				.int_pldif_8g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.int_pldif_8g_refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.int_pldif_8g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.int_pldif_g3_current_coeff(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff),
				.int_pldif_g3_current_rxpreset(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset),
				.int_pldif_krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.int_pldif_krfec_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.int_pldif_krfec_scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				.int_pldif_mem_atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.int_pldif_mem_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.int_pldif_pmaif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pldif_pmaif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pldif_pmaif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pldif_pmaif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pldif_pmaif_eye_monitor(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor),
				.int_pldif_pmaif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pldif_pmaif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pldif_pmaif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pldif_pmaif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pldif_pmaif_pcie_switch(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch),
				.int_pldif_pmaif_pma_reserved_out(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out),
				.int_pldif_pmaif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pldif_pmaif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pldif_pmaif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pldif_pmaif_rate(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate),
				.int_pldif_pmaif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pldif_pmaif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pldif_pmaif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pldif_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_pldif_pmaif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pldif_pmaif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pldif_pmaif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pldif_pmaif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pldif_pmaif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pldif_pmaif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pldif_pmaif_uhsif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.pld_pma_adapt_done(w_hssi_common_pld_pcs_interface_pld_pma_adapt_done),
				.pld_pma_clklow(w_hssi_common_pld_pcs_interface_pld_pma_clklow),
				.pld_pma_fref(w_hssi_common_pld_pcs_interface_pld_pma_fref),
				.pld_pma_hclk(w_hssi_common_pld_pcs_interface_pld_pma_hclk),
				.pld_pma_pcie_sw_done(w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done),
				.pld_pma_pfdmode_lock(w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock),
				.pld_pma_reserved_in(w_hssi_common_pld_pcs_interface_pld_pma_reserved_in),
				.pld_pma_rx_detect_valid(w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid),
				.pld_pma_rx_found(w_hssi_common_pld_pcs_interface_pld_pma_rx_found),
				.pld_pma_rxpll_lock(w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock),
				.pld_pma_testbus(w_hssi_common_pld_pcs_interface_pld_pma_testbus),
				.pld_pmaif_mask_tx_pll(w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll),
				.pld_reserved_out(w_hssi_common_pld_pcs_interface_pld_reserved_out),
				.pld_test_data(w_hssi_common_pld_pcs_interface_pld_test_data),
				.pld_uhsif_lock(w_hssi_common_pld_pcs_interface_pld_uhsif_lock),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.int_pldif_10g_test_data({w_hssi_10g_tx_pcs_tx_test_data[19], w_hssi_10g_tx_pcs_tx_test_data[18], w_hssi_10g_tx_pcs_tx_test_data[17], w_hssi_10g_tx_pcs_tx_test_data[16], w_hssi_10g_tx_pcs_tx_test_data[15], w_hssi_10g_tx_pcs_tx_test_data[14], w_hssi_10g_tx_pcs_tx_test_data[13], w_hssi_10g_tx_pcs_tx_test_data[12], w_hssi_10g_tx_pcs_tx_test_data[11], w_hssi_10g_tx_pcs_tx_test_data[10], w_hssi_10g_tx_pcs_tx_test_data[9], w_hssi_10g_tx_pcs_tx_test_data[8], w_hssi_10g_tx_pcs_tx_test_data[7], w_hssi_10g_tx_pcs_tx_test_data[6], w_hssi_10g_tx_pcs_tx_test_data[5], w_hssi_10g_tx_pcs_tx_test_data[4], w_hssi_10g_tx_pcs_tx_test_data[3], w_hssi_10g_tx_pcs_tx_test_data[2], w_hssi_10g_tx_pcs_tx_test_data[1], w_hssi_10g_tx_pcs_tx_test_data[0]}),
				.int_pldif_10g_tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.int_pldif_8g_chnl_test_bus_out({w_hssi_8g_rx_pcs_chnl_test_bus_out[19], w_hssi_8g_rx_pcs_chnl_test_bus_out[18], w_hssi_8g_rx_pcs_chnl_test_bus_out[17], w_hssi_8g_rx_pcs_chnl_test_bus_out[16], w_hssi_8g_rx_pcs_chnl_test_bus_out[15], w_hssi_8g_rx_pcs_chnl_test_bus_out[14], w_hssi_8g_rx_pcs_chnl_test_bus_out[13], w_hssi_8g_rx_pcs_chnl_test_bus_out[12], w_hssi_8g_rx_pcs_chnl_test_bus_out[11], w_hssi_8g_rx_pcs_chnl_test_bus_out[10], w_hssi_8g_rx_pcs_chnl_test_bus_out[9], w_hssi_8g_rx_pcs_chnl_test_bus_out[8], w_hssi_8g_rx_pcs_chnl_test_bus_out[7], w_hssi_8g_rx_pcs_chnl_test_bus_out[6], w_hssi_8g_rx_pcs_chnl_test_bus_out[5], w_hssi_8g_rx_pcs_chnl_test_bus_out[4], w_hssi_8g_rx_pcs_chnl_test_bus_out[3], w_hssi_8g_rx_pcs_chnl_test_bus_out[2], w_hssi_8g_rx_pcs_chnl_test_bus_out[1], w_hssi_8g_rx_pcs_chnl_test_bus_out[0]}),
				.int_pldif_8g_rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.int_pldif_8g_tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.int_pldif_g3_test_out({w_hssi_pipe_gen3_test_out[19], w_hssi_pipe_gen3_test_out[18], w_hssi_pipe_gen3_test_out[17], w_hssi_pipe_gen3_test_out[16], w_hssi_pipe_gen3_test_out[15], w_hssi_pipe_gen3_test_out[14], w_hssi_pipe_gen3_test_out[13], w_hssi_pipe_gen3_test_out[12], w_hssi_pipe_gen3_test_out[11], w_hssi_pipe_gen3_test_out[10], w_hssi_pipe_gen3_test_out[9], w_hssi_pipe_gen3_test_out[8], w_hssi_pipe_gen3_test_out[7], w_hssi_pipe_gen3_test_out[6], w_hssi_pipe_gen3_test_out[5], w_hssi_pipe_gen3_test_out[4], w_hssi_pipe_gen3_test_out[3], w_hssi_pipe_gen3_test_out[2], w_hssi_pipe_gen3_test_out[1], w_hssi_pipe_gen3_test_out[0]}),
				.int_pldif_krfec_test_data({w_hssi_krfec_tx_pcs_tx_test_data[19], w_hssi_krfec_tx_pcs_tx_test_data[18], w_hssi_krfec_tx_pcs_tx_test_data[17], w_hssi_krfec_tx_pcs_tx_test_data[16], w_hssi_krfec_tx_pcs_tx_test_data[15], w_hssi_krfec_tx_pcs_tx_test_data[14], w_hssi_krfec_tx_pcs_tx_test_data[13], w_hssi_krfec_tx_pcs_tx_test_data[12], w_hssi_krfec_tx_pcs_tx_test_data[11], w_hssi_krfec_tx_pcs_tx_test_data[10], w_hssi_krfec_tx_pcs_tx_test_data[9], w_hssi_krfec_tx_pcs_tx_test_data[8], w_hssi_krfec_tx_pcs_tx_test_data[7], w_hssi_krfec_tx_pcs_tx_test_data[6], w_hssi_krfec_tx_pcs_tx_test_data[5], w_hssi_krfec_tx_pcs_tx_test_data[4], w_hssi_krfec_tx_pcs_tx_test_data[3], w_hssi_krfec_tx_pcs_tx_test_data[2], w_hssi_krfec_tx_pcs_tx_test_data[1], w_hssi_krfec_tx_pcs_tx_test_data[0]}),
				.int_pldif_pmaif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pldif_pmaif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pldif_pmaif_pcie_sw_done({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0]}),
				.int_pldif_pmaif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pldif_pmaif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pldif_pmaif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pldif_pmaif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pldif_pmaif_pma_reserved_in({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0]}),
				.int_pldif_pmaif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pldif_pmaif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_test_out({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0]}),
				.int_pldif_pmaif_testbus({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0]}),
				.int_pldif_pmaif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.pld_8g_eidleinfersel({in_pld_8g_eidleinfersel[2], in_pld_8g_eidleinfersel[1], in_pld_8g_eidleinfersel[0]}),
				.pld_8g_refclk_dig2(in_pld_8g_refclk_dig2),
				.pld_atpg_los_en_n(in_pld_atpg_los_en_n),
				.pld_g3_current_coeff({in_pld_g3_current_coeff[17], in_pld_g3_current_coeff[16], in_pld_g3_current_coeff[15], in_pld_g3_current_coeff[14], in_pld_g3_current_coeff[13], in_pld_g3_current_coeff[12], in_pld_g3_current_coeff[11], in_pld_g3_current_coeff[10], in_pld_g3_current_coeff[9], in_pld_g3_current_coeff[8], in_pld_g3_current_coeff[7], in_pld_g3_current_coeff[6], in_pld_g3_current_coeff[5], in_pld_g3_current_coeff[4], in_pld_g3_current_coeff[3], in_pld_g3_current_coeff[2], in_pld_g3_current_coeff[1], in_pld_g3_current_coeff[0]}),
				.pld_g3_current_rxpreset({in_pld_g3_current_rxpreset[2], in_pld_g3_current_rxpreset[1], in_pld_g3_current_rxpreset[0]}),
				.pld_ltr(in_pld_ltr),
				.pld_mem_krfec_atpg_rst_n(in_pld_mem_krfec_atpg_rst_n),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pcs_refclk_dig(in_pld_pcs_refclk_dig),
				.pld_pma_adapt_start(in_pld_pma_adapt_start),
				.pld_pma_csr_test_dis(in_pld_pma_csr_test_dis),
				.pld_pma_early_eios(in_pld_pma_early_eios),
				.pld_pma_eye_monitor({in_pld_pma_eye_monitor[5], in_pld_pma_eye_monitor[4], in_pld_pma_eye_monitor[3], in_pld_pma_eye_monitor[2], in_pld_pma_eye_monitor[1], in_pld_pma_eye_monitor[0]}),
				.pld_pma_ltd_b(in_pld_pma_ltd_b),
				.pld_pma_nrpi_freeze(in_pld_pma_nrpi_freeze),
				.pld_pma_pcie_switch({in_pld_pma_pcie_switch[1], in_pld_pma_pcie_switch[0]}),
				.pld_pma_ppm_lock(in_pld_pma_ppm_lock),
				.pld_pma_reserved_out({in_pld_pma_reserved_out[4], in_pld_pma_reserved_out[3], in_pld_pma_reserved_out[2], in_pld_pma_reserved_out[1], in_pld_pma_reserved_out[0]}),
				.pld_pma_rs_lpbk_b(in_pld_pma_rs_lpbk_b),
				.pld_pma_rx_qpi_pullup(in_pld_pma_rx_qpi_pullup),
				.pld_pma_tx_bitslip(in_pld_pma_tx_bitslip),
				.pld_pma_tx_bonding_rstb(in_pld_pma_tx_bonding_rstb),
				.pld_pma_tx_qpi_pulldn(in_pld_pma_tx_qpi_pulldn),
				.pld_pma_tx_qpi_pullup(in_pld_pma_tx_qpi_pullup),
				.pld_pma_txdetectrx(in_pld_pma_txdetectrx),
				.pld_rate({in_pld_rate[1], in_pld_rate[0]}),
				.pld_reserved_in({in_pld_reserved_in[9], in_pld_reserved_in[8], in_pld_reserved_in[7], in_pld_reserved_in[6], in_pld_reserved_in[5], in_pld_reserved_in[4], in_pld_reserved_in[3], in_pld_reserved_in[2], in_pld_reserved_in[1], in_pld_reserved_in[0]}),
				.pld_scan_mode_n(in_pld_scan_mode_n),
				.pld_scan_shift_n(in_pld_scan_shift_n),
				
				// UNUSED
				.int_pldif_8g_ltr(),
				.int_pldif_avmm_pld_avmm1_request(),
				.int_pldif_avmm_pld_avmm2_request(),
				.int_pldif_avmm_refclk_dig_en(),
				.int_pldif_g3_scan_mode_n(),
				.pld_8g_eidleinfersel_fifo(),
				.pld_8g_eidleinfersel_reg(),
				.pld_partial_reconfig_fifo(),
				.pld_partial_reconfig_rx_div_by_2_rxclk_wire(),
				.pld_partial_reconfig_rx_div_by_2_txclk_wire(),
				.pld_partial_reconfig_rxclk_reg(),
				.pld_partial_reconfig_tx_div_by_2_wire(),
				.pld_partial_reconfig_txclk_reg(),
				.pld_rate_reg(),
				.pld_test_data_reg()
			);
		end // if generate
		else begin
				assign w_hssi_common_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_clk[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_npor = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_usermode = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2 = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_adapt_done = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_clklow = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_fref = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_hclk = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_found = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_testbus[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_reserved_out[9:0] = 10'b0;
				assign w_hssi_common_pld_pcs_interface_pld_test_data[19:0] = 20'b0;
				assign w_hssi_common_pld_pcs_interface_pld_uhsif_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_scan_mode_n = 1'b1;		// Override default tieoff
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_rx_pcs
			twentynm_hssi_fifo_rx_pcs #(
				.double_read_mode(hssi_fifo_rx_pcs_double_read_mode),
				.prot_mode(hssi_fifo_rx_pcs_prot_mode),
				.silicon_rev( "20nm4" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_rx_pcs_blockselect),
				.data_out2_10g(w_hssi_fifo_rx_pcs_data_out2_10g),
				.data_out2_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp),
				.data_out_10g(w_hssi_fifo_rx_pcs_data_out_10g),
				.data_out_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out_8g_clock_comp),
				.data_out_8g_phase_comp(w_hssi_fifo_rx_pcs_data_out_8g_phase_comp),
				.data_out_gen3(w_hssi_fifo_rx_pcs_data_out_gen3),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_data[73], w_hssi_10g_rx_pcs_rx_fifo_wr_data[72], w_hssi_10g_rx_pcs_rx_fifo_wr_data[71], w_hssi_10g_rx_pcs_rx_fifo_wr_data[70], w_hssi_10g_rx_pcs_rx_fifo_wr_data[69], w_hssi_10g_rx_pcs_rx_fifo_wr_data[68], w_hssi_10g_rx_pcs_rx_fifo_wr_data[67], w_hssi_10g_rx_pcs_rx_fifo_wr_data[66], w_hssi_10g_rx_pcs_rx_fifo_wr_data[65], w_hssi_10g_rx_pcs_rx_fifo_wr_data[64], w_hssi_10g_rx_pcs_rx_fifo_wr_data[63], w_hssi_10g_rx_pcs_rx_fifo_wr_data[62], w_hssi_10g_rx_pcs_rx_fifo_wr_data[61], w_hssi_10g_rx_pcs_rx_fifo_wr_data[60], w_hssi_10g_rx_pcs_rx_fifo_wr_data[59], w_hssi_10g_rx_pcs_rx_fifo_wr_data[58], w_hssi_10g_rx_pcs_rx_fifo_wr_data[57], w_hssi_10g_rx_pcs_rx_fifo_wr_data[56], w_hssi_10g_rx_pcs_rx_fifo_wr_data[55], w_hssi_10g_rx_pcs_rx_fifo_wr_data[54], w_hssi_10g_rx_pcs_rx_fifo_wr_data[53], w_hssi_10g_rx_pcs_rx_fifo_wr_data[52], w_hssi_10g_rx_pcs_rx_fifo_wr_data[51], w_hssi_10g_rx_pcs_rx_fifo_wr_data[50], w_hssi_10g_rx_pcs_rx_fifo_wr_data[49], w_hssi_10g_rx_pcs_rx_fifo_wr_data[48], w_hssi_10g_rx_pcs_rx_fifo_wr_data[47], w_hssi_10g_rx_pcs_rx_fifo_wr_data[46], w_hssi_10g_rx_pcs_rx_fifo_wr_data[45], w_hssi_10g_rx_pcs_rx_fifo_wr_data[44], w_hssi_10g_rx_pcs_rx_fifo_wr_data[43], w_hssi_10g_rx_pcs_rx_fifo_wr_data[42], w_hssi_10g_rx_pcs_rx_fifo_wr_data[41], w_hssi_10g_rx_pcs_rx_fifo_wr_data[40], w_hssi_10g_rx_pcs_rx_fifo_wr_data[39], w_hssi_10g_rx_pcs_rx_fifo_wr_data[38], w_hssi_10g_rx_pcs_rx_fifo_wr_data[37], w_hssi_10g_rx_pcs_rx_fifo_wr_data[36], w_hssi_10g_rx_pcs_rx_fifo_wr_data[35], w_hssi_10g_rx_pcs_rx_fifo_wr_data[34], w_hssi_10g_rx_pcs_rx_fifo_wr_data[33], w_hssi_10g_rx_pcs_rx_fifo_wr_data[32], w_hssi_10g_rx_pcs_rx_fifo_wr_data[31], w_hssi_10g_rx_pcs_rx_fifo_wr_data[30], w_hssi_10g_rx_pcs_rx_fifo_wr_data[29], w_hssi_10g_rx_pcs_rx_fifo_wr_data[28], w_hssi_10g_rx_pcs_rx_fifo_wr_data[27], w_hssi_10g_rx_pcs_rx_fifo_wr_data[26], w_hssi_10g_rx_pcs_rx_fifo_wr_data[25], w_hssi_10g_rx_pcs_rx_fifo_wr_data[24], w_hssi_10g_rx_pcs_rx_fifo_wr_data[23], w_hssi_10g_rx_pcs_rx_fifo_wr_data[22], w_hssi_10g_rx_pcs_rx_fifo_wr_data[21], w_hssi_10g_rx_pcs_rx_fifo_wr_data[20], w_hssi_10g_rx_pcs_rx_fifo_wr_data[19], w_hssi_10g_rx_pcs_rx_fifo_wr_data[18], w_hssi_10g_rx_pcs_rx_fifo_wr_data[17], w_hssi_10g_rx_pcs_rx_fifo_wr_data[16], w_hssi_10g_rx_pcs_rx_fifo_wr_data[15], w_hssi_10g_rx_pcs_rx_fifo_wr_data[14], w_hssi_10g_rx_pcs_rx_fifo_wr_data[13], w_hssi_10g_rx_pcs_rx_fifo_wr_data[12], w_hssi_10g_rx_pcs_rx_fifo_wr_data[11], w_hssi_10g_rx_pcs_rx_fifo_wr_data[10], w_hssi_10g_rx_pcs_rx_fifo_wr_data[9], w_hssi_10g_rx_pcs_rx_fifo_wr_data[8], w_hssi_10g_rx_pcs_rx_fifo_wr_data[7], w_hssi_10g_rx_pcs_rx_fifo_wr_data[6], w_hssi_10g_rx_pcs_rx_fifo_wr_data[5], w_hssi_10g_rx_pcs_rx_fifo_wr_data[4], w_hssi_10g_rx_pcs_rx_fifo_wr_data[3], w_hssi_10g_rx_pcs_rx_fifo_wr_data[2], w_hssi_10g_rx_pcs_rx_fifo_wr_data[1], w_hssi_10g_rx_pcs_rx_fifo_wr_data[0]}),
				.data_in_8g_clock_comp({w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0]}),
				.data_in_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr2_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0]}),
				.rd_ptr2_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0]}),
				.rd_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0]}),
				.rd_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.wr_clk_8g_clock_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_8g_clock_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.wr_en_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.wr_en_8g_clock_comp(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_en_8g_phase_comp(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.wr_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0]}),
				.wr_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0]}),
				.wr_rst_n_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.wr_rst_n_8g_clock_comp(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_n_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_rx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79:0] = 80'b0;
				assign w_hssi_fifo_rx_pcs_data_out_gen3[39:0] = 40'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_tx_pcs
			twentynm_hssi_fifo_tx_pcs #(
				.double_write_mode(hssi_fifo_tx_pcs_double_write_mode),
				.prot_mode(hssi_fifo_tx_pcs_prot_mode),
				.silicon_rev( "20nm4" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_tx_pcs_blockselect),
				.data_out_10g(w_hssi_fifo_tx_pcs_data_out_10g),
				.data_out_8g_phase_comp(w_hssi_fifo_tx_pcs_data_out_8g_phase_comp),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in2_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0]}),
				.data_in_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_en_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.wr_en_8g_phase_comp(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0]}),
				.wr_rst_n_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_tx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_tx_pcs_data_out_10g[72:0] = 73'b0;
				assign w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63:0] = 64'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_rx_pcs
			twentynm_hssi_gen3_rx_pcs #(
				.block_sync(hssi_gen3_rx_pcs_block_sync),
				.block_sync_sm(hssi_gen3_rx_pcs_block_sync_sm),
				.cdr_ctrl_force_unalgn(hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn),
				.lpbk_force(hssi_gen3_rx_pcs_lpbk_force),
				.mode(hssi_gen3_rx_pcs_mode),
				.rate_match_fifo(hssi_gen3_rx_pcs_rate_match_fifo),
				.rate_match_fifo_latency(hssi_gen3_rx_pcs_rate_match_fifo_latency),
				.reconfig_settings(hssi_gen3_rx_pcs_reconfig_settings),
				.reverse_lpbk(hssi_gen3_rx_pcs_reverse_lpbk),
				.rx_b4gb_par_lpbk(hssi_gen3_rx_pcs_rx_b4gb_par_lpbk),
				.rx_force_balign(hssi_gen3_rx_pcs_rx_force_balign),
				.rx_ins_del_one_skip(hssi_gen3_rx_pcs_rx_ins_del_one_skip),
				.rx_num_fixed_pat(hssi_gen3_rx_pcs_rx_num_fixed_pat),
				.rx_test_out_sel(hssi_gen3_rx_pcs_rx_test_out_sel),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_rx_pcs_sup_mode)
			) inst_twentynm_hssi_gen3_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_rx_pcs_avmmreaddata),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.blk_start(w_hssi_gen3_rx_pcs_blk_start),
				.blockselect(w_hssi_gen3_rx_pcs_blockselect),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.data_out(w_hssi_gen3_rx_pcs_data_out),
				.data_valid(w_hssi_gen3_rx_pcs_data_valid),
				.ei_det_int(w_hssi_gen3_rx_pcs_ei_det_int),
				.ei_partial_det_int(w_hssi_gen3_rx_pcs_ei_partial_det_int),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.i_det_int(w_hssi_gen3_rx_pcs_i_det_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data(w_hssi_gen3_rx_pcs_lpbk_data),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.mem_rx_fifo_rd_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr),
				.mem_rx_fifo_wr_clk(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.mem_rx_fifo_wr_data(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data),
				.mem_rx_fifo_wr_en(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.mem_rx_fifo_wr_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr),
				.mem_rx_fifo_wr_rst_n(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_test_out(w_hssi_gen3_rx_pcs_rx_test_out),
				.sync_hdr(w_hssi_gen3_rx_pcs_sync_hdr),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0]}),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.mem_rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_gen3[39], w_hssi_fifo_rx_pcs_data_out_gen3[38], w_hssi_fifo_rx_pcs_data_out_gen3[37], w_hssi_fifo_rx_pcs_data_out_gen3[36], w_hssi_fifo_rx_pcs_data_out_gen3[35], w_hssi_fifo_rx_pcs_data_out_gen3[34], w_hssi_fifo_rx_pcs_data_out_gen3[33], w_hssi_fifo_rx_pcs_data_out_gen3[32], w_hssi_fifo_rx_pcs_data_out_gen3[31], w_hssi_fifo_rx_pcs_data_out_gen3[30], w_hssi_fifo_rx_pcs_data_out_gen3[29], w_hssi_fifo_rx_pcs_data_out_gen3[28], w_hssi_fifo_rx_pcs_data_out_gen3[27], w_hssi_fifo_rx_pcs_data_out_gen3[26], w_hssi_fifo_rx_pcs_data_out_gen3[25], w_hssi_fifo_rx_pcs_data_out_gen3[24], w_hssi_fifo_rx_pcs_data_out_gen3[23], w_hssi_fifo_rx_pcs_data_out_gen3[22], w_hssi_fifo_rx_pcs_data_out_gen3[21], w_hssi_fifo_rx_pcs_data_out_gen3[20], w_hssi_fifo_rx_pcs_data_out_gen3[19], w_hssi_fifo_rx_pcs_data_out_gen3[18], w_hssi_fifo_rx_pcs_data_out_gen3[17], w_hssi_fifo_rx_pcs_data_out_gen3[16], w_hssi_fifo_rx_pcs_data_out_gen3[15], w_hssi_fifo_rx_pcs_data_out_gen3[14], w_hssi_fifo_rx_pcs_data_out_gen3[13], w_hssi_fifo_rx_pcs_data_out_gen3[12], w_hssi_fifo_rx_pcs_data_out_gen3[11], w_hssi_fifo_rx_pcs_data_out_gen3[10], w_hssi_fifo_rx_pcs_data_out_gen3[9], w_hssi_fifo_rx_pcs_data_out_gen3[8], w_hssi_fifo_rx_pcs_data_out_gen3[7], w_hssi_fifo_rx_pcs_data_out_gen3[6], w_hssi_fifo_rx_pcs_data_out_gen3[5], w_hssi_fifo_rx_pcs_data_out_gen3[4], w_hssi_fifo_rx_pcs_data_out_gen3[3], w_hssi_fifo_rx_pcs_data_out_gen3[2], w_hssi_fifo_rx_pcs_data_out_gen3[1], w_hssi_fifo_rx_pcs_data_out_gen3[0]}),
				.par_lpbk_b4gb_in({w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0]}),
				.par_lpbk_in({w_hssi_gen3_tx_pcs_par_lpbk_out[31], w_hssi_gen3_tx_pcs_par_lpbk_out[30], w_hssi_gen3_tx_pcs_par_lpbk_out[29], w_hssi_gen3_tx_pcs_par_lpbk_out[28], w_hssi_gen3_tx_pcs_par_lpbk_out[27], w_hssi_gen3_tx_pcs_par_lpbk_out[26], w_hssi_gen3_tx_pcs_par_lpbk_out[25], w_hssi_gen3_tx_pcs_par_lpbk_out[24], w_hssi_gen3_tx_pcs_par_lpbk_out[23], w_hssi_gen3_tx_pcs_par_lpbk_out[22], w_hssi_gen3_tx_pcs_par_lpbk_out[21], w_hssi_gen3_tx_pcs_par_lpbk_out[20], w_hssi_gen3_tx_pcs_par_lpbk_out[19], w_hssi_gen3_tx_pcs_par_lpbk_out[18], w_hssi_gen3_tx_pcs_par_lpbk_out[17], w_hssi_gen3_tx_pcs_par_lpbk_out[16], w_hssi_gen3_tx_pcs_par_lpbk_out[15], w_hssi_gen3_tx_pcs_par_lpbk_out[14], w_hssi_gen3_tx_pcs_par_lpbk_out[13], w_hssi_gen3_tx_pcs_par_lpbk_out[12], w_hssi_gen3_tx_pcs_par_lpbk_out[11], w_hssi_gen3_tx_pcs_par_lpbk_out[10], w_hssi_gen3_tx_pcs_par_lpbk_out[9], w_hssi_gen3_tx_pcs_par_lpbk_out[8], w_hssi_gen3_tx_pcs_par_lpbk_out[7], w_hssi_gen3_tx_pcs_par_lpbk_out[6], w_hssi_gen3_tx_pcs_par_lpbk_out[5], w_hssi_gen3_tx_pcs_par_lpbk_out[4], w_hssi_gen3_tx_pcs_par_lpbk_out[3], w_hssi_gen3_tx_pcs_par_lpbk_out[2], w_hssi_gen3_tx_pcs_par_lpbk_out[1], w_hssi_gen3_tx_pcs_par_lpbk_out[0]}),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.rcvd_clk(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_pma_clk(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.rxpolarity(w_hssi_pipe_gen3_rxpolarity_int),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.sync_sm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.txdatak_in({w_hssi_pipe_gen3_txdatak_int[3], w_hssi_pipe_gen3_txdatak_int[2], w_hssi_pipe_gen3_txdatak_int[1], w_hssi_pipe_gen3_txdatak_int[0]}),
				
				// UNUSED
				.blk_lockd_int(),
				.skp_det_int()
			);
		end // if generate
		else begin
				assign w_hssi_gen3_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_rx_pcs_blk_algnd_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_delete_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_insert_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_overfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_undfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_rx_pcs_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_partial_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_err_decode_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_i_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data[33:0] = 34'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39:0] = 40'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_rx_test_out[19:0] = 20'b0;
				assign w_hssi_gen3_rx_pcs_sync_hdr[1:0] = 2'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_tx_pcs
			twentynm_hssi_gen3_tx_pcs #(
				.mode(hssi_gen3_tx_pcs_mode),
				.reverse_lpbk(hssi_gen3_tx_pcs_reverse_lpbk),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_tx_pcs_sup_mode),
				.tx_bitslip(hssi_gen3_tx_pcs_tx_bitslip),
				.tx_gbox_byp(hssi_gen3_tx_pcs_tx_gbox_byp)
			) inst_twentynm_hssi_gen3_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_gen3_tx_pcs_blockselect),
				.data_out(w_hssi_gen3_tx_pcs_data_out),
				.par_lpbk_b4gb_out(w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out),
				.par_lpbk_out(w_hssi_gen3_tx_pcs_par_lpbk_out),
				.tx_test_out(w_hssi_gen3_tx_pcs_tx_test_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_start_in(w_hssi_pipe_gen3_tx_blk_start_int),
				.data_in({w_hssi_pipe_gen3_txdata_int[31], w_hssi_pipe_gen3_txdata_int[30], w_hssi_pipe_gen3_txdata_int[29], w_hssi_pipe_gen3_txdata_int[28], w_hssi_pipe_gen3_txdata_int[27], w_hssi_pipe_gen3_txdata_int[26], w_hssi_pipe_gen3_txdata_int[25], w_hssi_pipe_gen3_txdata_int[24], w_hssi_pipe_gen3_txdata_int[23], w_hssi_pipe_gen3_txdata_int[22], w_hssi_pipe_gen3_txdata_int[21], w_hssi_pipe_gen3_txdata_int[20], w_hssi_pipe_gen3_txdata_int[19], w_hssi_pipe_gen3_txdata_int[18], w_hssi_pipe_gen3_txdata_int[17], w_hssi_pipe_gen3_txdata_int[16], w_hssi_pipe_gen3_txdata_int[15], w_hssi_pipe_gen3_txdata_int[14], w_hssi_pipe_gen3_txdata_int[13], w_hssi_pipe_gen3_txdata_int[12], w_hssi_pipe_gen3_txdata_int[11], w_hssi_pipe_gen3_txdata_int[10], w_hssi_pipe_gen3_txdata_int[9], w_hssi_pipe_gen3_txdata_int[8], w_hssi_pipe_gen3_txdata_int[7], w_hssi_pipe_gen3_txdata_int[6], w_hssi_pipe_gen3_txdata_int[5], w_hssi_pipe_gen3_txdata_int[4], w_hssi_pipe_gen3_txdata_int[3], w_hssi_pipe_gen3_txdata_int[2], w_hssi_pipe_gen3_txdata_int[1], w_hssi_pipe_gen3_txdata_int[0]}),
				.data_valid(w_hssi_pipe_gen3_txdataskip_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data_in({w_hssi_gen3_rx_pcs_lpbk_data[33], w_hssi_gen3_rx_pcs_lpbk_data[32], w_hssi_gen3_rx_pcs_lpbk_data[31], w_hssi_gen3_rx_pcs_lpbk_data[30], w_hssi_gen3_rx_pcs_lpbk_data[29], w_hssi_gen3_rx_pcs_lpbk_data[28], w_hssi_gen3_rx_pcs_lpbk_data[27], w_hssi_gen3_rx_pcs_lpbk_data[26], w_hssi_gen3_rx_pcs_lpbk_data[25], w_hssi_gen3_rx_pcs_lpbk_data[24], w_hssi_gen3_rx_pcs_lpbk_data[23], w_hssi_gen3_rx_pcs_lpbk_data[22], w_hssi_gen3_rx_pcs_lpbk_data[21], w_hssi_gen3_rx_pcs_lpbk_data[20], w_hssi_gen3_rx_pcs_lpbk_data[19], w_hssi_gen3_rx_pcs_lpbk_data[18], w_hssi_gen3_rx_pcs_lpbk_data[17], w_hssi_gen3_rx_pcs_lpbk_data[16], w_hssi_gen3_rx_pcs_lpbk_data[15], w_hssi_gen3_rx_pcs_lpbk_data[14], w_hssi_gen3_rx_pcs_lpbk_data[13], w_hssi_gen3_rx_pcs_lpbk_data[12], w_hssi_gen3_rx_pcs_lpbk_data[11], w_hssi_gen3_rx_pcs_lpbk_data[10], w_hssi_gen3_rx_pcs_lpbk_data[9], w_hssi_gen3_rx_pcs_lpbk_data[8], w_hssi_gen3_rx_pcs_lpbk_data[7], w_hssi_gen3_rx_pcs_lpbk_data[6], w_hssi_gen3_rx_pcs_lpbk_data[5], w_hssi_gen3_rx_pcs_lpbk_data[4], w_hssi_gen3_rx_pcs_lpbk_data[3], w_hssi_gen3_rx_pcs_lpbk_data[2], w_hssi_gen3_rx_pcs_lpbk_data[1], w_hssi_gen3_rx_pcs_lpbk_data[0]}),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.sync_in({w_hssi_pipe_gen3_tx_sync_hdr_int[1], w_hssi_pipe_gen3_tx_sync_hdr_int[0]}),
				.tx_pma_clk(w_hssi_8g_tx_pcs_clk_out_gen3),
				.tx_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn)
			);
		end // if generate
		else begin
				assign w_hssi_gen3_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_tx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_tx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35:0] = 36'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_tx_test_out[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_rx_pcs
			twentynm_hssi_krfec_rx_pcs #(
				.blksync_cor_en(hssi_krfec_rx_pcs_blksync_cor_en),
				.bypass_gb(hssi_krfec_rx_pcs_bypass_gb),
				.clr_ctrl(hssi_krfec_rx_pcs_clr_ctrl),
				.ctrl_bit_reverse(hssi_krfec_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_rx_pcs_data_bit_reverse),
				.dv_start(hssi_krfec_rx_pcs_dv_start),
				.err_mark_type(hssi_krfec_rx_pcs_err_mark_type),
				.error_marking_en(hssi_krfec_rx_pcs_error_marking_en),
				.low_latency_en(hssi_krfec_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_krfec_rx_pcs_lpbk_mode),
				.parity_invalid_enum(hssi_krfec_rx_pcs_parity_invalid_enum),
				.parity_valid_num(hssi_krfec_rx_pcs_parity_valid_num),
				.pipeln_blksync(hssi_krfec_rx_pcs_pipeln_blksync),
				.pipeln_descrm(hssi_krfec_rx_pcs_pipeln_descrm),
				.pipeln_errcorrect(hssi_krfec_rx_pcs_pipeln_errcorrect),
				.pipeln_errtrap_ind(hssi_krfec_rx_pcs_pipeln_errtrap_ind),
				.pipeln_errtrap_lfsr(hssi_krfec_rx_pcs_pipeln_errtrap_lfsr),
				.pipeln_errtrap_loc(hssi_krfec_rx_pcs_pipeln_errtrap_loc),
				.pipeln_errtrap_pat(hssi_krfec_rx_pcs_pipeln_errtrap_pat),
				.pipeln_gearbox(hssi_krfec_rx_pcs_pipeln_gearbox),
				.pipeln_syndrm(hssi_krfec_rx_pcs_pipeln_syndrm),
				.pipeln_trans_dec(hssi_krfec_rx_pcs_pipeln_trans_dec),
				.prot_mode(hssi_krfec_rx_pcs_prot_mode),
				.receive_order(hssi_krfec_rx_pcs_receive_order),
				.reconfig_settings(hssi_krfec_rx_pcs_reconfig_settings),
				.rx_testbus_sel(hssi_krfec_rx_pcs_rx_testbus_sel),
				.signal_ok_en(hssi_krfec_rx_pcs_signal_ok_en),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_rx_pcs_sup_mode)
			) inst_twentynm_hssi_krfec_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_rx_pcs_blockselect),
				.rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.rx_control_out(w_hssi_krfec_rx_pcs_rx_control_out),
				.rx_data_out(w_hssi_krfec_rx_pcs_rx_data_out),
				.rx_data_status(w_hssi_krfec_rx_pcs_rx_data_status),
				.rx_data_valid_out(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.rx_signal_ok_out(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.rx_data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0]}),
				.rx_krfec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_krfec_reg(),
				.pld_10g_krfec_rx_blk_lock_krfec_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg(),
				.pld_10g_krfec_rx_frame_krfec_reg(),
				.pld_10g_krfec_rx_frame_krfec_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_rx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_block_lock = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_control_out[9:0] = 10'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_status[1:0] = 2'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_valid_out = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_frame = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_signal_ok_out = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_tx_pcs
			twentynm_hssi_krfec_tx_pcs #(
				.burst_err(hssi_krfec_tx_pcs_burst_err),
				.burst_err_len(hssi_krfec_tx_pcs_burst_err_len),
				.ctrl_bit_reverse(hssi_krfec_tx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_tx_pcs_data_bit_reverse),
				.enc_frame_query(hssi_krfec_tx_pcs_enc_frame_query),
				.low_latency_en(hssi_krfec_tx_pcs_low_latency_en),
				.pipeln_encoder(hssi_krfec_tx_pcs_pipeln_encoder),
				.pipeln_scrambler(hssi_krfec_tx_pcs_pipeln_scrambler),
				.prot_mode(hssi_krfec_tx_pcs_prot_mode),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_tx_pcs_sup_mode),
				.transcode_err(hssi_krfec_tx_pcs_transcode_err),
				.transmit_order(hssi_krfec_tx_pcs_transmit_order),
				.tx_testbus_sel(hssi_krfec_tx_pcs_tx_testbus_sel)
			) inst_twentynm_hssi_krfec_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_tx_pcs_blockselect),
				.tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.tx_data_out(w_hssi_krfec_tx_pcs_tx_data_out),
				.tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.tx_test_data(w_hssi_krfec_tx_pcs_tx_test_data),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.tx_control_in({w_hssi_10g_tx_pcs_tx_control_out_krfec[8], w_hssi_10g_tx_pcs_tx_control_out_krfec[7], w_hssi_10g_tx_pcs_tx_control_out_krfec[6], w_hssi_10g_tx_pcs_tx_control_out_krfec[5], w_hssi_10g_tx_pcs_tx_control_out_krfec[4], w_hssi_10g_tx_pcs_tx_control_out_krfec[3], w_hssi_10g_tx_pcs_tx_control_out_krfec[2], w_hssi_10g_tx_pcs_tx_control_out_krfec[1], w_hssi_10g_tx_pcs_tx_control_out_krfec[0]}),
				.tx_data_in({w_hssi_10g_tx_pcs_tx_data_out_krfec[63], w_hssi_10g_tx_pcs_tx_data_out_krfec[62], w_hssi_10g_tx_pcs_tx_data_out_krfec[61], w_hssi_10g_tx_pcs_tx_data_out_krfec[60], w_hssi_10g_tx_pcs_tx_data_out_krfec[59], w_hssi_10g_tx_pcs_tx_data_out_krfec[58], w_hssi_10g_tx_pcs_tx_data_out_krfec[57], w_hssi_10g_tx_pcs_tx_data_out_krfec[56], w_hssi_10g_tx_pcs_tx_data_out_krfec[55], w_hssi_10g_tx_pcs_tx_data_out_krfec[54], w_hssi_10g_tx_pcs_tx_data_out_krfec[53], w_hssi_10g_tx_pcs_tx_data_out_krfec[52], w_hssi_10g_tx_pcs_tx_data_out_krfec[51], w_hssi_10g_tx_pcs_tx_data_out_krfec[50], w_hssi_10g_tx_pcs_tx_data_out_krfec[49], w_hssi_10g_tx_pcs_tx_data_out_krfec[48], w_hssi_10g_tx_pcs_tx_data_out_krfec[47], w_hssi_10g_tx_pcs_tx_data_out_krfec[46], w_hssi_10g_tx_pcs_tx_data_out_krfec[45], w_hssi_10g_tx_pcs_tx_data_out_krfec[44], w_hssi_10g_tx_pcs_tx_data_out_krfec[43], w_hssi_10g_tx_pcs_tx_data_out_krfec[42], w_hssi_10g_tx_pcs_tx_data_out_krfec[41], w_hssi_10g_tx_pcs_tx_data_out_krfec[40], w_hssi_10g_tx_pcs_tx_data_out_krfec[39], w_hssi_10g_tx_pcs_tx_data_out_krfec[38], w_hssi_10g_tx_pcs_tx_data_out_krfec[37], w_hssi_10g_tx_pcs_tx_data_out_krfec[36], w_hssi_10g_tx_pcs_tx_data_out_krfec[35], w_hssi_10g_tx_pcs_tx_data_out_krfec[34], w_hssi_10g_tx_pcs_tx_data_out_krfec[33], w_hssi_10g_tx_pcs_tx_data_out_krfec[32], w_hssi_10g_tx_pcs_tx_data_out_krfec[31], w_hssi_10g_tx_pcs_tx_data_out_krfec[30], w_hssi_10g_tx_pcs_tx_data_out_krfec[29], w_hssi_10g_tx_pcs_tx_data_out_krfec[28], w_hssi_10g_tx_pcs_tx_data_out_krfec[27], w_hssi_10g_tx_pcs_tx_data_out_krfec[26], w_hssi_10g_tx_pcs_tx_data_out_krfec[25], w_hssi_10g_tx_pcs_tx_data_out_krfec[24], w_hssi_10g_tx_pcs_tx_data_out_krfec[23], w_hssi_10g_tx_pcs_tx_data_out_krfec[22], w_hssi_10g_tx_pcs_tx_data_out_krfec[21], w_hssi_10g_tx_pcs_tx_data_out_krfec[20], w_hssi_10g_tx_pcs_tx_data_out_krfec[19], w_hssi_10g_tx_pcs_tx_data_out_krfec[18], w_hssi_10g_tx_pcs_tx_data_out_krfec[17], w_hssi_10g_tx_pcs_tx_data_out_krfec[16], w_hssi_10g_tx_pcs_tx_data_out_krfec[15], w_hssi_10g_tx_pcs_tx_data_out_krfec[14], w_hssi_10g_tx_pcs_tx_data_out_krfec[13], w_hssi_10g_tx_pcs_tx_data_out_krfec[12], w_hssi_10g_tx_pcs_tx_data_out_krfec[11], w_hssi_10g_tx_pcs_tx_data_out_krfec[10], w_hssi_10g_tx_pcs_tx_data_out_krfec[9], w_hssi_10g_tx_pcs_tx_data_out_krfec[8], w_hssi_10g_tx_pcs_tx_data_out_krfec[7], w_hssi_10g_tx_pcs_tx_data_out_krfec[6], w_hssi_10g_tx_pcs_tx_data_out_krfec[5], w_hssi_10g_tx_pcs_tx_data_out_krfec[4], w_hssi_10g_tx_pcs_tx_data_out_krfec[3], w_hssi_10g_tx_pcs_tx_data_out_krfec[2], w_hssi_10g_tx_pcs_tx_data_out_krfec[1], w_hssi_10g_tx_pcs_tx_data_out_krfec[0]}),
				.tx_data_valid_in(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_krfec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_krfec_reg(),
				.pld_krfec_tx_alignment_plddirect_reg(),
				.pld_krfec_tx_alignment_reg()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_tx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_alignment = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_test_data[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen1_2
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen1_2
			twentynm_hssi_pipe_gen1_2 #(
				.elec_idle_delay_val(hssi_pipe_gen1_2_elec_idle_delay_val),
				.error_replace_pad(hssi_pipe_gen1_2_error_replace_pad),
				.hip_mode(hssi_pipe_gen1_2_hip_mode),
				.ind_error_reporting(hssi_pipe_gen1_2_ind_error_reporting),
				.phystatus_delay_val(hssi_pipe_gen1_2_phystatus_delay_val),
				.phystatus_rst_toggle(hssi_pipe_gen1_2_phystatus_rst_toggle),
				.pipe_byte_de_serializer_en(hssi_pipe_gen1_2_pipe_byte_de_serializer_en),
				.prot_mode(hssi_pipe_gen1_2_prot_mode),
				.reconfig_settings(hssi_pipe_gen1_2_reconfig_settings),
				.rx_pipe_enable(hssi_pipe_gen1_2_rx_pipe_enable),
				.rxdetect_bypass(hssi_pipe_gen1_2_rxdetect_bypass),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen1_2_sup_mode),
				.tx_pipe_enable(hssi_pipe_gen1_2_tx_pipe_enable),
				.txswing(hssi_pipe_gen1_2_txswing)
			) inst_twentynm_hssi_pipe_gen1_2 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen1_2_avmmreaddata),
				.blockselect(w_hssi_pipe_gen1_2_blockselect),
				.current_coeff(w_hssi_pipe_gen1_2_current_coeff),
				.phystatus(w_hssi_pipe_gen1_2_phystatus),
				.polarity_inversion_rx(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rev_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.rxelectricalidle_out(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxstatus(w_hssi_pipe_gen1_2_rxstatus),
				.rxvalid(w_hssi_pipe_gen1_2_rxvalid),
				.tx_elec_idle_out(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pipe_rx_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.power_state_transition_done_ena(1'b0),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rev_loopbk_pcs_gen3(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.revloopback(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.rx_pipe_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rxd({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxelectricalidle(w_hssi_8g_rx_pcs_eidle_detected),
				.rxelectricalidle_pcs_gen3(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.rxpolarity_pcs_gen3(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.tx_elec_idle_comp(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.txd_ch({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswingport(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.pld_8g_rxpolarity_pipe3_reg(),
				.rxd_ch(),
				.txd()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen1_2_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen1_2_blockselect = 1'b0;
				assign w_hssi_pipe_gen1_2_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen1_2_phystatus = 1'b0;
				assign w_hssi_pipe_gen1_2_polarity_inversion_rx = 1'b0;
				assign w_hssi_pipe_gen1_2_rev_loopbk = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelectricalidle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen1_2_rxvalid = 1'b0;
				assign w_hssi_pipe_gen1_2_tx_elec_idle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_txdetectrx = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen3
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen3
			twentynm_hssi_pipe_gen3 #(
				.bypass_rx_detection_enable(hssi_pipe_gen3_bypass_rx_detection_enable),
				.bypass_rx_preset(hssi_pipe_gen3_bypass_rx_preset),
				.bypass_rx_preset_enable(hssi_pipe_gen3_bypass_rx_preset_enable),
				.bypass_tx_coefficent(hssi_pipe_gen3_bypass_tx_coefficent),
				.bypass_tx_coefficent_enable(hssi_pipe_gen3_bypass_tx_coefficent_enable),
				.elecidle_delay_g3(hssi_pipe_gen3_elecidle_delay_g3),
				.ind_error_reporting(hssi_pipe_gen3_ind_error_reporting),
				.mode(hssi_pipe_gen3_mode),
				.phy_status_delay_g12(hssi_pipe_gen3_phy_status_delay_g12),
				.phy_status_delay_g3(hssi_pipe_gen3_phy_status_delay_g3),
				.phystatus_rst_toggle_g12(hssi_pipe_gen3_phystatus_rst_toggle_g12),
				.phystatus_rst_toggle_g3(hssi_pipe_gen3_phystatus_rst_toggle_g3),
				.rate_match_pad_insertion(hssi_pipe_gen3_rate_match_pad_insertion),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen3_sup_mode),
				.test_out_sel(hssi_pipe_gen3_test_out_sel)
			) inst_twentynm_hssi_pipe_gen3 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen3_avmmreaddata),
				.blockselect(w_hssi_pipe_gen3_blockselect),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.phystatus(w_hssi_pipe_gen3_phystatus),
				.pma_current_coeff(w_hssi_pipe_gen3_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_pipe_gen3_pma_current_rxpreset),
				.pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.rev_lpbk_8gpcs_out(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.rev_lpbk_int(w_hssi_pipe_gen3_rev_lpbk_int),
				.rx_blk_start(w_hssi_pipe_gen3_rx_blk_start),
				.rx_sync_hdr(w_hssi_pipe_gen3_rx_sync_hdr),
				.rxd_8gpcs_out(w_hssi_pipe_gen3_rxd_8gpcs_out),
				.rxdataskip(w_hssi_pipe_gen3_rxdataskip),
				.rxelecidle(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity_8gpcs_out(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.rxpolarity_int(w_hssi_pipe_gen3_rxpolarity_int),
				.rxstatus(w_hssi_pipe_gen3_rxstatus),
				.rxvalid(w_hssi_pipe_gen3_rxvalid),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.test_out(w_hssi_pipe_gen3_test_out),
				.tx_blk_start_int(w_hssi_pipe_gen3_tx_blk_start_int),
				.tx_sync_hdr_int(w_hssi_pipe_gen3_tx_sync_hdr_int),
				.txdata_int(w_hssi_pipe_gen3_txdata_int),
				.txdatak_int(w_hssi_pipe_gen3_txdatak_int),
				.txdataskip_int(w_hssi_pipe_gen3_txdataskip_int),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.current_coeff({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0]}),
				.current_rxpreset({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0]}),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.pcs_asn_bundling_in({w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0]}),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pipe_tx_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_blk_start_int(w_hssi_gen3_rx_pcs_blk_start),
				.rx_sync_hdr_int({w_hssi_gen3_rx_pcs_sync_hdr[1], w_hssi_gen3_rx_pcs_sync_hdr[0]}),
				.rx_test_out({w_hssi_gen3_rx_pcs_rx_test_out[19], w_hssi_gen3_rx_pcs_rx_test_out[18], w_hssi_gen3_rx_pcs_rx_test_out[17], w_hssi_gen3_rx_pcs_rx_test_out[16], w_hssi_gen3_rx_pcs_rx_test_out[15], w_hssi_gen3_rx_pcs_rx_test_out[14], w_hssi_gen3_rx_pcs_rx_test_out[13], w_hssi_gen3_rx_pcs_rx_test_out[12], w_hssi_gen3_rx_pcs_rx_test_out[11], w_hssi_gen3_rx_pcs_rx_test_out[10], w_hssi_gen3_rx_pcs_rx_test_out[9], w_hssi_gen3_rx_pcs_rx_test_out[8], w_hssi_gen3_rx_pcs_rx_test_out[7], w_hssi_gen3_rx_pcs_rx_test_out[6], w_hssi_gen3_rx_pcs_rx_test_out[5], w_hssi_gen3_rx_pcs_rx_test_out[4], w_hssi_gen3_rx_pcs_rx_test_out[3], w_hssi_gen3_rx_pcs_rx_test_out[2], w_hssi_gen3_rx_pcs_rx_test_out[1], w_hssi_gen3_rx_pcs_rx_test_out[0]}),
				.rxd_8gpcs_in({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxdata_int({w_hssi_gen3_rx_pcs_data_out[31], w_hssi_gen3_rx_pcs_data_out[30], w_hssi_gen3_rx_pcs_data_out[29], w_hssi_gen3_rx_pcs_data_out[28], w_hssi_gen3_rx_pcs_data_out[27], w_hssi_gen3_rx_pcs_data_out[26], w_hssi_gen3_rx_pcs_data_out[25], w_hssi_gen3_rx_pcs_data_out[24], w_hssi_gen3_rx_pcs_data_out[23], w_hssi_gen3_rx_pcs_data_out[22], w_hssi_gen3_rx_pcs_data_out[21], w_hssi_gen3_rx_pcs_data_out[20], w_hssi_gen3_rx_pcs_data_out[19], w_hssi_gen3_rx_pcs_data_out[18], w_hssi_gen3_rx_pcs_data_out[17], w_hssi_gen3_rx_pcs_data_out[16], w_hssi_gen3_rx_pcs_data_out[15], w_hssi_gen3_rx_pcs_data_out[14], w_hssi_gen3_rx_pcs_data_out[13], w_hssi_gen3_rx_pcs_data_out[12], w_hssi_gen3_rx_pcs_data_out[11], w_hssi_gen3_rx_pcs_data_out[10], w_hssi_gen3_rx_pcs_data_out[9], w_hssi_gen3_rx_pcs_data_out[8], w_hssi_gen3_rx_pcs_data_out[7], w_hssi_gen3_rx_pcs_data_out[6], w_hssi_gen3_rx_pcs_data_out[5], w_hssi_gen3_rx_pcs_data_out[4], w_hssi_gen3_rx_pcs_data_out[3], w_hssi_gen3_rx_pcs_data_out[2], w_hssi_gen3_rx_pcs_data_out[1], w_hssi_gen3_rx_pcs_data_out[0]}),
				.rxdatak_int({1'b0, 1'b0, 1'b0, 1'b0}),
				.rxdataskip_int(w_hssi_gen3_rx_pcs_data_valid),
				.rxelecidle_8gpcs_in(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.tx_blk_start(w_hssi_8g_tx_pcs_tx_blk_start_out[0]),
				.tx_sync_hdr({w_hssi_8g_tx_pcs_tx_sync_hdr_out[1], w_hssi_8g_tx_pcs_tx_sync_hdr_out[0]}),
				.tx_test_out({w_hssi_gen3_tx_pcs_tx_test_out[19], w_hssi_gen3_tx_pcs_tx_test_out[18], w_hssi_gen3_tx_pcs_tx_test_out[17], w_hssi_gen3_tx_pcs_tx_test_out[16], w_hssi_gen3_tx_pcs_tx_test_out[15], w_hssi_gen3_tx_pcs_tx_test_out[14], w_hssi_gen3_tx_pcs_tx_test_out[13], w_hssi_gen3_tx_pcs_tx_test_out[12], w_hssi_gen3_tx_pcs_tx_test_out[11], w_hssi_gen3_tx_pcs_tx_test_out[10], w_hssi_gen3_tx_pcs_tx_test_out[9], w_hssi_gen3_tx_pcs_tx_test_out[8], w_hssi_gen3_tx_pcs_tx_test_out[7], w_hssi_gen3_tx_pcs_tx_test_out[6], w_hssi_gen3_tx_pcs_tx_test_out[5], w_hssi_gen3_tx_pcs_tx_test_out[4], w_hssi_gen3_tx_pcs_tx_test_out[3], w_hssi_gen3_tx_pcs_tx_test_out[2], w_hssi_gen3_tx_pcs_tx_test_out[1], w_hssi_gen3_tx_pcs_tx_test_out[0]}),
				.txcompliance(w_hssi_8g_tx_pcs_txcompliance_out),
				.txdata({w_hssi_8g_tx_pcs_tx_data_out[31], w_hssi_8g_tx_pcs_tx_data_out[30], w_hssi_8g_tx_pcs_tx_data_out[29], w_hssi_8g_tx_pcs_tx_data_out[28], w_hssi_8g_tx_pcs_tx_data_out[27], w_hssi_8g_tx_pcs_tx_data_out[26], w_hssi_8g_tx_pcs_tx_data_out[25], w_hssi_8g_tx_pcs_tx_data_out[24], w_hssi_8g_tx_pcs_tx_data_out[23], w_hssi_8g_tx_pcs_tx_data_out[22], w_hssi_8g_tx_pcs_tx_data_out[21], w_hssi_8g_tx_pcs_tx_data_out[20], w_hssi_8g_tx_pcs_tx_data_out[19], w_hssi_8g_tx_pcs_tx_data_out[18], w_hssi_8g_tx_pcs_tx_data_out[17], w_hssi_8g_tx_pcs_tx_data_out[16], w_hssi_8g_tx_pcs_tx_data_out[15], w_hssi_8g_tx_pcs_tx_data_out[14], w_hssi_8g_tx_pcs_tx_data_out[13], w_hssi_8g_tx_pcs_tx_data_out[12], w_hssi_8g_tx_pcs_tx_data_out[11], w_hssi_8g_tx_pcs_tx_data_out[10], w_hssi_8g_tx_pcs_tx_data_out[9], w_hssi_8g_tx_pcs_tx_data_out[8], w_hssi_8g_tx_pcs_tx_data_out[7], w_hssi_8g_tx_pcs_tx_data_out[6], w_hssi_8g_tx_pcs_tx_data_out[5], w_hssi_8g_tx_pcs_tx_data_out[4], w_hssi_8g_tx_pcs_tx_data_out[3], w_hssi_8g_tx_pcs_tx_data_out[2], w_hssi_8g_tx_pcs_tx_data_out[1], w_hssi_8g_tx_pcs_tx_data_out[0]}),
				.txdatak({w_hssi_8g_tx_pcs_tx_datak_out[3], w_hssi_8g_tx_pcs_tx_datak_out[2], w_hssi_8g_tx_pcs_tx_datak_out[1], w_hssi_8g_tx_pcs_tx_datak_out[0]}),
				.txdataskip(w_hssi_8g_tx_pcs_tx_data_valid_out[0]),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_8g_tx_pcs_txelecidle_out),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.dis_pc_byte(),
				.pma_rx_det_pd(),
				.pma_txdeemph(),
				.pma_txmargin(),
				.pma_txswing(),
				.reset_pc_prts()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen3_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen3_blockselect = 1'b0;
				assign w_hssi_pipe_gen3_gen3_clk_sel = 1'b0;
				assign w_hssi_pipe_gen3_pcs_rst = 1'b0;
				assign w_hssi_pipe_gen3_phystatus = 1'b0;
				assign w_hssi_pipe_gen3_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen3_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_pma_tx_elec_idle = 1'b0;
				assign w_hssi_pipe_gen3_pma_txdetectrx = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_int = 1'b0;
				assign w_hssi_pipe_gen3_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_rxd_8gpcs_out[63:0] = 64'b0;
				assign w_hssi_pipe_gen3_rxdataskip[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_int = 1'b0;
				assign w_hssi_pipe_gen3_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_rxvalid = 1'b0;
				assign w_hssi_pipe_gen3_shutdown_clk = 1'b0;
				assign w_hssi_pipe_gen3_test_out[19:0] = 20'b0;
				assign w_hssi_pipe_gen3_tx_blk_start_int = 1'b0;
				assign w_hssi_pipe_gen3_tx_sync_hdr_int[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_txdata_int[31:0] = 32'b0;
				assign w_hssi_pipe_gen3_txdatak_int[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_txdataskip_int = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pcs_pma_interface
			twentynm_hssi_rx_pcs_pma_interface #(
				.block_sel(hssi_rx_pcs_pma_interface_block_sel),
				.channel_operation_mode(hssi_rx_pcs_pma_interface_channel_operation_mode),
				.clkslip_sel(hssi_rx_pcs_pma_interface_clkslip_sel),
				.lpbk_en(hssi_rx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_rx_pcs_pma_interface_master_clk_sel),
				.pldif_datawidth_mode(hssi_rx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_rx(hssi_rx_pcs_pma_interface_pma_dw_rx),
				.pma_if_dft_en(hssi_rx_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_rx_pcs_pma_interface_pma_if_dft_val),
				.prbs9_dwidth(hssi_rx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_rx_pcs_pma_interface_prbs_clken),
				.prbs_ver(hssi_rx_pcs_pma_interface_prbs_ver),
				.prot_mode_rx(hssi_rx_pcs_pma_interface_prot_mode_rx),
				.reconfig_settings(hssi_rx_pcs_pma_interface_reconfig_settings),
				.rx_dyn_polarity_inversion(hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion),
				.rx_lpbk_en(hssi_rx_pcs_pma_interface_rx_lpbk_en),
				.rx_prbs_force_signal_ok(hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok),
				.rx_prbs_mask(hssi_rx_pcs_pma_interface_rx_prbs_mask),
				.rx_prbs_mode(hssi_rx_pcs_pma_interface_rx_prbs_mode),
				.rx_signalok_signaldet_sel(hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel),
				.rx_static_polarity_inversion(hssi_rx_pcs_pma_interface_rx_static_polarity_inversion),
				.rx_uhsif_lpbk_en(hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sup_mode(hssi_rx_pcs_pma_interface_sup_mode)
			) inst_twentynm_hssi_rx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.int_pmaif_10g_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data),
				.int_pmaif_10g_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.int_pmaif_8g_pudi(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi),
				.int_pmaif_8g_rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.int_pmaif_8g_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.int_pmaif_8g_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.int_pmaif_8g_sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.int_pmaif_g3_pma_data_in(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in),
				.int_pmaif_g3_pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.int_pmaif_g3_pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.int_pmaif_g3_pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.int_pmaif_krfec_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data),
				.int_pmaif_krfec_rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.int_pmaif_pldif_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pmaif_pldif_prbs_err_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pmaif_pldif_rx_clkdiv(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pmaif_pldif_rx_clkdiv_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pmaif_pldif_rx_data(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data),
				.int_pmaif_pldif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pmaif_pldif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pmaif_pldif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pmaif_pldif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.pma_eye_monitor(w_hssi_rx_pcs_pma_interface_pma_eye_monitor),
				.pma_rx_clkslip(w_hssi_rx_pcs_pma_interface_pma_rx_clkslip),
				.pma_rxpma_rstb(w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb),
				.rx_pmaif_test_out(w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out),
				.rx_prbs_ver_test(w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.int_pmaif_8g_rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.int_pmaif_pldif_eye_monitor({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0]}),
				.int_pmaif_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pmaif_pldif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pmaif_pldif_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pmaif_pldif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pma_rx_clkdiv_user(in_pma_rx_clkdiv_user),
				.pma_rx_detect_valid(in_pma_rx_detect_valid),
				.pma_rx_found(in_pma_rx_found),
				.pma_rx_pma_clk(in_pma_rx_pma_clk),
				.pma_rx_pma_data({in_pma_rx_pma_data[63], in_pma_rx_pma_data[62], in_pma_rx_pma_data[61], in_pma_rx_pma_data[60], in_pma_rx_pma_data[59], in_pma_rx_pma_data[58], in_pma_rx_pma_data[57], in_pma_rx_pma_data[56], in_pma_rx_pma_data[55], in_pma_rx_pma_data[54], in_pma_rx_pma_data[53], in_pma_rx_pma_data[52], in_pma_rx_pma_data[51], in_pma_rx_pma_data[50], in_pma_rx_pma_data[49], in_pma_rx_pma_data[48], in_pma_rx_pma_data[47], in_pma_rx_pma_data[46], in_pma_rx_pma_data[45], in_pma_rx_pma_data[44], in_pma_rx_pma_data[43], in_pma_rx_pma_data[42], in_pma_rx_pma_data[41], in_pma_rx_pma_data[40], in_pma_rx_pma_data[39], in_pma_rx_pma_data[38], in_pma_rx_pma_data[37], in_pma_rx_pma_data[36], in_pma_rx_pma_data[35], in_pma_rx_pma_data[34], in_pma_rx_pma_data[33], in_pma_rx_pma_data[32], in_pma_rx_pma_data[31], in_pma_rx_pma_data[30], in_pma_rx_pma_data[29], in_pma_rx_pma_data[28], in_pma_rx_pma_data[27], in_pma_rx_pma_data[26], in_pma_rx_pma_data[25], in_pma_rx_pma_data[24], in_pma_rx_pma_data[23], in_pma_rx_pma_data[22], in_pma_rx_pma_data[21], in_pma_rx_pma_data[20], in_pma_rx_pma_data[19], in_pma_rx_pma_data[18], in_pma_rx_pma_data[17], in_pma_rx_pma_data[16], in_pma_rx_pma_data[15], in_pma_rx_pma_data[14], in_pma_rx_pma_data[13], in_pma_rx_pma_data[12], in_pma_rx_pma_data[11], in_pma_rx_pma_data[10], in_pma_rx_pma_data[9], in_pma_rx_pma_data[8], in_pma_rx_pma_data[7], in_pma_rx_pma_data[6], in_pma_rx_pma_data[5], in_pma_rx_pma_data[4], in_pma_rx_pma_data[3], in_pma_rx_pma_data[2], in_pma_rx_pma_data[1], in_pma_rx_pma_data[0]}),
				.pma_rx_signal_ok(in_pma_rx_signal_ok),
				.pma_rxpll_lock(in_pma_rxpll_lock),
				.pma_signal_det(in_pma_signal_det),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.tx_pma_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0]}),
				.tx_pma_uhsif_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0]}),
				
				// UNUSED
				.int_pmaif_g3_rcvd_clk(),
				.prbs_err_lt()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31:0] = 32'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5:0] = 6'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rx_clkslip = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pld_pcs_interface
			twentynm_hssi_rx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx),
				.hd_10g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx),
				.hd_10g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx),
				.hd_10g_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx),
				.hd_10g_lpbk_en(hssi_rx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx),
				.hd_10g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx),
				.hd_10g_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx),
				.hd_10g_test_bus_mode(hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode),
				.hd_8g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx),
				.hd_8g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx),
				.hd_8g_hip_mode(hssi_rx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_rx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx),
				.hd_8g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx),
				.hd_chnl_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_clklow_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz),
				.hd_chnl_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx),
				.hd_chnl_fref_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz),
				.hd_chnl_frequency_rules_en(hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_rx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_rx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx),
				.hd_chnl_lpbk_en(hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx),
				.hd_chnl_pld_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz),
				.hd_chnl_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx),
				.hd_chnl_pma_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz),
				.hd_chnl_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx),
				.hd_chnl_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx),
				.hd_chnl_transparent_pcs_rx(hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx),
				.hd_fifo_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx),
				.hd_fifo_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx),
				.hd_g3_prot_mode(hssi_rx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx),
				.hd_krfec_lpbk_en(hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx),
				.hd_krfec_test_bus_mode(hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode),
				.hd_pldif_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx),
				.hd_pmaif_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_lpbk_en(hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx),
				.hd_pmaif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx),
				.hd_pmaif_sim_mode(hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_rx_block_sel(hssi_rx_pld_pcs_interface_pcs_rx_block_sel),
				.pcs_rx_clk_out_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel),
				.pcs_rx_clk_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_sel),
				.pcs_rx_hip_clk_en(hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en),
				.pcs_rx_output_sel(hssi_rx_pld_pcs_interface_pcs_rx_output_sel),
				.reconfig_settings(hssi_rx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm4" )       //PARAM_HIDE
			) inst_twentynm_hssi_rx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pld_pcs_interface_blockselect),
				.hip_rx_ctrl(w_hssi_rx_pld_pcs_interface_hip_rx_ctrl),
				.hip_rx_data(w_hssi_rx_pld_pcs_interface_hip_rx_data),
				.int_pldif_10g_rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.int_pldif_10g_rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.int_pldif_10g_rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.int_pldif_10g_rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.int_pldif_10g_rx_control_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb),
				.int_pldif_10g_rx_data_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb),
				.int_pldif_10g_rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.int_pldif_10g_rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.int_pldif_10g_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.int_pldif_10g_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.int_pldif_10g_rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.int_pldif_8g_a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.int_pldif_8g_bitloc_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.int_pldif_8g_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.int_pldif_8g_byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.int_pldif_8g_encdt(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.int_pldif_8g_pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.int_pldif_8g_rdenable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.int_pldif_8g_rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.int_pldif_8g_rxurstpcs_n(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.int_pldif_8g_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.int_pldif_8g_wrdisable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.int_pldif_g3_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.int_pldif_krfec_rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.int_pldif_pmaif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pldif_pmaif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pldif_pmaif_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pldif_pmaif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pld_10g_krfec_rx_blk_lock(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock),
				.pld_10g_krfec_rx_diag_data_status(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status),
				.pld_10g_krfec_rx_frame(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame),
				.pld_10g_rx_align_val(w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val),
				.pld_10g_rx_crc32_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err),
				.pld_10g_rx_data_valid(w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid),
				.pld_10g_rx_empty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty),
				.pld_10g_rx_fifo_del(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del),
				.pld_10g_rx_fifo_insert(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert),
				.pld_10g_rx_fifo_num(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num),
				.pld_10g_rx_frame_lock(w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock),
				.pld_10g_rx_hi_ber(w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber),
				.pld_10g_rx_oflw_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err),
				.pld_10g_rx_pempty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty),
				.pld_10g_rx_pfull(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull),
				.pld_8g_a1a2_k1k2_flag(w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag),
				.pld_8g_empty_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf),
				.pld_8g_empty_rx(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx),
				.pld_8g_full_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf),
				.pld_8g_full_rx(w_hssi_rx_pld_pcs_interface_pld_8g_full_rx),
				.pld_8g_rxelecidle(w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle),
				.pld_8g_signal_detect_out(w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out),
				.pld_8g_wa_boundary(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary),
				.pld_pcs_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out),
				.pld_pma_clkdiv_rx_user(w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user),
				.pld_pma_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out),
				.pld_pma_signal_ok(w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok),
				.pld_rx_control(w_hssi_rx_pld_pcs_interface_pld_rx_control),
				.pld_rx_data(w_hssi_rx_pld_pcs_interface_pld_rx_data),
				.pld_rx_prbs_done(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done),
				.pld_rx_prbs_err(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.int_pldif_10g_rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.int_pldif_10g_rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.int_pldif_10g_rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_10g_rx_control({w_hssi_10g_rx_pcs_rx_control[19], w_hssi_10g_rx_pcs_rx_control[18], w_hssi_10g_rx_pcs_rx_control[17], w_hssi_10g_rx_pcs_rx_control[16], w_hssi_10g_rx_pcs_rx_control[15], w_hssi_10g_rx_pcs_rx_control[14], w_hssi_10g_rx_pcs_rx_control[13], w_hssi_10g_rx_pcs_rx_control[12], w_hssi_10g_rx_pcs_rx_control[11], w_hssi_10g_rx_pcs_rx_control[10], w_hssi_10g_rx_pcs_rx_control[9], w_hssi_10g_rx_pcs_rx_control[8], w_hssi_10g_rx_pcs_rx_control[7], w_hssi_10g_rx_pcs_rx_control[6], w_hssi_10g_rx_pcs_rx_control[5], w_hssi_10g_rx_pcs_rx_control[4], w_hssi_10g_rx_pcs_rx_control[3], w_hssi_10g_rx_pcs_rx_control[2], w_hssi_10g_rx_pcs_rx_control[1], w_hssi_10g_rx_pcs_rx_control[0]}),
				.int_pldif_10g_rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.int_pldif_10g_rx_data({w_hssi_10g_rx_pcs_rx_data[127], w_hssi_10g_rx_pcs_rx_data[126], w_hssi_10g_rx_pcs_rx_data[125], w_hssi_10g_rx_pcs_rx_data[124], w_hssi_10g_rx_pcs_rx_data[123], w_hssi_10g_rx_pcs_rx_data[122], w_hssi_10g_rx_pcs_rx_data[121], w_hssi_10g_rx_pcs_rx_data[120], w_hssi_10g_rx_pcs_rx_data[119], w_hssi_10g_rx_pcs_rx_data[118], w_hssi_10g_rx_pcs_rx_data[117], w_hssi_10g_rx_pcs_rx_data[116], w_hssi_10g_rx_pcs_rx_data[115], w_hssi_10g_rx_pcs_rx_data[114], w_hssi_10g_rx_pcs_rx_data[113], w_hssi_10g_rx_pcs_rx_data[112], w_hssi_10g_rx_pcs_rx_data[111], w_hssi_10g_rx_pcs_rx_data[110], w_hssi_10g_rx_pcs_rx_data[109], w_hssi_10g_rx_pcs_rx_data[108], w_hssi_10g_rx_pcs_rx_data[107], w_hssi_10g_rx_pcs_rx_data[106], w_hssi_10g_rx_pcs_rx_data[105], w_hssi_10g_rx_pcs_rx_data[104], w_hssi_10g_rx_pcs_rx_data[103], w_hssi_10g_rx_pcs_rx_data[102], w_hssi_10g_rx_pcs_rx_data[101], w_hssi_10g_rx_pcs_rx_data[100], w_hssi_10g_rx_pcs_rx_data[99], w_hssi_10g_rx_pcs_rx_data[98], w_hssi_10g_rx_pcs_rx_data[97], w_hssi_10g_rx_pcs_rx_data[96], w_hssi_10g_rx_pcs_rx_data[95], w_hssi_10g_rx_pcs_rx_data[94], w_hssi_10g_rx_pcs_rx_data[93], w_hssi_10g_rx_pcs_rx_data[92], w_hssi_10g_rx_pcs_rx_data[91], w_hssi_10g_rx_pcs_rx_data[90], w_hssi_10g_rx_pcs_rx_data[89], w_hssi_10g_rx_pcs_rx_data[88], w_hssi_10g_rx_pcs_rx_data[87], w_hssi_10g_rx_pcs_rx_data[86], w_hssi_10g_rx_pcs_rx_data[85], w_hssi_10g_rx_pcs_rx_data[84], w_hssi_10g_rx_pcs_rx_data[83], w_hssi_10g_rx_pcs_rx_data[82], w_hssi_10g_rx_pcs_rx_data[81], w_hssi_10g_rx_pcs_rx_data[80], w_hssi_10g_rx_pcs_rx_data[79], w_hssi_10g_rx_pcs_rx_data[78], w_hssi_10g_rx_pcs_rx_data[77], w_hssi_10g_rx_pcs_rx_data[76], w_hssi_10g_rx_pcs_rx_data[75], w_hssi_10g_rx_pcs_rx_data[74], w_hssi_10g_rx_pcs_rx_data[73], w_hssi_10g_rx_pcs_rx_data[72], w_hssi_10g_rx_pcs_rx_data[71], w_hssi_10g_rx_pcs_rx_data[70], w_hssi_10g_rx_pcs_rx_data[69], w_hssi_10g_rx_pcs_rx_data[68], w_hssi_10g_rx_pcs_rx_data[67], w_hssi_10g_rx_pcs_rx_data[66], w_hssi_10g_rx_pcs_rx_data[65], w_hssi_10g_rx_pcs_rx_data[64], w_hssi_10g_rx_pcs_rx_data[63], w_hssi_10g_rx_pcs_rx_data[62], w_hssi_10g_rx_pcs_rx_data[61], w_hssi_10g_rx_pcs_rx_data[60], w_hssi_10g_rx_pcs_rx_data[59], w_hssi_10g_rx_pcs_rx_data[58], w_hssi_10g_rx_pcs_rx_data[57], w_hssi_10g_rx_pcs_rx_data[56], w_hssi_10g_rx_pcs_rx_data[55], w_hssi_10g_rx_pcs_rx_data[54], w_hssi_10g_rx_pcs_rx_data[53], w_hssi_10g_rx_pcs_rx_data[52], w_hssi_10g_rx_pcs_rx_data[51], w_hssi_10g_rx_pcs_rx_data[50], w_hssi_10g_rx_pcs_rx_data[49], w_hssi_10g_rx_pcs_rx_data[48], w_hssi_10g_rx_pcs_rx_data[47], w_hssi_10g_rx_pcs_rx_data[46], w_hssi_10g_rx_pcs_rx_data[45], w_hssi_10g_rx_pcs_rx_data[44], w_hssi_10g_rx_pcs_rx_data[43], w_hssi_10g_rx_pcs_rx_data[42], w_hssi_10g_rx_pcs_rx_data[41], w_hssi_10g_rx_pcs_rx_data[40], w_hssi_10g_rx_pcs_rx_data[39], w_hssi_10g_rx_pcs_rx_data[38], w_hssi_10g_rx_pcs_rx_data[37], w_hssi_10g_rx_pcs_rx_data[36], w_hssi_10g_rx_pcs_rx_data[35], w_hssi_10g_rx_pcs_rx_data[34], w_hssi_10g_rx_pcs_rx_data[33], w_hssi_10g_rx_pcs_rx_data[32], w_hssi_10g_rx_pcs_rx_data[31], w_hssi_10g_rx_pcs_rx_data[30], w_hssi_10g_rx_pcs_rx_data[29], w_hssi_10g_rx_pcs_rx_data[28], w_hssi_10g_rx_pcs_rx_data[27], w_hssi_10g_rx_pcs_rx_data[26], w_hssi_10g_rx_pcs_rx_data[25], w_hssi_10g_rx_pcs_rx_data[24], w_hssi_10g_rx_pcs_rx_data[23], w_hssi_10g_rx_pcs_rx_data[22], w_hssi_10g_rx_pcs_rx_data[21], w_hssi_10g_rx_pcs_rx_data[20], w_hssi_10g_rx_pcs_rx_data[19], w_hssi_10g_rx_pcs_rx_data[18], w_hssi_10g_rx_pcs_rx_data[17], w_hssi_10g_rx_pcs_rx_data[16], w_hssi_10g_rx_pcs_rx_data[15], w_hssi_10g_rx_pcs_rx_data[14], w_hssi_10g_rx_pcs_rx_data[13], w_hssi_10g_rx_pcs_rx_data[12], w_hssi_10g_rx_pcs_rx_data[11], w_hssi_10g_rx_pcs_rx_data[10], w_hssi_10g_rx_pcs_rx_data[9], w_hssi_10g_rx_pcs_rx_data[8], w_hssi_10g_rx_pcs_rx_data[7], w_hssi_10g_rx_pcs_rx_data[6], w_hssi_10g_rx_pcs_rx_data[5], w_hssi_10g_rx_pcs_rx_data[4], w_hssi_10g_rx_pcs_rx_data[3], w_hssi_10g_rx_pcs_rx_data[2], w_hssi_10g_rx_pcs_rx_data[1], w_hssi_10g_rx_pcs_rx_data[0]}),
				.int_pldif_10g_rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.int_pldif_10g_rx_diag_status({w_hssi_10g_rx_pcs_rx_diag_status[1], w_hssi_10g_rx_pcs_rx_diag_status[0]}),
				.int_pldif_10g_rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.int_pldif_10g_rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.int_pldif_10g_rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.int_pldif_10g_rx_fifo_num({w_hssi_10g_rx_pcs_rx_fifo_num[4], w_hssi_10g_rx_pcs_rx_fifo_num[3], w_hssi_10g_rx_pcs_rx_fifo_num[2], w_hssi_10g_rx_pcs_rx_fifo_num[1], w_hssi_10g_rx_pcs_rx_fifo_num[0]}),
				.int_pldif_10g_rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.int_pldif_10g_rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.int_pldif_10g_rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.int_pldif_10g_rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.int_pldif_10g_rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.int_pldif_10g_rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				.int_pldif_8g_a1a2_k1k2_flag({w_hssi_8g_rx_pcs_a1a2k1k2flag[3], w_hssi_8g_rx_pcs_a1a2k1k2flag[2], w_hssi_8g_rx_pcs_a1a2k1k2flag[1], w_hssi_8g_rx_pcs_a1a2k1k2flag[0]}),
				.int_pldif_8g_empty_rmf(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.int_pldif_8g_empty_rx(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.int_pldif_8g_full_rmf(w_hssi_8g_rx_pcs_rm_fifo_full),
				.int_pldif_8g_full_rx(w_hssi_8g_rx_pcs_pcfifofull),
				.int_pldif_8g_phystatus(w_hssi_8g_rx_pcs_phystatus),
				.int_pldif_8g_rx_blk_start({w_hssi_8g_rx_pcs_rx_blk_start[3], w_hssi_8g_rx_pcs_rx_blk_start[2], w_hssi_8g_rx_pcs_rx_blk_start[1], w_hssi_8g_rx_pcs_rx_blk_start[0]}),
				.int_pldif_8g_rx_clk(w_hssi_8g_rx_pcs_clock_to_pld),
				.int_pldif_8g_rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_8g_rx_data_valid({w_hssi_8g_rx_pcs_rx_data_valid[3], w_hssi_8g_rx_pcs_rx_data_valid[2], w_hssi_8g_rx_pcs_rx_data_valid[1], w_hssi_8g_rx_pcs_rx_data_valid[0]}),
				.int_pldif_8g_rx_rstn_sync2wrfifo(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.int_pldif_8g_rx_sync_hdr({w_hssi_8g_rx_pcs_rx_sync_hdr[1], w_hssi_8g_rx_pcs_rx_sync_hdr[0]}),
				.int_pldif_8g_rxd({w_hssi_8g_rx_pcs_dataout[63], w_hssi_8g_rx_pcs_dataout[62], w_hssi_8g_rx_pcs_dataout[61], w_hssi_8g_rx_pcs_dataout[60], w_hssi_8g_rx_pcs_dataout[59], w_hssi_8g_rx_pcs_dataout[58], w_hssi_8g_rx_pcs_dataout[57], w_hssi_8g_rx_pcs_dataout[56], w_hssi_8g_rx_pcs_dataout[55], w_hssi_8g_rx_pcs_dataout[54], w_hssi_8g_rx_pcs_dataout[53], w_hssi_8g_rx_pcs_dataout[52], w_hssi_8g_rx_pcs_dataout[51], w_hssi_8g_rx_pcs_dataout[50], w_hssi_8g_rx_pcs_dataout[49], w_hssi_8g_rx_pcs_dataout[48], w_hssi_8g_rx_pcs_dataout[47], w_hssi_8g_rx_pcs_dataout[46], w_hssi_8g_rx_pcs_dataout[45], w_hssi_8g_rx_pcs_dataout[44], w_hssi_8g_rx_pcs_dataout[43], w_hssi_8g_rx_pcs_dataout[42], w_hssi_8g_rx_pcs_dataout[41], w_hssi_8g_rx_pcs_dataout[40], w_hssi_8g_rx_pcs_dataout[39], w_hssi_8g_rx_pcs_dataout[38], w_hssi_8g_rx_pcs_dataout[37], w_hssi_8g_rx_pcs_dataout[36], w_hssi_8g_rx_pcs_dataout[35], w_hssi_8g_rx_pcs_dataout[34], w_hssi_8g_rx_pcs_dataout[33], w_hssi_8g_rx_pcs_dataout[32], w_hssi_8g_rx_pcs_dataout[31], w_hssi_8g_rx_pcs_dataout[30], w_hssi_8g_rx_pcs_dataout[29], w_hssi_8g_rx_pcs_dataout[28], w_hssi_8g_rx_pcs_dataout[27], w_hssi_8g_rx_pcs_dataout[26], w_hssi_8g_rx_pcs_dataout[25], w_hssi_8g_rx_pcs_dataout[24], w_hssi_8g_rx_pcs_dataout[23], w_hssi_8g_rx_pcs_dataout[22], w_hssi_8g_rx_pcs_dataout[21], w_hssi_8g_rx_pcs_dataout[20], w_hssi_8g_rx_pcs_dataout[19], w_hssi_8g_rx_pcs_dataout[18], w_hssi_8g_rx_pcs_dataout[17], w_hssi_8g_rx_pcs_dataout[16], w_hssi_8g_rx_pcs_dataout[15], w_hssi_8g_rx_pcs_dataout[14], w_hssi_8g_rx_pcs_dataout[13], w_hssi_8g_rx_pcs_dataout[12], w_hssi_8g_rx_pcs_dataout[11], w_hssi_8g_rx_pcs_dataout[10], w_hssi_8g_rx_pcs_dataout[9], w_hssi_8g_rx_pcs_dataout[8], w_hssi_8g_rx_pcs_dataout[7], w_hssi_8g_rx_pcs_dataout[6], w_hssi_8g_rx_pcs_dataout[5], w_hssi_8g_rx_pcs_dataout[4], w_hssi_8g_rx_pcs_dataout[3], w_hssi_8g_rx_pcs_dataout[2], w_hssi_8g_rx_pcs_dataout[1], w_hssi_8g_rx_pcs_dataout[0]}),
				.int_pldif_8g_rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.int_pldif_8g_rxstatus({w_hssi_8g_rx_pcs_rxstatus[2], w_hssi_8g_rx_pcs_rxstatus[1], w_hssi_8g_rx_pcs_rxstatus[0]}),
				.int_pldif_8g_rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.int_pldif_8g_signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.int_pldif_8g_wa_boundary({w_hssi_8g_rx_pcs_word_align_boundary[4], w_hssi_8g_rx_pcs_word_align_boundary[3], w_hssi_8g_rx_pcs_word_align_boundary[2], w_hssi_8g_rx_pcs_word_align_boundary[1], w_hssi_8g_rx_pcs_word_align_boundary[0]}),
				.int_pldif_krfec_rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.int_pldif_krfec_rx_data_status({w_hssi_krfec_rx_pcs_rx_data_status[1], w_hssi_krfec_rx_pcs_rx_data_status[0]}),
				.int_pldif_krfec_rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.int_pldif_pmaif_clkdiv_rx(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pldif_pmaif_clkdiv_rx_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pldif_pmaif_rx_data({w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0]}),
				.int_pldif_pmaif_rx_prbs_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pldif_pmaif_rx_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.pld_10g_krfec_rx_clr_errblk_cnt(in_pld_10g_krfec_rx_clr_errblk_cnt),
				.pld_10g_krfec_rx_pld_rst_n(in_pld_10g_krfec_rx_pld_rst_n),
				.pld_10g_rx_align_clr(in_pld_10g_rx_align_clr),
				.pld_10g_rx_clr_ber_count(in_pld_10g_rx_clr_ber_count),
				.pld_10g_rx_rd_en(in_pld_10g_rx_rd_en),
				.pld_8g_a1a2_size(in_pld_8g_a1a2_size),
				.pld_8g_bitloc_rev_en(in_pld_8g_bitloc_rev_en),
				.pld_8g_byte_rev_en(in_pld_8g_byte_rev_en),
				.pld_8g_encdt(in_pld_8g_encdt),
				.pld_8g_g3_rx_pld_rst_n(in_pld_8g_g3_rx_pld_rst_n),
				.pld_8g_rdenable_rx(in_pld_8g_rdenable_rx),
				.pld_8g_rxpolarity(in_pld_8g_rxpolarity),
				.pld_8g_wrdisable_rx(in_pld_8g_wrdisable_rx),
				.pld_bitslip(in_pld_bitslip),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_rxpma_rstb(in_pld_pma_rxpma_rstb),
				.pld_pmaif_rx_pld_rst_n(in_pld_pmaif_rx_pld_rst_n),
				.pld_pmaif_rxclkslip(in_pld_pmaif_rxclkslip),
				.pld_polinv_rx(in_pld_polinv_rx),
				.pld_rx_clk(in_pld_rx_clk),
				.pld_rx_prbs_err_clr(in_pld_rx_prbs_err_clr),
				.pld_syncsm_en(in_pld_syncsm_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.int_pldif_pmaif_rx_pld_clk(),
				.pld_8g_wa_boundary_txclk_fastreg(),
				.pld_8g_wa_boundary_txclk_reg(),
				.pld_bitslip_10g_txclk_reg(),
				.pld_bitslip_8g_txclk_reg(),
				.pld_bitslip_rxclk_parallel_loopback_reg(),
				.pld_bitslip_rxclk_reg(),
				.pld_pcs_rx_clk_out_pcsdirect_wire(),
				.pld_pma_rx_clk_out_10g_or_pcsdirect_wire(),
				.pld_pma_rx_clk_out_8g_wire(),
				.pld_pmaif_rx_pld_rst_n_reg(),
				.pld_pmaif_tx_pld_rst_n_txclk_reg(),
				.pld_polinv_rx_reg(),
				.pld_rx_clk_fifo(),
				.pld_rx_control_fifo(),
				.pld_rx_control_pcsdirect_reg(),
				.pld_rx_data_fifo(),
				.pld_rx_data_pcsdirect_reg(),
				.pld_rx_prbs_done_reg(),
				.pld_rx_prbs_done_txclk_reg(),
				.pld_rx_prbs_err_clr_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_clr_reg(),
				.pld_rx_prbs_err_disprbs_reg(),
				.pld_rx_prbs_err_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_reg(),
				.pma_rx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_data[50:0] = 51'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3:0] = 4'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_control[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_data[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pcs_pma_interface
			twentynm_hssi_tx_pcs_pma_interface #(
				.bypass_pma_txelecidle(hssi_tx_pcs_pma_interface_bypass_pma_txelecidle),
				.channel_operation_mode(hssi_tx_pcs_pma_interface_channel_operation_mode),
				.lpbk_en(hssi_tx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_tx_pcs_pma_interface_master_clk_sel),
				.pcie_sub_prot_mode_tx(hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx),
				.pldif_datawidth_mode(hssi_tx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_tx(hssi_tx_pcs_pma_interface_pma_dw_tx),
				.pma_if_dft_en(hssi_tx_pcs_pma_interface_pma_if_dft_en),
				.pmagate_en(hssi_tx_pcs_pma_interface_pmagate_en),
				.prbs9_dwidth(hssi_tx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_tx_pcs_pma_interface_prbs_clken),
				.prbs_gen_pat(hssi_tx_pcs_pma_interface_prbs_gen_pat),
				.prot_mode_tx(hssi_tx_pcs_pma_interface_prot_mode_tx),
				.reconfig_settings(hssi_tx_pcs_pma_interface_reconfig_settings),
				.silicon_rev( "20nm4" ),       //PARAM_HIDE
				.sq_wave_num(hssi_tx_pcs_pma_interface_sq_wave_num),
				.sqwgen_clken(hssi_tx_pcs_pma_interface_sqwgen_clken),
				.sup_mode(hssi_tx_pcs_pma_interface_sup_mode),
				.tx_dyn_polarity_inversion(hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion),
				.tx_pma_data_sel(hssi_tx_pcs_pma_interface_tx_pma_data_sel),
				.tx_static_polarity_inversion(hssi_tx_pcs_pma_interface_tx_static_polarity_inversion),
				.uhsif_cnt_step_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock),
				.uhsif_cnt_thresh_filt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value),
				.uhsif_cnt_thresh_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock),
				.uhsif_dcn_test_update_period(hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period),
				.uhsif_dcn_testmode_enable(hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable),
				.uhsif_dead_zone_count_thresh(hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh),
				.uhsif_dead_zone_detection_enable(hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable),
				.uhsif_dead_zone_obser_window(hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window),
				.uhsif_dead_zone_skip_size(hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size),
				.uhsif_delay_cell_index_sel(hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel),
				.uhsif_delay_cell_margin(hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin),
				.uhsif_delay_cell_static_index_value(hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value),
				.uhsif_dft_dead_zone_control(hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control),
				.uhsif_dft_up_filt_control(hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control),
				.uhsif_enable(hssi_tx_pcs_pma_interface_uhsif_enable),
				.uhsif_lock_det_segsz_after_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock),
				.uhsif_lock_det_segsz_before_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock),
				.uhsif_lock_det_thresh_cnt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value),
				.uhsif_lock_det_thresh_cnt_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value),
				.uhsif_lock_det_thresh_diff_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value),
				.uhsif_lock_det_thresh_diff_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value)
			) inst_twentynm_hssi_tx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.int_pmaif_8g_txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.int_pmaif_pldif_tx_clkdiv(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pmaif_pldif_tx_clkdiv_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pmaif_pldif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.int_pmaif_pldif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.int_tx_dft_obsrv_clk(w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk),
				.pma_tx_elec_idle(w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle),
				.pma_tx_pma_data(w_hssi_tx_pcs_pma_interface_pma_tx_pma_data),
				.pma_txpma_rstb(w_hssi_tx_pcs_pma_interface_pma_txpma_rstb),
				.tx_pma_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback),
				.tx_pma_uhsif_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback),
				.tx_prbs_gen_test(w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test),
				.uhsif_test_out_1(w_hssi_tx_pcs_pma_interface_uhsif_test_out_1),
				.uhsif_test_out_2(w_hssi_tx_pcs_pma_interface_uhsif_test_out_2),
				.uhsif_test_out_3(w_hssi_tx_pcs_pma_interface_uhsif_test_out_3),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.int_pmaif_10g_tx_pma_data({w_hssi_10g_tx_pcs_tx_pma_data[63], w_hssi_10g_tx_pcs_tx_pma_data[62], w_hssi_10g_tx_pcs_tx_pma_data[61], w_hssi_10g_tx_pcs_tx_pma_data[60], w_hssi_10g_tx_pcs_tx_pma_data[59], w_hssi_10g_tx_pcs_tx_pma_data[58], w_hssi_10g_tx_pcs_tx_pma_data[57], w_hssi_10g_tx_pcs_tx_pma_data[56], w_hssi_10g_tx_pcs_tx_pma_data[55], w_hssi_10g_tx_pcs_tx_pma_data[54], w_hssi_10g_tx_pcs_tx_pma_data[53], w_hssi_10g_tx_pcs_tx_pma_data[52], w_hssi_10g_tx_pcs_tx_pma_data[51], w_hssi_10g_tx_pcs_tx_pma_data[50], w_hssi_10g_tx_pcs_tx_pma_data[49], w_hssi_10g_tx_pcs_tx_pma_data[48], w_hssi_10g_tx_pcs_tx_pma_data[47], w_hssi_10g_tx_pcs_tx_pma_data[46], w_hssi_10g_tx_pcs_tx_pma_data[45], w_hssi_10g_tx_pcs_tx_pma_data[44], w_hssi_10g_tx_pcs_tx_pma_data[43], w_hssi_10g_tx_pcs_tx_pma_data[42], w_hssi_10g_tx_pcs_tx_pma_data[41], w_hssi_10g_tx_pcs_tx_pma_data[40], w_hssi_10g_tx_pcs_tx_pma_data[39], w_hssi_10g_tx_pcs_tx_pma_data[38], w_hssi_10g_tx_pcs_tx_pma_data[37], w_hssi_10g_tx_pcs_tx_pma_data[36], w_hssi_10g_tx_pcs_tx_pma_data[35], w_hssi_10g_tx_pcs_tx_pma_data[34], w_hssi_10g_tx_pcs_tx_pma_data[33], w_hssi_10g_tx_pcs_tx_pma_data[32], w_hssi_10g_tx_pcs_tx_pma_data[31], w_hssi_10g_tx_pcs_tx_pma_data[30], w_hssi_10g_tx_pcs_tx_pma_data[29], w_hssi_10g_tx_pcs_tx_pma_data[28], w_hssi_10g_tx_pcs_tx_pma_data[27], w_hssi_10g_tx_pcs_tx_pma_data[26], w_hssi_10g_tx_pcs_tx_pma_data[25], w_hssi_10g_tx_pcs_tx_pma_data[24], w_hssi_10g_tx_pcs_tx_pma_data[23], w_hssi_10g_tx_pcs_tx_pma_data[22], w_hssi_10g_tx_pcs_tx_pma_data[21], w_hssi_10g_tx_pcs_tx_pma_data[20], w_hssi_10g_tx_pcs_tx_pma_data[19], w_hssi_10g_tx_pcs_tx_pma_data[18], w_hssi_10g_tx_pcs_tx_pma_data[17], w_hssi_10g_tx_pcs_tx_pma_data[16], w_hssi_10g_tx_pcs_tx_pma_data[15], w_hssi_10g_tx_pcs_tx_pma_data[14], w_hssi_10g_tx_pcs_tx_pma_data[13], w_hssi_10g_tx_pcs_tx_pma_data[12], w_hssi_10g_tx_pcs_tx_pma_data[11], w_hssi_10g_tx_pcs_tx_pma_data[10], w_hssi_10g_tx_pcs_tx_pma_data[9], w_hssi_10g_tx_pcs_tx_pma_data[8], w_hssi_10g_tx_pcs_tx_pma_data[7], w_hssi_10g_tx_pcs_tx_pma_data[6], w_hssi_10g_tx_pcs_tx_pma_data[5], w_hssi_10g_tx_pcs_tx_pma_data[4], w_hssi_10g_tx_pcs_tx_pma_data[3], w_hssi_10g_tx_pcs_tx_pma_data[2], w_hssi_10g_tx_pcs_tx_pma_data[1], w_hssi_10g_tx_pcs_tx_pma_data[0]}),
				.int_pmaif_10g_tx_pma_data_gate_val({w_hssi_10g_tx_pcs_tx_pma_gating_val[63], w_hssi_10g_tx_pcs_tx_pma_gating_val[62], w_hssi_10g_tx_pcs_tx_pma_gating_val[61], w_hssi_10g_tx_pcs_tx_pma_gating_val[60], w_hssi_10g_tx_pcs_tx_pma_gating_val[59], w_hssi_10g_tx_pcs_tx_pma_gating_val[58], w_hssi_10g_tx_pcs_tx_pma_gating_val[57], w_hssi_10g_tx_pcs_tx_pma_gating_val[56], w_hssi_10g_tx_pcs_tx_pma_gating_val[55], w_hssi_10g_tx_pcs_tx_pma_gating_val[54], w_hssi_10g_tx_pcs_tx_pma_gating_val[53], w_hssi_10g_tx_pcs_tx_pma_gating_val[52], w_hssi_10g_tx_pcs_tx_pma_gating_val[51], w_hssi_10g_tx_pcs_tx_pma_gating_val[50], w_hssi_10g_tx_pcs_tx_pma_gating_val[49], w_hssi_10g_tx_pcs_tx_pma_gating_val[48], w_hssi_10g_tx_pcs_tx_pma_gating_val[47], w_hssi_10g_tx_pcs_tx_pma_gating_val[46], w_hssi_10g_tx_pcs_tx_pma_gating_val[45], w_hssi_10g_tx_pcs_tx_pma_gating_val[44], w_hssi_10g_tx_pcs_tx_pma_gating_val[43], w_hssi_10g_tx_pcs_tx_pma_gating_val[42], w_hssi_10g_tx_pcs_tx_pma_gating_val[41], w_hssi_10g_tx_pcs_tx_pma_gating_val[40], w_hssi_10g_tx_pcs_tx_pma_gating_val[39], w_hssi_10g_tx_pcs_tx_pma_gating_val[38], w_hssi_10g_tx_pcs_tx_pma_gating_val[37], w_hssi_10g_tx_pcs_tx_pma_gating_val[36], w_hssi_10g_tx_pcs_tx_pma_gating_val[35], w_hssi_10g_tx_pcs_tx_pma_gating_val[34], w_hssi_10g_tx_pcs_tx_pma_gating_val[33], w_hssi_10g_tx_pcs_tx_pma_gating_val[32], w_hssi_10g_tx_pcs_tx_pma_gating_val[31], w_hssi_10g_tx_pcs_tx_pma_gating_val[30], w_hssi_10g_tx_pcs_tx_pma_gating_val[29], w_hssi_10g_tx_pcs_tx_pma_gating_val[28], w_hssi_10g_tx_pcs_tx_pma_gating_val[27], w_hssi_10g_tx_pcs_tx_pma_gating_val[26], w_hssi_10g_tx_pcs_tx_pma_gating_val[25], w_hssi_10g_tx_pcs_tx_pma_gating_val[24], w_hssi_10g_tx_pcs_tx_pma_gating_val[23], w_hssi_10g_tx_pcs_tx_pma_gating_val[22], w_hssi_10g_tx_pcs_tx_pma_gating_val[21], w_hssi_10g_tx_pcs_tx_pma_gating_val[20], w_hssi_10g_tx_pcs_tx_pma_gating_val[19], w_hssi_10g_tx_pcs_tx_pma_gating_val[18], w_hssi_10g_tx_pcs_tx_pma_gating_val[17], w_hssi_10g_tx_pcs_tx_pma_gating_val[16], w_hssi_10g_tx_pcs_tx_pma_gating_val[15], w_hssi_10g_tx_pcs_tx_pma_gating_val[14], w_hssi_10g_tx_pcs_tx_pma_gating_val[13], w_hssi_10g_tx_pcs_tx_pma_gating_val[12], w_hssi_10g_tx_pcs_tx_pma_gating_val[11], w_hssi_10g_tx_pcs_tx_pma_gating_val[10], w_hssi_10g_tx_pcs_tx_pma_gating_val[9], w_hssi_10g_tx_pcs_tx_pma_gating_val[8], w_hssi_10g_tx_pcs_tx_pma_gating_val[7], w_hssi_10g_tx_pcs_tx_pma_gating_val[6], w_hssi_10g_tx_pcs_tx_pma_gating_val[5], w_hssi_10g_tx_pcs_tx_pma_gating_val[4], w_hssi_10g_tx_pcs_tx_pma_gating_val[3], w_hssi_10g_tx_pcs_tx_pma_gating_val[2], w_hssi_10g_tx_pcs_tx_pma_gating_val[1], w_hssi_10g_tx_pcs_tx_pma_gating_val[0]}),
				.int_pmaif_8g_pudr({w_hssi_8g_tx_pcs_dataout[19], w_hssi_8g_tx_pcs_dataout[18], w_hssi_8g_tx_pcs_dataout[17], w_hssi_8g_tx_pcs_dataout[16], w_hssi_8g_tx_pcs_dataout[15], w_hssi_8g_tx_pcs_dataout[14], w_hssi_8g_tx_pcs_dataout[13], w_hssi_8g_tx_pcs_dataout[12], w_hssi_8g_tx_pcs_dataout[11], w_hssi_8g_tx_pcs_dataout[10], w_hssi_8g_tx_pcs_dataout[9], w_hssi_8g_tx_pcs_dataout[8], w_hssi_8g_tx_pcs_dataout[7], w_hssi_8g_tx_pcs_dataout[6], w_hssi_8g_tx_pcs_dataout[5], w_hssi_8g_tx_pcs_dataout[4], w_hssi_8g_tx_pcs_dataout[3], w_hssi_8g_tx_pcs_dataout[2], w_hssi_8g_tx_pcs_dataout[1], w_hssi_8g_tx_pcs_dataout[0]}),
				.int_pmaif_8g_tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.int_pmaif_8g_tx_elec_idle(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_pma_data_out({w_hssi_gen3_tx_pcs_data_out[31], w_hssi_gen3_tx_pcs_data_out[30], w_hssi_gen3_tx_pcs_data_out[29], w_hssi_gen3_tx_pcs_data_out[28], w_hssi_gen3_tx_pcs_data_out[27], w_hssi_gen3_tx_pcs_data_out[26], w_hssi_gen3_tx_pcs_data_out[25], w_hssi_gen3_tx_pcs_data_out[24], w_hssi_gen3_tx_pcs_data_out[23], w_hssi_gen3_tx_pcs_data_out[22], w_hssi_gen3_tx_pcs_data_out[21], w_hssi_gen3_tx_pcs_data_out[20], w_hssi_gen3_tx_pcs_data_out[19], w_hssi_gen3_tx_pcs_data_out[18], w_hssi_gen3_tx_pcs_data_out[17], w_hssi_gen3_tx_pcs_data_out[16], w_hssi_gen3_tx_pcs_data_out[15], w_hssi_gen3_tx_pcs_data_out[14], w_hssi_gen3_tx_pcs_data_out[13], w_hssi_gen3_tx_pcs_data_out[12], w_hssi_gen3_tx_pcs_data_out[11], w_hssi_gen3_tx_pcs_data_out[10], w_hssi_gen3_tx_pcs_data_out[9], w_hssi_gen3_tx_pcs_data_out[8], w_hssi_gen3_tx_pcs_data_out[7], w_hssi_gen3_tx_pcs_data_out[6], w_hssi_gen3_tx_pcs_data_out[5], w_hssi_gen3_tx_pcs_data_out[4], w_hssi_gen3_tx_pcs_data_out[3], w_hssi_gen3_tx_pcs_data_out[2], w_hssi_gen3_tx_pcs_data_out[1], w_hssi_gen3_tx_pcs_data_out[0]}),
				.int_pmaif_g3_pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.int_pmaif_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pmaif_pldif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pmaif_pldif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0]}),
				.int_pmaif_pldif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pmaif_pldif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.int_pmaif_pldif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pmaif_pldif_uhsif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0]}),
				.pma_tx_clkdiv_user(in_pma_tx_clkdiv_user),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.refclk_dig_uhsif(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.uhsif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.uhsif_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				
				// UNUSED
				.avmm_user_dataout(),
				.write_en(),
				.write_en_ack()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4:0] = 5'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_txpma_rstb = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pld_pcs_interface
			twentynm_hssi_tx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx),
				.hd_10g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx),
				.hd_10g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx),
				.hd_10g_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx),
				.hd_10g_lpbk_en(hssi_tx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx),
				.hd_10g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx),
				.hd_10g_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx),
				.hd_8g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx),
				.hd_8g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx),
				.hd_8g_hip_mode(hssi_tx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_tx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx),
				.hd_8g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx),
				.hd_chnl_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx),
				.hd_chnl_frequency_rules_en(hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_tx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_tx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx),
				.hd_chnl_lpbk_en(hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx),
				.hd_chnl_pld_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz),
				.hd_chnl_pld_uhsif_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz),
				.hd_chnl_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx),
				.hd_chnl_pma_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz),
				.hd_chnl_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx),
				.hd_chnl_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx),
				.hd_fifo_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx),
				.hd_fifo_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx),
				.hd_g3_prot_mode(hssi_tx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx),
				.hd_krfec_lpbk_en(hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx),
				.hd_pldif_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx),
				.hd_pmaif_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_ctrl_plane_bonding(hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding),
				.hd_pmaif_lpbk_en(hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx),
				.hd_pmaif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx),
				.hd_pmaif_sim_mode(hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_tx_clk_out_sel(hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel),
				.pcs_tx_clk_source(hssi_tx_pld_pcs_interface_pcs_tx_clk_source),
				.pcs_tx_data_source(hssi_tx_pld_pcs_interface_pcs_tx_data_source),
				.pcs_tx_delay1_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en),
				.pcs_tx_delay1_clk_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel),
				.pcs_tx_delay1_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl),
				.pcs_tx_delay1_data_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel),
				.pcs_tx_delay2_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en),
				.pcs_tx_delay2_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl),
				.pcs_tx_output_sel(hssi_tx_pld_pcs_interface_pcs_tx_output_sel),
				.reconfig_settings(hssi_tx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm4" )       //PARAM_HIDE
			) inst_twentynm_hssi_tx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pld_pcs_interface_blockselect),
				.hip_tx_clk(w_hssi_tx_pld_pcs_interface_hip_tx_clk),
				.int_pldif_10g_tx_bitslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip),
				.int_pldif_10g_tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.int_pldif_10g_tx_control(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control),
				.int_pldif_10g_tx_control_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg),
				.int_pldif_10g_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data),
				.int_pldif_10g_tx_data_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg),
				.int_pldif_10g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.int_pldif_10g_tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.int_pldif_10g_tx_diag_status(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status),
				.int_pldif_10g_tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.int_pldif_10g_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.int_pldif_10g_tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				.int_pldif_8g_pld_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.int_pldif_8g_powerdown(w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown),
				.int_pldif_8g_rddisable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.int_pldif_8g_rev_loopbk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.int_pldif_8g_tx_blk_start(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start),
				.int_pldif_8g_tx_boundary_sel(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel),
				.int_pldif_8g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid),
				.int_pldif_8g_tx_sync_hdr(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr),
				.int_pldif_8g_txd(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd),
				.int_pldif_8g_txd_fast_reg(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg),
				.int_pldif_8g_txdeemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.int_pldif_8g_txdetectrxloopback(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.int_pldif_8g_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.int_pldif_8g_txmargin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin),
				.int_pldif_8g_txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.int_pldif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.int_pldif_8g_wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				.int_pldif_pmaif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pldif_pmaif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pldif_pmaif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data),
				.int_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pldif_pmaif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pldif_pmaif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pldif_pmaif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pldif_pmaif_uhsif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data),
				.pld_10g_krfec_tx_frame(w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame),
				.pld_10g_tx_burst_en_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe),
				.pld_10g_tx_empty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty),
				.pld_10g_tx_fifo_num(w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num),
				.pld_10g_tx_full(w_hssi_tx_pld_pcs_interface_pld_10g_tx_full),
				.pld_10g_tx_pempty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty),
				.pld_10g_tx_pfull(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull),
				.pld_10g_tx_wordslip_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe),
				.pld_8g_empty_tx(w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx),
				.pld_8g_full_tx(w_hssi_tx_pld_pcs_interface_pld_8g_full_tx),
				.pld_krfec_tx_alignment(w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment),
				.pld_pcs_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out),
				.pld_pma_clkdiv_tx_user(w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user),
				.pld_pma_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out),
				.pld_uhsif_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.hip_tx_data({in_hip_tx_data[63], in_hip_tx_data[62], in_hip_tx_data[61], in_hip_tx_data[60], in_hip_tx_data[59], in_hip_tx_data[58], in_hip_tx_data[57], in_hip_tx_data[56], in_hip_tx_data[55], in_hip_tx_data[54], in_hip_tx_data[53], in_hip_tx_data[52], in_hip_tx_data[51], in_hip_tx_data[50], in_hip_tx_data[49], in_hip_tx_data[48], in_hip_tx_data[47], in_hip_tx_data[46], in_hip_tx_data[45], in_hip_tx_data[44], in_hip_tx_data[43], in_hip_tx_data[42], in_hip_tx_data[41], in_hip_tx_data[40], in_hip_tx_data[39], in_hip_tx_data[38], in_hip_tx_data[37], in_hip_tx_data[36], in_hip_tx_data[35], in_hip_tx_data[34], in_hip_tx_data[33], in_hip_tx_data[32], in_hip_tx_data[31], in_hip_tx_data[30], in_hip_tx_data[29], in_hip_tx_data[28], in_hip_tx_data[27], in_hip_tx_data[26], in_hip_tx_data[25], in_hip_tx_data[24], in_hip_tx_data[23], in_hip_tx_data[22], in_hip_tx_data[21], in_hip_tx_data[20], in_hip_tx_data[19], in_hip_tx_data[18], in_hip_tx_data[17], in_hip_tx_data[16], in_hip_tx_data[15], in_hip_tx_data[14], in_hip_tx_data[13], in_hip_tx_data[12], in_hip_tx_data[11], in_hip_tx_data[10], in_hip_tx_data[9], in_hip_tx_data[8], in_hip_tx_data[7], in_hip_tx_data[6], in_hip_tx_data[5], in_hip_tx_data[4], in_hip_tx_data[3], in_hip_tx_data[2], in_hip_tx_data[1], in_hip_tx_data[0]}),
				.int_pldif_10g_tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.int_pldif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.int_pldif_10g_tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_10g_tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.int_pldif_10g_tx_fifo_num({w_hssi_10g_tx_pcs_tx_fifo_num[3], w_hssi_10g_tx_pcs_tx_fifo_num[2], w_hssi_10g_tx_pcs_tx_fifo_num[1], w_hssi_10g_tx_pcs_tx_fifo_num[0]}),
				.int_pldif_10g_tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.int_pldif_10g_tx_full(w_hssi_10g_tx_pcs_tx_full),
				.int_pldif_10g_tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.int_pldif_10g_tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.int_pldif_10g_tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				.int_pldif_8g_empty_tx(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.int_pldif_8g_full_tx(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.int_pldif_8g_tx_clk_out(w_hssi_8g_tx_pcs_clk_out),
				.int_pldif_8g_tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_krfec_tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.int_pldif_krfec_tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.int_pldif_pmaif_clkdiv_tx(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pldif_pmaif_clkdiv_tx_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pldif_pmaif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.pld_10g_krfec_tx_pld_rst_n(in_pld_10g_krfec_tx_pld_rst_n),
				.pld_10g_tx_bitslip({in_pld_10g_tx_bitslip[6], in_pld_10g_tx_bitslip[5], in_pld_10g_tx_bitslip[4], in_pld_10g_tx_bitslip[3], in_pld_10g_tx_bitslip[2], in_pld_10g_tx_bitslip[1], in_pld_10g_tx_bitslip[0]}),
				.pld_10g_tx_burst_en(in_pld_10g_tx_burst_en),
				.pld_10g_tx_data_valid(in_pld_10g_tx_data_valid),
				.pld_10g_tx_diag_status({in_pld_10g_tx_diag_status[1], in_pld_10g_tx_diag_status[0]}),
				.pld_10g_tx_wordslip(in_pld_10g_tx_wordslip),
				.pld_8g_g3_tx_pld_rst_n(in_pld_8g_g3_tx_pld_rst_n),
				.pld_8g_rddisable_tx(in_pld_8g_rddisable_tx),
				.pld_8g_tx_boundary_sel({in_pld_8g_tx_boundary_sel[4], in_pld_8g_tx_boundary_sel[3], in_pld_8g_tx_boundary_sel[2], in_pld_8g_tx_boundary_sel[1], in_pld_8g_tx_boundary_sel[0]}),
				.pld_8g_wrenable_tx(in_pld_8g_wrenable_tx),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_txpma_rstb(in_pld_pma_txpma_rstb),
				.pld_pmaif_tx_pld_rst_n(in_pld_pmaif_tx_pld_rst_n),
				.pld_polinv_tx(in_pld_polinv_tx),
				.pld_tx_clk(in_pld_tx_clk),
				.pld_tx_control({in_pld_tx_control[17], in_pld_tx_control[16], in_pld_tx_control[15], in_pld_tx_control[14], in_pld_tx_control[13], in_pld_tx_control[12], in_pld_tx_control[11], in_pld_tx_control[10], in_pld_tx_control[9], in_pld_tx_control[8], in_pld_tx_control[7], in_pld_tx_control[6], in_pld_tx_control[5], in_pld_tx_control[4], in_pld_tx_control[3], in_pld_tx_control[2], in_pld_tx_control[1], in_pld_tx_control[0]}),
				.pld_tx_data({in_pld_tx_data[127], in_pld_tx_data[126], in_pld_tx_data[125], in_pld_tx_data[124], in_pld_tx_data[123], in_pld_tx_data[122], in_pld_tx_data[121], in_pld_tx_data[120], in_pld_tx_data[119], in_pld_tx_data[118], in_pld_tx_data[117], in_pld_tx_data[116], in_pld_tx_data[115], in_pld_tx_data[114], in_pld_tx_data[113], in_pld_tx_data[112], in_pld_tx_data[111], in_pld_tx_data[110], in_pld_tx_data[109], in_pld_tx_data[108], in_pld_tx_data[107], in_pld_tx_data[106], in_pld_tx_data[105], in_pld_tx_data[104], in_pld_tx_data[103], in_pld_tx_data[102], in_pld_tx_data[101], in_pld_tx_data[100], in_pld_tx_data[99], in_pld_tx_data[98], in_pld_tx_data[97], in_pld_tx_data[96], in_pld_tx_data[95], in_pld_tx_data[94], in_pld_tx_data[93], in_pld_tx_data[92], in_pld_tx_data[91], in_pld_tx_data[90], in_pld_tx_data[89], in_pld_tx_data[88], in_pld_tx_data[87], in_pld_tx_data[86], in_pld_tx_data[85], in_pld_tx_data[84], in_pld_tx_data[83], in_pld_tx_data[82], in_pld_tx_data[81], in_pld_tx_data[80], in_pld_tx_data[79], in_pld_tx_data[78], in_pld_tx_data[77], in_pld_tx_data[76], in_pld_tx_data[75], in_pld_tx_data[74], in_pld_tx_data[73], in_pld_tx_data[72], in_pld_tx_data[71], in_pld_tx_data[70], in_pld_tx_data[69], in_pld_tx_data[68], in_pld_tx_data[67], in_pld_tx_data[66], in_pld_tx_data[65], in_pld_tx_data[64], in_pld_tx_data[63], in_pld_tx_data[62], in_pld_tx_data[61], in_pld_tx_data[60], in_pld_tx_data[59], in_pld_tx_data[58], in_pld_tx_data[57], in_pld_tx_data[56], in_pld_tx_data[55], in_pld_tx_data[54], in_pld_tx_data[53], in_pld_tx_data[52], in_pld_tx_data[51], in_pld_tx_data[50], in_pld_tx_data[49], in_pld_tx_data[48], in_pld_tx_data[47], in_pld_tx_data[46], in_pld_tx_data[45], in_pld_tx_data[44], in_pld_tx_data[43], in_pld_tx_data[42], in_pld_tx_data[41], in_pld_tx_data[40], in_pld_tx_data[39], in_pld_tx_data[38], in_pld_tx_data[37], in_pld_tx_data[36], in_pld_tx_data[35], in_pld_tx_data[34], in_pld_tx_data[33], in_pld_tx_data[32], in_pld_tx_data[31], in_pld_tx_data[30], in_pld_tx_data[29], in_pld_tx_data[28], in_pld_tx_data[27], in_pld_tx_data[26], in_pld_tx_data[25], in_pld_tx_data[24], in_pld_tx_data[23], in_pld_tx_data[22], in_pld_tx_data[21], in_pld_tx_data[20], in_pld_tx_data[19], in_pld_tx_data[18], in_pld_tx_data[17], in_pld_tx_data[16], in_pld_tx_data[15], in_pld_tx_data[14], in_pld_tx_data[13], in_pld_tx_data[12], in_pld_tx_data[11], in_pld_tx_data[10], in_pld_tx_data[9], in_pld_tx_data[8], in_pld_tx_data[7], in_pld_tx_data[6], in_pld_tx_data[5], in_pld_tx_data[4], in_pld_tx_data[3], in_pld_tx_data[2], in_pld_tx_data[1], in_pld_tx_data[0]}),
				.pld_txelecidle(in_pld_txelecidle),
				.pld_uhsif_tx_clk(in_pld_uhsif_tx_clk),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.hip_clk_out_div_by_2_wire(),
				.hip_clk_out_wire(),
				.int_pldif_pmaif_tx_pld_clk(),
				.pld_10g_tx_burst_en_exe_10g_fastreg(),
				.pld_10g_tx_burst_en_exe_plddirect_reg(),
				.pld_10g_tx_data_valid_2ff_delay1_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay3_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg(),
				.pld_10g_tx_data_valid_fastreg(),
				.pld_10g_tx_data_valid_plddirect_fastreg(),
				.pld_pcs_tx_clk_out_pma_wire(),
				.pld_pma_tx_clk_out_wire(),
				.pld_pmaif_tx_pld_rst_n_reg(),
				.pld_polinv_tx_10g_pcsdirect_reg(),
				.pld_polinv_tx_8g_reg(),
				.pld_polinv_tx_pat_reg(),
				.pld_tx_clk_fifo(),
				.pld_tx_control_fifo(),
				.pld_tx_control_hi_10g_reg(),
				.pld_tx_control_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_10g_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_8g_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_control_lo_plddirect_fastreg(),
				.pld_tx_control_lo_plddirect_reg(),
				.pld_tx_data_hi_reg(),
				.pld_tx_data_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_10g_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_8g_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_data_lo_plddirect_fastreg(),
				.pld_tx_data_lo_plddirect_reg(),
				.pld_uhsif_reg(),
				.pma_tx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_hip_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6:0] = 7'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17:0] = 18'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8:0] = 9'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127:0] = 128'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4:0] = 5'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2:0] = 3'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_full = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_full_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out = 1'b0;
		end // if not generate
		
		//output assignments
		assign out_avmmreaddata_hssi_10g_rx_pcs = {w_hssi_10g_rx_pcs_avmmreaddata[7], w_hssi_10g_rx_pcs_avmmreaddata[6], w_hssi_10g_rx_pcs_avmmreaddata[5], w_hssi_10g_rx_pcs_avmmreaddata[4], w_hssi_10g_rx_pcs_avmmreaddata[3], w_hssi_10g_rx_pcs_avmmreaddata[2], w_hssi_10g_rx_pcs_avmmreaddata[1], w_hssi_10g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_10g_tx_pcs = {w_hssi_10g_tx_pcs_avmmreaddata[7], w_hssi_10g_tx_pcs_avmmreaddata[6], w_hssi_10g_tx_pcs_avmmreaddata[5], w_hssi_10g_tx_pcs_avmmreaddata[4], w_hssi_10g_tx_pcs_avmmreaddata[3], w_hssi_10g_tx_pcs_avmmreaddata[2], w_hssi_10g_tx_pcs_avmmreaddata[1], w_hssi_10g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_rx_pcs = {w_hssi_8g_rx_pcs_avmmreaddata[7], w_hssi_8g_rx_pcs_avmmreaddata[6], w_hssi_8g_rx_pcs_avmmreaddata[5], w_hssi_8g_rx_pcs_avmmreaddata[4], w_hssi_8g_rx_pcs_avmmreaddata[3], w_hssi_8g_rx_pcs_avmmreaddata[2], w_hssi_8g_rx_pcs_avmmreaddata[1], w_hssi_8g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_tx_pcs = {w_hssi_8g_tx_pcs_avmmreaddata[7], w_hssi_8g_tx_pcs_avmmreaddata[6], w_hssi_8g_tx_pcs_avmmreaddata[5], w_hssi_8g_tx_pcs_avmmreaddata[4], w_hssi_8g_tx_pcs_avmmreaddata[3], w_hssi_8g_tx_pcs_avmmreaddata[2], w_hssi_8g_tx_pcs_avmmreaddata[1], w_hssi_8g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pcs_pma_interface = {w_hssi_common_pcs_pma_interface_avmmreaddata[7], w_hssi_common_pcs_pma_interface_avmmreaddata[6], w_hssi_common_pcs_pma_interface_avmmreaddata[5], w_hssi_common_pcs_pma_interface_avmmreaddata[4], w_hssi_common_pcs_pma_interface_avmmreaddata[3], w_hssi_common_pcs_pma_interface_avmmreaddata[2], w_hssi_common_pcs_pma_interface_avmmreaddata[1], w_hssi_common_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pld_pcs_interface = {w_hssi_common_pld_pcs_interface_avmmreaddata[7], w_hssi_common_pld_pcs_interface_avmmreaddata[6], w_hssi_common_pld_pcs_interface_avmmreaddata[5], w_hssi_common_pld_pcs_interface_avmmreaddata[4], w_hssi_common_pld_pcs_interface_avmmreaddata[3], w_hssi_common_pld_pcs_interface_avmmreaddata[2], w_hssi_common_pld_pcs_interface_avmmreaddata[1], w_hssi_common_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_rx_pcs = {w_hssi_fifo_rx_pcs_avmmreaddata[7], w_hssi_fifo_rx_pcs_avmmreaddata[6], w_hssi_fifo_rx_pcs_avmmreaddata[5], w_hssi_fifo_rx_pcs_avmmreaddata[4], w_hssi_fifo_rx_pcs_avmmreaddata[3], w_hssi_fifo_rx_pcs_avmmreaddata[2], w_hssi_fifo_rx_pcs_avmmreaddata[1], w_hssi_fifo_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_tx_pcs = {w_hssi_fifo_tx_pcs_avmmreaddata[7], w_hssi_fifo_tx_pcs_avmmreaddata[6], w_hssi_fifo_tx_pcs_avmmreaddata[5], w_hssi_fifo_tx_pcs_avmmreaddata[4], w_hssi_fifo_tx_pcs_avmmreaddata[3], w_hssi_fifo_tx_pcs_avmmreaddata[2], w_hssi_fifo_tx_pcs_avmmreaddata[1], w_hssi_fifo_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_rx_pcs = {w_hssi_gen3_rx_pcs_avmmreaddata[7], w_hssi_gen3_rx_pcs_avmmreaddata[6], w_hssi_gen3_rx_pcs_avmmreaddata[5], w_hssi_gen3_rx_pcs_avmmreaddata[4], w_hssi_gen3_rx_pcs_avmmreaddata[3], w_hssi_gen3_rx_pcs_avmmreaddata[2], w_hssi_gen3_rx_pcs_avmmreaddata[1], w_hssi_gen3_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_tx_pcs = {w_hssi_gen3_tx_pcs_avmmreaddata[7], w_hssi_gen3_tx_pcs_avmmreaddata[6], w_hssi_gen3_tx_pcs_avmmreaddata[5], w_hssi_gen3_tx_pcs_avmmreaddata[4], w_hssi_gen3_tx_pcs_avmmreaddata[3], w_hssi_gen3_tx_pcs_avmmreaddata[2], w_hssi_gen3_tx_pcs_avmmreaddata[1], w_hssi_gen3_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_rx_pcs = {w_hssi_krfec_rx_pcs_avmmreaddata[7], w_hssi_krfec_rx_pcs_avmmreaddata[6], w_hssi_krfec_rx_pcs_avmmreaddata[5], w_hssi_krfec_rx_pcs_avmmreaddata[4], w_hssi_krfec_rx_pcs_avmmreaddata[3], w_hssi_krfec_rx_pcs_avmmreaddata[2], w_hssi_krfec_rx_pcs_avmmreaddata[1], w_hssi_krfec_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_tx_pcs = {w_hssi_krfec_tx_pcs_avmmreaddata[7], w_hssi_krfec_tx_pcs_avmmreaddata[6], w_hssi_krfec_tx_pcs_avmmreaddata[5], w_hssi_krfec_tx_pcs_avmmreaddata[4], w_hssi_krfec_tx_pcs_avmmreaddata[3], w_hssi_krfec_tx_pcs_avmmreaddata[2], w_hssi_krfec_tx_pcs_avmmreaddata[1], w_hssi_krfec_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen1_2 = {w_hssi_pipe_gen1_2_avmmreaddata[7], w_hssi_pipe_gen1_2_avmmreaddata[6], w_hssi_pipe_gen1_2_avmmreaddata[5], w_hssi_pipe_gen1_2_avmmreaddata[4], w_hssi_pipe_gen1_2_avmmreaddata[3], w_hssi_pipe_gen1_2_avmmreaddata[2], w_hssi_pipe_gen1_2_avmmreaddata[1], w_hssi_pipe_gen1_2_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen3 = {w_hssi_pipe_gen3_avmmreaddata[7], w_hssi_pipe_gen3_avmmreaddata[6], w_hssi_pipe_gen3_avmmreaddata[5], w_hssi_pipe_gen3_avmmreaddata[4], w_hssi_pipe_gen3_avmmreaddata[3], w_hssi_pipe_gen3_avmmreaddata[2], w_hssi_pipe_gen3_avmmreaddata[1], w_hssi_pipe_gen3_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pcs_pma_interface = {w_hssi_rx_pcs_pma_interface_avmmreaddata[7], w_hssi_rx_pcs_pma_interface_avmmreaddata[6], w_hssi_rx_pcs_pma_interface_avmmreaddata[5], w_hssi_rx_pcs_pma_interface_avmmreaddata[4], w_hssi_rx_pcs_pma_interface_avmmreaddata[3], w_hssi_rx_pcs_pma_interface_avmmreaddata[2], w_hssi_rx_pcs_pma_interface_avmmreaddata[1], w_hssi_rx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pld_pcs_interface = {w_hssi_rx_pld_pcs_interface_avmmreaddata[7], w_hssi_rx_pld_pcs_interface_avmmreaddata[6], w_hssi_rx_pld_pcs_interface_avmmreaddata[5], w_hssi_rx_pld_pcs_interface_avmmreaddata[4], w_hssi_rx_pld_pcs_interface_avmmreaddata[3], w_hssi_rx_pld_pcs_interface_avmmreaddata[2], w_hssi_rx_pld_pcs_interface_avmmreaddata[1], w_hssi_rx_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pcs_pma_interface = {w_hssi_tx_pcs_pma_interface_avmmreaddata[7], w_hssi_tx_pcs_pma_interface_avmmreaddata[6], w_hssi_tx_pcs_pma_interface_avmmreaddata[5], w_hssi_tx_pcs_pma_interface_avmmreaddata[4], w_hssi_tx_pcs_pma_interface_avmmreaddata[3], w_hssi_tx_pcs_pma_interface_avmmreaddata[2], w_hssi_tx_pcs_pma_interface_avmmreaddata[1], w_hssi_tx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pld_pcs_interface = {w_hssi_tx_pld_pcs_interface_avmmreaddata[7], w_hssi_tx_pld_pcs_interface_avmmreaddata[6], w_hssi_tx_pld_pcs_interface_avmmreaddata[5], w_hssi_tx_pld_pcs_interface_avmmreaddata[4], w_hssi_tx_pld_pcs_interface_avmmreaddata[3], w_hssi_tx_pld_pcs_interface_avmmreaddata[2], w_hssi_tx_pld_pcs_interface_avmmreaddata[1], w_hssi_tx_pld_pcs_interface_avmmreaddata[0]};
		assign out_blockselect_hssi_10g_rx_pcs = w_hssi_10g_rx_pcs_blockselect;
		assign out_blockselect_hssi_10g_tx_pcs = w_hssi_10g_tx_pcs_blockselect;
		assign out_blockselect_hssi_8g_rx_pcs = w_hssi_8g_rx_pcs_blockselect;
		assign out_blockselect_hssi_8g_tx_pcs = w_hssi_8g_tx_pcs_blockselect;
		assign out_blockselect_hssi_common_pcs_pma_interface = w_hssi_common_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_common_pld_pcs_interface = w_hssi_common_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_fifo_rx_pcs = w_hssi_fifo_rx_pcs_blockselect;
		assign out_blockselect_hssi_fifo_tx_pcs = w_hssi_fifo_tx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_rx_pcs = w_hssi_gen3_rx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_tx_pcs = w_hssi_gen3_tx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_rx_pcs = w_hssi_krfec_rx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_tx_pcs = w_hssi_krfec_tx_pcs_blockselect;
		assign out_blockselect_hssi_pipe_gen1_2 = w_hssi_pipe_gen1_2_blockselect;
		assign out_blockselect_hssi_pipe_gen3 = w_hssi_pipe_gen3_blockselect;
		assign out_blockselect_hssi_rx_pcs_pma_interface = w_hssi_rx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_rx_pld_pcs_interface = w_hssi_rx_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_tx_pcs_pma_interface = w_hssi_tx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_tx_pld_pcs_interface = w_hssi_tx_pld_pcs_interface_blockselect;
		assign out_bond_pcs10g_out_bot = {w_hssi_10g_tx_pcs_distdwn_out_rden, w_hssi_10g_tx_pcs_distdwn_out_wren, w_hssi_10g_tx_pcs_distdwn_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs10g_out_top = {w_hssi_10g_tx_pcs_distup_out_rden, w_hssi_10g_tx_pcs_distup_out_wren, w_hssi_10g_tx_pcs_distup_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs8g_out_bot = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down, w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_down, w_hssi_8g_tx_pcs_wr_enable_out_chnl_down, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_down, w_hssi_8g_rx_pcs_wr_enable_out_chnl_down, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[0]};
		assign out_bond_pcs8g_out_top = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up, w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_up, w_hssi_8g_tx_pcs_wr_enable_out_chnl_up, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_up, w_hssi_8g_rx_pcs_wr_enable_out_chnl_up, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[0]};
		assign out_bond_pmaif_out_bot = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[0]};
		assign out_bond_pmaif_out_top = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[0]};
		assign out_hip_clk_out = {w_hssi_common_pld_pcs_interface_hip_cmn_clk[1], w_hssi_common_pld_pcs_interface_hip_cmn_clk[0], w_hssi_tx_pld_pcs_interface_hip_tx_clk};
		assign out_hip_ctrl_out = {w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[4], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[3], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[2], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[1], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[0], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[0]};
		assign out_hip_iocsr_rdy = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
		assign out_hip_iocsr_rdy_dly = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
		assign out_hip_nfrzdrv = w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
		assign out_hip_npor = w_hssi_common_pld_pcs_interface_hip_npor;
		assign out_hip_rx_data = {w_hssi_rx_pld_pcs_interface_hip_rx_data[50], w_hssi_rx_pld_pcs_interface_hip_rx_data[49], w_hssi_rx_pld_pcs_interface_hip_rx_data[48], w_hssi_rx_pld_pcs_interface_hip_rx_data[47], w_hssi_rx_pld_pcs_interface_hip_rx_data[46], w_hssi_rx_pld_pcs_interface_hip_rx_data[45], w_hssi_rx_pld_pcs_interface_hip_rx_data[44], w_hssi_rx_pld_pcs_interface_hip_rx_data[43], w_hssi_rx_pld_pcs_interface_hip_rx_data[42], w_hssi_rx_pld_pcs_interface_hip_rx_data[41], w_hssi_rx_pld_pcs_interface_hip_rx_data[40], w_hssi_rx_pld_pcs_interface_hip_rx_data[39], w_hssi_rx_pld_pcs_interface_hip_rx_data[38], w_hssi_rx_pld_pcs_interface_hip_rx_data[37], w_hssi_rx_pld_pcs_interface_hip_rx_data[36], w_hssi_rx_pld_pcs_interface_hip_rx_data[35], w_hssi_rx_pld_pcs_interface_hip_rx_data[34], w_hssi_rx_pld_pcs_interface_hip_rx_data[33], w_hssi_rx_pld_pcs_interface_hip_rx_data[32], w_hssi_rx_pld_pcs_interface_hip_rx_data[31], w_hssi_rx_pld_pcs_interface_hip_rx_data[30], w_hssi_rx_pld_pcs_interface_hip_rx_data[29], w_hssi_rx_pld_pcs_interface_hip_rx_data[28], w_hssi_rx_pld_pcs_interface_hip_rx_data[27], w_hssi_rx_pld_pcs_interface_hip_rx_data[26], w_hssi_rx_pld_pcs_interface_hip_rx_data[25], w_hssi_rx_pld_pcs_interface_hip_rx_data[24], w_hssi_rx_pld_pcs_interface_hip_rx_data[23], w_hssi_rx_pld_pcs_interface_hip_rx_data[22], w_hssi_rx_pld_pcs_interface_hip_rx_data[21], w_hssi_rx_pld_pcs_interface_hip_rx_data[20], w_hssi_rx_pld_pcs_interface_hip_rx_data[19], w_hssi_rx_pld_pcs_interface_hip_rx_data[18], w_hssi_rx_pld_pcs_interface_hip_rx_data[17], w_hssi_rx_pld_pcs_interface_hip_rx_data[16], w_hssi_rx_pld_pcs_interface_hip_rx_data[15], w_hssi_rx_pld_pcs_interface_hip_rx_data[14], w_hssi_rx_pld_pcs_interface_hip_rx_data[13], w_hssi_rx_pld_pcs_interface_hip_rx_data[12], w_hssi_rx_pld_pcs_interface_hip_rx_data[11], w_hssi_rx_pld_pcs_interface_hip_rx_data[10], w_hssi_rx_pld_pcs_interface_hip_rx_data[9], w_hssi_rx_pld_pcs_interface_hip_rx_data[8], w_hssi_rx_pld_pcs_interface_hip_rx_data[7], w_hssi_rx_pld_pcs_interface_hip_rx_data[6], w_hssi_rx_pld_pcs_interface_hip_rx_data[5], w_hssi_rx_pld_pcs_interface_hip_rx_data[4], w_hssi_rx_pld_pcs_interface_hip_rx_data[3], w_hssi_rx_pld_pcs_interface_hip_rx_data[2], w_hssi_rx_pld_pcs_interface_hip_rx_data[1], w_hssi_rx_pld_pcs_interface_hip_rx_data[0]};
		assign out_hip_usermode = w_hssi_common_pld_pcs_interface_hip_usermode;
		assign out_pld_10g_krfec_rx_blk_lock = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
		assign out_pld_10g_krfec_rx_diag_data_status = {w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1], w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[0]};
		assign out_pld_10g_krfec_rx_frame = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
		assign out_pld_10g_krfec_tx_frame = w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
		assign out_pld_10g_rx_align_val = w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
		assign out_pld_10g_rx_crc32_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
		assign out_pld_10g_rx_data_valid = w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
		assign out_pld_10g_rx_empty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
		assign out_pld_10g_rx_fifo_del = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
		assign out_pld_10g_rx_fifo_insert = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
		assign out_pld_10g_rx_fifo_num = {w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[3], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[2], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[1], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[0]};
		assign out_pld_10g_rx_frame_lock = w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
		assign out_pld_10g_rx_hi_ber = w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
		assign out_pld_10g_rx_oflw_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
		assign out_pld_10g_rx_pempty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
		assign out_pld_10g_rx_pfull = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
		assign out_pld_10g_tx_burst_en_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
		assign out_pld_10g_tx_empty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
		assign out_pld_10g_tx_fifo_num = {w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[2], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[1], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[0]};
		assign out_pld_10g_tx_full = w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
		assign out_pld_10g_tx_pempty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
		assign out_pld_10g_tx_pfull = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
		assign out_pld_10g_tx_wordslip_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
		assign out_pld_8g_a1a2_k1k2_flag = {w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[2], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[1], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[0]};
		assign out_pld_8g_empty_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
		assign out_pld_8g_empty_rx = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
		assign out_pld_8g_empty_tx = w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
		assign out_pld_8g_full_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
		assign out_pld_8g_full_rx = w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
		assign out_pld_8g_full_tx = w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
		assign out_pld_8g_rxelecidle = w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
		assign out_pld_8g_signal_detect_out = w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
		assign out_pld_8g_wa_boundary = {w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0]};
		assign out_pld_krfec_tx_alignment = w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
		assign out_pld_pcs_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
		assign out_pld_pcs_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
		assign out_pld_pma_adapt_done = w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
		assign out_pld_pma_clkdiv_rx_user = w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
		assign out_pld_pma_clkdiv_tx_user = w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
		assign out_pld_pma_clklow = w_hssi_common_pld_pcs_interface_pld_pma_clklow;
		assign out_pld_pma_fref = w_hssi_common_pld_pcs_interface_pld_pma_fref;
		assign out_pld_pma_hclk = w_hssi_common_pld_pcs_interface_pld_pma_hclk;
		assign out_pld_pma_pcie_sw_done = {w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1], w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[0]};
		assign out_pld_pma_pfdmode_lock = w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
		assign out_pld_pma_reserved_in = {w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[3], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[2], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[1], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[0]};
		assign out_pld_pma_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
		assign out_pld_pma_rx_detect_valid = w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
		assign out_pld_pma_rx_found = w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
		assign out_pld_pma_rxpll_lock = w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
		assign out_pld_pma_signal_ok = w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
		assign out_pld_pma_testbus = {w_hssi_common_pld_pcs_interface_pld_pma_testbus[7], w_hssi_common_pld_pcs_interface_pld_pma_testbus[6], w_hssi_common_pld_pcs_interface_pld_pma_testbus[5], w_hssi_common_pld_pcs_interface_pld_pma_testbus[4], w_hssi_common_pld_pcs_interface_pld_pma_testbus[3], w_hssi_common_pld_pcs_interface_pld_pma_testbus[2], w_hssi_common_pld_pcs_interface_pld_pma_testbus[1], w_hssi_common_pld_pcs_interface_pld_pma_testbus[0]};
		assign out_pld_pma_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
		assign out_pld_pmaif_mask_tx_pll = w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
		assign out_pld_reserved_out = {w_hssi_common_pld_pcs_interface_pld_reserved_out[9], w_hssi_common_pld_pcs_interface_pld_reserved_out[8], w_hssi_common_pld_pcs_interface_pld_reserved_out[7], w_hssi_common_pld_pcs_interface_pld_reserved_out[6], w_hssi_common_pld_pcs_interface_pld_reserved_out[5], w_hssi_common_pld_pcs_interface_pld_reserved_out[4], w_hssi_common_pld_pcs_interface_pld_reserved_out[3], w_hssi_common_pld_pcs_interface_pld_reserved_out[2], w_hssi_common_pld_pcs_interface_pld_reserved_out[1], w_hssi_common_pld_pcs_interface_pld_reserved_out[0]};
		assign out_pld_rx_control = {w_hssi_rx_pld_pcs_interface_pld_rx_control[19], w_hssi_rx_pld_pcs_interface_pld_rx_control[18], w_hssi_rx_pld_pcs_interface_pld_rx_control[17], w_hssi_rx_pld_pcs_interface_pld_rx_control[16], w_hssi_rx_pld_pcs_interface_pld_rx_control[15], w_hssi_rx_pld_pcs_interface_pld_rx_control[14], w_hssi_rx_pld_pcs_interface_pld_rx_control[13], w_hssi_rx_pld_pcs_interface_pld_rx_control[12], w_hssi_rx_pld_pcs_interface_pld_rx_control[11], w_hssi_rx_pld_pcs_interface_pld_rx_control[10], w_hssi_rx_pld_pcs_interface_pld_rx_control[9], w_hssi_rx_pld_pcs_interface_pld_rx_control[8], w_hssi_rx_pld_pcs_interface_pld_rx_control[7], w_hssi_rx_pld_pcs_interface_pld_rx_control[6], w_hssi_rx_pld_pcs_interface_pld_rx_control[5], w_hssi_rx_pld_pcs_interface_pld_rx_control[4], w_hssi_rx_pld_pcs_interface_pld_rx_control[3], w_hssi_rx_pld_pcs_interface_pld_rx_control[2], w_hssi_rx_pld_pcs_interface_pld_rx_control[1], w_hssi_rx_pld_pcs_interface_pld_rx_control[0]};
		assign out_pld_rx_data = {w_hssi_rx_pld_pcs_interface_pld_rx_data[127], w_hssi_rx_pld_pcs_interface_pld_rx_data[126], w_hssi_rx_pld_pcs_interface_pld_rx_data[125], w_hssi_rx_pld_pcs_interface_pld_rx_data[124], w_hssi_rx_pld_pcs_interface_pld_rx_data[123], w_hssi_rx_pld_pcs_interface_pld_rx_data[122], w_hssi_rx_pld_pcs_interface_pld_rx_data[121], w_hssi_rx_pld_pcs_interface_pld_rx_data[120], w_hssi_rx_pld_pcs_interface_pld_rx_data[119], w_hssi_rx_pld_pcs_interface_pld_rx_data[118], w_hssi_rx_pld_pcs_interface_pld_rx_data[117], w_hssi_rx_pld_pcs_interface_pld_rx_data[116], w_hssi_rx_pld_pcs_interface_pld_rx_data[115], w_hssi_rx_pld_pcs_interface_pld_rx_data[114], w_hssi_rx_pld_pcs_interface_pld_rx_data[113], w_hssi_rx_pld_pcs_interface_pld_rx_data[112], w_hssi_rx_pld_pcs_interface_pld_rx_data[111], w_hssi_rx_pld_pcs_interface_pld_rx_data[110], w_hssi_rx_pld_pcs_interface_pld_rx_data[109], w_hssi_rx_pld_pcs_interface_pld_rx_data[108], w_hssi_rx_pld_pcs_interface_pld_rx_data[107], w_hssi_rx_pld_pcs_interface_pld_rx_data[106], w_hssi_rx_pld_pcs_interface_pld_rx_data[105], w_hssi_rx_pld_pcs_interface_pld_rx_data[104], w_hssi_rx_pld_pcs_interface_pld_rx_data[103], w_hssi_rx_pld_pcs_interface_pld_rx_data[102], w_hssi_rx_pld_pcs_interface_pld_rx_data[101], w_hssi_rx_pld_pcs_interface_pld_rx_data[100], w_hssi_rx_pld_pcs_interface_pld_rx_data[99], w_hssi_rx_pld_pcs_interface_pld_rx_data[98], w_hssi_rx_pld_pcs_interface_pld_rx_data[97], w_hssi_rx_pld_pcs_interface_pld_rx_data[96], w_hssi_rx_pld_pcs_interface_pld_rx_data[95], w_hssi_rx_pld_pcs_interface_pld_rx_data[94], w_hssi_rx_pld_pcs_interface_pld_rx_data[93], w_hssi_rx_pld_pcs_interface_pld_rx_data[92], w_hssi_rx_pld_pcs_interface_pld_rx_data[91], w_hssi_rx_pld_pcs_interface_pld_rx_data[90], w_hssi_rx_pld_pcs_interface_pld_rx_data[89], w_hssi_rx_pld_pcs_interface_pld_rx_data[88], w_hssi_rx_pld_pcs_interface_pld_rx_data[87], w_hssi_rx_pld_pcs_interface_pld_rx_data[86], w_hssi_rx_pld_pcs_interface_pld_rx_data[85], w_hssi_rx_pld_pcs_interface_pld_rx_data[84], w_hssi_rx_pld_pcs_interface_pld_rx_data[83], w_hssi_rx_pld_pcs_interface_pld_rx_data[82], w_hssi_rx_pld_pcs_interface_pld_rx_data[81], w_hssi_rx_pld_pcs_interface_pld_rx_data[80], w_hssi_rx_pld_pcs_interface_pld_rx_data[79], w_hssi_rx_pld_pcs_interface_pld_rx_data[78], w_hssi_rx_pld_pcs_interface_pld_rx_data[77], w_hssi_rx_pld_pcs_interface_pld_rx_data[76], w_hssi_rx_pld_pcs_interface_pld_rx_data[75], w_hssi_rx_pld_pcs_interface_pld_rx_data[74], w_hssi_rx_pld_pcs_interface_pld_rx_data[73], w_hssi_rx_pld_pcs_interface_pld_rx_data[72], w_hssi_rx_pld_pcs_interface_pld_rx_data[71], w_hssi_rx_pld_pcs_interface_pld_rx_data[70], w_hssi_rx_pld_pcs_interface_pld_rx_data[69], w_hssi_rx_pld_pcs_interface_pld_rx_data[68], w_hssi_rx_pld_pcs_interface_pld_rx_data[67], w_hssi_rx_pld_pcs_interface_pld_rx_data[66], w_hssi_rx_pld_pcs_interface_pld_rx_data[65], w_hssi_rx_pld_pcs_interface_pld_rx_data[64], w_hssi_rx_pld_pcs_interface_pld_rx_data[63], w_hssi_rx_pld_pcs_interface_pld_rx_data[62], w_hssi_rx_pld_pcs_interface_pld_rx_data[61], w_hssi_rx_pld_pcs_interface_pld_rx_data[60], w_hssi_rx_pld_pcs_interface_pld_rx_data[59], w_hssi_rx_pld_pcs_interface_pld_rx_data[58], w_hssi_rx_pld_pcs_interface_pld_rx_data[57], w_hssi_rx_pld_pcs_interface_pld_rx_data[56], w_hssi_rx_pld_pcs_interface_pld_rx_data[55], w_hssi_rx_pld_pcs_interface_pld_rx_data[54], w_hssi_rx_pld_pcs_interface_pld_rx_data[53], w_hssi_rx_pld_pcs_interface_pld_rx_data[52], w_hssi_rx_pld_pcs_interface_pld_rx_data[51], w_hssi_rx_pld_pcs_interface_pld_rx_data[50], w_hssi_rx_pld_pcs_interface_pld_rx_data[49], w_hssi_rx_pld_pcs_interface_pld_rx_data[48], w_hssi_rx_pld_pcs_interface_pld_rx_data[47], w_hssi_rx_pld_pcs_interface_pld_rx_data[46], w_hssi_rx_pld_pcs_interface_pld_rx_data[45], w_hssi_rx_pld_pcs_interface_pld_rx_data[44], w_hssi_rx_pld_pcs_interface_pld_rx_data[43], w_hssi_rx_pld_pcs_interface_pld_rx_data[42], w_hssi_rx_pld_pcs_interface_pld_rx_data[41], w_hssi_rx_pld_pcs_interface_pld_rx_data[40], w_hssi_rx_pld_pcs_interface_pld_rx_data[39], w_hssi_rx_pld_pcs_interface_pld_rx_data[38], w_hssi_rx_pld_pcs_interface_pld_rx_data[37], w_hssi_rx_pld_pcs_interface_pld_rx_data[36], w_hssi_rx_pld_pcs_interface_pld_rx_data[35], w_hssi_rx_pld_pcs_interface_pld_rx_data[34], w_hssi_rx_pld_pcs_interface_pld_rx_data[33], w_hssi_rx_pld_pcs_interface_pld_rx_data[32], w_hssi_rx_pld_pcs_interface_pld_rx_data[31], w_hssi_rx_pld_pcs_interface_pld_rx_data[30], w_hssi_rx_pld_pcs_interface_pld_rx_data[29], w_hssi_rx_pld_pcs_interface_pld_rx_data[28], w_hssi_rx_pld_pcs_interface_pld_rx_data[27], w_hssi_rx_pld_pcs_interface_pld_rx_data[26], w_hssi_rx_pld_pcs_interface_pld_rx_data[25], w_hssi_rx_pld_pcs_interface_pld_rx_data[24], w_hssi_rx_pld_pcs_interface_pld_rx_data[23], w_hssi_rx_pld_pcs_interface_pld_rx_data[22], w_hssi_rx_pld_pcs_interface_pld_rx_data[21], w_hssi_rx_pld_pcs_interface_pld_rx_data[20], w_hssi_rx_pld_pcs_interface_pld_rx_data[19], w_hssi_rx_pld_pcs_interface_pld_rx_data[18], w_hssi_rx_pld_pcs_interface_pld_rx_data[17], w_hssi_rx_pld_pcs_interface_pld_rx_data[16], w_hssi_rx_pld_pcs_interface_pld_rx_data[15], w_hssi_rx_pld_pcs_interface_pld_rx_data[14], w_hssi_rx_pld_pcs_interface_pld_rx_data[13], w_hssi_rx_pld_pcs_interface_pld_rx_data[12], w_hssi_rx_pld_pcs_interface_pld_rx_data[11], w_hssi_rx_pld_pcs_interface_pld_rx_data[10], w_hssi_rx_pld_pcs_interface_pld_rx_data[9], w_hssi_rx_pld_pcs_interface_pld_rx_data[8], w_hssi_rx_pld_pcs_interface_pld_rx_data[7], w_hssi_rx_pld_pcs_interface_pld_rx_data[6], w_hssi_rx_pld_pcs_interface_pld_rx_data[5], w_hssi_rx_pld_pcs_interface_pld_rx_data[4], w_hssi_rx_pld_pcs_interface_pld_rx_data[3], w_hssi_rx_pld_pcs_interface_pld_rx_data[2], w_hssi_rx_pld_pcs_interface_pld_rx_data[1], w_hssi_rx_pld_pcs_interface_pld_rx_data[0]};
		assign out_pld_rx_prbs_done = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
		assign out_pld_rx_prbs_err = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
		assign out_pld_test_data = {w_hssi_common_pld_pcs_interface_pld_test_data[19], w_hssi_common_pld_pcs_interface_pld_test_data[18], w_hssi_common_pld_pcs_interface_pld_test_data[17], w_hssi_common_pld_pcs_interface_pld_test_data[16], w_hssi_common_pld_pcs_interface_pld_test_data[15], w_hssi_common_pld_pcs_interface_pld_test_data[14], w_hssi_common_pld_pcs_interface_pld_test_data[13], w_hssi_common_pld_pcs_interface_pld_test_data[12], w_hssi_common_pld_pcs_interface_pld_test_data[11], w_hssi_common_pld_pcs_interface_pld_test_data[10], w_hssi_common_pld_pcs_interface_pld_test_data[9], w_hssi_common_pld_pcs_interface_pld_test_data[8], w_hssi_common_pld_pcs_interface_pld_test_data[7], w_hssi_common_pld_pcs_interface_pld_test_data[6], w_hssi_common_pld_pcs_interface_pld_test_data[5], w_hssi_common_pld_pcs_interface_pld_test_data[4], w_hssi_common_pld_pcs_interface_pld_test_data[3], w_hssi_common_pld_pcs_interface_pld_test_data[2], w_hssi_common_pld_pcs_interface_pld_test_data[1], w_hssi_common_pld_pcs_interface_pld_test_data[0]};
		assign out_pld_uhsif_lock = w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
		assign out_pld_uhsif_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
		assign out_pma_adapt_start = w_hssi_common_pcs_pma_interface_pma_adapt_start;
		assign out_pma_atpg_los_en_n = w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
		assign out_pma_csr_test_dis = w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
		assign out_pma_current_coeff = {w_hssi_common_pcs_pma_interface_pma_current_coeff[17], w_hssi_common_pcs_pma_interface_pma_current_coeff[16], w_hssi_common_pcs_pma_interface_pma_current_coeff[15], w_hssi_common_pcs_pma_interface_pma_current_coeff[14], w_hssi_common_pcs_pma_interface_pma_current_coeff[13], w_hssi_common_pcs_pma_interface_pma_current_coeff[12], w_hssi_common_pcs_pma_interface_pma_current_coeff[11], w_hssi_common_pcs_pma_interface_pma_current_coeff[10], w_hssi_common_pcs_pma_interface_pma_current_coeff[9], w_hssi_common_pcs_pma_interface_pma_current_coeff[8], w_hssi_common_pcs_pma_interface_pma_current_coeff[7], w_hssi_common_pcs_pma_interface_pma_current_coeff[6], w_hssi_common_pcs_pma_interface_pma_current_coeff[5], w_hssi_common_pcs_pma_interface_pma_current_coeff[4], w_hssi_common_pcs_pma_interface_pma_current_coeff[3], w_hssi_common_pcs_pma_interface_pma_current_coeff[2], w_hssi_common_pcs_pma_interface_pma_current_coeff[1], w_hssi_common_pcs_pma_interface_pma_current_coeff[0]};
		assign out_pma_current_rxpreset = {w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[1], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[0]};
		assign out_pma_early_eios = w_hssi_common_pcs_pma_interface_pma_early_eios;
		assign out_pma_eye_monitor = {w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0]};
		assign out_pma_interface_select = {w_hssi_common_pcs_pma_interface_pma_interface_select[1], w_hssi_common_pcs_pma_interface_pma_interface_select[0]};
		assign out_pma_ltd_b = w_hssi_common_pcs_pma_interface_pma_ltd_b;
		assign out_pma_ltr = w_hssi_common_pcs_pma_interface_pma_ltr;
		assign out_pma_nfrzdrv = w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
		assign out_pma_nrpi_freeze = w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
		assign out_pma_pcie_switch = {w_hssi_common_pcs_pma_interface_pma_pcie_switch[1], w_hssi_common_pcs_pma_interface_pma_pcie_switch[0]};
		assign out_pma_ppm_lock = w_hssi_common_pcs_pma_interface_pma_ppm_lock;
		assign out_pma_reserved_out = {w_hssi_common_pcs_pma_interface_pma_reserved_out[4], w_hssi_common_pcs_pma_interface_pma_reserved_out[3], w_hssi_common_pcs_pma_interface_pma_reserved_out[2], w_hssi_common_pcs_pma_interface_pma_reserved_out[1], w_hssi_common_pcs_pma_interface_pma_reserved_out[0]};
		assign out_pma_rs_lpbk_b = w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
		assign out_pma_rx_clkslip = w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
		assign out_pma_rx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
		assign out_pma_rxpma_rstb = w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
		assign out_pma_scan_mode_n = w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
		assign out_pma_scan_shift_n = w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
		assign out_pma_tx_bitslip = w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
		assign out_pma_tx_bonding_rstb = w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
		assign out_pma_tx_elec_idle = w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
		assign out_pma_tx_pma_data = {w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0]};
		assign out_pma_tx_qpi_pulldn = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
		assign out_pma_tx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
		assign out_pma_tx_txdetectrx = w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
		assign out_pma_txpma_rstb = w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	endgenerate
endmodule
module twentynm_pcs_rev_20nm5
	#(
	//PARAM_LIST_START
		parameter xcvr_native_mode = "mode_duplex",  // mode_duplex, mode_rx_only, mode_tx_only
		
		// parameters for twentynm_hssi_10g_rx_pcs
		parameter hssi_10g_rx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_align_del = "align_del_en", // align_del_dis|align_del_en
		parameter hssi_10g_rx_pcs_ber_bit_err_total_cnt = "bit_err_total_cnt_10g", // bit_err_total_cnt_10g
		parameter hssi_10g_rx_pcs_ber_clken = "ber_clk_dis", // ber_clk_dis|ber_clk_en
		parameter hssi_10g_rx_pcs_ber_xus_timer_window = 21'b100110001001010,
		parameter hssi_10g_rx_pcs_bitslip_mode = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_rx_pcs_blksync_bitslip_type = "bitslip_comb", // bitslip_comb|bitslip_reg
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_cnt = 3'b1,
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_type = "bitslip_match", // bitslip_match|bitslip_cnt
		parameter hssi_10g_rx_pcs_blksync_bypass = "blksync_bypass_dis", // blksync_bypass_dis|blksync_bypass_en
		parameter hssi_10g_rx_pcs_blksync_clken = "blksync_clk_dis", // blksync_clk_dis|blksync_clk_en
		parameter hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt = "enum_invalid_sh_cnt_10g", // enum_invalid_sh_cnt_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock = "knum_sh_cnt_postlock_10g", // knum_sh_cnt_postlock_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock = "knum_sh_cnt_prelock_10g", // knum_sh_cnt_prelock_10g
		parameter hssi_10g_rx_pcs_blksync_pipeln = "blksync_pipeln_dis", // blksync_pipeln_dis|blksync_pipeln_en
		parameter hssi_10g_rx_pcs_clr_errblk_cnt_en = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_control_del = "control_del_all", // control_del_all|control_del_none
		parameter hssi_10g_rx_pcs_crcchk_bypass = "crcchk_bypass_dis", // crcchk_bypass_dis|crcchk_bypass_en
		parameter hssi_10g_rx_pcs_crcchk_clken = "crcchk_clk_dis", // crcchk_clk_dis|crcchk_clk_en
		parameter hssi_10g_rx_pcs_crcchk_inv = "crcchk_inv_dis", // crcchk_inv_dis|crcchk_inv_en
		parameter hssi_10g_rx_pcs_crcchk_pipeln = "crcchk_pipeln_dis", // crcchk_pipeln_dis|crcchk_pipeln_en
		parameter hssi_10g_rx_pcs_crcflag_pipeln = "crcflag_pipeln_dis", // crcflag_pipeln_dis|crcflag_pipeln_en
		parameter hssi_10g_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_rx_pcs_dec64b66b_clken = "dec64b66b_clk_dis", // dec64b66b_clk_dis|dec64b66b_clk_en
		parameter hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass = "dec_64b66b_rxsm_bypass_dis", // dec_64b66b_rxsm_bypass_dis|dec_64b66b_rxsm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_bypass = "descrm_bypass_en", // descrm_bypass_dis|descrm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_clken = "descrm_clk_dis", // descrm_clk_dis|descrm_clk_en
		parameter hssi_10g_rx_pcs_descrm_mode = "async", // async|sync
		parameter hssi_10g_rx_pcs_descrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_dft_clk_out_sel = "rx_master_clk", // rx_master_clk|rx_gbexp_clk|rx_blksync_clk|rx_descrm_clk|rx_frmsync_clk|rx_64b66bdec_clk|rx_ber_clk|rx_rand_clk|rx_crcchk_clk|rx_wrfifo_clk|rx_rdfifo_clk|rx_fec_clk
		parameter hssi_10g_rx_pcs_dis_signal_ok = "dis_signal_ok_dis", // dis_signal_ok_dis|dis_signal_ok_en
		parameter hssi_10g_rx_pcs_dispchk_bypass = "dispchk_bypass_dis", // dispchk_bypass_dis|dispchk_bypass_en
		parameter hssi_10g_rx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_rx_pcs_fast_path = "fast_path_dis", // fast_path_dis|fast_path_en
		parameter hssi_10g_rx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_rx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_rx_pcs_fifo_double_read = "fifo_double_read_dis", // fifo_double_read_dis|fifo_double_read_en
		parameter hssi_10g_rx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_rx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_rx_pcs_force_align = "force_align_dis", // force_align_dis|force_align_en
		parameter hssi_10g_rx_pcs_frmsync_bypass = "frmsync_bypass_dis", // frmsync_bypass_dis|frmsync_bypass_en
		parameter hssi_10g_rx_pcs_frmsync_clken = "frmsync_clk_dis", // frmsync_clk_dis|frmsync_clk_en
		parameter hssi_10g_rx_pcs_frmsync_enum_scrm = "enum_scrm_default", // enum_scrm_default
		parameter hssi_10g_rx_pcs_frmsync_enum_sync = "enum_sync_default", // enum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_flag_type = "all_framing_words", // all_framing_words|location_only
		parameter hssi_10g_rx_pcs_frmsync_knum_sync = "knum_sync_default", // knum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_mfrm_length = 16'b100000000000,
		parameter hssi_10g_rx_pcs_frmsync_pipeln = "frmsync_pipeln_dis", // frmsync_pipeln_dis|frmsync_pipeln_en
		parameter hssi_10g_rx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_rx_pcs_gb_rx_idwidth = "width_32", // width_40|width_32|width_64
		parameter hssi_10g_rx_pcs_gb_rx_odwidth = "width_66", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_rx_pcs_gbexp_clken = "gbexp_clk_dis", // gbexp_clk_dis|gbexp_clk_en
		parameter hssi_10g_rx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_10g_rx_pcs_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_rx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_rx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_rx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_rx_pcs_pld_if_type = "fifo", // fifo|reg
		parameter hssi_10g_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_rx_pcs_rand_clken = "rand_clk_dis", // rand_clk_dis|rand_clk_en
		parameter hssi_10g_rx_pcs_rd_clk_sel = "rd_rx_pma_clk", // rd_rx_pld_clk|rd_rx_pma_clk|rd_refclk_dig
		parameter hssi_10g_rx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_rx_pcs_rx_fifo_write_ctrl = "blklock_stops", // blklock_stops|blklock_ignore
		parameter hssi_10g_rx_pcs_rx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_rx_pcs_rx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_rx_pcs_rx_signal_ok_sel = "synchronized_ver", // synchronized_ver|nonsync_ver
		parameter hssi_10g_rx_pcs_rx_sm_bypass = "rx_sm_bypass_dis", // rx_sm_bypass_dis|rx_sm_bypass_en
		parameter hssi_10g_rx_pcs_rx_sm_hiber = "rx_sm_hiber_en", // rx_sm_hiber_en|rx_sm_hiber_dis
		parameter hssi_10g_rx_pcs_rx_sm_pipeln = "rx_sm_pipeln_dis", // rx_sm_pipeln_dis|rx_sm_pipeln_en
		parameter hssi_10g_rx_pcs_rx_testbus_sel = "crc32_chk_testbus1", // crc32_chk_testbus1|crc32_chk_testbus2|frame_sync_testbus1|frame_sync_testbus2|dec64b66b_testbus|rxsm_testbus|ber_testbus|blksync_testbus1|blksync_testbus2|gearbox_exp_testbus|random_ver_testbus|descramble_testbus|blank_testbus|rx_fifo_testbus1|rx_fifo_testbus2
		parameter hssi_10g_rx_pcs_rx_true_b2b = "b2b", // single|b2b
		parameter hssi_10g_rx_pcs_rxfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_rx_pcs_rxfifo_full = "full_default", // full_default
		parameter hssi_10g_rx_pcs_rxfifo_mode = "phase_comp", // register_mode|clk_comp_10g|generic_interlaken|generic_basic|phase_comp|phase_comp_dv
		parameter hssi_10g_rx_pcs_rxfifo_pempty = 5'b10,
		parameter hssi_10g_rx_pcs_rxfifo_pfull = 5'b10111,
		parameter hssi_10g_rx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_rx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_rx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_10g_tx_pcs
		parameter hssi_10g_tx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_bitslip_en = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_10g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_10g_tx_pcs_comp_cnt = 8'b0,
		parameter hssi_10g_tx_pcs_compin_sel = "compin_master", // compin_master|compin_slave_top|compin_slave_bot|compin_default
		parameter hssi_10g_tx_pcs_crcgen_bypass = "crcgen_bypass_dis", // crcgen_bypass_dis|crcgen_bypass_en
		parameter hssi_10g_tx_pcs_crcgen_clken = "crcgen_clk_dis", // crcgen_clk_dis|crcgen_clk_en
		parameter hssi_10g_tx_pcs_crcgen_err = "crcgen_err_dis", // crcgen_err_dis|crcgen_err_en
		parameter hssi_10g_tx_pcs_crcgen_inv = "crcgen_inv_dis", // crcgen_inv_dis|crcgen_inv_en
		parameter hssi_10g_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_tx_pcs_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_10g_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_tx_pcs_dft_clk_out_sel = "tx_master_clk", // tx_master_clk|tx_rdfifo_clk|tx_frmgen_clk|tx_crcgen_clk|tx_64b66benc_txsm_clk|tx_scrm_clk|tx_dispgen_clk|tx_gbred_clk|tx_wrfifo_clk|tx_fec_clk
		parameter hssi_10g_tx_pcs_dispgen_bypass = "dispgen_bypass_dis", // dispgen_bypass_dis|dispgen_bypass_en
		parameter hssi_10g_tx_pcs_dispgen_clken = "dispgen_clk_dis", // dispgen_clk_dis|dispgen_clk_en
		parameter hssi_10g_tx_pcs_dispgen_err = "dispgen_err_dis", // dispgen_err_dis|dispgen_err_en
		parameter hssi_10g_tx_pcs_dispgen_pipeln = "dispgen_pipeln_dis", // dispgen_pipeln_dis|dispgen_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_bypass_pipeln = "distdwn_bypass_pipeln_dis", // distdwn_bypass_pipeln_dis|distdwn_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_master = "distdwn_master_en", // distdwn_master_en|distdwn_master_dis
		parameter hssi_10g_tx_pcs_distup_bypass_pipeln = "distup_bypass_pipeln_dis", // distup_bypass_pipeln_dis|distup_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distup_master = "distup_master_en", // distup_master_en|distup_master_dis
		parameter hssi_10g_tx_pcs_dv_bond = "dv_bond_dis", // dv_bond_en|dv_bond_dis
		parameter hssi_10g_tx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_tx_pcs_enc64b66b_txsm_clken = "enc64b66b_txsm_clk_dis", // enc64b66b_txsm_clk_dis|enc64b66b_txsm_clk_en
		parameter hssi_10g_tx_pcs_enc_64b66b_txsm_bypass = "enc_64b66b_txsm_bypass_dis", // enc_64b66b_txsm_bypass_dis|enc_64b66b_txsm_bypass_en
		parameter hssi_10g_tx_pcs_fastpath = "fastpath_dis", // fastpath_dis|fastpath_en
		parameter hssi_10g_tx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_tx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_tx_pcs_fifo_double_write = "fifo_double_write_dis", // fifo_double_write_dis|fifo_double_write_en
		parameter hssi_10g_tx_pcs_fifo_reg_fast = "fifo_reg_fast_dis", // fifo_reg_fast_dis|fifo_reg_fast_en
		parameter hssi_10g_tx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_tx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_tx_pcs_frmgen_burst = "frmgen_burst_dis", // frmgen_burst_dis|frmgen_burst_en
		parameter hssi_10g_tx_pcs_frmgen_bypass = "frmgen_bypass_dis", // frmgen_bypass_dis|frmgen_bypass_en
		parameter hssi_10g_tx_pcs_frmgen_clken = "frmgen_clk_dis", // frmgen_clk_dis|frmgen_clk_en
		parameter hssi_10g_tx_pcs_frmgen_mfrm_length = 16'b100000000000,
		parameter hssi_10g_tx_pcs_frmgen_pipeln = "frmgen_pipeln_dis", // frmgen_pipeln_dis|frmgen_pipeln_en
		parameter hssi_10g_tx_pcs_frmgen_pyld_ins = "frmgen_pyld_ins_dis", // frmgen_pyld_ins_dis|frmgen_pyld_ins_en
		parameter hssi_10g_tx_pcs_frmgen_wordslip = "frmgen_wordslip_dis", // frmgen_wordslip_dis|frmgen_wordslip_en
		parameter hssi_10g_tx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_tx_pcs_gb_pipeln_bypass = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_gb_tx_idwidth = "width_50", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_tx_pcs_gb_tx_odwidth = "width_32", // width_32|width_40|width_64
		parameter hssi_10g_tx_pcs_gbred_clken = "gbred_clk_dis", // gbred_clk_dis|gbred_clk_en
		parameter hssi_10g_tx_pcs_indv = "indv_en", // indv_en|indv_dis
		parameter hssi_10g_tx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_tx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_tx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_tx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del6|phcomp_rd_del5|phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_tx_pcs_pld_if_type = "fifo", // fifo|reg|fastreg
		parameter hssi_10g_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_tx_pcs_pseudo_random = "all_0", // two_lf|all_0
		parameter hssi_10g_tx_pcs_pseudo_seed_a = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_pseudo_seed_b = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_random_disp = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_tx_pcs_scrm_bypass = "scrm_bypass_dis", // scrm_bypass_dis|scrm_bypass_en
		parameter hssi_10g_tx_pcs_scrm_clken = "scrm_clk_dis", // scrm_clk_dis|scrm_clk_en
		parameter hssi_10g_tx_pcs_scrm_mode = "async", // async|sync
		parameter hssi_10g_tx_pcs_scrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_sh_err = "sh_err_dis", // sh_err_dis|sh_err_en
		parameter hssi_10g_tx_pcs_sop_mark = "sop_mark_dis", // sop_mark_en|sop_mark_dis
		parameter hssi_10g_tx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_tx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_tx_pcs_tx_scrm_err = "scrm_err_dis", // scrm_err_dis|scrm_err_en
		parameter hssi_10g_tx_pcs_tx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_tx_pcs_tx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_tx_pcs_tx_sm_bypass = "tx_sm_bypass_dis", // tx_sm_bypass_dis|tx_sm_bypass_en
		parameter hssi_10g_tx_pcs_tx_sm_pipeln = "tx_sm_pipeln_dis", // tx_sm_pipeln_dis|tx_sm_pipeln_en
		parameter hssi_10g_tx_pcs_tx_testbus_sel = "crc32_gen_testbus1", // crc32_gen_testbus1|crc32_gen_testbus2|disp_gen_testbus1|disp_gen_testbus2|frame_gen_testbus1|frame_gen_testbus2|enc64b66b_testbus|txsm_testbus|tx_cp_bond_testbus|gearbox_red_testbus|scramble_testbus|blank_testbus|tx_fifo_testbus1|tx_fifo_testbus2
		parameter hssi_10g_tx_pcs_txfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_tx_pcs_txfifo_full = "full_default", // full_default
		parameter hssi_10g_tx_pcs_txfifo_mode = "phase_comp", // register_mode|interlaken_generic|basic_generic|phase_comp
		parameter hssi_10g_tx_pcs_txfifo_pempty = 4'b10,
		parameter hssi_10g_tx_pcs_txfifo_pfull = 4'b1011,
		parameter hssi_10g_tx_pcs_wr_clk_sel = "wr_tx_pma_clk", // wr_tx_pld_clk|wr_tx_pma_clk|wr_refclk_dig
		parameter hssi_10g_tx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_8g_rx_pcs
		parameter hssi_8g_rx_pcs_auto_error_replacement = "dis_err_replace", // dis_err_replace|en_err_replace
		parameter hssi_8g_rx_pcs_auto_speed_nego = "dis_asn", // dis_asn|en_asn_g2_freq_scal
		parameter hssi_8g_rx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_rx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_rx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_rx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_rx_pcs_byte_deserializer = "dis_bds", // dis_bds|en_bds_by_2|en_bds_by_4|en_bds_by_2_det
		parameter hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask = "dis_rxvalid_mask", // dis_rxvalid_mask|en_rxvalid_mask
		parameter hssi_8g_rx_pcs_clkcmp_pattern_n = 20'b0,
		parameter hssi_8g_rx_pcs_clkcmp_pattern_p = 20'b0,
		parameter hssi_8g_rx_pcs_clock_gate_bds_dec_asn = "dis_bds_dec_asn_clk_gating", // dis_bds_dec_asn_clk_gating|en_bds_dec_asn_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_cdr_eidle = "dis_cdr_eidle_clk_gating", // dis_cdr_eidle_clk_gating|en_cdr_eidle_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk = "dis_dw_pc_wrclk_gating", // dis_dw_pc_wrclk_gating|en_dw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_rd = "dis_dw_rm_rdclk_gating", // dis_dw_rm_rdclk_gating|en_dw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_wr = "dis_dw_rm_wrclk_gating", // dis_dw_rm_wrclk_gating|en_dw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_wa = "dis_dw_wa_clk_gating", // dis_dw_wa_clk_gating|en_dw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_pc_rdclk = "dis_pc_rdclk_gating", // dis_pc_rdclk_gating|en_pc_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk = "dis_sw_pc_wrclk_gating", // dis_sw_pc_wrclk_gating|en_sw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_rd = "dis_sw_rm_rdclk_gating", // dis_sw_rm_rdclk_gating|en_sw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_wr = "dis_sw_rm_wrclk_gating", // dis_sw_rm_wrclk_gating|en_sw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_wa = "dis_sw_wa_clk_gating", // dis_sw_wa_clk_gating|en_sw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_observation_in_pld_core = "internal_sw_wa_clk", // internal_sw_wa_clk|internal_dw_wa_clk|internal_cdr_eidle_clk|internal_sm_rm_wr_clk|internal_dw_rm_wr_clk|internal_clk_2_b|internal_sw_rm_rd_clk|internal_dw_rm_rd_clk|internal_sw_rx_wr_clk|internal_dw_rx_wr_clk|internal_rx_rd_clk|internal_rx_pma_clk_gen3|internal_rx_rcvd_clk_gen3
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_rx_pcs_eidle_entry_eios = "dis_eidle_eios", // dis_eidle_eios|en_eidle_eios
		parameter hssi_8g_rx_pcs_eidle_entry_iei = "dis_eidle_iei", // dis_eidle_iei|en_eidle_iei
		parameter hssi_8g_rx_pcs_eidle_entry_sd = "dis_eidle_sd", // dis_eidle_sd|en_eidle_sd
		parameter hssi_8g_rx_pcs_eightb_tenb_decoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_rx_pcs_err_flags_sel = "err_flags_wa", // err_flags_wa|err_flags_8b10b
		parameter hssi_8g_rx_pcs_fixed_pat_det = "dis_fixed_patdet", // dis_fixed_patdet|en_fixed_patdet
		parameter hssi_8g_rx_pcs_fixed_pat_num = 4'b1111,
		parameter hssi_8g_rx_pcs_force_signal_detect = "en_force_signal_detect", // en_force_signal_detect|dis_force_signal_detect
		parameter hssi_8g_rx_pcs_gen3_clk_en = "disable_clk", // disable_clk|enable_clk
		parameter hssi_8g_rx_pcs_gen3_rx_clk_sel = "rcvd_clk", // en_dig_clk1_8g|rcvd_clk
		parameter hssi_8g_rx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // en_dig_clk2_8g|tx_pma_clk
		parameter hssi_8g_rx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_rx_pcs_ibm_invalid_code = "dis_ibm_invalid_code", // dis_ibm_invalid_code|en_ibm_invalid_code
		parameter hssi_8g_rx_pcs_invalid_code_flag_only = "dis_invalid_code_only", // dis_invalid_code_only|en_invalid_code_only
		parameter hssi_8g_rx_pcs_pad_or_edb_error_replace = "replace_edb", // replace_edb|replace_edb_dynamic|replace_pad
		parameter hssi_8g_rx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_rx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_rx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_rx_pcs_pipe_if_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_8g_rx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_rx_pcs_polinv_8b10b_dec = "dis_polinv_8b10b_dec", // dis_polinv_8b10b_dec|en_polinv_8b10b_dec
		parameter hssi_8g_rx_pcs_prot_mode = "gige", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic_rm_enable|basic_rm_disable|disabled_prot_mode
		parameter hssi_8g_rx_pcs_rate_match = "dis_rm", // dis_rm|gige_rm|pipe_rm|pipe_rm_0ppm|sw_basic_rm|dw_basic_rm
		parameter hssi_8g_rx_pcs_rate_match_del_thres = "dis_rm_del_thres", // dis_rm_del_thres|gige_rm_del_thres|pipe_rm_del_thres|pipe_rm_0ppm_del_thres|sw_basic_rm_del_thres|dw_basic_rm_del_thres
		parameter hssi_8g_rx_pcs_rate_match_empty_thres = "dis_rm_empty_thres", // dis_rm_empty_thres|gige_rm_empty_thres|pipe_rm_empty_thres|pipe_rm_0ppm_empty_thres|sw_basic_rm_empty_thres|dw_basic_rm_empty_thres
		parameter hssi_8g_rx_pcs_rate_match_full_thres = "dis_rm_full_thres", // dis_rm_full_thres|gige_rm_full_thres|pipe_rm_full_thres|pipe_rm_0ppm_full_thres|sw_basic_rm_full_thres|dw_basic_rm_full_thres
		parameter hssi_8g_rx_pcs_rate_match_ins_thres = "dis_rm_ins_thres", // dis_rm_ins_thres|gige_rm_ins_thres|pipe_rm_ins_thres|pipe_rm_0ppm_ins_thres|sw_basic_rm_ins_thres|dw_basic_rm_ins_thres
		parameter hssi_8g_rx_pcs_rate_match_start_thres = "dis_rm_start_thres", // dis_rm_start_thres|gige_rm_start_thres|pipe_rm_start_thres|pipe_rm_0ppm_start_thres|sw_basic_rm_start_thres|dw_basic_rm_start_thres
		parameter hssi_8g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_rx_pcs_rx_clk2 = "rcvd_clk_clk2", // rcvd_clk_clk2|tx_pma_clock_clk2|refclk_dig2_clk2
		parameter hssi_8g_rx_pcs_rx_clk_free_running = "en_rx_clk_free_run", // dis_rx_clk_free_run|en_rx_clk_free_run
		parameter hssi_8g_rx_pcs_rx_pcs_urst = "en_rx_pcs_urst", // dis_rx_pcs_urst|en_rx_pcs_urst
		parameter hssi_8g_rx_pcs_rx_rcvd_clk = "rcvd_clk_rcvd_clk", // rcvd_clk_rcvd_clk|tx_pma_clock_rcvd_clk
		parameter hssi_8g_rx_pcs_rx_rd_clk = "pld_rx_clk", // pld_rx_clk|rx_clk
		parameter hssi_8g_rx_pcs_rx_refclk = "dis_refclk_sel", // dis_refclk_sel|en_refclk_sel
		parameter hssi_8g_rx_pcs_rx_wr_clk = "rx_clk2_div_1_2_4", // rx_clk2_div_1_2_4|txfifo_rd_clk
		parameter hssi_8g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_rx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_rx_pcs_sync_sm_idle_eios = "dis_syncsm_idle", // dis_syncsm_idle|en_syncsm_idle
		parameter hssi_8g_rx_pcs_test_bus_sel = "tx_testbus", // tx_testbus|tx_ctrl_plane_testbus|wa_testbus|rm_testbus|rx_ctrl_testbus|pcie_ctrl_testbus|rx_ctrl_plane_testbus
		parameter hssi_8g_rx_pcs_tx_rx_parallel_loopback = "dis_plpbk", // dis_plpbk|en_plpbk
		parameter hssi_8g_rx_pcs_wa_boundary_lock_ctrl = "bit_slip", // bit_slip|sync_sm|deterministic_latency|auto_align_pld_ctrl
		parameter hssi_8g_rx_pcs_wa_clk_slip_spacing = 10'b10000,
		parameter hssi_8g_rx_pcs_wa_det_latency_sync_status_beh = "assert_sync_status_non_imm", // assert_sync_status_imm|assert_sync_status_non_imm|dont_care_assert_sync
		parameter hssi_8g_rx_pcs_wa_disp_err_flag = "dis_disp_err_flag", // dis_disp_err_flag|en_disp_err_flag
		parameter hssi_8g_rx_pcs_wa_kchar = "dis_kchar", // dis_kchar|en_kchar
		parameter hssi_8g_rx_pcs_wa_pd = "wa_pd_10", // wa_pd_7|wa_pd_10|wa_pd_20|wa_pd_40|wa_pd_8_sw|wa_pd_8_dw|wa_pd_16_sw|wa_pd_16_dw|wa_pd_32
		parameter hssi_8g_rx_pcs_wa_pd_data = 40'b0,
		parameter hssi_8g_rx_pcs_wa_pd_polarity = "dis_pd_both_pol", // dis_pd_both_pol|en_pd_both_pol|dont_care_both_pol
		parameter hssi_8g_rx_pcs_wa_pld_controlled = "dis_pld_ctrl", // dis_pld_ctrl|pld_ctrl_sw|rising_edge_sensitive_dw|level_sensitive_dw
		parameter hssi_8g_rx_pcs_wa_renumber_data = 6'b0,
		parameter hssi_8g_rx_pcs_wa_rgnumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rknumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rosnumber_data = 2'b0,
		parameter hssi_8g_rx_pcs_wa_rvnumber_data = 13'b0,
		parameter hssi_8g_rx_pcs_wa_sync_sm_ctrl = "gige_sync_sm", // gige_sync_sm|pipe_sync_sm|sw_basic_sync_sm|dw_basic_sync_sm|fibre_channel_sync_sm
		parameter hssi_8g_rx_pcs_wait_cnt = 12'b0,
		
		// parameters for twentynm_hssi_8g_tx_pcs
		parameter hssi_8g_tx_pcs_auto_speed_nego_gen2 = "dis_asn_g2", // dis_asn_g2|en_asn_g2_freq_scal
		parameter hssi_8g_tx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_tx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_tx_pcs_byte_serializer = "dis_bs", // dis_bs|en_bs_by_2|en_bs_by_4
		parameter hssi_8g_tx_pcs_clock_gate_bs_enc = "dis_bs_enc_clk_gating", // dis_bs_enc_clk_gating|en_bs_enc_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_dw_fifowr = "dis_dw_fifowr_clk_gating", // dis_dw_fifowr_clk_gating|en_dw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_fiford = "dis_fiford_clk_gating", // dis_fiford_clk_gating|en_fiford_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_sw_fifowr = "dis_sw_fifowr_clk_gating", // dis_sw_fifowr_clk_gating|en_sw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_observation_in_pld_core = "internal_refclk_b", // internal_refclk_b|internal_fifo_rd_clk|internal_sw_fifo_wr_clk|internal_dw_fifo_wr_clk|internal_tx_clk_out_gen3|internal_pipe_tx_clk_out_gen3
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_tx_pcs_data_selection_8b10b_encoder_input = "normal_data_path", // normal_data_path|gige_idle_conversion
		parameter hssi_8g_tx_pcs_dynamic_clk_switch = "dis_dyn_clk_switch", // dis_dyn_clk_switch|en_dyn_clk_switch
		parameter hssi_8g_tx_pcs_eightb_tenb_disp_ctrl = "dis_disp_ctrl", // dis_disp_ctrl|en_disp_ctrl|en_ib_disp_ctrl
		parameter hssi_8g_tx_pcs_eightb_tenb_encoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_tx_pcs_force_echar = "dis_force_echar", // dis_force_echar|en_force_echar
		parameter hssi_8g_tx_pcs_force_kchar = "dis_force_kchar", // dis_force_kchar|en_force_kchar
		parameter hssi_8g_tx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // dis_tx_clk|tx_pma_clk
		parameter hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel = "func_clk", // dis_tx_pipe_clk|func_clk
		parameter hssi_8g_tx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_tx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_tx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_tx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_tx_pcs_phfifo_write_clk_sel = "pld_tx_clk", // pld_tx_clk|tx_clk
		parameter hssi_8g_tx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_tx_pcs_prot_mode = "basic", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic|disabled_prot_mode
		parameter hssi_8g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_tx_pcs_refclk_b_clk_sel = "tx_pma_clock", // tx_pma_clock|refclk_dig
		parameter hssi_8g_tx_pcs_revloop_back_rm = "dis_rev_loopback_rx_rm", // dis_rev_loopback_rx_rm|en_rev_loopback_rx_rm
		parameter hssi_8g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_tx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_tx_pcs_tx_bitslip = "dis_tx_bitslip", // dis_tx_bitslip|en_tx_bitslip
		parameter hssi_8g_tx_pcs_tx_compliance_controlled_disparity = "dis_txcompliance", // dis_txcompliance|en_txcompliance_pipe2p0|en_txcompliance_pipe3p0
		parameter hssi_8g_tx_pcs_tx_fast_pld_reg = "dis_tx_fast_pld_reg", // dis_tx_fast_pld_reg|en_tx_fast_pld_reg
		parameter hssi_8g_tx_pcs_txclk_freerun = "dis_freerun_tx", // dis_freerun_tx|en_freerun_tx
		parameter hssi_8g_tx_pcs_txpcs_urst = "en_txpcs_urst", // dis_txpcs_urst|en_txpcs_urst
		
		// parameters for twentynm_hssi_common_pcs_pma_interface
		parameter hssi_common_pcs_pma_interface_asn_clk_enable = "false", // false|true
		parameter hssi_common_pcs_pma_interface_asn_enable = "dis_asn", // dis_asn|en_asn
		parameter hssi_common_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|pcie_gen3
		parameter hssi_common_pcs_pma_interface_bypass_early_eios = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pcie_switch = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_ltr = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_sw_done = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_ppm_lock = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_txdetectrx = "false", // false|true
		parameter hssi_common_pcs_pma_interface_cdr_control = "en_cdr_ctrl", // dis_cdr_ctrl|en_cdr_ctrl
		parameter hssi_common_pcs_pma_interface_cid_enable = "en_cid_mode", // dis_cid_mode|en_cid_mode
		parameter hssi_common_pcs_pma_interface_cp_cons_sel = "cp_cons_default", // cp_cons_master|cp_cons_slave_abv|cp_cons_slave_blw|cp_cons_default
		parameter hssi_common_pcs_pma_interface_cp_dwn_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_cp_up_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_blw|ctrl_slave_abv
		parameter hssi_common_pcs_pma_interface_data_mask_count = 16'b100111000100,
		parameter hssi_common_pcs_pma_interface_data_mask_count_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_dft_observation_clock_selection = "dft_clk_obsrv_tx0", // dft_clk_obsrv_tx0|dft_clk_obsrv_tx1|dft_clk_obsrv_tx2|dft_clk_obsrv_tx3|dft_clk_obsrv_tx4|dft_clk_obsrv_rx|dft_clk_obsrv_hclk|dft_clk_obsrv_fref|dft_clk_obsrv_clklow|dft_clk_obsrv_asn0|dft_clk_obsrv_asn1
		parameter hssi_common_pcs_pma_interface_early_eios_counter = 8'b110010,
		parameter hssi_common_pcs_pma_interface_force_freqdet = "force_freqdet_dis", // force_freqdet_dis|force1_freqdet_en|force0_freqdet_en
		parameter hssi_common_pcs_pma_interface_free_run_clk_enable = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ignore_sigdet_g23 = "false", // false|true
		parameter hssi_common_pcs_pma_interface_pc_en_counter = 7'b110111,
		parameter hssi_common_pcs_pma_interface_pc_rst_counter = 5'b10111,
		parameter hssi_common_pcs_pma_interface_pcie_hip_mode = "hip_disable", // hip_enable|hip_disable
		parameter hssi_common_pcs_pma_interface_ph_fifo_reg_mode = "phfifo_reg_mode_dis", // phfifo_reg_mode_dis|phfifo_reg_mode_en
		parameter hssi_common_pcs_pma_interface_phfifo_flush_wait = 6'b100100,
		parameter hssi_common_pcs_pma_interface_pipe_if_g3pcs = "pipe_if_8gpcs", // pipe_if_g3pcs|pipe_if_8gpcs
		parameter hssi_common_pcs_pma_interface_pma_done_counter = 18'b101010101110011000,
		parameter hssi_common_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_common_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_common_pcs_pma_interface_ppm_cnt_rst = "ppm_cnt_rst_dis", // ppm_cnt_rst_dis|ppm_cnt_rst_en
		parameter hssi_common_pcs_pma_interface_ppm_deassert_early = "deassert_early_dis", // deassert_early_dis|deassert_early_en
		parameter hssi_common_pcs_pma_interface_ppm_det_buckets = "ppm_100_bucket", // disable_prot|ppm_300_bucket|ppm_100_bucket|ppm_300_100_bucket
		parameter hssi_common_pcs_pma_interface_ppm_gen1_2_cnt = "cnt_32k", // cnt_32k|cnt_64k
		parameter hssi_common_pcs_pma_interface_ppm_post_eidle_delay = "cnt_200_cycles", // cnt_200_cycles|cnt_400_cycles
		parameter hssi_common_pcs_pma_interface_ppmsel = "ppmsel_300", // ppmsel_disable|ppmsel_5000|ppmsel_2500|ppmsel_1000|ppmsel_500|ppmsel_300|ppmsel_250|ppmsel_200|ppmsel_125|ppmsel_100|ppmsel_62p5|ppm_other
		parameter hssi_common_pcs_pma_interface_prot_mode = "disable_prot_mode", // disable_prot_mode|pipe_g12|pipe_g3|other_protocols
		parameter hssi_common_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_common_pcs_pma_interface_rxvalid_mask = "rxvalid_mask_en", // rxvalid_mask_dis|rxvalid_mask_en
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter = 12'b100111000100,
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_sim_mode = "disable", // disable|enable
		parameter hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en = "true", // false|true
		parameter hssi_common_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_common_pcs_pma_interface_testout_sel = "ppm_det_test", // ppm_det_test|asn_test|pma_pll_test|rxpmaif_test|prbs_gen_test|prbs_ver_test|uhsif_1_test|uhsif_2_test|uhsif_3_test
		parameter hssi_common_pcs_pma_interface_wait_clk_on_off_timer = 4'b100,
		parameter hssi_common_pcs_pma_interface_wait_pipe_synchronizing = 5'b10111,
		parameter hssi_common_pcs_pma_interface_wait_send_syncp_fbkp = 11'b11111010,
		
		// parameters for twentynm_hssi_common_pld_pcs_interface
		parameter hssi_common_pld_pcs_interface_dft_clk_out_en = "dft_clk_out_disable", // dft_clk_out_disable|dft_clk_out_enable
		parameter hssi_common_pld_pcs_interface_dft_clk_out_sel = "teng_rx_dft_clk", // teng_rx_dft_clk|teng_tx_dft_clk|eightg_rx_dft_clk|eightg_tx_dft_clk|pmaif_dft_clk
		parameter hssi_common_pld_pcs_interface_hrdrstctrl_en = "hrst_dis", // hrst_dis|hrst_en
		parameter hssi_common_pld_pcs_interface_pcs_testbus_block_sel = "eightg", // eightg|g3pcs|teng|krfec|pma_if
		parameter hssi_common_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_fifo_rx_pcs
		parameter hssi_fifo_rx_pcs_double_read_mode = "double_read_dis", // double_read_en|double_read_dis
		parameter hssi_fifo_rx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_fifo_tx_pcs
		parameter hssi_fifo_tx_pcs_double_write_mode = "double_write_dis", // double_write_en|double_write_dis
		parameter hssi_fifo_tx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_gen3_rx_pcs
		parameter hssi_gen3_rx_pcs_block_sync = "enable_block_sync", // bypass_block_sync|enable_block_sync
		parameter hssi_gen3_rx_pcs_block_sync_sm = "enable_blk_sync_sm", // disable_blk_sync_sm|enable_blk_sync_sm
		parameter hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn = "enable", // disable|enable
		parameter hssi_gen3_rx_pcs_lpbk_force = "lpbk_frce_dis", // lpbk_frce_dis|lpbk_frce_en
		parameter hssi_gen3_rx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_rx_pcs_rate_match_fifo = "enable_rm_fifo_600ppm", // bypass_rm_fifo|enable_rm_fifo_600ppm|enable_rm_fifo_0ppm
		parameter hssi_gen3_rx_pcs_rate_match_fifo_latency = "regular_latency", // regular_latency|low_latency
		parameter hssi_gen3_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_gen3_rx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_b4gb_par_lpbk = "b4gb_par_lpbk_dis", // b4gb_par_lpbk_dis|b4gb_par_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_force_balign = "en_force_balign", // en_force_balign|dis_force_balign
		parameter hssi_gen3_rx_pcs_rx_ins_del_one_skip = "ins_del_one_skip_en", // ins_del_one_skip_dis|ins_del_one_skip_en
		parameter hssi_gen3_rx_pcs_rx_num_fixed_pat = 4'b1000,
		parameter hssi_gen3_rx_pcs_rx_test_out_sel = "rx_test_out0", // rx_test_out0|rx_test_out1
		parameter hssi_gen3_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_gen3_tx_pcs
		parameter hssi_gen3_tx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_tx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_gen3_tx_pcs_tx_bitslip = 5'b0,
		parameter hssi_gen3_tx_pcs_tx_gbox_byp = "bypass_gbox", // bypass_gbox|enable_gbox
		
		// parameters for twentynm_hssi_krfec_rx_pcs
		parameter hssi_krfec_rx_pcs_blksync_cor_en = "detect", // detect|correct
		parameter hssi_krfec_rx_pcs_bypass_gb = "bypass_dis", // bypass_dis|bypass_en
		parameter hssi_krfec_rx_pcs_clr_ctrl = "both_enabled", // both_enabled|corr_cnt_only|uncorr_cnt_only
		parameter hssi_krfec_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_rx_pcs_dv_start = "with_blklock", // with_blksync|with_blklock
		parameter hssi_krfec_rx_pcs_err_mark_type = "err_mark_10g", // err_mark_10g|err_mark_40g
		parameter hssi_krfec_rx_pcs_error_marking_en = "err_mark_dis", // err_mark_dis|err_mark_en
		parameter hssi_krfec_rx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_krfec_rx_pcs_parity_invalid_enum = 8'b1000,
		parameter hssi_krfec_rx_pcs_parity_valid_num = 4'b100,
		parameter hssi_krfec_rx_pcs_pipeln_blksync = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_descrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errcorrect = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_ind = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_lfsr = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_loc = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_pat = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_gearbox = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_syndrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_trans_dec = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_rx_pcs_receive_order = "receive_lsb", // receive_lsb|receive_msb
		parameter hssi_krfec_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_krfec_rx_pcs_rx_testbus_sel = "overall", // overall|fast_search|fast_search_cntrs|blksync|blksync_cntrs|decoder_master_sm|decoder_master_sm_cntrs|syndrm_sm|syndrm1|syndrm2|errtrap_sm|errtrap_ind1|errtrap_ind2|errtrap_ind3|errtrap_ind4|errtrap_ind5|errtrap_loc|errtrap_pat1|errtrap_pat2|errtrap_pat3|errtrap_pat4|decoder_rd_sm|gb_and_trans
		parameter hssi_krfec_rx_pcs_signal_ok_en = "sig_ok_dis", // sig_ok_dis|sig_ok_en
		parameter hssi_krfec_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_krfec_tx_pcs
		parameter hssi_krfec_tx_pcs_burst_err = "burst_err_dis", // burst_err_dis|burst_err_en
		parameter hssi_krfec_tx_pcs_burst_err_len = "burst_err_len1", // burst_err_len1|burst_err_len2|burst_err_len3|burst_err_len4|burst_err_len5|burst_err_len6|burst_err_len7|burst_err_len8|burst_err_len9|burst_err_len10|burst_err_len11|burst_err_len12|burst_err_len13|burst_err_len14|burst_err_len15|burst_err_len16
		parameter hssi_krfec_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_tx_pcs_enc_frame_query = "enc_query_dis", // enc_query_dis|enc_query_en
		parameter hssi_krfec_tx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_encoder = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_scrambler = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_krfec_tx_pcs_transcode_err = "trans_err_dis", // trans_err_dis|trans_err_en
		parameter hssi_krfec_tx_pcs_transmit_order = "transmit_lsb", // transmit_lsb|transmit_msb
		parameter hssi_krfec_tx_pcs_tx_testbus_sel = "overall", // overall|encoder1|encoder2|scramble1|scramble2|scramble3|gearbox
		
		// parameters for twentynm_hssi_pipe_gen1_2
		parameter hssi_pipe_gen1_2_elec_idle_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_error_replace_pad = "replace_edb", // replace_edb|replace_pad
		parameter hssi_pipe_gen1_2_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_pipe_gen1_2_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen1_2_phystatus_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_phystatus_rst_toggle = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen1_2_pipe_byte_de_serializer_en = "dont_care_bds", // dis_bds|en_bds_by_2|dont_care_bds
		parameter hssi_pipe_gen1_2_prot_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|basic|disabled_prot_mode
		parameter hssi_pipe_gen1_2_reconfig_settings = "{}", // 
		parameter hssi_pipe_gen1_2_rx_pipe_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_pipe_gen1_2_rxdetect_bypass = "dis_rxdetect_bypass", // dis_rxdetect_bypass|en_rxdetect_bypass
		parameter hssi_pipe_gen1_2_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen1_2_tx_pipe_enable = "dis_pipe_tx", // dis_pipe_tx|en_pipe_tx|en_pipe3_tx
		parameter hssi_pipe_gen1_2_txswing = "dis_txswing", // dis_txswing|en_txswing
		
		// parameters for twentynm_hssi_pipe_gen3
		parameter hssi_pipe_gen3_bypass_rx_detection_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_rx_preset = 3'b0,
		parameter hssi_pipe_gen3_bypass_rx_preset_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_tx_coefficent = 18'b0,
		parameter hssi_pipe_gen3_bypass_tx_coefficent_enable = "false", // false|true
		parameter hssi_pipe_gen3_elecidle_delay_g3 = 3'b110,
		parameter hssi_pipe_gen3_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen3_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|disable_pcs
		parameter hssi_pipe_gen3_phy_status_delay_g12 = 3'b101,
		parameter hssi_pipe_gen3_phy_status_delay_g3 = 3'b101,
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g12 = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g3 = "dis_phystatus_rst_toggle_g3", // dis_phystatus_rst_toggle_g3|en_phystatus_rst_toggle_g3
		parameter hssi_pipe_gen3_rate_match_pad_insertion = "dis_rm_fifo_pad_ins", // dis_rm_fifo_pad_ins|en_rm_fifo_pad_ins
		parameter hssi_pipe_gen3_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen3_test_out_sel = "disable_test_out", // tx_test_out|rx_test_out|pipe_test_out1|pipe_test_out2|pipe_test_out3|pipe_ctrl_test_out|disable_test_out
		
		// parameters for twentynm_hssi_rx_pcs_pma_interface
		parameter hssi_rx_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|ten_g_pcs|direct_pld
		parameter hssi_rx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pcs_pma_interface_clkslip_sel = "pld", // pld|slip_eight_g_pcs
		parameter hssi_rx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pcs_pma_interface_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_rx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_rx_pcs_pma_interface_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_rx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_rx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_rx_pcs_pma_interface_prbs_ver = "prbs_off", // prbs_off|prbs_31|prbs_15|prbs_23|prbs_9|prbs_7
		parameter hssi_rx_pcs_pma_interface_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion = "rx_dyn_polinv_dis", // rx_dyn_polinv_dis|rx_dyn_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_lpbk_en = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok = "unforce_sig_ok", // unforce_sig_ok|force_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mask = "prbsmask128", // prbsmask128|prbsmask256|prbsmask512|prbsmask1024
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mode = "teng_mode", // teng_mode|eightg_mode
		parameter hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel = "sel_sig_det", // sel_sig_det|sel_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_static_polarity_inversion = "rx_stat_polinv_dis", // rx_stat_polinv_dis|rx_stat_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en = "uhsif_lpbk_dis", // uhsif_lpbk_dis|uhsif_lpbk_en
		parameter hssi_rx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_rx_pld_pcs_interface
		parameter hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx = "enable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx = "pma_64b_rx", // pma_32b_rx|pma_40b_rx|pma_64b_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_baser_mode_rx|interlaken_mode_rx|sfis_mode_rx|teng_sdi_mode_rx|basic_mode_rx|test_prp_mode_rx|test_prp_krfec_mode_rx|teng_1588_mode_rx|teng_baser_krfec_mode_rx|teng_1588_krfec_mode_rx|basic_krfec_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx = "disabled_prot_mode_rx", // pipe_g1_rx|pipe_g2_rx|pipe_g3_rx|cpri_rx|cpri_rx_tx_rx|gige_rx|gige_1588_rx|basic_rm_enable_rx|basic_rm_disable_rx|disabled_prot_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcie_g1_capable_rx|pcie_g2_capable_rx|pcie_g3_capable_rx|gige_rx|teng_baser_rx|teng_basekr_krfec_rx|fortyg_basekr_krfec_rx|cpri_8b10b_rx|interlaken_rx|sfis_rx|teng_sdi_rx|gige_1588_rx|teng_1588_baser_rx|teng_1588_basekr_krfec_rx|basic_8gpcs_rm_enable_rx|basic_8gpcs_rm_disable_rx|basic_10gpcs_rx|basic_10gpcs_krfec_rx|pcs_direct_rx|prp_rx|prp_krfec_rx|prbs_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx = "teng_mode_rx", // teng_mode_rx|non_teng_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_basekr_mode_rx|fortyg_basekr_mode_rx|teng_1588_basekr_mode_rx|basic_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|eightg_and_g3_pld_fifo_mode_rx|eightg_and_g3_reg_mode_rx|eightg_and_g3_reg_mode_hip_rx|teng_pld_fifo_mode_rx|teng_reg_mode_rx|teng_and_krfec_pld_fifo_mode_rx|teng_and_krfec_reg_mode_rx|pcs_direct_reg_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_block_sel = "pcs_direct", // eightg|teng|pcs_direct
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_rx_clk|pma_rx_clk_user
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_sel = "pld_rx_clk", // pld_rx_clk|pcs_rx_clk
		parameter hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en = "hip_rx_enable", // hip_rx_enable|hip_rx_disable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_rx_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_tx_pcs_pma_interface
		parameter hssi_tx_pcs_pma_interface_bypass_pma_txelecidle = "false", // false|true
		parameter hssi_tx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pcs_pma_interface_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx = "other_prot_mode", // pipe_g12|pipe_g3|other_prot_mode
		parameter hssi_tx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_tx_pcs_pma_interface_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_tx_pcs_pma_interface_pmagate_en = "pmagate_dis", // pmagate_dis|pmagate_en
		parameter hssi_tx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_tx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_tx_pcs_pma_interface_prbs_gen_pat = "prbs_gen_dis", // prbs_gen_dis|prbs_31|prbs_23|prbs_15|prbs_9|prbs_7
		parameter hssi_tx_pcs_pma_interface_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_tx_pcs_pma_interface_sq_wave_num = "sq_wave_4", // sq_wave_1|sq_wave_4|sq_wave_8|sq_wave_6|sq_wave_default
		parameter hssi_tx_pcs_pma_interface_sqwgen_clken = "sqwgen_clk_dis", // sqwgen_clk_dis|sqwgen_clk_en
		parameter hssi_tx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion = "tx_dyn_polinv_dis", // tx_dyn_polinv_dis|tx_dyn_polinv_en
		parameter hssi_tx_pcs_pma_interface_tx_pma_data_sel = "pld_dir", // pld_dir|pcie_gen3|eight_g_pcs|ten_g_pcs|prbs_pat|sq_wave_pat|block_sel_default|registered_uhsif_dat|directed_uhsif_dat
		parameter hssi_tx_pcs_pma_interface_tx_static_polarity_inversion = "tx_stat_polinv_dis", // tx_stat_polinv_dis|tx_stat_polinv_en
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock = "uhsif_filt_stepsz_b4lock_4", // uhsif_filt_stepsz_b4lock_2|uhsif_filt_stepsz_b4lock_4|uhsif_filt_stepsz_b4lock_6|uhsif_filt_stepsz_b4lock_8
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value = 4'b1011,
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock = "uhsif_filt_cntthr_b4lock_16", // uhsif_filt_cntthr_b4lock_8|uhsif_filt_cntthr_b4lock_16|uhsif_filt_cntthr_b4lock_24|uhsif_filt_cntthr_b4lock_32
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period = "uhsif_dcn_test_period_4", // uhsif_dcn_test_period_4|uhsif_dcn_test_period_8|uhsif_dcn_test_period_12|uhsif_dcn_test_period_16
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable = "uhsif_dcn_test_mode_disable", // uhsif_dcn_test_mode_enable|uhsif_dcn_test_mode_disable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh = "uhsif_dzt_cnt_thr_4", // uhsif_dzt_cnt_thr_2|uhsif_dzt_cnt_thr_4|uhsif_dzt_cnt_thr_6|uhsif_dzt_cnt_thr_8
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable = "uhsif_dzt_enable", // uhsif_dzt_disable|uhsif_dzt_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window = "uhsif_dzt_obr_win_32", // uhsif_dzt_obr_win_16|uhsif_dzt_obr_win_32|uhsif_dzt_obr_win_48|uhsif_dzt_obr_win_64
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size = "uhsif_dzt_skipsz_8", // uhsif_dzt_skipsz_4|uhsif_dzt_skipsz_8|uhsif_dzt_skipsz_12|uhsif_dzt_skipsz_16
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel = "uhsif_index_internal", // uhsif_index_internal|uhsif_index_cram
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin = "uhsif_dcn_margin_4", // uhsif_dcn_margin_2|uhsif_dcn_margin_3|uhsif_dcn_margin_4|uhsif_dcn_margin_5
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value = 8'b10000000,
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control = "uhsif_dft_dz_det_val_0", // uhsif_dft_dz_det_val_0|uhsif_dft_dz_det_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control = "uhsif_dft_up_val_0", // uhsif_dft_up_val_0|uhsif_dft_up_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_enable = "uhsif_disable", // uhsif_disable|uhsif_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock = "uhsif_lkd_segsz_aflock_2048", // uhsif_lkd_segsz_aflock_512|uhsif_lkd_segsz_aflock_1024|uhsif_lkd_segsz_aflock_2048|uhsif_lkd_segsz_aflock_4096
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock = "uhsif_lkd_segsz_b4lock_32", // uhsif_lkd_segsz_b4lock_16|uhsif_lkd_segsz_b4lock_32|uhsif_lkd_segsz_b4lock_64|uhsif_lkd_segsz_b4lock_128
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value = 4'b11,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value = 4'b11,
		
		// parameters for twentynm_hssi_tx_pld_pcs_interface
		parameter hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx = "enable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx = "pma_64b_tx", // pma_32b_tx|pma_40b_tx|pma_64b_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_baser_mode_tx|interlaken_mode_tx|sfis_mode_tx|teng_sdi_mode_tx|basic_mode_tx|test_prp_mode_tx|test_prp_krfec_mode_tx|teng_1588_mode_tx|teng_baser_krfec_mode_tx|teng_1588_krfec_mode_tx|basic_krfec_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx = "disabled_prot_mode_tx", // pipe_g1_tx|pipe_g2_tx|pipe_g3_tx|cpri_tx|cpri_rx_tx_tx|gige_tx|gige_1588_tx|basic_tx|disabled_prot_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcie_g1_capable_tx|pcie_g2_capable_tx|pcie_g3_capable_tx|gige_tx|teng_baser_tx|teng_basekr_krfec_tx|fortyg_basekr_krfec_tx|cpri_8b10b_tx|interlaken_tx|sfis_tx|teng_sdi_tx|gige_1588_tx|teng_1588_baser_tx|teng_1588_basekr_krfec_tx|basic_8gpcs_tx|basic_10gpcs_tx|basic_10gpcs_krfec_tx|pcs_direct_tx|uhsif_tx|prp_tx|prp_krfec_tx|prbs_tx|sqwave_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx = "teng_mode_tx", // teng_mode_tx|non_teng_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_basekr_mode_tx|fortyg_basekr_mode_tx|teng_1588_basekr_mode_tx|basic_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|eightg_and_g3_pld_fifo_mode_tx|eightg_and_g3_reg_mode_tx|eightg_and_g3_reg_mode_hip_tx|eightg_and_g3_fastreg_mode_tx|teng_pld_fifo_mode_tx|teng_reg_mode_tx|teng_fastreg_mode_tx|teng_and_krfec_pld_fifo_mode_tx|teng_and_krfec_reg_mode_tx|teng_and_krfec_fastreg_mode_tx|pcs_direct_fastreg_mode_tx|uhsif_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_tx_clk|pma_tx_clk_user
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_source = "teng", // eightg|teng|pma_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_data_source = "hip_disable", // hip_disable|hip_enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en = "delay1_clk_disable", // delay1_clk_enable|delay1_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel = "pld_tx_clk", // pld_tx_clk|pcs_tx_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl = "delay1_path0", // delay1_path0|delay1_path1|delay1_path2|delay1_path3|delay1_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel = "one_ff_delay", // one_ff_delay|two_ff_delay
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en = "delay2_clk_disable", // delay2_clk_enable|delay2_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl = "delay2_path0", // delay2_path0|delay2_path1|delay2_path2|delay2_path3|delay2_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_tx_pld_pcs_interface_reconfig_settings = "{}" // 
	//PARAM_LIST_END
	)
	(
	//PORT_LIST_START
		input wire	[8:0]	in_avmmaddress,
		input wire		in_avmmclk,
		input wire		in_avmmread,
		input wire		in_avmmrstn,
		input wire		in_avmmwrite,
		input wire	[7:0]	in_avmmwritedata,
		input wire	[4:0]	in_bond_pcs10g_in_bot,
		input wire	[4:0]	in_bond_pcs10g_in_top,
		input wire	[12:0]	in_bond_pcs8g_in_bot,
		input wire	[12:0]	in_bond_pcs8g_in_top,
		input wire	[11:0]	in_bond_pmaif_in_bot,
		input wire	[11:0]	in_bond_pmaif_in_top,
		input wire	[63:0]	in_hip_tx_data,
		input wire		in_iocsr_clk,
		input wire	[5:0]	in_iocsr_config,
		input wire		in_iocsr_rdy,
		input wire		in_iocsr_rdy_dly,
		input wire		in_pld_10g_krfec_rx_clr_errblk_cnt,
		input wire		in_pld_10g_krfec_rx_pld_rst_n,
		input wire		in_pld_10g_krfec_tx_pld_rst_n,
		input wire		in_pld_10g_rx_align_clr,
		input wire		in_pld_10g_rx_clr_ber_count,
		input wire		in_pld_10g_rx_rd_en,
		input wire	[6:0]	in_pld_10g_tx_bitslip,
		input wire		in_pld_10g_tx_burst_en,
		input wire		in_pld_10g_tx_data_valid,
		input wire	[1:0]	in_pld_10g_tx_diag_status,
		input wire		in_pld_10g_tx_wordslip,
		input wire		in_pld_8g_a1a2_size,
		input wire		in_pld_8g_bitloc_rev_en,
		input wire		in_pld_8g_byte_rev_en,
		input wire	[2:0]	in_pld_8g_eidleinfersel,
		input wire		in_pld_8g_encdt,
		input wire		in_pld_8g_g3_rx_pld_rst_n,
		input wire		in_pld_8g_g3_tx_pld_rst_n,
		input wire		in_pld_8g_rddisable_tx,
		input wire		in_pld_8g_rdenable_rx,
		input wire		in_pld_8g_refclk_dig2,
		input wire		in_pld_8g_rxpolarity,
		input wire	[4:0]	in_pld_8g_tx_boundary_sel,
		input wire		in_pld_8g_wrdisable_rx,
		input wire		in_pld_8g_wrenable_tx,
		input wire		in_pld_atpg_los_en_n,
		input wire		in_pld_bitslip,
		input wire	[17:0]	in_pld_g3_current_coeff,
		input wire	[2:0]	in_pld_g3_current_rxpreset,
		input wire		in_pld_ltr,
		input wire		in_pld_mem_krfec_atpg_rst_n,
		input wire		in_pld_partial_reconfig,
		input wire		in_pld_pcs_refclk_dig,
		input wire		in_pld_pma_adapt_start,
		input wire		in_pld_pma_csr_test_dis,
		input wire		in_pld_pma_early_eios,
		input wire	[5:0]	in_pld_pma_eye_monitor,
		input wire		in_pld_pma_ltd_b,
		input wire		in_pld_pma_nrpi_freeze,
		input wire	[1:0]	in_pld_pma_pcie_switch,
		input wire		in_pld_pma_ppm_lock,
		input wire	[4:0]	in_pld_pma_reserved_out,
		input wire		in_pld_pma_rs_lpbk_b,
		input wire		in_pld_pma_rx_qpi_pullup,
		input wire		in_pld_pma_rxpma_rstb,
		input wire		in_pld_pma_tx_bitslip,
		input wire		in_pld_pma_tx_bonding_rstb,
		input wire		in_pld_pma_tx_qpi_pulldn,
		input wire		in_pld_pma_tx_qpi_pullup,
		input wire		in_pld_pma_txdetectrx,
		input wire		in_pld_pma_txpma_rstb,
		input wire		in_pld_pmaif_rx_pld_rst_n,
		input wire		in_pld_pmaif_rxclkslip,
		input wire		in_pld_pmaif_tx_pld_rst_n,
		input wire		in_pld_polinv_rx,
		input wire		in_pld_polinv_tx,
		input wire	[1:0]	in_pld_rate,
		input wire	[9:0]	in_pld_reserved_in,
		input wire		in_pld_rx_clk,
		input wire		in_pld_rx_prbs_err_clr,
		input wire		in_pld_scan_mode_n,
		input wire		in_pld_scan_shift_n,
		input wire		in_pld_syncsm_en,
		input wire		in_pld_tx_clk,
		input wire	[17:0]	in_pld_tx_control,
		input wire	[127:0]	in_pld_tx_data,
		input wire		in_pld_txelecidle,
		input wire		in_pld_uhsif_tx_clk,
		input wire		in_pma_adapt_done,
		input wire		in_pma_clklow,
		input wire		in_pma_fref,
		input wire		in_pma_hclk,
		input wire	[1:0]	in_pma_pcie_sw_done,
		input wire		in_pma_pfdmode_lock,
		input wire	[4:0]	in_pma_reserved_in,
		input wire		in_pma_rx_clkdiv_user,
		input wire		in_pma_rx_detect_valid,
		input wire		in_pma_rx_found,
		input wire		in_pma_rx_pma_clk,
		input wire	[63:0]	in_pma_rx_pma_data,
		input wire		in_pma_rx_signal_ok,
		input wire		in_pma_rxpll_lock,
		input wire		in_pma_signal_det,
		input wire	[7:0]	in_pma_testbus,
		input wire		in_pma_tx_clkdiv_user,
		input wire		in_pma_tx_pma_clk,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen1_2,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen3,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pld_pcs_interface,
		output wire		out_blockselect_hssi_10g_rx_pcs,
		output wire		out_blockselect_hssi_10g_tx_pcs,
		output wire		out_blockselect_hssi_8g_rx_pcs,
		output wire		out_blockselect_hssi_8g_tx_pcs,
		output wire		out_blockselect_hssi_common_pcs_pma_interface,
		output wire		out_blockselect_hssi_common_pld_pcs_interface,
		output wire		out_blockselect_hssi_fifo_rx_pcs,
		output wire		out_blockselect_hssi_fifo_tx_pcs,
		output wire		out_blockselect_hssi_gen3_rx_pcs,
		output wire		out_blockselect_hssi_gen3_tx_pcs,
		output wire		out_blockselect_hssi_krfec_rx_pcs,
		output wire		out_blockselect_hssi_krfec_tx_pcs,
		output wire		out_blockselect_hssi_pipe_gen1_2,
		output wire		out_blockselect_hssi_pipe_gen3,
		output wire		out_blockselect_hssi_rx_pcs_pma_interface,
		output wire		out_blockselect_hssi_rx_pld_pcs_interface,
		output wire		out_blockselect_hssi_tx_pcs_pma_interface,
		output wire		out_blockselect_hssi_tx_pld_pcs_interface,
		output wire	[4:0]	out_bond_pcs10g_out_bot,
		output wire	[4:0]	out_bond_pcs10g_out_top,
		output wire	[12:0]	out_bond_pcs8g_out_bot,
		output wire	[12:0]	out_bond_pcs8g_out_top,
		output wire	[11:0]	out_bond_pmaif_out_bot,
		output wire	[11:0]	out_bond_pmaif_out_top,
		output wire	[2:0]	out_hip_clk_out,
		output wire	[7:0]	out_hip_ctrl_out,
		output wire		out_hip_iocsr_rdy,
		output wire		out_hip_iocsr_rdy_dly,
		output wire		out_hip_nfrzdrv,
		output wire		out_hip_npor,
		output wire	[50:0]	out_hip_rx_data,
		output wire		out_hip_usermode,
		output wire		out_pld_10g_krfec_rx_blk_lock,
		output wire	[1:0]	out_pld_10g_krfec_rx_diag_data_status,
		output wire		out_pld_10g_krfec_rx_frame,
		output wire		out_pld_10g_krfec_tx_frame,
		output wire		out_pld_10g_rx_align_val,
		output wire		out_pld_10g_rx_crc32_err,
		output wire		out_pld_10g_rx_data_valid,
		output wire		out_pld_10g_rx_empty,
		output wire		out_pld_10g_rx_fifo_del,
		output wire		out_pld_10g_rx_fifo_insert,
		output wire	[4:0]	out_pld_10g_rx_fifo_num,
		output wire		out_pld_10g_rx_frame_lock,
		output wire		out_pld_10g_rx_hi_ber,
		output wire		out_pld_10g_rx_oflw_err,
		output wire		out_pld_10g_rx_pempty,
		output wire		out_pld_10g_rx_pfull,
		output wire		out_pld_10g_tx_burst_en_exe,
		output wire		out_pld_10g_tx_empty,
		output wire	[3:0]	out_pld_10g_tx_fifo_num,
		output wire		out_pld_10g_tx_full,
		output wire		out_pld_10g_tx_pempty,
		output wire		out_pld_10g_tx_pfull,
		output wire		out_pld_10g_tx_wordslip_exe,
		output wire	[3:0]	out_pld_8g_a1a2_k1k2_flag,
		output wire		out_pld_8g_empty_rmf,
		output wire		out_pld_8g_empty_rx,
		output wire		out_pld_8g_empty_tx,
		output wire		out_pld_8g_full_rmf,
		output wire		out_pld_8g_full_rx,
		output wire		out_pld_8g_full_tx,
		output wire		out_pld_8g_rxelecidle,
		output wire		out_pld_8g_signal_detect_out,
		output wire	[4:0]	out_pld_8g_wa_boundary,
		output wire		out_pld_krfec_tx_alignment,
		output wire		out_pld_pcs_rx_clk_out,
		output wire		out_pld_pcs_tx_clk_out,
		output wire		out_pld_pma_adapt_done,
		output wire		out_pld_pma_clkdiv_rx_user,
		output wire		out_pld_pma_clkdiv_tx_user,
		output wire		out_pld_pma_clklow,
		output wire		out_pld_pma_fref,
		output wire		out_pld_pma_hclk,
		output wire	[1:0]	out_pld_pma_pcie_sw_done,
		output wire		out_pld_pma_pfdmode_lock,
		output wire	[4:0]	out_pld_pma_reserved_in,
		output wire		out_pld_pma_rx_clk_out,
		output wire		out_pld_pma_rx_detect_valid,
		output wire		out_pld_pma_rx_found,
		output wire		out_pld_pma_rxpll_lock,
		output wire		out_pld_pma_signal_ok,
		output wire	[7:0]	out_pld_pma_testbus,
		output wire		out_pld_pma_tx_clk_out,
		output wire		out_pld_pmaif_mask_tx_pll,
		output wire	[9:0]	out_pld_reserved_out,
		output wire	[19:0]	out_pld_rx_control,
		output wire	[127:0]	out_pld_rx_data,
		output wire		out_pld_rx_prbs_done,
		output wire		out_pld_rx_prbs_err,
		output wire	[19:0]	out_pld_test_data,
		output wire		out_pld_uhsif_lock,
		output wire		out_pld_uhsif_tx_clk_out,
		output wire		out_pma_adapt_start,
		output wire		out_pma_atpg_los_en_n,
		output wire		out_pma_csr_test_dis,
		output wire	[17:0]	out_pma_current_coeff,
		output wire	[2:0]	out_pma_current_rxpreset,
		output wire		out_pma_early_eios,
		output wire	[5:0]	out_pma_eye_monitor,
		output wire	[1:0]	out_pma_interface_select,
		output wire		out_pma_ltd_b,
		output wire		out_pma_ltr,
		output wire		out_pma_nfrzdrv,
		output wire		out_pma_nrpi_freeze,
		output wire	[1:0]	out_pma_pcie_switch,
		output wire		out_pma_ppm_lock,
		output wire	[4:0]	out_pma_reserved_out,
		output wire		out_pma_rs_lpbk_b,
		output wire		out_pma_rx_clkslip,
		output wire		out_pma_rx_qpi_pullup,
		output wire		out_pma_rxpma_rstb,
		output wire		out_pma_scan_mode_n,
		output wire		out_pma_scan_shift_n,
		output wire		out_pma_tx_bitslip,
		output wire		out_pma_tx_bonding_rstb,
		output wire		out_pma_tx_elec_idle,
		output wire	[63:0]	out_pma_tx_pma_data,
		output wire		out_pma_tx_qpi_pulldn,
		output wire		out_pma_tx_qpi_pullup,
		output wire		out_pma_tx_txdetectrx,
		output wire		out_pma_txpma_rstb
	//PORT_LIST_END
	);
	//wire declarations
	
	// wires for module twentynm_hssi_fifo_tx_pcs
	wire	[7:0]	w_hssi_fifo_tx_pcs_avmmreaddata;
	wire		w_hssi_fifo_tx_pcs_blockselect;
	wire	[72:0]	w_hssi_fifo_tx_pcs_data_out_10g;
	wire	[63:0]	w_hssi_fifo_tx_pcs_data_out_8g_phase_comp;
	
	// wires for module twentynm_hssi_gen3_rx_pcs
	wire	[7:0]	w_hssi_gen3_rx_pcs_avmmreaddata;
	wire		w_hssi_gen3_rx_pcs_blk_algnd_int;
	wire		w_hssi_gen3_rx_pcs_blk_start;
	wire		w_hssi_gen3_rx_pcs_blockselect;
	wire		w_hssi_gen3_rx_pcs_clkcomp_delete_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_insert_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_overfl_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_undfl_int;
	wire	[31:0]	w_hssi_gen3_rx_pcs_data_out;
	wire		w_hssi_gen3_rx_pcs_data_valid;
	wire		w_hssi_gen3_rx_pcs_ei_det_int;
	wire		w_hssi_gen3_rx_pcs_ei_partial_det_int;
	wire		w_hssi_gen3_rx_pcs_err_decode_int;
	wire		w_hssi_gen3_rx_pcs_i_det_int;
	wire		w_hssi_gen3_rx_pcs_lpbk_blk_start;
	wire	[33:0]	w_hssi_gen3_rx_pcs_lpbk_data;
	wire		w_hssi_gen3_rx_pcs_lpbk_data_valid;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk;
	wire	[39:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n;
	wire		w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int;
	wire	[19:0]	w_hssi_gen3_rx_pcs_rx_test_out;
	wire	[1:0]	w_hssi_gen3_rx_pcs_sync_hdr;
	
	// wires for module twentynm_hssi_krfec_tx_pcs
	wire	[7:0]	w_hssi_krfec_tx_pcs_avmmreaddata;
	wire		w_hssi_krfec_tx_pcs_blockselect;
	wire		w_hssi_krfec_tx_pcs_tx_alignment;
	wire	[63:0]	w_hssi_krfec_tx_pcs_tx_data_out;
	wire		w_hssi_krfec_tx_pcs_tx_frame;
	wire	[19:0]	w_hssi_krfec_tx_pcs_tx_test_data;
	
	// wires for module twentynm_hssi_krfec_rx_pcs
	wire	[7:0]	w_hssi_krfec_rx_pcs_avmmreaddata;
	wire		w_hssi_krfec_rx_pcs_blockselect;
	wire		w_hssi_krfec_rx_pcs_rx_block_lock;
	wire	[9:0]	w_hssi_krfec_rx_pcs_rx_control_out;
	wire	[63:0]	w_hssi_krfec_rx_pcs_rx_data_out;
	wire	[1:0]	w_hssi_krfec_rx_pcs_rx_data_status;
	wire		w_hssi_krfec_rx_pcs_rx_data_valid_out;
	wire		w_hssi_krfec_rx_pcs_rx_frame;
	wire		w_hssi_krfec_rx_pcs_rx_signal_ok_out;
	
	// wires for module twentynm_hssi_rx_pld_pcs_interface
	wire	[7:0]	w_hssi_rx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_rx_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_hip_rx_ctrl;
	wire	[50:0]	w_hssi_rx_pld_pcs_interface_hip_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
	wire	[3:0]	w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary;
	wire		w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_pld_rx_control;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_pld_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
	
	// wires for module twentynm_hssi_common_pld_pcs_interface
	wire	[7:0]	w_hssi_common_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_common_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_hip_cmn_clk;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_hip_cmn_ctrl;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
	wire		w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_hip_npor;
	wire		w_hssi_common_pld_pcs_interface_hip_usermode;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n;
	wire	[17:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel;
	wire		w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_clklow;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_fref;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_hclk;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_pld_pma_reserved_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
	wire	[7:0]	w_hssi_common_pld_pcs_interface_pld_pma_testbus;
	wire		w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
	wire	[9:0]	w_hssi_common_pld_pcs_interface_pld_reserved_out;
	wire	[19:0]	w_hssi_common_pld_pcs_interface_pld_test_data;
	wire		w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
	wire		w_hssi_common_pld_pcs_interface_scan_mode_n;
	
	// wires for module twentynm_hssi_10g_rx_pcs
	wire	[7:0]	w_hssi_10g_rx_pcs_avmmreaddata;
	wire		w_hssi_10g_rx_pcs_blockselect;
	wire		w_hssi_10g_rx_pcs_rx_align_val;
	wire		w_hssi_10g_rx_pcs_rx_blk_lock;
	wire		w_hssi_10g_rx_pcs_rx_clk_out;
	wire		w_hssi_10g_rx_pcs_rx_clk_out_pld_if;
	wire	[19:0]	w_hssi_10g_rx_pcs_rx_control;
	wire		w_hssi_10g_rx_pcs_rx_crc32_err;
	wire	[127:0]	w_hssi_10g_rx_pcs_rx_data;
	wire		w_hssi_10g_rx_pcs_rx_data_valid;
	wire		w_hssi_10g_rx_pcs_rx_dft_clk_out;
	wire	[1:0]	w_hssi_10g_rx_pcs_rx_diag_status;
	wire		w_hssi_10g_rx_pcs_rx_empty;
	wire		w_hssi_10g_rx_pcs_rx_fec_clk;
	wire		w_hssi_10g_rx_pcs_rx_fifo_del;
	wire		w_hssi_10g_rx_pcs_rx_fifo_insert;
	wire	[4:0]	w_hssi_10g_rx_pcs_rx_fifo_num;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_clk;
	wire	[73:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_data;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_en;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_ptr;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_frame_lock;
	wire		w_hssi_10g_rx_pcs_rx_hi_ber;
	wire		w_hssi_10g_rx_pcs_rx_master_clk;
	wire		w_hssi_10g_rx_pcs_rx_master_clk_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_oflw_err;
	wire		w_hssi_10g_rx_pcs_rx_pempty;
	wire		w_hssi_10g_rx_pcs_rx_pfull;
	wire		w_hssi_10g_rx_pcs_rx_random_err;
	wire		w_hssi_10g_rx_pcs_rx_rx_frame;
	
	// wires for module twentynm_hssi_tx_pld_pcs_interface
	wire	[7:0]	w_hssi_tx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_tx_pld_pcs_interface_blockselect;
	wire		w_hssi_tx_pld_pcs_interface_hip_tx_clk;
	wire	[6:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en;
	wire	[17:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control;
	wire	[8:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg;
	wire	[127:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start;
	wire	[4:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle;
	wire	[2:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
	wire		w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
	
	// wires for module twentynm_hssi_tx_pcs_pma_interface
	wire	[7:0]	w_hssi_tx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_tx_pcs_pma_interface_blockselect;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out;
	wire	[4:0]	w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk;
	wire		w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_pma_tx_pma_data;
	wire		w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_1;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_2;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_3;
	
	// wires for module twentynm_hssi_rx_pcs_pma_interface
	wire	[7:0]	w_hssi_rx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_rx_pcs_pma_interface_blockselect;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni;
	wire	[31:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok;
	wire		w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk;
	wire	[5:0]	w_hssi_rx_pcs_pma_interface_pma_eye_monitor;
	wire		w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
	wire		w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test;
	
	// wires for module twentynm_hssi_10g_tx_pcs
	wire	[7:0]	w_hssi_10g_tx_pcs_avmmreaddata;
	wire		w_hssi_10g_tx_pcs_blockselect;
	wire		w_hssi_10g_tx_pcs_distdwn_out_dv;
	wire		w_hssi_10g_tx_pcs_distdwn_out_rden;
	wire		w_hssi_10g_tx_pcs_distdwn_out_wren;
	wire		w_hssi_10g_tx_pcs_distup_out_dv;
	wire		w_hssi_10g_tx_pcs_distup_out_rden;
	wire		w_hssi_10g_tx_pcs_distup_out_wren;
	wire		w_hssi_10g_tx_pcs_tx_burst_en_exe;
	wire		w_hssi_10g_tx_pcs_tx_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pma_if;
	wire	[8:0]	w_hssi_10g_tx_pcs_tx_control_out_krfec;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_data_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_data_valid_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_dft_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_empty;
	wire		w_hssi_10g_tx_pcs_tx_fec_clk;
	wire	[3:0]	w_hssi_10g_tx_pcs_tx_fifo_num;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_rd_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_clk;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_en;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_frame;
	wire		w_hssi_10g_tx_pcs_tx_full;
	wire		w_hssi_10g_tx_pcs_tx_master_clk;
	wire		w_hssi_10g_tx_pcs_tx_master_clk_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_pempty;
	wire		w_hssi_10g_tx_pcs_tx_pfull;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_data;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_gating_val;
	wire	[19:0]	w_hssi_10g_tx_pcs_tx_test_data;
	wire		w_hssi_10g_tx_pcs_tx_wordslip_exe;
	
	// wires for module twentynm_hssi_8g_tx_pcs
	wire	[7:0]	w_hssi_8g_tx_pcs_avmmreaddata;
	wire		w_hssi_8g_tx_pcs_blockselect;
	wire		w_hssi_8g_tx_pcs_clk_out;
	wire		w_hssi_8g_tx_pcs_clk_out_gen3;
	wire	[19:0]	w_hssi_8g_tx_pcs_dataout;
	wire		w_hssi_8g_tx_pcs_dyn_clk_switch_n;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn;
	wire		w_hssi_8g_tx_pcs_g3_tx_pma_rstn;
	wire	[2:0]	w_hssi_8g_tx_pcs_non_gray_eidleinfersel;
	wire		w_hssi_8g_tx_pcs_ph_fifo_overflow;
	wire		w_hssi_8g_tx_pcs_ph_fifo_underflow;
	wire		w_hssi_8g_tx_pcs_phfifo_txdeemph;
	wire	[2:0]	w_hssi_8g_tx_pcs_phfifo_txmargin;
	wire		w_hssi_8g_tx_pcs_phfifo_txswing;
	wire		w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out;
	wire	[1:0]	w_hssi_8g_tx_pcs_pipe_power_down_out;
	wire		w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3;
	wire		w_hssi_8g_tx_pcs_pmaif_asn_rstn;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_refclk_b;
	wire		w_hssi_8g_tx_pcs_refclk_b_reset;
	wire		w_hssi_8g_tx_pcs_rxpolarity_int;
	wire		w_hssi_8g_tx_pcs_soft_reset_wclk1_n;
	wire		w_hssi_8g_tx_pcs_sw_fifo_wr_clk;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_blk_start_out;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_ctrlplane_testbus;
	wire	[31:0]	w_hssi_8g_tx_pcs_tx_data_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_data_valid_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_datak_out;
	wire		w_hssi_8g_tx_pcs_tx_detect_rxloopback_int;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_tx_pipe_clk;
	wire		w_hssi_8g_tx_pcs_tx_pipe_electidle;
	wire		w_hssi_8g_tx_pcs_tx_pipe_soft_reset;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_sync_hdr_out;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_testbus;
	wire		w_hssi_8g_tx_pcs_txcompliance_out;
	wire		w_hssi_8g_tx_pcs_txelecidle_out;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk;
	wire	[63:0]	w_hssi_8g_tx_pcs_wr_data_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_en_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo;
	
	// wires for module twentynm_hssi_pipe_gen3
	wire	[7:0]	w_hssi_pipe_gen3_avmmreaddata;
	wire		w_hssi_pipe_gen3_blockselect;
	wire		w_hssi_pipe_gen3_gen3_clk_sel;
	wire		w_hssi_pipe_gen3_pcs_rst;
	wire		w_hssi_pipe_gen3_phystatus;
	wire	[17:0]	w_hssi_pipe_gen3_pma_current_coeff;
	wire	[2:0]	w_hssi_pipe_gen3_pma_current_rxpreset;
	wire		w_hssi_pipe_gen3_pma_tx_elec_idle;
	wire		w_hssi_pipe_gen3_pma_txdetectrx;
	wire		w_hssi_pipe_gen3_rev_lpbk_8gpcs_out;
	wire		w_hssi_pipe_gen3_rev_lpbk_int;
	wire	[3:0]	w_hssi_pipe_gen3_rx_blk_start;
	wire	[1:0]	w_hssi_pipe_gen3_rx_sync_hdr;
	wire	[63:0]	w_hssi_pipe_gen3_rxd_8gpcs_out;
	wire	[3:0]	w_hssi_pipe_gen3_rxdataskip;
	wire		w_hssi_pipe_gen3_rxelecidle;
	wire		w_hssi_pipe_gen3_rxpolarity_8gpcs_out;
	wire		w_hssi_pipe_gen3_rxpolarity_int;
	wire	[2:0]	w_hssi_pipe_gen3_rxstatus;
	wire		w_hssi_pipe_gen3_rxvalid;
	wire		w_hssi_pipe_gen3_shutdown_clk;
	wire	[19:0]	w_hssi_pipe_gen3_test_out;
	wire		w_hssi_pipe_gen3_tx_blk_start_int;
	wire	[1:0]	w_hssi_pipe_gen3_tx_sync_hdr_int;
	wire	[31:0]	w_hssi_pipe_gen3_txdata_int;
	wire	[3:0]	w_hssi_pipe_gen3_txdatak_int;
	wire		w_hssi_pipe_gen3_txdataskip_int;
	
	// wires for module twentynm_hssi_pipe_gen1_2
	wire	[7:0]	w_hssi_pipe_gen1_2_avmmreaddata;
	wire		w_hssi_pipe_gen1_2_blockselect;
	wire	[17:0]	w_hssi_pipe_gen1_2_current_coeff;
	wire		w_hssi_pipe_gen1_2_phystatus;
	wire		w_hssi_pipe_gen1_2_polarity_inversion_rx;
	wire		w_hssi_pipe_gen1_2_rev_loopbk;
	wire		w_hssi_pipe_gen1_2_rxelecidle;
	wire		w_hssi_pipe_gen1_2_rxelectricalidle_out;
	wire	[2:0]	w_hssi_pipe_gen1_2_rxstatus;
	wire		w_hssi_pipe_gen1_2_rxvalid;
	wire		w_hssi_pipe_gen1_2_tx_elec_idle_out;
	wire		w_hssi_pipe_gen1_2_txdetectrx;
	
	// wires for module twentynm_hssi_gen3_tx_pcs
	wire	[7:0]	w_hssi_gen3_tx_pcs_avmmreaddata;
	wire		w_hssi_gen3_tx_pcs_blockselect;
	wire	[31:0]	w_hssi_gen3_tx_pcs_data_out;
	wire	[35:0]	w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out;
	wire	[31:0]	w_hssi_gen3_tx_pcs_par_lpbk_out;
	wire	[19:0]	w_hssi_gen3_tx_pcs_tx_test_out;
	
	// wires for module twentynm_hssi_8g_rx_pcs
	wire	[3:0]	w_hssi_8g_rx_pcs_a1a2k1k2flag;
	wire	[7:0]	w_hssi_8g_rx_pcs_avmmreaddata;
	wire		w_hssi_8g_rx_pcs_blockselect;
	wire	[19:0]	w_hssi_8g_rx_pcs_chnl_test_bus_out;
	wire		w_hssi_8g_rx_pcs_clock_to_pld;
	wire	[63:0]	w_hssi_8g_rx_pcs_dataout;
	wire		w_hssi_8g_rx_pcs_dis_pc_byte;
	wire		w_hssi_8g_rx_pcs_eidle_detected;
	wire	[2:0]	w_hssi_8g_rx_pcs_eios_det_cdr_ctrl;
	wire		w_hssi_8g_rx_pcs_g3_rx_pma_rstn;
	wire		w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn;
	wire		w_hssi_8g_rx_pcs_gen2ngen1;
	wire	[19:0]	w_hssi_8g_rx_pcs_parallel_rev_loopback;
	wire		w_hssi_8g_rx_pcs_pc_fifo_empty;
	wire		w_hssi_8g_rx_pcs_pcfifofull;
	wire		w_hssi_8g_rx_pcs_phystatus;
	wire	[63:0]	w_hssi_8g_rx_pcs_pipe_data;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_up;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo;
	wire	[7:0]	w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rm_fifo_empty;
	wire		w_hssi_8g_rx_pcs_rm_fifo_full;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_blk_start;
	wire		w_hssi_8g_rx_pcs_rx_clk_out_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clkslip;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_data_valid;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rx_pipe_clk;
	wire		w_hssi_8g_rx_pcs_rx_pipe_soft_reset;
	wire		w_hssi_8g_rx_pcs_rx_pma_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_sync_hdr;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_up;
	wire	[2:0]	w_hssi_8g_rx_pcs_rxstatus;
	wire		w_hssi_8g_rx_pcs_rxvalid;
	wire		w_hssi_8g_rx_pcs_signal_detect_out;
	wire	[4:0]	w_hssi_8g_rx_pcs_word_align_boundary;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk;
	wire	[79:0]	w_hssi_8g_rx_pcs_wr_data_rx_phfifo;
	wire	[31:0]	w_hssi_8g_rx_pcs_wr_data_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo;
	
	// wires for module twentynm_hssi_fifo_rx_pcs
	wire	[7:0]	w_hssi_fifo_rx_pcs_avmmreaddata;
	wire		w_hssi_fifo_rx_pcs_blockselect;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out2_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out_8g_clock_comp;
	wire	[79:0]	w_hssi_fifo_rx_pcs_data_out_8g_phase_comp;
	wire	[39:0]	w_hssi_fifo_rx_pcs_data_out_gen3;
	
	// wires for module twentynm_hssi_common_pcs_pma_interface
	wire	[7:0]	w_hssi_common_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_common_pcs_pma_interface_blockselect;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in;
	wire	[19:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out;
	wire	[7:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus;
	wire		w_hssi_common_pcs_pma_interface_pma_adapt_start;
	wire		w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
	wire		w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
	wire	[17:0]	w_hssi_common_pcs_pma_interface_pma_current_coeff;
	wire	[2:0]	w_hssi_common_pcs_pma_interface_pma_current_rxpreset;
	wire		w_hssi_common_pcs_pma_interface_pma_early_eios;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_interface_select;
	wire		w_hssi_common_pcs_pma_interface_pma_ltd_b;
	wire		w_hssi_common_pcs_pma_interface_pma_ltr;
	wire		w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
	wire		w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_pcie_switch;
	wire		w_hssi_common_pcs_pma_interface_pma_ppm_lock;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_pma_reserved_out;
	wire		w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
	wire		w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up;
	
	
	generate
		
		//module instantiations
		
		// instantiating twentynm_hssi_10g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_rx_pcs
			twentynm_hssi_10g_rx_pcs #(
				.advanced_user_mode(hssi_10g_rx_pcs_advanced_user_mode),
				.align_del(hssi_10g_rx_pcs_align_del),
				.ber_bit_err_total_cnt(hssi_10g_rx_pcs_ber_bit_err_total_cnt),
				.ber_clken(hssi_10g_rx_pcs_ber_clken),
				.ber_xus_timer_window(hssi_10g_rx_pcs_ber_xus_timer_window),
				.bitslip_mode(hssi_10g_rx_pcs_bitslip_mode),
				.blksync_bitslip_type(hssi_10g_rx_pcs_blksync_bitslip_type),
				.blksync_bitslip_wait_cnt(hssi_10g_rx_pcs_blksync_bitslip_wait_cnt),
				.blksync_bitslip_wait_type(hssi_10g_rx_pcs_blksync_bitslip_wait_type),
				.blksync_bypass(hssi_10g_rx_pcs_blksync_bypass),
				.blksync_clken(hssi_10g_rx_pcs_blksync_clken),
				.blksync_enum_invalid_sh_cnt(hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt),
				.blksync_knum_sh_cnt_postlock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock),
				.blksync_knum_sh_cnt_prelock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock),
				.blksync_pipeln(hssi_10g_rx_pcs_blksync_pipeln),
				.clr_errblk_cnt_en(hssi_10g_rx_pcs_clr_errblk_cnt_en),
				.control_del(hssi_10g_rx_pcs_control_del),
				.crcchk_bypass(hssi_10g_rx_pcs_crcchk_bypass),
				.crcchk_clken(hssi_10g_rx_pcs_crcchk_clken),
				.crcchk_inv(hssi_10g_rx_pcs_crcchk_inv),
				.crcchk_pipeln(hssi_10g_rx_pcs_crcchk_pipeln),
				.crcflag_pipeln(hssi_10g_rx_pcs_crcflag_pipeln),
				.ctrl_bit_reverse(hssi_10g_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_10g_rx_pcs_data_bit_reverse),
				.dec64b66b_clken(hssi_10g_rx_pcs_dec64b66b_clken),
				.dec_64b66b_rxsm_bypass(hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass),
				.descrm_bypass(hssi_10g_rx_pcs_descrm_bypass),
				.descrm_clken(hssi_10g_rx_pcs_descrm_clken),
				.descrm_mode(hssi_10g_rx_pcs_descrm_mode),
				.descrm_pipeln(hssi_10g_rx_pcs_descrm_pipeln),
				.dft_clk_out_sel(hssi_10g_rx_pcs_dft_clk_out_sel),
				.dis_signal_ok(hssi_10g_rx_pcs_dis_signal_ok),
				.dispchk_bypass(hssi_10g_rx_pcs_dispchk_bypass),
				.empty_flag_type(hssi_10g_rx_pcs_empty_flag_type),
				.fast_path(hssi_10g_rx_pcs_fast_path),
				.fec_clken(hssi_10g_rx_pcs_fec_clken),
				.fec_enable(hssi_10g_rx_pcs_fec_enable),
				.fifo_double_read(hssi_10g_rx_pcs_fifo_double_read),
				.fifo_stop_rd(hssi_10g_rx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_rx_pcs_fifo_stop_wr),
				.force_align(hssi_10g_rx_pcs_force_align),
				.frmsync_bypass(hssi_10g_rx_pcs_frmsync_bypass),
				.frmsync_clken(hssi_10g_rx_pcs_frmsync_clken),
				.frmsync_enum_scrm(hssi_10g_rx_pcs_frmsync_enum_scrm),
				.frmsync_enum_sync(hssi_10g_rx_pcs_frmsync_enum_sync),
				.frmsync_flag_type(hssi_10g_rx_pcs_frmsync_flag_type),
				.frmsync_knum_sync(hssi_10g_rx_pcs_frmsync_knum_sync),
				.frmsync_mfrm_length(hssi_10g_rx_pcs_frmsync_mfrm_length),
				.frmsync_pipeln(hssi_10g_rx_pcs_frmsync_pipeln),
				.full_flag_type(hssi_10g_rx_pcs_full_flag_type),
				.gb_rx_idwidth(hssi_10g_rx_pcs_gb_rx_idwidth),
				.gb_rx_odwidth(hssi_10g_rx_pcs_gb_rx_odwidth),
				.gbexp_clken(hssi_10g_rx_pcs_gbexp_clken),
				.low_latency_en(hssi_10g_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_10g_rx_pcs_lpbk_mode),
				.master_clk_sel(hssi_10g_rx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_rx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_rx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_rx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_rx_pcs_pld_if_type),
				.prot_mode(hssi_10g_rx_pcs_prot_mode),
				.rand_clken(hssi_10g_rx_pcs_rand_clken),
				.rd_clk_sel(hssi_10g_rx_pcs_rd_clk_sel),
				.rdfifo_clken(hssi_10g_rx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_rx_pcs_reconfig_settings),
				.rx_fifo_write_ctrl(hssi_10g_rx_pcs_rx_fifo_write_ctrl),
				.rx_scrm_width(hssi_10g_rx_pcs_rx_scrm_width),
				.rx_sh_location(hssi_10g_rx_pcs_rx_sh_location),
				.rx_signal_ok_sel(hssi_10g_rx_pcs_rx_signal_ok_sel),
				.rx_sm_bypass(hssi_10g_rx_pcs_rx_sm_bypass),
				.rx_sm_hiber(hssi_10g_rx_pcs_rx_sm_hiber),
				.rx_sm_pipeln(hssi_10g_rx_pcs_rx_sm_pipeln),
				.rx_testbus_sel(hssi_10g_rx_pcs_rx_testbus_sel),
				.rx_true_b2b(hssi_10g_rx_pcs_rx_true_b2b),
				.rxfifo_empty(hssi_10g_rx_pcs_rxfifo_empty),
				.rxfifo_full(hssi_10g_rx_pcs_rxfifo_full),
				.rxfifo_mode(hssi_10g_rx_pcs_rxfifo_mode),
				.rxfifo_pempty(hssi_10g_rx_pcs_rxfifo_pempty),
				.rxfifo_pfull(hssi_10g_rx_pcs_rxfifo_pfull),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.stretch_num_stages(hssi_10g_rx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_rx_pcs_sup_mode),
				.test_mode(hssi_10g_rx_pcs_test_mode),
				.wrfifo_clken(hssi_10g_rx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_rx_pcs_blockselect),
				.rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.rx_control(w_hssi_10g_rx_pcs_rx_control),
				.rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.rx_data(w_hssi_10g_rx_pcs_rx_data),
				.rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.rx_diag_status(w_hssi_10g_rx_pcs_rx_diag_status),
				.rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.rx_fec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.rx_fifo_num(w_hssi_10g_rx_pcs_rx_fifo_num),
				.rx_fifo_rd_ptr(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr),
				.rx_fifo_rd_ptr2(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2),
				.rx_fifo_wr_clk(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.rx_fifo_wr_data(w_hssi_10g_rx_pcs_rx_fifo_wr_data),
				.rx_fifo_wr_en(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.rx_fifo_wr_ptr(w_hssi_10g_rx_pcs_rx_fifo_wr_ptr),
				.rx_fifo_wr_rst_n(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.rx_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_rx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_rx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.rx_control_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0]}),
				.rx_control_in_krfec({w_hssi_krfec_rx_pcs_rx_control_out[9], w_hssi_krfec_rx_pcs_rx_control_out[8], w_hssi_krfec_rx_pcs_rx_control_out[7], w_hssi_krfec_rx_pcs_rx_control_out[6], w_hssi_krfec_rx_pcs_rx_control_out[5], w_hssi_krfec_rx_pcs_rx_control_out[4], w_hssi_krfec_rx_pcs_rx_control_out[3], w_hssi_krfec_rx_pcs_rx_control_out[2], w_hssi_krfec_rx_pcs_rx_control_out[1], w_hssi_krfec_rx_pcs_rx_control_out[0]}),
				.rx_data_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0]}),
				.rx_data_in_krfec({w_hssi_krfec_rx_pcs_rx_data_out[63], w_hssi_krfec_rx_pcs_rx_data_out[62], w_hssi_krfec_rx_pcs_rx_data_out[61], w_hssi_krfec_rx_pcs_rx_data_out[60], w_hssi_krfec_rx_pcs_rx_data_out[59], w_hssi_krfec_rx_pcs_rx_data_out[58], w_hssi_krfec_rx_pcs_rx_data_out[57], w_hssi_krfec_rx_pcs_rx_data_out[56], w_hssi_krfec_rx_pcs_rx_data_out[55], w_hssi_krfec_rx_pcs_rx_data_out[54], w_hssi_krfec_rx_pcs_rx_data_out[53], w_hssi_krfec_rx_pcs_rx_data_out[52], w_hssi_krfec_rx_pcs_rx_data_out[51], w_hssi_krfec_rx_pcs_rx_data_out[50], w_hssi_krfec_rx_pcs_rx_data_out[49], w_hssi_krfec_rx_pcs_rx_data_out[48], w_hssi_krfec_rx_pcs_rx_data_out[47], w_hssi_krfec_rx_pcs_rx_data_out[46], w_hssi_krfec_rx_pcs_rx_data_out[45], w_hssi_krfec_rx_pcs_rx_data_out[44], w_hssi_krfec_rx_pcs_rx_data_out[43], w_hssi_krfec_rx_pcs_rx_data_out[42], w_hssi_krfec_rx_pcs_rx_data_out[41], w_hssi_krfec_rx_pcs_rx_data_out[40], w_hssi_krfec_rx_pcs_rx_data_out[39], w_hssi_krfec_rx_pcs_rx_data_out[38], w_hssi_krfec_rx_pcs_rx_data_out[37], w_hssi_krfec_rx_pcs_rx_data_out[36], w_hssi_krfec_rx_pcs_rx_data_out[35], w_hssi_krfec_rx_pcs_rx_data_out[34], w_hssi_krfec_rx_pcs_rx_data_out[33], w_hssi_krfec_rx_pcs_rx_data_out[32], w_hssi_krfec_rx_pcs_rx_data_out[31], w_hssi_krfec_rx_pcs_rx_data_out[30], w_hssi_krfec_rx_pcs_rx_data_out[29], w_hssi_krfec_rx_pcs_rx_data_out[28], w_hssi_krfec_rx_pcs_rx_data_out[27], w_hssi_krfec_rx_pcs_rx_data_out[26], w_hssi_krfec_rx_pcs_rx_data_out[25], w_hssi_krfec_rx_pcs_rx_data_out[24], w_hssi_krfec_rx_pcs_rx_data_out[23], w_hssi_krfec_rx_pcs_rx_data_out[22], w_hssi_krfec_rx_pcs_rx_data_out[21], w_hssi_krfec_rx_pcs_rx_data_out[20], w_hssi_krfec_rx_pcs_rx_data_out[19], w_hssi_krfec_rx_pcs_rx_data_out[18], w_hssi_krfec_rx_pcs_rx_data_out[17], w_hssi_krfec_rx_pcs_rx_data_out[16], w_hssi_krfec_rx_pcs_rx_data_out[15], w_hssi_krfec_rx_pcs_rx_data_out[14], w_hssi_krfec_rx_pcs_rx_data_out[13], w_hssi_krfec_rx_pcs_rx_data_out[12], w_hssi_krfec_rx_pcs_rx_data_out[11], w_hssi_krfec_rx_pcs_rx_data_out[10], w_hssi_krfec_rx_pcs_rx_data_out[9], w_hssi_krfec_rx_pcs_rx_data_out[8], w_hssi_krfec_rx_pcs_rx_data_out[7], w_hssi_krfec_rx_pcs_rx_data_out[6], w_hssi_krfec_rx_pcs_rx_data_out[5], w_hssi_krfec_rx_pcs_rx_data_out[4], w_hssi_krfec_rx_pcs_rx_data_out[3], w_hssi_krfec_rx_pcs_rx_data_out[2], w_hssi_krfec_rx_pcs_rx_data_out[1], w_hssi_krfec_rx_pcs_rx_data_out[0]}),
				.rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.rx_data_valid_in_krfec(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_10g[73], w_hssi_fifo_rx_pcs_data_out_10g[72], w_hssi_fifo_rx_pcs_data_out_10g[71], w_hssi_fifo_rx_pcs_data_out_10g[70], w_hssi_fifo_rx_pcs_data_out_10g[69], w_hssi_fifo_rx_pcs_data_out_10g[68], w_hssi_fifo_rx_pcs_data_out_10g[67], w_hssi_fifo_rx_pcs_data_out_10g[66], w_hssi_fifo_rx_pcs_data_out_10g[65], w_hssi_fifo_rx_pcs_data_out_10g[64], w_hssi_fifo_rx_pcs_data_out_10g[63], w_hssi_fifo_rx_pcs_data_out_10g[62], w_hssi_fifo_rx_pcs_data_out_10g[61], w_hssi_fifo_rx_pcs_data_out_10g[60], w_hssi_fifo_rx_pcs_data_out_10g[59], w_hssi_fifo_rx_pcs_data_out_10g[58], w_hssi_fifo_rx_pcs_data_out_10g[57], w_hssi_fifo_rx_pcs_data_out_10g[56], w_hssi_fifo_rx_pcs_data_out_10g[55], w_hssi_fifo_rx_pcs_data_out_10g[54], w_hssi_fifo_rx_pcs_data_out_10g[53], w_hssi_fifo_rx_pcs_data_out_10g[52], w_hssi_fifo_rx_pcs_data_out_10g[51], w_hssi_fifo_rx_pcs_data_out_10g[50], w_hssi_fifo_rx_pcs_data_out_10g[49], w_hssi_fifo_rx_pcs_data_out_10g[48], w_hssi_fifo_rx_pcs_data_out_10g[47], w_hssi_fifo_rx_pcs_data_out_10g[46], w_hssi_fifo_rx_pcs_data_out_10g[45], w_hssi_fifo_rx_pcs_data_out_10g[44], w_hssi_fifo_rx_pcs_data_out_10g[43], w_hssi_fifo_rx_pcs_data_out_10g[42], w_hssi_fifo_rx_pcs_data_out_10g[41], w_hssi_fifo_rx_pcs_data_out_10g[40], w_hssi_fifo_rx_pcs_data_out_10g[39], w_hssi_fifo_rx_pcs_data_out_10g[38], w_hssi_fifo_rx_pcs_data_out_10g[37], w_hssi_fifo_rx_pcs_data_out_10g[36], w_hssi_fifo_rx_pcs_data_out_10g[35], w_hssi_fifo_rx_pcs_data_out_10g[34], w_hssi_fifo_rx_pcs_data_out_10g[33], w_hssi_fifo_rx_pcs_data_out_10g[32], w_hssi_fifo_rx_pcs_data_out_10g[31], w_hssi_fifo_rx_pcs_data_out_10g[30], w_hssi_fifo_rx_pcs_data_out_10g[29], w_hssi_fifo_rx_pcs_data_out_10g[28], w_hssi_fifo_rx_pcs_data_out_10g[27], w_hssi_fifo_rx_pcs_data_out_10g[26], w_hssi_fifo_rx_pcs_data_out_10g[25], w_hssi_fifo_rx_pcs_data_out_10g[24], w_hssi_fifo_rx_pcs_data_out_10g[23], w_hssi_fifo_rx_pcs_data_out_10g[22], w_hssi_fifo_rx_pcs_data_out_10g[21], w_hssi_fifo_rx_pcs_data_out_10g[20], w_hssi_fifo_rx_pcs_data_out_10g[19], w_hssi_fifo_rx_pcs_data_out_10g[18], w_hssi_fifo_rx_pcs_data_out_10g[17], w_hssi_fifo_rx_pcs_data_out_10g[16], w_hssi_fifo_rx_pcs_data_out_10g[15], w_hssi_fifo_rx_pcs_data_out_10g[14], w_hssi_fifo_rx_pcs_data_out_10g[13], w_hssi_fifo_rx_pcs_data_out_10g[12], w_hssi_fifo_rx_pcs_data_out_10g[11], w_hssi_fifo_rx_pcs_data_out_10g[10], w_hssi_fifo_rx_pcs_data_out_10g[9], w_hssi_fifo_rx_pcs_data_out_10g[8], w_hssi_fifo_rx_pcs_data_out_10g[7], w_hssi_fifo_rx_pcs_data_out_10g[6], w_hssi_fifo_rx_pcs_data_out_10g[5], w_hssi_fifo_rx_pcs_data_out_10g[4], w_hssi_fifo_rx_pcs_data_out_10g[3], w_hssi_fifo_rx_pcs_data_out_10g[2], w_hssi_fifo_rx_pcs_data_out_10g[1], w_hssi_fifo_rx_pcs_data_out_10g[0]}),
				.rx_fifo_rd_data_dw({w_hssi_fifo_rx_pcs_data_out2_10g[73], w_hssi_fifo_rx_pcs_data_out2_10g[72], w_hssi_fifo_rx_pcs_data_out2_10g[71], w_hssi_fifo_rx_pcs_data_out2_10g[70], w_hssi_fifo_rx_pcs_data_out2_10g[69], w_hssi_fifo_rx_pcs_data_out2_10g[68], w_hssi_fifo_rx_pcs_data_out2_10g[67], w_hssi_fifo_rx_pcs_data_out2_10g[66], w_hssi_fifo_rx_pcs_data_out2_10g[65], w_hssi_fifo_rx_pcs_data_out2_10g[64], w_hssi_fifo_rx_pcs_data_out2_10g[63], w_hssi_fifo_rx_pcs_data_out2_10g[62], w_hssi_fifo_rx_pcs_data_out2_10g[61], w_hssi_fifo_rx_pcs_data_out2_10g[60], w_hssi_fifo_rx_pcs_data_out2_10g[59], w_hssi_fifo_rx_pcs_data_out2_10g[58], w_hssi_fifo_rx_pcs_data_out2_10g[57], w_hssi_fifo_rx_pcs_data_out2_10g[56], w_hssi_fifo_rx_pcs_data_out2_10g[55], w_hssi_fifo_rx_pcs_data_out2_10g[54], w_hssi_fifo_rx_pcs_data_out2_10g[53], w_hssi_fifo_rx_pcs_data_out2_10g[52], w_hssi_fifo_rx_pcs_data_out2_10g[51], w_hssi_fifo_rx_pcs_data_out2_10g[50], w_hssi_fifo_rx_pcs_data_out2_10g[49], w_hssi_fifo_rx_pcs_data_out2_10g[48], w_hssi_fifo_rx_pcs_data_out2_10g[47], w_hssi_fifo_rx_pcs_data_out2_10g[46], w_hssi_fifo_rx_pcs_data_out2_10g[45], w_hssi_fifo_rx_pcs_data_out2_10g[44], w_hssi_fifo_rx_pcs_data_out2_10g[43], w_hssi_fifo_rx_pcs_data_out2_10g[42], w_hssi_fifo_rx_pcs_data_out2_10g[41], w_hssi_fifo_rx_pcs_data_out2_10g[40], w_hssi_fifo_rx_pcs_data_out2_10g[39], w_hssi_fifo_rx_pcs_data_out2_10g[38], w_hssi_fifo_rx_pcs_data_out2_10g[37], w_hssi_fifo_rx_pcs_data_out2_10g[36], w_hssi_fifo_rx_pcs_data_out2_10g[35], w_hssi_fifo_rx_pcs_data_out2_10g[34], w_hssi_fifo_rx_pcs_data_out2_10g[33], w_hssi_fifo_rx_pcs_data_out2_10g[32], w_hssi_fifo_rx_pcs_data_out2_10g[31], w_hssi_fifo_rx_pcs_data_out2_10g[30], w_hssi_fifo_rx_pcs_data_out2_10g[29], w_hssi_fifo_rx_pcs_data_out2_10g[28], w_hssi_fifo_rx_pcs_data_out2_10g[27], w_hssi_fifo_rx_pcs_data_out2_10g[26], w_hssi_fifo_rx_pcs_data_out2_10g[25], w_hssi_fifo_rx_pcs_data_out2_10g[24], w_hssi_fifo_rx_pcs_data_out2_10g[23], w_hssi_fifo_rx_pcs_data_out2_10g[22], w_hssi_fifo_rx_pcs_data_out2_10g[21], w_hssi_fifo_rx_pcs_data_out2_10g[20], w_hssi_fifo_rx_pcs_data_out2_10g[19], w_hssi_fifo_rx_pcs_data_out2_10g[18], w_hssi_fifo_rx_pcs_data_out2_10g[17], w_hssi_fifo_rx_pcs_data_out2_10g[16], w_hssi_fifo_rx_pcs_data_out2_10g[15], w_hssi_fifo_rx_pcs_data_out2_10g[14], w_hssi_fifo_rx_pcs_data_out2_10g[13], w_hssi_fifo_rx_pcs_data_out2_10g[12], w_hssi_fifo_rx_pcs_data_out2_10g[11], w_hssi_fifo_rx_pcs_data_out2_10g[10], w_hssi_fifo_rx_pcs_data_out2_10g[9], w_hssi_fifo_rx_pcs_data_out2_10g[8], w_hssi_fifo_rx_pcs_data_out2_10g[7], w_hssi_fifo_rx_pcs_data_out2_10g[6], w_hssi_fifo_rx_pcs_data_out2_10g[5], w_hssi_fifo_rx_pcs_data_out2_10g[4], w_hssi_fifo_rx_pcs_data_out2_10g[3], w_hssi_fifo_rx_pcs_data_out2_10g[2], w_hssi_fifo_rx_pcs_data_out2_10g[1], w_hssi_fifo_rx_pcs_data_out2_10g[0]}),
				.rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.rx_pma_data({w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0]}),
				.rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.signal_ok_krfec(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_10g_reg(),
				.pld_10g_krfec_rx_blk_lock_10g_txclk_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_txclk_reg(),
				.pld_10g_krfec_rx_frame_10g_reg(),
				.pld_10g_krfec_rx_frame_10g_txclk_reg(),
				.pld_10g_krfec_rx_pld_rst_n_fifo(),
				.pld_10g_krfec_rx_pld_rst_n_reg(),
				.pld_10g_krfec_rx_pld_rst_n_txclk_reg(),
				.pld_10g_rx_align_clr_fifo(),
				.pld_10g_rx_align_clr_reg(),
				.pld_10g_rx_align_clr_txclk_reg(),
				.pld_10g_rx_align_val_fifo(),
				.pld_10g_rx_align_val_reg(),
				.pld_10g_rx_align_val_txclk_reg(),
				.pld_10g_rx_clr_ber_count_reg(),
				.pld_10g_rx_clr_ber_count_txclk_reg(),
				.pld_10g_rx_crc32_err_reg(),
				.pld_10g_rx_crc32_err_txclk_reg(),
				.pld_10g_rx_data_valid_10g_reg(),
				.pld_10g_rx_data_valid_fifo(),
				.pld_10g_rx_data_valid_pcsdirect_reg(),
				.pld_10g_rx_data_valid_txclk_reg(),
				.pld_10g_rx_empty_fifo(),
				.pld_10g_rx_fifo_del_reg(),
				.pld_10g_rx_fifo_del_txclk_reg(),
				.pld_10g_rx_fifo_insert_fifo(),
				.pld_10g_rx_fifo_num_reg(),
				.pld_10g_rx_fifo_num_txclk_reg(),
				.pld_10g_rx_frame_lock_reg(),
				.pld_10g_rx_frame_lock_txclk_reg(),
				.pld_10g_rx_hi_ber_reg(),
				.pld_10g_rx_hi_ber_txclk_reg(),
				.pld_10g_rx_oflw_err_reg(),
				.pld_10g_rx_oflw_err_txclk_reg(),
				.pld_10g_rx_pempty_fifo(),
				.pld_10g_rx_pfull_reg(),
				.pld_10g_rx_pfull_txclk_reg(),
				.pld_10g_rx_rd_en_fifo(),
				.pld_pcs_rx_clk_out_10g_txclk_wire(),
				.pld_pcs_rx_clk_out_10g_wire(),
				.pld_rx_control_10g_reg(),
				.pld_rx_control_10g_txclk_reg(),
				.pld_rx_data_10g_reg(),
				.pld_rx_data_10g_txclk_reg(),
				.pld_rx_prbs_err_10g_txclk_reg(),
				.pld_rx_prbs_err_clr_10g_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_10g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_align_val = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_blk_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_control[19:0] = 20'b0;
				assign w_hssi_10g_rx_pcs_rx_crc32_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_data[127:0] = 128'b0;
				assign w_hssi_10g_rx_pcs_rx_data_valid = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_dft_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_diag_status[1:0] = 2'b0;
				assign w_hssi_10g_rx_pcs_rx_empty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fec_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_del = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_insert = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_data[73:0] = 74'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_frame_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_hi_ber = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_oflw_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pempty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pfull = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_random_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_rx_frame = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_10g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_tx_pcs
			twentynm_hssi_10g_tx_pcs #(
				.advanced_user_mode(hssi_10g_tx_pcs_advanced_user_mode),
				.bitslip_en(hssi_10g_tx_pcs_bitslip_en),
				.bonding_dft_en(hssi_10g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_10g_tx_pcs_bonding_dft_val),
				.comp_cnt(hssi_10g_tx_pcs_comp_cnt),
				.compin_sel(hssi_10g_tx_pcs_compin_sel),
				.crcgen_bypass(hssi_10g_tx_pcs_crcgen_bypass),
				.crcgen_clken(hssi_10g_tx_pcs_crcgen_clken),
				.crcgen_err(hssi_10g_tx_pcs_crcgen_err),
				.crcgen_inv(hssi_10g_tx_pcs_crcgen_inv),
				.ctrl_bit_reverse(hssi_10g_tx_pcs_ctrl_bit_reverse),
				.ctrl_plane_bonding(hssi_10g_tx_pcs_ctrl_plane_bonding),
				.data_bit_reverse(hssi_10g_tx_pcs_data_bit_reverse),
				.dft_clk_out_sel(hssi_10g_tx_pcs_dft_clk_out_sel),
				.dispgen_bypass(hssi_10g_tx_pcs_dispgen_bypass),
				.dispgen_clken(hssi_10g_tx_pcs_dispgen_clken),
				.dispgen_err(hssi_10g_tx_pcs_dispgen_err),
				.dispgen_pipeln(hssi_10g_tx_pcs_dispgen_pipeln),
				.distdwn_bypass_pipeln(hssi_10g_tx_pcs_distdwn_bypass_pipeln),
				.distdwn_master(hssi_10g_tx_pcs_distdwn_master),
				.distup_bypass_pipeln(hssi_10g_tx_pcs_distup_bypass_pipeln),
				.distup_master(hssi_10g_tx_pcs_distup_master),
				.dv_bond(hssi_10g_tx_pcs_dv_bond),
				.empty_flag_type(hssi_10g_tx_pcs_empty_flag_type),
				.enc64b66b_txsm_clken(hssi_10g_tx_pcs_enc64b66b_txsm_clken),
				.enc_64b66b_txsm_bypass(hssi_10g_tx_pcs_enc_64b66b_txsm_bypass),
				.fastpath(hssi_10g_tx_pcs_fastpath),
				.fec_clken(hssi_10g_tx_pcs_fec_clken),
				.fec_enable(hssi_10g_tx_pcs_fec_enable),
				.fifo_double_write(hssi_10g_tx_pcs_fifo_double_write),
				.fifo_reg_fast(hssi_10g_tx_pcs_fifo_reg_fast),
				.fifo_stop_rd(hssi_10g_tx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_tx_pcs_fifo_stop_wr),
				.frmgen_burst(hssi_10g_tx_pcs_frmgen_burst),
				.frmgen_bypass(hssi_10g_tx_pcs_frmgen_bypass),
				.frmgen_clken(hssi_10g_tx_pcs_frmgen_clken),
				.frmgen_mfrm_length(hssi_10g_tx_pcs_frmgen_mfrm_length),
				.frmgen_pipeln(hssi_10g_tx_pcs_frmgen_pipeln),
				.frmgen_pyld_ins(hssi_10g_tx_pcs_frmgen_pyld_ins),
				.frmgen_wordslip(hssi_10g_tx_pcs_frmgen_wordslip),
				.full_flag_type(hssi_10g_tx_pcs_full_flag_type),
				.gb_pipeln_bypass(hssi_10g_tx_pcs_gb_pipeln_bypass),
				.gb_tx_idwidth(hssi_10g_tx_pcs_gb_tx_idwidth),
				.gb_tx_odwidth(hssi_10g_tx_pcs_gb_tx_odwidth),
				.gbred_clken(hssi_10g_tx_pcs_gbred_clken),
				.indv(hssi_10g_tx_pcs_indv),
				.low_latency_en(hssi_10g_tx_pcs_low_latency_en),
				.master_clk_sel(hssi_10g_tx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_tx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_tx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_tx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_tx_pcs_pld_if_type),
				.prot_mode(hssi_10g_tx_pcs_prot_mode),
				.pseudo_random(hssi_10g_tx_pcs_pseudo_random),
				.pseudo_seed_a(hssi_10g_tx_pcs_pseudo_seed_a),
				.pseudo_seed_b(hssi_10g_tx_pcs_pseudo_seed_b),
				.random_disp(hssi_10g_tx_pcs_random_disp),
				.rdfifo_clken(hssi_10g_tx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_tx_pcs_reconfig_settings),
				.scrm_bypass(hssi_10g_tx_pcs_scrm_bypass),
				.scrm_clken(hssi_10g_tx_pcs_scrm_clken),
				.scrm_mode(hssi_10g_tx_pcs_scrm_mode),
				.scrm_pipeln(hssi_10g_tx_pcs_scrm_pipeln),
				.sh_err(hssi_10g_tx_pcs_sh_err),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sop_mark(hssi_10g_tx_pcs_sop_mark),
				.stretch_num_stages(hssi_10g_tx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_tx_pcs_sup_mode),
				.test_mode(hssi_10g_tx_pcs_test_mode),
				.tx_scrm_err(hssi_10g_tx_pcs_tx_scrm_err),
				.tx_scrm_width(hssi_10g_tx_pcs_tx_scrm_width),
				.tx_sh_location(hssi_10g_tx_pcs_tx_sh_location),
				.tx_sm_bypass(hssi_10g_tx_pcs_tx_sm_bypass),
				.tx_sm_pipeln(hssi_10g_tx_pcs_tx_sm_pipeln),
				.tx_testbus_sel(hssi_10g_tx_pcs_tx_testbus_sel),
				.txfifo_empty(hssi_10g_tx_pcs_txfifo_empty),
				.txfifo_full(hssi_10g_tx_pcs_txfifo_full),
				.txfifo_mode(hssi_10g_tx_pcs_txfifo_mode),
				.txfifo_pempty(hssi_10g_tx_pcs_txfifo_pempty),
				.txfifo_pfull(hssi_10g_tx_pcs_txfifo_pfull),
				.wr_clk_sel(hssi_10g_tx_pcs_wr_clk_sel),
				.wrfifo_clken(hssi_10g_tx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_tx_pcs_blockselect),
				.distdwn_out_dv(w_hssi_10g_tx_pcs_distdwn_out_dv),
				.distdwn_out_rden(w_hssi_10g_tx_pcs_distdwn_out_rden),
				.distdwn_out_wren(w_hssi_10g_tx_pcs_distdwn_out_wren),
				.distup_out_dv(w_hssi_10g_tx_pcs_distup_out_dv),
				.distup_out_rden(w_hssi_10g_tx_pcs_distup_out_rden),
				.distup_out_wren(w_hssi_10g_tx_pcs_distup_out_wren),
				.tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pma_if(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.tx_control_out_krfec(w_hssi_10g_tx_pcs_tx_control_out_krfec),
				.tx_data_out_krfec(w_hssi_10g_tx_pcs_tx_data_out_krfec),
				.tx_data_valid_out_krfec(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.tx_fec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_fifo_num(w_hssi_10g_tx_pcs_tx_fifo_num),
				.tx_fifo_rd_ptr(w_hssi_10g_tx_pcs_tx_fifo_rd_ptr),
				.tx_fifo_wr_clk(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.tx_fifo_wr_data(w_hssi_10g_tx_pcs_tx_fifo_wr_data),
				.tx_fifo_wr_data_dw(w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw),
				.tx_fifo_wr_en(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.tx_fifo_wr_ptr(w_hssi_10g_tx_pcs_tx_fifo_wr_ptr),
				.tx_fifo_wr_rst_n(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.tx_full(w_hssi_10g_tx_pcs_tx_full),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				.tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.tx_pma_data(w_hssi_10g_tx_pcs_tx_pma_data),
				.tx_pma_gating_val(w_hssi_10g_tx_pcs_tx_pma_gating_val),
				.tx_test_data(w_hssi_10g_tx_pcs_tx_test_data),
				.tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.distdwn_in_dv(in_bond_pcs10g_in_bot[2]),
				.distdwn_in_rden(in_bond_pcs10g_in_bot[4]),
				.distdwn_in_wren(in_bond_pcs10g_in_bot[3]),
				.distup_in_dv(in_bond_pcs10g_in_top[2]),
				.distup_in_rden(in_bond_pcs10g_in_top[4]),
				.distup_in_wren(in_bond_pcs10g_in_top[3]),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_tx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_tx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.tx_bitslip({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0]}),
				.tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.tx_control({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0]}),
				.tx_control_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0]}),
				.tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0]}),
				.tx_data_in_krfec({w_hssi_krfec_tx_pcs_tx_data_out[63], w_hssi_krfec_tx_pcs_tx_data_out[62], w_hssi_krfec_tx_pcs_tx_data_out[61], w_hssi_krfec_tx_pcs_tx_data_out[60], w_hssi_krfec_tx_pcs_tx_data_out[59], w_hssi_krfec_tx_pcs_tx_data_out[58], w_hssi_krfec_tx_pcs_tx_data_out[57], w_hssi_krfec_tx_pcs_tx_data_out[56], w_hssi_krfec_tx_pcs_tx_data_out[55], w_hssi_krfec_tx_pcs_tx_data_out[54], w_hssi_krfec_tx_pcs_tx_data_out[53], w_hssi_krfec_tx_pcs_tx_data_out[52], w_hssi_krfec_tx_pcs_tx_data_out[51], w_hssi_krfec_tx_pcs_tx_data_out[50], w_hssi_krfec_tx_pcs_tx_data_out[49], w_hssi_krfec_tx_pcs_tx_data_out[48], w_hssi_krfec_tx_pcs_tx_data_out[47], w_hssi_krfec_tx_pcs_tx_data_out[46], w_hssi_krfec_tx_pcs_tx_data_out[45], w_hssi_krfec_tx_pcs_tx_data_out[44], w_hssi_krfec_tx_pcs_tx_data_out[43], w_hssi_krfec_tx_pcs_tx_data_out[42], w_hssi_krfec_tx_pcs_tx_data_out[41], w_hssi_krfec_tx_pcs_tx_data_out[40], w_hssi_krfec_tx_pcs_tx_data_out[39], w_hssi_krfec_tx_pcs_tx_data_out[38], w_hssi_krfec_tx_pcs_tx_data_out[37], w_hssi_krfec_tx_pcs_tx_data_out[36], w_hssi_krfec_tx_pcs_tx_data_out[35], w_hssi_krfec_tx_pcs_tx_data_out[34], w_hssi_krfec_tx_pcs_tx_data_out[33], w_hssi_krfec_tx_pcs_tx_data_out[32], w_hssi_krfec_tx_pcs_tx_data_out[31], w_hssi_krfec_tx_pcs_tx_data_out[30], w_hssi_krfec_tx_pcs_tx_data_out[29], w_hssi_krfec_tx_pcs_tx_data_out[28], w_hssi_krfec_tx_pcs_tx_data_out[27], w_hssi_krfec_tx_pcs_tx_data_out[26], w_hssi_krfec_tx_pcs_tx_data_out[25], w_hssi_krfec_tx_pcs_tx_data_out[24], w_hssi_krfec_tx_pcs_tx_data_out[23], w_hssi_krfec_tx_pcs_tx_data_out[22], w_hssi_krfec_tx_pcs_tx_data_out[21], w_hssi_krfec_tx_pcs_tx_data_out[20], w_hssi_krfec_tx_pcs_tx_data_out[19], w_hssi_krfec_tx_pcs_tx_data_out[18], w_hssi_krfec_tx_pcs_tx_data_out[17], w_hssi_krfec_tx_pcs_tx_data_out[16], w_hssi_krfec_tx_pcs_tx_data_out[15], w_hssi_krfec_tx_pcs_tx_data_out[14], w_hssi_krfec_tx_pcs_tx_data_out[13], w_hssi_krfec_tx_pcs_tx_data_out[12], w_hssi_krfec_tx_pcs_tx_data_out[11], w_hssi_krfec_tx_pcs_tx_data_out[10], w_hssi_krfec_tx_pcs_tx_data_out[9], w_hssi_krfec_tx_pcs_tx_data_out[8], w_hssi_krfec_tx_pcs_tx_data_out[7], w_hssi_krfec_tx_pcs_tx_data_out[6], w_hssi_krfec_tx_pcs_tx_data_out[5], w_hssi_krfec_tx_pcs_tx_data_out[4], w_hssi_krfec_tx_pcs_tx_data_out[3], w_hssi_krfec_tx_pcs_tx_data_out[2], w_hssi_krfec_tx_pcs_tx_data_out[1], w_hssi_krfec_tx_pcs_tx_data_out[0]}),
				.tx_data_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0]}),
				.tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.tx_diag_status({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0]}),
				.tx_fifo_rd_data({w_hssi_fifo_tx_pcs_data_out_10g[72], w_hssi_fifo_tx_pcs_data_out_10g[71], w_hssi_fifo_tx_pcs_data_out_10g[70], w_hssi_fifo_tx_pcs_data_out_10g[69], w_hssi_fifo_tx_pcs_data_out_10g[68], w_hssi_fifo_tx_pcs_data_out_10g[67], w_hssi_fifo_tx_pcs_data_out_10g[66], w_hssi_fifo_tx_pcs_data_out_10g[65], w_hssi_fifo_tx_pcs_data_out_10g[64], w_hssi_fifo_tx_pcs_data_out_10g[63], w_hssi_fifo_tx_pcs_data_out_10g[62], w_hssi_fifo_tx_pcs_data_out_10g[61], w_hssi_fifo_tx_pcs_data_out_10g[60], w_hssi_fifo_tx_pcs_data_out_10g[59], w_hssi_fifo_tx_pcs_data_out_10g[58], w_hssi_fifo_tx_pcs_data_out_10g[57], w_hssi_fifo_tx_pcs_data_out_10g[56], w_hssi_fifo_tx_pcs_data_out_10g[55], w_hssi_fifo_tx_pcs_data_out_10g[54], w_hssi_fifo_tx_pcs_data_out_10g[53], w_hssi_fifo_tx_pcs_data_out_10g[52], w_hssi_fifo_tx_pcs_data_out_10g[51], w_hssi_fifo_tx_pcs_data_out_10g[50], w_hssi_fifo_tx_pcs_data_out_10g[49], w_hssi_fifo_tx_pcs_data_out_10g[48], w_hssi_fifo_tx_pcs_data_out_10g[47], w_hssi_fifo_tx_pcs_data_out_10g[46], w_hssi_fifo_tx_pcs_data_out_10g[45], w_hssi_fifo_tx_pcs_data_out_10g[44], w_hssi_fifo_tx_pcs_data_out_10g[43], w_hssi_fifo_tx_pcs_data_out_10g[42], w_hssi_fifo_tx_pcs_data_out_10g[41], w_hssi_fifo_tx_pcs_data_out_10g[40], w_hssi_fifo_tx_pcs_data_out_10g[39], w_hssi_fifo_tx_pcs_data_out_10g[38], w_hssi_fifo_tx_pcs_data_out_10g[37], w_hssi_fifo_tx_pcs_data_out_10g[36], w_hssi_fifo_tx_pcs_data_out_10g[35], w_hssi_fifo_tx_pcs_data_out_10g[34], w_hssi_fifo_tx_pcs_data_out_10g[33], w_hssi_fifo_tx_pcs_data_out_10g[32], w_hssi_fifo_tx_pcs_data_out_10g[31], w_hssi_fifo_tx_pcs_data_out_10g[30], w_hssi_fifo_tx_pcs_data_out_10g[29], w_hssi_fifo_tx_pcs_data_out_10g[28], w_hssi_fifo_tx_pcs_data_out_10g[27], w_hssi_fifo_tx_pcs_data_out_10g[26], w_hssi_fifo_tx_pcs_data_out_10g[25], w_hssi_fifo_tx_pcs_data_out_10g[24], w_hssi_fifo_tx_pcs_data_out_10g[23], w_hssi_fifo_tx_pcs_data_out_10g[22], w_hssi_fifo_tx_pcs_data_out_10g[21], w_hssi_fifo_tx_pcs_data_out_10g[20], w_hssi_fifo_tx_pcs_data_out_10g[19], w_hssi_fifo_tx_pcs_data_out_10g[18], w_hssi_fifo_tx_pcs_data_out_10g[17], w_hssi_fifo_tx_pcs_data_out_10g[16], w_hssi_fifo_tx_pcs_data_out_10g[15], w_hssi_fifo_tx_pcs_data_out_10g[14], w_hssi_fifo_tx_pcs_data_out_10g[13], w_hssi_fifo_tx_pcs_data_out_10g[12], w_hssi_fifo_tx_pcs_data_out_10g[11], w_hssi_fifo_tx_pcs_data_out_10g[10], w_hssi_fifo_tx_pcs_data_out_10g[9], w_hssi_fifo_tx_pcs_data_out_10g[8], w_hssi_fifo_tx_pcs_data_out_10g[7], w_hssi_fifo_tx_pcs_data_out_10g[6], w_hssi_fifo_tx_pcs_data_out_10g[5], w_hssi_fifo_tx_pcs_data_out_10g[4], w_hssi_fifo_tx_pcs_data_out_10g[3], w_hssi_fifo_tx_pcs_data_out_10g[2], w_hssi_fifo_tx_pcs_data_out_10g[1], w_hssi_fifo_tx_pcs_data_out_10g[0]}),
				.tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_10g_reg(),
				.pld_10g_krfec_tx_pld_rst_n_fifo(),
				.pld_10g_krfec_tx_pld_rst_n_reg(),
				.pld_10g_tx_bitslip_reg(),
				.pld_10g_tx_burst_en_exe_reg(),
				.pld_10g_tx_data_valid_10g_reg(),
				.pld_10g_tx_data_valid_fifo(),
				.pld_10g_tx_data_valid_reg(),
				.pld_10g_tx_diag_status_reg(),
				.pld_10g_tx_empty_reg(),
				.pld_10g_tx_fifo_num_reg(),
				.pld_10g_tx_full_fifo(),
				.pld_10g_tx_full_reg(),
				.pld_10g_tx_pempty_reg(),
				.pld_10g_tx_pfull_fifo(),
				.pld_10g_tx_wordslip_exe_reg(),
				.pld_10g_tx_wordslip_reg(),
				.pld_pcs_tx_clk_out_10g_wire(),
				.pld_tx_burst_en_reg(),
				.pld_tx_control_lo_10g_reg(),
				.pld_tx_data_10g_fifo(),
				.pld_tx_data_lo_10g_reg()
			);
		end // if generate
		else begin
				assign w_hssi_10g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_burst_en_exe = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pma_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_control_out_krfec[8:0] = 9'b0;
				assign w_hssi_10g_tx_pcs_tx_data_out_krfec[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_data_valid_out_krfec = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_dft_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_empty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fec_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_full = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_pempty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pfull = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_gating_val[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_test_data[19:0] = 20'b0;
				assign w_hssi_10g_tx_pcs_tx_wordslip_exe = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_rx_pcs
			twentynm_hssi_8g_rx_pcs #(
				.auto_error_replacement(hssi_8g_rx_pcs_auto_error_replacement),
				.auto_speed_nego(hssi_8g_rx_pcs_auto_speed_nego),
				.bit_reversal(hssi_8g_rx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_rx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_rx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_rx_pcs_bypass_pipeline_reg),
				.byte_deserializer(hssi_8g_rx_pcs_byte_deserializer),
				.cdr_ctrl_rxvalid_mask(hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask),
				.clkcmp_pattern_n(hssi_8g_rx_pcs_clkcmp_pattern_n),
				.clkcmp_pattern_p(hssi_8g_rx_pcs_clkcmp_pattern_p),
				.clock_gate_bds_dec_asn(hssi_8g_rx_pcs_clock_gate_bds_dec_asn),
				.clock_gate_cdr_eidle(hssi_8g_rx_pcs_clock_gate_cdr_eidle),
				.clock_gate_dw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk),
				.clock_gate_dw_rm_rd(hssi_8g_rx_pcs_clock_gate_dw_rm_rd),
				.clock_gate_dw_rm_wr(hssi_8g_rx_pcs_clock_gate_dw_rm_wr),
				.clock_gate_dw_wa(hssi_8g_rx_pcs_clock_gate_dw_wa),
				.clock_gate_pc_rdclk(hssi_8g_rx_pcs_clock_gate_pc_rdclk),
				.clock_gate_sw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk),
				.clock_gate_sw_rm_rd(hssi_8g_rx_pcs_clock_gate_sw_rm_rd),
				.clock_gate_sw_rm_wr(hssi_8g_rx_pcs_clock_gate_sw_rm_wr),
				.clock_gate_sw_wa(hssi_8g_rx_pcs_clock_gate_sw_wa),
				.clock_observation_in_pld_core(hssi_8g_rx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_rx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_rx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_rx_pcs_ctrl_plane_bonding_distribution),
				.eidle_entry_eios(hssi_8g_rx_pcs_eidle_entry_eios),
				.eidle_entry_iei(hssi_8g_rx_pcs_eidle_entry_iei),
				.eidle_entry_sd(hssi_8g_rx_pcs_eidle_entry_sd),
				.eightb_tenb_decoder(hssi_8g_rx_pcs_eightb_tenb_decoder),
				.err_flags_sel(hssi_8g_rx_pcs_err_flags_sel),
				.fixed_pat_det(hssi_8g_rx_pcs_fixed_pat_det),
				.fixed_pat_num(hssi_8g_rx_pcs_fixed_pat_num),
				.force_signal_detect(hssi_8g_rx_pcs_force_signal_detect),
				.gen3_clk_en(hssi_8g_rx_pcs_gen3_clk_en),
				.gen3_rx_clk_sel(hssi_8g_rx_pcs_gen3_rx_clk_sel),
				.gen3_tx_clk_sel(hssi_8g_rx_pcs_gen3_tx_clk_sel),
				.hip_mode(hssi_8g_rx_pcs_hip_mode),
				.ibm_invalid_code(hssi_8g_rx_pcs_ibm_invalid_code),
				.invalid_code_flag_only(hssi_8g_rx_pcs_invalid_code_flag_only),
				.pad_or_edb_error_replace(hssi_8g_rx_pcs_pad_or_edb_error_replace),
				.pcs_bypass(hssi_8g_rx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_rx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_rx_pcs_phase_compensation_fifo),
				.pipe_if_enable(hssi_8g_rx_pcs_pipe_if_enable),
				.pma_dw(hssi_8g_rx_pcs_pma_dw),
				.polinv_8b10b_dec(hssi_8g_rx_pcs_polinv_8b10b_dec),
				.prot_mode(hssi_8g_rx_pcs_prot_mode),
				.rate_match(hssi_8g_rx_pcs_rate_match),
				.rate_match_del_thres(hssi_8g_rx_pcs_rate_match_del_thres),
				.rate_match_empty_thres(hssi_8g_rx_pcs_rate_match_empty_thres),
				.rate_match_full_thres(hssi_8g_rx_pcs_rate_match_full_thres),
				.rate_match_ins_thres(hssi_8g_rx_pcs_rate_match_ins_thres),
				.rate_match_start_thres(hssi_8g_rx_pcs_rate_match_start_thres),
				.reconfig_settings(hssi_8g_rx_pcs_reconfig_settings),
				.rx_clk2(hssi_8g_rx_pcs_rx_clk2),
				.rx_clk_free_running(hssi_8g_rx_pcs_rx_clk_free_running),
				.rx_pcs_urst(hssi_8g_rx_pcs_rx_pcs_urst),
				.rx_rcvd_clk(hssi_8g_rx_pcs_rx_rcvd_clk),
				.rx_rd_clk(hssi_8g_rx_pcs_rx_rd_clk),
				.rx_refclk(hssi_8g_rx_pcs_rx_refclk),
				.rx_wr_clk(hssi_8g_rx_pcs_rx_wr_clk),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_rx_pcs_sup_mode),
				.symbol_swap(hssi_8g_rx_pcs_symbol_swap),
				.sync_sm_idle_eios(hssi_8g_rx_pcs_sync_sm_idle_eios),
				.test_bus_sel(hssi_8g_rx_pcs_test_bus_sel),
				.tx_rx_parallel_loopback(hssi_8g_rx_pcs_tx_rx_parallel_loopback),
				.wa_boundary_lock_ctrl(hssi_8g_rx_pcs_wa_boundary_lock_ctrl),
				.wa_clk_slip_spacing(hssi_8g_rx_pcs_wa_clk_slip_spacing),
				.wa_det_latency_sync_status_beh(hssi_8g_rx_pcs_wa_det_latency_sync_status_beh),
				.wa_disp_err_flag(hssi_8g_rx_pcs_wa_disp_err_flag),
				.wa_kchar(hssi_8g_rx_pcs_wa_kchar),
				.wa_pd(hssi_8g_rx_pcs_wa_pd),
				.wa_pd_data(hssi_8g_rx_pcs_wa_pd_data),
				.wa_pd_polarity(hssi_8g_rx_pcs_wa_pd_polarity),
				.wa_pld_controlled(hssi_8g_rx_pcs_wa_pld_controlled),
				.wa_renumber_data(hssi_8g_rx_pcs_wa_renumber_data),
				.wa_rgnumber_data(hssi_8g_rx_pcs_wa_rgnumber_data),
				.wa_rknumber_data(hssi_8g_rx_pcs_wa_rknumber_data),
				.wa_rosnumber_data(hssi_8g_rx_pcs_wa_rosnumber_data),
				.wa_rvnumber_data(hssi_8g_rx_pcs_wa_rvnumber_data),
				.wa_sync_sm_ctrl(hssi_8g_rx_pcs_wa_sync_sm_ctrl),
				.wait_cnt(hssi_8g_rx_pcs_wait_cnt)
			) inst_twentynm_hssi_8g_rx_pcs (
				// OUTPUTS
				.a1a2k1k2flag(w_hssi_8g_rx_pcs_a1a2k1k2flag),
				.avmmreaddata(w_hssi_8g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_rx_pcs_blockselect),
				.chnl_test_bus_out(w_hssi_8g_rx_pcs_chnl_test_bus_out),
				.clock_to_pld(w_hssi_8g_rx_pcs_clock_to_pld),
				.dataout(w_hssi_8g_rx_pcs_dataout),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidle_detected(w_hssi_8g_rx_pcs_eidle_detected),
				.eios_det_cdr_ctrl(w_hssi_8g_rx_pcs_eios_det_cdr_ctrl),
				.g3_rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.g3_rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.gen2ngen1(w_hssi_8g_rx_pcs_gen2ngen1),
				.parallel_rev_loopback(w_hssi_8g_rx_pcs_parallel_rev_loopback),
				.pc_fifo_empty(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.pcfifofull(w_hssi_8g_rx_pcs_pcfifofull),
				.phystatus(w_hssi_8g_rx_pcs_phystatus),
				.pipe_data(w_hssi_8g_rx_pcs_pipe_data),
				.rd_enable_out_chnl_down(w_hssi_8g_rx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_rx_pcs_rd_enable_out_chnl_up),
				.rd_ptr1_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo),
				.rd_ptr2_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo),
				.rd_ptr_rx_phfifo(w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.reset_pc_ptrs_out_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down),
				.reset_pc_ptrs_out_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up),
				.rm_fifo_empty(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.rm_fifo_full(w_hssi_8g_rx_pcs_rm_fifo_full),
				.rx_blk_start(w_hssi_8g_rx_pcs_rx_blk_start),
				.rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.rx_data_valid(w_hssi_8g_rx_pcs_rx_data_valid),
				.rx_div_sync_out_chnl_down(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down),
				.rx_div_sync_out_chnl_up(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up),
				.rx_pipe_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.rx_pipe_soft_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rx_pma_clk_gen3(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_rcvd_clk_gen3(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_rstn_sync2wrfifo_8g(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.rx_sync_hdr(w_hssi_8g_rx_pcs_rx_sync_hdr),
				.rx_we_out_chnl_down(w_hssi_8g_rx_pcs_rx_we_out_chnl_down),
				.rx_we_out_chnl_up(w_hssi_8g_rx_pcs_rx_we_out_chnl_up),
				.rxstatus(w_hssi_8g_rx_pcs_rxstatus),
				.rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.word_align_boundary(w_hssi_8g_rx_pcs_word_align_boundary),
				.wr_clk_rx_phfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_rx_phfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_rx_rmfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_rx_rmfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_data_rx_phfifo(w_hssi_8g_rx_pcs_wr_data_rx_phfifo),
				.wr_data_rx_rmfifo(w_hssi_8g_rx_pcs_wr_data_rx_rmfifo),
				.wr_en_rx_phfifo(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_rx_rmfifo(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_rx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_rx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_rx_phfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo),
				.wr_ptr_rx_rmfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo),
				.wr_rst_n_rx_phfifo(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_rx_rmfifo(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				// INPUTS
				.a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bit_reversal_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.datain({w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0]}),
				.disable_pc_fifo_byte_serdes(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4]),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.eidleinfersel({w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0]}),
				.eios_detected_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.enable_comma_detect(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.gen3_clk_sel(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.hrd_rst(1'b0),
				.inferred_rxvalid_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.pc_fifo_rd_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.pc_fifo_wrdisable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.phystatus_int(w_hssi_pipe_gen1_2_phystatus),
				.phystatus_pcs_gen3(w_hssi_pipe_gen3_phystatus),
				.pipe_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.polarity_inversion(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.rd_data1_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0]}),
				.rd_data2_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0]}),
				.rd_data_rx_phfifo({w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[3]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[3]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.reset_pc_ptrs_asn(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5]),
				.reset_pc_ptrs_in_chnl_down(in_bond_pcs8g_in_bot[12]),
				.reset_pc_ptrs_in_chnl_up(in_bond_pcs8g_in_top[12]),
				.reset_ppm_cntrs_pcs_pma(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7]),
				.rm_fifo_read_enable(1'b0),
				.rm_fifo_write_enable(1'b0),
				.rx_blk_start_pcs_gen3({w_hssi_pipe_gen3_rx_blk_start[3], w_hssi_pipe_gen3_rx_blk_start[2], w_hssi_pipe_gen3_rx_blk_start[1], w_hssi_pipe_gen3_rx_blk_start[0]}),
				.rx_data_pcs_gen3({w_hssi_pipe_gen3_rxd_8gpcs_out[63], w_hssi_pipe_gen3_rxd_8gpcs_out[62], w_hssi_pipe_gen3_rxd_8gpcs_out[61], w_hssi_pipe_gen3_rxd_8gpcs_out[60], w_hssi_pipe_gen3_rxd_8gpcs_out[59], w_hssi_pipe_gen3_rxd_8gpcs_out[58], w_hssi_pipe_gen3_rxd_8gpcs_out[57], w_hssi_pipe_gen3_rxd_8gpcs_out[56], w_hssi_pipe_gen3_rxd_8gpcs_out[55], w_hssi_pipe_gen3_rxd_8gpcs_out[54], w_hssi_pipe_gen3_rxd_8gpcs_out[53], w_hssi_pipe_gen3_rxd_8gpcs_out[52], w_hssi_pipe_gen3_rxd_8gpcs_out[51], w_hssi_pipe_gen3_rxd_8gpcs_out[50], w_hssi_pipe_gen3_rxd_8gpcs_out[49], w_hssi_pipe_gen3_rxd_8gpcs_out[48], w_hssi_pipe_gen3_rxd_8gpcs_out[47], w_hssi_pipe_gen3_rxd_8gpcs_out[46], w_hssi_pipe_gen3_rxd_8gpcs_out[45], w_hssi_pipe_gen3_rxd_8gpcs_out[44], w_hssi_pipe_gen3_rxd_8gpcs_out[43], w_hssi_pipe_gen3_rxd_8gpcs_out[42], w_hssi_pipe_gen3_rxd_8gpcs_out[41], w_hssi_pipe_gen3_rxd_8gpcs_out[40], w_hssi_pipe_gen3_rxd_8gpcs_out[39], w_hssi_pipe_gen3_rxd_8gpcs_out[38], w_hssi_pipe_gen3_rxd_8gpcs_out[37], w_hssi_pipe_gen3_rxd_8gpcs_out[36], w_hssi_pipe_gen3_rxd_8gpcs_out[35], w_hssi_pipe_gen3_rxd_8gpcs_out[34], w_hssi_pipe_gen3_rxd_8gpcs_out[33], w_hssi_pipe_gen3_rxd_8gpcs_out[32], w_hssi_pipe_gen3_rxd_8gpcs_out[31], w_hssi_pipe_gen3_rxd_8gpcs_out[30], w_hssi_pipe_gen3_rxd_8gpcs_out[29], w_hssi_pipe_gen3_rxd_8gpcs_out[28], w_hssi_pipe_gen3_rxd_8gpcs_out[27], w_hssi_pipe_gen3_rxd_8gpcs_out[26], w_hssi_pipe_gen3_rxd_8gpcs_out[25], w_hssi_pipe_gen3_rxd_8gpcs_out[24], w_hssi_pipe_gen3_rxd_8gpcs_out[23], w_hssi_pipe_gen3_rxd_8gpcs_out[22], w_hssi_pipe_gen3_rxd_8gpcs_out[21], w_hssi_pipe_gen3_rxd_8gpcs_out[20], w_hssi_pipe_gen3_rxd_8gpcs_out[19], w_hssi_pipe_gen3_rxd_8gpcs_out[18], w_hssi_pipe_gen3_rxd_8gpcs_out[17], w_hssi_pipe_gen3_rxd_8gpcs_out[16], w_hssi_pipe_gen3_rxd_8gpcs_out[15], w_hssi_pipe_gen3_rxd_8gpcs_out[14], w_hssi_pipe_gen3_rxd_8gpcs_out[13], w_hssi_pipe_gen3_rxd_8gpcs_out[12], w_hssi_pipe_gen3_rxd_8gpcs_out[11], w_hssi_pipe_gen3_rxd_8gpcs_out[10], w_hssi_pipe_gen3_rxd_8gpcs_out[9], w_hssi_pipe_gen3_rxd_8gpcs_out[8], w_hssi_pipe_gen3_rxd_8gpcs_out[7], w_hssi_pipe_gen3_rxd_8gpcs_out[6], w_hssi_pipe_gen3_rxd_8gpcs_out[5], w_hssi_pipe_gen3_rxd_8gpcs_out[4], w_hssi_pipe_gen3_rxd_8gpcs_out[3], w_hssi_pipe_gen3_rxd_8gpcs_out[2], w_hssi_pipe_gen3_rxd_8gpcs_out[1], w_hssi_pipe_gen3_rxd_8gpcs_out[0]}),
				.rx_data_valid_pcs_gen3({w_hssi_pipe_gen3_rxdataskip[3], w_hssi_pipe_gen3_rxdataskip[2], w_hssi_pipe_gen3_rxdataskip[1], w_hssi_pipe_gen3_rxdataskip[0]}),
				.rx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[1], in_bond_pcs8g_in_bot[0]}),
				.rx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[1], in_bond_pcs8g_in_top[0]}),
				.rx_pcs_rst(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.rx_sync_hdr_pcs_gen3({w_hssi_pipe_gen3_rx_sync_hdr[1], w_hssi_pipe_gen3_rx_sync_hdr[0]}),
				.rx_we_in_chnl_down({in_bond_pcs8g_in_bot[5], in_bond_pcs8g_in_bot[4]}),
				.rx_we_in_chnl_up({in_bond_pcs8g_in_top[5], in_bond_pcs8g_in_top[4]}),
				.rxstatus_int({w_hssi_pipe_gen1_2_rxstatus[2], w_hssi_pipe_gen1_2_rxstatus[1], w_hssi_pipe_gen1_2_rxstatus[0]}),
				.rxstatus_pcs_gen3({w_hssi_pipe_gen3_rxstatus[2], w_hssi_pipe_gen3_rxstatus[1], w_hssi_pipe_gen3_rxstatus[0]}),
				.rxvalid_int(w_hssi_pipe_gen1_2_rxvalid),
				.rxvalid_pcs_gen3(w_hssi_pipe_gen3_rxvalid),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.sig_det_from_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_ctrlplane_testbus({w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0]}),
				.tx_div_sync({w_hssi_8g_tx_pcs_tx_div_sync[1], w_hssi_8g_tx_pcs_tx_div_sync[0]}),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.tx_testbus({w_hssi_8g_tx_pcs_tx_testbus[19], w_hssi_8g_tx_pcs_tx_testbus[18], w_hssi_8g_tx_pcs_tx_testbus[17], w_hssi_8g_tx_pcs_tx_testbus[16], w_hssi_8g_tx_pcs_tx_testbus[15], w_hssi_8g_tx_pcs_tx_testbus[14], w_hssi_8g_tx_pcs_tx_testbus[13], w_hssi_8g_tx_pcs_tx_testbus[12], w_hssi_8g_tx_pcs_tx_testbus[11], w_hssi_8g_tx_pcs_tx_testbus[10], w_hssi_8g_tx_pcs_tx_testbus[9], w_hssi_8g_tx_pcs_tx_testbus[8], w_hssi_8g_tx_pcs_tx_testbus[7], w_hssi_8g_tx_pcs_tx_testbus[6], w_hssi_8g_tx_pcs_tx_testbus[5], w_hssi_8g_tx_pcs_tx_testbus[4], w_hssi_8g_tx_pcs_tx_testbus[3], w_hssi_8g_tx_pcs_tx_testbus[2], w_hssi_8g_tx_pcs_tx_testbus[1], w_hssi_8g_tx_pcs_tx_testbus[0]}),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[2]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[2]),
				
				// UNUSED
				.byte_deserializer_pcs_clk_div_by_2_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_wire(),
				.byte_deserializer_pcs_clk_div_by_2_wire(),
				.byte_deserializer_pcs_clk_div_by_4_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_2_reg(),
				.byte_deserializer_pld_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_4_txclk_reg(),
				.pld_8g_a1a2_k1k2_flag_reg(),
				.pld_8g_a1a2_k1k2_flag_txclk_reg(),
				.pld_8g_a1a2_size_reg(),
				.pld_8g_a1a2_size_txclk_reg(),
				.pld_8g_bitloc_rev_en_reg(),
				.pld_8g_bitloc_rev_en_txclk_reg(),
				.pld_8g_byte_rev_en_reg(),
				.pld_8g_byte_rev_en_txclk_reg(),
				.pld_8g_elecidle_reg(),
				.pld_8g_empty_rmf_lowlatency_reg(),
				.pld_8g_empty_rmf_lowlatency_txclk_reg(),
				.pld_8g_empty_rmf_reg(),
				.pld_8g_empty_rmf_txclk_reg(),
				.pld_8g_empty_rx_fifo(),
				.pld_8g_empty_rx_reg(),
				.pld_8g_empty_rx_txclk_reg(),
				.pld_8g_encdt_reg(),
				.pld_8g_encdt_txclk_reg(),
				.pld_8g_full_rmf_reg(),
				.pld_8g_full_rmf_txclk_reg(),
				.pld_8g_full_rx_fifo(),
				.pld_8g_full_rx_reg(),
				.pld_8g_full_rx_txclk_reg(),
				.pld_8g_g3_rx_pld_rst_n_reg(),
				.pld_8g_g3_rx_pld_rst_n_txclk_reg(),
				.pld_8g_rxelecidle_txclk_reg(),
				.pld_8g_rxpolarity_reg(),
				.pld_8g_rxpolarity_txclk_reg(),
				.pld_8g_wa_boundary_reg(),
				.pld_8g_wrdisable_rx_reg(),
				.pld_8g_wrdisable_rx_txclk_reg(),
				.pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_rx_clk_out_8g_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_wire(),
				.pld_rx_control_8g_reg(),
				.pld_rx_control_8g_txclk_reg(),
				.pld_rx_data_8g_reg(),
				.pld_rx_data_8g_txclk_reg(),
				.pld_syncsm_en_reg(),
				.pld_syncsm_en_txclk_reg(),
				.rm_fifo_partial_empty(),
				.rm_fifo_partial_full(),
				.sta_rx_clk2_by2_1(),
				.sta_rx_clk2_by2_1_out(),
				.sta_rx_clk2_by2_2(),
				.sta_rx_clk2_by2_2_out(),
				.sta_rx_clk2_by4_1(),
				.sta_rx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_rx_pcs_a1a2k1k2flag[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_rx_pcs_chnl_test_bus_out[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_clock_to_pld = 1'b0;
				assign w_hssi_8g_rx_pcs_dataout[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_dis_pc_byte = 1'b0;
				assign w_hssi_8g_rx_pcs_eidle_detected = 1'b0;
				assign w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_pma_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_gen2ngen1 = 1'b0;
				assign w_hssi_8g_rx_pcs_parallel_rev_loopback[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_pc_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_pcfifofull = 1'b0;
				assign w_hssi_8g_rx_pcs_phystatus = 1'b0;
				assign w_hssi_8g_rx_pcs_pipe_data[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_full = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clkslip = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_data_valid[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pma_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rxstatus[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_rxvalid = 1'b0;
				assign w_hssi_8g_rx_pcs_signal_detect_out = 1'b0;
				assign w_hssi_8g_rx_pcs_word_align_boundary[4:0] = 5'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79:0] = 80'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31:0] = 32'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_rmfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_tx_pcs
			twentynm_hssi_8g_tx_pcs #(
				.auto_speed_nego_gen2(hssi_8g_tx_pcs_auto_speed_nego_gen2),
				.bit_reversal(hssi_8g_tx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_tx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_tx_pcs_bypass_pipeline_reg),
				.byte_serializer(hssi_8g_tx_pcs_byte_serializer),
				.clock_gate_bs_enc(hssi_8g_tx_pcs_clock_gate_bs_enc),
				.clock_gate_dw_fifowr(hssi_8g_tx_pcs_clock_gate_dw_fifowr),
				.clock_gate_fiford(hssi_8g_tx_pcs_clock_gate_fiford),
				.clock_gate_sw_fifowr(hssi_8g_tx_pcs_clock_gate_sw_fifowr),
				.clock_observation_in_pld_core(hssi_8g_tx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_tx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_tx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_tx_pcs_ctrl_plane_bonding_distribution),
				.data_selection_8b10b_encoder_input(hssi_8g_tx_pcs_data_selection_8b10b_encoder_input),
				.dynamic_clk_switch(hssi_8g_tx_pcs_dynamic_clk_switch),
				.eightb_tenb_disp_ctrl(hssi_8g_tx_pcs_eightb_tenb_disp_ctrl),
				.eightb_tenb_encoder(hssi_8g_tx_pcs_eightb_tenb_encoder),
				.force_echar(hssi_8g_tx_pcs_force_echar),
				.force_kchar(hssi_8g_tx_pcs_force_kchar),
				.gen3_tx_clk_sel(hssi_8g_tx_pcs_gen3_tx_clk_sel),
				.gen3_tx_pipe_clk_sel(hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel),
				.hip_mode(hssi_8g_tx_pcs_hip_mode),
				.pcs_bypass(hssi_8g_tx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_tx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_tx_pcs_phase_compensation_fifo),
				.phfifo_write_clk_sel(hssi_8g_tx_pcs_phfifo_write_clk_sel),
				.pma_dw(hssi_8g_tx_pcs_pma_dw),
				.prot_mode(hssi_8g_tx_pcs_prot_mode),
				.reconfig_settings(hssi_8g_tx_pcs_reconfig_settings),
				.refclk_b_clk_sel(hssi_8g_tx_pcs_refclk_b_clk_sel),
				.revloop_back_rm(hssi_8g_tx_pcs_revloop_back_rm),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_tx_pcs_sup_mode),
				.symbol_swap(hssi_8g_tx_pcs_symbol_swap),
				.tx_bitslip(hssi_8g_tx_pcs_tx_bitslip),
				.tx_compliance_controlled_disparity(hssi_8g_tx_pcs_tx_compliance_controlled_disparity),
				.tx_fast_pld_reg(hssi_8g_tx_pcs_tx_fast_pld_reg),
				.txclk_freerun(hssi_8g_tx_pcs_txclk_freerun),
				.txpcs_urst(hssi_8g_tx_pcs_txpcs_urst)
			) inst_twentynm_hssi_8g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_8g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_tx_pcs_blockselect),
				.clk_out(w_hssi_8g_tx_pcs_clk_out),
				.clk_out_gen3(w_hssi_8g_tx_pcs_clk_out_gen3),
				.dataout(w_hssi_8g_tx_pcs_dataout),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.fifo_select_out_chnl_down(w_hssi_8g_tx_pcs_fifo_select_out_chnl_down),
				.fifo_select_out_chnl_up(w_hssi_8g_tx_pcs_fifo_select_out_chnl_up),
				.g3_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.g3_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
				.non_gray_eidleinfersel(w_hssi_8g_tx_pcs_non_gray_eidleinfersel),
				.ph_fifo_overflow(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.ph_fifo_underflow(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.phfifo_txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.phfifo_txmargin(w_hssi_8g_tx_pcs_phfifo_txmargin),
				.phfifo_txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				.pipe_en_rev_parallel_lpbk_out(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.pipe_power_down_out(w_hssi_8g_tx_pcs_pipe_power_down_out),
				.pipe_tx_clk_out_gen3(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pmaif_asn_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.rd_enable_out_chnl_down(w_hssi_8g_tx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_tx_pcs_rd_enable_out_chnl_up),
				.rd_ptr_tx_phfifo(w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rxpolarity_int(w_hssi_8g_tx_pcs_rxpolarity_int),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.tx_blk_start_out(w_hssi_8g_tx_pcs_tx_blk_start_out),
				.tx_clk_out_8g_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.tx_ctrlplane_testbus(w_hssi_8g_tx_pcs_tx_ctrlplane_testbus),
				.tx_data_out(w_hssi_8g_tx_pcs_tx_data_out),
				.tx_data_valid_out(w_hssi_8g_tx_pcs_tx_data_valid_out),
				.tx_datak_out(w_hssi_8g_tx_pcs_tx_datak_out),
				.tx_detect_rxloopback_int(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.tx_div_sync(w_hssi_8g_tx_pcs_tx_div_sync),
				.tx_div_sync_out_chnl_down(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down),
				.tx_div_sync_out_chnl_up(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up),
				.tx_pipe_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.tx_pipe_electidle(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_soft_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.tx_sync_hdr_out(w_hssi_8g_tx_pcs_tx_sync_hdr_out),
				.tx_testbus(w_hssi_8g_tx_pcs_tx_testbus),
				.txcompliance_out(w_hssi_8g_tx_pcs_txcompliance_out),
				.txelecidle_out(w_hssi_8g_tx_pcs_txelecidle_out),
				.wr_clk_tx_phfifo_dw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_tx_phfifo_sw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_data_tx_phfifo(w_hssi_8g_tx_pcs_wr_data_tx_phfifo),
				.wr_en_tx_phfifo(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_tx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_tx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_tx_phfifo(w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo),
				.wr_rst_n_tx_phfifo(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bitslip_boundary_select({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0]}),
				.clk_sel_gen3(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.coreclk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.datain({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.detectrxloopin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidleinfersel({w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0]}),
				.en_rev_parallel_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.fifo_select_in_chnl_down({in_bond_pcs8g_in_bot[11], in_bond_pcs8g_in_bot[10]}),
				.fifo_select_in_chnl_up({in_bond_pcs8g_in_top[11], in_bond_pcs8g_in_top[10]}),
				.hrdrst(1'b0),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.ph_fifo_rd_disable(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.pipe_en_rev_parallel_lpbk_in(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.pipe_tx_deemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.pipe_tx_margin({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0]}),
				.powerdn({w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0]}),
				.rate_switch(w_hssi_8g_rx_pcs_gen2ngen1),
				.rd_data_tx_phfifo({w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[9]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[9]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.rev_parallel_lpbk_data({w_hssi_8g_rx_pcs_parallel_rev_loopback[19], w_hssi_8g_rx_pcs_parallel_rev_loopback[18], w_hssi_8g_rx_pcs_parallel_rev_loopback[17], w_hssi_8g_rx_pcs_parallel_rev_loopback[16], w_hssi_8g_rx_pcs_parallel_rev_loopback[15], w_hssi_8g_rx_pcs_parallel_rev_loopback[14], w_hssi_8g_rx_pcs_parallel_rev_loopback[13], w_hssi_8g_rx_pcs_parallel_rev_loopback[12], w_hssi_8g_rx_pcs_parallel_rev_loopback[11], w_hssi_8g_rx_pcs_parallel_rev_loopback[10], w_hssi_8g_rx_pcs_parallel_rev_loopback[9], w_hssi_8g_rx_pcs_parallel_rev_loopback[8], w_hssi_8g_rx_pcs_parallel_rev_loopback[7], w_hssi_8g_rx_pcs_parallel_rev_loopback[6], w_hssi_8g_rx_pcs_parallel_rev_loopback[5], w_hssi_8g_rx_pcs_parallel_rev_loopback[4], w_hssi_8g_rx_pcs_parallel_rev_loopback[3], w_hssi_8g_rx_pcs_parallel_rev_loopback[2], w_hssi_8g_rx_pcs_parallel_rev_loopback[1], w_hssi_8g_rx_pcs_parallel_rev_loopback[0]}),
				.rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.tx_blk_start({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0]}),
				.tx_data_valid({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0]}),
				.tx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[7], in_bond_pcs8g_in_bot[6]}),
				.tx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[7], in_bond_pcs8g_in_top[6]}),
				.tx_pcs_reset(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.tx_sync_hdr({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0]}),
				.txd_fast_reg({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0]}),
				.txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[8]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[8]),
				.wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				
				// UNUSED
				.byte_serializer_pcs_clk_div_by_2_reg(),
				.byte_serializer_pcs_clk_div_by_2_wire(),
				.byte_serializer_pcs_clk_div_by_4_reg(),
				.byte_serializer_pld_clk_div_by_2_reg(),
				.byte_serializer_pld_clk_div_by_4_reg(),
				.pld_8g_empty_tx_fifo(),
				.pld_8g_empty_tx_reg(),
				.pld_8g_full_tx_fifo(),
				.pld_8g_full_tx_reg(),
				.pld_8g_g3_tx_pld_rst_n_reg(),
				.pld_8g_rddisable_tx_reg(),
				.pld_8g_tx_boundary_sel_reg(),
				.pld_pcs_tx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_tx_clk_out_8g_wire(),
				.pld_tx_data_8g_fifo(),
				.pld_tx_data_lo_8g_reg(),
				.sta_tx_clk2_by2_1(),
				.sta_tx_clk2_by2_1_out(),
				.sta_tx_clk2_by4_1(),
				.sta_tx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_dataout[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_dyn_clk_switch_n = 1'b1;		// Override default tieoff
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_g3_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_overflow = 1'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_underflow = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txdeemph = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txmargin[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txswing = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_power_down_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_pmaif_asn_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_refclk_b = 1'b0;
				assign w_hssi_8g_tx_pcs_refclk_b_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_rxpolarity_int = 1'b0;
				assign w_hssi_8g_tx_pcs_soft_reset_wclk1_n = 1'b0;
				assign w_hssi_8g_tx_pcs_sw_fifo_wr_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_blk_start_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_tx_data_out[31:0] = 32'b0;
				assign w_hssi_8g_tx_pcs_tx_data_valid_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_datak_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_detect_rxloopback_int = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_electidle = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_sync_hdr_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_txcompliance_out = 1'b0;
				assign w_hssi_8g_tx_pcs_txelecidle_out = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63:0] = 64'b0;
				assign w_hssi_8g_tx_pcs_wr_en_tx_phfifo = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pcs_pma_interface
			twentynm_hssi_common_pcs_pma_interface #(
				.asn_clk_enable(hssi_common_pcs_pma_interface_asn_clk_enable),
				.asn_enable(hssi_common_pcs_pma_interface_asn_enable),
				.block_sel(hssi_common_pcs_pma_interface_block_sel),
				.bypass_early_eios(hssi_common_pcs_pma_interface_bypass_early_eios),
				.bypass_pcie_switch(hssi_common_pcs_pma_interface_bypass_pcie_switch),
				.bypass_pma_ltr(hssi_common_pcs_pma_interface_bypass_pma_ltr),
				.bypass_pma_sw_done(hssi_common_pcs_pma_interface_bypass_pma_sw_done),
				.bypass_ppm_lock(hssi_common_pcs_pma_interface_bypass_ppm_lock),
				.bypass_send_syncp_fbkp(hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp),
				.bypass_txdetectrx(hssi_common_pcs_pma_interface_bypass_txdetectrx),
				.cdr_control(hssi_common_pcs_pma_interface_cdr_control),
				.cid_enable(hssi_common_pcs_pma_interface_cid_enable),
				.cp_cons_sel(hssi_common_pcs_pma_interface_cp_cons_sel),
				.cp_dwn_mstr(hssi_common_pcs_pma_interface_cp_dwn_mstr),
				.cp_up_mstr(hssi_common_pcs_pma_interface_cp_up_mstr),
				.ctrl_plane_bonding(hssi_common_pcs_pma_interface_ctrl_plane_bonding),
				.data_mask_count(hssi_common_pcs_pma_interface_data_mask_count),
				.data_mask_count_multi(hssi_common_pcs_pma_interface_data_mask_count_multi),
				.dft_observation_clock_selection(hssi_common_pcs_pma_interface_dft_observation_clock_selection),
				.early_eios_counter(hssi_common_pcs_pma_interface_early_eios_counter),
				.force_freqdet(hssi_common_pcs_pma_interface_force_freqdet),
				.free_run_clk_enable(hssi_common_pcs_pma_interface_free_run_clk_enable),
				.ignore_sigdet_g23(hssi_common_pcs_pma_interface_ignore_sigdet_g23),
				.pc_en_counter(hssi_common_pcs_pma_interface_pc_en_counter),
				.pc_rst_counter(hssi_common_pcs_pma_interface_pc_rst_counter),
				.pcie_hip_mode(hssi_common_pcs_pma_interface_pcie_hip_mode),
				.ph_fifo_reg_mode(hssi_common_pcs_pma_interface_ph_fifo_reg_mode),
				.phfifo_flush_wait(hssi_common_pcs_pma_interface_phfifo_flush_wait),
				.pipe_if_g3pcs(hssi_common_pcs_pma_interface_pipe_if_g3pcs),
				.pma_done_counter(hssi_common_pcs_pma_interface_pma_done_counter),
				.pma_if_dft_en(hssi_common_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_common_pcs_pma_interface_pma_if_dft_val),
				.ppm_cnt_rst(hssi_common_pcs_pma_interface_ppm_cnt_rst),
				.ppm_deassert_early(hssi_common_pcs_pma_interface_ppm_deassert_early),
				.ppm_det_buckets(hssi_common_pcs_pma_interface_ppm_det_buckets),
				.ppm_gen1_2_cnt(hssi_common_pcs_pma_interface_ppm_gen1_2_cnt),
				.ppm_post_eidle_delay(hssi_common_pcs_pma_interface_ppm_post_eidle_delay),
				.ppmsel(hssi_common_pcs_pma_interface_ppmsel),
				.prot_mode(hssi_common_pcs_pma_interface_prot_mode),
				.reconfig_settings(hssi_common_pcs_pma_interface_reconfig_settings),
				.rxvalid_mask(hssi_common_pcs_pma_interface_rxvalid_mask),
				.sigdet_wait_counter(hssi_common_pcs_pma_interface_sigdet_wait_counter),
				.sigdet_wait_counter_multi(hssi_common_pcs_pma_interface_sigdet_wait_counter_multi),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sim_mode(hssi_common_pcs_pma_interface_sim_mode),
				.spd_chg_rst_wait_cnt_en(hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en),
				.sup_mode(hssi_common_pcs_pma_interface_sup_mode),
				.testout_sel(hssi_common_pcs_pma_interface_testout_sel),
				.wait_clk_on_off_timer(hssi_common_pcs_pma_interface_wait_clk_on_off_timer),
				.wait_pipe_synchronizing(hssi_common_pcs_pma_interface_wait_pipe_synchronizing),
				.wait_send_syncp_fbkp(hssi_common_pcs_pma_interface_wait_send_syncp_fbkp)
			) inst_twentynm_hssi_common_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_common_pcs_pma_interface_blockselect),
				.int_pmaif_8g_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in),
				.int_pmaif_8g_eios_detected(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.int_pmaif_8g_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.int_pmaif_8g_power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.int_pmaif_g3_pcs_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in),
				.int_pmaif_pldif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pmaif_pldif_pcie_sw_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done),
				.int_pmaif_pldif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pmaif_pldif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pmaif_pldif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pmaif_pldif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pmaif_pldif_pma_reserved_in(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in),
				.int_pmaif_pldif_test_out(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out),
				.int_pmaif_pldif_testbus(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus),
				.pma_adapt_start(w_hssi_common_pcs_pma_interface_pma_adapt_start),
				.pma_atpg_los_en_n(w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n),
				.pma_csr_test_dis(w_hssi_common_pcs_pma_interface_pma_csr_test_dis),
				.pma_current_coeff(w_hssi_common_pcs_pma_interface_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_common_pcs_pma_interface_pma_current_rxpreset),
				.pma_early_eios(w_hssi_common_pcs_pma_interface_pma_early_eios),
				.pma_interface_select(w_hssi_common_pcs_pma_interface_pma_interface_select),
				.pma_ltd_b(w_hssi_common_pcs_pma_interface_pma_ltd_b),
				.pma_ltr(w_hssi_common_pcs_pma_interface_pma_ltr),
				.pma_nfrzdrv(w_hssi_common_pcs_pma_interface_pma_nfrzdrv),
				.pma_nrpi_freeze(w_hssi_common_pcs_pma_interface_pma_nrpi_freeze),
				.pma_pcie_switch(w_hssi_common_pcs_pma_interface_pma_pcie_switch),
				.pma_ppm_lock(w_hssi_common_pcs_pma_interface_pma_ppm_lock),
				.pma_reserved_out(w_hssi_common_pcs_pma_interface_pma_reserved_out),
				.pma_rs_lpbk_b(w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b),
				.pma_rx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup),
				.pma_scan_mode_n(w_hssi_common_pcs_pma_interface_pma_scan_mode_n),
				.pma_scan_shift_n(w_hssi_common_pcs_pma_interface_pma_scan_shift_n),
				.pma_tx_bitslip(w_hssi_common_pcs_pma_interface_pma_tx_bitslip),
				.pma_tx_bonding_rstb(w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb),
				.pma_tx_qpi_pulldn(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn),
				.pma_tx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup),
				.pma_tx_txdetectrx(w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx),
				.pmaif_bundling_out_down(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down),
				.pmaif_bundling_out_up(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_8g_current_coeff({w_hssi_pipe_gen1_2_current_coeff[17], w_hssi_pipe_gen1_2_current_coeff[16], w_hssi_pipe_gen1_2_current_coeff[15], w_hssi_pipe_gen1_2_current_coeff[14], w_hssi_pipe_gen1_2_current_coeff[13], w_hssi_pipe_gen1_2_current_coeff[12], w_hssi_pipe_gen1_2_current_coeff[11], w_hssi_pipe_gen1_2_current_coeff[10], w_hssi_pipe_gen1_2_current_coeff[9], w_hssi_pipe_gen1_2_current_coeff[8], w_hssi_pipe_gen1_2_current_coeff[7], w_hssi_pipe_gen1_2_current_coeff[6], w_hssi_pipe_gen1_2_current_coeff[5], w_hssi_pipe_gen1_2_current_coeff[4], w_hssi_pipe_gen1_2_current_coeff[3], w_hssi_pipe_gen1_2_current_coeff[2], w_hssi_pipe_gen1_2_current_coeff[1], w_hssi_pipe_gen1_2_current_coeff[0]}),
				.int_pmaif_8g_eios_det({w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0]}),
				.int_pmaif_8g_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.int_pmaif_8g_rev_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.int_pmaif_8g_tx_clk_out_gen3(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.int_pmaif_8g_txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				.int_pmaif_g3_eios_det({w_hssi_gen3_rx_pcs_ei_det_int, w_hssi_gen3_rx_pcs_ei_partial_det_int, w_hssi_gen3_rx_pcs_i_det_int}),
				.int_pmaif_g3_pma_current_coeff({w_hssi_pipe_gen3_pma_current_coeff[17], w_hssi_pipe_gen3_pma_current_coeff[16], w_hssi_pipe_gen3_pma_current_coeff[15], w_hssi_pipe_gen3_pma_current_coeff[14], w_hssi_pipe_gen3_pma_current_coeff[13], w_hssi_pipe_gen3_pma_current_coeff[12], w_hssi_pipe_gen3_pma_current_coeff[11], w_hssi_pipe_gen3_pma_current_coeff[10], w_hssi_pipe_gen3_pma_current_coeff[9], w_hssi_pipe_gen3_pma_current_coeff[8], w_hssi_pipe_gen3_pma_current_coeff[7], w_hssi_pipe_gen3_pma_current_coeff[6], w_hssi_pipe_gen3_pma_current_coeff[5], w_hssi_pipe_gen3_pma_current_coeff[4], w_hssi_pipe_gen3_pma_current_coeff[3], w_hssi_pipe_gen3_pma_current_coeff[2], w_hssi_pipe_gen3_pma_current_coeff[1], w_hssi_pipe_gen3_pma_current_coeff[0]}),
				.int_pmaif_g3_pma_current_rxpreset({w_hssi_pipe_gen3_pma_current_rxpreset[2], w_hssi_pipe_gen3_pma_current_rxpreset[1], w_hssi_pipe_gen3_pma_current_rxpreset[0]}),
				.int_pmaif_g3_pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.int_pmaif_g3_rev_lpbk(w_hssi_pipe_gen3_rev_lpbk_int),
				.int_pmaif_pldif_8g_tx_pld_rstn(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pmaif_pldif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pmaif_pldif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pmaif_pldif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pmaif_pldif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pmaif_pldif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pmaif_pldif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pmaif_pldif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pmaif_pldif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pmaif_pldif_pcie_switch({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0]}),
				.int_pmaif_pldif_pma_reserved_out({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0]}),
				.int_pmaif_pldif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pmaif_pldif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pmaif_pldif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pmaif_pldif_rate({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0]}),
				.int_pmaif_pldif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pmaif_pldif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pmaif_pldif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.int_pmaif_pldif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pmaif_pldif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pmaif_pldif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pmaif_pldif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pmaif_pldif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pmaif_pldif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.int_tx_dft_obsrv_clk({w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0]}),
				.iocsr_clk(in_iocsr_clk),
				.iocsr_config({in_iocsr_config[5], in_iocsr_config[4], in_iocsr_config[3], in_iocsr_config[2], in_iocsr_config[1], in_iocsr_config[0]}),
				.iocsr_rdy(in_iocsr_rdy),
				.iocsr_rdy_dly(in_iocsr_rdy_dly),
				.pma_adapt_done(in_pma_adapt_done),
				.pma_clklow(in_pma_clklow),
				.pma_fref(in_pma_fref),
				.pma_hclk(in_pma_hclk),
				.pma_pcie_sw_done({in_pma_pcie_sw_done[1], in_pma_pcie_sw_done[0]}),
				.pma_pfdmode_lock(in_pma_pfdmode_lock),
				.pma_reserved_in({in_pma_reserved_in[4], in_pma_reserved_in[3], in_pma_reserved_in[2], in_pma_reserved_in[1], in_pma_reserved_in[0]}),
				.pma_signal_det(in_pma_signal_det),
				.pma_testbus({in_pma_testbus[7], in_pma_testbus[6], in_pma_testbus[5], in_pma_testbus[4], in_pma_testbus[3], in_pma_testbus[2], in_pma_testbus[1], in_pma_testbus[0]}),
				.pmaif_bundling_in_down({in_bond_pmaif_in_bot[11], in_bond_pmaif_in_bot[10], in_bond_pmaif_in_bot[9], in_bond_pmaif_in_bot[8], in_bond_pmaif_in_bot[7], in_bond_pmaif_in_bot[6], in_bond_pmaif_in_bot[5], in_bond_pmaif_in_bot[4], in_bond_pmaif_in_bot[3], in_bond_pmaif_in_bot[2], in_bond_pmaif_in_bot[1], in_bond_pmaif_in_bot[0]}),
				.pmaif_bundling_in_up({in_bond_pmaif_in_top[11], in_bond_pmaif_in_top[10], in_bond_pmaif_in_top[9], in_bond_pmaif_in_top[8], in_bond_pmaif_in_top[7], in_bond_pmaif_in_top[6], in_bond_pmaif_in_top[5], in_bond_pmaif_in_top[4], in_bond_pmaif_in_top[3], in_bond_pmaif_in_top[2], in_bond_pmaif_in_top[1], in_bond_pmaif_in_top[0]}),
				.rx_pmaif_test_out({w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0]}),
				.rx_prbs_ver_test({w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0]}),
				.tx_prbs_gen_test({w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0]}),
				.uhsif_test_out_1({w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0]}),
				.uhsif_test_out_2({w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0]}),
				.uhsif_test_out_3({w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0]}),
				
				// UNUSED
				.int_pmaif_avmm_iocsr_clk(),
				.int_pmaif_avmm_iocsr_config(),
				.int_pmaif_avmm_iocsr_rdy(),
				.int_pmaif_avmm_iocsr_rdy_dly(),
				.int_pmaif_pldif_interface_select(),
				.pma_tx_pma_syncp(),
				.sta_pma_hclk_by2()
			);
		end // if generate
		else begin
				assign w_hssi_common_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19:0] = 20'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_pma_adapt_start = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_csr_test_dis = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pcs_pma_interface_pma_early_eios = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_interface_select[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltd_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltr = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nfrzdrv = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nrpi_freeze = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ppm_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_tx_bitslip = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx = in_pld_pma_txdetectrx;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11:0] = 12'b0;
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11:0] = 12'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pld_pcs_interface
			twentynm_hssi_common_pld_pcs_interface #(
				.dft_clk_out_en(hssi_common_pld_pcs_interface_dft_clk_out_en),
				.dft_clk_out_sel(hssi_common_pld_pcs_interface_dft_clk_out_sel),
				.hrdrstctrl_en(hssi_common_pld_pcs_interface_hrdrstctrl_en),
				.pcs_testbus_block_sel(hssi_common_pld_pcs_interface_pcs_testbus_block_sel),
				.reconfig_settings(hssi_common_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm5" )       //PARAM_HIDE
			) inst_twentynm_hssi_common_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_common_pld_pcs_interface_blockselect),
				.hip_cmn_clk(w_hssi_common_pld_pcs_interface_hip_cmn_clk),
				.hip_cmn_ctrl(w_hssi_common_pld_pcs_interface_hip_cmn_ctrl),
				.hip_iocsr_rdy(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy),
				.hip_iocsr_rdy_dly(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly),
				.hip_nfrzdrv(w_hssi_common_pld_pcs_interface_hip_nfrzdrv),
				.hip_npor(w_hssi_common_pld_pcs_interface_hip_npor),
				.hip_usermode(w_hssi_common_pld_pcs_interface_hip_usermode),
				.int_pldif_10g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.int_pldif_10g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.int_pldif_8g_eidleinfersel(w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel),
				.int_pldif_8g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.int_pldif_8g_refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.int_pldif_8g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.int_pldif_g3_current_coeff(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff),
				.int_pldif_g3_current_rxpreset(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset),
				.int_pldif_krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.int_pldif_krfec_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.int_pldif_krfec_scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				.int_pldif_mem_atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.int_pldif_mem_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.int_pldif_pmaif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pldif_pmaif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pldif_pmaif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pldif_pmaif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pldif_pmaif_eye_monitor(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor),
				.int_pldif_pmaif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pldif_pmaif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pldif_pmaif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pldif_pmaif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pldif_pmaif_pcie_switch(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch),
				.int_pldif_pmaif_pma_reserved_out(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out),
				.int_pldif_pmaif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pldif_pmaif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pldif_pmaif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pldif_pmaif_rate(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate),
				.int_pldif_pmaif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pldif_pmaif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pldif_pmaif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pldif_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_pldif_pmaif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pldif_pmaif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pldif_pmaif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pldif_pmaif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pldif_pmaif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pldif_pmaif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pldif_pmaif_uhsif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.pld_pma_adapt_done(w_hssi_common_pld_pcs_interface_pld_pma_adapt_done),
				.pld_pma_clklow(w_hssi_common_pld_pcs_interface_pld_pma_clklow),
				.pld_pma_fref(w_hssi_common_pld_pcs_interface_pld_pma_fref),
				.pld_pma_hclk(w_hssi_common_pld_pcs_interface_pld_pma_hclk),
				.pld_pma_pcie_sw_done(w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done),
				.pld_pma_pfdmode_lock(w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock),
				.pld_pma_reserved_in(w_hssi_common_pld_pcs_interface_pld_pma_reserved_in),
				.pld_pma_rx_detect_valid(w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid),
				.pld_pma_rx_found(w_hssi_common_pld_pcs_interface_pld_pma_rx_found),
				.pld_pma_rxpll_lock(w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock),
				.pld_pma_testbus(w_hssi_common_pld_pcs_interface_pld_pma_testbus),
				.pld_pmaif_mask_tx_pll(w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll),
				.pld_reserved_out(w_hssi_common_pld_pcs_interface_pld_reserved_out),
				.pld_test_data(w_hssi_common_pld_pcs_interface_pld_test_data),
				.pld_uhsif_lock(w_hssi_common_pld_pcs_interface_pld_uhsif_lock),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.int_pldif_10g_test_data({w_hssi_10g_tx_pcs_tx_test_data[19], w_hssi_10g_tx_pcs_tx_test_data[18], w_hssi_10g_tx_pcs_tx_test_data[17], w_hssi_10g_tx_pcs_tx_test_data[16], w_hssi_10g_tx_pcs_tx_test_data[15], w_hssi_10g_tx_pcs_tx_test_data[14], w_hssi_10g_tx_pcs_tx_test_data[13], w_hssi_10g_tx_pcs_tx_test_data[12], w_hssi_10g_tx_pcs_tx_test_data[11], w_hssi_10g_tx_pcs_tx_test_data[10], w_hssi_10g_tx_pcs_tx_test_data[9], w_hssi_10g_tx_pcs_tx_test_data[8], w_hssi_10g_tx_pcs_tx_test_data[7], w_hssi_10g_tx_pcs_tx_test_data[6], w_hssi_10g_tx_pcs_tx_test_data[5], w_hssi_10g_tx_pcs_tx_test_data[4], w_hssi_10g_tx_pcs_tx_test_data[3], w_hssi_10g_tx_pcs_tx_test_data[2], w_hssi_10g_tx_pcs_tx_test_data[1], w_hssi_10g_tx_pcs_tx_test_data[0]}),
				.int_pldif_10g_tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.int_pldif_8g_chnl_test_bus_out({w_hssi_8g_rx_pcs_chnl_test_bus_out[19], w_hssi_8g_rx_pcs_chnl_test_bus_out[18], w_hssi_8g_rx_pcs_chnl_test_bus_out[17], w_hssi_8g_rx_pcs_chnl_test_bus_out[16], w_hssi_8g_rx_pcs_chnl_test_bus_out[15], w_hssi_8g_rx_pcs_chnl_test_bus_out[14], w_hssi_8g_rx_pcs_chnl_test_bus_out[13], w_hssi_8g_rx_pcs_chnl_test_bus_out[12], w_hssi_8g_rx_pcs_chnl_test_bus_out[11], w_hssi_8g_rx_pcs_chnl_test_bus_out[10], w_hssi_8g_rx_pcs_chnl_test_bus_out[9], w_hssi_8g_rx_pcs_chnl_test_bus_out[8], w_hssi_8g_rx_pcs_chnl_test_bus_out[7], w_hssi_8g_rx_pcs_chnl_test_bus_out[6], w_hssi_8g_rx_pcs_chnl_test_bus_out[5], w_hssi_8g_rx_pcs_chnl_test_bus_out[4], w_hssi_8g_rx_pcs_chnl_test_bus_out[3], w_hssi_8g_rx_pcs_chnl_test_bus_out[2], w_hssi_8g_rx_pcs_chnl_test_bus_out[1], w_hssi_8g_rx_pcs_chnl_test_bus_out[0]}),
				.int_pldif_8g_rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.int_pldif_8g_tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.int_pldif_g3_test_out({w_hssi_pipe_gen3_test_out[19], w_hssi_pipe_gen3_test_out[18], w_hssi_pipe_gen3_test_out[17], w_hssi_pipe_gen3_test_out[16], w_hssi_pipe_gen3_test_out[15], w_hssi_pipe_gen3_test_out[14], w_hssi_pipe_gen3_test_out[13], w_hssi_pipe_gen3_test_out[12], w_hssi_pipe_gen3_test_out[11], w_hssi_pipe_gen3_test_out[10], w_hssi_pipe_gen3_test_out[9], w_hssi_pipe_gen3_test_out[8], w_hssi_pipe_gen3_test_out[7], w_hssi_pipe_gen3_test_out[6], w_hssi_pipe_gen3_test_out[5], w_hssi_pipe_gen3_test_out[4], w_hssi_pipe_gen3_test_out[3], w_hssi_pipe_gen3_test_out[2], w_hssi_pipe_gen3_test_out[1], w_hssi_pipe_gen3_test_out[0]}),
				.int_pldif_krfec_test_data({w_hssi_krfec_tx_pcs_tx_test_data[19], w_hssi_krfec_tx_pcs_tx_test_data[18], w_hssi_krfec_tx_pcs_tx_test_data[17], w_hssi_krfec_tx_pcs_tx_test_data[16], w_hssi_krfec_tx_pcs_tx_test_data[15], w_hssi_krfec_tx_pcs_tx_test_data[14], w_hssi_krfec_tx_pcs_tx_test_data[13], w_hssi_krfec_tx_pcs_tx_test_data[12], w_hssi_krfec_tx_pcs_tx_test_data[11], w_hssi_krfec_tx_pcs_tx_test_data[10], w_hssi_krfec_tx_pcs_tx_test_data[9], w_hssi_krfec_tx_pcs_tx_test_data[8], w_hssi_krfec_tx_pcs_tx_test_data[7], w_hssi_krfec_tx_pcs_tx_test_data[6], w_hssi_krfec_tx_pcs_tx_test_data[5], w_hssi_krfec_tx_pcs_tx_test_data[4], w_hssi_krfec_tx_pcs_tx_test_data[3], w_hssi_krfec_tx_pcs_tx_test_data[2], w_hssi_krfec_tx_pcs_tx_test_data[1], w_hssi_krfec_tx_pcs_tx_test_data[0]}),
				.int_pldif_pmaif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pldif_pmaif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pldif_pmaif_pcie_sw_done({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0]}),
				.int_pldif_pmaif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pldif_pmaif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pldif_pmaif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pldif_pmaif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pldif_pmaif_pma_reserved_in({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0]}),
				.int_pldif_pmaif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pldif_pmaif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_test_out({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0]}),
				.int_pldif_pmaif_testbus({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0]}),
				.int_pldif_pmaif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.pld_8g_eidleinfersel({in_pld_8g_eidleinfersel[2], in_pld_8g_eidleinfersel[1], in_pld_8g_eidleinfersel[0]}),
				.pld_8g_refclk_dig2(in_pld_8g_refclk_dig2),
				.pld_atpg_los_en_n(in_pld_atpg_los_en_n),
				.pld_g3_current_coeff({in_pld_g3_current_coeff[17], in_pld_g3_current_coeff[16], in_pld_g3_current_coeff[15], in_pld_g3_current_coeff[14], in_pld_g3_current_coeff[13], in_pld_g3_current_coeff[12], in_pld_g3_current_coeff[11], in_pld_g3_current_coeff[10], in_pld_g3_current_coeff[9], in_pld_g3_current_coeff[8], in_pld_g3_current_coeff[7], in_pld_g3_current_coeff[6], in_pld_g3_current_coeff[5], in_pld_g3_current_coeff[4], in_pld_g3_current_coeff[3], in_pld_g3_current_coeff[2], in_pld_g3_current_coeff[1], in_pld_g3_current_coeff[0]}),
				.pld_g3_current_rxpreset({in_pld_g3_current_rxpreset[2], in_pld_g3_current_rxpreset[1], in_pld_g3_current_rxpreset[0]}),
				.pld_ltr(in_pld_ltr),
				.pld_mem_krfec_atpg_rst_n(in_pld_mem_krfec_atpg_rst_n),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pcs_refclk_dig(in_pld_pcs_refclk_dig),
				.pld_pma_adapt_start(in_pld_pma_adapt_start),
				.pld_pma_csr_test_dis(in_pld_pma_csr_test_dis),
				.pld_pma_early_eios(in_pld_pma_early_eios),
				.pld_pma_eye_monitor({in_pld_pma_eye_monitor[5], in_pld_pma_eye_monitor[4], in_pld_pma_eye_monitor[3], in_pld_pma_eye_monitor[2], in_pld_pma_eye_monitor[1], in_pld_pma_eye_monitor[0]}),
				.pld_pma_ltd_b(in_pld_pma_ltd_b),
				.pld_pma_nrpi_freeze(in_pld_pma_nrpi_freeze),
				.pld_pma_pcie_switch({in_pld_pma_pcie_switch[1], in_pld_pma_pcie_switch[0]}),
				.pld_pma_ppm_lock(in_pld_pma_ppm_lock),
				.pld_pma_reserved_out({in_pld_pma_reserved_out[4], in_pld_pma_reserved_out[3], in_pld_pma_reserved_out[2], in_pld_pma_reserved_out[1], in_pld_pma_reserved_out[0]}),
				.pld_pma_rs_lpbk_b(in_pld_pma_rs_lpbk_b),
				.pld_pma_rx_qpi_pullup(in_pld_pma_rx_qpi_pullup),
				.pld_pma_tx_bitslip(in_pld_pma_tx_bitslip),
				.pld_pma_tx_bonding_rstb(in_pld_pma_tx_bonding_rstb),
				.pld_pma_tx_qpi_pulldn(in_pld_pma_tx_qpi_pulldn),
				.pld_pma_tx_qpi_pullup(in_pld_pma_tx_qpi_pullup),
				.pld_pma_txdetectrx(in_pld_pma_txdetectrx),
				.pld_rate({in_pld_rate[1], in_pld_rate[0]}),
				.pld_reserved_in({in_pld_reserved_in[9], in_pld_reserved_in[8], in_pld_reserved_in[7], in_pld_reserved_in[6], in_pld_reserved_in[5], in_pld_reserved_in[4], in_pld_reserved_in[3], in_pld_reserved_in[2], in_pld_reserved_in[1], in_pld_reserved_in[0]}),
				.pld_scan_mode_n(in_pld_scan_mode_n),
				.pld_scan_shift_n(in_pld_scan_shift_n),
				
				// UNUSED
				.int_pldif_8g_ltr(),
				.int_pldif_avmm_pld_avmm1_request(),
				.int_pldif_avmm_pld_avmm2_request(),
				.int_pldif_avmm_refclk_dig_en(),
				.int_pldif_g3_scan_mode_n(),
				.pld_8g_eidleinfersel_fifo(),
				.pld_8g_eidleinfersel_reg(),
				.pld_partial_reconfig_fifo(),
				.pld_partial_reconfig_rx_div_by_2_rxclk_wire(),
				.pld_partial_reconfig_rx_div_by_2_txclk_wire(),
				.pld_partial_reconfig_rxclk_reg(),
				.pld_partial_reconfig_tx_div_by_2_wire(),
				.pld_partial_reconfig_txclk_reg(),
				.pld_rate_reg(),
				.pld_test_data_reg()
			);
		end // if generate
		else begin
				assign w_hssi_common_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_clk[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_npor = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_usermode = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2 = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_adapt_done = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_clklow = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_fref = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_hclk = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_found = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_testbus[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_reserved_out[9:0] = 10'b0;
				assign w_hssi_common_pld_pcs_interface_pld_test_data[19:0] = 20'b0;
				assign w_hssi_common_pld_pcs_interface_pld_uhsif_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_scan_mode_n = 1'b1;		// Override default tieoff
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_rx_pcs
			twentynm_hssi_fifo_rx_pcs #(
				.double_read_mode(hssi_fifo_rx_pcs_double_read_mode),
				.prot_mode(hssi_fifo_rx_pcs_prot_mode),
				.silicon_rev( "20nm5" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_rx_pcs_blockselect),
				.data_out2_10g(w_hssi_fifo_rx_pcs_data_out2_10g),
				.data_out2_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp),
				.data_out_10g(w_hssi_fifo_rx_pcs_data_out_10g),
				.data_out_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out_8g_clock_comp),
				.data_out_8g_phase_comp(w_hssi_fifo_rx_pcs_data_out_8g_phase_comp),
				.data_out_gen3(w_hssi_fifo_rx_pcs_data_out_gen3),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_data[73], w_hssi_10g_rx_pcs_rx_fifo_wr_data[72], w_hssi_10g_rx_pcs_rx_fifo_wr_data[71], w_hssi_10g_rx_pcs_rx_fifo_wr_data[70], w_hssi_10g_rx_pcs_rx_fifo_wr_data[69], w_hssi_10g_rx_pcs_rx_fifo_wr_data[68], w_hssi_10g_rx_pcs_rx_fifo_wr_data[67], w_hssi_10g_rx_pcs_rx_fifo_wr_data[66], w_hssi_10g_rx_pcs_rx_fifo_wr_data[65], w_hssi_10g_rx_pcs_rx_fifo_wr_data[64], w_hssi_10g_rx_pcs_rx_fifo_wr_data[63], w_hssi_10g_rx_pcs_rx_fifo_wr_data[62], w_hssi_10g_rx_pcs_rx_fifo_wr_data[61], w_hssi_10g_rx_pcs_rx_fifo_wr_data[60], w_hssi_10g_rx_pcs_rx_fifo_wr_data[59], w_hssi_10g_rx_pcs_rx_fifo_wr_data[58], w_hssi_10g_rx_pcs_rx_fifo_wr_data[57], w_hssi_10g_rx_pcs_rx_fifo_wr_data[56], w_hssi_10g_rx_pcs_rx_fifo_wr_data[55], w_hssi_10g_rx_pcs_rx_fifo_wr_data[54], w_hssi_10g_rx_pcs_rx_fifo_wr_data[53], w_hssi_10g_rx_pcs_rx_fifo_wr_data[52], w_hssi_10g_rx_pcs_rx_fifo_wr_data[51], w_hssi_10g_rx_pcs_rx_fifo_wr_data[50], w_hssi_10g_rx_pcs_rx_fifo_wr_data[49], w_hssi_10g_rx_pcs_rx_fifo_wr_data[48], w_hssi_10g_rx_pcs_rx_fifo_wr_data[47], w_hssi_10g_rx_pcs_rx_fifo_wr_data[46], w_hssi_10g_rx_pcs_rx_fifo_wr_data[45], w_hssi_10g_rx_pcs_rx_fifo_wr_data[44], w_hssi_10g_rx_pcs_rx_fifo_wr_data[43], w_hssi_10g_rx_pcs_rx_fifo_wr_data[42], w_hssi_10g_rx_pcs_rx_fifo_wr_data[41], w_hssi_10g_rx_pcs_rx_fifo_wr_data[40], w_hssi_10g_rx_pcs_rx_fifo_wr_data[39], w_hssi_10g_rx_pcs_rx_fifo_wr_data[38], w_hssi_10g_rx_pcs_rx_fifo_wr_data[37], w_hssi_10g_rx_pcs_rx_fifo_wr_data[36], w_hssi_10g_rx_pcs_rx_fifo_wr_data[35], w_hssi_10g_rx_pcs_rx_fifo_wr_data[34], w_hssi_10g_rx_pcs_rx_fifo_wr_data[33], w_hssi_10g_rx_pcs_rx_fifo_wr_data[32], w_hssi_10g_rx_pcs_rx_fifo_wr_data[31], w_hssi_10g_rx_pcs_rx_fifo_wr_data[30], w_hssi_10g_rx_pcs_rx_fifo_wr_data[29], w_hssi_10g_rx_pcs_rx_fifo_wr_data[28], w_hssi_10g_rx_pcs_rx_fifo_wr_data[27], w_hssi_10g_rx_pcs_rx_fifo_wr_data[26], w_hssi_10g_rx_pcs_rx_fifo_wr_data[25], w_hssi_10g_rx_pcs_rx_fifo_wr_data[24], w_hssi_10g_rx_pcs_rx_fifo_wr_data[23], w_hssi_10g_rx_pcs_rx_fifo_wr_data[22], w_hssi_10g_rx_pcs_rx_fifo_wr_data[21], w_hssi_10g_rx_pcs_rx_fifo_wr_data[20], w_hssi_10g_rx_pcs_rx_fifo_wr_data[19], w_hssi_10g_rx_pcs_rx_fifo_wr_data[18], w_hssi_10g_rx_pcs_rx_fifo_wr_data[17], w_hssi_10g_rx_pcs_rx_fifo_wr_data[16], w_hssi_10g_rx_pcs_rx_fifo_wr_data[15], w_hssi_10g_rx_pcs_rx_fifo_wr_data[14], w_hssi_10g_rx_pcs_rx_fifo_wr_data[13], w_hssi_10g_rx_pcs_rx_fifo_wr_data[12], w_hssi_10g_rx_pcs_rx_fifo_wr_data[11], w_hssi_10g_rx_pcs_rx_fifo_wr_data[10], w_hssi_10g_rx_pcs_rx_fifo_wr_data[9], w_hssi_10g_rx_pcs_rx_fifo_wr_data[8], w_hssi_10g_rx_pcs_rx_fifo_wr_data[7], w_hssi_10g_rx_pcs_rx_fifo_wr_data[6], w_hssi_10g_rx_pcs_rx_fifo_wr_data[5], w_hssi_10g_rx_pcs_rx_fifo_wr_data[4], w_hssi_10g_rx_pcs_rx_fifo_wr_data[3], w_hssi_10g_rx_pcs_rx_fifo_wr_data[2], w_hssi_10g_rx_pcs_rx_fifo_wr_data[1], w_hssi_10g_rx_pcs_rx_fifo_wr_data[0]}),
				.data_in_8g_clock_comp({w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0]}),
				.data_in_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr2_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0]}),
				.rd_ptr2_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0]}),
				.rd_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0]}),
				.rd_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.wr_clk_8g_clock_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_8g_clock_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.wr_en_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.wr_en_8g_clock_comp(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_en_8g_phase_comp(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.wr_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0]}),
				.wr_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0]}),
				.wr_rst_n_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.wr_rst_n_8g_clock_comp(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_n_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_rx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79:0] = 80'b0;
				assign w_hssi_fifo_rx_pcs_data_out_gen3[39:0] = 40'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_tx_pcs
			twentynm_hssi_fifo_tx_pcs #(
				.double_write_mode(hssi_fifo_tx_pcs_double_write_mode),
				.prot_mode(hssi_fifo_tx_pcs_prot_mode),
				.silicon_rev( "20nm5" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_tx_pcs_blockselect),
				.data_out_10g(w_hssi_fifo_tx_pcs_data_out_10g),
				.data_out_8g_phase_comp(w_hssi_fifo_tx_pcs_data_out_8g_phase_comp),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in2_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0]}),
				.data_in_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_en_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.wr_en_8g_phase_comp(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0]}),
				.wr_rst_n_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_tx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_tx_pcs_data_out_10g[72:0] = 73'b0;
				assign w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63:0] = 64'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_rx_pcs
			twentynm_hssi_gen3_rx_pcs #(
				.block_sync(hssi_gen3_rx_pcs_block_sync),
				.block_sync_sm(hssi_gen3_rx_pcs_block_sync_sm),
				.cdr_ctrl_force_unalgn(hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn),
				.lpbk_force(hssi_gen3_rx_pcs_lpbk_force),
				.mode(hssi_gen3_rx_pcs_mode),
				.rate_match_fifo(hssi_gen3_rx_pcs_rate_match_fifo),
				.rate_match_fifo_latency(hssi_gen3_rx_pcs_rate_match_fifo_latency),
				.reconfig_settings(hssi_gen3_rx_pcs_reconfig_settings),
				.reverse_lpbk(hssi_gen3_rx_pcs_reverse_lpbk),
				.rx_b4gb_par_lpbk(hssi_gen3_rx_pcs_rx_b4gb_par_lpbk),
				.rx_force_balign(hssi_gen3_rx_pcs_rx_force_balign),
				.rx_ins_del_one_skip(hssi_gen3_rx_pcs_rx_ins_del_one_skip),
				.rx_num_fixed_pat(hssi_gen3_rx_pcs_rx_num_fixed_pat),
				.rx_test_out_sel(hssi_gen3_rx_pcs_rx_test_out_sel),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_rx_pcs_sup_mode)
			) inst_twentynm_hssi_gen3_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_rx_pcs_avmmreaddata),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.blk_start(w_hssi_gen3_rx_pcs_blk_start),
				.blockselect(w_hssi_gen3_rx_pcs_blockselect),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.data_out(w_hssi_gen3_rx_pcs_data_out),
				.data_valid(w_hssi_gen3_rx_pcs_data_valid),
				.ei_det_int(w_hssi_gen3_rx_pcs_ei_det_int),
				.ei_partial_det_int(w_hssi_gen3_rx_pcs_ei_partial_det_int),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.i_det_int(w_hssi_gen3_rx_pcs_i_det_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data(w_hssi_gen3_rx_pcs_lpbk_data),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.mem_rx_fifo_rd_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr),
				.mem_rx_fifo_wr_clk(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.mem_rx_fifo_wr_data(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data),
				.mem_rx_fifo_wr_en(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.mem_rx_fifo_wr_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr),
				.mem_rx_fifo_wr_rst_n(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_test_out(w_hssi_gen3_rx_pcs_rx_test_out),
				.sync_hdr(w_hssi_gen3_rx_pcs_sync_hdr),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0]}),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.mem_rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_gen3[39], w_hssi_fifo_rx_pcs_data_out_gen3[38], w_hssi_fifo_rx_pcs_data_out_gen3[37], w_hssi_fifo_rx_pcs_data_out_gen3[36], w_hssi_fifo_rx_pcs_data_out_gen3[35], w_hssi_fifo_rx_pcs_data_out_gen3[34], w_hssi_fifo_rx_pcs_data_out_gen3[33], w_hssi_fifo_rx_pcs_data_out_gen3[32], w_hssi_fifo_rx_pcs_data_out_gen3[31], w_hssi_fifo_rx_pcs_data_out_gen3[30], w_hssi_fifo_rx_pcs_data_out_gen3[29], w_hssi_fifo_rx_pcs_data_out_gen3[28], w_hssi_fifo_rx_pcs_data_out_gen3[27], w_hssi_fifo_rx_pcs_data_out_gen3[26], w_hssi_fifo_rx_pcs_data_out_gen3[25], w_hssi_fifo_rx_pcs_data_out_gen3[24], w_hssi_fifo_rx_pcs_data_out_gen3[23], w_hssi_fifo_rx_pcs_data_out_gen3[22], w_hssi_fifo_rx_pcs_data_out_gen3[21], w_hssi_fifo_rx_pcs_data_out_gen3[20], w_hssi_fifo_rx_pcs_data_out_gen3[19], w_hssi_fifo_rx_pcs_data_out_gen3[18], w_hssi_fifo_rx_pcs_data_out_gen3[17], w_hssi_fifo_rx_pcs_data_out_gen3[16], w_hssi_fifo_rx_pcs_data_out_gen3[15], w_hssi_fifo_rx_pcs_data_out_gen3[14], w_hssi_fifo_rx_pcs_data_out_gen3[13], w_hssi_fifo_rx_pcs_data_out_gen3[12], w_hssi_fifo_rx_pcs_data_out_gen3[11], w_hssi_fifo_rx_pcs_data_out_gen3[10], w_hssi_fifo_rx_pcs_data_out_gen3[9], w_hssi_fifo_rx_pcs_data_out_gen3[8], w_hssi_fifo_rx_pcs_data_out_gen3[7], w_hssi_fifo_rx_pcs_data_out_gen3[6], w_hssi_fifo_rx_pcs_data_out_gen3[5], w_hssi_fifo_rx_pcs_data_out_gen3[4], w_hssi_fifo_rx_pcs_data_out_gen3[3], w_hssi_fifo_rx_pcs_data_out_gen3[2], w_hssi_fifo_rx_pcs_data_out_gen3[1], w_hssi_fifo_rx_pcs_data_out_gen3[0]}),
				.par_lpbk_b4gb_in({w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0]}),
				.par_lpbk_in({w_hssi_gen3_tx_pcs_par_lpbk_out[31], w_hssi_gen3_tx_pcs_par_lpbk_out[30], w_hssi_gen3_tx_pcs_par_lpbk_out[29], w_hssi_gen3_tx_pcs_par_lpbk_out[28], w_hssi_gen3_tx_pcs_par_lpbk_out[27], w_hssi_gen3_tx_pcs_par_lpbk_out[26], w_hssi_gen3_tx_pcs_par_lpbk_out[25], w_hssi_gen3_tx_pcs_par_lpbk_out[24], w_hssi_gen3_tx_pcs_par_lpbk_out[23], w_hssi_gen3_tx_pcs_par_lpbk_out[22], w_hssi_gen3_tx_pcs_par_lpbk_out[21], w_hssi_gen3_tx_pcs_par_lpbk_out[20], w_hssi_gen3_tx_pcs_par_lpbk_out[19], w_hssi_gen3_tx_pcs_par_lpbk_out[18], w_hssi_gen3_tx_pcs_par_lpbk_out[17], w_hssi_gen3_tx_pcs_par_lpbk_out[16], w_hssi_gen3_tx_pcs_par_lpbk_out[15], w_hssi_gen3_tx_pcs_par_lpbk_out[14], w_hssi_gen3_tx_pcs_par_lpbk_out[13], w_hssi_gen3_tx_pcs_par_lpbk_out[12], w_hssi_gen3_tx_pcs_par_lpbk_out[11], w_hssi_gen3_tx_pcs_par_lpbk_out[10], w_hssi_gen3_tx_pcs_par_lpbk_out[9], w_hssi_gen3_tx_pcs_par_lpbk_out[8], w_hssi_gen3_tx_pcs_par_lpbk_out[7], w_hssi_gen3_tx_pcs_par_lpbk_out[6], w_hssi_gen3_tx_pcs_par_lpbk_out[5], w_hssi_gen3_tx_pcs_par_lpbk_out[4], w_hssi_gen3_tx_pcs_par_lpbk_out[3], w_hssi_gen3_tx_pcs_par_lpbk_out[2], w_hssi_gen3_tx_pcs_par_lpbk_out[1], w_hssi_gen3_tx_pcs_par_lpbk_out[0]}),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.rcvd_clk(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_pma_clk(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.rxpolarity(w_hssi_pipe_gen3_rxpolarity_int),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.sync_sm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.txdatak_in({w_hssi_pipe_gen3_txdatak_int[3], w_hssi_pipe_gen3_txdatak_int[2], w_hssi_pipe_gen3_txdatak_int[1], w_hssi_pipe_gen3_txdatak_int[0]}),
				
				// UNUSED
				.blk_lockd_int(),
				.skp_det_int()
			);
		end // if generate
		else begin
				assign w_hssi_gen3_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_rx_pcs_blk_algnd_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_delete_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_insert_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_overfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_undfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_rx_pcs_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_partial_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_err_decode_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_i_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data[33:0] = 34'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39:0] = 40'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_rx_test_out[19:0] = 20'b0;
				assign w_hssi_gen3_rx_pcs_sync_hdr[1:0] = 2'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_tx_pcs
			twentynm_hssi_gen3_tx_pcs #(
				.mode(hssi_gen3_tx_pcs_mode),
				.reverse_lpbk(hssi_gen3_tx_pcs_reverse_lpbk),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_tx_pcs_sup_mode),
				.tx_bitslip(hssi_gen3_tx_pcs_tx_bitslip),
				.tx_gbox_byp(hssi_gen3_tx_pcs_tx_gbox_byp)
			) inst_twentynm_hssi_gen3_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_gen3_tx_pcs_blockselect),
				.data_out(w_hssi_gen3_tx_pcs_data_out),
				.par_lpbk_b4gb_out(w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out),
				.par_lpbk_out(w_hssi_gen3_tx_pcs_par_lpbk_out),
				.tx_test_out(w_hssi_gen3_tx_pcs_tx_test_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_start_in(w_hssi_pipe_gen3_tx_blk_start_int),
				.data_in({w_hssi_pipe_gen3_txdata_int[31], w_hssi_pipe_gen3_txdata_int[30], w_hssi_pipe_gen3_txdata_int[29], w_hssi_pipe_gen3_txdata_int[28], w_hssi_pipe_gen3_txdata_int[27], w_hssi_pipe_gen3_txdata_int[26], w_hssi_pipe_gen3_txdata_int[25], w_hssi_pipe_gen3_txdata_int[24], w_hssi_pipe_gen3_txdata_int[23], w_hssi_pipe_gen3_txdata_int[22], w_hssi_pipe_gen3_txdata_int[21], w_hssi_pipe_gen3_txdata_int[20], w_hssi_pipe_gen3_txdata_int[19], w_hssi_pipe_gen3_txdata_int[18], w_hssi_pipe_gen3_txdata_int[17], w_hssi_pipe_gen3_txdata_int[16], w_hssi_pipe_gen3_txdata_int[15], w_hssi_pipe_gen3_txdata_int[14], w_hssi_pipe_gen3_txdata_int[13], w_hssi_pipe_gen3_txdata_int[12], w_hssi_pipe_gen3_txdata_int[11], w_hssi_pipe_gen3_txdata_int[10], w_hssi_pipe_gen3_txdata_int[9], w_hssi_pipe_gen3_txdata_int[8], w_hssi_pipe_gen3_txdata_int[7], w_hssi_pipe_gen3_txdata_int[6], w_hssi_pipe_gen3_txdata_int[5], w_hssi_pipe_gen3_txdata_int[4], w_hssi_pipe_gen3_txdata_int[3], w_hssi_pipe_gen3_txdata_int[2], w_hssi_pipe_gen3_txdata_int[1], w_hssi_pipe_gen3_txdata_int[0]}),
				.data_valid(w_hssi_pipe_gen3_txdataskip_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data_in({w_hssi_gen3_rx_pcs_lpbk_data[33], w_hssi_gen3_rx_pcs_lpbk_data[32], w_hssi_gen3_rx_pcs_lpbk_data[31], w_hssi_gen3_rx_pcs_lpbk_data[30], w_hssi_gen3_rx_pcs_lpbk_data[29], w_hssi_gen3_rx_pcs_lpbk_data[28], w_hssi_gen3_rx_pcs_lpbk_data[27], w_hssi_gen3_rx_pcs_lpbk_data[26], w_hssi_gen3_rx_pcs_lpbk_data[25], w_hssi_gen3_rx_pcs_lpbk_data[24], w_hssi_gen3_rx_pcs_lpbk_data[23], w_hssi_gen3_rx_pcs_lpbk_data[22], w_hssi_gen3_rx_pcs_lpbk_data[21], w_hssi_gen3_rx_pcs_lpbk_data[20], w_hssi_gen3_rx_pcs_lpbk_data[19], w_hssi_gen3_rx_pcs_lpbk_data[18], w_hssi_gen3_rx_pcs_lpbk_data[17], w_hssi_gen3_rx_pcs_lpbk_data[16], w_hssi_gen3_rx_pcs_lpbk_data[15], w_hssi_gen3_rx_pcs_lpbk_data[14], w_hssi_gen3_rx_pcs_lpbk_data[13], w_hssi_gen3_rx_pcs_lpbk_data[12], w_hssi_gen3_rx_pcs_lpbk_data[11], w_hssi_gen3_rx_pcs_lpbk_data[10], w_hssi_gen3_rx_pcs_lpbk_data[9], w_hssi_gen3_rx_pcs_lpbk_data[8], w_hssi_gen3_rx_pcs_lpbk_data[7], w_hssi_gen3_rx_pcs_lpbk_data[6], w_hssi_gen3_rx_pcs_lpbk_data[5], w_hssi_gen3_rx_pcs_lpbk_data[4], w_hssi_gen3_rx_pcs_lpbk_data[3], w_hssi_gen3_rx_pcs_lpbk_data[2], w_hssi_gen3_rx_pcs_lpbk_data[1], w_hssi_gen3_rx_pcs_lpbk_data[0]}),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.sync_in({w_hssi_pipe_gen3_tx_sync_hdr_int[1], w_hssi_pipe_gen3_tx_sync_hdr_int[0]}),
				.tx_pma_clk(w_hssi_8g_tx_pcs_clk_out_gen3),
				.tx_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn)
			);
		end // if generate
		else begin
				assign w_hssi_gen3_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_tx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_tx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35:0] = 36'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_tx_test_out[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_rx_pcs
			twentynm_hssi_krfec_rx_pcs #(
				.blksync_cor_en(hssi_krfec_rx_pcs_blksync_cor_en),
				.bypass_gb(hssi_krfec_rx_pcs_bypass_gb),
				.clr_ctrl(hssi_krfec_rx_pcs_clr_ctrl),
				.ctrl_bit_reverse(hssi_krfec_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_rx_pcs_data_bit_reverse),
				.dv_start(hssi_krfec_rx_pcs_dv_start),
				.err_mark_type(hssi_krfec_rx_pcs_err_mark_type),
				.error_marking_en(hssi_krfec_rx_pcs_error_marking_en),
				.low_latency_en(hssi_krfec_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_krfec_rx_pcs_lpbk_mode),
				.parity_invalid_enum(hssi_krfec_rx_pcs_parity_invalid_enum),
				.parity_valid_num(hssi_krfec_rx_pcs_parity_valid_num),
				.pipeln_blksync(hssi_krfec_rx_pcs_pipeln_blksync),
				.pipeln_descrm(hssi_krfec_rx_pcs_pipeln_descrm),
				.pipeln_errcorrect(hssi_krfec_rx_pcs_pipeln_errcorrect),
				.pipeln_errtrap_ind(hssi_krfec_rx_pcs_pipeln_errtrap_ind),
				.pipeln_errtrap_lfsr(hssi_krfec_rx_pcs_pipeln_errtrap_lfsr),
				.pipeln_errtrap_loc(hssi_krfec_rx_pcs_pipeln_errtrap_loc),
				.pipeln_errtrap_pat(hssi_krfec_rx_pcs_pipeln_errtrap_pat),
				.pipeln_gearbox(hssi_krfec_rx_pcs_pipeln_gearbox),
				.pipeln_syndrm(hssi_krfec_rx_pcs_pipeln_syndrm),
				.pipeln_trans_dec(hssi_krfec_rx_pcs_pipeln_trans_dec),
				.prot_mode(hssi_krfec_rx_pcs_prot_mode),
				.receive_order(hssi_krfec_rx_pcs_receive_order),
				.reconfig_settings(hssi_krfec_rx_pcs_reconfig_settings),
				.rx_testbus_sel(hssi_krfec_rx_pcs_rx_testbus_sel),
				.signal_ok_en(hssi_krfec_rx_pcs_signal_ok_en),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_rx_pcs_sup_mode)
			) inst_twentynm_hssi_krfec_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_rx_pcs_blockselect),
				.rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.rx_control_out(w_hssi_krfec_rx_pcs_rx_control_out),
				.rx_data_out(w_hssi_krfec_rx_pcs_rx_data_out),
				.rx_data_status(w_hssi_krfec_rx_pcs_rx_data_status),
				.rx_data_valid_out(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.rx_signal_ok_out(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.rx_data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0]}),
				.rx_krfec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_krfec_reg(),
				.pld_10g_krfec_rx_blk_lock_krfec_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg(),
				.pld_10g_krfec_rx_frame_krfec_reg(),
				.pld_10g_krfec_rx_frame_krfec_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_rx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_block_lock = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_control_out[9:0] = 10'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_status[1:0] = 2'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_valid_out = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_frame = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_signal_ok_out = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_tx_pcs
			twentynm_hssi_krfec_tx_pcs #(
				.burst_err(hssi_krfec_tx_pcs_burst_err),
				.burst_err_len(hssi_krfec_tx_pcs_burst_err_len),
				.ctrl_bit_reverse(hssi_krfec_tx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_tx_pcs_data_bit_reverse),
				.enc_frame_query(hssi_krfec_tx_pcs_enc_frame_query),
				.low_latency_en(hssi_krfec_tx_pcs_low_latency_en),
				.pipeln_encoder(hssi_krfec_tx_pcs_pipeln_encoder),
				.pipeln_scrambler(hssi_krfec_tx_pcs_pipeln_scrambler),
				.prot_mode(hssi_krfec_tx_pcs_prot_mode),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_tx_pcs_sup_mode),
				.transcode_err(hssi_krfec_tx_pcs_transcode_err),
				.transmit_order(hssi_krfec_tx_pcs_transmit_order),
				.tx_testbus_sel(hssi_krfec_tx_pcs_tx_testbus_sel)
			) inst_twentynm_hssi_krfec_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_tx_pcs_blockselect),
				.tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.tx_data_out(w_hssi_krfec_tx_pcs_tx_data_out),
				.tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.tx_test_data(w_hssi_krfec_tx_pcs_tx_test_data),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.tx_control_in({w_hssi_10g_tx_pcs_tx_control_out_krfec[8], w_hssi_10g_tx_pcs_tx_control_out_krfec[7], w_hssi_10g_tx_pcs_tx_control_out_krfec[6], w_hssi_10g_tx_pcs_tx_control_out_krfec[5], w_hssi_10g_tx_pcs_tx_control_out_krfec[4], w_hssi_10g_tx_pcs_tx_control_out_krfec[3], w_hssi_10g_tx_pcs_tx_control_out_krfec[2], w_hssi_10g_tx_pcs_tx_control_out_krfec[1], w_hssi_10g_tx_pcs_tx_control_out_krfec[0]}),
				.tx_data_in({w_hssi_10g_tx_pcs_tx_data_out_krfec[63], w_hssi_10g_tx_pcs_tx_data_out_krfec[62], w_hssi_10g_tx_pcs_tx_data_out_krfec[61], w_hssi_10g_tx_pcs_tx_data_out_krfec[60], w_hssi_10g_tx_pcs_tx_data_out_krfec[59], w_hssi_10g_tx_pcs_tx_data_out_krfec[58], w_hssi_10g_tx_pcs_tx_data_out_krfec[57], w_hssi_10g_tx_pcs_tx_data_out_krfec[56], w_hssi_10g_tx_pcs_tx_data_out_krfec[55], w_hssi_10g_tx_pcs_tx_data_out_krfec[54], w_hssi_10g_tx_pcs_tx_data_out_krfec[53], w_hssi_10g_tx_pcs_tx_data_out_krfec[52], w_hssi_10g_tx_pcs_tx_data_out_krfec[51], w_hssi_10g_tx_pcs_tx_data_out_krfec[50], w_hssi_10g_tx_pcs_tx_data_out_krfec[49], w_hssi_10g_tx_pcs_tx_data_out_krfec[48], w_hssi_10g_tx_pcs_tx_data_out_krfec[47], w_hssi_10g_tx_pcs_tx_data_out_krfec[46], w_hssi_10g_tx_pcs_tx_data_out_krfec[45], w_hssi_10g_tx_pcs_tx_data_out_krfec[44], w_hssi_10g_tx_pcs_tx_data_out_krfec[43], w_hssi_10g_tx_pcs_tx_data_out_krfec[42], w_hssi_10g_tx_pcs_tx_data_out_krfec[41], w_hssi_10g_tx_pcs_tx_data_out_krfec[40], w_hssi_10g_tx_pcs_tx_data_out_krfec[39], w_hssi_10g_tx_pcs_tx_data_out_krfec[38], w_hssi_10g_tx_pcs_tx_data_out_krfec[37], w_hssi_10g_tx_pcs_tx_data_out_krfec[36], w_hssi_10g_tx_pcs_tx_data_out_krfec[35], w_hssi_10g_tx_pcs_tx_data_out_krfec[34], w_hssi_10g_tx_pcs_tx_data_out_krfec[33], w_hssi_10g_tx_pcs_tx_data_out_krfec[32], w_hssi_10g_tx_pcs_tx_data_out_krfec[31], w_hssi_10g_tx_pcs_tx_data_out_krfec[30], w_hssi_10g_tx_pcs_tx_data_out_krfec[29], w_hssi_10g_tx_pcs_tx_data_out_krfec[28], w_hssi_10g_tx_pcs_tx_data_out_krfec[27], w_hssi_10g_tx_pcs_tx_data_out_krfec[26], w_hssi_10g_tx_pcs_tx_data_out_krfec[25], w_hssi_10g_tx_pcs_tx_data_out_krfec[24], w_hssi_10g_tx_pcs_tx_data_out_krfec[23], w_hssi_10g_tx_pcs_tx_data_out_krfec[22], w_hssi_10g_tx_pcs_tx_data_out_krfec[21], w_hssi_10g_tx_pcs_tx_data_out_krfec[20], w_hssi_10g_tx_pcs_tx_data_out_krfec[19], w_hssi_10g_tx_pcs_tx_data_out_krfec[18], w_hssi_10g_tx_pcs_tx_data_out_krfec[17], w_hssi_10g_tx_pcs_tx_data_out_krfec[16], w_hssi_10g_tx_pcs_tx_data_out_krfec[15], w_hssi_10g_tx_pcs_tx_data_out_krfec[14], w_hssi_10g_tx_pcs_tx_data_out_krfec[13], w_hssi_10g_tx_pcs_tx_data_out_krfec[12], w_hssi_10g_tx_pcs_tx_data_out_krfec[11], w_hssi_10g_tx_pcs_tx_data_out_krfec[10], w_hssi_10g_tx_pcs_tx_data_out_krfec[9], w_hssi_10g_tx_pcs_tx_data_out_krfec[8], w_hssi_10g_tx_pcs_tx_data_out_krfec[7], w_hssi_10g_tx_pcs_tx_data_out_krfec[6], w_hssi_10g_tx_pcs_tx_data_out_krfec[5], w_hssi_10g_tx_pcs_tx_data_out_krfec[4], w_hssi_10g_tx_pcs_tx_data_out_krfec[3], w_hssi_10g_tx_pcs_tx_data_out_krfec[2], w_hssi_10g_tx_pcs_tx_data_out_krfec[1], w_hssi_10g_tx_pcs_tx_data_out_krfec[0]}),
				.tx_data_valid_in(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_krfec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_krfec_reg(),
				.pld_krfec_tx_alignment_plddirect_reg(),
				.pld_krfec_tx_alignment_reg()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_tx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_alignment = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_test_data[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen1_2
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen1_2
			twentynm_hssi_pipe_gen1_2 #(
				.elec_idle_delay_val(hssi_pipe_gen1_2_elec_idle_delay_val),
				.error_replace_pad(hssi_pipe_gen1_2_error_replace_pad),
				.hip_mode(hssi_pipe_gen1_2_hip_mode),
				.ind_error_reporting(hssi_pipe_gen1_2_ind_error_reporting),
				.phystatus_delay_val(hssi_pipe_gen1_2_phystatus_delay_val),
				.phystatus_rst_toggle(hssi_pipe_gen1_2_phystatus_rst_toggle),
				.pipe_byte_de_serializer_en(hssi_pipe_gen1_2_pipe_byte_de_serializer_en),
				.prot_mode(hssi_pipe_gen1_2_prot_mode),
				.reconfig_settings(hssi_pipe_gen1_2_reconfig_settings),
				.rx_pipe_enable(hssi_pipe_gen1_2_rx_pipe_enable),
				.rxdetect_bypass(hssi_pipe_gen1_2_rxdetect_bypass),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen1_2_sup_mode),
				.tx_pipe_enable(hssi_pipe_gen1_2_tx_pipe_enable),
				.txswing(hssi_pipe_gen1_2_txswing)
			) inst_twentynm_hssi_pipe_gen1_2 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen1_2_avmmreaddata),
				.blockselect(w_hssi_pipe_gen1_2_blockselect),
				.current_coeff(w_hssi_pipe_gen1_2_current_coeff),
				.phystatus(w_hssi_pipe_gen1_2_phystatus),
				.polarity_inversion_rx(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rev_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.rxelectricalidle_out(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxstatus(w_hssi_pipe_gen1_2_rxstatus),
				.rxvalid(w_hssi_pipe_gen1_2_rxvalid),
				.tx_elec_idle_out(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pipe_rx_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.power_state_transition_done_ena(1'b0),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rev_loopbk_pcs_gen3(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.revloopback(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.rx_pipe_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rxd({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxelectricalidle(w_hssi_8g_rx_pcs_eidle_detected),
				.rxelectricalidle_pcs_gen3(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.rxpolarity_pcs_gen3(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.tx_elec_idle_comp(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.txd_ch({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswingport(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.pld_8g_rxpolarity_pipe3_reg(),
				.rxd_ch(),
				.txd()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen1_2_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen1_2_blockselect = 1'b0;
				assign w_hssi_pipe_gen1_2_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen1_2_phystatus = 1'b0;
				assign w_hssi_pipe_gen1_2_polarity_inversion_rx = 1'b0;
				assign w_hssi_pipe_gen1_2_rev_loopbk = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelectricalidle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen1_2_rxvalid = 1'b0;
				assign w_hssi_pipe_gen1_2_tx_elec_idle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_txdetectrx = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen3
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen3
			twentynm_hssi_pipe_gen3 #(
				.bypass_rx_detection_enable(hssi_pipe_gen3_bypass_rx_detection_enable),
				.bypass_rx_preset(hssi_pipe_gen3_bypass_rx_preset),
				.bypass_rx_preset_enable(hssi_pipe_gen3_bypass_rx_preset_enable),
				.bypass_tx_coefficent(hssi_pipe_gen3_bypass_tx_coefficent),
				.bypass_tx_coefficent_enable(hssi_pipe_gen3_bypass_tx_coefficent_enable),
				.elecidle_delay_g3(hssi_pipe_gen3_elecidle_delay_g3),
				.ind_error_reporting(hssi_pipe_gen3_ind_error_reporting),
				.mode(hssi_pipe_gen3_mode),
				.phy_status_delay_g12(hssi_pipe_gen3_phy_status_delay_g12),
				.phy_status_delay_g3(hssi_pipe_gen3_phy_status_delay_g3),
				.phystatus_rst_toggle_g12(hssi_pipe_gen3_phystatus_rst_toggle_g12),
				.phystatus_rst_toggle_g3(hssi_pipe_gen3_phystatus_rst_toggle_g3),
				.rate_match_pad_insertion(hssi_pipe_gen3_rate_match_pad_insertion),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen3_sup_mode),
				.test_out_sel(hssi_pipe_gen3_test_out_sel)
			) inst_twentynm_hssi_pipe_gen3 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen3_avmmreaddata),
				.blockselect(w_hssi_pipe_gen3_blockselect),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.phystatus(w_hssi_pipe_gen3_phystatus),
				.pma_current_coeff(w_hssi_pipe_gen3_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_pipe_gen3_pma_current_rxpreset),
				.pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.rev_lpbk_8gpcs_out(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.rev_lpbk_int(w_hssi_pipe_gen3_rev_lpbk_int),
				.rx_blk_start(w_hssi_pipe_gen3_rx_blk_start),
				.rx_sync_hdr(w_hssi_pipe_gen3_rx_sync_hdr),
				.rxd_8gpcs_out(w_hssi_pipe_gen3_rxd_8gpcs_out),
				.rxdataskip(w_hssi_pipe_gen3_rxdataskip),
				.rxelecidle(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity_8gpcs_out(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.rxpolarity_int(w_hssi_pipe_gen3_rxpolarity_int),
				.rxstatus(w_hssi_pipe_gen3_rxstatus),
				.rxvalid(w_hssi_pipe_gen3_rxvalid),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.test_out(w_hssi_pipe_gen3_test_out),
				.tx_blk_start_int(w_hssi_pipe_gen3_tx_blk_start_int),
				.tx_sync_hdr_int(w_hssi_pipe_gen3_tx_sync_hdr_int),
				.txdata_int(w_hssi_pipe_gen3_txdata_int),
				.txdatak_int(w_hssi_pipe_gen3_txdatak_int),
				.txdataskip_int(w_hssi_pipe_gen3_txdataskip_int),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.current_coeff({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0]}),
				.current_rxpreset({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0]}),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.pcs_asn_bundling_in({w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0]}),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pipe_tx_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_blk_start_int(w_hssi_gen3_rx_pcs_blk_start),
				.rx_sync_hdr_int({w_hssi_gen3_rx_pcs_sync_hdr[1], w_hssi_gen3_rx_pcs_sync_hdr[0]}),
				.rx_test_out({w_hssi_gen3_rx_pcs_rx_test_out[19], w_hssi_gen3_rx_pcs_rx_test_out[18], w_hssi_gen3_rx_pcs_rx_test_out[17], w_hssi_gen3_rx_pcs_rx_test_out[16], w_hssi_gen3_rx_pcs_rx_test_out[15], w_hssi_gen3_rx_pcs_rx_test_out[14], w_hssi_gen3_rx_pcs_rx_test_out[13], w_hssi_gen3_rx_pcs_rx_test_out[12], w_hssi_gen3_rx_pcs_rx_test_out[11], w_hssi_gen3_rx_pcs_rx_test_out[10], w_hssi_gen3_rx_pcs_rx_test_out[9], w_hssi_gen3_rx_pcs_rx_test_out[8], w_hssi_gen3_rx_pcs_rx_test_out[7], w_hssi_gen3_rx_pcs_rx_test_out[6], w_hssi_gen3_rx_pcs_rx_test_out[5], w_hssi_gen3_rx_pcs_rx_test_out[4], w_hssi_gen3_rx_pcs_rx_test_out[3], w_hssi_gen3_rx_pcs_rx_test_out[2], w_hssi_gen3_rx_pcs_rx_test_out[1], w_hssi_gen3_rx_pcs_rx_test_out[0]}),
				.rxd_8gpcs_in({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxdata_int({w_hssi_gen3_rx_pcs_data_out[31], w_hssi_gen3_rx_pcs_data_out[30], w_hssi_gen3_rx_pcs_data_out[29], w_hssi_gen3_rx_pcs_data_out[28], w_hssi_gen3_rx_pcs_data_out[27], w_hssi_gen3_rx_pcs_data_out[26], w_hssi_gen3_rx_pcs_data_out[25], w_hssi_gen3_rx_pcs_data_out[24], w_hssi_gen3_rx_pcs_data_out[23], w_hssi_gen3_rx_pcs_data_out[22], w_hssi_gen3_rx_pcs_data_out[21], w_hssi_gen3_rx_pcs_data_out[20], w_hssi_gen3_rx_pcs_data_out[19], w_hssi_gen3_rx_pcs_data_out[18], w_hssi_gen3_rx_pcs_data_out[17], w_hssi_gen3_rx_pcs_data_out[16], w_hssi_gen3_rx_pcs_data_out[15], w_hssi_gen3_rx_pcs_data_out[14], w_hssi_gen3_rx_pcs_data_out[13], w_hssi_gen3_rx_pcs_data_out[12], w_hssi_gen3_rx_pcs_data_out[11], w_hssi_gen3_rx_pcs_data_out[10], w_hssi_gen3_rx_pcs_data_out[9], w_hssi_gen3_rx_pcs_data_out[8], w_hssi_gen3_rx_pcs_data_out[7], w_hssi_gen3_rx_pcs_data_out[6], w_hssi_gen3_rx_pcs_data_out[5], w_hssi_gen3_rx_pcs_data_out[4], w_hssi_gen3_rx_pcs_data_out[3], w_hssi_gen3_rx_pcs_data_out[2], w_hssi_gen3_rx_pcs_data_out[1], w_hssi_gen3_rx_pcs_data_out[0]}),
				.rxdatak_int({1'b0, 1'b0, 1'b0, 1'b0}),
				.rxdataskip_int(w_hssi_gen3_rx_pcs_data_valid),
				.rxelecidle_8gpcs_in(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.tx_blk_start(w_hssi_8g_tx_pcs_tx_blk_start_out[0]),
				.tx_sync_hdr({w_hssi_8g_tx_pcs_tx_sync_hdr_out[1], w_hssi_8g_tx_pcs_tx_sync_hdr_out[0]}),
				.tx_test_out({w_hssi_gen3_tx_pcs_tx_test_out[19], w_hssi_gen3_tx_pcs_tx_test_out[18], w_hssi_gen3_tx_pcs_tx_test_out[17], w_hssi_gen3_tx_pcs_tx_test_out[16], w_hssi_gen3_tx_pcs_tx_test_out[15], w_hssi_gen3_tx_pcs_tx_test_out[14], w_hssi_gen3_tx_pcs_tx_test_out[13], w_hssi_gen3_tx_pcs_tx_test_out[12], w_hssi_gen3_tx_pcs_tx_test_out[11], w_hssi_gen3_tx_pcs_tx_test_out[10], w_hssi_gen3_tx_pcs_tx_test_out[9], w_hssi_gen3_tx_pcs_tx_test_out[8], w_hssi_gen3_tx_pcs_tx_test_out[7], w_hssi_gen3_tx_pcs_tx_test_out[6], w_hssi_gen3_tx_pcs_tx_test_out[5], w_hssi_gen3_tx_pcs_tx_test_out[4], w_hssi_gen3_tx_pcs_tx_test_out[3], w_hssi_gen3_tx_pcs_tx_test_out[2], w_hssi_gen3_tx_pcs_tx_test_out[1], w_hssi_gen3_tx_pcs_tx_test_out[0]}),
				.txcompliance(w_hssi_8g_tx_pcs_txcompliance_out),
				.txdata({w_hssi_8g_tx_pcs_tx_data_out[31], w_hssi_8g_tx_pcs_tx_data_out[30], w_hssi_8g_tx_pcs_tx_data_out[29], w_hssi_8g_tx_pcs_tx_data_out[28], w_hssi_8g_tx_pcs_tx_data_out[27], w_hssi_8g_tx_pcs_tx_data_out[26], w_hssi_8g_tx_pcs_tx_data_out[25], w_hssi_8g_tx_pcs_tx_data_out[24], w_hssi_8g_tx_pcs_tx_data_out[23], w_hssi_8g_tx_pcs_tx_data_out[22], w_hssi_8g_tx_pcs_tx_data_out[21], w_hssi_8g_tx_pcs_tx_data_out[20], w_hssi_8g_tx_pcs_tx_data_out[19], w_hssi_8g_tx_pcs_tx_data_out[18], w_hssi_8g_tx_pcs_tx_data_out[17], w_hssi_8g_tx_pcs_tx_data_out[16], w_hssi_8g_tx_pcs_tx_data_out[15], w_hssi_8g_tx_pcs_tx_data_out[14], w_hssi_8g_tx_pcs_tx_data_out[13], w_hssi_8g_tx_pcs_tx_data_out[12], w_hssi_8g_tx_pcs_tx_data_out[11], w_hssi_8g_tx_pcs_tx_data_out[10], w_hssi_8g_tx_pcs_tx_data_out[9], w_hssi_8g_tx_pcs_tx_data_out[8], w_hssi_8g_tx_pcs_tx_data_out[7], w_hssi_8g_tx_pcs_tx_data_out[6], w_hssi_8g_tx_pcs_tx_data_out[5], w_hssi_8g_tx_pcs_tx_data_out[4], w_hssi_8g_tx_pcs_tx_data_out[3], w_hssi_8g_tx_pcs_tx_data_out[2], w_hssi_8g_tx_pcs_tx_data_out[1], w_hssi_8g_tx_pcs_tx_data_out[0]}),
				.txdatak({w_hssi_8g_tx_pcs_tx_datak_out[3], w_hssi_8g_tx_pcs_tx_datak_out[2], w_hssi_8g_tx_pcs_tx_datak_out[1], w_hssi_8g_tx_pcs_tx_datak_out[0]}),
				.txdataskip(w_hssi_8g_tx_pcs_tx_data_valid_out[0]),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_8g_tx_pcs_txelecidle_out),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.dis_pc_byte(),
				.pma_rx_det_pd(),
				.pma_txdeemph(),
				.pma_txmargin(),
				.pma_txswing(),
				.reset_pc_prts()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen3_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen3_blockselect = 1'b0;
				assign w_hssi_pipe_gen3_gen3_clk_sel = 1'b0;
				assign w_hssi_pipe_gen3_pcs_rst = 1'b0;
				assign w_hssi_pipe_gen3_phystatus = 1'b0;
				assign w_hssi_pipe_gen3_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen3_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_pma_tx_elec_idle = 1'b0;
				assign w_hssi_pipe_gen3_pma_txdetectrx = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_int = 1'b0;
				assign w_hssi_pipe_gen3_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_rxd_8gpcs_out[63:0] = 64'b0;
				assign w_hssi_pipe_gen3_rxdataskip[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_int = 1'b0;
				assign w_hssi_pipe_gen3_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_rxvalid = 1'b0;
				assign w_hssi_pipe_gen3_shutdown_clk = 1'b0;
				assign w_hssi_pipe_gen3_test_out[19:0] = 20'b0;
				assign w_hssi_pipe_gen3_tx_blk_start_int = 1'b0;
				assign w_hssi_pipe_gen3_tx_sync_hdr_int[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_txdata_int[31:0] = 32'b0;
				assign w_hssi_pipe_gen3_txdatak_int[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_txdataskip_int = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pcs_pma_interface
			twentynm_hssi_rx_pcs_pma_interface #(
				.block_sel(hssi_rx_pcs_pma_interface_block_sel),
				.channel_operation_mode(hssi_rx_pcs_pma_interface_channel_operation_mode),
				.clkslip_sel(hssi_rx_pcs_pma_interface_clkslip_sel),
				.lpbk_en(hssi_rx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_rx_pcs_pma_interface_master_clk_sel),
				.pldif_datawidth_mode(hssi_rx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_rx(hssi_rx_pcs_pma_interface_pma_dw_rx),
				.pma_if_dft_en(hssi_rx_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_rx_pcs_pma_interface_pma_if_dft_val),
				.prbs9_dwidth(hssi_rx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_rx_pcs_pma_interface_prbs_clken),
				.prbs_ver(hssi_rx_pcs_pma_interface_prbs_ver),
				.prot_mode_rx(hssi_rx_pcs_pma_interface_prot_mode_rx),
				.reconfig_settings(hssi_rx_pcs_pma_interface_reconfig_settings),
				.rx_dyn_polarity_inversion(hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion),
				.rx_lpbk_en(hssi_rx_pcs_pma_interface_rx_lpbk_en),
				.rx_prbs_force_signal_ok(hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok),
				.rx_prbs_mask(hssi_rx_pcs_pma_interface_rx_prbs_mask),
				.rx_prbs_mode(hssi_rx_pcs_pma_interface_rx_prbs_mode),
				.rx_signalok_signaldet_sel(hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel),
				.rx_static_polarity_inversion(hssi_rx_pcs_pma_interface_rx_static_polarity_inversion),
				.rx_uhsif_lpbk_en(hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sup_mode(hssi_rx_pcs_pma_interface_sup_mode)
			) inst_twentynm_hssi_rx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.int_pmaif_10g_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data),
				.int_pmaif_10g_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.int_pmaif_8g_pudi(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi),
				.int_pmaif_8g_rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.int_pmaif_8g_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.int_pmaif_8g_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.int_pmaif_8g_sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.int_pmaif_g3_pma_data_in(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in),
				.int_pmaif_g3_pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.int_pmaif_g3_pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.int_pmaif_g3_pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.int_pmaif_krfec_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data),
				.int_pmaif_krfec_rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.int_pmaif_pldif_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pmaif_pldif_prbs_err_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pmaif_pldif_rx_clkdiv(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pmaif_pldif_rx_clkdiv_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pmaif_pldif_rx_data(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data),
				.int_pmaif_pldif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pmaif_pldif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pmaif_pldif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pmaif_pldif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.pma_eye_monitor(w_hssi_rx_pcs_pma_interface_pma_eye_monitor),
				.pma_rx_clkslip(w_hssi_rx_pcs_pma_interface_pma_rx_clkslip),
				.pma_rxpma_rstb(w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb),
				.rx_pmaif_test_out(w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out),
				.rx_prbs_ver_test(w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.int_pmaif_8g_rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.int_pmaif_pldif_eye_monitor({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0]}),
				.int_pmaif_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pmaif_pldif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pmaif_pldif_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pmaif_pldif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pma_rx_clkdiv_user(in_pma_rx_clkdiv_user),
				.pma_rx_detect_valid(in_pma_rx_detect_valid),
				.pma_rx_found(in_pma_rx_found),
				.pma_rx_pma_clk(in_pma_rx_pma_clk),
				.pma_rx_pma_data({in_pma_rx_pma_data[63], in_pma_rx_pma_data[62], in_pma_rx_pma_data[61], in_pma_rx_pma_data[60], in_pma_rx_pma_data[59], in_pma_rx_pma_data[58], in_pma_rx_pma_data[57], in_pma_rx_pma_data[56], in_pma_rx_pma_data[55], in_pma_rx_pma_data[54], in_pma_rx_pma_data[53], in_pma_rx_pma_data[52], in_pma_rx_pma_data[51], in_pma_rx_pma_data[50], in_pma_rx_pma_data[49], in_pma_rx_pma_data[48], in_pma_rx_pma_data[47], in_pma_rx_pma_data[46], in_pma_rx_pma_data[45], in_pma_rx_pma_data[44], in_pma_rx_pma_data[43], in_pma_rx_pma_data[42], in_pma_rx_pma_data[41], in_pma_rx_pma_data[40], in_pma_rx_pma_data[39], in_pma_rx_pma_data[38], in_pma_rx_pma_data[37], in_pma_rx_pma_data[36], in_pma_rx_pma_data[35], in_pma_rx_pma_data[34], in_pma_rx_pma_data[33], in_pma_rx_pma_data[32], in_pma_rx_pma_data[31], in_pma_rx_pma_data[30], in_pma_rx_pma_data[29], in_pma_rx_pma_data[28], in_pma_rx_pma_data[27], in_pma_rx_pma_data[26], in_pma_rx_pma_data[25], in_pma_rx_pma_data[24], in_pma_rx_pma_data[23], in_pma_rx_pma_data[22], in_pma_rx_pma_data[21], in_pma_rx_pma_data[20], in_pma_rx_pma_data[19], in_pma_rx_pma_data[18], in_pma_rx_pma_data[17], in_pma_rx_pma_data[16], in_pma_rx_pma_data[15], in_pma_rx_pma_data[14], in_pma_rx_pma_data[13], in_pma_rx_pma_data[12], in_pma_rx_pma_data[11], in_pma_rx_pma_data[10], in_pma_rx_pma_data[9], in_pma_rx_pma_data[8], in_pma_rx_pma_data[7], in_pma_rx_pma_data[6], in_pma_rx_pma_data[5], in_pma_rx_pma_data[4], in_pma_rx_pma_data[3], in_pma_rx_pma_data[2], in_pma_rx_pma_data[1], in_pma_rx_pma_data[0]}),
				.pma_rx_signal_ok(in_pma_rx_signal_ok),
				.pma_rxpll_lock(in_pma_rxpll_lock),
				.pma_signal_det(in_pma_signal_det),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.tx_pma_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0]}),
				.tx_pma_uhsif_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0]}),
				
				// UNUSED
				.int_pmaif_g3_rcvd_clk(),
				.prbs_err_lt()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31:0] = 32'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5:0] = 6'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rx_clkslip = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pld_pcs_interface
			twentynm_hssi_rx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx),
				.hd_10g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx),
				.hd_10g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx),
				.hd_10g_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx),
				.hd_10g_lpbk_en(hssi_rx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx),
				.hd_10g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx),
				.hd_10g_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx),
				.hd_10g_test_bus_mode(hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode),
				.hd_8g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx),
				.hd_8g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx),
				.hd_8g_hip_mode(hssi_rx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_rx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx),
				.hd_8g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx),
				.hd_chnl_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_clklow_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz),
				.hd_chnl_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx),
				.hd_chnl_fref_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz),
				.hd_chnl_frequency_rules_en(hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_rx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_rx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx),
				.hd_chnl_lpbk_en(hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx),
				.hd_chnl_pld_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz),
				.hd_chnl_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx),
				.hd_chnl_pma_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz),
				.hd_chnl_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx),
				.hd_chnl_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx),
				.hd_chnl_transparent_pcs_rx(hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx),
				.hd_fifo_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx),
				.hd_fifo_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx),
				.hd_g3_prot_mode(hssi_rx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx),
				.hd_krfec_lpbk_en(hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx),
				.hd_krfec_test_bus_mode(hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode),
				.hd_pldif_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx),
				.hd_pmaif_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_lpbk_en(hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx),
				.hd_pmaif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx),
				.hd_pmaif_sim_mode(hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_rx_block_sel(hssi_rx_pld_pcs_interface_pcs_rx_block_sel),
				.pcs_rx_clk_out_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel),
				.pcs_rx_clk_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_sel),
				.pcs_rx_hip_clk_en(hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en),
				.pcs_rx_output_sel(hssi_rx_pld_pcs_interface_pcs_rx_output_sel),
				.reconfig_settings(hssi_rx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm5" )       //PARAM_HIDE
			) inst_twentynm_hssi_rx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pld_pcs_interface_blockselect),
				.hip_rx_ctrl(w_hssi_rx_pld_pcs_interface_hip_rx_ctrl),
				.hip_rx_data(w_hssi_rx_pld_pcs_interface_hip_rx_data),
				.int_pldif_10g_rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.int_pldif_10g_rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.int_pldif_10g_rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.int_pldif_10g_rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.int_pldif_10g_rx_control_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb),
				.int_pldif_10g_rx_data_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb),
				.int_pldif_10g_rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.int_pldif_10g_rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.int_pldif_10g_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.int_pldif_10g_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.int_pldif_10g_rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.int_pldif_8g_a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.int_pldif_8g_bitloc_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.int_pldif_8g_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.int_pldif_8g_byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.int_pldif_8g_encdt(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.int_pldif_8g_pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.int_pldif_8g_rdenable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.int_pldif_8g_rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.int_pldif_8g_rxurstpcs_n(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.int_pldif_8g_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.int_pldif_8g_wrdisable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.int_pldif_g3_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.int_pldif_krfec_rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.int_pldif_pmaif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pldif_pmaif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pldif_pmaif_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pldif_pmaif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pld_10g_krfec_rx_blk_lock(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock),
				.pld_10g_krfec_rx_diag_data_status(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status),
				.pld_10g_krfec_rx_frame(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame),
				.pld_10g_rx_align_val(w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val),
				.pld_10g_rx_crc32_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err),
				.pld_10g_rx_data_valid(w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid),
				.pld_10g_rx_empty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty),
				.pld_10g_rx_fifo_del(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del),
				.pld_10g_rx_fifo_insert(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert),
				.pld_10g_rx_fifo_num(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num),
				.pld_10g_rx_frame_lock(w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock),
				.pld_10g_rx_hi_ber(w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber),
				.pld_10g_rx_oflw_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err),
				.pld_10g_rx_pempty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty),
				.pld_10g_rx_pfull(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull),
				.pld_8g_a1a2_k1k2_flag(w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag),
				.pld_8g_empty_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf),
				.pld_8g_empty_rx(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx),
				.pld_8g_full_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf),
				.pld_8g_full_rx(w_hssi_rx_pld_pcs_interface_pld_8g_full_rx),
				.pld_8g_rxelecidle(w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle),
				.pld_8g_signal_detect_out(w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out),
				.pld_8g_wa_boundary(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary),
				.pld_pcs_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out),
				.pld_pma_clkdiv_rx_user(w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user),
				.pld_pma_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out),
				.pld_pma_signal_ok(w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok),
				.pld_rx_control(w_hssi_rx_pld_pcs_interface_pld_rx_control),
				.pld_rx_data(w_hssi_rx_pld_pcs_interface_pld_rx_data),
				.pld_rx_prbs_done(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done),
				.pld_rx_prbs_err(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.int_pldif_10g_rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.int_pldif_10g_rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.int_pldif_10g_rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_10g_rx_control({w_hssi_10g_rx_pcs_rx_control[19], w_hssi_10g_rx_pcs_rx_control[18], w_hssi_10g_rx_pcs_rx_control[17], w_hssi_10g_rx_pcs_rx_control[16], w_hssi_10g_rx_pcs_rx_control[15], w_hssi_10g_rx_pcs_rx_control[14], w_hssi_10g_rx_pcs_rx_control[13], w_hssi_10g_rx_pcs_rx_control[12], w_hssi_10g_rx_pcs_rx_control[11], w_hssi_10g_rx_pcs_rx_control[10], w_hssi_10g_rx_pcs_rx_control[9], w_hssi_10g_rx_pcs_rx_control[8], w_hssi_10g_rx_pcs_rx_control[7], w_hssi_10g_rx_pcs_rx_control[6], w_hssi_10g_rx_pcs_rx_control[5], w_hssi_10g_rx_pcs_rx_control[4], w_hssi_10g_rx_pcs_rx_control[3], w_hssi_10g_rx_pcs_rx_control[2], w_hssi_10g_rx_pcs_rx_control[1], w_hssi_10g_rx_pcs_rx_control[0]}),
				.int_pldif_10g_rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.int_pldif_10g_rx_data({w_hssi_10g_rx_pcs_rx_data[127], w_hssi_10g_rx_pcs_rx_data[126], w_hssi_10g_rx_pcs_rx_data[125], w_hssi_10g_rx_pcs_rx_data[124], w_hssi_10g_rx_pcs_rx_data[123], w_hssi_10g_rx_pcs_rx_data[122], w_hssi_10g_rx_pcs_rx_data[121], w_hssi_10g_rx_pcs_rx_data[120], w_hssi_10g_rx_pcs_rx_data[119], w_hssi_10g_rx_pcs_rx_data[118], w_hssi_10g_rx_pcs_rx_data[117], w_hssi_10g_rx_pcs_rx_data[116], w_hssi_10g_rx_pcs_rx_data[115], w_hssi_10g_rx_pcs_rx_data[114], w_hssi_10g_rx_pcs_rx_data[113], w_hssi_10g_rx_pcs_rx_data[112], w_hssi_10g_rx_pcs_rx_data[111], w_hssi_10g_rx_pcs_rx_data[110], w_hssi_10g_rx_pcs_rx_data[109], w_hssi_10g_rx_pcs_rx_data[108], w_hssi_10g_rx_pcs_rx_data[107], w_hssi_10g_rx_pcs_rx_data[106], w_hssi_10g_rx_pcs_rx_data[105], w_hssi_10g_rx_pcs_rx_data[104], w_hssi_10g_rx_pcs_rx_data[103], w_hssi_10g_rx_pcs_rx_data[102], w_hssi_10g_rx_pcs_rx_data[101], w_hssi_10g_rx_pcs_rx_data[100], w_hssi_10g_rx_pcs_rx_data[99], w_hssi_10g_rx_pcs_rx_data[98], w_hssi_10g_rx_pcs_rx_data[97], w_hssi_10g_rx_pcs_rx_data[96], w_hssi_10g_rx_pcs_rx_data[95], w_hssi_10g_rx_pcs_rx_data[94], w_hssi_10g_rx_pcs_rx_data[93], w_hssi_10g_rx_pcs_rx_data[92], w_hssi_10g_rx_pcs_rx_data[91], w_hssi_10g_rx_pcs_rx_data[90], w_hssi_10g_rx_pcs_rx_data[89], w_hssi_10g_rx_pcs_rx_data[88], w_hssi_10g_rx_pcs_rx_data[87], w_hssi_10g_rx_pcs_rx_data[86], w_hssi_10g_rx_pcs_rx_data[85], w_hssi_10g_rx_pcs_rx_data[84], w_hssi_10g_rx_pcs_rx_data[83], w_hssi_10g_rx_pcs_rx_data[82], w_hssi_10g_rx_pcs_rx_data[81], w_hssi_10g_rx_pcs_rx_data[80], w_hssi_10g_rx_pcs_rx_data[79], w_hssi_10g_rx_pcs_rx_data[78], w_hssi_10g_rx_pcs_rx_data[77], w_hssi_10g_rx_pcs_rx_data[76], w_hssi_10g_rx_pcs_rx_data[75], w_hssi_10g_rx_pcs_rx_data[74], w_hssi_10g_rx_pcs_rx_data[73], w_hssi_10g_rx_pcs_rx_data[72], w_hssi_10g_rx_pcs_rx_data[71], w_hssi_10g_rx_pcs_rx_data[70], w_hssi_10g_rx_pcs_rx_data[69], w_hssi_10g_rx_pcs_rx_data[68], w_hssi_10g_rx_pcs_rx_data[67], w_hssi_10g_rx_pcs_rx_data[66], w_hssi_10g_rx_pcs_rx_data[65], w_hssi_10g_rx_pcs_rx_data[64], w_hssi_10g_rx_pcs_rx_data[63], w_hssi_10g_rx_pcs_rx_data[62], w_hssi_10g_rx_pcs_rx_data[61], w_hssi_10g_rx_pcs_rx_data[60], w_hssi_10g_rx_pcs_rx_data[59], w_hssi_10g_rx_pcs_rx_data[58], w_hssi_10g_rx_pcs_rx_data[57], w_hssi_10g_rx_pcs_rx_data[56], w_hssi_10g_rx_pcs_rx_data[55], w_hssi_10g_rx_pcs_rx_data[54], w_hssi_10g_rx_pcs_rx_data[53], w_hssi_10g_rx_pcs_rx_data[52], w_hssi_10g_rx_pcs_rx_data[51], w_hssi_10g_rx_pcs_rx_data[50], w_hssi_10g_rx_pcs_rx_data[49], w_hssi_10g_rx_pcs_rx_data[48], w_hssi_10g_rx_pcs_rx_data[47], w_hssi_10g_rx_pcs_rx_data[46], w_hssi_10g_rx_pcs_rx_data[45], w_hssi_10g_rx_pcs_rx_data[44], w_hssi_10g_rx_pcs_rx_data[43], w_hssi_10g_rx_pcs_rx_data[42], w_hssi_10g_rx_pcs_rx_data[41], w_hssi_10g_rx_pcs_rx_data[40], w_hssi_10g_rx_pcs_rx_data[39], w_hssi_10g_rx_pcs_rx_data[38], w_hssi_10g_rx_pcs_rx_data[37], w_hssi_10g_rx_pcs_rx_data[36], w_hssi_10g_rx_pcs_rx_data[35], w_hssi_10g_rx_pcs_rx_data[34], w_hssi_10g_rx_pcs_rx_data[33], w_hssi_10g_rx_pcs_rx_data[32], w_hssi_10g_rx_pcs_rx_data[31], w_hssi_10g_rx_pcs_rx_data[30], w_hssi_10g_rx_pcs_rx_data[29], w_hssi_10g_rx_pcs_rx_data[28], w_hssi_10g_rx_pcs_rx_data[27], w_hssi_10g_rx_pcs_rx_data[26], w_hssi_10g_rx_pcs_rx_data[25], w_hssi_10g_rx_pcs_rx_data[24], w_hssi_10g_rx_pcs_rx_data[23], w_hssi_10g_rx_pcs_rx_data[22], w_hssi_10g_rx_pcs_rx_data[21], w_hssi_10g_rx_pcs_rx_data[20], w_hssi_10g_rx_pcs_rx_data[19], w_hssi_10g_rx_pcs_rx_data[18], w_hssi_10g_rx_pcs_rx_data[17], w_hssi_10g_rx_pcs_rx_data[16], w_hssi_10g_rx_pcs_rx_data[15], w_hssi_10g_rx_pcs_rx_data[14], w_hssi_10g_rx_pcs_rx_data[13], w_hssi_10g_rx_pcs_rx_data[12], w_hssi_10g_rx_pcs_rx_data[11], w_hssi_10g_rx_pcs_rx_data[10], w_hssi_10g_rx_pcs_rx_data[9], w_hssi_10g_rx_pcs_rx_data[8], w_hssi_10g_rx_pcs_rx_data[7], w_hssi_10g_rx_pcs_rx_data[6], w_hssi_10g_rx_pcs_rx_data[5], w_hssi_10g_rx_pcs_rx_data[4], w_hssi_10g_rx_pcs_rx_data[3], w_hssi_10g_rx_pcs_rx_data[2], w_hssi_10g_rx_pcs_rx_data[1], w_hssi_10g_rx_pcs_rx_data[0]}),
				.int_pldif_10g_rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.int_pldif_10g_rx_diag_status({w_hssi_10g_rx_pcs_rx_diag_status[1], w_hssi_10g_rx_pcs_rx_diag_status[0]}),
				.int_pldif_10g_rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.int_pldif_10g_rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.int_pldif_10g_rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.int_pldif_10g_rx_fifo_num({w_hssi_10g_rx_pcs_rx_fifo_num[4], w_hssi_10g_rx_pcs_rx_fifo_num[3], w_hssi_10g_rx_pcs_rx_fifo_num[2], w_hssi_10g_rx_pcs_rx_fifo_num[1], w_hssi_10g_rx_pcs_rx_fifo_num[0]}),
				.int_pldif_10g_rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.int_pldif_10g_rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.int_pldif_10g_rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.int_pldif_10g_rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.int_pldif_10g_rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.int_pldif_10g_rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				.int_pldif_8g_a1a2_k1k2_flag({w_hssi_8g_rx_pcs_a1a2k1k2flag[3], w_hssi_8g_rx_pcs_a1a2k1k2flag[2], w_hssi_8g_rx_pcs_a1a2k1k2flag[1], w_hssi_8g_rx_pcs_a1a2k1k2flag[0]}),
				.int_pldif_8g_empty_rmf(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.int_pldif_8g_empty_rx(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.int_pldif_8g_full_rmf(w_hssi_8g_rx_pcs_rm_fifo_full),
				.int_pldif_8g_full_rx(w_hssi_8g_rx_pcs_pcfifofull),
				.int_pldif_8g_phystatus(w_hssi_8g_rx_pcs_phystatus),
				.int_pldif_8g_rx_blk_start({w_hssi_8g_rx_pcs_rx_blk_start[3], w_hssi_8g_rx_pcs_rx_blk_start[2], w_hssi_8g_rx_pcs_rx_blk_start[1], w_hssi_8g_rx_pcs_rx_blk_start[0]}),
				.int_pldif_8g_rx_clk(w_hssi_8g_rx_pcs_clock_to_pld),
				.int_pldif_8g_rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_8g_rx_data_valid({w_hssi_8g_rx_pcs_rx_data_valid[3], w_hssi_8g_rx_pcs_rx_data_valid[2], w_hssi_8g_rx_pcs_rx_data_valid[1], w_hssi_8g_rx_pcs_rx_data_valid[0]}),
				.int_pldif_8g_rx_rstn_sync2wrfifo(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.int_pldif_8g_rx_sync_hdr({w_hssi_8g_rx_pcs_rx_sync_hdr[1], w_hssi_8g_rx_pcs_rx_sync_hdr[0]}),
				.int_pldif_8g_rxd({w_hssi_8g_rx_pcs_dataout[63], w_hssi_8g_rx_pcs_dataout[62], w_hssi_8g_rx_pcs_dataout[61], w_hssi_8g_rx_pcs_dataout[60], w_hssi_8g_rx_pcs_dataout[59], w_hssi_8g_rx_pcs_dataout[58], w_hssi_8g_rx_pcs_dataout[57], w_hssi_8g_rx_pcs_dataout[56], w_hssi_8g_rx_pcs_dataout[55], w_hssi_8g_rx_pcs_dataout[54], w_hssi_8g_rx_pcs_dataout[53], w_hssi_8g_rx_pcs_dataout[52], w_hssi_8g_rx_pcs_dataout[51], w_hssi_8g_rx_pcs_dataout[50], w_hssi_8g_rx_pcs_dataout[49], w_hssi_8g_rx_pcs_dataout[48], w_hssi_8g_rx_pcs_dataout[47], w_hssi_8g_rx_pcs_dataout[46], w_hssi_8g_rx_pcs_dataout[45], w_hssi_8g_rx_pcs_dataout[44], w_hssi_8g_rx_pcs_dataout[43], w_hssi_8g_rx_pcs_dataout[42], w_hssi_8g_rx_pcs_dataout[41], w_hssi_8g_rx_pcs_dataout[40], w_hssi_8g_rx_pcs_dataout[39], w_hssi_8g_rx_pcs_dataout[38], w_hssi_8g_rx_pcs_dataout[37], w_hssi_8g_rx_pcs_dataout[36], w_hssi_8g_rx_pcs_dataout[35], w_hssi_8g_rx_pcs_dataout[34], w_hssi_8g_rx_pcs_dataout[33], w_hssi_8g_rx_pcs_dataout[32], w_hssi_8g_rx_pcs_dataout[31], w_hssi_8g_rx_pcs_dataout[30], w_hssi_8g_rx_pcs_dataout[29], w_hssi_8g_rx_pcs_dataout[28], w_hssi_8g_rx_pcs_dataout[27], w_hssi_8g_rx_pcs_dataout[26], w_hssi_8g_rx_pcs_dataout[25], w_hssi_8g_rx_pcs_dataout[24], w_hssi_8g_rx_pcs_dataout[23], w_hssi_8g_rx_pcs_dataout[22], w_hssi_8g_rx_pcs_dataout[21], w_hssi_8g_rx_pcs_dataout[20], w_hssi_8g_rx_pcs_dataout[19], w_hssi_8g_rx_pcs_dataout[18], w_hssi_8g_rx_pcs_dataout[17], w_hssi_8g_rx_pcs_dataout[16], w_hssi_8g_rx_pcs_dataout[15], w_hssi_8g_rx_pcs_dataout[14], w_hssi_8g_rx_pcs_dataout[13], w_hssi_8g_rx_pcs_dataout[12], w_hssi_8g_rx_pcs_dataout[11], w_hssi_8g_rx_pcs_dataout[10], w_hssi_8g_rx_pcs_dataout[9], w_hssi_8g_rx_pcs_dataout[8], w_hssi_8g_rx_pcs_dataout[7], w_hssi_8g_rx_pcs_dataout[6], w_hssi_8g_rx_pcs_dataout[5], w_hssi_8g_rx_pcs_dataout[4], w_hssi_8g_rx_pcs_dataout[3], w_hssi_8g_rx_pcs_dataout[2], w_hssi_8g_rx_pcs_dataout[1], w_hssi_8g_rx_pcs_dataout[0]}),
				.int_pldif_8g_rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.int_pldif_8g_rxstatus({w_hssi_8g_rx_pcs_rxstatus[2], w_hssi_8g_rx_pcs_rxstatus[1], w_hssi_8g_rx_pcs_rxstatus[0]}),
				.int_pldif_8g_rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.int_pldif_8g_signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.int_pldif_8g_wa_boundary({w_hssi_8g_rx_pcs_word_align_boundary[4], w_hssi_8g_rx_pcs_word_align_boundary[3], w_hssi_8g_rx_pcs_word_align_boundary[2], w_hssi_8g_rx_pcs_word_align_boundary[1], w_hssi_8g_rx_pcs_word_align_boundary[0]}),
				.int_pldif_krfec_rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.int_pldif_krfec_rx_data_status({w_hssi_krfec_rx_pcs_rx_data_status[1], w_hssi_krfec_rx_pcs_rx_data_status[0]}),
				.int_pldif_krfec_rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.int_pldif_pmaif_clkdiv_rx(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pldif_pmaif_clkdiv_rx_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pldif_pmaif_rx_data({w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0]}),
				.int_pldif_pmaif_rx_prbs_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pldif_pmaif_rx_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.pld_10g_krfec_rx_clr_errblk_cnt(in_pld_10g_krfec_rx_clr_errblk_cnt),
				.pld_10g_krfec_rx_pld_rst_n(in_pld_10g_krfec_rx_pld_rst_n),
				.pld_10g_rx_align_clr(in_pld_10g_rx_align_clr),
				.pld_10g_rx_clr_ber_count(in_pld_10g_rx_clr_ber_count),
				.pld_10g_rx_rd_en(in_pld_10g_rx_rd_en),
				.pld_8g_a1a2_size(in_pld_8g_a1a2_size),
				.pld_8g_bitloc_rev_en(in_pld_8g_bitloc_rev_en),
				.pld_8g_byte_rev_en(in_pld_8g_byte_rev_en),
				.pld_8g_encdt(in_pld_8g_encdt),
				.pld_8g_g3_rx_pld_rst_n(in_pld_8g_g3_rx_pld_rst_n),
				.pld_8g_rdenable_rx(in_pld_8g_rdenable_rx),
				.pld_8g_rxpolarity(in_pld_8g_rxpolarity),
				.pld_8g_wrdisable_rx(in_pld_8g_wrdisable_rx),
				.pld_bitslip(in_pld_bitslip),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_rxpma_rstb(in_pld_pma_rxpma_rstb),
				.pld_pmaif_rx_pld_rst_n(in_pld_pmaif_rx_pld_rst_n),
				.pld_pmaif_rxclkslip(in_pld_pmaif_rxclkslip),
				.pld_polinv_rx(in_pld_polinv_rx),
				.pld_rx_clk(in_pld_rx_clk),
				.pld_rx_prbs_err_clr(in_pld_rx_prbs_err_clr),
				.pld_syncsm_en(in_pld_syncsm_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.int_pldif_pmaif_rx_pld_clk(),
				.pld_8g_wa_boundary_txclk_fastreg(),
				.pld_8g_wa_boundary_txclk_reg(),
				.pld_bitslip_10g_txclk_reg(),
				.pld_bitslip_8g_txclk_reg(),
				.pld_bitslip_rxclk_parallel_loopback_reg(),
				.pld_bitslip_rxclk_reg(),
				.pld_pcs_rx_clk_out_pcsdirect_wire(),
				.pld_pma_rx_clk_out_10g_or_pcsdirect_wire(),
				.pld_pma_rx_clk_out_8g_wire(),
				.pld_pmaif_rx_pld_rst_n_reg(),
				.pld_pmaif_tx_pld_rst_n_txclk_reg(),
				.pld_polinv_rx_reg(),
				.pld_rx_clk_fifo(),
				.pld_rx_control_fifo(),
				.pld_rx_control_pcsdirect_reg(),
				.pld_rx_data_fifo(),
				.pld_rx_data_pcsdirect_reg(),
				.pld_rx_prbs_done_reg(),
				.pld_rx_prbs_done_txclk_reg(),
				.pld_rx_prbs_err_clr_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_clr_reg(),
				.pld_rx_prbs_err_disprbs_reg(),
				.pld_rx_prbs_err_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_reg(),
				.pma_rx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_data[50:0] = 51'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3:0] = 4'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_control[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_data[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pcs_pma_interface
			twentynm_hssi_tx_pcs_pma_interface #(
				.bypass_pma_txelecidle(hssi_tx_pcs_pma_interface_bypass_pma_txelecidle),
				.channel_operation_mode(hssi_tx_pcs_pma_interface_channel_operation_mode),
				.lpbk_en(hssi_tx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_tx_pcs_pma_interface_master_clk_sel),
				.pcie_sub_prot_mode_tx(hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx),
				.pldif_datawidth_mode(hssi_tx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_tx(hssi_tx_pcs_pma_interface_pma_dw_tx),
				.pma_if_dft_en(hssi_tx_pcs_pma_interface_pma_if_dft_en),
				.pmagate_en(hssi_tx_pcs_pma_interface_pmagate_en),
				.prbs9_dwidth(hssi_tx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_tx_pcs_pma_interface_prbs_clken),
				.prbs_gen_pat(hssi_tx_pcs_pma_interface_prbs_gen_pat),
				.prot_mode_tx(hssi_tx_pcs_pma_interface_prot_mode_tx),
				.reconfig_settings(hssi_tx_pcs_pma_interface_reconfig_settings),
				.silicon_rev( "20nm5" ),       //PARAM_HIDE
				.sq_wave_num(hssi_tx_pcs_pma_interface_sq_wave_num),
				.sqwgen_clken(hssi_tx_pcs_pma_interface_sqwgen_clken),
				.sup_mode(hssi_tx_pcs_pma_interface_sup_mode),
				.tx_dyn_polarity_inversion(hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion),
				.tx_pma_data_sel(hssi_tx_pcs_pma_interface_tx_pma_data_sel),
				.tx_static_polarity_inversion(hssi_tx_pcs_pma_interface_tx_static_polarity_inversion),
				.uhsif_cnt_step_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock),
				.uhsif_cnt_thresh_filt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value),
				.uhsif_cnt_thresh_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock),
				.uhsif_dcn_test_update_period(hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period),
				.uhsif_dcn_testmode_enable(hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable),
				.uhsif_dead_zone_count_thresh(hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh),
				.uhsif_dead_zone_detection_enable(hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable),
				.uhsif_dead_zone_obser_window(hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window),
				.uhsif_dead_zone_skip_size(hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size),
				.uhsif_delay_cell_index_sel(hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel),
				.uhsif_delay_cell_margin(hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin),
				.uhsif_delay_cell_static_index_value(hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value),
				.uhsif_dft_dead_zone_control(hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control),
				.uhsif_dft_up_filt_control(hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control),
				.uhsif_enable(hssi_tx_pcs_pma_interface_uhsif_enable),
				.uhsif_lock_det_segsz_after_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock),
				.uhsif_lock_det_segsz_before_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock),
				.uhsif_lock_det_thresh_cnt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value),
				.uhsif_lock_det_thresh_cnt_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value),
				.uhsif_lock_det_thresh_diff_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value),
				.uhsif_lock_det_thresh_diff_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value)
			) inst_twentynm_hssi_tx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.int_pmaif_8g_txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.int_pmaif_pldif_tx_clkdiv(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pmaif_pldif_tx_clkdiv_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pmaif_pldif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.int_pmaif_pldif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.int_tx_dft_obsrv_clk(w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk),
				.pma_tx_elec_idle(w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle),
				.pma_tx_pma_data(w_hssi_tx_pcs_pma_interface_pma_tx_pma_data),
				.pma_txpma_rstb(w_hssi_tx_pcs_pma_interface_pma_txpma_rstb),
				.tx_pma_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback),
				.tx_pma_uhsif_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback),
				.tx_prbs_gen_test(w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test),
				.uhsif_test_out_1(w_hssi_tx_pcs_pma_interface_uhsif_test_out_1),
				.uhsif_test_out_2(w_hssi_tx_pcs_pma_interface_uhsif_test_out_2),
				.uhsif_test_out_3(w_hssi_tx_pcs_pma_interface_uhsif_test_out_3),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.int_pmaif_10g_tx_pma_data({w_hssi_10g_tx_pcs_tx_pma_data[63], w_hssi_10g_tx_pcs_tx_pma_data[62], w_hssi_10g_tx_pcs_tx_pma_data[61], w_hssi_10g_tx_pcs_tx_pma_data[60], w_hssi_10g_tx_pcs_tx_pma_data[59], w_hssi_10g_tx_pcs_tx_pma_data[58], w_hssi_10g_tx_pcs_tx_pma_data[57], w_hssi_10g_tx_pcs_tx_pma_data[56], w_hssi_10g_tx_pcs_tx_pma_data[55], w_hssi_10g_tx_pcs_tx_pma_data[54], w_hssi_10g_tx_pcs_tx_pma_data[53], w_hssi_10g_tx_pcs_tx_pma_data[52], w_hssi_10g_tx_pcs_tx_pma_data[51], w_hssi_10g_tx_pcs_tx_pma_data[50], w_hssi_10g_tx_pcs_tx_pma_data[49], w_hssi_10g_tx_pcs_tx_pma_data[48], w_hssi_10g_tx_pcs_tx_pma_data[47], w_hssi_10g_tx_pcs_tx_pma_data[46], w_hssi_10g_tx_pcs_tx_pma_data[45], w_hssi_10g_tx_pcs_tx_pma_data[44], w_hssi_10g_tx_pcs_tx_pma_data[43], w_hssi_10g_tx_pcs_tx_pma_data[42], w_hssi_10g_tx_pcs_tx_pma_data[41], w_hssi_10g_tx_pcs_tx_pma_data[40], w_hssi_10g_tx_pcs_tx_pma_data[39], w_hssi_10g_tx_pcs_tx_pma_data[38], w_hssi_10g_tx_pcs_tx_pma_data[37], w_hssi_10g_tx_pcs_tx_pma_data[36], w_hssi_10g_tx_pcs_tx_pma_data[35], w_hssi_10g_tx_pcs_tx_pma_data[34], w_hssi_10g_tx_pcs_tx_pma_data[33], w_hssi_10g_tx_pcs_tx_pma_data[32], w_hssi_10g_tx_pcs_tx_pma_data[31], w_hssi_10g_tx_pcs_tx_pma_data[30], w_hssi_10g_tx_pcs_tx_pma_data[29], w_hssi_10g_tx_pcs_tx_pma_data[28], w_hssi_10g_tx_pcs_tx_pma_data[27], w_hssi_10g_tx_pcs_tx_pma_data[26], w_hssi_10g_tx_pcs_tx_pma_data[25], w_hssi_10g_tx_pcs_tx_pma_data[24], w_hssi_10g_tx_pcs_tx_pma_data[23], w_hssi_10g_tx_pcs_tx_pma_data[22], w_hssi_10g_tx_pcs_tx_pma_data[21], w_hssi_10g_tx_pcs_tx_pma_data[20], w_hssi_10g_tx_pcs_tx_pma_data[19], w_hssi_10g_tx_pcs_tx_pma_data[18], w_hssi_10g_tx_pcs_tx_pma_data[17], w_hssi_10g_tx_pcs_tx_pma_data[16], w_hssi_10g_tx_pcs_tx_pma_data[15], w_hssi_10g_tx_pcs_tx_pma_data[14], w_hssi_10g_tx_pcs_tx_pma_data[13], w_hssi_10g_tx_pcs_tx_pma_data[12], w_hssi_10g_tx_pcs_tx_pma_data[11], w_hssi_10g_tx_pcs_tx_pma_data[10], w_hssi_10g_tx_pcs_tx_pma_data[9], w_hssi_10g_tx_pcs_tx_pma_data[8], w_hssi_10g_tx_pcs_tx_pma_data[7], w_hssi_10g_tx_pcs_tx_pma_data[6], w_hssi_10g_tx_pcs_tx_pma_data[5], w_hssi_10g_tx_pcs_tx_pma_data[4], w_hssi_10g_tx_pcs_tx_pma_data[3], w_hssi_10g_tx_pcs_tx_pma_data[2], w_hssi_10g_tx_pcs_tx_pma_data[1], w_hssi_10g_tx_pcs_tx_pma_data[0]}),
				.int_pmaif_10g_tx_pma_data_gate_val({w_hssi_10g_tx_pcs_tx_pma_gating_val[63], w_hssi_10g_tx_pcs_tx_pma_gating_val[62], w_hssi_10g_tx_pcs_tx_pma_gating_val[61], w_hssi_10g_tx_pcs_tx_pma_gating_val[60], w_hssi_10g_tx_pcs_tx_pma_gating_val[59], w_hssi_10g_tx_pcs_tx_pma_gating_val[58], w_hssi_10g_tx_pcs_tx_pma_gating_val[57], w_hssi_10g_tx_pcs_tx_pma_gating_val[56], w_hssi_10g_tx_pcs_tx_pma_gating_val[55], w_hssi_10g_tx_pcs_tx_pma_gating_val[54], w_hssi_10g_tx_pcs_tx_pma_gating_val[53], w_hssi_10g_tx_pcs_tx_pma_gating_val[52], w_hssi_10g_tx_pcs_tx_pma_gating_val[51], w_hssi_10g_tx_pcs_tx_pma_gating_val[50], w_hssi_10g_tx_pcs_tx_pma_gating_val[49], w_hssi_10g_tx_pcs_tx_pma_gating_val[48], w_hssi_10g_tx_pcs_tx_pma_gating_val[47], w_hssi_10g_tx_pcs_tx_pma_gating_val[46], w_hssi_10g_tx_pcs_tx_pma_gating_val[45], w_hssi_10g_tx_pcs_tx_pma_gating_val[44], w_hssi_10g_tx_pcs_tx_pma_gating_val[43], w_hssi_10g_tx_pcs_tx_pma_gating_val[42], w_hssi_10g_tx_pcs_tx_pma_gating_val[41], w_hssi_10g_tx_pcs_tx_pma_gating_val[40], w_hssi_10g_tx_pcs_tx_pma_gating_val[39], w_hssi_10g_tx_pcs_tx_pma_gating_val[38], w_hssi_10g_tx_pcs_tx_pma_gating_val[37], w_hssi_10g_tx_pcs_tx_pma_gating_val[36], w_hssi_10g_tx_pcs_tx_pma_gating_val[35], w_hssi_10g_tx_pcs_tx_pma_gating_val[34], w_hssi_10g_tx_pcs_tx_pma_gating_val[33], w_hssi_10g_tx_pcs_tx_pma_gating_val[32], w_hssi_10g_tx_pcs_tx_pma_gating_val[31], w_hssi_10g_tx_pcs_tx_pma_gating_val[30], w_hssi_10g_tx_pcs_tx_pma_gating_val[29], w_hssi_10g_tx_pcs_tx_pma_gating_val[28], w_hssi_10g_tx_pcs_tx_pma_gating_val[27], w_hssi_10g_tx_pcs_tx_pma_gating_val[26], w_hssi_10g_tx_pcs_tx_pma_gating_val[25], w_hssi_10g_tx_pcs_tx_pma_gating_val[24], w_hssi_10g_tx_pcs_tx_pma_gating_val[23], w_hssi_10g_tx_pcs_tx_pma_gating_val[22], w_hssi_10g_tx_pcs_tx_pma_gating_val[21], w_hssi_10g_tx_pcs_tx_pma_gating_val[20], w_hssi_10g_tx_pcs_tx_pma_gating_val[19], w_hssi_10g_tx_pcs_tx_pma_gating_val[18], w_hssi_10g_tx_pcs_tx_pma_gating_val[17], w_hssi_10g_tx_pcs_tx_pma_gating_val[16], w_hssi_10g_tx_pcs_tx_pma_gating_val[15], w_hssi_10g_tx_pcs_tx_pma_gating_val[14], w_hssi_10g_tx_pcs_tx_pma_gating_val[13], w_hssi_10g_tx_pcs_tx_pma_gating_val[12], w_hssi_10g_tx_pcs_tx_pma_gating_val[11], w_hssi_10g_tx_pcs_tx_pma_gating_val[10], w_hssi_10g_tx_pcs_tx_pma_gating_val[9], w_hssi_10g_tx_pcs_tx_pma_gating_val[8], w_hssi_10g_tx_pcs_tx_pma_gating_val[7], w_hssi_10g_tx_pcs_tx_pma_gating_val[6], w_hssi_10g_tx_pcs_tx_pma_gating_val[5], w_hssi_10g_tx_pcs_tx_pma_gating_val[4], w_hssi_10g_tx_pcs_tx_pma_gating_val[3], w_hssi_10g_tx_pcs_tx_pma_gating_val[2], w_hssi_10g_tx_pcs_tx_pma_gating_val[1], w_hssi_10g_tx_pcs_tx_pma_gating_val[0]}),
				.int_pmaif_8g_pudr({w_hssi_8g_tx_pcs_dataout[19], w_hssi_8g_tx_pcs_dataout[18], w_hssi_8g_tx_pcs_dataout[17], w_hssi_8g_tx_pcs_dataout[16], w_hssi_8g_tx_pcs_dataout[15], w_hssi_8g_tx_pcs_dataout[14], w_hssi_8g_tx_pcs_dataout[13], w_hssi_8g_tx_pcs_dataout[12], w_hssi_8g_tx_pcs_dataout[11], w_hssi_8g_tx_pcs_dataout[10], w_hssi_8g_tx_pcs_dataout[9], w_hssi_8g_tx_pcs_dataout[8], w_hssi_8g_tx_pcs_dataout[7], w_hssi_8g_tx_pcs_dataout[6], w_hssi_8g_tx_pcs_dataout[5], w_hssi_8g_tx_pcs_dataout[4], w_hssi_8g_tx_pcs_dataout[3], w_hssi_8g_tx_pcs_dataout[2], w_hssi_8g_tx_pcs_dataout[1], w_hssi_8g_tx_pcs_dataout[0]}),
				.int_pmaif_8g_tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.int_pmaif_8g_tx_elec_idle(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_pma_data_out({w_hssi_gen3_tx_pcs_data_out[31], w_hssi_gen3_tx_pcs_data_out[30], w_hssi_gen3_tx_pcs_data_out[29], w_hssi_gen3_tx_pcs_data_out[28], w_hssi_gen3_tx_pcs_data_out[27], w_hssi_gen3_tx_pcs_data_out[26], w_hssi_gen3_tx_pcs_data_out[25], w_hssi_gen3_tx_pcs_data_out[24], w_hssi_gen3_tx_pcs_data_out[23], w_hssi_gen3_tx_pcs_data_out[22], w_hssi_gen3_tx_pcs_data_out[21], w_hssi_gen3_tx_pcs_data_out[20], w_hssi_gen3_tx_pcs_data_out[19], w_hssi_gen3_tx_pcs_data_out[18], w_hssi_gen3_tx_pcs_data_out[17], w_hssi_gen3_tx_pcs_data_out[16], w_hssi_gen3_tx_pcs_data_out[15], w_hssi_gen3_tx_pcs_data_out[14], w_hssi_gen3_tx_pcs_data_out[13], w_hssi_gen3_tx_pcs_data_out[12], w_hssi_gen3_tx_pcs_data_out[11], w_hssi_gen3_tx_pcs_data_out[10], w_hssi_gen3_tx_pcs_data_out[9], w_hssi_gen3_tx_pcs_data_out[8], w_hssi_gen3_tx_pcs_data_out[7], w_hssi_gen3_tx_pcs_data_out[6], w_hssi_gen3_tx_pcs_data_out[5], w_hssi_gen3_tx_pcs_data_out[4], w_hssi_gen3_tx_pcs_data_out[3], w_hssi_gen3_tx_pcs_data_out[2], w_hssi_gen3_tx_pcs_data_out[1], w_hssi_gen3_tx_pcs_data_out[0]}),
				.int_pmaif_g3_pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.int_pmaif_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pmaif_pldif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pmaif_pldif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0]}),
				.int_pmaif_pldif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pmaif_pldif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.int_pmaif_pldif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pmaif_pldif_uhsif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0]}),
				.pma_tx_clkdiv_user(in_pma_tx_clkdiv_user),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.refclk_dig_uhsif(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.uhsif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.uhsif_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				
				// UNUSED
				.avmm_user_dataout(),
				.write_en(),
				.write_en_ack()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4:0] = 5'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_txpma_rstb = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pld_pcs_interface
			twentynm_hssi_tx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx),
				.hd_10g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx),
				.hd_10g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx),
				.hd_10g_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx),
				.hd_10g_lpbk_en(hssi_tx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx),
				.hd_10g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx),
				.hd_10g_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx),
				.hd_8g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx),
				.hd_8g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx),
				.hd_8g_hip_mode(hssi_tx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_tx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx),
				.hd_8g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx),
				.hd_chnl_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx),
				.hd_chnl_frequency_rules_en(hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_tx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_tx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx),
				.hd_chnl_lpbk_en(hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx),
				.hd_chnl_pld_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz),
				.hd_chnl_pld_uhsif_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz),
				.hd_chnl_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx),
				.hd_chnl_pma_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz),
				.hd_chnl_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx),
				.hd_chnl_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx),
				.hd_fifo_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx),
				.hd_fifo_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx),
				.hd_g3_prot_mode(hssi_tx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx),
				.hd_krfec_lpbk_en(hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx),
				.hd_pldif_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx),
				.hd_pmaif_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_ctrl_plane_bonding(hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding),
				.hd_pmaif_lpbk_en(hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx),
				.hd_pmaif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx),
				.hd_pmaif_sim_mode(hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_tx_clk_out_sel(hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel),
				.pcs_tx_clk_source(hssi_tx_pld_pcs_interface_pcs_tx_clk_source),
				.pcs_tx_data_source(hssi_tx_pld_pcs_interface_pcs_tx_data_source),
				.pcs_tx_delay1_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en),
				.pcs_tx_delay1_clk_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel),
				.pcs_tx_delay1_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl),
				.pcs_tx_delay1_data_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel),
				.pcs_tx_delay2_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en),
				.pcs_tx_delay2_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl),
				.pcs_tx_output_sel(hssi_tx_pld_pcs_interface_pcs_tx_output_sel),
				.reconfig_settings(hssi_tx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm5" )       //PARAM_HIDE
			) inst_twentynm_hssi_tx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pld_pcs_interface_blockselect),
				.hip_tx_clk(w_hssi_tx_pld_pcs_interface_hip_tx_clk),
				.int_pldif_10g_tx_bitslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip),
				.int_pldif_10g_tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.int_pldif_10g_tx_control(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control),
				.int_pldif_10g_tx_control_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg),
				.int_pldif_10g_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data),
				.int_pldif_10g_tx_data_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg),
				.int_pldif_10g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.int_pldif_10g_tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.int_pldif_10g_tx_diag_status(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status),
				.int_pldif_10g_tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.int_pldif_10g_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.int_pldif_10g_tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				.int_pldif_8g_pld_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.int_pldif_8g_powerdown(w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown),
				.int_pldif_8g_rddisable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.int_pldif_8g_rev_loopbk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.int_pldif_8g_tx_blk_start(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start),
				.int_pldif_8g_tx_boundary_sel(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel),
				.int_pldif_8g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid),
				.int_pldif_8g_tx_sync_hdr(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr),
				.int_pldif_8g_txd(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd),
				.int_pldif_8g_txd_fast_reg(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg),
				.int_pldif_8g_txdeemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.int_pldif_8g_txdetectrxloopback(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.int_pldif_8g_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.int_pldif_8g_txmargin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin),
				.int_pldif_8g_txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.int_pldif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.int_pldif_8g_wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				.int_pldif_pmaif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pldif_pmaif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pldif_pmaif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data),
				.int_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pldif_pmaif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pldif_pmaif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pldif_pmaif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pldif_pmaif_uhsif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data),
				.pld_10g_krfec_tx_frame(w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame),
				.pld_10g_tx_burst_en_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe),
				.pld_10g_tx_empty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty),
				.pld_10g_tx_fifo_num(w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num),
				.pld_10g_tx_full(w_hssi_tx_pld_pcs_interface_pld_10g_tx_full),
				.pld_10g_tx_pempty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty),
				.pld_10g_tx_pfull(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull),
				.pld_10g_tx_wordslip_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe),
				.pld_8g_empty_tx(w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx),
				.pld_8g_full_tx(w_hssi_tx_pld_pcs_interface_pld_8g_full_tx),
				.pld_krfec_tx_alignment(w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment),
				.pld_pcs_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out),
				.pld_pma_clkdiv_tx_user(w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user),
				.pld_pma_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out),
				.pld_uhsif_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.hip_tx_data({in_hip_tx_data[63], in_hip_tx_data[62], in_hip_tx_data[61], in_hip_tx_data[60], in_hip_tx_data[59], in_hip_tx_data[58], in_hip_tx_data[57], in_hip_tx_data[56], in_hip_tx_data[55], in_hip_tx_data[54], in_hip_tx_data[53], in_hip_tx_data[52], in_hip_tx_data[51], in_hip_tx_data[50], in_hip_tx_data[49], in_hip_tx_data[48], in_hip_tx_data[47], in_hip_tx_data[46], in_hip_tx_data[45], in_hip_tx_data[44], in_hip_tx_data[43], in_hip_tx_data[42], in_hip_tx_data[41], in_hip_tx_data[40], in_hip_tx_data[39], in_hip_tx_data[38], in_hip_tx_data[37], in_hip_tx_data[36], in_hip_tx_data[35], in_hip_tx_data[34], in_hip_tx_data[33], in_hip_tx_data[32], in_hip_tx_data[31], in_hip_tx_data[30], in_hip_tx_data[29], in_hip_tx_data[28], in_hip_tx_data[27], in_hip_tx_data[26], in_hip_tx_data[25], in_hip_tx_data[24], in_hip_tx_data[23], in_hip_tx_data[22], in_hip_tx_data[21], in_hip_tx_data[20], in_hip_tx_data[19], in_hip_tx_data[18], in_hip_tx_data[17], in_hip_tx_data[16], in_hip_tx_data[15], in_hip_tx_data[14], in_hip_tx_data[13], in_hip_tx_data[12], in_hip_tx_data[11], in_hip_tx_data[10], in_hip_tx_data[9], in_hip_tx_data[8], in_hip_tx_data[7], in_hip_tx_data[6], in_hip_tx_data[5], in_hip_tx_data[4], in_hip_tx_data[3], in_hip_tx_data[2], in_hip_tx_data[1], in_hip_tx_data[0]}),
				.int_pldif_10g_tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.int_pldif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.int_pldif_10g_tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_10g_tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.int_pldif_10g_tx_fifo_num({w_hssi_10g_tx_pcs_tx_fifo_num[3], w_hssi_10g_tx_pcs_tx_fifo_num[2], w_hssi_10g_tx_pcs_tx_fifo_num[1], w_hssi_10g_tx_pcs_tx_fifo_num[0]}),
				.int_pldif_10g_tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.int_pldif_10g_tx_full(w_hssi_10g_tx_pcs_tx_full),
				.int_pldif_10g_tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.int_pldif_10g_tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.int_pldif_10g_tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				.int_pldif_8g_empty_tx(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.int_pldif_8g_full_tx(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.int_pldif_8g_tx_clk_out(w_hssi_8g_tx_pcs_clk_out),
				.int_pldif_8g_tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_krfec_tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.int_pldif_krfec_tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.int_pldif_pmaif_clkdiv_tx(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pldif_pmaif_clkdiv_tx_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pldif_pmaif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.pld_10g_krfec_tx_pld_rst_n(in_pld_10g_krfec_tx_pld_rst_n),
				.pld_10g_tx_bitslip({in_pld_10g_tx_bitslip[6], in_pld_10g_tx_bitslip[5], in_pld_10g_tx_bitslip[4], in_pld_10g_tx_bitslip[3], in_pld_10g_tx_bitslip[2], in_pld_10g_tx_bitslip[1], in_pld_10g_tx_bitslip[0]}),
				.pld_10g_tx_burst_en(in_pld_10g_tx_burst_en),
				.pld_10g_tx_data_valid(in_pld_10g_tx_data_valid),
				.pld_10g_tx_diag_status({in_pld_10g_tx_diag_status[1], in_pld_10g_tx_diag_status[0]}),
				.pld_10g_tx_wordslip(in_pld_10g_tx_wordslip),
				.pld_8g_g3_tx_pld_rst_n(in_pld_8g_g3_tx_pld_rst_n),
				.pld_8g_rddisable_tx(in_pld_8g_rddisable_tx),
				.pld_8g_tx_boundary_sel({in_pld_8g_tx_boundary_sel[4], in_pld_8g_tx_boundary_sel[3], in_pld_8g_tx_boundary_sel[2], in_pld_8g_tx_boundary_sel[1], in_pld_8g_tx_boundary_sel[0]}),
				.pld_8g_wrenable_tx(in_pld_8g_wrenable_tx),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_txpma_rstb(in_pld_pma_txpma_rstb),
				.pld_pmaif_tx_pld_rst_n(in_pld_pmaif_tx_pld_rst_n),
				.pld_polinv_tx(in_pld_polinv_tx),
				.pld_tx_clk(in_pld_tx_clk),
				.pld_tx_control({in_pld_tx_control[17], in_pld_tx_control[16], in_pld_tx_control[15], in_pld_tx_control[14], in_pld_tx_control[13], in_pld_tx_control[12], in_pld_tx_control[11], in_pld_tx_control[10], in_pld_tx_control[9], in_pld_tx_control[8], in_pld_tx_control[7], in_pld_tx_control[6], in_pld_tx_control[5], in_pld_tx_control[4], in_pld_tx_control[3], in_pld_tx_control[2], in_pld_tx_control[1], in_pld_tx_control[0]}),
				.pld_tx_data({in_pld_tx_data[127], in_pld_tx_data[126], in_pld_tx_data[125], in_pld_tx_data[124], in_pld_tx_data[123], in_pld_tx_data[122], in_pld_tx_data[121], in_pld_tx_data[120], in_pld_tx_data[119], in_pld_tx_data[118], in_pld_tx_data[117], in_pld_tx_data[116], in_pld_tx_data[115], in_pld_tx_data[114], in_pld_tx_data[113], in_pld_tx_data[112], in_pld_tx_data[111], in_pld_tx_data[110], in_pld_tx_data[109], in_pld_tx_data[108], in_pld_tx_data[107], in_pld_tx_data[106], in_pld_tx_data[105], in_pld_tx_data[104], in_pld_tx_data[103], in_pld_tx_data[102], in_pld_tx_data[101], in_pld_tx_data[100], in_pld_tx_data[99], in_pld_tx_data[98], in_pld_tx_data[97], in_pld_tx_data[96], in_pld_tx_data[95], in_pld_tx_data[94], in_pld_tx_data[93], in_pld_tx_data[92], in_pld_tx_data[91], in_pld_tx_data[90], in_pld_tx_data[89], in_pld_tx_data[88], in_pld_tx_data[87], in_pld_tx_data[86], in_pld_tx_data[85], in_pld_tx_data[84], in_pld_tx_data[83], in_pld_tx_data[82], in_pld_tx_data[81], in_pld_tx_data[80], in_pld_tx_data[79], in_pld_tx_data[78], in_pld_tx_data[77], in_pld_tx_data[76], in_pld_tx_data[75], in_pld_tx_data[74], in_pld_tx_data[73], in_pld_tx_data[72], in_pld_tx_data[71], in_pld_tx_data[70], in_pld_tx_data[69], in_pld_tx_data[68], in_pld_tx_data[67], in_pld_tx_data[66], in_pld_tx_data[65], in_pld_tx_data[64], in_pld_tx_data[63], in_pld_tx_data[62], in_pld_tx_data[61], in_pld_tx_data[60], in_pld_tx_data[59], in_pld_tx_data[58], in_pld_tx_data[57], in_pld_tx_data[56], in_pld_tx_data[55], in_pld_tx_data[54], in_pld_tx_data[53], in_pld_tx_data[52], in_pld_tx_data[51], in_pld_tx_data[50], in_pld_tx_data[49], in_pld_tx_data[48], in_pld_tx_data[47], in_pld_tx_data[46], in_pld_tx_data[45], in_pld_tx_data[44], in_pld_tx_data[43], in_pld_tx_data[42], in_pld_tx_data[41], in_pld_tx_data[40], in_pld_tx_data[39], in_pld_tx_data[38], in_pld_tx_data[37], in_pld_tx_data[36], in_pld_tx_data[35], in_pld_tx_data[34], in_pld_tx_data[33], in_pld_tx_data[32], in_pld_tx_data[31], in_pld_tx_data[30], in_pld_tx_data[29], in_pld_tx_data[28], in_pld_tx_data[27], in_pld_tx_data[26], in_pld_tx_data[25], in_pld_tx_data[24], in_pld_tx_data[23], in_pld_tx_data[22], in_pld_tx_data[21], in_pld_tx_data[20], in_pld_tx_data[19], in_pld_tx_data[18], in_pld_tx_data[17], in_pld_tx_data[16], in_pld_tx_data[15], in_pld_tx_data[14], in_pld_tx_data[13], in_pld_tx_data[12], in_pld_tx_data[11], in_pld_tx_data[10], in_pld_tx_data[9], in_pld_tx_data[8], in_pld_tx_data[7], in_pld_tx_data[6], in_pld_tx_data[5], in_pld_tx_data[4], in_pld_tx_data[3], in_pld_tx_data[2], in_pld_tx_data[1], in_pld_tx_data[0]}),
				.pld_txelecidle(in_pld_txelecidle),
				.pld_uhsif_tx_clk(in_pld_uhsif_tx_clk),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.hip_clk_out_div_by_2_wire(),
				.hip_clk_out_wire(),
				.int_pldif_pmaif_tx_pld_clk(),
				.pld_10g_tx_burst_en_exe_10g_fastreg(),
				.pld_10g_tx_burst_en_exe_plddirect_reg(),
				.pld_10g_tx_data_valid_2ff_delay1_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay3_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg(),
				.pld_10g_tx_data_valid_fastreg(),
				.pld_10g_tx_data_valid_plddirect_fastreg(),
				.pld_pcs_tx_clk_out_pma_wire(),
				.pld_pma_tx_clk_out_wire(),
				.pld_pmaif_tx_pld_rst_n_reg(),
				.pld_polinv_tx_10g_pcsdirect_reg(),
				.pld_polinv_tx_8g_reg(),
				.pld_polinv_tx_pat_reg(),
				.pld_tx_clk_fifo(),
				.pld_tx_control_fifo(),
				.pld_tx_control_hi_10g_reg(),
				.pld_tx_control_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_10g_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_8g_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_control_lo_plddirect_fastreg(),
				.pld_tx_control_lo_plddirect_reg(),
				.pld_tx_data_hi_reg(),
				.pld_tx_data_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_10g_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_8g_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_data_lo_plddirect_fastreg(),
				.pld_tx_data_lo_plddirect_reg(),
				.pld_uhsif_reg(),
				.pma_tx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_hip_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6:0] = 7'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17:0] = 18'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8:0] = 9'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127:0] = 128'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4:0] = 5'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2:0] = 3'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_full = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_full_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out = 1'b0;
		end // if not generate
		
		//output assignments
		assign out_avmmreaddata_hssi_10g_rx_pcs = {w_hssi_10g_rx_pcs_avmmreaddata[7], w_hssi_10g_rx_pcs_avmmreaddata[6], w_hssi_10g_rx_pcs_avmmreaddata[5], w_hssi_10g_rx_pcs_avmmreaddata[4], w_hssi_10g_rx_pcs_avmmreaddata[3], w_hssi_10g_rx_pcs_avmmreaddata[2], w_hssi_10g_rx_pcs_avmmreaddata[1], w_hssi_10g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_10g_tx_pcs = {w_hssi_10g_tx_pcs_avmmreaddata[7], w_hssi_10g_tx_pcs_avmmreaddata[6], w_hssi_10g_tx_pcs_avmmreaddata[5], w_hssi_10g_tx_pcs_avmmreaddata[4], w_hssi_10g_tx_pcs_avmmreaddata[3], w_hssi_10g_tx_pcs_avmmreaddata[2], w_hssi_10g_tx_pcs_avmmreaddata[1], w_hssi_10g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_rx_pcs = {w_hssi_8g_rx_pcs_avmmreaddata[7], w_hssi_8g_rx_pcs_avmmreaddata[6], w_hssi_8g_rx_pcs_avmmreaddata[5], w_hssi_8g_rx_pcs_avmmreaddata[4], w_hssi_8g_rx_pcs_avmmreaddata[3], w_hssi_8g_rx_pcs_avmmreaddata[2], w_hssi_8g_rx_pcs_avmmreaddata[1], w_hssi_8g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_tx_pcs = {w_hssi_8g_tx_pcs_avmmreaddata[7], w_hssi_8g_tx_pcs_avmmreaddata[6], w_hssi_8g_tx_pcs_avmmreaddata[5], w_hssi_8g_tx_pcs_avmmreaddata[4], w_hssi_8g_tx_pcs_avmmreaddata[3], w_hssi_8g_tx_pcs_avmmreaddata[2], w_hssi_8g_tx_pcs_avmmreaddata[1], w_hssi_8g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pcs_pma_interface = {w_hssi_common_pcs_pma_interface_avmmreaddata[7], w_hssi_common_pcs_pma_interface_avmmreaddata[6], w_hssi_common_pcs_pma_interface_avmmreaddata[5], w_hssi_common_pcs_pma_interface_avmmreaddata[4], w_hssi_common_pcs_pma_interface_avmmreaddata[3], w_hssi_common_pcs_pma_interface_avmmreaddata[2], w_hssi_common_pcs_pma_interface_avmmreaddata[1], w_hssi_common_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pld_pcs_interface = {w_hssi_common_pld_pcs_interface_avmmreaddata[7], w_hssi_common_pld_pcs_interface_avmmreaddata[6], w_hssi_common_pld_pcs_interface_avmmreaddata[5], w_hssi_common_pld_pcs_interface_avmmreaddata[4], w_hssi_common_pld_pcs_interface_avmmreaddata[3], w_hssi_common_pld_pcs_interface_avmmreaddata[2], w_hssi_common_pld_pcs_interface_avmmreaddata[1], w_hssi_common_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_rx_pcs = {w_hssi_fifo_rx_pcs_avmmreaddata[7], w_hssi_fifo_rx_pcs_avmmreaddata[6], w_hssi_fifo_rx_pcs_avmmreaddata[5], w_hssi_fifo_rx_pcs_avmmreaddata[4], w_hssi_fifo_rx_pcs_avmmreaddata[3], w_hssi_fifo_rx_pcs_avmmreaddata[2], w_hssi_fifo_rx_pcs_avmmreaddata[1], w_hssi_fifo_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_tx_pcs = {w_hssi_fifo_tx_pcs_avmmreaddata[7], w_hssi_fifo_tx_pcs_avmmreaddata[6], w_hssi_fifo_tx_pcs_avmmreaddata[5], w_hssi_fifo_tx_pcs_avmmreaddata[4], w_hssi_fifo_tx_pcs_avmmreaddata[3], w_hssi_fifo_tx_pcs_avmmreaddata[2], w_hssi_fifo_tx_pcs_avmmreaddata[1], w_hssi_fifo_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_rx_pcs = {w_hssi_gen3_rx_pcs_avmmreaddata[7], w_hssi_gen3_rx_pcs_avmmreaddata[6], w_hssi_gen3_rx_pcs_avmmreaddata[5], w_hssi_gen3_rx_pcs_avmmreaddata[4], w_hssi_gen3_rx_pcs_avmmreaddata[3], w_hssi_gen3_rx_pcs_avmmreaddata[2], w_hssi_gen3_rx_pcs_avmmreaddata[1], w_hssi_gen3_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_tx_pcs = {w_hssi_gen3_tx_pcs_avmmreaddata[7], w_hssi_gen3_tx_pcs_avmmreaddata[6], w_hssi_gen3_tx_pcs_avmmreaddata[5], w_hssi_gen3_tx_pcs_avmmreaddata[4], w_hssi_gen3_tx_pcs_avmmreaddata[3], w_hssi_gen3_tx_pcs_avmmreaddata[2], w_hssi_gen3_tx_pcs_avmmreaddata[1], w_hssi_gen3_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_rx_pcs = {w_hssi_krfec_rx_pcs_avmmreaddata[7], w_hssi_krfec_rx_pcs_avmmreaddata[6], w_hssi_krfec_rx_pcs_avmmreaddata[5], w_hssi_krfec_rx_pcs_avmmreaddata[4], w_hssi_krfec_rx_pcs_avmmreaddata[3], w_hssi_krfec_rx_pcs_avmmreaddata[2], w_hssi_krfec_rx_pcs_avmmreaddata[1], w_hssi_krfec_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_tx_pcs = {w_hssi_krfec_tx_pcs_avmmreaddata[7], w_hssi_krfec_tx_pcs_avmmreaddata[6], w_hssi_krfec_tx_pcs_avmmreaddata[5], w_hssi_krfec_tx_pcs_avmmreaddata[4], w_hssi_krfec_tx_pcs_avmmreaddata[3], w_hssi_krfec_tx_pcs_avmmreaddata[2], w_hssi_krfec_tx_pcs_avmmreaddata[1], w_hssi_krfec_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen1_2 = {w_hssi_pipe_gen1_2_avmmreaddata[7], w_hssi_pipe_gen1_2_avmmreaddata[6], w_hssi_pipe_gen1_2_avmmreaddata[5], w_hssi_pipe_gen1_2_avmmreaddata[4], w_hssi_pipe_gen1_2_avmmreaddata[3], w_hssi_pipe_gen1_2_avmmreaddata[2], w_hssi_pipe_gen1_2_avmmreaddata[1], w_hssi_pipe_gen1_2_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen3 = {w_hssi_pipe_gen3_avmmreaddata[7], w_hssi_pipe_gen3_avmmreaddata[6], w_hssi_pipe_gen3_avmmreaddata[5], w_hssi_pipe_gen3_avmmreaddata[4], w_hssi_pipe_gen3_avmmreaddata[3], w_hssi_pipe_gen3_avmmreaddata[2], w_hssi_pipe_gen3_avmmreaddata[1], w_hssi_pipe_gen3_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pcs_pma_interface = {w_hssi_rx_pcs_pma_interface_avmmreaddata[7], w_hssi_rx_pcs_pma_interface_avmmreaddata[6], w_hssi_rx_pcs_pma_interface_avmmreaddata[5], w_hssi_rx_pcs_pma_interface_avmmreaddata[4], w_hssi_rx_pcs_pma_interface_avmmreaddata[3], w_hssi_rx_pcs_pma_interface_avmmreaddata[2], w_hssi_rx_pcs_pma_interface_avmmreaddata[1], w_hssi_rx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pld_pcs_interface = {w_hssi_rx_pld_pcs_interface_avmmreaddata[7], w_hssi_rx_pld_pcs_interface_avmmreaddata[6], w_hssi_rx_pld_pcs_interface_avmmreaddata[5], w_hssi_rx_pld_pcs_interface_avmmreaddata[4], w_hssi_rx_pld_pcs_interface_avmmreaddata[3], w_hssi_rx_pld_pcs_interface_avmmreaddata[2], w_hssi_rx_pld_pcs_interface_avmmreaddata[1], w_hssi_rx_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pcs_pma_interface = {w_hssi_tx_pcs_pma_interface_avmmreaddata[7], w_hssi_tx_pcs_pma_interface_avmmreaddata[6], w_hssi_tx_pcs_pma_interface_avmmreaddata[5], w_hssi_tx_pcs_pma_interface_avmmreaddata[4], w_hssi_tx_pcs_pma_interface_avmmreaddata[3], w_hssi_tx_pcs_pma_interface_avmmreaddata[2], w_hssi_tx_pcs_pma_interface_avmmreaddata[1], w_hssi_tx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pld_pcs_interface = {w_hssi_tx_pld_pcs_interface_avmmreaddata[7], w_hssi_tx_pld_pcs_interface_avmmreaddata[6], w_hssi_tx_pld_pcs_interface_avmmreaddata[5], w_hssi_tx_pld_pcs_interface_avmmreaddata[4], w_hssi_tx_pld_pcs_interface_avmmreaddata[3], w_hssi_tx_pld_pcs_interface_avmmreaddata[2], w_hssi_tx_pld_pcs_interface_avmmreaddata[1], w_hssi_tx_pld_pcs_interface_avmmreaddata[0]};
		assign out_blockselect_hssi_10g_rx_pcs = w_hssi_10g_rx_pcs_blockselect;
		assign out_blockselect_hssi_10g_tx_pcs = w_hssi_10g_tx_pcs_blockselect;
		assign out_blockselect_hssi_8g_rx_pcs = w_hssi_8g_rx_pcs_blockselect;
		assign out_blockselect_hssi_8g_tx_pcs = w_hssi_8g_tx_pcs_blockselect;
		assign out_blockselect_hssi_common_pcs_pma_interface = w_hssi_common_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_common_pld_pcs_interface = w_hssi_common_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_fifo_rx_pcs = w_hssi_fifo_rx_pcs_blockselect;
		assign out_blockselect_hssi_fifo_tx_pcs = w_hssi_fifo_tx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_rx_pcs = w_hssi_gen3_rx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_tx_pcs = w_hssi_gen3_tx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_rx_pcs = w_hssi_krfec_rx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_tx_pcs = w_hssi_krfec_tx_pcs_blockselect;
		assign out_blockselect_hssi_pipe_gen1_2 = w_hssi_pipe_gen1_2_blockselect;
		assign out_blockselect_hssi_pipe_gen3 = w_hssi_pipe_gen3_blockselect;
		assign out_blockselect_hssi_rx_pcs_pma_interface = w_hssi_rx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_rx_pld_pcs_interface = w_hssi_rx_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_tx_pcs_pma_interface = w_hssi_tx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_tx_pld_pcs_interface = w_hssi_tx_pld_pcs_interface_blockselect;
		assign out_bond_pcs10g_out_bot = {w_hssi_10g_tx_pcs_distdwn_out_rden, w_hssi_10g_tx_pcs_distdwn_out_wren, w_hssi_10g_tx_pcs_distdwn_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs10g_out_top = {w_hssi_10g_tx_pcs_distup_out_rden, w_hssi_10g_tx_pcs_distup_out_wren, w_hssi_10g_tx_pcs_distup_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs8g_out_bot = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down, w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_down, w_hssi_8g_tx_pcs_wr_enable_out_chnl_down, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_down, w_hssi_8g_rx_pcs_wr_enable_out_chnl_down, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[0]};
		assign out_bond_pcs8g_out_top = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up, w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_up, w_hssi_8g_tx_pcs_wr_enable_out_chnl_up, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_up, w_hssi_8g_rx_pcs_wr_enable_out_chnl_up, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[0]};
		assign out_bond_pmaif_out_bot = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[0]};
		assign out_bond_pmaif_out_top = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[0]};
		assign out_hip_clk_out = {w_hssi_common_pld_pcs_interface_hip_cmn_clk[1], w_hssi_common_pld_pcs_interface_hip_cmn_clk[0], w_hssi_tx_pld_pcs_interface_hip_tx_clk};
		assign out_hip_ctrl_out = {w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[4], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[3], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[2], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[1], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[0], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[0]};
		assign out_hip_iocsr_rdy = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
		assign out_hip_iocsr_rdy_dly = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
		assign out_hip_nfrzdrv = w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
		assign out_hip_npor = w_hssi_common_pld_pcs_interface_hip_npor;
		assign out_hip_rx_data = {w_hssi_rx_pld_pcs_interface_hip_rx_data[50], w_hssi_rx_pld_pcs_interface_hip_rx_data[49], w_hssi_rx_pld_pcs_interface_hip_rx_data[48], w_hssi_rx_pld_pcs_interface_hip_rx_data[47], w_hssi_rx_pld_pcs_interface_hip_rx_data[46], w_hssi_rx_pld_pcs_interface_hip_rx_data[45], w_hssi_rx_pld_pcs_interface_hip_rx_data[44], w_hssi_rx_pld_pcs_interface_hip_rx_data[43], w_hssi_rx_pld_pcs_interface_hip_rx_data[42], w_hssi_rx_pld_pcs_interface_hip_rx_data[41], w_hssi_rx_pld_pcs_interface_hip_rx_data[40], w_hssi_rx_pld_pcs_interface_hip_rx_data[39], w_hssi_rx_pld_pcs_interface_hip_rx_data[38], w_hssi_rx_pld_pcs_interface_hip_rx_data[37], w_hssi_rx_pld_pcs_interface_hip_rx_data[36], w_hssi_rx_pld_pcs_interface_hip_rx_data[35], w_hssi_rx_pld_pcs_interface_hip_rx_data[34], w_hssi_rx_pld_pcs_interface_hip_rx_data[33], w_hssi_rx_pld_pcs_interface_hip_rx_data[32], w_hssi_rx_pld_pcs_interface_hip_rx_data[31], w_hssi_rx_pld_pcs_interface_hip_rx_data[30], w_hssi_rx_pld_pcs_interface_hip_rx_data[29], w_hssi_rx_pld_pcs_interface_hip_rx_data[28], w_hssi_rx_pld_pcs_interface_hip_rx_data[27], w_hssi_rx_pld_pcs_interface_hip_rx_data[26], w_hssi_rx_pld_pcs_interface_hip_rx_data[25], w_hssi_rx_pld_pcs_interface_hip_rx_data[24], w_hssi_rx_pld_pcs_interface_hip_rx_data[23], w_hssi_rx_pld_pcs_interface_hip_rx_data[22], w_hssi_rx_pld_pcs_interface_hip_rx_data[21], w_hssi_rx_pld_pcs_interface_hip_rx_data[20], w_hssi_rx_pld_pcs_interface_hip_rx_data[19], w_hssi_rx_pld_pcs_interface_hip_rx_data[18], w_hssi_rx_pld_pcs_interface_hip_rx_data[17], w_hssi_rx_pld_pcs_interface_hip_rx_data[16], w_hssi_rx_pld_pcs_interface_hip_rx_data[15], w_hssi_rx_pld_pcs_interface_hip_rx_data[14], w_hssi_rx_pld_pcs_interface_hip_rx_data[13], w_hssi_rx_pld_pcs_interface_hip_rx_data[12], w_hssi_rx_pld_pcs_interface_hip_rx_data[11], w_hssi_rx_pld_pcs_interface_hip_rx_data[10], w_hssi_rx_pld_pcs_interface_hip_rx_data[9], w_hssi_rx_pld_pcs_interface_hip_rx_data[8], w_hssi_rx_pld_pcs_interface_hip_rx_data[7], w_hssi_rx_pld_pcs_interface_hip_rx_data[6], w_hssi_rx_pld_pcs_interface_hip_rx_data[5], w_hssi_rx_pld_pcs_interface_hip_rx_data[4], w_hssi_rx_pld_pcs_interface_hip_rx_data[3], w_hssi_rx_pld_pcs_interface_hip_rx_data[2], w_hssi_rx_pld_pcs_interface_hip_rx_data[1], w_hssi_rx_pld_pcs_interface_hip_rx_data[0]};
		assign out_hip_usermode = w_hssi_common_pld_pcs_interface_hip_usermode;
		assign out_pld_10g_krfec_rx_blk_lock = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
		assign out_pld_10g_krfec_rx_diag_data_status = {w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1], w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[0]};
		assign out_pld_10g_krfec_rx_frame = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
		assign out_pld_10g_krfec_tx_frame = w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
		assign out_pld_10g_rx_align_val = w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
		assign out_pld_10g_rx_crc32_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
		assign out_pld_10g_rx_data_valid = w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
		assign out_pld_10g_rx_empty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
		assign out_pld_10g_rx_fifo_del = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
		assign out_pld_10g_rx_fifo_insert = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
		assign out_pld_10g_rx_fifo_num = {w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[3], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[2], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[1], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[0]};
		assign out_pld_10g_rx_frame_lock = w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
		assign out_pld_10g_rx_hi_ber = w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
		assign out_pld_10g_rx_oflw_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
		assign out_pld_10g_rx_pempty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
		assign out_pld_10g_rx_pfull = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
		assign out_pld_10g_tx_burst_en_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
		assign out_pld_10g_tx_empty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
		assign out_pld_10g_tx_fifo_num = {w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[2], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[1], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[0]};
		assign out_pld_10g_tx_full = w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
		assign out_pld_10g_tx_pempty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
		assign out_pld_10g_tx_pfull = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
		assign out_pld_10g_tx_wordslip_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
		assign out_pld_8g_a1a2_k1k2_flag = {w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[2], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[1], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[0]};
		assign out_pld_8g_empty_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
		assign out_pld_8g_empty_rx = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
		assign out_pld_8g_empty_tx = w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
		assign out_pld_8g_full_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
		assign out_pld_8g_full_rx = w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
		assign out_pld_8g_full_tx = w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
		assign out_pld_8g_rxelecidle = w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
		assign out_pld_8g_signal_detect_out = w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
		assign out_pld_8g_wa_boundary = {w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0]};
		assign out_pld_krfec_tx_alignment = w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
		assign out_pld_pcs_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
		assign out_pld_pcs_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
		assign out_pld_pma_adapt_done = w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
		assign out_pld_pma_clkdiv_rx_user = w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
		assign out_pld_pma_clkdiv_tx_user = w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
		assign out_pld_pma_clklow = w_hssi_common_pld_pcs_interface_pld_pma_clklow;
		assign out_pld_pma_fref = w_hssi_common_pld_pcs_interface_pld_pma_fref;
		assign out_pld_pma_hclk = w_hssi_common_pld_pcs_interface_pld_pma_hclk;
		assign out_pld_pma_pcie_sw_done = {w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1], w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[0]};
		assign out_pld_pma_pfdmode_lock = w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
		assign out_pld_pma_reserved_in = {w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[3], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[2], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[1], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[0]};
		assign out_pld_pma_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
		assign out_pld_pma_rx_detect_valid = w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
		assign out_pld_pma_rx_found = w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
		assign out_pld_pma_rxpll_lock = w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
		assign out_pld_pma_signal_ok = w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
		assign out_pld_pma_testbus = {w_hssi_common_pld_pcs_interface_pld_pma_testbus[7], w_hssi_common_pld_pcs_interface_pld_pma_testbus[6], w_hssi_common_pld_pcs_interface_pld_pma_testbus[5], w_hssi_common_pld_pcs_interface_pld_pma_testbus[4], w_hssi_common_pld_pcs_interface_pld_pma_testbus[3], w_hssi_common_pld_pcs_interface_pld_pma_testbus[2], w_hssi_common_pld_pcs_interface_pld_pma_testbus[1], w_hssi_common_pld_pcs_interface_pld_pma_testbus[0]};
		assign out_pld_pma_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
		assign out_pld_pmaif_mask_tx_pll = w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
		assign out_pld_reserved_out = {w_hssi_common_pld_pcs_interface_pld_reserved_out[9], w_hssi_common_pld_pcs_interface_pld_reserved_out[8], w_hssi_common_pld_pcs_interface_pld_reserved_out[7], w_hssi_common_pld_pcs_interface_pld_reserved_out[6], w_hssi_common_pld_pcs_interface_pld_reserved_out[5], w_hssi_common_pld_pcs_interface_pld_reserved_out[4], w_hssi_common_pld_pcs_interface_pld_reserved_out[3], w_hssi_common_pld_pcs_interface_pld_reserved_out[2], w_hssi_common_pld_pcs_interface_pld_reserved_out[1], w_hssi_common_pld_pcs_interface_pld_reserved_out[0]};
		assign out_pld_rx_control = {w_hssi_rx_pld_pcs_interface_pld_rx_control[19], w_hssi_rx_pld_pcs_interface_pld_rx_control[18], w_hssi_rx_pld_pcs_interface_pld_rx_control[17], w_hssi_rx_pld_pcs_interface_pld_rx_control[16], w_hssi_rx_pld_pcs_interface_pld_rx_control[15], w_hssi_rx_pld_pcs_interface_pld_rx_control[14], w_hssi_rx_pld_pcs_interface_pld_rx_control[13], w_hssi_rx_pld_pcs_interface_pld_rx_control[12], w_hssi_rx_pld_pcs_interface_pld_rx_control[11], w_hssi_rx_pld_pcs_interface_pld_rx_control[10], w_hssi_rx_pld_pcs_interface_pld_rx_control[9], w_hssi_rx_pld_pcs_interface_pld_rx_control[8], w_hssi_rx_pld_pcs_interface_pld_rx_control[7], w_hssi_rx_pld_pcs_interface_pld_rx_control[6], w_hssi_rx_pld_pcs_interface_pld_rx_control[5], w_hssi_rx_pld_pcs_interface_pld_rx_control[4], w_hssi_rx_pld_pcs_interface_pld_rx_control[3], w_hssi_rx_pld_pcs_interface_pld_rx_control[2], w_hssi_rx_pld_pcs_interface_pld_rx_control[1], w_hssi_rx_pld_pcs_interface_pld_rx_control[0]};
		assign out_pld_rx_data = {w_hssi_rx_pld_pcs_interface_pld_rx_data[127], w_hssi_rx_pld_pcs_interface_pld_rx_data[126], w_hssi_rx_pld_pcs_interface_pld_rx_data[125], w_hssi_rx_pld_pcs_interface_pld_rx_data[124], w_hssi_rx_pld_pcs_interface_pld_rx_data[123], w_hssi_rx_pld_pcs_interface_pld_rx_data[122], w_hssi_rx_pld_pcs_interface_pld_rx_data[121], w_hssi_rx_pld_pcs_interface_pld_rx_data[120], w_hssi_rx_pld_pcs_interface_pld_rx_data[119], w_hssi_rx_pld_pcs_interface_pld_rx_data[118], w_hssi_rx_pld_pcs_interface_pld_rx_data[117], w_hssi_rx_pld_pcs_interface_pld_rx_data[116], w_hssi_rx_pld_pcs_interface_pld_rx_data[115], w_hssi_rx_pld_pcs_interface_pld_rx_data[114], w_hssi_rx_pld_pcs_interface_pld_rx_data[113], w_hssi_rx_pld_pcs_interface_pld_rx_data[112], w_hssi_rx_pld_pcs_interface_pld_rx_data[111], w_hssi_rx_pld_pcs_interface_pld_rx_data[110], w_hssi_rx_pld_pcs_interface_pld_rx_data[109], w_hssi_rx_pld_pcs_interface_pld_rx_data[108], w_hssi_rx_pld_pcs_interface_pld_rx_data[107], w_hssi_rx_pld_pcs_interface_pld_rx_data[106], w_hssi_rx_pld_pcs_interface_pld_rx_data[105], w_hssi_rx_pld_pcs_interface_pld_rx_data[104], w_hssi_rx_pld_pcs_interface_pld_rx_data[103], w_hssi_rx_pld_pcs_interface_pld_rx_data[102], w_hssi_rx_pld_pcs_interface_pld_rx_data[101], w_hssi_rx_pld_pcs_interface_pld_rx_data[100], w_hssi_rx_pld_pcs_interface_pld_rx_data[99], w_hssi_rx_pld_pcs_interface_pld_rx_data[98], w_hssi_rx_pld_pcs_interface_pld_rx_data[97], w_hssi_rx_pld_pcs_interface_pld_rx_data[96], w_hssi_rx_pld_pcs_interface_pld_rx_data[95], w_hssi_rx_pld_pcs_interface_pld_rx_data[94], w_hssi_rx_pld_pcs_interface_pld_rx_data[93], w_hssi_rx_pld_pcs_interface_pld_rx_data[92], w_hssi_rx_pld_pcs_interface_pld_rx_data[91], w_hssi_rx_pld_pcs_interface_pld_rx_data[90], w_hssi_rx_pld_pcs_interface_pld_rx_data[89], w_hssi_rx_pld_pcs_interface_pld_rx_data[88], w_hssi_rx_pld_pcs_interface_pld_rx_data[87], w_hssi_rx_pld_pcs_interface_pld_rx_data[86], w_hssi_rx_pld_pcs_interface_pld_rx_data[85], w_hssi_rx_pld_pcs_interface_pld_rx_data[84], w_hssi_rx_pld_pcs_interface_pld_rx_data[83], w_hssi_rx_pld_pcs_interface_pld_rx_data[82], w_hssi_rx_pld_pcs_interface_pld_rx_data[81], w_hssi_rx_pld_pcs_interface_pld_rx_data[80], w_hssi_rx_pld_pcs_interface_pld_rx_data[79], w_hssi_rx_pld_pcs_interface_pld_rx_data[78], w_hssi_rx_pld_pcs_interface_pld_rx_data[77], w_hssi_rx_pld_pcs_interface_pld_rx_data[76], w_hssi_rx_pld_pcs_interface_pld_rx_data[75], w_hssi_rx_pld_pcs_interface_pld_rx_data[74], w_hssi_rx_pld_pcs_interface_pld_rx_data[73], w_hssi_rx_pld_pcs_interface_pld_rx_data[72], w_hssi_rx_pld_pcs_interface_pld_rx_data[71], w_hssi_rx_pld_pcs_interface_pld_rx_data[70], w_hssi_rx_pld_pcs_interface_pld_rx_data[69], w_hssi_rx_pld_pcs_interface_pld_rx_data[68], w_hssi_rx_pld_pcs_interface_pld_rx_data[67], w_hssi_rx_pld_pcs_interface_pld_rx_data[66], w_hssi_rx_pld_pcs_interface_pld_rx_data[65], w_hssi_rx_pld_pcs_interface_pld_rx_data[64], w_hssi_rx_pld_pcs_interface_pld_rx_data[63], w_hssi_rx_pld_pcs_interface_pld_rx_data[62], w_hssi_rx_pld_pcs_interface_pld_rx_data[61], w_hssi_rx_pld_pcs_interface_pld_rx_data[60], w_hssi_rx_pld_pcs_interface_pld_rx_data[59], w_hssi_rx_pld_pcs_interface_pld_rx_data[58], w_hssi_rx_pld_pcs_interface_pld_rx_data[57], w_hssi_rx_pld_pcs_interface_pld_rx_data[56], w_hssi_rx_pld_pcs_interface_pld_rx_data[55], w_hssi_rx_pld_pcs_interface_pld_rx_data[54], w_hssi_rx_pld_pcs_interface_pld_rx_data[53], w_hssi_rx_pld_pcs_interface_pld_rx_data[52], w_hssi_rx_pld_pcs_interface_pld_rx_data[51], w_hssi_rx_pld_pcs_interface_pld_rx_data[50], w_hssi_rx_pld_pcs_interface_pld_rx_data[49], w_hssi_rx_pld_pcs_interface_pld_rx_data[48], w_hssi_rx_pld_pcs_interface_pld_rx_data[47], w_hssi_rx_pld_pcs_interface_pld_rx_data[46], w_hssi_rx_pld_pcs_interface_pld_rx_data[45], w_hssi_rx_pld_pcs_interface_pld_rx_data[44], w_hssi_rx_pld_pcs_interface_pld_rx_data[43], w_hssi_rx_pld_pcs_interface_pld_rx_data[42], w_hssi_rx_pld_pcs_interface_pld_rx_data[41], w_hssi_rx_pld_pcs_interface_pld_rx_data[40], w_hssi_rx_pld_pcs_interface_pld_rx_data[39], w_hssi_rx_pld_pcs_interface_pld_rx_data[38], w_hssi_rx_pld_pcs_interface_pld_rx_data[37], w_hssi_rx_pld_pcs_interface_pld_rx_data[36], w_hssi_rx_pld_pcs_interface_pld_rx_data[35], w_hssi_rx_pld_pcs_interface_pld_rx_data[34], w_hssi_rx_pld_pcs_interface_pld_rx_data[33], w_hssi_rx_pld_pcs_interface_pld_rx_data[32], w_hssi_rx_pld_pcs_interface_pld_rx_data[31], w_hssi_rx_pld_pcs_interface_pld_rx_data[30], w_hssi_rx_pld_pcs_interface_pld_rx_data[29], w_hssi_rx_pld_pcs_interface_pld_rx_data[28], w_hssi_rx_pld_pcs_interface_pld_rx_data[27], w_hssi_rx_pld_pcs_interface_pld_rx_data[26], w_hssi_rx_pld_pcs_interface_pld_rx_data[25], w_hssi_rx_pld_pcs_interface_pld_rx_data[24], w_hssi_rx_pld_pcs_interface_pld_rx_data[23], w_hssi_rx_pld_pcs_interface_pld_rx_data[22], w_hssi_rx_pld_pcs_interface_pld_rx_data[21], w_hssi_rx_pld_pcs_interface_pld_rx_data[20], w_hssi_rx_pld_pcs_interface_pld_rx_data[19], w_hssi_rx_pld_pcs_interface_pld_rx_data[18], w_hssi_rx_pld_pcs_interface_pld_rx_data[17], w_hssi_rx_pld_pcs_interface_pld_rx_data[16], w_hssi_rx_pld_pcs_interface_pld_rx_data[15], w_hssi_rx_pld_pcs_interface_pld_rx_data[14], w_hssi_rx_pld_pcs_interface_pld_rx_data[13], w_hssi_rx_pld_pcs_interface_pld_rx_data[12], w_hssi_rx_pld_pcs_interface_pld_rx_data[11], w_hssi_rx_pld_pcs_interface_pld_rx_data[10], w_hssi_rx_pld_pcs_interface_pld_rx_data[9], w_hssi_rx_pld_pcs_interface_pld_rx_data[8], w_hssi_rx_pld_pcs_interface_pld_rx_data[7], w_hssi_rx_pld_pcs_interface_pld_rx_data[6], w_hssi_rx_pld_pcs_interface_pld_rx_data[5], w_hssi_rx_pld_pcs_interface_pld_rx_data[4], w_hssi_rx_pld_pcs_interface_pld_rx_data[3], w_hssi_rx_pld_pcs_interface_pld_rx_data[2], w_hssi_rx_pld_pcs_interface_pld_rx_data[1], w_hssi_rx_pld_pcs_interface_pld_rx_data[0]};
		assign out_pld_rx_prbs_done = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
		assign out_pld_rx_prbs_err = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
		assign out_pld_test_data = {w_hssi_common_pld_pcs_interface_pld_test_data[19], w_hssi_common_pld_pcs_interface_pld_test_data[18], w_hssi_common_pld_pcs_interface_pld_test_data[17], w_hssi_common_pld_pcs_interface_pld_test_data[16], w_hssi_common_pld_pcs_interface_pld_test_data[15], w_hssi_common_pld_pcs_interface_pld_test_data[14], w_hssi_common_pld_pcs_interface_pld_test_data[13], w_hssi_common_pld_pcs_interface_pld_test_data[12], w_hssi_common_pld_pcs_interface_pld_test_data[11], w_hssi_common_pld_pcs_interface_pld_test_data[10], w_hssi_common_pld_pcs_interface_pld_test_data[9], w_hssi_common_pld_pcs_interface_pld_test_data[8], w_hssi_common_pld_pcs_interface_pld_test_data[7], w_hssi_common_pld_pcs_interface_pld_test_data[6], w_hssi_common_pld_pcs_interface_pld_test_data[5], w_hssi_common_pld_pcs_interface_pld_test_data[4], w_hssi_common_pld_pcs_interface_pld_test_data[3], w_hssi_common_pld_pcs_interface_pld_test_data[2], w_hssi_common_pld_pcs_interface_pld_test_data[1], w_hssi_common_pld_pcs_interface_pld_test_data[0]};
		assign out_pld_uhsif_lock = w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
		assign out_pld_uhsif_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
		assign out_pma_adapt_start = w_hssi_common_pcs_pma_interface_pma_adapt_start;
		assign out_pma_atpg_los_en_n = w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
		assign out_pma_csr_test_dis = w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
		assign out_pma_current_coeff = {w_hssi_common_pcs_pma_interface_pma_current_coeff[17], w_hssi_common_pcs_pma_interface_pma_current_coeff[16], w_hssi_common_pcs_pma_interface_pma_current_coeff[15], w_hssi_common_pcs_pma_interface_pma_current_coeff[14], w_hssi_common_pcs_pma_interface_pma_current_coeff[13], w_hssi_common_pcs_pma_interface_pma_current_coeff[12], w_hssi_common_pcs_pma_interface_pma_current_coeff[11], w_hssi_common_pcs_pma_interface_pma_current_coeff[10], w_hssi_common_pcs_pma_interface_pma_current_coeff[9], w_hssi_common_pcs_pma_interface_pma_current_coeff[8], w_hssi_common_pcs_pma_interface_pma_current_coeff[7], w_hssi_common_pcs_pma_interface_pma_current_coeff[6], w_hssi_common_pcs_pma_interface_pma_current_coeff[5], w_hssi_common_pcs_pma_interface_pma_current_coeff[4], w_hssi_common_pcs_pma_interface_pma_current_coeff[3], w_hssi_common_pcs_pma_interface_pma_current_coeff[2], w_hssi_common_pcs_pma_interface_pma_current_coeff[1], w_hssi_common_pcs_pma_interface_pma_current_coeff[0]};
		assign out_pma_current_rxpreset = {w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[1], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[0]};
		assign out_pma_early_eios = w_hssi_common_pcs_pma_interface_pma_early_eios;
		assign out_pma_eye_monitor = {w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0]};
		assign out_pma_interface_select = {w_hssi_common_pcs_pma_interface_pma_interface_select[1], w_hssi_common_pcs_pma_interface_pma_interface_select[0]};
		assign out_pma_ltd_b = w_hssi_common_pcs_pma_interface_pma_ltd_b;
		assign out_pma_ltr = w_hssi_common_pcs_pma_interface_pma_ltr;
		assign out_pma_nfrzdrv = w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
		assign out_pma_nrpi_freeze = w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
		assign out_pma_pcie_switch = {w_hssi_common_pcs_pma_interface_pma_pcie_switch[1], w_hssi_common_pcs_pma_interface_pma_pcie_switch[0]};
		assign out_pma_ppm_lock = w_hssi_common_pcs_pma_interface_pma_ppm_lock;
		assign out_pma_reserved_out = {w_hssi_common_pcs_pma_interface_pma_reserved_out[4], w_hssi_common_pcs_pma_interface_pma_reserved_out[3], w_hssi_common_pcs_pma_interface_pma_reserved_out[2], w_hssi_common_pcs_pma_interface_pma_reserved_out[1], w_hssi_common_pcs_pma_interface_pma_reserved_out[0]};
		assign out_pma_rs_lpbk_b = w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
		assign out_pma_rx_clkslip = w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
		assign out_pma_rx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
		assign out_pma_rxpma_rstb = w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
		assign out_pma_scan_mode_n = w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
		assign out_pma_scan_shift_n = w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
		assign out_pma_tx_bitslip = w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
		assign out_pma_tx_bonding_rstb = w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
		assign out_pma_tx_elec_idle = w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
		assign out_pma_tx_pma_data = {w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0]};
		assign out_pma_tx_qpi_pulldn = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
		assign out_pma_tx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
		assign out_pma_tx_txdetectrx = w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
		assign out_pma_txpma_rstb = w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	endgenerate
endmodule
module twentynm_pcs_rev_20nm5es
	#(
	//PARAM_LIST_START
		parameter xcvr_native_mode = "mode_duplex",  // mode_duplex, mode_rx_only, mode_tx_only
		
		// parameters for twentynm_hssi_10g_rx_pcs
		parameter hssi_10g_rx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_align_del = "align_del_en", // align_del_dis|align_del_en
		parameter hssi_10g_rx_pcs_ber_bit_err_total_cnt = "bit_err_total_cnt_10g", // bit_err_total_cnt_10g
		parameter hssi_10g_rx_pcs_ber_clken = "ber_clk_dis", // ber_clk_dis|ber_clk_en
		parameter hssi_10g_rx_pcs_ber_xus_timer_window = 21'b100110001001010,
		parameter hssi_10g_rx_pcs_bitslip_mode = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_rx_pcs_blksync_bitslip_type = "bitslip_comb", // bitslip_comb|bitslip_reg
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_cnt = 3'b1,
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_type = "bitslip_match", // bitslip_match|bitslip_cnt
		parameter hssi_10g_rx_pcs_blksync_bypass = "blksync_bypass_dis", // blksync_bypass_dis|blksync_bypass_en
		parameter hssi_10g_rx_pcs_blksync_clken = "blksync_clk_dis", // blksync_clk_dis|blksync_clk_en
		parameter hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt = "enum_invalid_sh_cnt_10g", // enum_invalid_sh_cnt_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock = "knum_sh_cnt_postlock_10g", // knum_sh_cnt_postlock_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock = "knum_sh_cnt_prelock_10g", // knum_sh_cnt_prelock_10g
		parameter hssi_10g_rx_pcs_blksync_pipeln = "blksync_pipeln_dis", // blksync_pipeln_dis|blksync_pipeln_en
		parameter hssi_10g_rx_pcs_clr_errblk_cnt_en = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_control_del = "control_del_all", // control_del_all|control_del_none
		parameter hssi_10g_rx_pcs_crcchk_bypass = "crcchk_bypass_dis", // crcchk_bypass_dis|crcchk_bypass_en
		parameter hssi_10g_rx_pcs_crcchk_clken = "crcchk_clk_dis", // crcchk_clk_dis|crcchk_clk_en
		parameter hssi_10g_rx_pcs_crcchk_inv = "crcchk_inv_dis", // crcchk_inv_dis|crcchk_inv_en
		parameter hssi_10g_rx_pcs_crcchk_pipeln = "crcchk_pipeln_dis", // crcchk_pipeln_dis|crcchk_pipeln_en
		parameter hssi_10g_rx_pcs_crcflag_pipeln = "crcflag_pipeln_dis", // crcflag_pipeln_dis|crcflag_pipeln_en
		parameter hssi_10g_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_rx_pcs_dec64b66b_clken = "dec64b66b_clk_dis", // dec64b66b_clk_dis|dec64b66b_clk_en
		parameter hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass = "dec_64b66b_rxsm_bypass_dis", // dec_64b66b_rxsm_bypass_dis|dec_64b66b_rxsm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_bypass = "descrm_bypass_en", // descrm_bypass_dis|descrm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_clken = "descrm_clk_dis", // descrm_clk_dis|descrm_clk_en
		parameter hssi_10g_rx_pcs_descrm_mode = "async", // async|sync
		parameter hssi_10g_rx_pcs_descrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_dft_clk_out_sel = "rx_master_clk", // rx_master_clk|rx_gbexp_clk|rx_blksync_clk|rx_descrm_clk|rx_frmsync_clk|rx_64b66bdec_clk|rx_ber_clk|rx_rand_clk|rx_crcchk_clk|rx_wrfifo_clk|rx_rdfifo_clk|rx_fec_clk
		parameter hssi_10g_rx_pcs_dis_signal_ok = "dis_signal_ok_dis", // dis_signal_ok_dis|dis_signal_ok_en
		parameter hssi_10g_rx_pcs_dispchk_bypass = "dispchk_bypass_dis", // dispchk_bypass_dis|dispchk_bypass_en
		parameter hssi_10g_rx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_rx_pcs_fast_path = "fast_path_dis", // fast_path_dis|fast_path_en
		parameter hssi_10g_rx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_rx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_rx_pcs_fifo_double_read = "fifo_double_read_dis", // fifo_double_read_dis|fifo_double_read_en
		parameter hssi_10g_rx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_rx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_rx_pcs_force_align = "force_align_dis", // force_align_dis|force_align_en
		parameter hssi_10g_rx_pcs_frmsync_bypass = "frmsync_bypass_dis", // frmsync_bypass_dis|frmsync_bypass_en
		parameter hssi_10g_rx_pcs_frmsync_clken = "frmsync_clk_dis", // frmsync_clk_dis|frmsync_clk_en
		parameter hssi_10g_rx_pcs_frmsync_enum_scrm = "enum_scrm_default", // enum_scrm_default
		parameter hssi_10g_rx_pcs_frmsync_enum_sync = "enum_sync_default", // enum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_flag_type = "all_framing_words", // all_framing_words|location_only
		parameter hssi_10g_rx_pcs_frmsync_knum_sync = "knum_sync_default", // knum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_mfrm_length = 16'b100000000000,
		parameter hssi_10g_rx_pcs_frmsync_pipeln = "frmsync_pipeln_dis", // frmsync_pipeln_dis|frmsync_pipeln_en
		parameter hssi_10g_rx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_rx_pcs_gb_rx_idwidth = "width_32", // width_40|width_32|width_64
		parameter hssi_10g_rx_pcs_gb_rx_odwidth = "width_66", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_rx_pcs_gbexp_clken = "gbexp_clk_dis", // gbexp_clk_dis|gbexp_clk_en
		parameter hssi_10g_rx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_10g_rx_pcs_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_rx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_rx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_rx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_rx_pcs_pld_if_type = "fifo", // fifo|reg
		parameter hssi_10g_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_rx_pcs_rand_clken = "rand_clk_dis", // rand_clk_dis|rand_clk_en
		parameter hssi_10g_rx_pcs_rd_clk_sel = "rd_rx_pma_clk", // rd_rx_pld_clk|rd_rx_pma_clk|rd_refclk_dig
		parameter hssi_10g_rx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_rx_pcs_rx_fifo_write_ctrl = "blklock_stops", // blklock_stops|blklock_ignore
		parameter hssi_10g_rx_pcs_rx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_rx_pcs_rx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_rx_pcs_rx_signal_ok_sel = "synchronized_ver", // synchronized_ver|nonsync_ver
		parameter hssi_10g_rx_pcs_rx_sm_bypass = "rx_sm_bypass_dis", // rx_sm_bypass_dis|rx_sm_bypass_en
		parameter hssi_10g_rx_pcs_rx_sm_hiber = "rx_sm_hiber_en", // rx_sm_hiber_en|rx_sm_hiber_dis
		parameter hssi_10g_rx_pcs_rx_sm_pipeln = "rx_sm_pipeln_dis", // rx_sm_pipeln_dis|rx_sm_pipeln_en
		parameter hssi_10g_rx_pcs_rx_testbus_sel = "crc32_chk_testbus1", // crc32_chk_testbus1|crc32_chk_testbus2|frame_sync_testbus1|frame_sync_testbus2|dec64b66b_testbus|rxsm_testbus|ber_testbus|blksync_testbus1|blksync_testbus2|gearbox_exp_testbus|random_ver_testbus|descramble_testbus|blank_testbus|rx_fifo_testbus1|rx_fifo_testbus2
		parameter hssi_10g_rx_pcs_rx_true_b2b = "b2b", // single|b2b
		parameter hssi_10g_rx_pcs_rxfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_rx_pcs_rxfifo_full = "full_default", // full_default
		parameter hssi_10g_rx_pcs_rxfifo_mode = "phase_comp", // register_mode|clk_comp_10g|generic_interlaken|generic_basic|phase_comp|phase_comp_dv
		parameter hssi_10g_rx_pcs_rxfifo_pempty = 5'b10,
		parameter hssi_10g_rx_pcs_rxfifo_pfull = 5'b10111,
		parameter hssi_10g_rx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_rx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_rx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_10g_tx_pcs
		parameter hssi_10g_tx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_bitslip_en = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_10g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_10g_tx_pcs_comp_cnt = 8'b0,
		parameter hssi_10g_tx_pcs_compin_sel = "compin_master", // compin_master|compin_slave_top|compin_slave_bot|compin_default
		parameter hssi_10g_tx_pcs_crcgen_bypass = "crcgen_bypass_dis", // crcgen_bypass_dis|crcgen_bypass_en
		parameter hssi_10g_tx_pcs_crcgen_clken = "crcgen_clk_dis", // crcgen_clk_dis|crcgen_clk_en
		parameter hssi_10g_tx_pcs_crcgen_err = "crcgen_err_dis", // crcgen_err_dis|crcgen_err_en
		parameter hssi_10g_tx_pcs_crcgen_inv = "crcgen_inv_dis", // crcgen_inv_dis|crcgen_inv_en
		parameter hssi_10g_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_tx_pcs_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_10g_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_tx_pcs_dft_clk_out_sel = "tx_master_clk", // tx_master_clk|tx_rdfifo_clk|tx_frmgen_clk|tx_crcgen_clk|tx_64b66benc_txsm_clk|tx_scrm_clk|tx_dispgen_clk|tx_gbred_clk|tx_wrfifo_clk|tx_fec_clk
		parameter hssi_10g_tx_pcs_dispgen_bypass = "dispgen_bypass_dis", // dispgen_bypass_dis|dispgen_bypass_en
		parameter hssi_10g_tx_pcs_dispgen_clken = "dispgen_clk_dis", // dispgen_clk_dis|dispgen_clk_en
		parameter hssi_10g_tx_pcs_dispgen_err = "dispgen_err_dis", // dispgen_err_dis|dispgen_err_en
		parameter hssi_10g_tx_pcs_dispgen_pipeln = "dispgen_pipeln_dis", // dispgen_pipeln_dis|dispgen_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_bypass_pipeln = "distdwn_bypass_pipeln_dis", // distdwn_bypass_pipeln_dis|distdwn_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_master = "distdwn_master_en", // distdwn_master_en|distdwn_master_dis
		parameter hssi_10g_tx_pcs_distup_bypass_pipeln = "distup_bypass_pipeln_dis", // distup_bypass_pipeln_dis|distup_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distup_master = "distup_master_en", // distup_master_en|distup_master_dis
		parameter hssi_10g_tx_pcs_dv_bond = "dv_bond_dis", // dv_bond_en|dv_bond_dis
		parameter hssi_10g_tx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_tx_pcs_enc64b66b_txsm_clken = "enc64b66b_txsm_clk_dis", // enc64b66b_txsm_clk_dis|enc64b66b_txsm_clk_en
		parameter hssi_10g_tx_pcs_enc_64b66b_txsm_bypass = "enc_64b66b_txsm_bypass_dis", // enc_64b66b_txsm_bypass_dis|enc_64b66b_txsm_bypass_en
		parameter hssi_10g_tx_pcs_fastpath = "fastpath_dis", // fastpath_dis|fastpath_en
		parameter hssi_10g_tx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_tx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_tx_pcs_fifo_double_write = "fifo_double_write_dis", // fifo_double_write_dis|fifo_double_write_en
		parameter hssi_10g_tx_pcs_fifo_reg_fast = "fifo_reg_fast_dis", // fifo_reg_fast_dis|fifo_reg_fast_en
		parameter hssi_10g_tx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_tx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_tx_pcs_frmgen_burst = "frmgen_burst_dis", // frmgen_burst_dis|frmgen_burst_en
		parameter hssi_10g_tx_pcs_frmgen_bypass = "frmgen_bypass_dis", // frmgen_bypass_dis|frmgen_bypass_en
		parameter hssi_10g_tx_pcs_frmgen_clken = "frmgen_clk_dis", // frmgen_clk_dis|frmgen_clk_en
		parameter hssi_10g_tx_pcs_frmgen_mfrm_length = 16'b100000000000,
		parameter hssi_10g_tx_pcs_frmgen_pipeln = "frmgen_pipeln_dis", // frmgen_pipeln_dis|frmgen_pipeln_en
		parameter hssi_10g_tx_pcs_frmgen_pyld_ins = "frmgen_pyld_ins_dis", // frmgen_pyld_ins_dis|frmgen_pyld_ins_en
		parameter hssi_10g_tx_pcs_frmgen_wordslip = "frmgen_wordslip_dis", // frmgen_wordslip_dis|frmgen_wordslip_en
		parameter hssi_10g_tx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_tx_pcs_gb_pipeln_bypass = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_gb_tx_idwidth = "width_50", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_tx_pcs_gb_tx_odwidth = "width_32", // width_32|width_40|width_64
		parameter hssi_10g_tx_pcs_gbred_clken = "gbred_clk_dis", // gbred_clk_dis|gbred_clk_en
		parameter hssi_10g_tx_pcs_indv = "indv_en", // indv_en|indv_dis
		parameter hssi_10g_tx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_tx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_tx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_tx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del6|phcomp_rd_del5|phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_tx_pcs_pld_if_type = "fifo", // fifo|reg|fastreg
		parameter hssi_10g_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_tx_pcs_pseudo_random = "all_0", // two_lf|all_0
		parameter hssi_10g_tx_pcs_pseudo_seed_a = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_pseudo_seed_b = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_random_disp = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_tx_pcs_scrm_bypass = "scrm_bypass_dis", // scrm_bypass_dis|scrm_bypass_en
		parameter hssi_10g_tx_pcs_scrm_clken = "scrm_clk_dis", // scrm_clk_dis|scrm_clk_en
		parameter hssi_10g_tx_pcs_scrm_mode = "async", // async|sync
		parameter hssi_10g_tx_pcs_scrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_sh_err = "sh_err_dis", // sh_err_dis|sh_err_en
		parameter hssi_10g_tx_pcs_sop_mark = "sop_mark_dis", // sop_mark_en|sop_mark_dis
		parameter hssi_10g_tx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_tx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_tx_pcs_tx_scrm_err = "scrm_err_dis", // scrm_err_dis|scrm_err_en
		parameter hssi_10g_tx_pcs_tx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_tx_pcs_tx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_tx_pcs_tx_sm_bypass = "tx_sm_bypass_dis", // tx_sm_bypass_dis|tx_sm_bypass_en
		parameter hssi_10g_tx_pcs_tx_sm_pipeln = "tx_sm_pipeln_dis", // tx_sm_pipeln_dis|tx_sm_pipeln_en
		parameter hssi_10g_tx_pcs_tx_testbus_sel = "crc32_gen_testbus1", // crc32_gen_testbus1|crc32_gen_testbus2|disp_gen_testbus1|disp_gen_testbus2|frame_gen_testbus1|frame_gen_testbus2|enc64b66b_testbus|txsm_testbus|tx_cp_bond_testbus|gearbox_red_testbus|scramble_testbus|blank_testbus|tx_fifo_testbus1|tx_fifo_testbus2
		parameter hssi_10g_tx_pcs_txfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_tx_pcs_txfifo_full = "full_default", // full_default
		parameter hssi_10g_tx_pcs_txfifo_mode = "phase_comp", // register_mode|interlaken_generic|basic_generic|phase_comp
		parameter hssi_10g_tx_pcs_txfifo_pempty = 4'b10,
		parameter hssi_10g_tx_pcs_txfifo_pfull = 4'b1011,
		parameter hssi_10g_tx_pcs_wr_clk_sel = "wr_tx_pma_clk", // wr_tx_pld_clk|wr_tx_pma_clk|wr_refclk_dig
		parameter hssi_10g_tx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_8g_rx_pcs
		parameter hssi_8g_rx_pcs_auto_error_replacement = "dis_err_replace", // dis_err_replace|en_err_replace
		parameter hssi_8g_rx_pcs_auto_speed_nego = "dis_asn", // dis_asn|en_asn_g2_freq_scal
		parameter hssi_8g_rx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_rx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_rx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_rx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_rx_pcs_byte_deserializer = "dis_bds", // dis_bds|en_bds_by_2|en_bds_by_4|en_bds_by_2_det
		parameter hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask = "dis_rxvalid_mask", // dis_rxvalid_mask|en_rxvalid_mask
		parameter hssi_8g_rx_pcs_clkcmp_pattern_n = 20'b0,
		parameter hssi_8g_rx_pcs_clkcmp_pattern_p = 20'b0,
		parameter hssi_8g_rx_pcs_clock_gate_bds_dec_asn = "dis_bds_dec_asn_clk_gating", // dis_bds_dec_asn_clk_gating|en_bds_dec_asn_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_cdr_eidle = "dis_cdr_eidle_clk_gating", // dis_cdr_eidle_clk_gating|en_cdr_eidle_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk = "dis_dw_pc_wrclk_gating", // dis_dw_pc_wrclk_gating|en_dw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_rd = "dis_dw_rm_rdclk_gating", // dis_dw_rm_rdclk_gating|en_dw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_wr = "dis_dw_rm_wrclk_gating", // dis_dw_rm_wrclk_gating|en_dw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_wa = "dis_dw_wa_clk_gating", // dis_dw_wa_clk_gating|en_dw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_pc_rdclk = "dis_pc_rdclk_gating", // dis_pc_rdclk_gating|en_pc_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk = "dis_sw_pc_wrclk_gating", // dis_sw_pc_wrclk_gating|en_sw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_rd = "dis_sw_rm_rdclk_gating", // dis_sw_rm_rdclk_gating|en_sw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_wr = "dis_sw_rm_wrclk_gating", // dis_sw_rm_wrclk_gating|en_sw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_wa = "dis_sw_wa_clk_gating", // dis_sw_wa_clk_gating|en_sw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_observation_in_pld_core = "internal_sw_wa_clk", // internal_sw_wa_clk|internal_dw_wa_clk|internal_cdr_eidle_clk|internal_sm_rm_wr_clk|internal_dw_rm_wr_clk|internal_clk_2_b|internal_sw_rm_rd_clk|internal_dw_rm_rd_clk|internal_sw_rx_wr_clk|internal_dw_rx_wr_clk|internal_rx_rd_clk|internal_rx_pma_clk_gen3|internal_rx_rcvd_clk_gen3
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_rx_pcs_eidle_entry_eios = "dis_eidle_eios", // dis_eidle_eios|en_eidle_eios
		parameter hssi_8g_rx_pcs_eidle_entry_iei = "dis_eidle_iei", // dis_eidle_iei|en_eidle_iei
		parameter hssi_8g_rx_pcs_eidle_entry_sd = "dis_eidle_sd", // dis_eidle_sd|en_eidle_sd
		parameter hssi_8g_rx_pcs_eightb_tenb_decoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_rx_pcs_err_flags_sel = "err_flags_wa", // err_flags_wa|err_flags_8b10b
		parameter hssi_8g_rx_pcs_fixed_pat_det = "dis_fixed_patdet", // dis_fixed_patdet|en_fixed_patdet
		parameter hssi_8g_rx_pcs_fixed_pat_num = 4'b1111,
		parameter hssi_8g_rx_pcs_force_signal_detect = "en_force_signal_detect", // en_force_signal_detect|dis_force_signal_detect
		parameter hssi_8g_rx_pcs_gen3_clk_en = "disable_clk", // disable_clk|enable_clk
		parameter hssi_8g_rx_pcs_gen3_rx_clk_sel = "rcvd_clk", // en_dig_clk1_8g|rcvd_clk
		parameter hssi_8g_rx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // en_dig_clk2_8g|tx_pma_clk
		parameter hssi_8g_rx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_rx_pcs_ibm_invalid_code = "dis_ibm_invalid_code", // dis_ibm_invalid_code|en_ibm_invalid_code
		parameter hssi_8g_rx_pcs_invalid_code_flag_only = "dis_invalid_code_only", // dis_invalid_code_only|en_invalid_code_only
		parameter hssi_8g_rx_pcs_pad_or_edb_error_replace = "replace_edb", // replace_edb|replace_edb_dynamic|replace_pad
		parameter hssi_8g_rx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_rx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_rx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_rx_pcs_pipe_if_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_8g_rx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_rx_pcs_polinv_8b10b_dec = "dis_polinv_8b10b_dec", // dis_polinv_8b10b_dec|en_polinv_8b10b_dec
		parameter hssi_8g_rx_pcs_prot_mode = "gige", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic_rm_enable|basic_rm_disable|disabled_prot_mode
		parameter hssi_8g_rx_pcs_rate_match = "dis_rm", // dis_rm|gige_rm|pipe_rm|pipe_rm_0ppm|sw_basic_rm|dw_basic_rm
		parameter hssi_8g_rx_pcs_rate_match_del_thres = "dis_rm_del_thres", // dis_rm_del_thres|gige_rm_del_thres|pipe_rm_del_thres|pipe_rm_0ppm_del_thres|sw_basic_rm_del_thres|dw_basic_rm_del_thres
		parameter hssi_8g_rx_pcs_rate_match_empty_thres = "dis_rm_empty_thres", // dis_rm_empty_thres|gige_rm_empty_thres|pipe_rm_empty_thres|pipe_rm_0ppm_empty_thres|sw_basic_rm_empty_thres|dw_basic_rm_empty_thres
		parameter hssi_8g_rx_pcs_rate_match_full_thres = "dis_rm_full_thres", // dis_rm_full_thres|gige_rm_full_thres|pipe_rm_full_thres|pipe_rm_0ppm_full_thres|sw_basic_rm_full_thres|dw_basic_rm_full_thres
		parameter hssi_8g_rx_pcs_rate_match_ins_thres = "dis_rm_ins_thres", // dis_rm_ins_thres|gige_rm_ins_thres|pipe_rm_ins_thres|pipe_rm_0ppm_ins_thres|sw_basic_rm_ins_thres|dw_basic_rm_ins_thres
		parameter hssi_8g_rx_pcs_rate_match_start_thres = "dis_rm_start_thres", // dis_rm_start_thres|gige_rm_start_thres|pipe_rm_start_thres|pipe_rm_0ppm_start_thres|sw_basic_rm_start_thres|dw_basic_rm_start_thres
		parameter hssi_8g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_rx_pcs_rx_clk2 = "rcvd_clk_clk2", // rcvd_clk_clk2|tx_pma_clock_clk2|refclk_dig2_clk2
		parameter hssi_8g_rx_pcs_rx_clk_free_running = "en_rx_clk_free_run", // dis_rx_clk_free_run|en_rx_clk_free_run
		parameter hssi_8g_rx_pcs_rx_pcs_urst = "en_rx_pcs_urst", // dis_rx_pcs_urst|en_rx_pcs_urst
		parameter hssi_8g_rx_pcs_rx_rcvd_clk = "rcvd_clk_rcvd_clk", // rcvd_clk_rcvd_clk|tx_pma_clock_rcvd_clk
		parameter hssi_8g_rx_pcs_rx_rd_clk = "pld_rx_clk", // pld_rx_clk|rx_clk
		parameter hssi_8g_rx_pcs_rx_refclk = "dis_refclk_sel", // dis_refclk_sel|en_refclk_sel
		parameter hssi_8g_rx_pcs_rx_wr_clk = "rx_clk2_div_1_2_4", // rx_clk2_div_1_2_4|txfifo_rd_clk
		parameter hssi_8g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_rx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_rx_pcs_sync_sm_idle_eios = "dis_syncsm_idle", // dis_syncsm_idle|en_syncsm_idle
		parameter hssi_8g_rx_pcs_test_bus_sel = "tx_testbus", // tx_testbus|tx_ctrl_plane_testbus|wa_testbus|rm_testbus|rx_ctrl_testbus|pcie_ctrl_testbus|rx_ctrl_plane_testbus
		parameter hssi_8g_rx_pcs_tx_rx_parallel_loopback = "dis_plpbk", // dis_plpbk|en_plpbk
		parameter hssi_8g_rx_pcs_wa_boundary_lock_ctrl = "bit_slip", // bit_slip|sync_sm|deterministic_latency|auto_align_pld_ctrl
		parameter hssi_8g_rx_pcs_wa_clk_slip_spacing = 10'b10000,
		parameter hssi_8g_rx_pcs_wa_det_latency_sync_status_beh = "assert_sync_status_non_imm", // assert_sync_status_imm|assert_sync_status_non_imm|dont_care_assert_sync
		parameter hssi_8g_rx_pcs_wa_disp_err_flag = "dis_disp_err_flag", // dis_disp_err_flag|en_disp_err_flag
		parameter hssi_8g_rx_pcs_wa_kchar = "dis_kchar", // dis_kchar|en_kchar
		parameter hssi_8g_rx_pcs_wa_pd = "wa_pd_10", // wa_pd_7|wa_pd_10|wa_pd_20|wa_pd_40|wa_pd_8_sw|wa_pd_8_dw|wa_pd_16_sw|wa_pd_16_dw|wa_pd_32
		parameter hssi_8g_rx_pcs_wa_pd_data = 40'b0,
		parameter hssi_8g_rx_pcs_wa_pd_polarity = "dis_pd_both_pol", // dis_pd_both_pol|en_pd_both_pol|dont_care_both_pol
		parameter hssi_8g_rx_pcs_wa_pld_controlled = "dis_pld_ctrl", // dis_pld_ctrl|pld_ctrl_sw|rising_edge_sensitive_dw|level_sensitive_dw
		parameter hssi_8g_rx_pcs_wa_renumber_data = 6'b0,
		parameter hssi_8g_rx_pcs_wa_rgnumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rknumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rosnumber_data = 2'b0,
		parameter hssi_8g_rx_pcs_wa_rvnumber_data = 13'b0,
		parameter hssi_8g_rx_pcs_wa_sync_sm_ctrl = "gige_sync_sm", // gige_sync_sm|pipe_sync_sm|sw_basic_sync_sm|dw_basic_sync_sm|fibre_channel_sync_sm
		parameter hssi_8g_rx_pcs_wait_cnt = 12'b0,
		
		// parameters for twentynm_hssi_8g_tx_pcs
		parameter hssi_8g_tx_pcs_auto_speed_nego_gen2 = "dis_asn_g2", // dis_asn_g2|en_asn_g2_freq_scal
		parameter hssi_8g_tx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_tx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_tx_pcs_byte_serializer = "dis_bs", // dis_bs|en_bs_by_2|en_bs_by_4
		parameter hssi_8g_tx_pcs_clock_gate_bs_enc = "dis_bs_enc_clk_gating", // dis_bs_enc_clk_gating|en_bs_enc_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_dw_fifowr = "dis_dw_fifowr_clk_gating", // dis_dw_fifowr_clk_gating|en_dw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_fiford = "dis_fiford_clk_gating", // dis_fiford_clk_gating|en_fiford_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_sw_fifowr = "dis_sw_fifowr_clk_gating", // dis_sw_fifowr_clk_gating|en_sw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_observation_in_pld_core = "internal_refclk_b", // internal_refclk_b|internal_fifo_rd_clk|internal_sw_fifo_wr_clk|internal_dw_fifo_wr_clk|internal_tx_clk_out_gen3|internal_pipe_tx_clk_out_gen3
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_tx_pcs_data_selection_8b10b_encoder_input = "normal_data_path", // normal_data_path|gige_idle_conversion
		parameter hssi_8g_tx_pcs_dynamic_clk_switch = "dis_dyn_clk_switch", // dis_dyn_clk_switch|en_dyn_clk_switch
		parameter hssi_8g_tx_pcs_eightb_tenb_disp_ctrl = "dis_disp_ctrl", // dis_disp_ctrl|en_disp_ctrl|en_ib_disp_ctrl
		parameter hssi_8g_tx_pcs_eightb_tenb_encoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_tx_pcs_force_echar = "dis_force_echar", // dis_force_echar|en_force_echar
		parameter hssi_8g_tx_pcs_force_kchar = "dis_force_kchar", // dis_force_kchar|en_force_kchar
		parameter hssi_8g_tx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // dis_tx_clk|tx_pma_clk
		parameter hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel = "func_clk", // dis_tx_pipe_clk|func_clk
		parameter hssi_8g_tx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_tx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_tx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_tx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_tx_pcs_phfifo_write_clk_sel = "pld_tx_clk", // pld_tx_clk|tx_clk
		parameter hssi_8g_tx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_tx_pcs_prot_mode = "basic", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic|disabled_prot_mode
		parameter hssi_8g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_tx_pcs_refclk_b_clk_sel = "tx_pma_clock", // tx_pma_clock|refclk_dig
		parameter hssi_8g_tx_pcs_revloop_back_rm = "dis_rev_loopback_rx_rm", // dis_rev_loopback_rx_rm|en_rev_loopback_rx_rm
		parameter hssi_8g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_tx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_tx_pcs_tx_bitslip = "dis_tx_bitslip", // dis_tx_bitslip|en_tx_bitslip
		parameter hssi_8g_tx_pcs_tx_compliance_controlled_disparity = "dis_txcompliance", // dis_txcompliance|en_txcompliance_pipe2p0|en_txcompliance_pipe3p0
		parameter hssi_8g_tx_pcs_tx_fast_pld_reg = "dis_tx_fast_pld_reg", // dis_tx_fast_pld_reg|en_tx_fast_pld_reg
		parameter hssi_8g_tx_pcs_txclk_freerun = "dis_freerun_tx", // dis_freerun_tx|en_freerun_tx
		parameter hssi_8g_tx_pcs_txpcs_urst = "en_txpcs_urst", // dis_txpcs_urst|en_txpcs_urst
		
		// parameters for twentynm_hssi_common_pcs_pma_interface
		parameter hssi_common_pcs_pma_interface_asn_clk_enable = "false", // false|true
		parameter hssi_common_pcs_pma_interface_asn_enable = "dis_asn", // dis_asn|en_asn
		parameter hssi_common_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|pcie_gen3
		parameter hssi_common_pcs_pma_interface_bypass_early_eios = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pcie_switch = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_ltr = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_sw_done = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_ppm_lock = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_txdetectrx = "false", // false|true
		parameter hssi_common_pcs_pma_interface_cdr_control = "en_cdr_ctrl", // dis_cdr_ctrl|en_cdr_ctrl
		parameter hssi_common_pcs_pma_interface_cid_enable = "en_cid_mode", // dis_cid_mode|en_cid_mode
		parameter hssi_common_pcs_pma_interface_cp_cons_sel = "cp_cons_default", // cp_cons_master|cp_cons_slave_abv|cp_cons_slave_blw|cp_cons_default
		parameter hssi_common_pcs_pma_interface_cp_dwn_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_cp_up_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_blw|ctrl_slave_abv
		parameter hssi_common_pcs_pma_interface_data_mask_count = 16'b100111000100,
		parameter hssi_common_pcs_pma_interface_data_mask_count_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_dft_observation_clock_selection = "dft_clk_obsrv_tx0", // dft_clk_obsrv_tx0|dft_clk_obsrv_tx1|dft_clk_obsrv_tx2|dft_clk_obsrv_tx3|dft_clk_obsrv_tx4|dft_clk_obsrv_rx|dft_clk_obsrv_hclk|dft_clk_obsrv_fref|dft_clk_obsrv_clklow|dft_clk_obsrv_asn0|dft_clk_obsrv_asn1
		parameter hssi_common_pcs_pma_interface_early_eios_counter = 8'b110010,
		parameter hssi_common_pcs_pma_interface_force_freqdet = "force_freqdet_dis", // force_freqdet_dis|force1_freqdet_en|force0_freqdet_en
		parameter hssi_common_pcs_pma_interface_free_run_clk_enable = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ignore_sigdet_g23 = "false", // false|true
		parameter hssi_common_pcs_pma_interface_pc_en_counter = 7'b110111,
		parameter hssi_common_pcs_pma_interface_pc_rst_counter = 5'b10111,
		parameter hssi_common_pcs_pma_interface_pcie_hip_mode = "hip_disable", // hip_enable|hip_disable
		parameter hssi_common_pcs_pma_interface_ph_fifo_reg_mode = "phfifo_reg_mode_dis", // phfifo_reg_mode_dis|phfifo_reg_mode_en
		parameter hssi_common_pcs_pma_interface_phfifo_flush_wait = 6'b100100,
		parameter hssi_common_pcs_pma_interface_pipe_if_g3pcs = "pipe_if_8gpcs", // pipe_if_g3pcs|pipe_if_8gpcs
		parameter hssi_common_pcs_pma_interface_pma_done_counter = 18'b101010101110011000,
		parameter hssi_common_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_common_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_common_pcs_pma_interface_ppm_cnt_rst = "ppm_cnt_rst_dis", // ppm_cnt_rst_dis|ppm_cnt_rst_en
		parameter hssi_common_pcs_pma_interface_ppm_deassert_early = "deassert_early_dis", // deassert_early_dis|deassert_early_en
		parameter hssi_common_pcs_pma_interface_ppm_det_buckets = "ppm_100_bucket", // disable_prot|ppm_300_bucket|ppm_100_bucket|ppm_300_100_bucket
		parameter hssi_common_pcs_pma_interface_ppm_gen1_2_cnt = "cnt_32k", // cnt_32k|cnt_64k
		parameter hssi_common_pcs_pma_interface_ppm_post_eidle_delay = "cnt_200_cycles", // cnt_200_cycles|cnt_400_cycles
		parameter hssi_common_pcs_pma_interface_ppmsel = "ppmsel_300", // ppmsel_disable|ppmsel_5000|ppmsel_2500|ppmsel_1000|ppmsel_500|ppmsel_300|ppmsel_250|ppmsel_200|ppmsel_125|ppmsel_100|ppmsel_62p5|ppm_other
		parameter hssi_common_pcs_pma_interface_prot_mode = "disable_prot_mode", // disable_prot_mode|pipe_g12|pipe_g3|other_protocols
		parameter hssi_common_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_common_pcs_pma_interface_rxvalid_mask = "rxvalid_mask_en", // rxvalid_mask_dis|rxvalid_mask_en
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter = 12'b100111000100,
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_sim_mode = "disable", // disable|enable
		parameter hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en = "true", // false|true
		parameter hssi_common_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_common_pcs_pma_interface_testout_sel = "ppm_det_test", // ppm_det_test|asn_test|pma_pll_test|rxpmaif_test|prbs_gen_test|prbs_ver_test|uhsif_1_test|uhsif_2_test|uhsif_3_test
		parameter hssi_common_pcs_pma_interface_wait_clk_on_off_timer = 4'b100,
		parameter hssi_common_pcs_pma_interface_wait_pipe_synchronizing = 5'b10111,
		parameter hssi_common_pcs_pma_interface_wait_send_syncp_fbkp = 11'b11111010,
		
		// parameters for twentynm_hssi_common_pld_pcs_interface
		parameter hssi_common_pld_pcs_interface_dft_clk_out_en = "dft_clk_out_disable", // dft_clk_out_disable|dft_clk_out_enable
		parameter hssi_common_pld_pcs_interface_dft_clk_out_sel = "teng_rx_dft_clk", // teng_rx_dft_clk|teng_tx_dft_clk|eightg_rx_dft_clk|eightg_tx_dft_clk|pmaif_dft_clk
		parameter hssi_common_pld_pcs_interface_hrdrstctrl_en = "hrst_dis", // hrst_dis|hrst_en
		parameter hssi_common_pld_pcs_interface_pcs_testbus_block_sel = "eightg", // eightg|g3pcs|teng|krfec|pma_if
		parameter hssi_common_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_fifo_rx_pcs
		parameter hssi_fifo_rx_pcs_double_read_mode = "double_read_dis", // double_read_en|double_read_dis
		parameter hssi_fifo_rx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_fifo_tx_pcs
		parameter hssi_fifo_tx_pcs_double_write_mode = "double_write_dis", // double_write_en|double_write_dis
		parameter hssi_fifo_tx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_gen3_rx_pcs
		parameter hssi_gen3_rx_pcs_block_sync = "enable_block_sync", // bypass_block_sync|enable_block_sync
		parameter hssi_gen3_rx_pcs_block_sync_sm = "enable_blk_sync_sm", // disable_blk_sync_sm|enable_blk_sync_sm
		parameter hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn = "enable", // disable|enable
		parameter hssi_gen3_rx_pcs_lpbk_force = "lpbk_frce_dis", // lpbk_frce_dis|lpbk_frce_en
		parameter hssi_gen3_rx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_rx_pcs_rate_match_fifo = "enable_rm_fifo_600ppm", // bypass_rm_fifo|enable_rm_fifo_600ppm|enable_rm_fifo_0ppm
		parameter hssi_gen3_rx_pcs_rate_match_fifo_latency = "regular_latency", // regular_latency|low_latency
		parameter hssi_gen3_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_gen3_rx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_b4gb_par_lpbk = "b4gb_par_lpbk_dis", // b4gb_par_lpbk_dis|b4gb_par_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_force_balign = "en_force_balign", // en_force_balign|dis_force_balign
		parameter hssi_gen3_rx_pcs_rx_ins_del_one_skip = "ins_del_one_skip_en", // ins_del_one_skip_dis|ins_del_one_skip_en
		parameter hssi_gen3_rx_pcs_rx_num_fixed_pat = 4'b1000,
		parameter hssi_gen3_rx_pcs_rx_test_out_sel = "rx_test_out0", // rx_test_out0|rx_test_out1
		parameter hssi_gen3_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_gen3_tx_pcs
		parameter hssi_gen3_tx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_tx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_gen3_tx_pcs_tx_bitslip = 5'b0,
		parameter hssi_gen3_tx_pcs_tx_gbox_byp = "bypass_gbox", // bypass_gbox|enable_gbox
		
		// parameters for twentynm_hssi_krfec_rx_pcs
		parameter hssi_krfec_rx_pcs_blksync_cor_en = "detect", // detect|correct
		parameter hssi_krfec_rx_pcs_bypass_gb = "bypass_dis", // bypass_dis|bypass_en
		parameter hssi_krfec_rx_pcs_clr_ctrl = "both_enabled", // both_enabled|corr_cnt_only|uncorr_cnt_only
		parameter hssi_krfec_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_rx_pcs_dv_start = "with_blklock", // with_blksync|with_blklock
		parameter hssi_krfec_rx_pcs_err_mark_type = "err_mark_10g", // err_mark_10g|err_mark_40g
		parameter hssi_krfec_rx_pcs_error_marking_en = "err_mark_dis", // err_mark_dis|err_mark_en
		parameter hssi_krfec_rx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_krfec_rx_pcs_parity_invalid_enum = 8'b1000,
		parameter hssi_krfec_rx_pcs_parity_valid_num = 4'b100,
		parameter hssi_krfec_rx_pcs_pipeln_blksync = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_descrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errcorrect = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_ind = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_lfsr = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_loc = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_pat = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_gearbox = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_syndrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_trans_dec = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_rx_pcs_receive_order = "receive_lsb", // receive_lsb|receive_msb
		parameter hssi_krfec_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_krfec_rx_pcs_rx_testbus_sel = "overall", // overall|fast_search|fast_search_cntrs|blksync|blksync_cntrs|decoder_master_sm|decoder_master_sm_cntrs|syndrm_sm|syndrm1|syndrm2|errtrap_sm|errtrap_ind1|errtrap_ind2|errtrap_ind3|errtrap_ind4|errtrap_ind5|errtrap_loc|errtrap_pat1|errtrap_pat2|errtrap_pat3|errtrap_pat4|decoder_rd_sm|gb_and_trans
		parameter hssi_krfec_rx_pcs_signal_ok_en = "sig_ok_dis", // sig_ok_dis|sig_ok_en
		parameter hssi_krfec_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_krfec_tx_pcs
		parameter hssi_krfec_tx_pcs_burst_err = "burst_err_dis", // burst_err_dis|burst_err_en
		parameter hssi_krfec_tx_pcs_burst_err_len = "burst_err_len1", // burst_err_len1|burst_err_len2|burst_err_len3|burst_err_len4|burst_err_len5|burst_err_len6|burst_err_len7|burst_err_len8|burst_err_len9|burst_err_len10|burst_err_len11|burst_err_len12|burst_err_len13|burst_err_len14|burst_err_len15|burst_err_len16
		parameter hssi_krfec_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_tx_pcs_enc_frame_query = "enc_query_dis", // enc_query_dis|enc_query_en
		parameter hssi_krfec_tx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_encoder = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_scrambler = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_krfec_tx_pcs_transcode_err = "trans_err_dis", // trans_err_dis|trans_err_en
		parameter hssi_krfec_tx_pcs_transmit_order = "transmit_lsb", // transmit_lsb|transmit_msb
		parameter hssi_krfec_tx_pcs_tx_testbus_sel = "overall", // overall|encoder1|encoder2|scramble1|scramble2|scramble3|gearbox
		
		// parameters for twentynm_hssi_pipe_gen1_2
		parameter hssi_pipe_gen1_2_elec_idle_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_error_replace_pad = "replace_edb", // replace_edb|replace_pad
		parameter hssi_pipe_gen1_2_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_pipe_gen1_2_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen1_2_phystatus_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_phystatus_rst_toggle = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen1_2_pipe_byte_de_serializer_en = "dont_care_bds", // dis_bds|en_bds_by_2|dont_care_bds
		parameter hssi_pipe_gen1_2_prot_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|basic|disabled_prot_mode
		parameter hssi_pipe_gen1_2_reconfig_settings = "{}", // 
		parameter hssi_pipe_gen1_2_rx_pipe_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_pipe_gen1_2_rxdetect_bypass = "dis_rxdetect_bypass", // dis_rxdetect_bypass|en_rxdetect_bypass
		parameter hssi_pipe_gen1_2_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen1_2_tx_pipe_enable = "dis_pipe_tx", // dis_pipe_tx|en_pipe_tx|en_pipe3_tx
		parameter hssi_pipe_gen1_2_txswing = "dis_txswing", // dis_txswing|en_txswing
		
		// parameters for twentynm_hssi_pipe_gen3
		parameter hssi_pipe_gen3_bypass_rx_detection_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_rx_preset = 3'b0,
		parameter hssi_pipe_gen3_bypass_rx_preset_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_tx_coefficent = 18'b0,
		parameter hssi_pipe_gen3_bypass_tx_coefficent_enable = "false", // false|true
		parameter hssi_pipe_gen3_elecidle_delay_g3 = 3'b110,
		parameter hssi_pipe_gen3_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen3_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|disable_pcs
		parameter hssi_pipe_gen3_phy_status_delay_g12 = 3'b101,
		parameter hssi_pipe_gen3_phy_status_delay_g3 = 3'b101,
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g12 = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g3 = "dis_phystatus_rst_toggle_g3", // dis_phystatus_rst_toggle_g3|en_phystatus_rst_toggle_g3
		parameter hssi_pipe_gen3_rate_match_pad_insertion = "dis_rm_fifo_pad_ins", // dis_rm_fifo_pad_ins|en_rm_fifo_pad_ins
		parameter hssi_pipe_gen3_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen3_test_out_sel = "disable_test_out", // tx_test_out|rx_test_out|pipe_test_out1|pipe_test_out2|pipe_test_out3|pipe_ctrl_test_out|disable_test_out
		
		// parameters for twentynm_hssi_rx_pcs_pma_interface
		parameter hssi_rx_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|ten_g_pcs|direct_pld
		parameter hssi_rx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pcs_pma_interface_clkslip_sel = "pld", // pld|slip_eight_g_pcs
		parameter hssi_rx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pcs_pma_interface_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_rx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_rx_pcs_pma_interface_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_rx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_rx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_rx_pcs_pma_interface_prbs_ver = "prbs_off", // prbs_off|prbs_31|prbs_15|prbs_23|prbs_9|prbs_7
		parameter hssi_rx_pcs_pma_interface_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion = "rx_dyn_polinv_dis", // rx_dyn_polinv_dis|rx_dyn_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_lpbk_en = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok = "unforce_sig_ok", // unforce_sig_ok|force_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mask = "prbsmask128", // prbsmask128|prbsmask256|prbsmask512|prbsmask1024
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mode = "teng_mode", // teng_mode|eightg_mode
		parameter hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel = "sel_sig_det", // sel_sig_det|sel_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_static_polarity_inversion = "rx_stat_polinv_dis", // rx_stat_polinv_dis|rx_stat_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en = "uhsif_lpbk_dis", // uhsif_lpbk_dis|uhsif_lpbk_en
		parameter hssi_rx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_rx_pld_pcs_interface
		parameter hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx = "enable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx = "pma_64b_rx", // pma_32b_rx|pma_40b_rx|pma_64b_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_baser_mode_rx|interlaken_mode_rx|sfis_mode_rx|teng_sdi_mode_rx|basic_mode_rx|test_prp_mode_rx|test_prp_krfec_mode_rx|teng_1588_mode_rx|teng_baser_krfec_mode_rx|teng_1588_krfec_mode_rx|basic_krfec_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx = "disabled_prot_mode_rx", // pipe_g1_rx|pipe_g2_rx|pipe_g3_rx|cpri_rx|cpri_rx_tx_rx|gige_rx|gige_1588_rx|basic_rm_enable_rx|basic_rm_disable_rx|disabled_prot_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcie_g1_capable_rx|pcie_g2_capable_rx|pcie_g3_capable_rx|gige_rx|teng_baser_rx|teng_basekr_krfec_rx|fortyg_basekr_krfec_rx|cpri_8b10b_rx|interlaken_rx|sfis_rx|teng_sdi_rx|gige_1588_rx|teng_1588_baser_rx|teng_1588_basekr_krfec_rx|basic_8gpcs_rm_enable_rx|basic_8gpcs_rm_disable_rx|basic_10gpcs_rx|basic_10gpcs_krfec_rx|pcs_direct_rx|prp_rx|prp_krfec_rx|prbs_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx = "teng_mode_rx", // teng_mode_rx|non_teng_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_basekr_mode_rx|fortyg_basekr_mode_rx|teng_1588_basekr_mode_rx|basic_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|eightg_and_g3_pld_fifo_mode_rx|eightg_and_g3_reg_mode_rx|eightg_and_g3_reg_mode_hip_rx|teng_pld_fifo_mode_rx|teng_reg_mode_rx|teng_and_krfec_pld_fifo_mode_rx|teng_and_krfec_reg_mode_rx|pcs_direct_reg_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_block_sel = "pcs_direct", // eightg|teng|pcs_direct
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_rx_clk|pma_rx_clk_user
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_sel = "pld_rx_clk", // pld_rx_clk|pcs_rx_clk
		parameter hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en = "hip_rx_enable", // hip_rx_enable|hip_rx_disable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_rx_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_tx_pcs_pma_interface
		parameter hssi_tx_pcs_pma_interface_bypass_pma_txelecidle = "false", // false|true
		parameter hssi_tx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pcs_pma_interface_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx = "other_prot_mode", // pipe_g12|pipe_g3|other_prot_mode
		parameter hssi_tx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_tx_pcs_pma_interface_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_tx_pcs_pma_interface_pmagate_en = "pmagate_dis", // pmagate_dis|pmagate_en
		parameter hssi_tx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_tx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_tx_pcs_pma_interface_prbs_gen_pat = "prbs_gen_dis", // prbs_gen_dis|prbs_31|prbs_23|prbs_15|prbs_9|prbs_7
		parameter hssi_tx_pcs_pma_interface_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_tx_pcs_pma_interface_sq_wave_num = "sq_wave_4", // sq_wave_1|sq_wave_4|sq_wave_8|sq_wave_6|sq_wave_default
		parameter hssi_tx_pcs_pma_interface_sqwgen_clken = "sqwgen_clk_dis", // sqwgen_clk_dis|sqwgen_clk_en
		parameter hssi_tx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion = "tx_dyn_polinv_dis", // tx_dyn_polinv_dis|tx_dyn_polinv_en
		parameter hssi_tx_pcs_pma_interface_tx_pma_data_sel = "pld_dir", // pld_dir|pcie_gen3|eight_g_pcs|ten_g_pcs|prbs_pat|sq_wave_pat|block_sel_default|registered_uhsif_dat|directed_uhsif_dat
		parameter hssi_tx_pcs_pma_interface_tx_static_polarity_inversion = "tx_stat_polinv_dis", // tx_stat_polinv_dis|tx_stat_polinv_en
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock = "uhsif_filt_stepsz_b4lock_4", // uhsif_filt_stepsz_b4lock_2|uhsif_filt_stepsz_b4lock_4|uhsif_filt_stepsz_b4lock_6|uhsif_filt_stepsz_b4lock_8
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value = 4'b1011,
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock = "uhsif_filt_cntthr_b4lock_16", // uhsif_filt_cntthr_b4lock_8|uhsif_filt_cntthr_b4lock_16|uhsif_filt_cntthr_b4lock_24|uhsif_filt_cntthr_b4lock_32
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period = "uhsif_dcn_test_period_4", // uhsif_dcn_test_period_4|uhsif_dcn_test_period_8|uhsif_dcn_test_period_12|uhsif_dcn_test_period_16
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable = "uhsif_dcn_test_mode_disable", // uhsif_dcn_test_mode_enable|uhsif_dcn_test_mode_disable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh = "uhsif_dzt_cnt_thr_4", // uhsif_dzt_cnt_thr_2|uhsif_dzt_cnt_thr_4|uhsif_dzt_cnt_thr_6|uhsif_dzt_cnt_thr_8
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable = "uhsif_dzt_enable", // uhsif_dzt_disable|uhsif_dzt_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window = "uhsif_dzt_obr_win_32", // uhsif_dzt_obr_win_16|uhsif_dzt_obr_win_32|uhsif_dzt_obr_win_48|uhsif_dzt_obr_win_64
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size = "uhsif_dzt_skipsz_8", // uhsif_dzt_skipsz_4|uhsif_dzt_skipsz_8|uhsif_dzt_skipsz_12|uhsif_dzt_skipsz_16
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel = "uhsif_index_internal", // uhsif_index_internal|uhsif_index_cram
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin = "uhsif_dcn_margin_4", // uhsif_dcn_margin_2|uhsif_dcn_margin_3|uhsif_dcn_margin_4|uhsif_dcn_margin_5
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value = 8'b10000000,
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control = "uhsif_dft_dz_det_val_0", // uhsif_dft_dz_det_val_0|uhsif_dft_dz_det_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control = "uhsif_dft_up_val_0", // uhsif_dft_up_val_0|uhsif_dft_up_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_enable = "uhsif_disable", // uhsif_disable|uhsif_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock = "uhsif_lkd_segsz_aflock_2048", // uhsif_lkd_segsz_aflock_512|uhsif_lkd_segsz_aflock_1024|uhsif_lkd_segsz_aflock_2048|uhsif_lkd_segsz_aflock_4096
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock = "uhsif_lkd_segsz_b4lock_32", // uhsif_lkd_segsz_b4lock_16|uhsif_lkd_segsz_b4lock_32|uhsif_lkd_segsz_b4lock_64|uhsif_lkd_segsz_b4lock_128
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value = 4'b11,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value = 4'b11,
		
		// parameters for twentynm_hssi_tx_pld_pcs_interface
		parameter hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx = "enable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx = "pma_64b_tx", // pma_32b_tx|pma_40b_tx|pma_64b_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_baser_mode_tx|interlaken_mode_tx|sfis_mode_tx|teng_sdi_mode_tx|basic_mode_tx|test_prp_mode_tx|test_prp_krfec_mode_tx|teng_1588_mode_tx|teng_baser_krfec_mode_tx|teng_1588_krfec_mode_tx|basic_krfec_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx = "disabled_prot_mode_tx", // pipe_g1_tx|pipe_g2_tx|pipe_g3_tx|cpri_tx|cpri_rx_tx_tx|gige_tx|gige_1588_tx|basic_tx|disabled_prot_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcie_g1_capable_tx|pcie_g2_capable_tx|pcie_g3_capable_tx|gige_tx|teng_baser_tx|teng_basekr_krfec_tx|fortyg_basekr_krfec_tx|cpri_8b10b_tx|interlaken_tx|sfis_tx|teng_sdi_tx|gige_1588_tx|teng_1588_baser_tx|teng_1588_basekr_krfec_tx|basic_8gpcs_tx|basic_10gpcs_tx|basic_10gpcs_krfec_tx|pcs_direct_tx|uhsif_tx|prp_tx|prp_krfec_tx|prbs_tx|sqwave_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx = "teng_mode_tx", // teng_mode_tx|non_teng_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_basekr_mode_tx|fortyg_basekr_mode_tx|teng_1588_basekr_mode_tx|basic_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|eightg_and_g3_pld_fifo_mode_tx|eightg_and_g3_reg_mode_tx|eightg_and_g3_reg_mode_hip_tx|eightg_and_g3_fastreg_mode_tx|teng_pld_fifo_mode_tx|teng_reg_mode_tx|teng_fastreg_mode_tx|teng_and_krfec_pld_fifo_mode_tx|teng_and_krfec_reg_mode_tx|teng_and_krfec_fastreg_mode_tx|pcs_direct_fastreg_mode_tx|uhsif_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_tx_clk|pma_tx_clk_user
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_source = "teng", // eightg|teng|pma_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_data_source = "hip_disable", // hip_disable|hip_enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en = "delay1_clk_disable", // delay1_clk_enable|delay1_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel = "pld_tx_clk", // pld_tx_clk|pcs_tx_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl = "delay1_path0", // delay1_path0|delay1_path1|delay1_path2|delay1_path3|delay1_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel = "one_ff_delay", // one_ff_delay|two_ff_delay
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en = "delay2_clk_disable", // delay2_clk_enable|delay2_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl = "delay2_path0", // delay2_path0|delay2_path1|delay2_path2|delay2_path3|delay2_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_tx_pld_pcs_interface_reconfig_settings = "{}" // 
	//PARAM_LIST_END
	)
	(
	//PORT_LIST_START
		input wire	[8:0]	in_avmmaddress,
		input wire		in_avmmclk,
		input wire		in_avmmread,
		input wire		in_avmmrstn,
		input wire		in_avmmwrite,
		input wire	[7:0]	in_avmmwritedata,
		input wire	[4:0]	in_bond_pcs10g_in_bot,
		input wire	[4:0]	in_bond_pcs10g_in_top,
		input wire	[12:0]	in_bond_pcs8g_in_bot,
		input wire	[12:0]	in_bond_pcs8g_in_top,
		input wire	[11:0]	in_bond_pmaif_in_bot,
		input wire	[11:0]	in_bond_pmaif_in_top,
		input wire	[63:0]	in_hip_tx_data,
		input wire		in_iocsr_clk,
		input wire	[5:0]	in_iocsr_config,
		input wire		in_iocsr_rdy,
		input wire		in_iocsr_rdy_dly,
		input wire		in_pld_10g_krfec_rx_clr_errblk_cnt,
		input wire		in_pld_10g_krfec_rx_pld_rst_n,
		input wire		in_pld_10g_krfec_tx_pld_rst_n,
		input wire		in_pld_10g_rx_align_clr,
		input wire		in_pld_10g_rx_clr_ber_count,
		input wire		in_pld_10g_rx_rd_en,
		input wire	[6:0]	in_pld_10g_tx_bitslip,
		input wire		in_pld_10g_tx_burst_en,
		input wire		in_pld_10g_tx_data_valid,
		input wire	[1:0]	in_pld_10g_tx_diag_status,
		input wire		in_pld_10g_tx_wordslip,
		input wire		in_pld_8g_a1a2_size,
		input wire		in_pld_8g_bitloc_rev_en,
		input wire		in_pld_8g_byte_rev_en,
		input wire	[2:0]	in_pld_8g_eidleinfersel,
		input wire		in_pld_8g_encdt,
		input wire		in_pld_8g_g3_rx_pld_rst_n,
		input wire		in_pld_8g_g3_tx_pld_rst_n,
		input wire		in_pld_8g_rddisable_tx,
		input wire		in_pld_8g_rdenable_rx,
		input wire		in_pld_8g_refclk_dig2,
		input wire		in_pld_8g_rxpolarity,
		input wire	[4:0]	in_pld_8g_tx_boundary_sel,
		input wire		in_pld_8g_wrdisable_rx,
		input wire		in_pld_8g_wrenable_tx,
		input wire		in_pld_atpg_los_en_n,
		input wire		in_pld_bitslip,
		input wire	[17:0]	in_pld_g3_current_coeff,
		input wire	[2:0]	in_pld_g3_current_rxpreset,
		input wire		in_pld_ltr,
		input wire		in_pld_mem_krfec_atpg_rst_n,
		input wire		in_pld_partial_reconfig,
		input wire		in_pld_pcs_refclk_dig,
		input wire		in_pld_pma_adapt_start,
		input wire		in_pld_pma_csr_test_dis,
		input wire		in_pld_pma_early_eios,
		input wire	[5:0]	in_pld_pma_eye_monitor,
		input wire		in_pld_pma_ltd_b,
		input wire		in_pld_pma_nrpi_freeze,
		input wire	[1:0]	in_pld_pma_pcie_switch,
		input wire		in_pld_pma_ppm_lock,
		input wire	[4:0]	in_pld_pma_reserved_out,
		input wire		in_pld_pma_rs_lpbk_b,
		input wire		in_pld_pma_rx_qpi_pullup,
		input wire		in_pld_pma_rxpma_rstb,
		input wire		in_pld_pma_tx_bitslip,
		input wire		in_pld_pma_tx_bonding_rstb,
		input wire		in_pld_pma_tx_qpi_pulldn,
		input wire		in_pld_pma_tx_qpi_pullup,
		input wire		in_pld_pma_txdetectrx,
		input wire		in_pld_pma_txpma_rstb,
		input wire		in_pld_pmaif_rx_pld_rst_n,
		input wire		in_pld_pmaif_rxclkslip,
		input wire		in_pld_pmaif_tx_pld_rst_n,
		input wire		in_pld_polinv_rx,
		input wire		in_pld_polinv_tx,
		input wire	[1:0]	in_pld_rate,
		input wire	[9:0]	in_pld_reserved_in,
		input wire		in_pld_rx_clk,
		input wire		in_pld_rx_prbs_err_clr,
		input wire		in_pld_scan_mode_n,
		input wire		in_pld_scan_shift_n,
		input wire		in_pld_syncsm_en,
		input wire		in_pld_tx_clk,
		input wire	[17:0]	in_pld_tx_control,
		input wire	[127:0]	in_pld_tx_data,
		input wire		in_pld_txelecidle,
		input wire		in_pld_uhsif_tx_clk,
		input wire		in_pma_adapt_done,
		input wire		in_pma_clklow,
		input wire		in_pma_fref,
		input wire		in_pma_hclk,
		input wire	[1:0]	in_pma_pcie_sw_done,
		input wire		in_pma_pfdmode_lock,
		input wire	[4:0]	in_pma_reserved_in,
		input wire		in_pma_rx_clkdiv_user,
		input wire		in_pma_rx_detect_valid,
		input wire		in_pma_rx_found,
		input wire		in_pma_rx_pma_clk,
		input wire	[63:0]	in_pma_rx_pma_data,
		input wire		in_pma_rx_signal_ok,
		input wire		in_pma_rxpll_lock,
		input wire		in_pma_signal_det,
		input wire	[7:0]	in_pma_testbus,
		input wire		in_pma_tx_clkdiv_user,
		input wire		in_pma_tx_pma_clk,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen1_2,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen3,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pld_pcs_interface,
		output wire		out_blockselect_hssi_10g_rx_pcs,
		output wire		out_blockselect_hssi_10g_tx_pcs,
		output wire		out_blockselect_hssi_8g_rx_pcs,
		output wire		out_blockselect_hssi_8g_tx_pcs,
		output wire		out_blockselect_hssi_common_pcs_pma_interface,
		output wire		out_blockselect_hssi_common_pld_pcs_interface,
		output wire		out_blockselect_hssi_fifo_rx_pcs,
		output wire		out_blockselect_hssi_fifo_tx_pcs,
		output wire		out_blockselect_hssi_gen3_rx_pcs,
		output wire		out_blockselect_hssi_gen3_tx_pcs,
		output wire		out_blockselect_hssi_krfec_rx_pcs,
		output wire		out_blockselect_hssi_krfec_tx_pcs,
		output wire		out_blockselect_hssi_pipe_gen1_2,
		output wire		out_blockselect_hssi_pipe_gen3,
		output wire		out_blockselect_hssi_rx_pcs_pma_interface,
		output wire		out_blockselect_hssi_rx_pld_pcs_interface,
		output wire		out_blockselect_hssi_tx_pcs_pma_interface,
		output wire		out_blockselect_hssi_tx_pld_pcs_interface,
		output wire	[4:0]	out_bond_pcs10g_out_bot,
		output wire	[4:0]	out_bond_pcs10g_out_top,
		output wire	[12:0]	out_bond_pcs8g_out_bot,
		output wire	[12:0]	out_bond_pcs8g_out_top,
		output wire	[11:0]	out_bond_pmaif_out_bot,
		output wire	[11:0]	out_bond_pmaif_out_top,
		output wire	[2:0]	out_hip_clk_out,
		output wire	[7:0]	out_hip_ctrl_out,
		output wire		out_hip_iocsr_rdy,
		output wire		out_hip_iocsr_rdy_dly,
		output wire		out_hip_nfrzdrv,
		output wire		out_hip_npor,
		output wire	[50:0]	out_hip_rx_data,
		output wire		out_hip_usermode,
		output wire		out_pld_10g_krfec_rx_blk_lock,
		output wire	[1:0]	out_pld_10g_krfec_rx_diag_data_status,
		output wire		out_pld_10g_krfec_rx_frame,
		output wire		out_pld_10g_krfec_tx_frame,
		output wire		out_pld_10g_rx_align_val,
		output wire		out_pld_10g_rx_crc32_err,
		output wire		out_pld_10g_rx_data_valid,
		output wire		out_pld_10g_rx_empty,
		output wire		out_pld_10g_rx_fifo_del,
		output wire		out_pld_10g_rx_fifo_insert,
		output wire	[4:0]	out_pld_10g_rx_fifo_num,
		output wire		out_pld_10g_rx_frame_lock,
		output wire		out_pld_10g_rx_hi_ber,
		output wire		out_pld_10g_rx_oflw_err,
		output wire		out_pld_10g_rx_pempty,
		output wire		out_pld_10g_rx_pfull,
		output wire		out_pld_10g_tx_burst_en_exe,
		output wire		out_pld_10g_tx_empty,
		output wire	[3:0]	out_pld_10g_tx_fifo_num,
		output wire		out_pld_10g_tx_full,
		output wire		out_pld_10g_tx_pempty,
		output wire		out_pld_10g_tx_pfull,
		output wire		out_pld_10g_tx_wordslip_exe,
		output wire	[3:0]	out_pld_8g_a1a2_k1k2_flag,
		output wire		out_pld_8g_empty_rmf,
		output wire		out_pld_8g_empty_rx,
		output wire		out_pld_8g_empty_tx,
		output wire		out_pld_8g_full_rmf,
		output wire		out_pld_8g_full_rx,
		output wire		out_pld_8g_full_tx,
		output wire		out_pld_8g_rxelecidle,
		output wire		out_pld_8g_signal_detect_out,
		output wire	[4:0]	out_pld_8g_wa_boundary,
		output wire		out_pld_krfec_tx_alignment,
		output wire		out_pld_pcs_rx_clk_out,
		output wire		out_pld_pcs_tx_clk_out,
		output wire		out_pld_pma_adapt_done,
		output wire		out_pld_pma_clkdiv_rx_user,
		output wire		out_pld_pma_clkdiv_tx_user,
		output wire		out_pld_pma_clklow,
		output wire		out_pld_pma_fref,
		output wire		out_pld_pma_hclk,
		output wire	[1:0]	out_pld_pma_pcie_sw_done,
		output wire		out_pld_pma_pfdmode_lock,
		output wire	[4:0]	out_pld_pma_reserved_in,
		output wire		out_pld_pma_rx_clk_out,
		output wire		out_pld_pma_rx_detect_valid,
		output wire		out_pld_pma_rx_found,
		output wire		out_pld_pma_rxpll_lock,
		output wire		out_pld_pma_signal_ok,
		output wire	[7:0]	out_pld_pma_testbus,
		output wire		out_pld_pma_tx_clk_out,
		output wire		out_pld_pmaif_mask_tx_pll,
		output wire	[9:0]	out_pld_reserved_out,
		output wire	[19:0]	out_pld_rx_control,
		output wire	[127:0]	out_pld_rx_data,
		output wire		out_pld_rx_prbs_done,
		output wire		out_pld_rx_prbs_err,
		output wire	[19:0]	out_pld_test_data,
		output wire		out_pld_uhsif_lock,
		output wire		out_pld_uhsif_tx_clk_out,
		output wire		out_pma_adapt_start,
		output wire		out_pma_atpg_los_en_n,
		output wire		out_pma_csr_test_dis,
		output wire	[17:0]	out_pma_current_coeff,
		output wire	[2:0]	out_pma_current_rxpreset,
		output wire		out_pma_early_eios,
		output wire	[5:0]	out_pma_eye_monitor,
		output wire	[1:0]	out_pma_interface_select,
		output wire		out_pma_ltd_b,
		output wire		out_pma_ltr,
		output wire		out_pma_nfrzdrv,
		output wire		out_pma_nrpi_freeze,
		output wire	[1:0]	out_pma_pcie_switch,
		output wire		out_pma_ppm_lock,
		output wire	[4:0]	out_pma_reserved_out,
		output wire		out_pma_rs_lpbk_b,
		output wire		out_pma_rx_clkslip,
		output wire		out_pma_rx_qpi_pullup,
		output wire		out_pma_rxpma_rstb,
		output wire		out_pma_scan_mode_n,
		output wire		out_pma_scan_shift_n,
		output wire		out_pma_tx_bitslip,
		output wire		out_pma_tx_bonding_rstb,
		output wire		out_pma_tx_elec_idle,
		output wire	[63:0]	out_pma_tx_pma_data,
		output wire		out_pma_tx_qpi_pulldn,
		output wire		out_pma_tx_qpi_pullup,
		output wire		out_pma_tx_txdetectrx,
		output wire		out_pma_txpma_rstb
	//PORT_LIST_END
	);
	//wire declarations
	
	// wires for module twentynm_hssi_fifo_tx_pcs
	wire	[7:0]	w_hssi_fifo_tx_pcs_avmmreaddata;
	wire		w_hssi_fifo_tx_pcs_blockselect;
	wire	[72:0]	w_hssi_fifo_tx_pcs_data_out_10g;
	wire	[63:0]	w_hssi_fifo_tx_pcs_data_out_8g_phase_comp;
	
	// wires for module twentynm_hssi_gen3_rx_pcs
	wire	[7:0]	w_hssi_gen3_rx_pcs_avmmreaddata;
	wire		w_hssi_gen3_rx_pcs_blk_algnd_int;
	wire		w_hssi_gen3_rx_pcs_blk_start;
	wire		w_hssi_gen3_rx_pcs_blockselect;
	wire		w_hssi_gen3_rx_pcs_clkcomp_delete_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_insert_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_overfl_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_undfl_int;
	wire	[31:0]	w_hssi_gen3_rx_pcs_data_out;
	wire		w_hssi_gen3_rx_pcs_data_valid;
	wire		w_hssi_gen3_rx_pcs_ei_det_int;
	wire		w_hssi_gen3_rx_pcs_ei_partial_det_int;
	wire		w_hssi_gen3_rx_pcs_err_decode_int;
	wire		w_hssi_gen3_rx_pcs_i_det_int;
	wire		w_hssi_gen3_rx_pcs_lpbk_blk_start;
	wire	[33:0]	w_hssi_gen3_rx_pcs_lpbk_data;
	wire		w_hssi_gen3_rx_pcs_lpbk_data_valid;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk;
	wire	[39:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n;
	wire		w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int;
	wire	[19:0]	w_hssi_gen3_rx_pcs_rx_test_out;
	wire	[1:0]	w_hssi_gen3_rx_pcs_sync_hdr;
	
	// wires for module twentynm_hssi_krfec_tx_pcs
	wire	[7:0]	w_hssi_krfec_tx_pcs_avmmreaddata;
	wire		w_hssi_krfec_tx_pcs_blockselect;
	wire		w_hssi_krfec_tx_pcs_tx_alignment;
	wire	[63:0]	w_hssi_krfec_tx_pcs_tx_data_out;
	wire		w_hssi_krfec_tx_pcs_tx_frame;
	wire	[19:0]	w_hssi_krfec_tx_pcs_tx_test_data;
	
	// wires for module twentynm_hssi_krfec_rx_pcs
	wire	[7:0]	w_hssi_krfec_rx_pcs_avmmreaddata;
	wire		w_hssi_krfec_rx_pcs_blockselect;
	wire		w_hssi_krfec_rx_pcs_rx_block_lock;
	wire	[9:0]	w_hssi_krfec_rx_pcs_rx_control_out;
	wire	[63:0]	w_hssi_krfec_rx_pcs_rx_data_out;
	wire	[1:0]	w_hssi_krfec_rx_pcs_rx_data_status;
	wire		w_hssi_krfec_rx_pcs_rx_data_valid_out;
	wire		w_hssi_krfec_rx_pcs_rx_frame;
	wire		w_hssi_krfec_rx_pcs_rx_signal_ok_out;
	
	// wires for module twentynm_hssi_rx_pld_pcs_interface
	wire	[7:0]	w_hssi_rx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_rx_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_hip_rx_ctrl;
	wire	[50:0]	w_hssi_rx_pld_pcs_interface_hip_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
	wire	[3:0]	w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary;
	wire		w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_pld_rx_control;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_pld_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
	
	// wires for module twentynm_hssi_common_pld_pcs_interface
	wire	[7:0]	w_hssi_common_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_common_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_hip_cmn_clk;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_hip_cmn_ctrl;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
	wire		w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_hip_npor;
	wire		w_hssi_common_pld_pcs_interface_hip_usermode;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n;
	wire	[17:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel;
	wire		w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_clklow;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_fref;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_hclk;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_pld_pma_reserved_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
	wire	[7:0]	w_hssi_common_pld_pcs_interface_pld_pma_testbus;
	wire		w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
	wire	[9:0]	w_hssi_common_pld_pcs_interface_pld_reserved_out;
	wire	[19:0]	w_hssi_common_pld_pcs_interface_pld_test_data;
	wire		w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
	wire		w_hssi_common_pld_pcs_interface_scan_mode_n;
	
	// wires for module twentynm_hssi_10g_rx_pcs
	wire	[7:0]	w_hssi_10g_rx_pcs_avmmreaddata;
	wire		w_hssi_10g_rx_pcs_blockselect;
	wire		w_hssi_10g_rx_pcs_rx_align_val;
	wire		w_hssi_10g_rx_pcs_rx_blk_lock;
	wire		w_hssi_10g_rx_pcs_rx_clk_out;
	wire		w_hssi_10g_rx_pcs_rx_clk_out_pld_if;
	wire	[19:0]	w_hssi_10g_rx_pcs_rx_control;
	wire		w_hssi_10g_rx_pcs_rx_crc32_err;
	wire	[127:0]	w_hssi_10g_rx_pcs_rx_data;
	wire		w_hssi_10g_rx_pcs_rx_data_valid;
	wire		w_hssi_10g_rx_pcs_rx_dft_clk_out;
	wire	[1:0]	w_hssi_10g_rx_pcs_rx_diag_status;
	wire		w_hssi_10g_rx_pcs_rx_empty;
	wire		w_hssi_10g_rx_pcs_rx_fec_clk;
	wire		w_hssi_10g_rx_pcs_rx_fifo_del;
	wire		w_hssi_10g_rx_pcs_rx_fifo_insert;
	wire	[4:0]	w_hssi_10g_rx_pcs_rx_fifo_num;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_clk;
	wire	[73:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_data;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_en;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_ptr;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_frame_lock;
	wire		w_hssi_10g_rx_pcs_rx_hi_ber;
	wire		w_hssi_10g_rx_pcs_rx_master_clk;
	wire		w_hssi_10g_rx_pcs_rx_master_clk_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_oflw_err;
	wire		w_hssi_10g_rx_pcs_rx_pempty;
	wire		w_hssi_10g_rx_pcs_rx_pfull;
	wire		w_hssi_10g_rx_pcs_rx_random_err;
	wire		w_hssi_10g_rx_pcs_rx_rx_frame;
	
	// wires for module twentynm_hssi_tx_pld_pcs_interface
	wire	[7:0]	w_hssi_tx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_tx_pld_pcs_interface_blockselect;
	wire		w_hssi_tx_pld_pcs_interface_hip_tx_clk;
	wire	[6:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en;
	wire	[17:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control;
	wire	[8:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg;
	wire	[127:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start;
	wire	[4:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle;
	wire	[2:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
	wire		w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
	
	// wires for module twentynm_hssi_tx_pcs_pma_interface
	wire	[7:0]	w_hssi_tx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_tx_pcs_pma_interface_blockselect;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out;
	wire	[4:0]	w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk;
	wire		w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_pma_tx_pma_data;
	wire		w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_1;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_2;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_3;
	
	// wires for module twentynm_hssi_rx_pcs_pma_interface
	wire	[7:0]	w_hssi_rx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_rx_pcs_pma_interface_blockselect;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni;
	wire	[31:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok;
	wire		w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk;
	wire	[5:0]	w_hssi_rx_pcs_pma_interface_pma_eye_monitor;
	wire		w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
	wire		w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test;
	
	// wires for module twentynm_hssi_10g_tx_pcs
	wire	[7:0]	w_hssi_10g_tx_pcs_avmmreaddata;
	wire		w_hssi_10g_tx_pcs_blockselect;
	wire		w_hssi_10g_tx_pcs_distdwn_out_dv;
	wire		w_hssi_10g_tx_pcs_distdwn_out_rden;
	wire		w_hssi_10g_tx_pcs_distdwn_out_wren;
	wire		w_hssi_10g_tx_pcs_distup_out_dv;
	wire		w_hssi_10g_tx_pcs_distup_out_rden;
	wire		w_hssi_10g_tx_pcs_distup_out_wren;
	wire		w_hssi_10g_tx_pcs_tx_burst_en_exe;
	wire		w_hssi_10g_tx_pcs_tx_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pma_if;
	wire	[8:0]	w_hssi_10g_tx_pcs_tx_control_out_krfec;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_data_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_data_valid_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_dft_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_empty;
	wire		w_hssi_10g_tx_pcs_tx_fec_clk;
	wire	[3:0]	w_hssi_10g_tx_pcs_tx_fifo_num;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_rd_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_clk;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_en;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_frame;
	wire		w_hssi_10g_tx_pcs_tx_full;
	wire		w_hssi_10g_tx_pcs_tx_master_clk;
	wire		w_hssi_10g_tx_pcs_tx_master_clk_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_pempty;
	wire		w_hssi_10g_tx_pcs_tx_pfull;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_data;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_gating_val;
	wire	[19:0]	w_hssi_10g_tx_pcs_tx_test_data;
	wire		w_hssi_10g_tx_pcs_tx_wordslip_exe;
	
	// wires for module twentynm_hssi_8g_tx_pcs
	wire	[7:0]	w_hssi_8g_tx_pcs_avmmreaddata;
	wire		w_hssi_8g_tx_pcs_blockselect;
	wire		w_hssi_8g_tx_pcs_clk_out;
	wire		w_hssi_8g_tx_pcs_clk_out_gen3;
	wire	[19:0]	w_hssi_8g_tx_pcs_dataout;
	wire		w_hssi_8g_tx_pcs_dyn_clk_switch_n;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn;
	wire		w_hssi_8g_tx_pcs_g3_tx_pma_rstn;
	wire	[2:0]	w_hssi_8g_tx_pcs_non_gray_eidleinfersel;
	wire		w_hssi_8g_tx_pcs_ph_fifo_overflow;
	wire		w_hssi_8g_tx_pcs_ph_fifo_underflow;
	wire		w_hssi_8g_tx_pcs_phfifo_txdeemph;
	wire	[2:0]	w_hssi_8g_tx_pcs_phfifo_txmargin;
	wire		w_hssi_8g_tx_pcs_phfifo_txswing;
	wire		w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out;
	wire	[1:0]	w_hssi_8g_tx_pcs_pipe_power_down_out;
	wire		w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3;
	wire		w_hssi_8g_tx_pcs_pmaif_asn_rstn;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_refclk_b;
	wire		w_hssi_8g_tx_pcs_refclk_b_reset;
	wire		w_hssi_8g_tx_pcs_rxpolarity_int;
	wire		w_hssi_8g_tx_pcs_soft_reset_wclk1_n;
	wire		w_hssi_8g_tx_pcs_sw_fifo_wr_clk;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_blk_start_out;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_ctrlplane_testbus;
	wire	[31:0]	w_hssi_8g_tx_pcs_tx_data_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_data_valid_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_datak_out;
	wire		w_hssi_8g_tx_pcs_tx_detect_rxloopback_int;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_tx_pipe_clk;
	wire		w_hssi_8g_tx_pcs_tx_pipe_electidle;
	wire		w_hssi_8g_tx_pcs_tx_pipe_soft_reset;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_sync_hdr_out;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_testbus;
	wire		w_hssi_8g_tx_pcs_txcompliance_out;
	wire		w_hssi_8g_tx_pcs_txelecidle_out;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk;
	wire	[63:0]	w_hssi_8g_tx_pcs_wr_data_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_en_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo;
	
	// wires for module twentynm_hssi_pipe_gen3
	wire	[7:0]	w_hssi_pipe_gen3_avmmreaddata;
	wire		w_hssi_pipe_gen3_blockselect;
	wire		w_hssi_pipe_gen3_gen3_clk_sel;
	wire		w_hssi_pipe_gen3_pcs_rst;
	wire		w_hssi_pipe_gen3_phystatus;
	wire	[17:0]	w_hssi_pipe_gen3_pma_current_coeff;
	wire	[2:0]	w_hssi_pipe_gen3_pma_current_rxpreset;
	wire		w_hssi_pipe_gen3_pma_tx_elec_idle;
	wire		w_hssi_pipe_gen3_pma_txdetectrx;
	wire		w_hssi_pipe_gen3_rev_lpbk_8gpcs_out;
	wire		w_hssi_pipe_gen3_rev_lpbk_int;
	wire	[3:0]	w_hssi_pipe_gen3_rx_blk_start;
	wire	[1:0]	w_hssi_pipe_gen3_rx_sync_hdr;
	wire	[63:0]	w_hssi_pipe_gen3_rxd_8gpcs_out;
	wire	[3:0]	w_hssi_pipe_gen3_rxdataskip;
	wire		w_hssi_pipe_gen3_rxelecidle;
	wire		w_hssi_pipe_gen3_rxpolarity_8gpcs_out;
	wire		w_hssi_pipe_gen3_rxpolarity_int;
	wire	[2:0]	w_hssi_pipe_gen3_rxstatus;
	wire		w_hssi_pipe_gen3_rxvalid;
	wire		w_hssi_pipe_gen3_shutdown_clk;
	wire	[19:0]	w_hssi_pipe_gen3_test_out;
	wire		w_hssi_pipe_gen3_tx_blk_start_int;
	wire	[1:0]	w_hssi_pipe_gen3_tx_sync_hdr_int;
	wire	[31:0]	w_hssi_pipe_gen3_txdata_int;
	wire	[3:0]	w_hssi_pipe_gen3_txdatak_int;
	wire		w_hssi_pipe_gen3_txdataskip_int;
	
	// wires for module twentynm_hssi_pipe_gen1_2
	wire	[7:0]	w_hssi_pipe_gen1_2_avmmreaddata;
	wire		w_hssi_pipe_gen1_2_blockselect;
	wire	[17:0]	w_hssi_pipe_gen1_2_current_coeff;
	wire		w_hssi_pipe_gen1_2_phystatus;
	wire		w_hssi_pipe_gen1_2_polarity_inversion_rx;
	wire		w_hssi_pipe_gen1_2_rev_loopbk;
	wire		w_hssi_pipe_gen1_2_rxelecidle;
	wire		w_hssi_pipe_gen1_2_rxelectricalidle_out;
	wire	[2:0]	w_hssi_pipe_gen1_2_rxstatus;
	wire		w_hssi_pipe_gen1_2_rxvalid;
	wire		w_hssi_pipe_gen1_2_tx_elec_idle_out;
	wire		w_hssi_pipe_gen1_2_txdetectrx;
	
	// wires for module twentynm_hssi_gen3_tx_pcs
	wire	[7:0]	w_hssi_gen3_tx_pcs_avmmreaddata;
	wire		w_hssi_gen3_tx_pcs_blockselect;
	wire	[31:0]	w_hssi_gen3_tx_pcs_data_out;
	wire	[35:0]	w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out;
	wire	[31:0]	w_hssi_gen3_tx_pcs_par_lpbk_out;
	wire	[19:0]	w_hssi_gen3_tx_pcs_tx_test_out;
	
	// wires for module twentynm_hssi_8g_rx_pcs
	wire	[3:0]	w_hssi_8g_rx_pcs_a1a2k1k2flag;
	wire	[7:0]	w_hssi_8g_rx_pcs_avmmreaddata;
	wire		w_hssi_8g_rx_pcs_blockselect;
	wire	[19:0]	w_hssi_8g_rx_pcs_chnl_test_bus_out;
	wire		w_hssi_8g_rx_pcs_clock_to_pld;
	wire	[63:0]	w_hssi_8g_rx_pcs_dataout;
	wire		w_hssi_8g_rx_pcs_dis_pc_byte;
	wire		w_hssi_8g_rx_pcs_eidle_detected;
	wire	[2:0]	w_hssi_8g_rx_pcs_eios_det_cdr_ctrl;
	wire		w_hssi_8g_rx_pcs_g3_rx_pma_rstn;
	wire		w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn;
	wire		w_hssi_8g_rx_pcs_gen2ngen1;
	wire	[19:0]	w_hssi_8g_rx_pcs_parallel_rev_loopback;
	wire		w_hssi_8g_rx_pcs_pc_fifo_empty;
	wire		w_hssi_8g_rx_pcs_pcfifofull;
	wire		w_hssi_8g_rx_pcs_phystatus;
	wire	[63:0]	w_hssi_8g_rx_pcs_pipe_data;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_up;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo;
	wire	[7:0]	w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rm_fifo_empty;
	wire		w_hssi_8g_rx_pcs_rm_fifo_full;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_blk_start;
	wire		w_hssi_8g_rx_pcs_rx_clk_out_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clkslip;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_data_valid;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rx_pipe_clk;
	wire		w_hssi_8g_rx_pcs_rx_pipe_soft_reset;
	wire		w_hssi_8g_rx_pcs_rx_pma_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_sync_hdr;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_up;
	wire	[2:0]	w_hssi_8g_rx_pcs_rxstatus;
	wire		w_hssi_8g_rx_pcs_rxvalid;
	wire		w_hssi_8g_rx_pcs_signal_detect_out;
	wire	[4:0]	w_hssi_8g_rx_pcs_word_align_boundary;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk;
	wire	[79:0]	w_hssi_8g_rx_pcs_wr_data_rx_phfifo;
	wire	[31:0]	w_hssi_8g_rx_pcs_wr_data_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo;
	
	// wires for module twentynm_hssi_fifo_rx_pcs
	wire	[7:0]	w_hssi_fifo_rx_pcs_avmmreaddata;
	wire		w_hssi_fifo_rx_pcs_blockselect;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out2_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out_8g_clock_comp;
	wire	[79:0]	w_hssi_fifo_rx_pcs_data_out_8g_phase_comp;
	wire	[39:0]	w_hssi_fifo_rx_pcs_data_out_gen3;
	
	// wires for module twentynm_hssi_common_pcs_pma_interface
	wire	[7:0]	w_hssi_common_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_common_pcs_pma_interface_blockselect;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in;
	wire	[19:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out;
	wire	[7:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus;
	wire		w_hssi_common_pcs_pma_interface_pma_adapt_start;
	wire		w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
	wire		w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
	wire	[17:0]	w_hssi_common_pcs_pma_interface_pma_current_coeff;
	wire	[2:0]	w_hssi_common_pcs_pma_interface_pma_current_rxpreset;
	wire		w_hssi_common_pcs_pma_interface_pma_early_eios;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_interface_select;
	wire		w_hssi_common_pcs_pma_interface_pma_ltd_b;
	wire		w_hssi_common_pcs_pma_interface_pma_ltr;
	wire		w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
	wire		w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_pcie_switch;
	wire		w_hssi_common_pcs_pma_interface_pma_ppm_lock;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_pma_reserved_out;
	wire		w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
	wire		w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up;
	
	
	generate
		
		//module instantiations
		
		// instantiating twentynm_hssi_10g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_rx_pcs
			twentynm_hssi_10g_rx_pcs #(
				.advanced_user_mode(hssi_10g_rx_pcs_advanced_user_mode),
				.align_del(hssi_10g_rx_pcs_align_del),
				.ber_bit_err_total_cnt(hssi_10g_rx_pcs_ber_bit_err_total_cnt),
				.ber_clken(hssi_10g_rx_pcs_ber_clken),
				.ber_xus_timer_window(hssi_10g_rx_pcs_ber_xus_timer_window),
				.bitslip_mode(hssi_10g_rx_pcs_bitslip_mode),
				.blksync_bitslip_type(hssi_10g_rx_pcs_blksync_bitslip_type),
				.blksync_bitslip_wait_cnt(hssi_10g_rx_pcs_blksync_bitslip_wait_cnt),
				.blksync_bitslip_wait_type(hssi_10g_rx_pcs_blksync_bitslip_wait_type),
				.blksync_bypass(hssi_10g_rx_pcs_blksync_bypass),
				.blksync_clken(hssi_10g_rx_pcs_blksync_clken),
				.blksync_enum_invalid_sh_cnt(hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt),
				.blksync_knum_sh_cnt_postlock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock),
				.blksync_knum_sh_cnt_prelock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock),
				.blksync_pipeln(hssi_10g_rx_pcs_blksync_pipeln),
				.clr_errblk_cnt_en(hssi_10g_rx_pcs_clr_errblk_cnt_en),
				.control_del(hssi_10g_rx_pcs_control_del),
				.crcchk_bypass(hssi_10g_rx_pcs_crcchk_bypass),
				.crcchk_clken(hssi_10g_rx_pcs_crcchk_clken),
				.crcchk_inv(hssi_10g_rx_pcs_crcchk_inv),
				.crcchk_pipeln(hssi_10g_rx_pcs_crcchk_pipeln),
				.crcflag_pipeln(hssi_10g_rx_pcs_crcflag_pipeln),
				.ctrl_bit_reverse(hssi_10g_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_10g_rx_pcs_data_bit_reverse),
				.dec64b66b_clken(hssi_10g_rx_pcs_dec64b66b_clken),
				.dec_64b66b_rxsm_bypass(hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass),
				.descrm_bypass(hssi_10g_rx_pcs_descrm_bypass),
				.descrm_clken(hssi_10g_rx_pcs_descrm_clken),
				.descrm_mode(hssi_10g_rx_pcs_descrm_mode),
				.descrm_pipeln(hssi_10g_rx_pcs_descrm_pipeln),
				.dft_clk_out_sel(hssi_10g_rx_pcs_dft_clk_out_sel),
				.dis_signal_ok(hssi_10g_rx_pcs_dis_signal_ok),
				.dispchk_bypass(hssi_10g_rx_pcs_dispchk_bypass),
				.empty_flag_type(hssi_10g_rx_pcs_empty_flag_type),
				.fast_path(hssi_10g_rx_pcs_fast_path),
				.fec_clken(hssi_10g_rx_pcs_fec_clken),
				.fec_enable(hssi_10g_rx_pcs_fec_enable),
				.fifo_double_read(hssi_10g_rx_pcs_fifo_double_read),
				.fifo_stop_rd(hssi_10g_rx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_rx_pcs_fifo_stop_wr),
				.force_align(hssi_10g_rx_pcs_force_align),
				.frmsync_bypass(hssi_10g_rx_pcs_frmsync_bypass),
				.frmsync_clken(hssi_10g_rx_pcs_frmsync_clken),
				.frmsync_enum_scrm(hssi_10g_rx_pcs_frmsync_enum_scrm),
				.frmsync_enum_sync(hssi_10g_rx_pcs_frmsync_enum_sync),
				.frmsync_flag_type(hssi_10g_rx_pcs_frmsync_flag_type),
				.frmsync_knum_sync(hssi_10g_rx_pcs_frmsync_knum_sync),
				.frmsync_mfrm_length(hssi_10g_rx_pcs_frmsync_mfrm_length),
				.frmsync_pipeln(hssi_10g_rx_pcs_frmsync_pipeln),
				.full_flag_type(hssi_10g_rx_pcs_full_flag_type),
				.gb_rx_idwidth(hssi_10g_rx_pcs_gb_rx_idwidth),
				.gb_rx_odwidth(hssi_10g_rx_pcs_gb_rx_odwidth),
				.gbexp_clken(hssi_10g_rx_pcs_gbexp_clken),
				.low_latency_en(hssi_10g_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_10g_rx_pcs_lpbk_mode),
				.master_clk_sel(hssi_10g_rx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_rx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_rx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_rx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_rx_pcs_pld_if_type),
				.prot_mode(hssi_10g_rx_pcs_prot_mode),
				.rand_clken(hssi_10g_rx_pcs_rand_clken),
				.rd_clk_sel(hssi_10g_rx_pcs_rd_clk_sel),
				.rdfifo_clken(hssi_10g_rx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_rx_pcs_reconfig_settings),
				.rx_fifo_write_ctrl(hssi_10g_rx_pcs_rx_fifo_write_ctrl),
				.rx_scrm_width(hssi_10g_rx_pcs_rx_scrm_width),
				.rx_sh_location(hssi_10g_rx_pcs_rx_sh_location),
				.rx_signal_ok_sel(hssi_10g_rx_pcs_rx_signal_ok_sel),
				.rx_sm_bypass(hssi_10g_rx_pcs_rx_sm_bypass),
				.rx_sm_hiber(hssi_10g_rx_pcs_rx_sm_hiber),
				.rx_sm_pipeln(hssi_10g_rx_pcs_rx_sm_pipeln),
				.rx_testbus_sel(hssi_10g_rx_pcs_rx_testbus_sel),
				.rx_true_b2b(hssi_10g_rx_pcs_rx_true_b2b),
				.rxfifo_empty(hssi_10g_rx_pcs_rxfifo_empty),
				.rxfifo_full(hssi_10g_rx_pcs_rxfifo_full),
				.rxfifo_mode(hssi_10g_rx_pcs_rxfifo_mode),
				.rxfifo_pempty(hssi_10g_rx_pcs_rxfifo_pempty),
				.rxfifo_pfull(hssi_10g_rx_pcs_rxfifo_pfull),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.stretch_num_stages(hssi_10g_rx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_rx_pcs_sup_mode),
				.test_mode(hssi_10g_rx_pcs_test_mode),
				.wrfifo_clken(hssi_10g_rx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_rx_pcs_blockselect),
				.rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.rx_control(w_hssi_10g_rx_pcs_rx_control),
				.rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.rx_data(w_hssi_10g_rx_pcs_rx_data),
				.rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.rx_diag_status(w_hssi_10g_rx_pcs_rx_diag_status),
				.rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.rx_fec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.rx_fifo_num(w_hssi_10g_rx_pcs_rx_fifo_num),
				.rx_fifo_rd_ptr(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr),
				.rx_fifo_rd_ptr2(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2),
				.rx_fifo_wr_clk(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.rx_fifo_wr_data(w_hssi_10g_rx_pcs_rx_fifo_wr_data),
				.rx_fifo_wr_en(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.rx_fifo_wr_ptr(w_hssi_10g_rx_pcs_rx_fifo_wr_ptr),
				.rx_fifo_wr_rst_n(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.rx_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_rx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_rx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.rx_control_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0]}),
				.rx_control_in_krfec({w_hssi_krfec_rx_pcs_rx_control_out[9], w_hssi_krfec_rx_pcs_rx_control_out[8], w_hssi_krfec_rx_pcs_rx_control_out[7], w_hssi_krfec_rx_pcs_rx_control_out[6], w_hssi_krfec_rx_pcs_rx_control_out[5], w_hssi_krfec_rx_pcs_rx_control_out[4], w_hssi_krfec_rx_pcs_rx_control_out[3], w_hssi_krfec_rx_pcs_rx_control_out[2], w_hssi_krfec_rx_pcs_rx_control_out[1], w_hssi_krfec_rx_pcs_rx_control_out[0]}),
				.rx_data_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0]}),
				.rx_data_in_krfec({w_hssi_krfec_rx_pcs_rx_data_out[63], w_hssi_krfec_rx_pcs_rx_data_out[62], w_hssi_krfec_rx_pcs_rx_data_out[61], w_hssi_krfec_rx_pcs_rx_data_out[60], w_hssi_krfec_rx_pcs_rx_data_out[59], w_hssi_krfec_rx_pcs_rx_data_out[58], w_hssi_krfec_rx_pcs_rx_data_out[57], w_hssi_krfec_rx_pcs_rx_data_out[56], w_hssi_krfec_rx_pcs_rx_data_out[55], w_hssi_krfec_rx_pcs_rx_data_out[54], w_hssi_krfec_rx_pcs_rx_data_out[53], w_hssi_krfec_rx_pcs_rx_data_out[52], w_hssi_krfec_rx_pcs_rx_data_out[51], w_hssi_krfec_rx_pcs_rx_data_out[50], w_hssi_krfec_rx_pcs_rx_data_out[49], w_hssi_krfec_rx_pcs_rx_data_out[48], w_hssi_krfec_rx_pcs_rx_data_out[47], w_hssi_krfec_rx_pcs_rx_data_out[46], w_hssi_krfec_rx_pcs_rx_data_out[45], w_hssi_krfec_rx_pcs_rx_data_out[44], w_hssi_krfec_rx_pcs_rx_data_out[43], w_hssi_krfec_rx_pcs_rx_data_out[42], w_hssi_krfec_rx_pcs_rx_data_out[41], w_hssi_krfec_rx_pcs_rx_data_out[40], w_hssi_krfec_rx_pcs_rx_data_out[39], w_hssi_krfec_rx_pcs_rx_data_out[38], w_hssi_krfec_rx_pcs_rx_data_out[37], w_hssi_krfec_rx_pcs_rx_data_out[36], w_hssi_krfec_rx_pcs_rx_data_out[35], w_hssi_krfec_rx_pcs_rx_data_out[34], w_hssi_krfec_rx_pcs_rx_data_out[33], w_hssi_krfec_rx_pcs_rx_data_out[32], w_hssi_krfec_rx_pcs_rx_data_out[31], w_hssi_krfec_rx_pcs_rx_data_out[30], w_hssi_krfec_rx_pcs_rx_data_out[29], w_hssi_krfec_rx_pcs_rx_data_out[28], w_hssi_krfec_rx_pcs_rx_data_out[27], w_hssi_krfec_rx_pcs_rx_data_out[26], w_hssi_krfec_rx_pcs_rx_data_out[25], w_hssi_krfec_rx_pcs_rx_data_out[24], w_hssi_krfec_rx_pcs_rx_data_out[23], w_hssi_krfec_rx_pcs_rx_data_out[22], w_hssi_krfec_rx_pcs_rx_data_out[21], w_hssi_krfec_rx_pcs_rx_data_out[20], w_hssi_krfec_rx_pcs_rx_data_out[19], w_hssi_krfec_rx_pcs_rx_data_out[18], w_hssi_krfec_rx_pcs_rx_data_out[17], w_hssi_krfec_rx_pcs_rx_data_out[16], w_hssi_krfec_rx_pcs_rx_data_out[15], w_hssi_krfec_rx_pcs_rx_data_out[14], w_hssi_krfec_rx_pcs_rx_data_out[13], w_hssi_krfec_rx_pcs_rx_data_out[12], w_hssi_krfec_rx_pcs_rx_data_out[11], w_hssi_krfec_rx_pcs_rx_data_out[10], w_hssi_krfec_rx_pcs_rx_data_out[9], w_hssi_krfec_rx_pcs_rx_data_out[8], w_hssi_krfec_rx_pcs_rx_data_out[7], w_hssi_krfec_rx_pcs_rx_data_out[6], w_hssi_krfec_rx_pcs_rx_data_out[5], w_hssi_krfec_rx_pcs_rx_data_out[4], w_hssi_krfec_rx_pcs_rx_data_out[3], w_hssi_krfec_rx_pcs_rx_data_out[2], w_hssi_krfec_rx_pcs_rx_data_out[1], w_hssi_krfec_rx_pcs_rx_data_out[0]}),
				.rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.rx_data_valid_in_krfec(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_10g[73], w_hssi_fifo_rx_pcs_data_out_10g[72], w_hssi_fifo_rx_pcs_data_out_10g[71], w_hssi_fifo_rx_pcs_data_out_10g[70], w_hssi_fifo_rx_pcs_data_out_10g[69], w_hssi_fifo_rx_pcs_data_out_10g[68], w_hssi_fifo_rx_pcs_data_out_10g[67], w_hssi_fifo_rx_pcs_data_out_10g[66], w_hssi_fifo_rx_pcs_data_out_10g[65], w_hssi_fifo_rx_pcs_data_out_10g[64], w_hssi_fifo_rx_pcs_data_out_10g[63], w_hssi_fifo_rx_pcs_data_out_10g[62], w_hssi_fifo_rx_pcs_data_out_10g[61], w_hssi_fifo_rx_pcs_data_out_10g[60], w_hssi_fifo_rx_pcs_data_out_10g[59], w_hssi_fifo_rx_pcs_data_out_10g[58], w_hssi_fifo_rx_pcs_data_out_10g[57], w_hssi_fifo_rx_pcs_data_out_10g[56], w_hssi_fifo_rx_pcs_data_out_10g[55], w_hssi_fifo_rx_pcs_data_out_10g[54], w_hssi_fifo_rx_pcs_data_out_10g[53], w_hssi_fifo_rx_pcs_data_out_10g[52], w_hssi_fifo_rx_pcs_data_out_10g[51], w_hssi_fifo_rx_pcs_data_out_10g[50], w_hssi_fifo_rx_pcs_data_out_10g[49], w_hssi_fifo_rx_pcs_data_out_10g[48], w_hssi_fifo_rx_pcs_data_out_10g[47], w_hssi_fifo_rx_pcs_data_out_10g[46], w_hssi_fifo_rx_pcs_data_out_10g[45], w_hssi_fifo_rx_pcs_data_out_10g[44], w_hssi_fifo_rx_pcs_data_out_10g[43], w_hssi_fifo_rx_pcs_data_out_10g[42], w_hssi_fifo_rx_pcs_data_out_10g[41], w_hssi_fifo_rx_pcs_data_out_10g[40], w_hssi_fifo_rx_pcs_data_out_10g[39], w_hssi_fifo_rx_pcs_data_out_10g[38], w_hssi_fifo_rx_pcs_data_out_10g[37], w_hssi_fifo_rx_pcs_data_out_10g[36], w_hssi_fifo_rx_pcs_data_out_10g[35], w_hssi_fifo_rx_pcs_data_out_10g[34], w_hssi_fifo_rx_pcs_data_out_10g[33], w_hssi_fifo_rx_pcs_data_out_10g[32], w_hssi_fifo_rx_pcs_data_out_10g[31], w_hssi_fifo_rx_pcs_data_out_10g[30], w_hssi_fifo_rx_pcs_data_out_10g[29], w_hssi_fifo_rx_pcs_data_out_10g[28], w_hssi_fifo_rx_pcs_data_out_10g[27], w_hssi_fifo_rx_pcs_data_out_10g[26], w_hssi_fifo_rx_pcs_data_out_10g[25], w_hssi_fifo_rx_pcs_data_out_10g[24], w_hssi_fifo_rx_pcs_data_out_10g[23], w_hssi_fifo_rx_pcs_data_out_10g[22], w_hssi_fifo_rx_pcs_data_out_10g[21], w_hssi_fifo_rx_pcs_data_out_10g[20], w_hssi_fifo_rx_pcs_data_out_10g[19], w_hssi_fifo_rx_pcs_data_out_10g[18], w_hssi_fifo_rx_pcs_data_out_10g[17], w_hssi_fifo_rx_pcs_data_out_10g[16], w_hssi_fifo_rx_pcs_data_out_10g[15], w_hssi_fifo_rx_pcs_data_out_10g[14], w_hssi_fifo_rx_pcs_data_out_10g[13], w_hssi_fifo_rx_pcs_data_out_10g[12], w_hssi_fifo_rx_pcs_data_out_10g[11], w_hssi_fifo_rx_pcs_data_out_10g[10], w_hssi_fifo_rx_pcs_data_out_10g[9], w_hssi_fifo_rx_pcs_data_out_10g[8], w_hssi_fifo_rx_pcs_data_out_10g[7], w_hssi_fifo_rx_pcs_data_out_10g[6], w_hssi_fifo_rx_pcs_data_out_10g[5], w_hssi_fifo_rx_pcs_data_out_10g[4], w_hssi_fifo_rx_pcs_data_out_10g[3], w_hssi_fifo_rx_pcs_data_out_10g[2], w_hssi_fifo_rx_pcs_data_out_10g[1], w_hssi_fifo_rx_pcs_data_out_10g[0]}),
				.rx_fifo_rd_data_dw({w_hssi_fifo_rx_pcs_data_out2_10g[73], w_hssi_fifo_rx_pcs_data_out2_10g[72], w_hssi_fifo_rx_pcs_data_out2_10g[71], w_hssi_fifo_rx_pcs_data_out2_10g[70], w_hssi_fifo_rx_pcs_data_out2_10g[69], w_hssi_fifo_rx_pcs_data_out2_10g[68], w_hssi_fifo_rx_pcs_data_out2_10g[67], w_hssi_fifo_rx_pcs_data_out2_10g[66], w_hssi_fifo_rx_pcs_data_out2_10g[65], w_hssi_fifo_rx_pcs_data_out2_10g[64], w_hssi_fifo_rx_pcs_data_out2_10g[63], w_hssi_fifo_rx_pcs_data_out2_10g[62], w_hssi_fifo_rx_pcs_data_out2_10g[61], w_hssi_fifo_rx_pcs_data_out2_10g[60], w_hssi_fifo_rx_pcs_data_out2_10g[59], w_hssi_fifo_rx_pcs_data_out2_10g[58], w_hssi_fifo_rx_pcs_data_out2_10g[57], w_hssi_fifo_rx_pcs_data_out2_10g[56], w_hssi_fifo_rx_pcs_data_out2_10g[55], w_hssi_fifo_rx_pcs_data_out2_10g[54], w_hssi_fifo_rx_pcs_data_out2_10g[53], w_hssi_fifo_rx_pcs_data_out2_10g[52], w_hssi_fifo_rx_pcs_data_out2_10g[51], w_hssi_fifo_rx_pcs_data_out2_10g[50], w_hssi_fifo_rx_pcs_data_out2_10g[49], w_hssi_fifo_rx_pcs_data_out2_10g[48], w_hssi_fifo_rx_pcs_data_out2_10g[47], w_hssi_fifo_rx_pcs_data_out2_10g[46], w_hssi_fifo_rx_pcs_data_out2_10g[45], w_hssi_fifo_rx_pcs_data_out2_10g[44], w_hssi_fifo_rx_pcs_data_out2_10g[43], w_hssi_fifo_rx_pcs_data_out2_10g[42], w_hssi_fifo_rx_pcs_data_out2_10g[41], w_hssi_fifo_rx_pcs_data_out2_10g[40], w_hssi_fifo_rx_pcs_data_out2_10g[39], w_hssi_fifo_rx_pcs_data_out2_10g[38], w_hssi_fifo_rx_pcs_data_out2_10g[37], w_hssi_fifo_rx_pcs_data_out2_10g[36], w_hssi_fifo_rx_pcs_data_out2_10g[35], w_hssi_fifo_rx_pcs_data_out2_10g[34], w_hssi_fifo_rx_pcs_data_out2_10g[33], w_hssi_fifo_rx_pcs_data_out2_10g[32], w_hssi_fifo_rx_pcs_data_out2_10g[31], w_hssi_fifo_rx_pcs_data_out2_10g[30], w_hssi_fifo_rx_pcs_data_out2_10g[29], w_hssi_fifo_rx_pcs_data_out2_10g[28], w_hssi_fifo_rx_pcs_data_out2_10g[27], w_hssi_fifo_rx_pcs_data_out2_10g[26], w_hssi_fifo_rx_pcs_data_out2_10g[25], w_hssi_fifo_rx_pcs_data_out2_10g[24], w_hssi_fifo_rx_pcs_data_out2_10g[23], w_hssi_fifo_rx_pcs_data_out2_10g[22], w_hssi_fifo_rx_pcs_data_out2_10g[21], w_hssi_fifo_rx_pcs_data_out2_10g[20], w_hssi_fifo_rx_pcs_data_out2_10g[19], w_hssi_fifo_rx_pcs_data_out2_10g[18], w_hssi_fifo_rx_pcs_data_out2_10g[17], w_hssi_fifo_rx_pcs_data_out2_10g[16], w_hssi_fifo_rx_pcs_data_out2_10g[15], w_hssi_fifo_rx_pcs_data_out2_10g[14], w_hssi_fifo_rx_pcs_data_out2_10g[13], w_hssi_fifo_rx_pcs_data_out2_10g[12], w_hssi_fifo_rx_pcs_data_out2_10g[11], w_hssi_fifo_rx_pcs_data_out2_10g[10], w_hssi_fifo_rx_pcs_data_out2_10g[9], w_hssi_fifo_rx_pcs_data_out2_10g[8], w_hssi_fifo_rx_pcs_data_out2_10g[7], w_hssi_fifo_rx_pcs_data_out2_10g[6], w_hssi_fifo_rx_pcs_data_out2_10g[5], w_hssi_fifo_rx_pcs_data_out2_10g[4], w_hssi_fifo_rx_pcs_data_out2_10g[3], w_hssi_fifo_rx_pcs_data_out2_10g[2], w_hssi_fifo_rx_pcs_data_out2_10g[1], w_hssi_fifo_rx_pcs_data_out2_10g[0]}),
				.rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.rx_pma_data({w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0]}),
				.rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.signal_ok_krfec(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_10g_reg(),
				.pld_10g_krfec_rx_blk_lock_10g_txclk_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_txclk_reg(),
				.pld_10g_krfec_rx_frame_10g_reg(),
				.pld_10g_krfec_rx_frame_10g_txclk_reg(),
				.pld_10g_krfec_rx_pld_rst_n_fifo(),
				.pld_10g_krfec_rx_pld_rst_n_reg(),
				.pld_10g_krfec_rx_pld_rst_n_txclk_reg(),
				.pld_10g_rx_align_clr_fifo(),
				.pld_10g_rx_align_clr_reg(),
				.pld_10g_rx_align_clr_txclk_reg(),
				.pld_10g_rx_align_val_fifo(),
				.pld_10g_rx_align_val_reg(),
				.pld_10g_rx_align_val_txclk_reg(),
				.pld_10g_rx_clr_ber_count_reg(),
				.pld_10g_rx_clr_ber_count_txclk_reg(),
				.pld_10g_rx_crc32_err_reg(),
				.pld_10g_rx_crc32_err_txclk_reg(),
				.pld_10g_rx_data_valid_10g_reg(),
				.pld_10g_rx_data_valid_fifo(),
				.pld_10g_rx_data_valid_pcsdirect_reg(),
				.pld_10g_rx_data_valid_txclk_reg(),
				.pld_10g_rx_empty_fifo(),
				.pld_10g_rx_fifo_del_reg(),
				.pld_10g_rx_fifo_del_txclk_reg(),
				.pld_10g_rx_fifo_insert_fifo(),
				.pld_10g_rx_fifo_num_reg(),
				.pld_10g_rx_fifo_num_txclk_reg(),
				.pld_10g_rx_frame_lock_reg(),
				.pld_10g_rx_frame_lock_txclk_reg(),
				.pld_10g_rx_hi_ber_reg(),
				.pld_10g_rx_hi_ber_txclk_reg(),
				.pld_10g_rx_oflw_err_reg(),
				.pld_10g_rx_oflw_err_txclk_reg(),
				.pld_10g_rx_pempty_fifo(),
				.pld_10g_rx_pfull_reg(),
				.pld_10g_rx_pfull_txclk_reg(),
				.pld_10g_rx_rd_en_fifo(),
				.pld_pcs_rx_clk_out_10g_txclk_wire(),
				.pld_pcs_rx_clk_out_10g_wire(),
				.pld_rx_control_10g_reg(),
				.pld_rx_control_10g_txclk_reg(),
				.pld_rx_data_10g_reg(),
				.pld_rx_data_10g_txclk_reg(),
				.pld_rx_prbs_err_10g_txclk_reg(),
				.pld_rx_prbs_err_clr_10g_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_10g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_align_val = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_blk_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_control[19:0] = 20'b0;
				assign w_hssi_10g_rx_pcs_rx_crc32_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_data[127:0] = 128'b0;
				assign w_hssi_10g_rx_pcs_rx_data_valid = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_dft_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_diag_status[1:0] = 2'b0;
				assign w_hssi_10g_rx_pcs_rx_empty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fec_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_del = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_insert = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_data[73:0] = 74'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_frame_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_hi_ber = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_oflw_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pempty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pfull = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_random_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_rx_frame = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_10g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_tx_pcs
			twentynm_hssi_10g_tx_pcs #(
				.advanced_user_mode(hssi_10g_tx_pcs_advanced_user_mode),
				.bitslip_en(hssi_10g_tx_pcs_bitslip_en),
				.bonding_dft_en(hssi_10g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_10g_tx_pcs_bonding_dft_val),
				.comp_cnt(hssi_10g_tx_pcs_comp_cnt),
				.compin_sel(hssi_10g_tx_pcs_compin_sel),
				.crcgen_bypass(hssi_10g_tx_pcs_crcgen_bypass),
				.crcgen_clken(hssi_10g_tx_pcs_crcgen_clken),
				.crcgen_err(hssi_10g_tx_pcs_crcgen_err),
				.crcgen_inv(hssi_10g_tx_pcs_crcgen_inv),
				.ctrl_bit_reverse(hssi_10g_tx_pcs_ctrl_bit_reverse),
				.ctrl_plane_bonding(hssi_10g_tx_pcs_ctrl_plane_bonding),
				.data_bit_reverse(hssi_10g_tx_pcs_data_bit_reverse),
				.dft_clk_out_sel(hssi_10g_tx_pcs_dft_clk_out_sel),
				.dispgen_bypass(hssi_10g_tx_pcs_dispgen_bypass),
				.dispgen_clken(hssi_10g_tx_pcs_dispgen_clken),
				.dispgen_err(hssi_10g_tx_pcs_dispgen_err),
				.dispgen_pipeln(hssi_10g_tx_pcs_dispgen_pipeln),
				.distdwn_bypass_pipeln(hssi_10g_tx_pcs_distdwn_bypass_pipeln),
				.distdwn_master(hssi_10g_tx_pcs_distdwn_master),
				.distup_bypass_pipeln(hssi_10g_tx_pcs_distup_bypass_pipeln),
				.distup_master(hssi_10g_tx_pcs_distup_master),
				.dv_bond(hssi_10g_tx_pcs_dv_bond),
				.empty_flag_type(hssi_10g_tx_pcs_empty_flag_type),
				.enc64b66b_txsm_clken(hssi_10g_tx_pcs_enc64b66b_txsm_clken),
				.enc_64b66b_txsm_bypass(hssi_10g_tx_pcs_enc_64b66b_txsm_bypass),
				.fastpath(hssi_10g_tx_pcs_fastpath),
				.fec_clken(hssi_10g_tx_pcs_fec_clken),
				.fec_enable(hssi_10g_tx_pcs_fec_enable),
				.fifo_double_write(hssi_10g_tx_pcs_fifo_double_write),
				.fifo_reg_fast(hssi_10g_tx_pcs_fifo_reg_fast),
				.fifo_stop_rd(hssi_10g_tx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_tx_pcs_fifo_stop_wr),
				.frmgen_burst(hssi_10g_tx_pcs_frmgen_burst),
				.frmgen_bypass(hssi_10g_tx_pcs_frmgen_bypass),
				.frmgen_clken(hssi_10g_tx_pcs_frmgen_clken),
				.frmgen_mfrm_length(hssi_10g_tx_pcs_frmgen_mfrm_length),
				.frmgen_pipeln(hssi_10g_tx_pcs_frmgen_pipeln),
				.frmgen_pyld_ins(hssi_10g_tx_pcs_frmgen_pyld_ins),
				.frmgen_wordslip(hssi_10g_tx_pcs_frmgen_wordslip),
				.full_flag_type(hssi_10g_tx_pcs_full_flag_type),
				.gb_pipeln_bypass(hssi_10g_tx_pcs_gb_pipeln_bypass),
				.gb_tx_idwidth(hssi_10g_tx_pcs_gb_tx_idwidth),
				.gb_tx_odwidth(hssi_10g_tx_pcs_gb_tx_odwidth),
				.gbred_clken(hssi_10g_tx_pcs_gbred_clken),
				.indv(hssi_10g_tx_pcs_indv),
				.low_latency_en(hssi_10g_tx_pcs_low_latency_en),
				.master_clk_sel(hssi_10g_tx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_tx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_tx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_tx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_tx_pcs_pld_if_type),
				.prot_mode(hssi_10g_tx_pcs_prot_mode),
				.pseudo_random(hssi_10g_tx_pcs_pseudo_random),
				.pseudo_seed_a(hssi_10g_tx_pcs_pseudo_seed_a),
				.pseudo_seed_b(hssi_10g_tx_pcs_pseudo_seed_b),
				.random_disp(hssi_10g_tx_pcs_random_disp),
				.rdfifo_clken(hssi_10g_tx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_tx_pcs_reconfig_settings),
				.scrm_bypass(hssi_10g_tx_pcs_scrm_bypass),
				.scrm_clken(hssi_10g_tx_pcs_scrm_clken),
				.scrm_mode(hssi_10g_tx_pcs_scrm_mode),
				.scrm_pipeln(hssi_10g_tx_pcs_scrm_pipeln),
				.sh_err(hssi_10g_tx_pcs_sh_err),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sop_mark(hssi_10g_tx_pcs_sop_mark),
				.stretch_num_stages(hssi_10g_tx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_tx_pcs_sup_mode),
				.test_mode(hssi_10g_tx_pcs_test_mode),
				.tx_scrm_err(hssi_10g_tx_pcs_tx_scrm_err),
				.tx_scrm_width(hssi_10g_tx_pcs_tx_scrm_width),
				.tx_sh_location(hssi_10g_tx_pcs_tx_sh_location),
				.tx_sm_bypass(hssi_10g_tx_pcs_tx_sm_bypass),
				.tx_sm_pipeln(hssi_10g_tx_pcs_tx_sm_pipeln),
				.tx_testbus_sel(hssi_10g_tx_pcs_tx_testbus_sel),
				.txfifo_empty(hssi_10g_tx_pcs_txfifo_empty),
				.txfifo_full(hssi_10g_tx_pcs_txfifo_full),
				.txfifo_mode(hssi_10g_tx_pcs_txfifo_mode),
				.txfifo_pempty(hssi_10g_tx_pcs_txfifo_pempty),
				.txfifo_pfull(hssi_10g_tx_pcs_txfifo_pfull),
				.wr_clk_sel(hssi_10g_tx_pcs_wr_clk_sel),
				.wrfifo_clken(hssi_10g_tx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_tx_pcs_blockselect),
				.distdwn_out_dv(w_hssi_10g_tx_pcs_distdwn_out_dv),
				.distdwn_out_rden(w_hssi_10g_tx_pcs_distdwn_out_rden),
				.distdwn_out_wren(w_hssi_10g_tx_pcs_distdwn_out_wren),
				.distup_out_dv(w_hssi_10g_tx_pcs_distup_out_dv),
				.distup_out_rden(w_hssi_10g_tx_pcs_distup_out_rden),
				.distup_out_wren(w_hssi_10g_tx_pcs_distup_out_wren),
				.tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pma_if(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.tx_control_out_krfec(w_hssi_10g_tx_pcs_tx_control_out_krfec),
				.tx_data_out_krfec(w_hssi_10g_tx_pcs_tx_data_out_krfec),
				.tx_data_valid_out_krfec(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.tx_fec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_fifo_num(w_hssi_10g_tx_pcs_tx_fifo_num),
				.tx_fifo_rd_ptr(w_hssi_10g_tx_pcs_tx_fifo_rd_ptr),
				.tx_fifo_wr_clk(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.tx_fifo_wr_data(w_hssi_10g_tx_pcs_tx_fifo_wr_data),
				.tx_fifo_wr_data_dw(w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw),
				.tx_fifo_wr_en(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.tx_fifo_wr_ptr(w_hssi_10g_tx_pcs_tx_fifo_wr_ptr),
				.tx_fifo_wr_rst_n(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.tx_full(w_hssi_10g_tx_pcs_tx_full),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				.tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.tx_pma_data(w_hssi_10g_tx_pcs_tx_pma_data),
				.tx_pma_gating_val(w_hssi_10g_tx_pcs_tx_pma_gating_val),
				.tx_test_data(w_hssi_10g_tx_pcs_tx_test_data),
				.tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.distdwn_in_dv(in_bond_pcs10g_in_bot[2]),
				.distdwn_in_rden(in_bond_pcs10g_in_bot[4]),
				.distdwn_in_wren(in_bond_pcs10g_in_bot[3]),
				.distup_in_dv(in_bond_pcs10g_in_top[2]),
				.distup_in_rden(in_bond_pcs10g_in_top[4]),
				.distup_in_wren(in_bond_pcs10g_in_top[3]),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_tx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_tx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.tx_bitslip({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0]}),
				.tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.tx_control({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0]}),
				.tx_control_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0]}),
				.tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0]}),
				.tx_data_in_krfec({w_hssi_krfec_tx_pcs_tx_data_out[63], w_hssi_krfec_tx_pcs_tx_data_out[62], w_hssi_krfec_tx_pcs_tx_data_out[61], w_hssi_krfec_tx_pcs_tx_data_out[60], w_hssi_krfec_tx_pcs_tx_data_out[59], w_hssi_krfec_tx_pcs_tx_data_out[58], w_hssi_krfec_tx_pcs_tx_data_out[57], w_hssi_krfec_tx_pcs_tx_data_out[56], w_hssi_krfec_tx_pcs_tx_data_out[55], w_hssi_krfec_tx_pcs_tx_data_out[54], w_hssi_krfec_tx_pcs_tx_data_out[53], w_hssi_krfec_tx_pcs_tx_data_out[52], w_hssi_krfec_tx_pcs_tx_data_out[51], w_hssi_krfec_tx_pcs_tx_data_out[50], w_hssi_krfec_tx_pcs_tx_data_out[49], w_hssi_krfec_tx_pcs_tx_data_out[48], w_hssi_krfec_tx_pcs_tx_data_out[47], w_hssi_krfec_tx_pcs_tx_data_out[46], w_hssi_krfec_tx_pcs_tx_data_out[45], w_hssi_krfec_tx_pcs_tx_data_out[44], w_hssi_krfec_tx_pcs_tx_data_out[43], w_hssi_krfec_tx_pcs_tx_data_out[42], w_hssi_krfec_tx_pcs_tx_data_out[41], w_hssi_krfec_tx_pcs_tx_data_out[40], w_hssi_krfec_tx_pcs_tx_data_out[39], w_hssi_krfec_tx_pcs_tx_data_out[38], w_hssi_krfec_tx_pcs_tx_data_out[37], w_hssi_krfec_tx_pcs_tx_data_out[36], w_hssi_krfec_tx_pcs_tx_data_out[35], w_hssi_krfec_tx_pcs_tx_data_out[34], w_hssi_krfec_tx_pcs_tx_data_out[33], w_hssi_krfec_tx_pcs_tx_data_out[32], w_hssi_krfec_tx_pcs_tx_data_out[31], w_hssi_krfec_tx_pcs_tx_data_out[30], w_hssi_krfec_tx_pcs_tx_data_out[29], w_hssi_krfec_tx_pcs_tx_data_out[28], w_hssi_krfec_tx_pcs_tx_data_out[27], w_hssi_krfec_tx_pcs_tx_data_out[26], w_hssi_krfec_tx_pcs_tx_data_out[25], w_hssi_krfec_tx_pcs_tx_data_out[24], w_hssi_krfec_tx_pcs_tx_data_out[23], w_hssi_krfec_tx_pcs_tx_data_out[22], w_hssi_krfec_tx_pcs_tx_data_out[21], w_hssi_krfec_tx_pcs_tx_data_out[20], w_hssi_krfec_tx_pcs_tx_data_out[19], w_hssi_krfec_tx_pcs_tx_data_out[18], w_hssi_krfec_tx_pcs_tx_data_out[17], w_hssi_krfec_tx_pcs_tx_data_out[16], w_hssi_krfec_tx_pcs_tx_data_out[15], w_hssi_krfec_tx_pcs_tx_data_out[14], w_hssi_krfec_tx_pcs_tx_data_out[13], w_hssi_krfec_tx_pcs_tx_data_out[12], w_hssi_krfec_tx_pcs_tx_data_out[11], w_hssi_krfec_tx_pcs_tx_data_out[10], w_hssi_krfec_tx_pcs_tx_data_out[9], w_hssi_krfec_tx_pcs_tx_data_out[8], w_hssi_krfec_tx_pcs_tx_data_out[7], w_hssi_krfec_tx_pcs_tx_data_out[6], w_hssi_krfec_tx_pcs_tx_data_out[5], w_hssi_krfec_tx_pcs_tx_data_out[4], w_hssi_krfec_tx_pcs_tx_data_out[3], w_hssi_krfec_tx_pcs_tx_data_out[2], w_hssi_krfec_tx_pcs_tx_data_out[1], w_hssi_krfec_tx_pcs_tx_data_out[0]}),
				.tx_data_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0]}),
				.tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.tx_diag_status({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0]}),
				.tx_fifo_rd_data({w_hssi_fifo_tx_pcs_data_out_10g[72], w_hssi_fifo_tx_pcs_data_out_10g[71], w_hssi_fifo_tx_pcs_data_out_10g[70], w_hssi_fifo_tx_pcs_data_out_10g[69], w_hssi_fifo_tx_pcs_data_out_10g[68], w_hssi_fifo_tx_pcs_data_out_10g[67], w_hssi_fifo_tx_pcs_data_out_10g[66], w_hssi_fifo_tx_pcs_data_out_10g[65], w_hssi_fifo_tx_pcs_data_out_10g[64], w_hssi_fifo_tx_pcs_data_out_10g[63], w_hssi_fifo_tx_pcs_data_out_10g[62], w_hssi_fifo_tx_pcs_data_out_10g[61], w_hssi_fifo_tx_pcs_data_out_10g[60], w_hssi_fifo_tx_pcs_data_out_10g[59], w_hssi_fifo_tx_pcs_data_out_10g[58], w_hssi_fifo_tx_pcs_data_out_10g[57], w_hssi_fifo_tx_pcs_data_out_10g[56], w_hssi_fifo_tx_pcs_data_out_10g[55], w_hssi_fifo_tx_pcs_data_out_10g[54], w_hssi_fifo_tx_pcs_data_out_10g[53], w_hssi_fifo_tx_pcs_data_out_10g[52], w_hssi_fifo_tx_pcs_data_out_10g[51], w_hssi_fifo_tx_pcs_data_out_10g[50], w_hssi_fifo_tx_pcs_data_out_10g[49], w_hssi_fifo_tx_pcs_data_out_10g[48], w_hssi_fifo_tx_pcs_data_out_10g[47], w_hssi_fifo_tx_pcs_data_out_10g[46], w_hssi_fifo_tx_pcs_data_out_10g[45], w_hssi_fifo_tx_pcs_data_out_10g[44], w_hssi_fifo_tx_pcs_data_out_10g[43], w_hssi_fifo_tx_pcs_data_out_10g[42], w_hssi_fifo_tx_pcs_data_out_10g[41], w_hssi_fifo_tx_pcs_data_out_10g[40], w_hssi_fifo_tx_pcs_data_out_10g[39], w_hssi_fifo_tx_pcs_data_out_10g[38], w_hssi_fifo_tx_pcs_data_out_10g[37], w_hssi_fifo_tx_pcs_data_out_10g[36], w_hssi_fifo_tx_pcs_data_out_10g[35], w_hssi_fifo_tx_pcs_data_out_10g[34], w_hssi_fifo_tx_pcs_data_out_10g[33], w_hssi_fifo_tx_pcs_data_out_10g[32], w_hssi_fifo_tx_pcs_data_out_10g[31], w_hssi_fifo_tx_pcs_data_out_10g[30], w_hssi_fifo_tx_pcs_data_out_10g[29], w_hssi_fifo_tx_pcs_data_out_10g[28], w_hssi_fifo_tx_pcs_data_out_10g[27], w_hssi_fifo_tx_pcs_data_out_10g[26], w_hssi_fifo_tx_pcs_data_out_10g[25], w_hssi_fifo_tx_pcs_data_out_10g[24], w_hssi_fifo_tx_pcs_data_out_10g[23], w_hssi_fifo_tx_pcs_data_out_10g[22], w_hssi_fifo_tx_pcs_data_out_10g[21], w_hssi_fifo_tx_pcs_data_out_10g[20], w_hssi_fifo_tx_pcs_data_out_10g[19], w_hssi_fifo_tx_pcs_data_out_10g[18], w_hssi_fifo_tx_pcs_data_out_10g[17], w_hssi_fifo_tx_pcs_data_out_10g[16], w_hssi_fifo_tx_pcs_data_out_10g[15], w_hssi_fifo_tx_pcs_data_out_10g[14], w_hssi_fifo_tx_pcs_data_out_10g[13], w_hssi_fifo_tx_pcs_data_out_10g[12], w_hssi_fifo_tx_pcs_data_out_10g[11], w_hssi_fifo_tx_pcs_data_out_10g[10], w_hssi_fifo_tx_pcs_data_out_10g[9], w_hssi_fifo_tx_pcs_data_out_10g[8], w_hssi_fifo_tx_pcs_data_out_10g[7], w_hssi_fifo_tx_pcs_data_out_10g[6], w_hssi_fifo_tx_pcs_data_out_10g[5], w_hssi_fifo_tx_pcs_data_out_10g[4], w_hssi_fifo_tx_pcs_data_out_10g[3], w_hssi_fifo_tx_pcs_data_out_10g[2], w_hssi_fifo_tx_pcs_data_out_10g[1], w_hssi_fifo_tx_pcs_data_out_10g[0]}),
				.tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_10g_reg(),
				.pld_10g_krfec_tx_pld_rst_n_fifo(),
				.pld_10g_krfec_tx_pld_rst_n_reg(),
				.pld_10g_tx_bitslip_reg(),
				.pld_10g_tx_burst_en_exe_reg(),
				.pld_10g_tx_data_valid_10g_reg(),
				.pld_10g_tx_data_valid_fifo(),
				.pld_10g_tx_data_valid_reg(),
				.pld_10g_tx_diag_status_reg(),
				.pld_10g_tx_empty_reg(),
				.pld_10g_tx_fifo_num_reg(),
				.pld_10g_tx_full_fifo(),
				.pld_10g_tx_full_reg(),
				.pld_10g_tx_pempty_reg(),
				.pld_10g_tx_pfull_fifo(),
				.pld_10g_tx_wordslip_exe_reg(),
				.pld_10g_tx_wordslip_reg(),
				.pld_pcs_tx_clk_out_10g_wire(),
				.pld_tx_burst_en_reg(),
				.pld_tx_control_lo_10g_reg(),
				.pld_tx_data_10g_fifo(),
				.pld_tx_data_lo_10g_reg()
			);
		end // if generate
		else begin
				assign w_hssi_10g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_burst_en_exe = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pma_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_control_out_krfec[8:0] = 9'b0;
				assign w_hssi_10g_tx_pcs_tx_data_out_krfec[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_data_valid_out_krfec = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_dft_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_empty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fec_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_full = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_pempty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pfull = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_gating_val[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_test_data[19:0] = 20'b0;
				assign w_hssi_10g_tx_pcs_tx_wordslip_exe = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_rx_pcs
			twentynm_hssi_8g_rx_pcs #(
				.auto_error_replacement(hssi_8g_rx_pcs_auto_error_replacement),
				.auto_speed_nego(hssi_8g_rx_pcs_auto_speed_nego),
				.bit_reversal(hssi_8g_rx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_rx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_rx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_rx_pcs_bypass_pipeline_reg),
				.byte_deserializer(hssi_8g_rx_pcs_byte_deserializer),
				.cdr_ctrl_rxvalid_mask(hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask),
				.clkcmp_pattern_n(hssi_8g_rx_pcs_clkcmp_pattern_n),
				.clkcmp_pattern_p(hssi_8g_rx_pcs_clkcmp_pattern_p),
				.clock_gate_bds_dec_asn(hssi_8g_rx_pcs_clock_gate_bds_dec_asn),
				.clock_gate_cdr_eidle(hssi_8g_rx_pcs_clock_gate_cdr_eidle),
				.clock_gate_dw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk),
				.clock_gate_dw_rm_rd(hssi_8g_rx_pcs_clock_gate_dw_rm_rd),
				.clock_gate_dw_rm_wr(hssi_8g_rx_pcs_clock_gate_dw_rm_wr),
				.clock_gate_dw_wa(hssi_8g_rx_pcs_clock_gate_dw_wa),
				.clock_gate_pc_rdclk(hssi_8g_rx_pcs_clock_gate_pc_rdclk),
				.clock_gate_sw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk),
				.clock_gate_sw_rm_rd(hssi_8g_rx_pcs_clock_gate_sw_rm_rd),
				.clock_gate_sw_rm_wr(hssi_8g_rx_pcs_clock_gate_sw_rm_wr),
				.clock_gate_sw_wa(hssi_8g_rx_pcs_clock_gate_sw_wa),
				.clock_observation_in_pld_core(hssi_8g_rx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_rx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_rx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_rx_pcs_ctrl_plane_bonding_distribution),
				.eidle_entry_eios(hssi_8g_rx_pcs_eidle_entry_eios),
				.eidle_entry_iei(hssi_8g_rx_pcs_eidle_entry_iei),
				.eidle_entry_sd(hssi_8g_rx_pcs_eidle_entry_sd),
				.eightb_tenb_decoder(hssi_8g_rx_pcs_eightb_tenb_decoder),
				.err_flags_sel(hssi_8g_rx_pcs_err_flags_sel),
				.fixed_pat_det(hssi_8g_rx_pcs_fixed_pat_det),
				.fixed_pat_num(hssi_8g_rx_pcs_fixed_pat_num),
				.force_signal_detect(hssi_8g_rx_pcs_force_signal_detect),
				.gen3_clk_en(hssi_8g_rx_pcs_gen3_clk_en),
				.gen3_rx_clk_sel(hssi_8g_rx_pcs_gen3_rx_clk_sel),
				.gen3_tx_clk_sel(hssi_8g_rx_pcs_gen3_tx_clk_sel),
				.hip_mode(hssi_8g_rx_pcs_hip_mode),
				.ibm_invalid_code(hssi_8g_rx_pcs_ibm_invalid_code),
				.invalid_code_flag_only(hssi_8g_rx_pcs_invalid_code_flag_only),
				.pad_or_edb_error_replace(hssi_8g_rx_pcs_pad_or_edb_error_replace),
				.pcs_bypass(hssi_8g_rx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_rx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_rx_pcs_phase_compensation_fifo),
				.pipe_if_enable(hssi_8g_rx_pcs_pipe_if_enable),
				.pma_dw(hssi_8g_rx_pcs_pma_dw),
				.polinv_8b10b_dec(hssi_8g_rx_pcs_polinv_8b10b_dec),
				.prot_mode(hssi_8g_rx_pcs_prot_mode),
				.rate_match(hssi_8g_rx_pcs_rate_match),
				.rate_match_del_thres(hssi_8g_rx_pcs_rate_match_del_thres),
				.rate_match_empty_thres(hssi_8g_rx_pcs_rate_match_empty_thres),
				.rate_match_full_thres(hssi_8g_rx_pcs_rate_match_full_thres),
				.rate_match_ins_thres(hssi_8g_rx_pcs_rate_match_ins_thres),
				.rate_match_start_thres(hssi_8g_rx_pcs_rate_match_start_thres),
				.reconfig_settings(hssi_8g_rx_pcs_reconfig_settings),
				.rx_clk2(hssi_8g_rx_pcs_rx_clk2),
				.rx_clk_free_running(hssi_8g_rx_pcs_rx_clk_free_running),
				.rx_pcs_urst(hssi_8g_rx_pcs_rx_pcs_urst),
				.rx_rcvd_clk(hssi_8g_rx_pcs_rx_rcvd_clk),
				.rx_rd_clk(hssi_8g_rx_pcs_rx_rd_clk),
				.rx_refclk(hssi_8g_rx_pcs_rx_refclk),
				.rx_wr_clk(hssi_8g_rx_pcs_rx_wr_clk),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_rx_pcs_sup_mode),
				.symbol_swap(hssi_8g_rx_pcs_symbol_swap),
				.sync_sm_idle_eios(hssi_8g_rx_pcs_sync_sm_idle_eios),
				.test_bus_sel(hssi_8g_rx_pcs_test_bus_sel),
				.tx_rx_parallel_loopback(hssi_8g_rx_pcs_tx_rx_parallel_loopback),
				.wa_boundary_lock_ctrl(hssi_8g_rx_pcs_wa_boundary_lock_ctrl),
				.wa_clk_slip_spacing(hssi_8g_rx_pcs_wa_clk_slip_spacing),
				.wa_det_latency_sync_status_beh(hssi_8g_rx_pcs_wa_det_latency_sync_status_beh),
				.wa_disp_err_flag(hssi_8g_rx_pcs_wa_disp_err_flag),
				.wa_kchar(hssi_8g_rx_pcs_wa_kchar),
				.wa_pd(hssi_8g_rx_pcs_wa_pd),
				.wa_pd_data(hssi_8g_rx_pcs_wa_pd_data),
				.wa_pd_polarity(hssi_8g_rx_pcs_wa_pd_polarity),
				.wa_pld_controlled(hssi_8g_rx_pcs_wa_pld_controlled),
				.wa_renumber_data(hssi_8g_rx_pcs_wa_renumber_data),
				.wa_rgnumber_data(hssi_8g_rx_pcs_wa_rgnumber_data),
				.wa_rknumber_data(hssi_8g_rx_pcs_wa_rknumber_data),
				.wa_rosnumber_data(hssi_8g_rx_pcs_wa_rosnumber_data),
				.wa_rvnumber_data(hssi_8g_rx_pcs_wa_rvnumber_data),
				.wa_sync_sm_ctrl(hssi_8g_rx_pcs_wa_sync_sm_ctrl),
				.wait_cnt(hssi_8g_rx_pcs_wait_cnt)
			) inst_twentynm_hssi_8g_rx_pcs (
				// OUTPUTS
				.a1a2k1k2flag(w_hssi_8g_rx_pcs_a1a2k1k2flag),
				.avmmreaddata(w_hssi_8g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_rx_pcs_blockselect),
				.chnl_test_bus_out(w_hssi_8g_rx_pcs_chnl_test_bus_out),
				.clock_to_pld(w_hssi_8g_rx_pcs_clock_to_pld),
				.dataout(w_hssi_8g_rx_pcs_dataout),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidle_detected(w_hssi_8g_rx_pcs_eidle_detected),
				.eios_det_cdr_ctrl(w_hssi_8g_rx_pcs_eios_det_cdr_ctrl),
				.g3_rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.g3_rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.gen2ngen1(w_hssi_8g_rx_pcs_gen2ngen1),
				.parallel_rev_loopback(w_hssi_8g_rx_pcs_parallel_rev_loopback),
				.pc_fifo_empty(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.pcfifofull(w_hssi_8g_rx_pcs_pcfifofull),
				.phystatus(w_hssi_8g_rx_pcs_phystatus),
				.pipe_data(w_hssi_8g_rx_pcs_pipe_data),
				.rd_enable_out_chnl_down(w_hssi_8g_rx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_rx_pcs_rd_enable_out_chnl_up),
				.rd_ptr1_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo),
				.rd_ptr2_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo),
				.rd_ptr_rx_phfifo(w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.reset_pc_ptrs_out_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down),
				.reset_pc_ptrs_out_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up),
				.rm_fifo_empty(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.rm_fifo_full(w_hssi_8g_rx_pcs_rm_fifo_full),
				.rx_blk_start(w_hssi_8g_rx_pcs_rx_blk_start),
				.rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.rx_data_valid(w_hssi_8g_rx_pcs_rx_data_valid),
				.rx_div_sync_out_chnl_down(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down),
				.rx_div_sync_out_chnl_up(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up),
				.rx_pipe_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.rx_pipe_soft_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rx_pma_clk_gen3(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_rcvd_clk_gen3(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_rstn_sync2wrfifo_8g(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.rx_sync_hdr(w_hssi_8g_rx_pcs_rx_sync_hdr),
				.rx_we_out_chnl_down(w_hssi_8g_rx_pcs_rx_we_out_chnl_down),
				.rx_we_out_chnl_up(w_hssi_8g_rx_pcs_rx_we_out_chnl_up),
				.rxstatus(w_hssi_8g_rx_pcs_rxstatus),
				.rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.word_align_boundary(w_hssi_8g_rx_pcs_word_align_boundary),
				.wr_clk_rx_phfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_rx_phfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_rx_rmfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_rx_rmfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_data_rx_phfifo(w_hssi_8g_rx_pcs_wr_data_rx_phfifo),
				.wr_data_rx_rmfifo(w_hssi_8g_rx_pcs_wr_data_rx_rmfifo),
				.wr_en_rx_phfifo(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_rx_rmfifo(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_rx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_rx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_rx_phfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo),
				.wr_ptr_rx_rmfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo),
				.wr_rst_n_rx_phfifo(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_rx_rmfifo(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				// INPUTS
				.a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bit_reversal_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.datain({w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0]}),
				.disable_pc_fifo_byte_serdes(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4]),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.eidleinfersel({w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0]}),
				.eios_detected_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.enable_comma_detect(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.gen3_clk_sel(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.hrd_rst(1'b0),
				.inferred_rxvalid_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.pc_fifo_rd_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.pc_fifo_wrdisable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.phystatus_int(w_hssi_pipe_gen1_2_phystatus),
				.phystatus_pcs_gen3(w_hssi_pipe_gen3_phystatus),
				.pipe_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.polarity_inversion(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.rd_data1_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0]}),
				.rd_data2_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0]}),
				.rd_data_rx_phfifo({w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[3]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[3]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.reset_pc_ptrs_asn(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5]),
				.reset_pc_ptrs_in_chnl_down(in_bond_pcs8g_in_bot[12]),
				.reset_pc_ptrs_in_chnl_up(in_bond_pcs8g_in_top[12]),
				.reset_ppm_cntrs_pcs_pma(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7]),
				.rm_fifo_read_enable(1'b0),
				.rm_fifo_write_enable(1'b0),
				.rx_blk_start_pcs_gen3({w_hssi_pipe_gen3_rx_blk_start[3], w_hssi_pipe_gen3_rx_blk_start[2], w_hssi_pipe_gen3_rx_blk_start[1], w_hssi_pipe_gen3_rx_blk_start[0]}),
				.rx_data_pcs_gen3({w_hssi_pipe_gen3_rxd_8gpcs_out[63], w_hssi_pipe_gen3_rxd_8gpcs_out[62], w_hssi_pipe_gen3_rxd_8gpcs_out[61], w_hssi_pipe_gen3_rxd_8gpcs_out[60], w_hssi_pipe_gen3_rxd_8gpcs_out[59], w_hssi_pipe_gen3_rxd_8gpcs_out[58], w_hssi_pipe_gen3_rxd_8gpcs_out[57], w_hssi_pipe_gen3_rxd_8gpcs_out[56], w_hssi_pipe_gen3_rxd_8gpcs_out[55], w_hssi_pipe_gen3_rxd_8gpcs_out[54], w_hssi_pipe_gen3_rxd_8gpcs_out[53], w_hssi_pipe_gen3_rxd_8gpcs_out[52], w_hssi_pipe_gen3_rxd_8gpcs_out[51], w_hssi_pipe_gen3_rxd_8gpcs_out[50], w_hssi_pipe_gen3_rxd_8gpcs_out[49], w_hssi_pipe_gen3_rxd_8gpcs_out[48], w_hssi_pipe_gen3_rxd_8gpcs_out[47], w_hssi_pipe_gen3_rxd_8gpcs_out[46], w_hssi_pipe_gen3_rxd_8gpcs_out[45], w_hssi_pipe_gen3_rxd_8gpcs_out[44], w_hssi_pipe_gen3_rxd_8gpcs_out[43], w_hssi_pipe_gen3_rxd_8gpcs_out[42], w_hssi_pipe_gen3_rxd_8gpcs_out[41], w_hssi_pipe_gen3_rxd_8gpcs_out[40], w_hssi_pipe_gen3_rxd_8gpcs_out[39], w_hssi_pipe_gen3_rxd_8gpcs_out[38], w_hssi_pipe_gen3_rxd_8gpcs_out[37], w_hssi_pipe_gen3_rxd_8gpcs_out[36], w_hssi_pipe_gen3_rxd_8gpcs_out[35], w_hssi_pipe_gen3_rxd_8gpcs_out[34], w_hssi_pipe_gen3_rxd_8gpcs_out[33], w_hssi_pipe_gen3_rxd_8gpcs_out[32], w_hssi_pipe_gen3_rxd_8gpcs_out[31], w_hssi_pipe_gen3_rxd_8gpcs_out[30], w_hssi_pipe_gen3_rxd_8gpcs_out[29], w_hssi_pipe_gen3_rxd_8gpcs_out[28], w_hssi_pipe_gen3_rxd_8gpcs_out[27], w_hssi_pipe_gen3_rxd_8gpcs_out[26], w_hssi_pipe_gen3_rxd_8gpcs_out[25], w_hssi_pipe_gen3_rxd_8gpcs_out[24], w_hssi_pipe_gen3_rxd_8gpcs_out[23], w_hssi_pipe_gen3_rxd_8gpcs_out[22], w_hssi_pipe_gen3_rxd_8gpcs_out[21], w_hssi_pipe_gen3_rxd_8gpcs_out[20], w_hssi_pipe_gen3_rxd_8gpcs_out[19], w_hssi_pipe_gen3_rxd_8gpcs_out[18], w_hssi_pipe_gen3_rxd_8gpcs_out[17], w_hssi_pipe_gen3_rxd_8gpcs_out[16], w_hssi_pipe_gen3_rxd_8gpcs_out[15], w_hssi_pipe_gen3_rxd_8gpcs_out[14], w_hssi_pipe_gen3_rxd_8gpcs_out[13], w_hssi_pipe_gen3_rxd_8gpcs_out[12], w_hssi_pipe_gen3_rxd_8gpcs_out[11], w_hssi_pipe_gen3_rxd_8gpcs_out[10], w_hssi_pipe_gen3_rxd_8gpcs_out[9], w_hssi_pipe_gen3_rxd_8gpcs_out[8], w_hssi_pipe_gen3_rxd_8gpcs_out[7], w_hssi_pipe_gen3_rxd_8gpcs_out[6], w_hssi_pipe_gen3_rxd_8gpcs_out[5], w_hssi_pipe_gen3_rxd_8gpcs_out[4], w_hssi_pipe_gen3_rxd_8gpcs_out[3], w_hssi_pipe_gen3_rxd_8gpcs_out[2], w_hssi_pipe_gen3_rxd_8gpcs_out[1], w_hssi_pipe_gen3_rxd_8gpcs_out[0]}),
				.rx_data_valid_pcs_gen3({w_hssi_pipe_gen3_rxdataskip[3], w_hssi_pipe_gen3_rxdataskip[2], w_hssi_pipe_gen3_rxdataskip[1], w_hssi_pipe_gen3_rxdataskip[0]}),
				.rx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[1], in_bond_pcs8g_in_bot[0]}),
				.rx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[1], in_bond_pcs8g_in_top[0]}),
				.rx_pcs_rst(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.rx_sync_hdr_pcs_gen3({w_hssi_pipe_gen3_rx_sync_hdr[1], w_hssi_pipe_gen3_rx_sync_hdr[0]}),
				.rx_we_in_chnl_down({in_bond_pcs8g_in_bot[5], in_bond_pcs8g_in_bot[4]}),
				.rx_we_in_chnl_up({in_bond_pcs8g_in_top[5], in_bond_pcs8g_in_top[4]}),
				.rxstatus_int({w_hssi_pipe_gen1_2_rxstatus[2], w_hssi_pipe_gen1_2_rxstatus[1], w_hssi_pipe_gen1_2_rxstatus[0]}),
				.rxstatus_pcs_gen3({w_hssi_pipe_gen3_rxstatus[2], w_hssi_pipe_gen3_rxstatus[1], w_hssi_pipe_gen3_rxstatus[0]}),
				.rxvalid_int(w_hssi_pipe_gen1_2_rxvalid),
				.rxvalid_pcs_gen3(w_hssi_pipe_gen3_rxvalid),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.sig_det_from_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_ctrlplane_testbus({w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0]}),
				.tx_div_sync({w_hssi_8g_tx_pcs_tx_div_sync[1], w_hssi_8g_tx_pcs_tx_div_sync[0]}),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.tx_testbus({w_hssi_8g_tx_pcs_tx_testbus[19], w_hssi_8g_tx_pcs_tx_testbus[18], w_hssi_8g_tx_pcs_tx_testbus[17], w_hssi_8g_tx_pcs_tx_testbus[16], w_hssi_8g_tx_pcs_tx_testbus[15], w_hssi_8g_tx_pcs_tx_testbus[14], w_hssi_8g_tx_pcs_tx_testbus[13], w_hssi_8g_tx_pcs_tx_testbus[12], w_hssi_8g_tx_pcs_tx_testbus[11], w_hssi_8g_tx_pcs_tx_testbus[10], w_hssi_8g_tx_pcs_tx_testbus[9], w_hssi_8g_tx_pcs_tx_testbus[8], w_hssi_8g_tx_pcs_tx_testbus[7], w_hssi_8g_tx_pcs_tx_testbus[6], w_hssi_8g_tx_pcs_tx_testbus[5], w_hssi_8g_tx_pcs_tx_testbus[4], w_hssi_8g_tx_pcs_tx_testbus[3], w_hssi_8g_tx_pcs_tx_testbus[2], w_hssi_8g_tx_pcs_tx_testbus[1], w_hssi_8g_tx_pcs_tx_testbus[0]}),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[2]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[2]),
				
				// UNUSED
				.byte_deserializer_pcs_clk_div_by_2_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_wire(),
				.byte_deserializer_pcs_clk_div_by_2_wire(),
				.byte_deserializer_pcs_clk_div_by_4_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_2_reg(),
				.byte_deserializer_pld_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_4_txclk_reg(),
				.pld_8g_a1a2_k1k2_flag_reg(),
				.pld_8g_a1a2_k1k2_flag_txclk_reg(),
				.pld_8g_a1a2_size_reg(),
				.pld_8g_a1a2_size_txclk_reg(),
				.pld_8g_bitloc_rev_en_reg(),
				.pld_8g_bitloc_rev_en_txclk_reg(),
				.pld_8g_byte_rev_en_reg(),
				.pld_8g_byte_rev_en_txclk_reg(),
				.pld_8g_elecidle_reg(),
				.pld_8g_empty_rmf_lowlatency_reg(),
				.pld_8g_empty_rmf_lowlatency_txclk_reg(),
				.pld_8g_empty_rmf_reg(),
				.pld_8g_empty_rmf_txclk_reg(),
				.pld_8g_empty_rx_fifo(),
				.pld_8g_empty_rx_reg(),
				.pld_8g_empty_rx_txclk_reg(),
				.pld_8g_encdt_reg(),
				.pld_8g_encdt_txclk_reg(),
				.pld_8g_full_rmf_reg(),
				.pld_8g_full_rmf_txclk_reg(),
				.pld_8g_full_rx_fifo(),
				.pld_8g_full_rx_reg(),
				.pld_8g_full_rx_txclk_reg(),
				.pld_8g_g3_rx_pld_rst_n_reg(),
				.pld_8g_g3_rx_pld_rst_n_txclk_reg(),
				.pld_8g_rxelecidle_txclk_reg(),
				.pld_8g_rxpolarity_reg(),
				.pld_8g_rxpolarity_txclk_reg(),
				.pld_8g_wa_boundary_reg(),
				.pld_8g_wrdisable_rx_reg(),
				.pld_8g_wrdisable_rx_txclk_reg(),
				.pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_rx_clk_out_8g_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_wire(),
				.pld_rx_control_8g_reg(),
				.pld_rx_control_8g_txclk_reg(),
				.pld_rx_data_8g_reg(),
				.pld_rx_data_8g_txclk_reg(),
				.pld_syncsm_en_reg(),
				.pld_syncsm_en_txclk_reg(),
				.rm_fifo_partial_empty(),
				.rm_fifo_partial_full(),
				.sta_rx_clk2_by2_1(),
				.sta_rx_clk2_by2_1_out(),
				.sta_rx_clk2_by2_2(),
				.sta_rx_clk2_by2_2_out(),
				.sta_rx_clk2_by4_1(),
				.sta_rx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_rx_pcs_a1a2k1k2flag[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_rx_pcs_chnl_test_bus_out[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_clock_to_pld = 1'b0;
				assign w_hssi_8g_rx_pcs_dataout[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_dis_pc_byte = 1'b0;
				assign w_hssi_8g_rx_pcs_eidle_detected = 1'b0;
				assign w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_pma_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_gen2ngen1 = 1'b0;
				assign w_hssi_8g_rx_pcs_parallel_rev_loopback[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_pc_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_pcfifofull = 1'b0;
				assign w_hssi_8g_rx_pcs_phystatus = 1'b0;
				assign w_hssi_8g_rx_pcs_pipe_data[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_full = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clkslip = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_data_valid[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pma_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rxstatus[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_rxvalid = 1'b0;
				assign w_hssi_8g_rx_pcs_signal_detect_out = 1'b0;
				assign w_hssi_8g_rx_pcs_word_align_boundary[4:0] = 5'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79:0] = 80'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31:0] = 32'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_rmfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_tx_pcs
			twentynm_hssi_8g_tx_pcs #(
				.auto_speed_nego_gen2(hssi_8g_tx_pcs_auto_speed_nego_gen2),
				.bit_reversal(hssi_8g_tx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_tx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_tx_pcs_bypass_pipeline_reg),
				.byte_serializer(hssi_8g_tx_pcs_byte_serializer),
				.clock_gate_bs_enc(hssi_8g_tx_pcs_clock_gate_bs_enc),
				.clock_gate_dw_fifowr(hssi_8g_tx_pcs_clock_gate_dw_fifowr),
				.clock_gate_fiford(hssi_8g_tx_pcs_clock_gate_fiford),
				.clock_gate_sw_fifowr(hssi_8g_tx_pcs_clock_gate_sw_fifowr),
				.clock_observation_in_pld_core(hssi_8g_tx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_tx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_tx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_tx_pcs_ctrl_plane_bonding_distribution),
				.data_selection_8b10b_encoder_input(hssi_8g_tx_pcs_data_selection_8b10b_encoder_input),
				.dynamic_clk_switch(hssi_8g_tx_pcs_dynamic_clk_switch),
				.eightb_tenb_disp_ctrl(hssi_8g_tx_pcs_eightb_tenb_disp_ctrl),
				.eightb_tenb_encoder(hssi_8g_tx_pcs_eightb_tenb_encoder),
				.force_echar(hssi_8g_tx_pcs_force_echar),
				.force_kchar(hssi_8g_tx_pcs_force_kchar),
				.gen3_tx_clk_sel(hssi_8g_tx_pcs_gen3_tx_clk_sel),
				.gen3_tx_pipe_clk_sel(hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel),
				.hip_mode(hssi_8g_tx_pcs_hip_mode),
				.pcs_bypass(hssi_8g_tx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_tx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_tx_pcs_phase_compensation_fifo),
				.phfifo_write_clk_sel(hssi_8g_tx_pcs_phfifo_write_clk_sel),
				.pma_dw(hssi_8g_tx_pcs_pma_dw),
				.prot_mode(hssi_8g_tx_pcs_prot_mode),
				.reconfig_settings(hssi_8g_tx_pcs_reconfig_settings),
				.refclk_b_clk_sel(hssi_8g_tx_pcs_refclk_b_clk_sel),
				.revloop_back_rm(hssi_8g_tx_pcs_revloop_back_rm),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_tx_pcs_sup_mode),
				.symbol_swap(hssi_8g_tx_pcs_symbol_swap),
				.tx_bitslip(hssi_8g_tx_pcs_tx_bitslip),
				.tx_compliance_controlled_disparity(hssi_8g_tx_pcs_tx_compliance_controlled_disparity),
				.tx_fast_pld_reg(hssi_8g_tx_pcs_tx_fast_pld_reg),
				.txclk_freerun(hssi_8g_tx_pcs_txclk_freerun),
				.txpcs_urst(hssi_8g_tx_pcs_txpcs_urst)
			) inst_twentynm_hssi_8g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_8g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_tx_pcs_blockselect),
				.clk_out(w_hssi_8g_tx_pcs_clk_out),
				.clk_out_gen3(w_hssi_8g_tx_pcs_clk_out_gen3),
				.dataout(w_hssi_8g_tx_pcs_dataout),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.fifo_select_out_chnl_down(w_hssi_8g_tx_pcs_fifo_select_out_chnl_down),
				.fifo_select_out_chnl_up(w_hssi_8g_tx_pcs_fifo_select_out_chnl_up),
				.g3_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.g3_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
				.non_gray_eidleinfersel(w_hssi_8g_tx_pcs_non_gray_eidleinfersel),
				.ph_fifo_overflow(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.ph_fifo_underflow(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.phfifo_txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.phfifo_txmargin(w_hssi_8g_tx_pcs_phfifo_txmargin),
				.phfifo_txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				.pipe_en_rev_parallel_lpbk_out(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.pipe_power_down_out(w_hssi_8g_tx_pcs_pipe_power_down_out),
				.pipe_tx_clk_out_gen3(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pmaif_asn_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.rd_enable_out_chnl_down(w_hssi_8g_tx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_tx_pcs_rd_enable_out_chnl_up),
				.rd_ptr_tx_phfifo(w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rxpolarity_int(w_hssi_8g_tx_pcs_rxpolarity_int),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.tx_blk_start_out(w_hssi_8g_tx_pcs_tx_blk_start_out),
				.tx_clk_out_8g_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.tx_ctrlplane_testbus(w_hssi_8g_tx_pcs_tx_ctrlplane_testbus),
				.tx_data_out(w_hssi_8g_tx_pcs_tx_data_out),
				.tx_data_valid_out(w_hssi_8g_tx_pcs_tx_data_valid_out),
				.tx_datak_out(w_hssi_8g_tx_pcs_tx_datak_out),
				.tx_detect_rxloopback_int(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.tx_div_sync(w_hssi_8g_tx_pcs_tx_div_sync),
				.tx_div_sync_out_chnl_down(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down),
				.tx_div_sync_out_chnl_up(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up),
				.tx_pipe_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.tx_pipe_electidle(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_soft_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.tx_sync_hdr_out(w_hssi_8g_tx_pcs_tx_sync_hdr_out),
				.tx_testbus(w_hssi_8g_tx_pcs_tx_testbus),
				.txcompliance_out(w_hssi_8g_tx_pcs_txcompliance_out),
				.txelecidle_out(w_hssi_8g_tx_pcs_txelecidle_out),
				.wr_clk_tx_phfifo_dw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_tx_phfifo_sw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_data_tx_phfifo(w_hssi_8g_tx_pcs_wr_data_tx_phfifo),
				.wr_en_tx_phfifo(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_tx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_tx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_tx_phfifo(w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo),
				.wr_rst_n_tx_phfifo(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bitslip_boundary_select({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0]}),
				.clk_sel_gen3(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.coreclk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.datain({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.detectrxloopin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidleinfersel({w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0]}),
				.en_rev_parallel_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.fifo_select_in_chnl_down({in_bond_pcs8g_in_bot[11], in_bond_pcs8g_in_bot[10]}),
				.fifo_select_in_chnl_up({in_bond_pcs8g_in_top[11], in_bond_pcs8g_in_top[10]}),
				.hrdrst(1'b0),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.ph_fifo_rd_disable(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.pipe_en_rev_parallel_lpbk_in(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.pipe_tx_deemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.pipe_tx_margin({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0]}),
				.powerdn({w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0]}),
				.rate_switch(w_hssi_8g_rx_pcs_gen2ngen1),
				.rd_data_tx_phfifo({w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[9]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[9]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.rev_parallel_lpbk_data({w_hssi_8g_rx_pcs_parallel_rev_loopback[19], w_hssi_8g_rx_pcs_parallel_rev_loopback[18], w_hssi_8g_rx_pcs_parallel_rev_loopback[17], w_hssi_8g_rx_pcs_parallel_rev_loopback[16], w_hssi_8g_rx_pcs_parallel_rev_loopback[15], w_hssi_8g_rx_pcs_parallel_rev_loopback[14], w_hssi_8g_rx_pcs_parallel_rev_loopback[13], w_hssi_8g_rx_pcs_parallel_rev_loopback[12], w_hssi_8g_rx_pcs_parallel_rev_loopback[11], w_hssi_8g_rx_pcs_parallel_rev_loopback[10], w_hssi_8g_rx_pcs_parallel_rev_loopback[9], w_hssi_8g_rx_pcs_parallel_rev_loopback[8], w_hssi_8g_rx_pcs_parallel_rev_loopback[7], w_hssi_8g_rx_pcs_parallel_rev_loopback[6], w_hssi_8g_rx_pcs_parallel_rev_loopback[5], w_hssi_8g_rx_pcs_parallel_rev_loopback[4], w_hssi_8g_rx_pcs_parallel_rev_loopback[3], w_hssi_8g_rx_pcs_parallel_rev_loopback[2], w_hssi_8g_rx_pcs_parallel_rev_loopback[1], w_hssi_8g_rx_pcs_parallel_rev_loopback[0]}),
				.rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.tx_blk_start({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0]}),
				.tx_data_valid({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0]}),
				.tx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[7], in_bond_pcs8g_in_bot[6]}),
				.tx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[7], in_bond_pcs8g_in_top[6]}),
				.tx_pcs_reset(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.tx_sync_hdr({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0]}),
				.txd_fast_reg({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0]}),
				.txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[8]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[8]),
				.wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				
				// UNUSED
				.byte_serializer_pcs_clk_div_by_2_reg(),
				.byte_serializer_pcs_clk_div_by_2_wire(),
				.byte_serializer_pcs_clk_div_by_4_reg(),
				.byte_serializer_pld_clk_div_by_2_reg(),
				.byte_serializer_pld_clk_div_by_4_reg(),
				.pld_8g_empty_tx_fifo(),
				.pld_8g_empty_tx_reg(),
				.pld_8g_full_tx_fifo(),
				.pld_8g_full_tx_reg(),
				.pld_8g_g3_tx_pld_rst_n_reg(),
				.pld_8g_rddisable_tx_reg(),
				.pld_8g_tx_boundary_sel_reg(),
				.pld_pcs_tx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_tx_clk_out_8g_wire(),
				.pld_tx_data_8g_fifo(),
				.pld_tx_data_lo_8g_reg(),
				.sta_tx_clk2_by2_1(),
				.sta_tx_clk2_by2_1_out(),
				.sta_tx_clk2_by4_1(),
				.sta_tx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_dataout[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_dyn_clk_switch_n = 1'b1;		// Override default tieoff
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_g3_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_overflow = 1'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_underflow = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txdeemph = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txmargin[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txswing = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_power_down_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_pmaif_asn_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_refclk_b = 1'b0;
				assign w_hssi_8g_tx_pcs_refclk_b_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_rxpolarity_int = 1'b0;
				assign w_hssi_8g_tx_pcs_soft_reset_wclk1_n = 1'b0;
				assign w_hssi_8g_tx_pcs_sw_fifo_wr_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_blk_start_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_tx_data_out[31:0] = 32'b0;
				assign w_hssi_8g_tx_pcs_tx_data_valid_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_datak_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_detect_rxloopback_int = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_electidle = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_sync_hdr_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_txcompliance_out = 1'b0;
				assign w_hssi_8g_tx_pcs_txelecidle_out = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63:0] = 64'b0;
				assign w_hssi_8g_tx_pcs_wr_en_tx_phfifo = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pcs_pma_interface
			twentynm_hssi_common_pcs_pma_interface #(
				.asn_clk_enable(hssi_common_pcs_pma_interface_asn_clk_enable),
				.asn_enable(hssi_common_pcs_pma_interface_asn_enable),
				.block_sel(hssi_common_pcs_pma_interface_block_sel),
				.bypass_early_eios(hssi_common_pcs_pma_interface_bypass_early_eios),
				.bypass_pcie_switch(hssi_common_pcs_pma_interface_bypass_pcie_switch),
				.bypass_pma_ltr(hssi_common_pcs_pma_interface_bypass_pma_ltr),
				.bypass_pma_sw_done(hssi_common_pcs_pma_interface_bypass_pma_sw_done),
				.bypass_ppm_lock(hssi_common_pcs_pma_interface_bypass_ppm_lock),
				.bypass_send_syncp_fbkp(hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp),
				.bypass_txdetectrx(hssi_common_pcs_pma_interface_bypass_txdetectrx),
				.cdr_control(hssi_common_pcs_pma_interface_cdr_control),
				.cid_enable(hssi_common_pcs_pma_interface_cid_enable),
				.cp_cons_sel(hssi_common_pcs_pma_interface_cp_cons_sel),
				.cp_dwn_mstr(hssi_common_pcs_pma_interface_cp_dwn_mstr),
				.cp_up_mstr(hssi_common_pcs_pma_interface_cp_up_mstr),
				.ctrl_plane_bonding(hssi_common_pcs_pma_interface_ctrl_plane_bonding),
				.data_mask_count(hssi_common_pcs_pma_interface_data_mask_count),
				.data_mask_count_multi(hssi_common_pcs_pma_interface_data_mask_count_multi),
				.dft_observation_clock_selection(hssi_common_pcs_pma_interface_dft_observation_clock_selection),
				.early_eios_counter(hssi_common_pcs_pma_interface_early_eios_counter),
				.force_freqdet(hssi_common_pcs_pma_interface_force_freqdet),
				.free_run_clk_enable(hssi_common_pcs_pma_interface_free_run_clk_enable),
				.ignore_sigdet_g23(hssi_common_pcs_pma_interface_ignore_sigdet_g23),
				.pc_en_counter(hssi_common_pcs_pma_interface_pc_en_counter),
				.pc_rst_counter(hssi_common_pcs_pma_interface_pc_rst_counter),
				.pcie_hip_mode(hssi_common_pcs_pma_interface_pcie_hip_mode),
				.ph_fifo_reg_mode(hssi_common_pcs_pma_interface_ph_fifo_reg_mode),
				.phfifo_flush_wait(hssi_common_pcs_pma_interface_phfifo_flush_wait),
				.pipe_if_g3pcs(hssi_common_pcs_pma_interface_pipe_if_g3pcs),
				.pma_done_counter(hssi_common_pcs_pma_interface_pma_done_counter),
				.pma_if_dft_en(hssi_common_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_common_pcs_pma_interface_pma_if_dft_val),
				.ppm_cnt_rst(hssi_common_pcs_pma_interface_ppm_cnt_rst),
				.ppm_deassert_early(hssi_common_pcs_pma_interface_ppm_deassert_early),
				.ppm_det_buckets(hssi_common_pcs_pma_interface_ppm_det_buckets),
				.ppm_gen1_2_cnt(hssi_common_pcs_pma_interface_ppm_gen1_2_cnt),
				.ppm_post_eidle_delay(hssi_common_pcs_pma_interface_ppm_post_eidle_delay),
				.ppmsel(hssi_common_pcs_pma_interface_ppmsel),
				.prot_mode(hssi_common_pcs_pma_interface_prot_mode),
				.reconfig_settings(hssi_common_pcs_pma_interface_reconfig_settings),
				.rxvalid_mask(hssi_common_pcs_pma_interface_rxvalid_mask),
				.sigdet_wait_counter(hssi_common_pcs_pma_interface_sigdet_wait_counter),
				.sigdet_wait_counter_multi(hssi_common_pcs_pma_interface_sigdet_wait_counter_multi),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sim_mode(hssi_common_pcs_pma_interface_sim_mode),
				.spd_chg_rst_wait_cnt_en(hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en),
				.sup_mode(hssi_common_pcs_pma_interface_sup_mode),
				.testout_sel(hssi_common_pcs_pma_interface_testout_sel),
				.wait_clk_on_off_timer(hssi_common_pcs_pma_interface_wait_clk_on_off_timer),
				.wait_pipe_synchronizing(hssi_common_pcs_pma_interface_wait_pipe_synchronizing),
				.wait_send_syncp_fbkp(hssi_common_pcs_pma_interface_wait_send_syncp_fbkp)
			) inst_twentynm_hssi_common_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_common_pcs_pma_interface_blockselect),
				.int_pmaif_8g_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in),
				.int_pmaif_8g_eios_detected(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.int_pmaif_8g_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.int_pmaif_8g_power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.int_pmaif_g3_pcs_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in),
				.int_pmaif_pldif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pmaif_pldif_pcie_sw_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done),
				.int_pmaif_pldif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pmaif_pldif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pmaif_pldif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pmaif_pldif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pmaif_pldif_pma_reserved_in(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in),
				.int_pmaif_pldif_test_out(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out),
				.int_pmaif_pldif_testbus(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus),
				.pma_adapt_start(w_hssi_common_pcs_pma_interface_pma_adapt_start),
				.pma_atpg_los_en_n(w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n),
				.pma_csr_test_dis(w_hssi_common_pcs_pma_interface_pma_csr_test_dis),
				.pma_current_coeff(w_hssi_common_pcs_pma_interface_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_common_pcs_pma_interface_pma_current_rxpreset),
				.pma_early_eios(w_hssi_common_pcs_pma_interface_pma_early_eios),
				.pma_interface_select(w_hssi_common_pcs_pma_interface_pma_interface_select),
				.pma_ltd_b(w_hssi_common_pcs_pma_interface_pma_ltd_b),
				.pma_ltr(w_hssi_common_pcs_pma_interface_pma_ltr),
				.pma_nfrzdrv(w_hssi_common_pcs_pma_interface_pma_nfrzdrv),
				.pma_nrpi_freeze(w_hssi_common_pcs_pma_interface_pma_nrpi_freeze),
				.pma_pcie_switch(w_hssi_common_pcs_pma_interface_pma_pcie_switch),
				.pma_ppm_lock(w_hssi_common_pcs_pma_interface_pma_ppm_lock),
				.pma_reserved_out(w_hssi_common_pcs_pma_interface_pma_reserved_out),
				.pma_rs_lpbk_b(w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b),
				.pma_rx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup),
				.pma_scan_mode_n(w_hssi_common_pcs_pma_interface_pma_scan_mode_n),
				.pma_scan_shift_n(w_hssi_common_pcs_pma_interface_pma_scan_shift_n),
				.pma_tx_bitslip(w_hssi_common_pcs_pma_interface_pma_tx_bitslip),
				.pma_tx_bonding_rstb(w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb),
				.pma_tx_qpi_pulldn(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn),
				.pma_tx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup),
				.pma_tx_txdetectrx(w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx),
				.pmaif_bundling_out_down(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down),
				.pmaif_bundling_out_up(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_8g_current_coeff({w_hssi_pipe_gen1_2_current_coeff[17], w_hssi_pipe_gen1_2_current_coeff[16], w_hssi_pipe_gen1_2_current_coeff[15], w_hssi_pipe_gen1_2_current_coeff[14], w_hssi_pipe_gen1_2_current_coeff[13], w_hssi_pipe_gen1_2_current_coeff[12], w_hssi_pipe_gen1_2_current_coeff[11], w_hssi_pipe_gen1_2_current_coeff[10], w_hssi_pipe_gen1_2_current_coeff[9], w_hssi_pipe_gen1_2_current_coeff[8], w_hssi_pipe_gen1_2_current_coeff[7], w_hssi_pipe_gen1_2_current_coeff[6], w_hssi_pipe_gen1_2_current_coeff[5], w_hssi_pipe_gen1_2_current_coeff[4], w_hssi_pipe_gen1_2_current_coeff[3], w_hssi_pipe_gen1_2_current_coeff[2], w_hssi_pipe_gen1_2_current_coeff[1], w_hssi_pipe_gen1_2_current_coeff[0]}),
				.int_pmaif_8g_eios_det({w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0]}),
				.int_pmaif_8g_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.int_pmaif_8g_rev_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.int_pmaif_8g_tx_clk_out_gen3(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.int_pmaif_8g_txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				.int_pmaif_g3_eios_det({w_hssi_gen3_rx_pcs_ei_det_int, w_hssi_gen3_rx_pcs_ei_partial_det_int, w_hssi_gen3_rx_pcs_i_det_int}),
				.int_pmaif_g3_pma_current_coeff({w_hssi_pipe_gen3_pma_current_coeff[17], w_hssi_pipe_gen3_pma_current_coeff[16], w_hssi_pipe_gen3_pma_current_coeff[15], w_hssi_pipe_gen3_pma_current_coeff[14], w_hssi_pipe_gen3_pma_current_coeff[13], w_hssi_pipe_gen3_pma_current_coeff[12], w_hssi_pipe_gen3_pma_current_coeff[11], w_hssi_pipe_gen3_pma_current_coeff[10], w_hssi_pipe_gen3_pma_current_coeff[9], w_hssi_pipe_gen3_pma_current_coeff[8], w_hssi_pipe_gen3_pma_current_coeff[7], w_hssi_pipe_gen3_pma_current_coeff[6], w_hssi_pipe_gen3_pma_current_coeff[5], w_hssi_pipe_gen3_pma_current_coeff[4], w_hssi_pipe_gen3_pma_current_coeff[3], w_hssi_pipe_gen3_pma_current_coeff[2], w_hssi_pipe_gen3_pma_current_coeff[1], w_hssi_pipe_gen3_pma_current_coeff[0]}),
				.int_pmaif_g3_pma_current_rxpreset({w_hssi_pipe_gen3_pma_current_rxpreset[2], w_hssi_pipe_gen3_pma_current_rxpreset[1], w_hssi_pipe_gen3_pma_current_rxpreset[0]}),
				.int_pmaif_g3_pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.int_pmaif_g3_rev_lpbk(w_hssi_pipe_gen3_rev_lpbk_int),
				.int_pmaif_pldif_8g_tx_pld_rstn(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pmaif_pldif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pmaif_pldif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pmaif_pldif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pmaif_pldif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pmaif_pldif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pmaif_pldif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pmaif_pldif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pmaif_pldif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pmaif_pldif_pcie_switch({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0]}),
				.int_pmaif_pldif_pma_reserved_out({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0]}),
				.int_pmaif_pldif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pmaif_pldif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pmaif_pldif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pmaif_pldif_rate({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0]}),
				.int_pmaif_pldif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pmaif_pldif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pmaif_pldif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.int_pmaif_pldif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pmaif_pldif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pmaif_pldif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pmaif_pldif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pmaif_pldif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pmaif_pldif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.int_tx_dft_obsrv_clk({w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0]}),
				.iocsr_clk(in_iocsr_clk),
				.iocsr_config({in_iocsr_config[5], in_iocsr_config[4], in_iocsr_config[3], in_iocsr_config[2], in_iocsr_config[1], in_iocsr_config[0]}),
				.iocsr_rdy(in_iocsr_rdy),
				.iocsr_rdy_dly(in_iocsr_rdy_dly),
				.pma_adapt_done(in_pma_adapt_done),
				.pma_clklow(in_pma_clklow),
				.pma_fref(in_pma_fref),
				.pma_hclk(in_pma_hclk),
				.pma_pcie_sw_done({in_pma_pcie_sw_done[1], in_pma_pcie_sw_done[0]}),
				.pma_pfdmode_lock(in_pma_pfdmode_lock),
				.pma_reserved_in({in_pma_reserved_in[4], in_pma_reserved_in[3], in_pma_reserved_in[2], in_pma_reserved_in[1], in_pma_reserved_in[0]}),
				.pma_signal_det(in_pma_signal_det),
				.pma_testbus({in_pma_testbus[7], in_pma_testbus[6], in_pma_testbus[5], in_pma_testbus[4], in_pma_testbus[3], in_pma_testbus[2], in_pma_testbus[1], in_pma_testbus[0]}),
				.pmaif_bundling_in_down({in_bond_pmaif_in_bot[11], in_bond_pmaif_in_bot[10], in_bond_pmaif_in_bot[9], in_bond_pmaif_in_bot[8], in_bond_pmaif_in_bot[7], in_bond_pmaif_in_bot[6], in_bond_pmaif_in_bot[5], in_bond_pmaif_in_bot[4], in_bond_pmaif_in_bot[3], in_bond_pmaif_in_bot[2], in_bond_pmaif_in_bot[1], in_bond_pmaif_in_bot[0]}),
				.pmaif_bundling_in_up({in_bond_pmaif_in_top[11], in_bond_pmaif_in_top[10], in_bond_pmaif_in_top[9], in_bond_pmaif_in_top[8], in_bond_pmaif_in_top[7], in_bond_pmaif_in_top[6], in_bond_pmaif_in_top[5], in_bond_pmaif_in_top[4], in_bond_pmaif_in_top[3], in_bond_pmaif_in_top[2], in_bond_pmaif_in_top[1], in_bond_pmaif_in_top[0]}),
				.rx_pmaif_test_out({w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0]}),
				.rx_prbs_ver_test({w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0]}),
				.tx_prbs_gen_test({w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0]}),
				.uhsif_test_out_1({w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0]}),
				.uhsif_test_out_2({w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0]}),
				.uhsif_test_out_3({w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0]}),
				
				// UNUSED
				.int_pmaif_avmm_iocsr_clk(),
				.int_pmaif_avmm_iocsr_config(),
				.int_pmaif_avmm_iocsr_rdy(),
				.int_pmaif_avmm_iocsr_rdy_dly(),
				.int_pmaif_pldif_interface_select(),
				.pma_tx_pma_syncp(),
				.sta_pma_hclk_by2()
			);
		end // if generate
		else begin
				assign w_hssi_common_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19:0] = 20'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_pma_adapt_start = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_csr_test_dis = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pcs_pma_interface_pma_early_eios = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_interface_select[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltd_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltr = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nfrzdrv = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nrpi_freeze = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ppm_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_tx_bitslip = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx = in_pld_pma_txdetectrx;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11:0] = 12'b0;
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11:0] = 12'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pld_pcs_interface
			twentynm_hssi_common_pld_pcs_interface #(
				.dft_clk_out_en(hssi_common_pld_pcs_interface_dft_clk_out_en),
				.dft_clk_out_sel(hssi_common_pld_pcs_interface_dft_clk_out_sel),
				.hrdrstctrl_en(hssi_common_pld_pcs_interface_hrdrstctrl_en),
				.pcs_testbus_block_sel(hssi_common_pld_pcs_interface_pcs_testbus_block_sel),
				.reconfig_settings(hssi_common_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm5es" )       //PARAM_HIDE
			) inst_twentynm_hssi_common_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_common_pld_pcs_interface_blockselect),
				.hip_cmn_clk(w_hssi_common_pld_pcs_interface_hip_cmn_clk),
				.hip_cmn_ctrl(w_hssi_common_pld_pcs_interface_hip_cmn_ctrl),
				.hip_iocsr_rdy(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy),
				.hip_iocsr_rdy_dly(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly),
				.hip_nfrzdrv(w_hssi_common_pld_pcs_interface_hip_nfrzdrv),
				.hip_npor(w_hssi_common_pld_pcs_interface_hip_npor),
				.hip_usermode(w_hssi_common_pld_pcs_interface_hip_usermode),
				.int_pldif_10g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.int_pldif_10g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.int_pldif_8g_eidleinfersel(w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel),
				.int_pldif_8g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.int_pldif_8g_refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.int_pldif_8g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.int_pldif_g3_current_coeff(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff),
				.int_pldif_g3_current_rxpreset(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset),
				.int_pldif_krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.int_pldif_krfec_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.int_pldif_krfec_scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				.int_pldif_mem_atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.int_pldif_mem_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.int_pldif_pmaif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pldif_pmaif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pldif_pmaif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pldif_pmaif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pldif_pmaif_eye_monitor(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor),
				.int_pldif_pmaif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pldif_pmaif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pldif_pmaif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pldif_pmaif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pldif_pmaif_pcie_switch(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch),
				.int_pldif_pmaif_pma_reserved_out(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out),
				.int_pldif_pmaif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pldif_pmaif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pldif_pmaif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pldif_pmaif_rate(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate),
				.int_pldif_pmaif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pldif_pmaif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pldif_pmaif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pldif_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_pldif_pmaif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pldif_pmaif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pldif_pmaif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pldif_pmaif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pldif_pmaif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pldif_pmaif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pldif_pmaif_uhsif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.pld_pma_adapt_done(w_hssi_common_pld_pcs_interface_pld_pma_adapt_done),
				.pld_pma_clklow(w_hssi_common_pld_pcs_interface_pld_pma_clklow),
				.pld_pma_fref(w_hssi_common_pld_pcs_interface_pld_pma_fref),
				.pld_pma_hclk(w_hssi_common_pld_pcs_interface_pld_pma_hclk),
				.pld_pma_pcie_sw_done(w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done),
				.pld_pma_pfdmode_lock(w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock),
				.pld_pma_reserved_in(w_hssi_common_pld_pcs_interface_pld_pma_reserved_in),
				.pld_pma_rx_detect_valid(w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid),
				.pld_pma_rx_found(w_hssi_common_pld_pcs_interface_pld_pma_rx_found),
				.pld_pma_rxpll_lock(w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock),
				.pld_pma_testbus(w_hssi_common_pld_pcs_interface_pld_pma_testbus),
				.pld_pmaif_mask_tx_pll(w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll),
				.pld_reserved_out(w_hssi_common_pld_pcs_interface_pld_reserved_out),
				.pld_test_data(w_hssi_common_pld_pcs_interface_pld_test_data),
				.pld_uhsif_lock(w_hssi_common_pld_pcs_interface_pld_uhsif_lock),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.int_pldif_10g_test_data({w_hssi_10g_tx_pcs_tx_test_data[19], w_hssi_10g_tx_pcs_tx_test_data[18], w_hssi_10g_tx_pcs_tx_test_data[17], w_hssi_10g_tx_pcs_tx_test_data[16], w_hssi_10g_tx_pcs_tx_test_data[15], w_hssi_10g_tx_pcs_tx_test_data[14], w_hssi_10g_tx_pcs_tx_test_data[13], w_hssi_10g_tx_pcs_tx_test_data[12], w_hssi_10g_tx_pcs_tx_test_data[11], w_hssi_10g_tx_pcs_tx_test_data[10], w_hssi_10g_tx_pcs_tx_test_data[9], w_hssi_10g_tx_pcs_tx_test_data[8], w_hssi_10g_tx_pcs_tx_test_data[7], w_hssi_10g_tx_pcs_tx_test_data[6], w_hssi_10g_tx_pcs_tx_test_data[5], w_hssi_10g_tx_pcs_tx_test_data[4], w_hssi_10g_tx_pcs_tx_test_data[3], w_hssi_10g_tx_pcs_tx_test_data[2], w_hssi_10g_tx_pcs_tx_test_data[1], w_hssi_10g_tx_pcs_tx_test_data[0]}),
				.int_pldif_10g_tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.int_pldif_8g_chnl_test_bus_out({w_hssi_8g_rx_pcs_chnl_test_bus_out[19], w_hssi_8g_rx_pcs_chnl_test_bus_out[18], w_hssi_8g_rx_pcs_chnl_test_bus_out[17], w_hssi_8g_rx_pcs_chnl_test_bus_out[16], w_hssi_8g_rx_pcs_chnl_test_bus_out[15], w_hssi_8g_rx_pcs_chnl_test_bus_out[14], w_hssi_8g_rx_pcs_chnl_test_bus_out[13], w_hssi_8g_rx_pcs_chnl_test_bus_out[12], w_hssi_8g_rx_pcs_chnl_test_bus_out[11], w_hssi_8g_rx_pcs_chnl_test_bus_out[10], w_hssi_8g_rx_pcs_chnl_test_bus_out[9], w_hssi_8g_rx_pcs_chnl_test_bus_out[8], w_hssi_8g_rx_pcs_chnl_test_bus_out[7], w_hssi_8g_rx_pcs_chnl_test_bus_out[6], w_hssi_8g_rx_pcs_chnl_test_bus_out[5], w_hssi_8g_rx_pcs_chnl_test_bus_out[4], w_hssi_8g_rx_pcs_chnl_test_bus_out[3], w_hssi_8g_rx_pcs_chnl_test_bus_out[2], w_hssi_8g_rx_pcs_chnl_test_bus_out[1], w_hssi_8g_rx_pcs_chnl_test_bus_out[0]}),
				.int_pldif_8g_rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.int_pldif_8g_tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.int_pldif_g3_test_out({w_hssi_pipe_gen3_test_out[19], w_hssi_pipe_gen3_test_out[18], w_hssi_pipe_gen3_test_out[17], w_hssi_pipe_gen3_test_out[16], w_hssi_pipe_gen3_test_out[15], w_hssi_pipe_gen3_test_out[14], w_hssi_pipe_gen3_test_out[13], w_hssi_pipe_gen3_test_out[12], w_hssi_pipe_gen3_test_out[11], w_hssi_pipe_gen3_test_out[10], w_hssi_pipe_gen3_test_out[9], w_hssi_pipe_gen3_test_out[8], w_hssi_pipe_gen3_test_out[7], w_hssi_pipe_gen3_test_out[6], w_hssi_pipe_gen3_test_out[5], w_hssi_pipe_gen3_test_out[4], w_hssi_pipe_gen3_test_out[3], w_hssi_pipe_gen3_test_out[2], w_hssi_pipe_gen3_test_out[1], w_hssi_pipe_gen3_test_out[0]}),
				.int_pldif_krfec_test_data({w_hssi_krfec_tx_pcs_tx_test_data[19], w_hssi_krfec_tx_pcs_tx_test_data[18], w_hssi_krfec_tx_pcs_tx_test_data[17], w_hssi_krfec_tx_pcs_tx_test_data[16], w_hssi_krfec_tx_pcs_tx_test_data[15], w_hssi_krfec_tx_pcs_tx_test_data[14], w_hssi_krfec_tx_pcs_tx_test_data[13], w_hssi_krfec_tx_pcs_tx_test_data[12], w_hssi_krfec_tx_pcs_tx_test_data[11], w_hssi_krfec_tx_pcs_tx_test_data[10], w_hssi_krfec_tx_pcs_tx_test_data[9], w_hssi_krfec_tx_pcs_tx_test_data[8], w_hssi_krfec_tx_pcs_tx_test_data[7], w_hssi_krfec_tx_pcs_tx_test_data[6], w_hssi_krfec_tx_pcs_tx_test_data[5], w_hssi_krfec_tx_pcs_tx_test_data[4], w_hssi_krfec_tx_pcs_tx_test_data[3], w_hssi_krfec_tx_pcs_tx_test_data[2], w_hssi_krfec_tx_pcs_tx_test_data[1], w_hssi_krfec_tx_pcs_tx_test_data[0]}),
				.int_pldif_pmaif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pldif_pmaif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pldif_pmaif_pcie_sw_done({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0]}),
				.int_pldif_pmaif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pldif_pmaif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pldif_pmaif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pldif_pmaif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pldif_pmaif_pma_reserved_in({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0]}),
				.int_pldif_pmaif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pldif_pmaif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_test_out({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0]}),
				.int_pldif_pmaif_testbus({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0]}),
				.int_pldif_pmaif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.pld_8g_eidleinfersel({in_pld_8g_eidleinfersel[2], in_pld_8g_eidleinfersel[1], in_pld_8g_eidleinfersel[0]}),
				.pld_8g_refclk_dig2(in_pld_8g_refclk_dig2),
				.pld_atpg_los_en_n(in_pld_atpg_los_en_n),
				.pld_g3_current_coeff({in_pld_g3_current_coeff[17], in_pld_g3_current_coeff[16], in_pld_g3_current_coeff[15], in_pld_g3_current_coeff[14], in_pld_g3_current_coeff[13], in_pld_g3_current_coeff[12], in_pld_g3_current_coeff[11], in_pld_g3_current_coeff[10], in_pld_g3_current_coeff[9], in_pld_g3_current_coeff[8], in_pld_g3_current_coeff[7], in_pld_g3_current_coeff[6], in_pld_g3_current_coeff[5], in_pld_g3_current_coeff[4], in_pld_g3_current_coeff[3], in_pld_g3_current_coeff[2], in_pld_g3_current_coeff[1], in_pld_g3_current_coeff[0]}),
				.pld_g3_current_rxpreset({in_pld_g3_current_rxpreset[2], in_pld_g3_current_rxpreset[1], in_pld_g3_current_rxpreset[0]}),
				.pld_ltr(in_pld_ltr),
				.pld_mem_krfec_atpg_rst_n(in_pld_mem_krfec_atpg_rst_n),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pcs_refclk_dig(in_pld_pcs_refclk_dig),
				.pld_pma_adapt_start(in_pld_pma_adapt_start),
				.pld_pma_csr_test_dis(in_pld_pma_csr_test_dis),
				.pld_pma_early_eios(in_pld_pma_early_eios),
				.pld_pma_eye_monitor({in_pld_pma_eye_monitor[5], in_pld_pma_eye_monitor[4], in_pld_pma_eye_monitor[3], in_pld_pma_eye_monitor[2], in_pld_pma_eye_monitor[1], in_pld_pma_eye_monitor[0]}),
				.pld_pma_ltd_b(in_pld_pma_ltd_b),
				.pld_pma_nrpi_freeze(in_pld_pma_nrpi_freeze),
				.pld_pma_pcie_switch({in_pld_pma_pcie_switch[1], in_pld_pma_pcie_switch[0]}),
				.pld_pma_ppm_lock(in_pld_pma_ppm_lock),
				.pld_pma_reserved_out({in_pld_pma_reserved_out[4], in_pld_pma_reserved_out[3], in_pld_pma_reserved_out[2], in_pld_pma_reserved_out[1], in_pld_pma_reserved_out[0]}),
				.pld_pma_rs_lpbk_b(in_pld_pma_rs_lpbk_b),
				.pld_pma_rx_qpi_pullup(in_pld_pma_rx_qpi_pullup),
				.pld_pma_tx_bitslip(in_pld_pma_tx_bitslip),
				.pld_pma_tx_bonding_rstb(in_pld_pma_tx_bonding_rstb),
				.pld_pma_tx_qpi_pulldn(in_pld_pma_tx_qpi_pulldn),
				.pld_pma_tx_qpi_pullup(in_pld_pma_tx_qpi_pullup),
				.pld_pma_txdetectrx(in_pld_pma_txdetectrx),
				.pld_rate({in_pld_rate[1], in_pld_rate[0]}),
				.pld_reserved_in({in_pld_reserved_in[9], in_pld_reserved_in[8], in_pld_reserved_in[7], in_pld_reserved_in[6], in_pld_reserved_in[5], in_pld_reserved_in[4], in_pld_reserved_in[3], in_pld_reserved_in[2], in_pld_reserved_in[1], in_pld_reserved_in[0]}),
				.pld_scan_mode_n(in_pld_scan_mode_n),
				.pld_scan_shift_n(in_pld_scan_shift_n),
				
				// UNUSED
				.int_pldif_8g_ltr(),
				.int_pldif_avmm_pld_avmm1_request(),
				.int_pldif_avmm_pld_avmm2_request(),
				.int_pldif_avmm_refclk_dig_en(),
				.int_pldif_g3_scan_mode_n(),
				.pld_8g_eidleinfersel_fifo(),
				.pld_8g_eidleinfersel_reg(),
				.pld_partial_reconfig_fifo(),
				.pld_partial_reconfig_rx_div_by_2_rxclk_wire(),
				.pld_partial_reconfig_rx_div_by_2_txclk_wire(),
				.pld_partial_reconfig_rxclk_reg(),
				.pld_partial_reconfig_tx_div_by_2_wire(),
				.pld_partial_reconfig_txclk_reg(),
				.pld_rate_reg(),
				.pld_test_data_reg()
			);
		end // if generate
		else begin
				assign w_hssi_common_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_clk[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_npor = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_usermode = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2 = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_adapt_done = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_clklow = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_fref = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_hclk = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_found = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_testbus[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_reserved_out[9:0] = 10'b0;
				assign w_hssi_common_pld_pcs_interface_pld_test_data[19:0] = 20'b0;
				assign w_hssi_common_pld_pcs_interface_pld_uhsif_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_scan_mode_n = 1'b1;		// Override default tieoff
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_rx_pcs
			twentynm_hssi_fifo_rx_pcs #(
				.double_read_mode(hssi_fifo_rx_pcs_double_read_mode),
				.prot_mode(hssi_fifo_rx_pcs_prot_mode),
				.silicon_rev( "20nm5es" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_rx_pcs_blockselect),
				.data_out2_10g(w_hssi_fifo_rx_pcs_data_out2_10g),
				.data_out2_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp),
				.data_out_10g(w_hssi_fifo_rx_pcs_data_out_10g),
				.data_out_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out_8g_clock_comp),
				.data_out_8g_phase_comp(w_hssi_fifo_rx_pcs_data_out_8g_phase_comp),
				.data_out_gen3(w_hssi_fifo_rx_pcs_data_out_gen3),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_data[73], w_hssi_10g_rx_pcs_rx_fifo_wr_data[72], w_hssi_10g_rx_pcs_rx_fifo_wr_data[71], w_hssi_10g_rx_pcs_rx_fifo_wr_data[70], w_hssi_10g_rx_pcs_rx_fifo_wr_data[69], w_hssi_10g_rx_pcs_rx_fifo_wr_data[68], w_hssi_10g_rx_pcs_rx_fifo_wr_data[67], w_hssi_10g_rx_pcs_rx_fifo_wr_data[66], w_hssi_10g_rx_pcs_rx_fifo_wr_data[65], w_hssi_10g_rx_pcs_rx_fifo_wr_data[64], w_hssi_10g_rx_pcs_rx_fifo_wr_data[63], w_hssi_10g_rx_pcs_rx_fifo_wr_data[62], w_hssi_10g_rx_pcs_rx_fifo_wr_data[61], w_hssi_10g_rx_pcs_rx_fifo_wr_data[60], w_hssi_10g_rx_pcs_rx_fifo_wr_data[59], w_hssi_10g_rx_pcs_rx_fifo_wr_data[58], w_hssi_10g_rx_pcs_rx_fifo_wr_data[57], w_hssi_10g_rx_pcs_rx_fifo_wr_data[56], w_hssi_10g_rx_pcs_rx_fifo_wr_data[55], w_hssi_10g_rx_pcs_rx_fifo_wr_data[54], w_hssi_10g_rx_pcs_rx_fifo_wr_data[53], w_hssi_10g_rx_pcs_rx_fifo_wr_data[52], w_hssi_10g_rx_pcs_rx_fifo_wr_data[51], w_hssi_10g_rx_pcs_rx_fifo_wr_data[50], w_hssi_10g_rx_pcs_rx_fifo_wr_data[49], w_hssi_10g_rx_pcs_rx_fifo_wr_data[48], w_hssi_10g_rx_pcs_rx_fifo_wr_data[47], w_hssi_10g_rx_pcs_rx_fifo_wr_data[46], w_hssi_10g_rx_pcs_rx_fifo_wr_data[45], w_hssi_10g_rx_pcs_rx_fifo_wr_data[44], w_hssi_10g_rx_pcs_rx_fifo_wr_data[43], w_hssi_10g_rx_pcs_rx_fifo_wr_data[42], w_hssi_10g_rx_pcs_rx_fifo_wr_data[41], w_hssi_10g_rx_pcs_rx_fifo_wr_data[40], w_hssi_10g_rx_pcs_rx_fifo_wr_data[39], w_hssi_10g_rx_pcs_rx_fifo_wr_data[38], w_hssi_10g_rx_pcs_rx_fifo_wr_data[37], w_hssi_10g_rx_pcs_rx_fifo_wr_data[36], w_hssi_10g_rx_pcs_rx_fifo_wr_data[35], w_hssi_10g_rx_pcs_rx_fifo_wr_data[34], w_hssi_10g_rx_pcs_rx_fifo_wr_data[33], w_hssi_10g_rx_pcs_rx_fifo_wr_data[32], w_hssi_10g_rx_pcs_rx_fifo_wr_data[31], w_hssi_10g_rx_pcs_rx_fifo_wr_data[30], w_hssi_10g_rx_pcs_rx_fifo_wr_data[29], w_hssi_10g_rx_pcs_rx_fifo_wr_data[28], w_hssi_10g_rx_pcs_rx_fifo_wr_data[27], w_hssi_10g_rx_pcs_rx_fifo_wr_data[26], w_hssi_10g_rx_pcs_rx_fifo_wr_data[25], w_hssi_10g_rx_pcs_rx_fifo_wr_data[24], w_hssi_10g_rx_pcs_rx_fifo_wr_data[23], w_hssi_10g_rx_pcs_rx_fifo_wr_data[22], w_hssi_10g_rx_pcs_rx_fifo_wr_data[21], w_hssi_10g_rx_pcs_rx_fifo_wr_data[20], w_hssi_10g_rx_pcs_rx_fifo_wr_data[19], w_hssi_10g_rx_pcs_rx_fifo_wr_data[18], w_hssi_10g_rx_pcs_rx_fifo_wr_data[17], w_hssi_10g_rx_pcs_rx_fifo_wr_data[16], w_hssi_10g_rx_pcs_rx_fifo_wr_data[15], w_hssi_10g_rx_pcs_rx_fifo_wr_data[14], w_hssi_10g_rx_pcs_rx_fifo_wr_data[13], w_hssi_10g_rx_pcs_rx_fifo_wr_data[12], w_hssi_10g_rx_pcs_rx_fifo_wr_data[11], w_hssi_10g_rx_pcs_rx_fifo_wr_data[10], w_hssi_10g_rx_pcs_rx_fifo_wr_data[9], w_hssi_10g_rx_pcs_rx_fifo_wr_data[8], w_hssi_10g_rx_pcs_rx_fifo_wr_data[7], w_hssi_10g_rx_pcs_rx_fifo_wr_data[6], w_hssi_10g_rx_pcs_rx_fifo_wr_data[5], w_hssi_10g_rx_pcs_rx_fifo_wr_data[4], w_hssi_10g_rx_pcs_rx_fifo_wr_data[3], w_hssi_10g_rx_pcs_rx_fifo_wr_data[2], w_hssi_10g_rx_pcs_rx_fifo_wr_data[1], w_hssi_10g_rx_pcs_rx_fifo_wr_data[0]}),
				.data_in_8g_clock_comp({w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0]}),
				.data_in_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr2_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0]}),
				.rd_ptr2_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0]}),
				.rd_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0]}),
				.rd_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.wr_clk_8g_clock_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_8g_clock_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.wr_en_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.wr_en_8g_clock_comp(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_en_8g_phase_comp(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.wr_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0]}),
				.wr_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0]}),
				.wr_rst_n_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.wr_rst_n_8g_clock_comp(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_n_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_rx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79:0] = 80'b0;
				assign w_hssi_fifo_rx_pcs_data_out_gen3[39:0] = 40'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_tx_pcs
			twentynm_hssi_fifo_tx_pcs #(
				.double_write_mode(hssi_fifo_tx_pcs_double_write_mode),
				.prot_mode(hssi_fifo_tx_pcs_prot_mode),
				.silicon_rev( "20nm5es" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_tx_pcs_blockselect),
				.data_out_10g(w_hssi_fifo_tx_pcs_data_out_10g),
				.data_out_8g_phase_comp(w_hssi_fifo_tx_pcs_data_out_8g_phase_comp),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in2_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0]}),
				.data_in_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_en_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.wr_en_8g_phase_comp(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0]}),
				.wr_rst_n_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_tx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_tx_pcs_data_out_10g[72:0] = 73'b0;
				assign w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63:0] = 64'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_rx_pcs
			twentynm_hssi_gen3_rx_pcs #(
				.block_sync(hssi_gen3_rx_pcs_block_sync),
				.block_sync_sm(hssi_gen3_rx_pcs_block_sync_sm),
				.cdr_ctrl_force_unalgn(hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn),
				.lpbk_force(hssi_gen3_rx_pcs_lpbk_force),
				.mode(hssi_gen3_rx_pcs_mode),
				.rate_match_fifo(hssi_gen3_rx_pcs_rate_match_fifo),
				.rate_match_fifo_latency(hssi_gen3_rx_pcs_rate_match_fifo_latency),
				.reconfig_settings(hssi_gen3_rx_pcs_reconfig_settings),
				.reverse_lpbk(hssi_gen3_rx_pcs_reverse_lpbk),
				.rx_b4gb_par_lpbk(hssi_gen3_rx_pcs_rx_b4gb_par_lpbk),
				.rx_force_balign(hssi_gen3_rx_pcs_rx_force_balign),
				.rx_ins_del_one_skip(hssi_gen3_rx_pcs_rx_ins_del_one_skip),
				.rx_num_fixed_pat(hssi_gen3_rx_pcs_rx_num_fixed_pat),
				.rx_test_out_sel(hssi_gen3_rx_pcs_rx_test_out_sel),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_rx_pcs_sup_mode)
			) inst_twentynm_hssi_gen3_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_rx_pcs_avmmreaddata),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.blk_start(w_hssi_gen3_rx_pcs_blk_start),
				.blockselect(w_hssi_gen3_rx_pcs_blockselect),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.data_out(w_hssi_gen3_rx_pcs_data_out),
				.data_valid(w_hssi_gen3_rx_pcs_data_valid),
				.ei_det_int(w_hssi_gen3_rx_pcs_ei_det_int),
				.ei_partial_det_int(w_hssi_gen3_rx_pcs_ei_partial_det_int),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.i_det_int(w_hssi_gen3_rx_pcs_i_det_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data(w_hssi_gen3_rx_pcs_lpbk_data),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.mem_rx_fifo_rd_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr),
				.mem_rx_fifo_wr_clk(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.mem_rx_fifo_wr_data(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data),
				.mem_rx_fifo_wr_en(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.mem_rx_fifo_wr_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr),
				.mem_rx_fifo_wr_rst_n(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_test_out(w_hssi_gen3_rx_pcs_rx_test_out),
				.sync_hdr(w_hssi_gen3_rx_pcs_sync_hdr),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0]}),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.mem_rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_gen3[39], w_hssi_fifo_rx_pcs_data_out_gen3[38], w_hssi_fifo_rx_pcs_data_out_gen3[37], w_hssi_fifo_rx_pcs_data_out_gen3[36], w_hssi_fifo_rx_pcs_data_out_gen3[35], w_hssi_fifo_rx_pcs_data_out_gen3[34], w_hssi_fifo_rx_pcs_data_out_gen3[33], w_hssi_fifo_rx_pcs_data_out_gen3[32], w_hssi_fifo_rx_pcs_data_out_gen3[31], w_hssi_fifo_rx_pcs_data_out_gen3[30], w_hssi_fifo_rx_pcs_data_out_gen3[29], w_hssi_fifo_rx_pcs_data_out_gen3[28], w_hssi_fifo_rx_pcs_data_out_gen3[27], w_hssi_fifo_rx_pcs_data_out_gen3[26], w_hssi_fifo_rx_pcs_data_out_gen3[25], w_hssi_fifo_rx_pcs_data_out_gen3[24], w_hssi_fifo_rx_pcs_data_out_gen3[23], w_hssi_fifo_rx_pcs_data_out_gen3[22], w_hssi_fifo_rx_pcs_data_out_gen3[21], w_hssi_fifo_rx_pcs_data_out_gen3[20], w_hssi_fifo_rx_pcs_data_out_gen3[19], w_hssi_fifo_rx_pcs_data_out_gen3[18], w_hssi_fifo_rx_pcs_data_out_gen3[17], w_hssi_fifo_rx_pcs_data_out_gen3[16], w_hssi_fifo_rx_pcs_data_out_gen3[15], w_hssi_fifo_rx_pcs_data_out_gen3[14], w_hssi_fifo_rx_pcs_data_out_gen3[13], w_hssi_fifo_rx_pcs_data_out_gen3[12], w_hssi_fifo_rx_pcs_data_out_gen3[11], w_hssi_fifo_rx_pcs_data_out_gen3[10], w_hssi_fifo_rx_pcs_data_out_gen3[9], w_hssi_fifo_rx_pcs_data_out_gen3[8], w_hssi_fifo_rx_pcs_data_out_gen3[7], w_hssi_fifo_rx_pcs_data_out_gen3[6], w_hssi_fifo_rx_pcs_data_out_gen3[5], w_hssi_fifo_rx_pcs_data_out_gen3[4], w_hssi_fifo_rx_pcs_data_out_gen3[3], w_hssi_fifo_rx_pcs_data_out_gen3[2], w_hssi_fifo_rx_pcs_data_out_gen3[1], w_hssi_fifo_rx_pcs_data_out_gen3[0]}),
				.par_lpbk_b4gb_in({w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0]}),
				.par_lpbk_in({w_hssi_gen3_tx_pcs_par_lpbk_out[31], w_hssi_gen3_tx_pcs_par_lpbk_out[30], w_hssi_gen3_tx_pcs_par_lpbk_out[29], w_hssi_gen3_tx_pcs_par_lpbk_out[28], w_hssi_gen3_tx_pcs_par_lpbk_out[27], w_hssi_gen3_tx_pcs_par_lpbk_out[26], w_hssi_gen3_tx_pcs_par_lpbk_out[25], w_hssi_gen3_tx_pcs_par_lpbk_out[24], w_hssi_gen3_tx_pcs_par_lpbk_out[23], w_hssi_gen3_tx_pcs_par_lpbk_out[22], w_hssi_gen3_tx_pcs_par_lpbk_out[21], w_hssi_gen3_tx_pcs_par_lpbk_out[20], w_hssi_gen3_tx_pcs_par_lpbk_out[19], w_hssi_gen3_tx_pcs_par_lpbk_out[18], w_hssi_gen3_tx_pcs_par_lpbk_out[17], w_hssi_gen3_tx_pcs_par_lpbk_out[16], w_hssi_gen3_tx_pcs_par_lpbk_out[15], w_hssi_gen3_tx_pcs_par_lpbk_out[14], w_hssi_gen3_tx_pcs_par_lpbk_out[13], w_hssi_gen3_tx_pcs_par_lpbk_out[12], w_hssi_gen3_tx_pcs_par_lpbk_out[11], w_hssi_gen3_tx_pcs_par_lpbk_out[10], w_hssi_gen3_tx_pcs_par_lpbk_out[9], w_hssi_gen3_tx_pcs_par_lpbk_out[8], w_hssi_gen3_tx_pcs_par_lpbk_out[7], w_hssi_gen3_tx_pcs_par_lpbk_out[6], w_hssi_gen3_tx_pcs_par_lpbk_out[5], w_hssi_gen3_tx_pcs_par_lpbk_out[4], w_hssi_gen3_tx_pcs_par_lpbk_out[3], w_hssi_gen3_tx_pcs_par_lpbk_out[2], w_hssi_gen3_tx_pcs_par_lpbk_out[1], w_hssi_gen3_tx_pcs_par_lpbk_out[0]}),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.rcvd_clk(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_pma_clk(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.rxpolarity(w_hssi_pipe_gen3_rxpolarity_int),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.sync_sm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.txdatak_in({w_hssi_pipe_gen3_txdatak_int[3], w_hssi_pipe_gen3_txdatak_int[2], w_hssi_pipe_gen3_txdatak_int[1], w_hssi_pipe_gen3_txdatak_int[0]}),
				
				// UNUSED
				.blk_lockd_int(),
				.skp_det_int()
			);
		end // if generate
		else begin
				assign w_hssi_gen3_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_rx_pcs_blk_algnd_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_delete_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_insert_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_overfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_undfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_rx_pcs_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_partial_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_err_decode_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_i_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data[33:0] = 34'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39:0] = 40'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_rx_test_out[19:0] = 20'b0;
				assign w_hssi_gen3_rx_pcs_sync_hdr[1:0] = 2'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_tx_pcs
			twentynm_hssi_gen3_tx_pcs #(
				.mode(hssi_gen3_tx_pcs_mode),
				.reverse_lpbk(hssi_gen3_tx_pcs_reverse_lpbk),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_tx_pcs_sup_mode),
				.tx_bitslip(hssi_gen3_tx_pcs_tx_bitslip),
				.tx_gbox_byp(hssi_gen3_tx_pcs_tx_gbox_byp)
			) inst_twentynm_hssi_gen3_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_gen3_tx_pcs_blockselect),
				.data_out(w_hssi_gen3_tx_pcs_data_out),
				.par_lpbk_b4gb_out(w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out),
				.par_lpbk_out(w_hssi_gen3_tx_pcs_par_lpbk_out),
				.tx_test_out(w_hssi_gen3_tx_pcs_tx_test_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_start_in(w_hssi_pipe_gen3_tx_blk_start_int),
				.data_in({w_hssi_pipe_gen3_txdata_int[31], w_hssi_pipe_gen3_txdata_int[30], w_hssi_pipe_gen3_txdata_int[29], w_hssi_pipe_gen3_txdata_int[28], w_hssi_pipe_gen3_txdata_int[27], w_hssi_pipe_gen3_txdata_int[26], w_hssi_pipe_gen3_txdata_int[25], w_hssi_pipe_gen3_txdata_int[24], w_hssi_pipe_gen3_txdata_int[23], w_hssi_pipe_gen3_txdata_int[22], w_hssi_pipe_gen3_txdata_int[21], w_hssi_pipe_gen3_txdata_int[20], w_hssi_pipe_gen3_txdata_int[19], w_hssi_pipe_gen3_txdata_int[18], w_hssi_pipe_gen3_txdata_int[17], w_hssi_pipe_gen3_txdata_int[16], w_hssi_pipe_gen3_txdata_int[15], w_hssi_pipe_gen3_txdata_int[14], w_hssi_pipe_gen3_txdata_int[13], w_hssi_pipe_gen3_txdata_int[12], w_hssi_pipe_gen3_txdata_int[11], w_hssi_pipe_gen3_txdata_int[10], w_hssi_pipe_gen3_txdata_int[9], w_hssi_pipe_gen3_txdata_int[8], w_hssi_pipe_gen3_txdata_int[7], w_hssi_pipe_gen3_txdata_int[6], w_hssi_pipe_gen3_txdata_int[5], w_hssi_pipe_gen3_txdata_int[4], w_hssi_pipe_gen3_txdata_int[3], w_hssi_pipe_gen3_txdata_int[2], w_hssi_pipe_gen3_txdata_int[1], w_hssi_pipe_gen3_txdata_int[0]}),
				.data_valid(w_hssi_pipe_gen3_txdataskip_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data_in({w_hssi_gen3_rx_pcs_lpbk_data[33], w_hssi_gen3_rx_pcs_lpbk_data[32], w_hssi_gen3_rx_pcs_lpbk_data[31], w_hssi_gen3_rx_pcs_lpbk_data[30], w_hssi_gen3_rx_pcs_lpbk_data[29], w_hssi_gen3_rx_pcs_lpbk_data[28], w_hssi_gen3_rx_pcs_lpbk_data[27], w_hssi_gen3_rx_pcs_lpbk_data[26], w_hssi_gen3_rx_pcs_lpbk_data[25], w_hssi_gen3_rx_pcs_lpbk_data[24], w_hssi_gen3_rx_pcs_lpbk_data[23], w_hssi_gen3_rx_pcs_lpbk_data[22], w_hssi_gen3_rx_pcs_lpbk_data[21], w_hssi_gen3_rx_pcs_lpbk_data[20], w_hssi_gen3_rx_pcs_lpbk_data[19], w_hssi_gen3_rx_pcs_lpbk_data[18], w_hssi_gen3_rx_pcs_lpbk_data[17], w_hssi_gen3_rx_pcs_lpbk_data[16], w_hssi_gen3_rx_pcs_lpbk_data[15], w_hssi_gen3_rx_pcs_lpbk_data[14], w_hssi_gen3_rx_pcs_lpbk_data[13], w_hssi_gen3_rx_pcs_lpbk_data[12], w_hssi_gen3_rx_pcs_lpbk_data[11], w_hssi_gen3_rx_pcs_lpbk_data[10], w_hssi_gen3_rx_pcs_lpbk_data[9], w_hssi_gen3_rx_pcs_lpbk_data[8], w_hssi_gen3_rx_pcs_lpbk_data[7], w_hssi_gen3_rx_pcs_lpbk_data[6], w_hssi_gen3_rx_pcs_lpbk_data[5], w_hssi_gen3_rx_pcs_lpbk_data[4], w_hssi_gen3_rx_pcs_lpbk_data[3], w_hssi_gen3_rx_pcs_lpbk_data[2], w_hssi_gen3_rx_pcs_lpbk_data[1], w_hssi_gen3_rx_pcs_lpbk_data[0]}),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.sync_in({w_hssi_pipe_gen3_tx_sync_hdr_int[1], w_hssi_pipe_gen3_tx_sync_hdr_int[0]}),
				.tx_pma_clk(w_hssi_8g_tx_pcs_clk_out_gen3),
				.tx_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn)
			);
		end // if generate
		else begin
				assign w_hssi_gen3_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_tx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_tx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35:0] = 36'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_tx_test_out[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_rx_pcs
			twentynm_hssi_krfec_rx_pcs #(
				.blksync_cor_en(hssi_krfec_rx_pcs_blksync_cor_en),
				.bypass_gb(hssi_krfec_rx_pcs_bypass_gb),
				.clr_ctrl(hssi_krfec_rx_pcs_clr_ctrl),
				.ctrl_bit_reverse(hssi_krfec_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_rx_pcs_data_bit_reverse),
				.dv_start(hssi_krfec_rx_pcs_dv_start),
				.err_mark_type(hssi_krfec_rx_pcs_err_mark_type),
				.error_marking_en(hssi_krfec_rx_pcs_error_marking_en),
				.low_latency_en(hssi_krfec_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_krfec_rx_pcs_lpbk_mode),
				.parity_invalid_enum(hssi_krfec_rx_pcs_parity_invalid_enum),
				.parity_valid_num(hssi_krfec_rx_pcs_parity_valid_num),
				.pipeln_blksync(hssi_krfec_rx_pcs_pipeln_blksync),
				.pipeln_descrm(hssi_krfec_rx_pcs_pipeln_descrm),
				.pipeln_errcorrect(hssi_krfec_rx_pcs_pipeln_errcorrect),
				.pipeln_errtrap_ind(hssi_krfec_rx_pcs_pipeln_errtrap_ind),
				.pipeln_errtrap_lfsr(hssi_krfec_rx_pcs_pipeln_errtrap_lfsr),
				.pipeln_errtrap_loc(hssi_krfec_rx_pcs_pipeln_errtrap_loc),
				.pipeln_errtrap_pat(hssi_krfec_rx_pcs_pipeln_errtrap_pat),
				.pipeln_gearbox(hssi_krfec_rx_pcs_pipeln_gearbox),
				.pipeln_syndrm(hssi_krfec_rx_pcs_pipeln_syndrm),
				.pipeln_trans_dec(hssi_krfec_rx_pcs_pipeln_trans_dec),
				.prot_mode(hssi_krfec_rx_pcs_prot_mode),
				.receive_order(hssi_krfec_rx_pcs_receive_order),
				.reconfig_settings(hssi_krfec_rx_pcs_reconfig_settings),
				.rx_testbus_sel(hssi_krfec_rx_pcs_rx_testbus_sel),
				.signal_ok_en(hssi_krfec_rx_pcs_signal_ok_en),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_rx_pcs_sup_mode)
			) inst_twentynm_hssi_krfec_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_rx_pcs_blockselect),
				.rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.rx_control_out(w_hssi_krfec_rx_pcs_rx_control_out),
				.rx_data_out(w_hssi_krfec_rx_pcs_rx_data_out),
				.rx_data_status(w_hssi_krfec_rx_pcs_rx_data_status),
				.rx_data_valid_out(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.rx_signal_ok_out(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.rx_data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0]}),
				.rx_krfec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_krfec_reg(),
				.pld_10g_krfec_rx_blk_lock_krfec_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg(),
				.pld_10g_krfec_rx_frame_krfec_reg(),
				.pld_10g_krfec_rx_frame_krfec_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_rx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_block_lock = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_control_out[9:0] = 10'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_status[1:0] = 2'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_valid_out = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_frame = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_signal_ok_out = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_tx_pcs
			twentynm_hssi_krfec_tx_pcs #(
				.burst_err(hssi_krfec_tx_pcs_burst_err),
				.burst_err_len(hssi_krfec_tx_pcs_burst_err_len),
				.ctrl_bit_reverse(hssi_krfec_tx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_tx_pcs_data_bit_reverse),
				.enc_frame_query(hssi_krfec_tx_pcs_enc_frame_query),
				.low_latency_en(hssi_krfec_tx_pcs_low_latency_en),
				.pipeln_encoder(hssi_krfec_tx_pcs_pipeln_encoder),
				.pipeln_scrambler(hssi_krfec_tx_pcs_pipeln_scrambler),
				.prot_mode(hssi_krfec_tx_pcs_prot_mode),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_tx_pcs_sup_mode),
				.transcode_err(hssi_krfec_tx_pcs_transcode_err),
				.transmit_order(hssi_krfec_tx_pcs_transmit_order),
				.tx_testbus_sel(hssi_krfec_tx_pcs_tx_testbus_sel)
			) inst_twentynm_hssi_krfec_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_tx_pcs_blockselect),
				.tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.tx_data_out(w_hssi_krfec_tx_pcs_tx_data_out),
				.tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.tx_test_data(w_hssi_krfec_tx_pcs_tx_test_data),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.tx_control_in({w_hssi_10g_tx_pcs_tx_control_out_krfec[8], w_hssi_10g_tx_pcs_tx_control_out_krfec[7], w_hssi_10g_tx_pcs_tx_control_out_krfec[6], w_hssi_10g_tx_pcs_tx_control_out_krfec[5], w_hssi_10g_tx_pcs_tx_control_out_krfec[4], w_hssi_10g_tx_pcs_tx_control_out_krfec[3], w_hssi_10g_tx_pcs_tx_control_out_krfec[2], w_hssi_10g_tx_pcs_tx_control_out_krfec[1], w_hssi_10g_tx_pcs_tx_control_out_krfec[0]}),
				.tx_data_in({w_hssi_10g_tx_pcs_tx_data_out_krfec[63], w_hssi_10g_tx_pcs_tx_data_out_krfec[62], w_hssi_10g_tx_pcs_tx_data_out_krfec[61], w_hssi_10g_tx_pcs_tx_data_out_krfec[60], w_hssi_10g_tx_pcs_tx_data_out_krfec[59], w_hssi_10g_tx_pcs_tx_data_out_krfec[58], w_hssi_10g_tx_pcs_tx_data_out_krfec[57], w_hssi_10g_tx_pcs_tx_data_out_krfec[56], w_hssi_10g_tx_pcs_tx_data_out_krfec[55], w_hssi_10g_tx_pcs_tx_data_out_krfec[54], w_hssi_10g_tx_pcs_tx_data_out_krfec[53], w_hssi_10g_tx_pcs_tx_data_out_krfec[52], w_hssi_10g_tx_pcs_tx_data_out_krfec[51], w_hssi_10g_tx_pcs_tx_data_out_krfec[50], w_hssi_10g_tx_pcs_tx_data_out_krfec[49], w_hssi_10g_tx_pcs_tx_data_out_krfec[48], w_hssi_10g_tx_pcs_tx_data_out_krfec[47], w_hssi_10g_tx_pcs_tx_data_out_krfec[46], w_hssi_10g_tx_pcs_tx_data_out_krfec[45], w_hssi_10g_tx_pcs_tx_data_out_krfec[44], w_hssi_10g_tx_pcs_tx_data_out_krfec[43], w_hssi_10g_tx_pcs_tx_data_out_krfec[42], w_hssi_10g_tx_pcs_tx_data_out_krfec[41], w_hssi_10g_tx_pcs_tx_data_out_krfec[40], w_hssi_10g_tx_pcs_tx_data_out_krfec[39], w_hssi_10g_tx_pcs_tx_data_out_krfec[38], w_hssi_10g_tx_pcs_tx_data_out_krfec[37], w_hssi_10g_tx_pcs_tx_data_out_krfec[36], w_hssi_10g_tx_pcs_tx_data_out_krfec[35], w_hssi_10g_tx_pcs_tx_data_out_krfec[34], w_hssi_10g_tx_pcs_tx_data_out_krfec[33], w_hssi_10g_tx_pcs_tx_data_out_krfec[32], w_hssi_10g_tx_pcs_tx_data_out_krfec[31], w_hssi_10g_tx_pcs_tx_data_out_krfec[30], w_hssi_10g_tx_pcs_tx_data_out_krfec[29], w_hssi_10g_tx_pcs_tx_data_out_krfec[28], w_hssi_10g_tx_pcs_tx_data_out_krfec[27], w_hssi_10g_tx_pcs_tx_data_out_krfec[26], w_hssi_10g_tx_pcs_tx_data_out_krfec[25], w_hssi_10g_tx_pcs_tx_data_out_krfec[24], w_hssi_10g_tx_pcs_tx_data_out_krfec[23], w_hssi_10g_tx_pcs_tx_data_out_krfec[22], w_hssi_10g_tx_pcs_tx_data_out_krfec[21], w_hssi_10g_tx_pcs_tx_data_out_krfec[20], w_hssi_10g_tx_pcs_tx_data_out_krfec[19], w_hssi_10g_tx_pcs_tx_data_out_krfec[18], w_hssi_10g_tx_pcs_tx_data_out_krfec[17], w_hssi_10g_tx_pcs_tx_data_out_krfec[16], w_hssi_10g_tx_pcs_tx_data_out_krfec[15], w_hssi_10g_tx_pcs_tx_data_out_krfec[14], w_hssi_10g_tx_pcs_tx_data_out_krfec[13], w_hssi_10g_tx_pcs_tx_data_out_krfec[12], w_hssi_10g_tx_pcs_tx_data_out_krfec[11], w_hssi_10g_tx_pcs_tx_data_out_krfec[10], w_hssi_10g_tx_pcs_tx_data_out_krfec[9], w_hssi_10g_tx_pcs_tx_data_out_krfec[8], w_hssi_10g_tx_pcs_tx_data_out_krfec[7], w_hssi_10g_tx_pcs_tx_data_out_krfec[6], w_hssi_10g_tx_pcs_tx_data_out_krfec[5], w_hssi_10g_tx_pcs_tx_data_out_krfec[4], w_hssi_10g_tx_pcs_tx_data_out_krfec[3], w_hssi_10g_tx_pcs_tx_data_out_krfec[2], w_hssi_10g_tx_pcs_tx_data_out_krfec[1], w_hssi_10g_tx_pcs_tx_data_out_krfec[0]}),
				.tx_data_valid_in(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_krfec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_krfec_reg(),
				.pld_krfec_tx_alignment_plddirect_reg(),
				.pld_krfec_tx_alignment_reg()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_tx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_alignment = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_test_data[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen1_2
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen1_2
			twentynm_hssi_pipe_gen1_2 #(
				.elec_idle_delay_val(hssi_pipe_gen1_2_elec_idle_delay_val),
				.error_replace_pad(hssi_pipe_gen1_2_error_replace_pad),
				.hip_mode(hssi_pipe_gen1_2_hip_mode),
				.ind_error_reporting(hssi_pipe_gen1_2_ind_error_reporting),
				.phystatus_delay_val(hssi_pipe_gen1_2_phystatus_delay_val),
				.phystatus_rst_toggle(hssi_pipe_gen1_2_phystatus_rst_toggle),
				.pipe_byte_de_serializer_en(hssi_pipe_gen1_2_pipe_byte_de_serializer_en),
				.prot_mode(hssi_pipe_gen1_2_prot_mode),
				.reconfig_settings(hssi_pipe_gen1_2_reconfig_settings),
				.rx_pipe_enable(hssi_pipe_gen1_2_rx_pipe_enable),
				.rxdetect_bypass(hssi_pipe_gen1_2_rxdetect_bypass),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen1_2_sup_mode),
				.tx_pipe_enable(hssi_pipe_gen1_2_tx_pipe_enable),
				.txswing(hssi_pipe_gen1_2_txswing)
			) inst_twentynm_hssi_pipe_gen1_2 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen1_2_avmmreaddata),
				.blockselect(w_hssi_pipe_gen1_2_blockselect),
				.current_coeff(w_hssi_pipe_gen1_2_current_coeff),
				.phystatus(w_hssi_pipe_gen1_2_phystatus),
				.polarity_inversion_rx(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rev_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.rxelectricalidle_out(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxstatus(w_hssi_pipe_gen1_2_rxstatus),
				.rxvalid(w_hssi_pipe_gen1_2_rxvalid),
				.tx_elec_idle_out(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pipe_rx_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.power_state_transition_done_ena(1'b0),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rev_loopbk_pcs_gen3(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.revloopback(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.rx_pipe_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rxd({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxelectricalidle(w_hssi_8g_rx_pcs_eidle_detected),
				.rxelectricalidle_pcs_gen3(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.rxpolarity_pcs_gen3(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.tx_elec_idle_comp(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.txd_ch({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswingport(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.pld_8g_rxpolarity_pipe3_reg(),
				.rxd_ch(),
				.txd()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen1_2_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen1_2_blockselect = 1'b0;
				assign w_hssi_pipe_gen1_2_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen1_2_phystatus = 1'b0;
				assign w_hssi_pipe_gen1_2_polarity_inversion_rx = 1'b0;
				assign w_hssi_pipe_gen1_2_rev_loopbk = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelectricalidle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen1_2_rxvalid = 1'b0;
				assign w_hssi_pipe_gen1_2_tx_elec_idle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_txdetectrx = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen3
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen3
			twentynm_hssi_pipe_gen3 #(
				.bypass_rx_detection_enable(hssi_pipe_gen3_bypass_rx_detection_enable),
				.bypass_rx_preset(hssi_pipe_gen3_bypass_rx_preset),
				.bypass_rx_preset_enable(hssi_pipe_gen3_bypass_rx_preset_enable),
				.bypass_tx_coefficent(hssi_pipe_gen3_bypass_tx_coefficent),
				.bypass_tx_coefficent_enable(hssi_pipe_gen3_bypass_tx_coefficent_enable),
				.elecidle_delay_g3(hssi_pipe_gen3_elecidle_delay_g3),
				.ind_error_reporting(hssi_pipe_gen3_ind_error_reporting),
				.mode(hssi_pipe_gen3_mode),
				.phy_status_delay_g12(hssi_pipe_gen3_phy_status_delay_g12),
				.phy_status_delay_g3(hssi_pipe_gen3_phy_status_delay_g3),
				.phystatus_rst_toggle_g12(hssi_pipe_gen3_phystatus_rst_toggle_g12),
				.phystatus_rst_toggle_g3(hssi_pipe_gen3_phystatus_rst_toggle_g3),
				.rate_match_pad_insertion(hssi_pipe_gen3_rate_match_pad_insertion),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen3_sup_mode),
				.test_out_sel(hssi_pipe_gen3_test_out_sel)
			) inst_twentynm_hssi_pipe_gen3 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen3_avmmreaddata),
				.blockselect(w_hssi_pipe_gen3_blockselect),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.phystatus(w_hssi_pipe_gen3_phystatus),
				.pma_current_coeff(w_hssi_pipe_gen3_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_pipe_gen3_pma_current_rxpreset),
				.pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.rev_lpbk_8gpcs_out(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.rev_lpbk_int(w_hssi_pipe_gen3_rev_lpbk_int),
				.rx_blk_start(w_hssi_pipe_gen3_rx_blk_start),
				.rx_sync_hdr(w_hssi_pipe_gen3_rx_sync_hdr),
				.rxd_8gpcs_out(w_hssi_pipe_gen3_rxd_8gpcs_out),
				.rxdataskip(w_hssi_pipe_gen3_rxdataskip),
				.rxelecidle(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity_8gpcs_out(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.rxpolarity_int(w_hssi_pipe_gen3_rxpolarity_int),
				.rxstatus(w_hssi_pipe_gen3_rxstatus),
				.rxvalid(w_hssi_pipe_gen3_rxvalid),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.test_out(w_hssi_pipe_gen3_test_out),
				.tx_blk_start_int(w_hssi_pipe_gen3_tx_blk_start_int),
				.tx_sync_hdr_int(w_hssi_pipe_gen3_tx_sync_hdr_int),
				.txdata_int(w_hssi_pipe_gen3_txdata_int),
				.txdatak_int(w_hssi_pipe_gen3_txdatak_int),
				.txdataskip_int(w_hssi_pipe_gen3_txdataskip_int),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.current_coeff({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0]}),
				.current_rxpreset({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0]}),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.pcs_asn_bundling_in({w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0]}),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pipe_tx_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_blk_start_int(w_hssi_gen3_rx_pcs_blk_start),
				.rx_sync_hdr_int({w_hssi_gen3_rx_pcs_sync_hdr[1], w_hssi_gen3_rx_pcs_sync_hdr[0]}),
				.rx_test_out({w_hssi_gen3_rx_pcs_rx_test_out[19], w_hssi_gen3_rx_pcs_rx_test_out[18], w_hssi_gen3_rx_pcs_rx_test_out[17], w_hssi_gen3_rx_pcs_rx_test_out[16], w_hssi_gen3_rx_pcs_rx_test_out[15], w_hssi_gen3_rx_pcs_rx_test_out[14], w_hssi_gen3_rx_pcs_rx_test_out[13], w_hssi_gen3_rx_pcs_rx_test_out[12], w_hssi_gen3_rx_pcs_rx_test_out[11], w_hssi_gen3_rx_pcs_rx_test_out[10], w_hssi_gen3_rx_pcs_rx_test_out[9], w_hssi_gen3_rx_pcs_rx_test_out[8], w_hssi_gen3_rx_pcs_rx_test_out[7], w_hssi_gen3_rx_pcs_rx_test_out[6], w_hssi_gen3_rx_pcs_rx_test_out[5], w_hssi_gen3_rx_pcs_rx_test_out[4], w_hssi_gen3_rx_pcs_rx_test_out[3], w_hssi_gen3_rx_pcs_rx_test_out[2], w_hssi_gen3_rx_pcs_rx_test_out[1], w_hssi_gen3_rx_pcs_rx_test_out[0]}),
				.rxd_8gpcs_in({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxdata_int({w_hssi_gen3_rx_pcs_data_out[31], w_hssi_gen3_rx_pcs_data_out[30], w_hssi_gen3_rx_pcs_data_out[29], w_hssi_gen3_rx_pcs_data_out[28], w_hssi_gen3_rx_pcs_data_out[27], w_hssi_gen3_rx_pcs_data_out[26], w_hssi_gen3_rx_pcs_data_out[25], w_hssi_gen3_rx_pcs_data_out[24], w_hssi_gen3_rx_pcs_data_out[23], w_hssi_gen3_rx_pcs_data_out[22], w_hssi_gen3_rx_pcs_data_out[21], w_hssi_gen3_rx_pcs_data_out[20], w_hssi_gen3_rx_pcs_data_out[19], w_hssi_gen3_rx_pcs_data_out[18], w_hssi_gen3_rx_pcs_data_out[17], w_hssi_gen3_rx_pcs_data_out[16], w_hssi_gen3_rx_pcs_data_out[15], w_hssi_gen3_rx_pcs_data_out[14], w_hssi_gen3_rx_pcs_data_out[13], w_hssi_gen3_rx_pcs_data_out[12], w_hssi_gen3_rx_pcs_data_out[11], w_hssi_gen3_rx_pcs_data_out[10], w_hssi_gen3_rx_pcs_data_out[9], w_hssi_gen3_rx_pcs_data_out[8], w_hssi_gen3_rx_pcs_data_out[7], w_hssi_gen3_rx_pcs_data_out[6], w_hssi_gen3_rx_pcs_data_out[5], w_hssi_gen3_rx_pcs_data_out[4], w_hssi_gen3_rx_pcs_data_out[3], w_hssi_gen3_rx_pcs_data_out[2], w_hssi_gen3_rx_pcs_data_out[1], w_hssi_gen3_rx_pcs_data_out[0]}),
				.rxdatak_int({1'b0, 1'b0, 1'b0, 1'b0}),
				.rxdataskip_int(w_hssi_gen3_rx_pcs_data_valid),
				.rxelecidle_8gpcs_in(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.tx_blk_start(w_hssi_8g_tx_pcs_tx_blk_start_out[0]),
				.tx_sync_hdr({w_hssi_8g_tx_pcs_tx_sync_hdr_out[1], w_hssi_8g_tx_pcs_tx_sync_hdr_out[0]}),
				.tx_test_out({w_hssi_gen3_tx_pcs_tx_test_out[19], w_hssi_gen3_tx_pcs_tx_test_out[18], w_hssi_gen3_tx_pcs_tx_test_out[17], w_hssi_gen3_tx_pcs_tx_test_out[16], w_hssi_gen3_tx_pcs_tx_test_out[15], w_hssi_gen3_tx_pcs_tx_test_out[14], w_hssi_gen3_tx_pcs_tx_test_out[13], w_hssi_gen3_tx_pcs_tx_test_out[12], w_hssi_gen3_tx_pcs_tx_test_out[11], w_hssi_gen3_tx_pcs_tx_test_out[10], w_hssi_gen3_tx_pcs_tx_test_out[9], w_hssi_gen3_tx_pcs_tx_test_out[8], w_hssi_gen3_tx_pcs_tx_test_out[7], w_hssi_gen3_tx_pcs_tx_test_out[6], w_hssi_gen3_tx_pcs_tx_test_out[5], w_hssi_gen3_tx_pcs_tx_test_out[4], w_hssi_gen3_tx_pcs_tx_test_out[3], w_hssi_gen3_tx_pcs_tx_test_out[2], w_hssi_gen3_tx_pcs_tx_test_out[1], w_hssi_gen3_tx_pcs_tx_test_out[0]}),
				.txcompliance(w_hssi_8g_tx_pcs_txcompliance_out),
				.txdata({w_hssi_8g_tx_pcs_tx_data_out[31], w_hssi_8g_tx_pcs_tx_data_out[30], w_hssi_8g_tx_pcs_tx_data_out[29], w_hssi_8g_tx_pcs_tx_data_out[28], w_hssi_8g_tx_pcs_tx_data_out[27], w_hssi_8g_tx_pcs_tx_data_out[26], w_hssi_8g_tx_pcs_tx_data_out[25], w_hssi_8g_tx_pcs_tx_data_out[24], w_hssi_8g_tx_pcs_tx_data_out[23], w_hssi_8g_tx_pcs_tx_data_out[22], w_hssi_8g_tx_pcs_tx_data_out[21], w_hssi_8g_tx_pcs_tx_data_out[20], w_hssi_8g_tx_pcs_tx_data_out[19], w_hssi_8g_tx_pcs_tx_data_out[18], w_hssi_8g_tx_pcs_tx_data_out[17], w_hssi_8g_tx_pcs_tx_data_out[16], w_hssi_8g_tx_pcs_tx_data_out[15], w_hssi_8g_tx_pcs_tx_data_out[14], w_hssi_8g_tx_pcs_tx_data_out[13], w_hssi_8g_tx_pcs_tx_data_out[12], w_hssi_8g_tx_pcs_tx_data_out[11], w_hssi_8g_tx_pcs_tx_data_out[10], w_hssi_8g_tx_pcs_tx_data_out[9], w_hssi_8g_tx_pcs_tx_data_out[8], w_hssi_8g_tx_pcs_tx_data_out[7], w_hssi_8g_tx_pcs_tx_data_out[6], w_hssi_8g_tx_pcs_tx_data_out[5], w_hssi_8g_tx_pcs_tx_data_out[4], w_hssi_8g_tx_pcs_tx_data_out[3], w_hssi_8g_tx_pcs_tx_data_out[2], w_hssi_8g_tx_pcs_tx_data_out[1], w_hssi_8g_tx_pcs_tx_data_out[0]}),
				.txdatak({w_hssi_8g_tx_pcs_tx_datak_out[3], w_hssi_8g_tx_pcs_tx_datak_out[2], w_hssi_8g_tx_pcs_tx_datak_out[1], w_hssi_8g_tx_pcs_tx_datak_out[0]}),
				.txdataskip(w_hssi_8g_tx_pcs_tx_data_valid_out[0]),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_8g_tx_pcs_txelecidle_out),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.dis_pc_byte(),
				.pma_rx_det_pd(),
				.pma_txdeemph(),
				.pma_txmargin(),
				.pma_txswing(),
				.reset_pc_prts()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen3_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen3_blockselect = 1'b0;
				assign w_hssi_pipe_gen3_gen3_clk_sel = 1'b0;
				assign w_hssi_pipe_gen3_pcs_rst = 1'b0;
				assign w_hssi_pipe_gen3_phystatus = 1'b0;
				assign w_hssi_pipe_gen3_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen3_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_pma_tx_elec_idle = 1'b0;
				assign w_hssi_pipe_gen3_pma_txdetectrx = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_int = 1'b0;
				assign w_hssi_pipe_gen3_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_rxd_8gpcs_out[63:0] = 64'b0;
				assign w_hssi_pipe_gen3_rxdataskip[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_int = 1'b0;
				assign w_hssi_pipe_gen3_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_rxvalid = 1'b0;
				assign w_hssi_pipe_gen3_shutdown_clk = 1'b0;
				assign w_hssi_pipe_gen3_test_out[19:0] = 20'b0;
				assign w_hssi_pipe_gen3_tx_blk_start_int = 1'b0;
				assign w_hssi_pipe_gen3_tx_sync_hdr_int[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_txdata_int[31:0] = 32'b0;
				assign w_hssi_pipe_gen3_txdatak_int[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_txdataskip_int = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pcs_pma_interface
			twentynm_hssi_rx_pcs_pma_interface #(
				.block_sel(hssi_rx_pcs_pma_interface_block_sel),
				.channel_operation_mode(hssi_rx_pcs_pma_interface_channel_operation_mode),
				.clkslip_sel(hssi_rx_pcs_pma_interface_clkslip_sel),
				.lpbk_en(hssi_rx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_rx_pcs_pma_interface_master_clk_sel),
				.pldif_datawidth_mode(hssi_rx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_rx(hssi_rx_pcs_pma_interface_pma_dw_rx),
				.pma_if_dft_en(hssi_rx_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_rx_pcs_pma_interface_pma_if_dft_val),
				.prbs9_dwidth(hssi_rx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_rx_pcs_pma_interface_prbs_clken),
				.prbs_ver(hssi_rx_pcs_pma_interface_prbs_ver),
				.prot_mode_rx(hssi_rx_pcs_pma_interface_prot_mode_rx),
				.reconfig_settings(hssi_rx_pcs_pma_interface_reconfig_settings),
				.rx_dyn_polarity_inversion(hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion),
				.rx_lpbk_en(hssi_rx_pcs_pma_interface_rx_lpbk_en),
				.rx_prbs_force_signal_ok(hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok),
				.rx_prbs_mask(hssi_rx_pcs_pma_interface_rx_prbs_mask),
				.rx_prbs_mode(hssi_rx_pcs_pma_interface_rx_prbs_mode),
				.rx_signalok_signaldet_sel(hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel),
				.rx_static_polarity_inversion(hssi_rx_pcs_pma_interface_rx_static_polarity_inversion),
				.rx_uhsif_lpbk_en(hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sup_mode(hssi_rx_pcs_pma_interface_sup_mode)
			) inst_twentynm_hssi_rx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.int_pmaif_10g_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data),
				.int_pmaif_10g_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.int_pmaif_8g_pudi(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi),
				.int_pmaif_8g_rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.int_pmaif_8g_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.int_pmaif_8g_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.int_pmaif_8g_sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.int_pmaif_g3_pma_data_in(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in),
				.int_pmaif_g3_pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.int_pmaif_g3_pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.int_pmaif_g3_pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.int_pmaif_krfec_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data),
				.int_pmaif_krfec_rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.int_pmaif_pldif_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pmaif_pldif_prbs_err_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pmaif_pldif_rx_clkdiv(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pmaif_pldif_rx_clkdiv_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pmaif_pldif_rx_data(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data),
				.int_pmaif_pldif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pmaif_pldif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pmaif_pldif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pmaif_pldif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.pma_eye_monitor(w_hssi_rx_pcs_pma_interface_pma_eye_monitor),
				.pma_rx_clkslip(w_hssi_rx_pcs_pma_interface_pma_rx_clkslip),
				.pma_rxpma_rstb(w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb),
				.rx_pmaif_test_out(w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out),
				.rx_prbs_ver_test(w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.int_pmaif_8g_rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.int_pmaif_pldif_eye_monitor({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0]}),
				.int_pmaif_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pmaif_pldif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pmaif_pldif_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pmaif_pldif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pma_rx_clkdiv_user(in_pma_rx_clkdiv_user),
				.pma_rx_detect_valid(in_pma_rx_detect_valid),
				.pma_rx_found(in_pma_rx_found),
				.pma_rx_pma_clk(in_pma_rx_pma_clk),
				.pma_rx_pma_data({in_pma_rx_pma_data[63], in_pma_rx_pma_data[62], in_pma_rx_pma_data[61], in_pma_rx_pma_data[60], in_pma_rx_pma_data[59], in_pma_rx_pma_data[58], in_pma_rx_pma_data[57], in_pma_rx_pma_data[56], in_pma_rx_pma_data[55], in_pma_rx_pma_data[54], in_pma_rx_pma_data[53], in_pma_rx_pma_data[52], in_pma_rx_pma_data[51], in_pma_rx_pma_data[50], in_pma_rx_pma_data[49], in_pma_rx_pma_data[48], in_pma_rx_pma_data[47], in_pma_rx_pma_data[46], in_pma_rx_pma_data[45], in_pma_rx_pma_data[44], in_pma_rx_pma_data[43], in_pma_rx_pma_data[42], in_pma_rx_pma_data[41], in_pma_rx_pma_data[40], in_pma_rx_pma_data[39], in_pma_rx_pma_data[38], in_pma_rx_pma_data[37], in_pma_rx_pma_data[36], in_pma_rx_pma_data[35], in_pma_rx_pma_data[34], in_pma_rx_pma_data[33], in_pma_rx_pma_data[32], in_pma_rx_pma_data[31], in_pma_rx_pma_data[30], in_pma_rx_pma_data[29], in_pma_rx_pma_data[28], in_pma_rx_pma_data[27], in_pma_rx_pma_data[26], in_pma_rx_pma_data[25], in_pma_rx_pma_data[24], in_pma_rx_pma_data[23], in_pma_rx_pma_data[22], in_pma_rx_pma_data[21], in_pma_rx_pma_data[20], in_pma_rx_pma_data[19], in_pma_rx_pma_data[18], in_pma_rx_pma_data[17], in_pma_rx_pma_data[16], in_pma_rx_pma_data[15], in_pma_rx_pma_data[14], in_pma_rx_pma_data[13], in_pma_rx_pma_data[12], in_pma_rx_pma_data[11], in_pma_rx_pma_data[10], in_pma_rx_pma_data[9], in_pma_rx_pma_data[8], in_pma_rx_pma_data[7], in_pma_rx_pma_data[6], in_pma_rx_pma_data[5], in_pma_rx_pma_data[4], in_pma_rx_pma_data[3], in_pma_rx_pma_data[2], in_pma_rx_pma_data[1], in_pma_rx_pma_data[0]}),
				.pma_rx_signal_ok(in_pma_rx_signal_ok),
				.pma_rxpll_lock(in_pma_rxpll_lock),
				.pma_signal_det(in_pma_signal_det),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.tx_pma_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0]}),
				.tx_pma_uhsif_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0]}),
				
				// UNUSED
				.int_pmaif_g3_rcvd_clk(),
				.prbs_err_lt()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31:0] = 32'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5:0] = 6'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rx_clkslip = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pld_pcs_interface
			twentynm_hssi_rx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx),
				.hd_10g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx),
				.hd_10g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx),
				.hd_10g_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx),
				.hd_10g_lpbk_en(hssi_rx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx),
				.hd_10g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx),
				.hd_10g_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx),
				.hd_10g_test_bus_mode(hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode),
				.hd_8g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx),
				.hd_8g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx),
				.hd_8g_hip_mode(hssi_rx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_rx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx),
				.hd_8g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx),
				.hd_chnl_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_clklow_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz),
				.hd_chnl_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx),
				.hd_chnl_fref_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz),
				.hd_chnl_frequency_rules_en(hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_rx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_rx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx),
				.hd_chnl_lpbk_en(hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx),
				.hd_chnl_pld_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz),
				.hd_chnl_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx),
				.hd_chnl_pma_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz),
				.hd_chnl_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx),
				.hd_chnl_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx),
				.hd_chnl_transparent_pcs_rx(hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx),
				.hd_fifo_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx),
				.hd_fifo_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx),
				.hd_g3_prot_mode(hssi_rx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx),
				.hd_krfec_lpbk_en(hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx),
				.hd_krfec_test_bus_mode(hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode),
				.hd_pldif_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx),
				.hd_pmaif_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_lpbk_en(hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx),
				.hd_pmaif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx),
				.hd_pmaif_sim_mode(hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_rx_block_sel(hssi_rx_pld_pcs_interface_pcs_rx_block_sel),
				.pcs_rx_clk_out_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel),
				.pcs_rx_clk_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_sel),
				.pcs_rx_hip_clk_en(hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en),
				.pcs_rx_output_sel(hssi_rx_pld_pcs_interface_pcs_rx_output_sel),
				.reconfig_settings(hssi_rx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm5es" )       //PARAM_HIDE
			) inst_twentynm_hssi_rx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pld_pcs_interface_blockselect),
				.hip_rx_ctrl(w_hssi_rx_pld_pcs_interface_hip_rx_ctrl),
				.hip_rx_data(w_hssi_rx_pld_pcs_interface_hip_rx_data),
				.int_pldif_10g_rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.int_pldif_10g_rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.int_pldif_10g_rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.int_pldif_10g_rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.int_pldif_10g_rx_control_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb),
				.int_pldif_10g_rx_data_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb),
				.int_pldif_10g_rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.int_pldif_10g_rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.int_pldif_10g_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.int_pldif_10g_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.int_pldif_10g_rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.int_pldif_8g_a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.int_pldif_8g_bitloc_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.int_pldif_8g_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.int_pldif_8g_byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.int_pldif_8g_encdt(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.int_pldif_8g_pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.int_pldif_8g_rdenable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.int_pldif_8g_rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.int_pldif_8g_rxurstpcs_n(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.int_pldif_8g_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.int_pldif_8g_wrdisable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.int_pldif_g3_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.int_pldif_krfec_rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.int_pldif_pmaif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pldif_pmaif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pldif_pmaif_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pldif_pmaif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pld_10g_krfec_rx_blk_lock(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock),
				.pld_10g_krfec_rx_diag_data_status(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status),
				.pld_10g_krfec_rx_frame(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame),
				.pld_10g_rx_align_val(w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val),
				.pld_10g_rx_crc32_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err),
				.pld_10g_rx_data_valid(w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid),
				.pld_10g_rx_empty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty),
				.pld_10g_rx_fifo_del(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del),
				.pld_10g_rx_fifo_insert(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert),
				.pld_10g_rx_fifo_num(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num),
				.pld_10g_rx_frame_lock(w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock),
				.pld_10g_rx_hi_ber(w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber),
				.pld_10g_rx_oflw_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err),
				.pld_10g_rx_pempty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty),
				.pld_10g_rx_pfull(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull),
				.pld_8g_a1a2_k1k2_flag(w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag),
				.pld_8g_empty_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf),
				.pld_8g_empty_rx(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx),
				.pld_8g_full_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf),
				.pld_8g_full_rx(w_hssi_rx_pld_pcs_interface_pld_8g_full_rx),
				.pld_8g_rxelecidle(w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle),
				.pld_8g_signal_detect_out(w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out),
				.pld_8g_wa_boundary(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary),
				.pld_pcs_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out),
				.pld_pma_clkdiv_rx_user(w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user),
				.pld_pma_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out),
				.pld_pma_signal_ok(w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok),
				.pld_rx_control(w_hssi_rx_pld_pcs_interface_pld_rx_control),
				.pld_rx_data(w_hssi_rx_pld_pcs_interface_pld_rx_data),
				.pld_rx_prbs_done(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done),
				.pld_rx_prbs_err(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.int_pldif_10g_rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.int_pldif_10g_rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.int_pldif_10g_rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_10g_rx_control({w_hssi_10g_rx_pcs_rx_control[19], w_hssi_10g_rx_pcs_rx_control[18], w_hssi_10g_rx_pcs_rx_control[17], w_hssi_10g_rx_pcs_rx_control[16], w_hssi_10g_rx_pcs_rx_control[15], w_hssi_10g_rx_pcs_rx_control[14], w_hssi_10g_rx_pcs_rx_control[13], w_hssi_10g_rx_pcs_rx_control[12], w_hssi_10g_rx_pcs_rx_control[11], w_hssi_10g_rx_pcs_rx_control[10], w_hssi_10g_rx_pcs_rx_control[9], w_hssi_10g_rx_pcs_rx_control[8], w_hssi_10g_rx_pcs_rx_control[7], w_hssi_10g_rx_pcs_rx_control[6], w_hssi_10g_rx_pcs_rx_control[5], w_hssi_10g_rx_pcs_rx_control[4], w_hssi_10g_rx_pcs_rx_control[3], w_hssi_10g_rx_pcs_rx_control[2], w_hssi_10g_rx_pcs_rx_control[1], w_hssi_10g_rx_pcs_rx_control[0]}),
				.int_pldif_10g_rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.int_pldif_10g_rx_data({w_hssi_10g_rx_pcs_rx_data[127], w_hssi_10g_rx_pcs_rx_data[126], w_hssi_10g_rx_pcs_rx_data[125], w_hssi_10g_rx_pcs_rx_data[124], w_hssi_10g_rx_pcs_rx_data[123], w_hssi_10g_rx_pcs_rx_data[122], w_hssi_10g_rx_pcs_rx_data[121], w_hssi_10g_rx_pcs_rx_data[120], w_hssi_10g_rx_pcs_rx_data[119], w_hssi_10g_rx_pcs_rx_data[118], w_hssi_10g_rx_pcs_rx_data[117], w_hssi_10g_rx_pcs_rx_data[116], w_hssi_10g_rx_pcs_rx_data[115], w_hssi_10g_rx_pcs_rx_data[114], w_hssi_10g_rx_pcs_rx_data[113], w_hssi_10g_rx_pcs_rx_data[112], w_hssi_10g_rx_pcs_rx_data[111], w_hssi_10g_rx_pcs_rx_data[110], w_hssi_10g_rx_pcs_rx_data[109], w_hssi_10g_rx_pcs_rx_data[108], w_hssi_10g_rx_pcs_rx_data[107], w_hssi_10g_rx_pcs_rx_data[106], w_hssi_10g_rx_pcs_rx_data[105], w_hssi_10g_rx_pcs_rx_data[104], w_hssi_10g_rx_pcs_rx_data[103], w_hssi_10g_rx_pcs_rx_data[102], w_hssi_10g_rx_pcs_rx_data[101], w_hssi_10g_rx_pcs_rx_data[100], w_hssi_10g_rx_pcs_rx_data[99], w_hssi_10g_rx_pcs_rx_data[98], w_hssi_10g_rx_pcs_rx_data[97], w_hssi_10g_rx_pcs_rx_data[96], w_hssi_10g_rx_pcs_rx_data[95], w_hssi_10g_rx_pcs_rx_data[94], w_hssi_10g_rx_pcs_rx_data[93], w_hssi_10g_rx_pcs_rx_data[92], w_hssi_10g_rx_pcs_rx_data[91], w_hssi_10g_rx_pcs_rx_data[90], w_hssi_10g_rx_pcs_rx_data[89], w_hssi_10g_rx_pcs_rx_data[88], w_hssi_10g_rx_pcs_rx_data[87], w_hssi_10g_rx_pcs_rx_data[86], w_hssi_10g_rx_pcs_rx_data[85], w_hssi_10g_rx_pcs_rx_data[84], w_hssi_10g_rx_pcs_rx_data[83], w_hssi_10g_rx_pcs_rx_data[82], w_hssi_10g_rx_pcs_rx_data[81], w_hssi_10g_rx_pcs_rx_data[80], w_hssi_10g_rx_pcs_rx_data[79], w_hssi_10g_rx_pcs_rx_data[78], w_hssi_10g_rx_pcs_rx_data[77], w_hssi_10g_rx_pcs_rx_data[76], w_hssi_10g_rx_pcs_rx_data[75], w_hssi_10g_rx_pcs_rx_data[74], w_hssi_10g_rx_pcs_rx_data[73], w_hssi_10g_rx_pcs_rx_data[72], w_hssi_10g_rx_pcs_rx_data[71], w_hssi_10g_rx_pcs_rx_data[70], w_hssi_10g_rx_pcs_rx_data[69], w_hssi_10g_rx_pcs_rx_data[68], w_hssi_10g_rx_pcs_rx_data[67], w_hssi_10g_rx_pcs_rx_data[66], w_hssi_10g_rx_pcs_rx_data[65], w_hssi_10g_rx_pcs_rx_data[64], w_hssi_10g_rx_pcs_rx_data[63], w_hssi_10g_rx_pcs_rx_data[62], w_hssi_10g_rx_pcs_rx_data[61], w_hssi_10g_rx_pcs_rx_data[60], w_hssi_10g_rx_pcs_rx_data[59], w_hssi_10g_rx_pcs_rx_data[58], w_hssi_10g_rx_pcs_rx_data[57], w_hssi_10g_rx_pcs_rx_data[56], w_hssi_10g_rx_pcs_rx_data[55], w_hssi_10g_rx_pcs_rx_data[54], w_hssi_10g_rx_pcs_rx_data[53], w_hssi_10g_rx_pcs_rx_data[52], w_hssi_10g_rx_pcs_rx_data[51], w_hssi_10g_rx_pcs_rx_data[50], w_hssi_10g_rx_pcs_rx_data[49], w_hssi_10g_rx_pcs_rx_data[48], w_hssi_10g_rx_pcs_rx_data[47], w_hssi_10g_rx_pcs_rx_data[46], w_hssi_10g_rx_pcs_rx_data[45], w_hssi_10g_rx_pcs_rx_data[44], w_hssi_10g_rx_pcs_rx_data[43], w_hssi_10g_rx_pcs_rx_data[42], w_hssi_10g_rx_pcs_rx_data[41], w_hssi_10g_rx_pcs_rx_data[40], w_hssi_10g_rx_pcs_rx_data[39], w_hssi_10g_rx_pcs_rx_data[38], w_hssi_10g_rx_pcs_rx_data[37], w_hssi_10g_rx_pcs_rx_data[36], w_hssi_10g_rx_pcs_rx_data[35], w_hssi_10g_rx_pcs_rx_data[34], w_hssi_10g_rx_pcs_rx_data[33], w_hssi_10g_rx_pcs_rx_data[32], w_hssi_10g_rx_pcs_rx_data[31], w_hssi_10g_rx_pcs_rx_data[30], w_hssi_10g_rx_pcs_rx_data[29], w_hssi_10g_rx_pcs_rx_data[28], w_hssi_10g_rx_pcs_rx_data[27], w_hssi_10g_rx_pcs_rx_data[26], w_hssi_10g_rx_pcs_rx_data[25], w_hssi_10g_rx_pcs_rx_data[24], w_hssi_10g_rx_pcs_rx_data[23], w_hssi_10g_rx_pcs_rx_data[22], w_hssi_10g_rx_pcs_rx_data[21], w_hssi_10g_rx_pcs_rx_data[20], w_hssi_10g_rx_pcs_rx_data[19], w_hssi_10g_rx_pcs_rx_data[18], w_hssi_10g_rx_pcs_rx_data[17], w_hssi_10g_rx_pcs_rx_data[16], w_hssi_10g_rx_pcs_rx_data[15], w_hssi_10g_rx_pcs_rx_data[14], w_hssi_10g_rx_pcs_rx_data[13], w_hssi_10g_rx_pcs_rx_data[12], w_hssi_10g_rx_pcs_rx_data[11], w_hssi_10g_rx_pcs_rx_data[10], w_hssi_10g_rx_pcs_rx_data[9], w_hssi_10g_rx_pcs_rx_data[8], w_hssi_10g_rx_pcs_rx_data[7], w_hssi_10g_rx_pcs_rx_data[6], w_hssi_10g_rx_pcs_rx_data[5], w_hssi_10g_rx_pcs_rx_data[4], w_hssi_10g_rx_pcs_rx_data[3], w_hssi_10g_rx_pcs_rx_data[2], w_hssi_10g_rx_pcs_rx_data[1], w_hssi_10g_rx_pcs_rx_data[0]}),
				.int_pldif_10g_rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.int_pldif_10g_rx_diag_status({w_hssi_10g_rx_pcs_rx_diag_status[1], w_hssi_10g_rx_pcs_rx_diag_status[0]}),
				.int_pldif_10g_rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.int_pldif_10g_rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.int_pldif_10g_rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.int_pldif_10g_rx_fifo_num({w_hssi_10g_rx_pcs_rx_fifo_num[4], w_hssi_10g_rx_pcs_rx_fifo_num[3], w_hssi_10g_rx_pcs_rx_fifo_num[2], w_hssi_10g_rx_pcs_rx_fifo_num[1], w_hssi_10g_rx_pcs_rx_fifo_num[0]}),
				.int_pldif_10g_rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.int_pldif_10g_rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.int_pldif_10g_rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.int_pldif_10g_rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.int_pldif_10g_rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.int_pldif_10g_rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				.int_pldif_8g_a1a2_k1k2_flag({w_hssi_8g_rx_pcs_a1a2k1k2flag[3], w_hssi_8g_rx_pcs_a1a2k1k2flag[2], w_hssi_8g_rx_pcs_a1a2k1k2flag[1], w_hssi_8g_rx_pcs_a1a2k1k2flag[0]}),
				.int_pldif_8g_empty_rmf(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.int_pldif_8g_empty_rx(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.int_pldif_8g_full_rmf(w_hssi_8g_rx_pcs_rm_fifo_full),
				.int_pldif_8g_full_rx(w_hssi_8g_rx_pcs_pcfifofull),
				.int_pldif_8g_phystatus(w_hssi_8g_rx_pcs_phystatus),
				.int_pldif_8g_rx_blk_start({w_hssi_8g_rx_pcs_rx_blk_start[3], w_hssi_8g_rx_pcs_rx_blk_start[2], w_hssi_8g_rx_pcs_rx_blk_start[1], w_hssi_8g_rx_pcs_rx_blk_start[0]}),
				.int_pldif_8g_rx_clk(w_hssi_8g_rx_pcs_clock_to_pld),
				.int_pldif_8g_rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_8g_rx_data_valid({w_hssi_8g_rx_pcs_rx_data_valid[3], w_hssi_8g_rx_pcs_rx_data_valid[2], w_hssi_8g_rx_pcs_rx_data_valid[1], w_hssi_8g_rx_pcs_rx_data_valid[0]}),
				.int_pldif_8g_rx_rstn_sync2wrfifo(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.int_pldif_8g_rx_sync_hdr({w_hssi_8g_rx_pcs_rx_sync_hdr[1], w_hssi_8g_rx_pcs_rx_sync_hdr[0]}),
				.int_pldif_8g_rxd({w_hssi_8g_rx_pcs_dataout[63], w_hssi_8g_rx_pcs_dataout[62], w_hssi_8g_rx_pcs_dataout[61], w_hssi_8g_rx_pcs_dataout[60], w_hssi_8g_rx_pcs_dataout[59], w_hssi_8g_rx_pcs_dataout[58], w_hssi_8g_rx_pcs_dataout[57], w_hssi_8g_rx_pcs_dataout[56], w_hssi_8g_rx_pcs_dataout[55], w_hssi_8g_rx_pcs_dataout[54], w_hssi_8g_rx_pcs_dataout[53], w_hssi_8g_rx_pcs_dataout[52], w_hssi_8g_rx_pcs_dataout[51], w_hssi_8g_rx_pcs_dataout[50], w_hssi_8g_rx_pcs_dataout[49], w_hssi_8g_rx_pcs_dataout[48], w_hssi_8g_rx_pcs_dataout[47], w_hssi_8g_rx_pcs_dataout[46], w_hssi_8g_rx_pcs_dataout[45], w_hssi_8g_rx_pcs_dataout[44], w_hssi_8g_rx_pcs_dataout[43], w_hssi_8g_rx_pcs_dataout[42], w_hssi_8g_rx_pcs_dataout[41], w_hssi_8g_rx_pcs_dataout[40], w_hssi_8g_rx_pcs_dataout[39], w_hssi_8g_rx_pcs_dataout[38], w_hssi_8g_rx_pcs_dataout[37], w_hssi_8g_rx_pcs_dataout[36], w_hssi_8g_rx_pcs_dataout[35], w_hssi_8g_rx_pcs_dataout[34], w_hssi_8g_rx_pcs_dataout[33], w_hssi_8g_rx_pcs_dataout[32], w_hssi_8g_rx_pcs_dataout[31], w_hssi_8g_rx_pcs_dataout[30], w_hssi_8g_rx_pcs_dataout[29], w_hssi_8g_rx_pcs_dataout[28], w_hssi_8g_rx_pcs_dataout[27], w_hssi_8g_rx_pcs_dataout[26], w_hssi_8g_rx_pcs_dataout[25], w_hssi_8g_rx_pcs_dataout[24], w_hssi_8g_rx_pcs_dataout[23], w_hssi_8g_rx_pcs_dataout[22], w_hssi_8g_rx_pcs_dataout[21], w_hssi_8g_rx_pcs_dataout[20], w_hssi_8g_rx_pcs_dataout[19], w_hssi_8g_rx_pcs_dataout[18], w_hssi_8g_rx_pcs_dataout[17], w_hssi_8g_rx_pcs_dataout[16], w_hssi_8g_rx_pcs_dataout[15], w_hssi_8g_rx_pcs_dataout[14], w_hssi_8g_rx_pcs_dataout[13], w_hssi_8g_rx_pcs_dataout[12], w_hssi_8g_rx_pcs_dataout[11], w_hssi_8g_rx_pcs_dataout[10], w_hssi_8g_rx_pcs_dataout[9], w_hssi_8g_rx_pcs_dataout[8], w_hssi_8g_rx_pcs_dataout[7], w_hssi_8g_rx_pcs_dataout[6], w_hssi_8g_rx_pcs_dataout[5], w_hssi_8g_rx_pcs_dataout[4], w_hssi_8g_rx_pcs_dataout[3], w_hssi_8g_rx_pcs_dataout[2], w_hssi_8g_rx_pcs_dataout[1], w_hssi_8g_rx_pcs_dataout[0]}),
				.int_pldif_8g_rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.int_pldif_8g_rxstatus({w_hssi_8g_rx_pcs_rxstatus[2], w_hssi_8g_rx_pcs_rxstatus[1], w_hssi_8g_rx_pcs_rxstatus[0]}),
				.int_pldif_8g_rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.int_pldif_8g_signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.int_pldif_8g_wa_boundary({w_hssi_8g_rx_pcs_word_align_boundary[4], w_hssi_8g_rx_pcs_word_align_boundary[3], w_hssi_8g_rx_pcs_word_align_boundary[2], w_hssi_8g_rx_pcs_word_align_boundary[1], w_hssi_8g_rx_pcs_word_align_boundary[0]}),
				.int_pldif_krfec_rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.int_pldif_krfec_rx_data_status({w_hssi_krfec_rx_pcs_rx_data_status[1], w_hssi_krfec_rx_pcs_rx_data_status[0]}),
				.int_pldif_krfec_rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.int_pldif_pmaif_clkdiv_rx(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pldif_pmaif_clkdiv_rx_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pldif_pmaif_rx_data({w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0]}),
				.int_pldif_pmaif_rx_prbs_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pldif_pmaif_rx_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.pld_10g_krfec_rx_clr_errblk_cnt(in_pld_10g_krfec_rx_clr_errblk_cnt),
				.pld_10g_krfec_rx_pld_rst_n(in_pld_10g_krfec_rx_pld_rst_n),
				.pld_10g_rx_align_clr(in_pld_10g_rx_align_clr),
				.pld_10g_rx_clr_ber_count(in_pld_10g_rx_clr_ber_count),
				.pld_10g_rx_rd_en(in_pld_10g_rx_rd_en),
				.pld_8g_a1a2_size(in_pld_8g_a1a2_size),
				.pld_8g_bitloc_rev_en(in_pld_8g_bitloc_rev_en),
				.pld_8g_byte_rev_en(in_pld_8g_byte_rev_en),
				.pld_8g_encdt(in_pld_8g_encdt),
				.pld_8g_g3_rx_pld_rst_n(in_pld_8g_g3_rx_pld_rst_n),
				.pld_8g_rdenable_rx(in_pld_8g_rdenable_rx),
				.pld_8g_rxpolarity(in_pld_8g_rxpolarity),
				.pld_8g_wrdisable_rx(in_pld_8g_wrdisable_rx),
				.pld_bitslip(in_pld_bitslip),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_rxpma_rstb(in_pld_pma_rxpma_rstb),
				.pld_pmaif_rx_pld_rst_n(in_pld_pmaif_rx_pld_rst_n),
				.pld_pmaif_rxclkslip(in_pld_pmaif_rxclkslip),
				.pld_polinv_rx(in_pld_polinv_rx),
				.pld_rx_clk(in_pld_rx_clk),
				.pld_rx_prbs_err_clr(in_pld_rx_prbs_err_clr),
				.pld_syncsm_en(in_pld_syncsm_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.int_pldif_pmaif_rx_pld_clk(),
				.pld_8g_wa_boundary_txclk_fastreg(),
				.pld_8g_wa_boundary_txclk_reg(),
				.pld_bitslip_10g_txclk_reg(),
				.pld_bitslip_8g_txclk_reg(),
				.pld_bitslip_rxclk_parallel_loopback_reg(),
				.pld_bitslip_rxclk_reg(),
				.pld_pcs_rx_clk_out_pcsdirect_wire(),
				.pld_pma_rx_clk_out_10g_or_pcsdirect_wire(),
				.pld_pma_rx_clk_out_8g_wire(),
				.pld_pmaif_rx_pld_rst_n_reg(),
				.pld_pmaif_tx_pld_rst_n_txclk_reg(),
				.pld_polinv_rx_reg(),
				.pld_rx_clk_fifo(),
				.pld_rx_control_fifo(),
				.pld_rx_control_pcsdirect_reg(),
				.pld_rx_data_fifo(),
				.pld_rx_data_pcsdirect_reg(),
				.pld_rx_prbs_done_reg(),
				.pld_rx_prbs_done_txclk_reg(),
				.pld_rx_prbs_err_clr_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_clr_reg(),
				.pld_rx_prbs_err_disprbs_reg(),
				.pld_rx_prbs_err_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_reg(),
				.pma_rx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_data[50:0] = 51'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3:0] = 4'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_control[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_data[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pcs_pma_interface
			twentynm_hssi_tx_pcs_pma_interface #(
				.bypass_pma_txelecidle(hssi_tx_pcs_pma_interface_bypass_pma_txelecidle),
				.channel_operation_mode(hssi_tx_pcs_pma_interface_channel_operation_mode),
				.lpbk_en(hssi_tx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_tx_pcs_pma_interface_master_clk_sel),
				.pcie_sub_prot_mode_tx(hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx),
				.pldif_datawidth_mode(hssi_tx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_tx(hssi_tx_pcs_pma_interface_pma_dw_tx),
				.pma_if_dft_en(hssi_tx_pcs_pma_interface_pma_if_dft_en),
				.pmagate_en(hssi_tx_pcs_pma_interface_pmagate_en),
				.prbs9_dwidth(hssi_tx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_tx_pcs_pma_interface_prbs_clken),
				.prbs_gen_pat(hssi_tx_pcs_pma_interface_prbs_gen_pat),
				.prot_mode_tx(hssi_tx_pcs_pma_interface_prot_mode_tx),
				.reconfig_settings(hssi_tx_pcs_pma_interface_reconfig_settings),
				.silicon_rev( "20nm5es" ),       //PARAM_HIDE
				.sq_wave_num(hssi_tx_pcs_pma_interface_sq_wave_num),
				.sqwgen_clken(hssi_tx_pcs_pma_interface_sqwgen_clken),
				.sup_mode(hssi_tx_pcs_pma_interface_sup_mode),
				.tx_dyn_polarity_inversion(hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion),
				.tx_pma_data_sel(hssi_tx_pcs_pma_interface_tx_pma_data_sel),
				.tx_static_polarity_inversion(hssi_tx_pcs_pma_interface_tx_static_polarity_inversion),
				.uhsif_cnt_step_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock),
				.uhsif_cnt_thresh_filt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value),
				.uhsif_cnt_thresh_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock),
				.uhsif_dcn_test_update_period(hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period),
				.uhsif_dcn_testmode_enable(hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable),
				.uhsif_dead_zone_count_thresh(hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh),
				.uhsif_dead_zone_detection_enable(hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable),
				.uhsif_dead_zone_obser_window(hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window),
				.uhsif_dead_zone_skip_size(hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size),
				.uhsif_delay_cell_index_sel(hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel),
				.uhsif_delay_cell_margin(hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin),
				.uhsif_delay_cell_static_index_value(hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value),
				.uhsif_dft_dead_zone_control(hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control),
				.uhsif_dft_up_filt_control(hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control),
				.uhsif_enable(hssi_tx_pcs_pma_interface_uhsif_enable),
				.uhsif_lock_det_segsz_after_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock),
				.uhsif_lock_det_segsz_before_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock),
				.uhsif_lock_det_thresh_cnt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value),
				.uhsif_lock_det_thresh_cnt_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value),
				.uhsif_lock_det_thresh_diff_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value),
				.uhsif_lock_det_thresh_diff_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value)
			) inst_twentynm_hssi_tx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.int_pmaif_8g_txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.int_pmaif_pldif_tx_clkdiv(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pmaif_pldif_tx_clkdiv_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pmaif_pldif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.int_pmaif_pldif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.int_tx_dft_obsrv_clk(w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk),
				.pma_tx_elec_idle(w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle),
				.pma_tx_pma_data(w_hssi_tx_pcs_pma_interface_pma_tx_pma_data),
				.pma_txpma_rstb(w_hssi_tx_pcs_pma_interface_pma_txpma_rstb),
				.tx_pma_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback),
				.tx_pma_uhsif_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback),
				.tx_prbs_gen_test(w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test),
				.uhsif_test_out_1(w_hssi_tx_pcs_pma_interface_uhsif_test_out_1),
				.uhsif_test_out_2(w_hssi_tx_pcs_pma_interface_uhsif_test_out_2),
				.uhsif_test_out_3(w_hssi_tx_pcs_pma_interface_uhsif_test_out_3),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.int_pmaif_10g_tx_pma_data({w_hssi_10g_tx_pcs_tx_pma_data[63], w_hssi_10g_tx_pcs_tx_pma_data[62], w_hssi_10g_tx_pcs_tx_pma_data[61], w_hssi_10g_tx_pcs_tx_pma_data[60], w_hssi_10g_tx_pcs_tx_pma_data[59], w_hssi_10g_tx_pcs_tx_pma_data[58], w_hssi_10g_tx_pcs_tx_pma_data[57], w_hssi_10g_tx_pcs_tx_pma_data[56], w_hssi_10g_tx_pcs_tx_pma_data[55], w_hssi_10g_tx_pcs_tx_pma_data[54], w_hssi_10g_tx_pcs_tx_pma_data[53], w_hssi_10g_tx_pcs_tx_pma_data[52], w_hssi_10g_tx_pcs_tx_pma_data[51], w_hssi_10g_tx_pcs_tx_pma_data[50], w_hssi_10g_tx_pcs_tx_pma_data[49], w_hssi_10g_tx_pcs_tx_pma_data[48], w_hssi_10g_tx_pcs_tx_pma_data[47], w_hssi_10g_tx_pcs_tx_pma_data[46], w_hssi_10g_tx_pcs_tx_pma_data[45], w_hssi_10g_tx_pcs_tx_pma_data[44], w_hssi_10g_tx_pcs_tx_pma_data[43], w_hssi_10g_tx_pcs_tx_pma_data[42], w_hssi_10g_tx_pcs_tx_pma_data[41], w_hssi_10g_tx_pcs_tx_pma_data[40], w_hssi_10g_tx_pcs_tx_pma_data[39], w_hssi_10g_tx_pcs_tx_pma_data[38], w_hssi_10g_tx_pcs_tx_pma_data[37], w_hssi_10g_tx_pcs_tx_pma_data[36], w_hssi_10g_tx_pcs_tx_pma_data[35], w_hssi_10g_tx_pcs_tx_pma_data[34], w_hssi_10g_tx_pcs_tx_pma_data[33], w_hssi_10g_tx_pcs_tx_pma_data[32], w_hssi_10g_tx_pcs_tx_pma_data[31], w_hssi_10g_tx_pcs_tx_pma_data[30], w_hssi_10g_tx_pcs_tx_pma_data[29], w_hssi_10g_tx_pcs_tx_pma_data[28], w_hssi_10g_tx_pcs_tx_pma_data[27], w_hssi_10g_tx_pcs_tx_pma_data[26], w_hssi_10g_tx_pcs_tx_pma_data[25], w_hssi_10g_tx_pcs_tx_pma_data[24], w_hssi_10g_tx_pcs_tx_pma_data[23], w_hssi_10g_tx_pcs_tx_pma_data[22], w_hssi_10g_tx_pcs_tx_pma_data[21], w_hssi_10g_tx_pcs_tx_pma_data[20], w_hssi_10g_tx_pcs_tx_pma_data[19], w_hssi_10g_tx_pcs_tx_pma_data[18], w_hssi_10g_tx_pcs_tx_pma_data[17], w_hssi_10g_tx_pcs_tx_pma_data[16], w_hssi_10g_tx_pcs_tx_pma_data[15], w_hssi_10g_tx_pcs_tx_pma_data[14], w_hssi_10g_tx_pcs_tx_pma_data[13], w_hssi_10g_tx_pcs_tx_pma_data[12], w_hssi_10g_tx_pcs_tx_pma_data[11], w_hssi_10g_tx_pcs_tx_pma_data[10], w_hssi_10g_tx_pcs_tx_pma_data[9], w_hssi_10g_tx_pcs_tx_pma_data[8], w_hssi_10g_tx_pcs_tx_pma_data[7], w_hssi_10g_tx_pcs_tx_pma_data[6], w_hssi_10g_tx_pcs_tx_pma_data[5], w_hssi_10g_tx_pcs_tx_pma_data[4], w_hssi_10g_tx_pcs_tx_pma_data[3], w_hssi_10g_tx_pcs_tx_pma_data[2], w_hssi_10g_tx_pcs_tx_pma_data[1], w_hssi_10g_tx_pcs_tx_pma_data[0]}),
				.int_pmaif_10g_tx_pma_data_gate_val({w_hssi_10g_tx_pcs_tx_pma_gating_val[63], w_hssi_10g_tx_pcs_tx_pma_gating_val[62], w_hssi_10g_tx_pcs_tx_pma_gating_val[61], w_hssi_10g_tx_pcs_tx_pma_gating_val[60], w_hssi_10g_tx_pcs_tx_pma_gating_val[59], w_hssi_10g_tx_pcs_tx_pma_gating_val[58], w_hssi_10g_tx_pcs_tx_pma_gating_val[57], w_hssi_10g_tx_pcs_tx_pma_gating_val[56], w_hssi_10g_tx_pcs_tx_pma_gating_val[55], w_hssi_10g_tx_pcs_tx_pma_gating_val[54], w_hssi_10g_tx_pcs_tx_pma_gating_val[53], w_hssi_10g_tx_pcs_tx_pma_gating_val[52], w_hssi_10g_tx_pcs_tx_pma_gating_val[51], w_hssi_10g_tx_pcs_tx_pma_gating_val[50], w_hssi_10g_tx_pcs_tx_pma_gating_val[49], w_hssi_10g_tx_pcs_tx_pma_gating_val[48], w_hssi_10g_tx_pcs_tx_pma_gating_val[47], w_hssi_10g_tx_pcs_tx_pma_gating_val[46], w_hssi_10g_tx_pcs_tx_pma_gating_val[45], w_hssi_10g_tx_pcs_tx_pma_gating_val[44], w_hssi_10g_tx_pcs_tx_pma_gating_val[43], w_hssi_10g_tx_pcs_tx_pma_gating_val[42], w_hssi_10g_tx_pcs_tx_pma_gating_val[41], w_hssi_10g_tx_pcs_tx_pma_gating_val[40], w_hssi_10g_tx_pcs_tx_pma_gating_val[39], w_hssi_10g_tx_pcs_tx_pma_gating_val[38], w_hssi_10g_tx_pcs_tx_pma_gating_val[37], w_hssi_10g_tx_pcs_tx_pma_gating_val[36], w_hssi_10g_tx_pcs_tx_pma_gating_val[35], w_hssi_10g_tx_pcs_tx_pma_gating_val[34], w_hssi_10g_tx_pcs_tx_pma_gating_val[33], w_hssi_10g_tx_pcs_tx_pma_gating_val[32], w_hssi_10g_tx_pcs_tx_pma_gating_val[31], w_hssi_10g_tx_pcs_tx_pma_gating_val[30], w_hssi_10g_tx_pcs_tx_pma_gating_val[29], w_hssi_10g_tx_pcs_tx_pma_gating_val[28], w_hssi_10g_tx_pcs_tx_pma_gating_val[27], w_hssi_10g_tx_pcs_tx_pma_gating_val[26], w_hssi_10g_tx_pcs_tx_pma_gating_val[25], w_hssi_10g_tx_pcs_tx_pma_gating_val[24], w_hssi_10g_tx_pcs_tx_pma_gating_val[23], w_hssi_10g_tx_pcs_tx_pma_gating_val[22], w_hssi_10g_tx_pcs_tx_pma_gating_val[21], w_hssi_10g_tx_pcs_tx_pma_gating_val[20], w_hssi_10g_tx_pcs_tx_pma_gating_val[19], w_hssi_10g_tx_pcs_tx_pma_gating_val[18], w_hssi_10g_tx_pcs_tx_pma_gating_val[17], w_hssi_10g_tx_pcs_tx_pma_gating_val[16], w_hssi_10g_tx_pcs_tx_pma_gating_val[15], w_hssi_10g_tx_pcs_tx_pma_gating_val[14], w_hssi_10g_tx_pcs_tx_pma_gating_val[13], w_hssi_10g_tx_pcs_tx_pma_gating_val[12], w_hssi_10g_tx_pcs_tx_pma_gating_val[11], w_hssi_10g_tx_pcs_tx_pma_gating_val[10], w_hssi_10g_tx_pcs_tx_pma_gating_val[9], w_hssi_10g_tx_pcs_tx_pma_gating_val[8], w_hssi_10g_tx_pcs_tx_pma_gating_val[7], w_hssi_10g_tx_pcs_tx_pma_gating_val[6], w_hssi_10g_tx_pcs_tx_pma_gating_val[5], w_hssi_10g_tx_pcs_tx_pma_gating_val[4], w_hssi_10g_tx_pcs_tx_pma_gating_val[3], w_hssi_10g_tx_pcs_tx_pma_gating_val[2], w_hssi_10g_tx_pcs_tx_pma_gating_val[1], w_hssi_10g_tx_pcs_tx_pma_gating_val[0]}),
				.int_pmaif_8g_pudr({w_hssi_8g_tx_pcs_dataout[19], w_hssi_8g_tx_pcs_dataout[18], w_hssi_8g_tx_pcs_dataout[17], w_hssi_8g_tx_pcs_dataout[16], w_hssi_8g_tx_pcs_dataout[15], w_hssi_8g_tx_pcs_dataout[14], w_hssi_8g_tx_pcs_dataout[13], w_hssi_8g_tx_pcs_dataout[12], w_hssi_8g_tx_pcs_dataout[11], w_hssi_8g_tx_pcs_dataout[10], w_hssi_8g_tx_pcs_dataout[9], w_hssi_8g_tx_pcs_dataout[8], w_hssi_8g_tx_pcs_dataout[7], w_hssi_8g_tx_pcs_dataout[6], w_hssi_8g_tx_pcs_dataout[5], w_hssi_8g_tx_pcs_dataout[4], w_hssi_8g_tx_pcs_dataout[3], w_hssi_8g_tx_pcs_dataout[2], w_hssi_8g_tx_pcs_dataout[1], w_hssi_8g_tx_pcs_dataout[0]}),
				.int_pmaif_8g_tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.int_pmaif_8g_tx_elec_idle(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_pma_data_out({w_hssi_gen3_tx_pcs_data_out[31], w_hssi_gen3_tx_pcs_data_out[30], w_hssi_gen3_tx_pcs_data_out[29], w_hssi_gen3_tx_pcs_data_out[28], w_hssi_gen3_tx_pcs_data_out[27], w_hssi_gen3_tx_pcs_data_out[26], w_hssi_gen3_tx_pcs_data_out[25], w_hssi_gen3_tx_pcs_data_out[24], w_hssi_gen3_tx_pcs_data_out[23], w_hssi_gen3_tx_pcs_data_out[22], w_hssi_gen3_tx_pcs_data_out[21], w_hssi_gen3_tx_pcs_data_out[20], w_hssi_gen3_tx_pcs_data_out[19], w_hssi_gen3_tx_pcs_data_out[18], w_hssi_gen3_tx_pcs_data_out[17], w_hssi_gen3_tx_pcs_data_out[16], w_hssi_gen3_tx_pcs_data_out[15], w_hssi_gen3_tx_pcs_data_out[14], w_hssi_gen3_tx_pcs_data_out[13], w_hssi_gen3_tx_pcs_data_out[12], w_hssi_gen3_tx_pcs_data_out[11], w_hssi_gen3_tx_pcs_data_out[10], w_hssi_gen3_tx_pcs_data_out[9], w_hssi_gen3_tx_pcs_data_out[8], w_hssi_gen3_tx_pcs_data_out[7], w_hssi_gen3_tx_pcs_data_out[6], w_hssi_gen3_tx_pcs_data_out[5], w_hssi_gen3_tx_pcs_data_out[4], w_hssi_gen3_tx_pcs_data_out[3], w_hssi_gen3_tx_pcs_data_out[2], w_hssi_gen3_tx_pcs_data_out[1], w_hssi_gen3_tx_pcs_data_out[0]}),
				.int_pmaif_g3_pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.int_pmaif_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pmaif_pldif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pmaif_pldif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0]}),
				.int_pmaif_pldif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pmaif_pldif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.int_pmaif_pldif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pmaif_pldif_uhsif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0]}),
				.pma_tx_clkdiv_user(in_pma_tx_clkdiv_user),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.refclk_dig_uhsif(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.uhsif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.uhsif_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				
				// UNUSED
				.avmm_user_dataout(),
				.write_en(),
				.write_en_ack()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4:0] = 5'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_txpma_rstb = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pld_pcs_interface
			twentynm_hssi_tx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx),
				.hd_10g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx),
				.hd_10g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx),
				.hd_10g_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx),
				.hd_10g_lpbk_en(hssi_tx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx),
				.hd_10g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx),
				.hd_10g_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx),
				.hd_8g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx),
				.hd_8g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx),
				.hd_8g_hip_mode(hssi_tx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_tx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx),
				.hd_8g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx),
				.hd_chnl_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx),
				.hd_chnl_frequency_rules_en(hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_tx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_tx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx),
				.hd_chnl_lpbk_en(hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx),
				.hd_chnl_pld_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz),
				.hd_chnl_pld_uhsif_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz),
				.hd_chnl_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx),
				.hd_chnl_pma_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz),
				.hd_chnl_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx),
				.hd_chnl_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx),
				.hd_fifo_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx),
				.hd_fifo_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx),
				.hd_g3_prot_mode(hssi_tx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx),
				.hd_krfec_lpbk_en(hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx),
				.hd_pldif_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx),
				.hd_pmaif_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_ctrl_plane_bonding(hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding),
				.hd_pmaif_lpbk_en(hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx),
				.hd_pmaif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx),
				.hd_pmaif_sim_mode(hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_tx_clk_out_sel(hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel),
				.pcs_tx_clk_source(hssi_tx_pld_pcs_interface_pcs_tx_clk_source),
				.pcs_tx_data_source(hssi_tx_pld_pcs_interface_pcs_tx_data_source),
				.pcs_tx_delay1_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en),
				.pcs_tx_delay1_clk_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel),
				.pcs_tx_delay1_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl),
				.pcs_tx_delay1_data_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel),
				.pcs_tx_delay2_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en),
				.pcs_tx_delay2_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl),
				.pcs_tx_output_sel(hssi_tx_pld_pcs_interface_pcs_tx_output_sel),
				.reconfig_settings(hssi_tx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm5es" )       //PARAM_HIDE
			) inst_twentynm_hssi_tx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pld_pcs_interface_blockselect),
				.hip_tx_clk(w_hssi_tx_pld_pcs_interface_hip_tx_clk),
				.int_pldif_10g_tx_bitslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip),
				.int_pldif_10g_tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.int_pldif_10g_tx_control(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control),
				.int_pldif_10g_tx_control_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg),
				.int_pldif_10g_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data),
				.int_pldif_10g_tx_data_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg),
				.int_pldif_10g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.int_pldif_10g_tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.int_pldif_10g_tx_diag_status(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status),
				.int_pldif_10g_tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.int_pldif_10g_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.int_pldif_10g_tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				.int_pldif_8g_pld_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.int_pldif_8g_powerdown(w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown),
				.int_pldif_8g_rddisable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.int_pldif_8g_rev_loopbk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.int_pldif_8g_tx_blk_start(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start),
				.int_pldif_8g_tx_boundary_sel(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel),
				.int_pldif_8g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid),
				.int_pldif_8g_tx_sync_hdr(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr),
				.int_pldif_8g_txd(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd),
				.int_pldif_8g_txd_fast_reg(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg),
				.int_pldif_8g_txdeemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.int_pldif_8g_txdetectrxloopback(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.int_pldif_8g_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.int_pldif_8g_txmargin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin),
				.int_pldif_8g_txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.int_pldif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.int_pldif_8g_wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				.int_pldif_pmaif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pldif_pmaif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pldif_pmaif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data),
				.int_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pldif_pmaif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pldif_pmaif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pldif_pmaif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pldif_pmaif_uhsif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data),
				.pld_10g_krfec_tx_frame(w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame),
				.pld_10g_tx_burst_en_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe),
				.pld_10g_tx_empty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty),
				.pld_10g_tx_fifo_num(w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num),
				.pld_10g_tx_full(w_hssi_tx_pld_pcs_interface_pld_10g_tx_full),
				.pld_10g_tx_pempty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty),
				.pld_10g_tx_pfull(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull),
				.pld_10g_tx_wordslip_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe),
				.pld_8g_empty_tx(w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx),
				.pld_8g_full_tx(w_hssi_tx_pld_pcs_interface_pld_8g_full_tx),
				.pld_krfec_tx_alignment(w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment),
				.pld_pcs_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out),
				.pld_pma_clkdiv_tx_user(w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user),
				.pld_pma_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out),
				.pld_uhsif_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.hip_tx_data({in_hip_tx_data[63], in_hip_tx_data[62], in_hip_tx_data[61], in_hip_tx_data[60], in_hip_tx_data[59], in_hip_tx_data[58], in_hip_tx_data[57], in_hip_tx_data[56], in_hip_tx_data[55], in_hip_tx_data[54], in_hip_tx_data[53], in_hip_tx_data[52], in_hip_tx_data[51], in_hip_tx_data[50], in_hip_tx_data[49], in_hip_tx_data[48], in_hip_tx_data[47], in_hip_tx_data[46], in_hip_tx_data[45], in_hip_tx_data[44], in_hip_tx_data[43], in_hip_tx_data[42], in_hip_tx_data[41], in_hip_tx_data[40], in_hip_tx_data[39], in_hip_tx_data[38], in_hip_tx_data[37], in_hip_tx_data[36], in_hip_tx_data[35], in_hip_tx_data[34], in_hip_tx_data[33], in_hip_tx_data[32], in_hip_tx_data[31], in_hip_tx_data[30], in_hip_tx_data[29], in_hip_tx_data[28], in_hip_tx_data[27], in_hip_tx_data[26], in_hip_tx_data[25], in_hip_tx_data[24], in_hip_tx_data[23], in_hip_tx_data[22], in_hip_tx_data[21], in_hip_tx_data[20], in_hip_tx_data[19], in_hip_tx_data[18], in_hip_tx_data[17], in_hip_tx_data[16], in_hip_tx_data[15], in_hip_tx_data[14], in_hip_tx_data[13], in_hip_tx_data[12], in_hip_tx_data[11], in_hip_tx_data[10], in_hip_tx_data[9], in_hip_tx_data[8], in_hip_tx_data[7], in_hip_tx_data[6], in_hip_tx_data[5], in_hip_tx_data[4], in_hip_tx_data[3], in_hip_tx_data[2], in_hip_tx_data[1], in_hip_tx_data[0]}),
				.int_pldif_10g_tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.int_pldif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.int_pldif_10g_tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_10g_tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.int_pldif_10g_tx_fifo_num({w_hssi_10g_tx_pcs_tx_fifo_num[3], w_hssi_10g_tx_pcs_tx_fifo_num[2], w_hssi_10g_tx_pcs_tx_fifo_num[1], w_hssi_10g_tx_pcs_tx_fifo_num[0]}),
				.int_pldif_10g_tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.int_pldif_10g_tx_full(w_hssi_10g_tx_pcs_tx_full),
				.int_pldif_10g_tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.int_pldif_10g_tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.int_pldif_10g_tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				.int_pldif_8g_empty_tx(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.int_pldif_8g_full_tx(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.int_pldif_8g_tx_clk_out(w_hssi_8g_tx_pcs_clk_out),
				.int_pldif_8g_tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_krfec_tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.int_pldif_krfec_tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.int_pldif_pmaif_clkdiv_tx(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pldif_pmaif_clkdiv_tx_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pldif_pmaif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.pld_10g_krfec_tx_pld_rst_n(in_pld_10g_krfec_tx_pld_rst_n),
				.pld_10g_tx_bitslip({in_pld_10g_tx_bitslip[6], in_pld_10g_tx_bitslip[5], in_pld_10g_tx_bitslip[4], in_pld_10g_tx_bitslip[3], in_pld_10g_tx_bitslip[2], in_pld_10g_tx_bitslip[1], in_pld_10g_tx_bitslip[0]}),
				.pld_10g_tx_burst_en(in_pld_10g_tx_burst_en),
				.pld_10g_tx_data_valid(in_pld_10g_tx_data_valid),
				.pld_10g_tx_diag_status({in_pld_10g_tx_diag_status[1], in_pld_10g_tx_diag_status[0]}),
				.pld_10g_tx_wordslip(in_pld_10g_tx_wordslip),
				.pld_8g_g3_tx_pld_rst_n(in_pld_8g_g3_tx_pld_rst_n),
				.pld_8g_rddisable_tx(in_pld_8g_rddisable_tx),
				.pld_8g_tx_boundary_sel({in_pld_8g_tx_boundary_sel[4], in_pld_8g_tx_boundary_sel[3], in_pld_8g_tx_boundary_sel[2], in_pld_8g_tx_boundary_sel[1], in_pld_8g_tx_boundary_sel[0]}),
				.pld_8g_wrenable_tx(in_pld_8g_wrenable_tx),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_txpma_rstb(in_pld_pma_txpma_rstb),
				.pld_pmaif_tx_pld_rst_n(in_pld_pmaif_tx_pld_rst_n),
				.pld_polinv_tx(in_pld_polinv_tx),
				.pld_tx_clk(in_pld_tx_clk),
				.pld_tx_control({in_pld_tx_control[17], in_pld_tx_control[16], in_pld_tx_control[15], in_pld_tx_control[14], in_pld_tx_control[13], in_pld_tx_control[12], in_pld_tx_control[11], in_pld_tx_control[10], in_pld_tx_control[9], in_pld_tx_control[8], in_pld_tx_control[7], in_pld_tx_control[6], in_pld_tx_control[5], in_pld_tx_control[4], in_pld_tx_control[3], in_pld_tx_control[2], in_pld_tx_control[1], in_pld_tx_control[0]}),
				.pld_tx_data({in_pld_tx_data[127], in_pld_tx_data[126], in_pld_tx_data[125], in_pld_tx_data[124], in_pld_tx_data[123], in_pld_tx_data[122], in_pld_tx_data[121], in_pld_tx_data[120], in_pld_tx_data[119], in_pld_tx_data[118], in_pld_tx_data[117], in_pld_tx_data[116], in_pld_tx_data[115], in_pld_tx_data[114], in_pld_tx_data[113], in_pld_tx_data[112], in_pld_tx_data[111], in_pld_tx_data[110], in_pld_tx_data[109], in_pld_tx_data[108], in_pld_tx_data[107], in_pld_tx_data[106], in_pld_tx_data[105], in_pld_tx_data[104], in_pld_tx_data[103], in_pld_tx_data[102], in_pld_tx_data[101], in_pld_tx_data[100], in_pld_tx_data[99], in_pld_tx_data[98], in_pld_tx_data[97], in_pld_tx_data[96], in_pld_tx_data[95], in_pld_tx_data[94], in_pld_tx_data[93], in_pld_tx_data[92], in_pld_tx_data[91], in_pld_tx_data[90], in_pld_tx_data[89], in_pld_tx_data[88], in_pld_tx_data[87], in_pld_tx_data[86], in_pld_tx_data[85], in_pld_tx_data[84], in_pld_tx_data[83], in_pld_tx_data[82], in_pld_tx_data[81], in_pld_tx_data[80], in_pld_tx_data[79], in_pld_tx_data[78], in_pld_tx_data[77], in_pld_tx_data[76], in_pld_tx_data[75], in_pld_tx_data[74], in_pld_tx_data[73], in_pld_tx_data[72], in_pld_tx_data[71], in_pld_tx_data[70], in_pld_tx_data[69], in_pld_tx_data[68], in_pld_tx_data[67], in_pld_tx_data[66], in_pld_tx_data[65], in_pld_tx_data[64], in_pld_tx_data[63], in_pld_tx_data[62], in_pld_tx_data[61], in_pld_tx_data[60], in_pld_tx_data[59], in_pld_tx_data[58], in_pld_tx_data[57], in_pld_tx_data[56], in_pld_tx_data[55], in_pld_tx_data[54], in_pld_tx_data[53], in_pld_tx_data[52], in_pld_tx_data[51], in_pld_tx_data[50], in_pld_tx_data[49], in_pld_tx_data[48], in_pld_tx_data[47], in_pld_tx_data[46], in_pld_tx_data[45], in_pld_tx_data[44], in_pld_tx_data[43], in_pld_tx_data[42], in_pld_tx_data[41], in_pld_tx_data[40], in_pld_tx_data[39], in_pld_tx_data[38], in_pld_tx_data[37], in_pld_tx_data[36], in_pld_tx_data[35], in_pld_tx_data[34], in_pld_tx_data[33], in_pld_tx_data[32], in_pld_tx_data[31], in_pld_tx_data[30], in_pld_tx_data[29], in_pld_tx_data[28], in_pld_tx_data[27], in_pld_tx_data[26], in_pld_tx_data[25], in_pld_tx_data[24], in_pld_tx_data[23], in_pld_tx_data[22], in_pld_tx_data[21], in_pld_tx_data[20], in_pld_tx_data[19], in_pld_tx_data[18], in_pld_tx_data[17], in_pld_tx_data[16], in_pld_tx_data[15], in_pld_tx_data[14], in_pld_tx_data[13], in_pld_tx_data[12], in_pld_tx_data[11], in_pld_tx_data[10], in_pld_tx_data[9], in_pld_tx_data[8], in_pld_tx_data[7], in_pld_tx_data[6], in_pld_tx_data[5], in_pld_tx_data[4], in_pld_tx_data[3], in_pld_tx_data[2], in_pld_tx_data[1], in_pld_tx_data[0]}),
				.pld_txelecidle(in_pld_txelecidle),
				.pld_uhsif_tx_clk(in_pld_uhsif_tx_clk),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.hip_clk_out_div_by_2_wire(),
				.hip_clk_out_wire(),
				.int_pldif_pmaif_tx_pld_clk(),
				.pld_10g_tx_burst_en_exe_10g_fastreg(),
				.pld_10g_tx_burst_en_exe_plddirect_reg(),
				.pld_10g_tx_data_valid_2ff_delay1_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay3_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg(),
				.pld_10g_tx_data_valid_fastreg(),
				.pld_10g_tx_data_valid_plddirect_fastreg(),
				.pld_pcs_tx_clk_out_pma_wire(),
				.pld_pma_tx_clk_out_wire(),
				.pld_pmaif_tx_pld_rst_n_reg(),
				.pld_polinv_tx_10g_pcsdirect_reg(),
				.pld_polinv_tx_8g_reg(),
				.pld_polinv_tx_pat_reg(),
				.pld_tx_clk_fifo(),
				.pld_tx_control_fifo(),
				.pld_tx_control_hi_10g_reg(),
				.pld_tx_control_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_10g_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_8g_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_control_lo_plddirect_fastreg(),
				.pld_tx_control_lo_plddirect_reg(),
				.pld_tx_data_hi_reg(),
				.pld_tx_data_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_10g_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_8g_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_data_lo_plddirect_fastreg(),
				.pld_tx_data_lo_plddirect_reg(),
				.pld_uhsif_reg(),
				.pma_tx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_hip_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6:0] = 7'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17:0] = 18'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8:0] = 9'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127:0] = 128'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4:0] = 5'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2:0] = 3'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_full = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_full_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out = 1'b0;
		end // if not generate
		
		//output assignments
		assign out_avmmreaddata_hssi_10g_rx_pcs = {w_hssi_10g_rx_pcs_avmmreaddata[7], w_hssi_10g_rx_pcs_avmmreaddata[6], w_hssi_10g_rx_pcs_avmmreaddata[5], w_hssi_10g_rx_pcs_avmmreaddata[4], w_hssi_10g_rx_pcs_avmmreaddata[3], w_hssi_10g_rx_pcs_avmmreaddata[2], w_hssi_10g_rx_pcs_avmmreaddata[1], w_hssi_10g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_10g_tx_pcs = {w_hssi_10g_tx_pcs_avmmreaddata[7], w_hssi_10g_tx_pcs_avmmreaddata[6], w_hssi_10g_tx_pcs_avmmreaddata[5], w_hssi_10g_tx_pcs_avmmreaddata[4], w_hssi_10g_tx_pcs_avmmreaddata[3], w_hssi_10g_tx_pcs_avmmreaddata[2], w_hssi_10g_tx_pcs_avmmreaddata[1], w_hssi_10g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_rx_pcs = {w_hssi_8g_rx_pcs_avmmreaddata[7], w_hssi_8g_rx_pcs_avmmreaddata[6], w_hssi_8g_rx_pcs_avmmreaddata[5], w_hssi_8g_rx_pcs_avmmreaddata[4], w_hssi_8g_rx_pcs_avmmreaddata[3], w_hssi_8g_rx_pcs_avmmreaddata[2], w_hssi_8g_rx_pcs_avmmreaddata[1], w_hssi_8g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_tx_pcs = {w_hssi_8g_tx_pcs_avmmreaddata[7], w_hssi_8g_tx_pcs_avmmreaddata[6], w_hssi_8g_tx_pcs_avmmreaddata[5], w_hssi_8g_tx_pcs_avmmreaddata[4], w_hssi_8g_tx_pcs_avmmreaddata[3], w_hssi_8g_tx_pcs_avmmreaddata[2], w_hssi_8g_tx_pcs_avmmreaddata[1], w_hssi_8g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pcs_pma_interface = {w_hssi_common_pcs_pma_interface_avmmreaddata[7], w_hssi_common_pcs_pma_interface_avmmreaddata[6], w_hssi_common_pcs_pma_interface_avmmreaddata[5], w_hssi_common_pcs_pma_interface_avmmreaddata[4], w_hssi_common_pcs_pma_interface_avmmreaddata[3], w_hssi_common_pcs_pma_interface_avmmreaddata[2], w_hssi_common_pcs_pma_interface_avmmreaddata[1], w_hssi_common_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pld_pcs_interface = {w_hssi_common_pld_pcs_interface_avmmreaddata[7], w_hssi_common_pld_pcs_interface_avmmreaddata[6], w_hssi_common_pld_pcs_interface_avmmreaddata[5], w_hssi_common_pld_pcs_interface_avmmreaddata[4], w_hssi_common_pld_pcs_interface_avmmreaddata[3], w_hssi_common_pld_pcs_interface_avmmreaddata[2], w_hssi_common_pld_pcs_interface_avmmreaddata[1], w_hssi_common_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_rx_pcs = {w_hssi_fifo_rx_pcs_avmmreaddata[7], w_hssi_fifo_rx_pcs_avmmreaddata[6], w_hssi_fifo_rx_pcs_avmmreaddata[5], w_hssi_fifo_rx_pcs_avmmreaddata[4], w_hssi_fifo_rx_pcs_avmmreaddata[3], w_hssi_fifo_rx_pcs_avmmreaddata[2], w_hssi_fifo_rx_pcs_avmmreaddata[1], w_hssi_fifo_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_tx_pcs = {w_hssi_fifo_tx_pcs_avmmreaddata[7], w_hssi_fifo_tx_pcs_avmmreaddata[6], w_hssi_fifo_tx_pcs_avmmreaddata[5], w_hssi_fifo_tx_pcs_avmmreaddata[4], w_hssi_fifo_tx_pcs_avmmreaddata[3], w_hssi_fifo_tx_pcs_avmmreaddata[2], w_hssi_fifo_tx_pcs_avmmreaddata[1], w_hssi_fifo_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_rx_pcs = {w_hssi_gen3_rx_pcs_avmmreaddata[7], w_hssi_gen3_rx_pcs_avmmreaddata[6], w_hssi_gen3_rx_pcs_avmmreaddata[5], w_hssi_gen3_rx_pcs_avmmreaddata[4], w_hssi_gen3_rx_pcs_avmmreaddata[3], w_hssi_gen3_rx_pcs_avmmreaddata[2], w_hssi_gen3_rx_pcs_avmmreaddata[1], w_hssi_gen3_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_tx_pcs = {w_hssi_gen3_tx_pcs_avmmreaddata[7], w_hssi_gen3_tx_pcs_avmmreaddata[6], w_hssi_gen3_tx_pcs_avmmreaddata[5], w_hssi_gen3_tx_pcs_avmmreaddata[4], w_hssi_gen3_tx_pcs_avmmreaddata[3], w_hssi_gen3_tx_pcs_avmmreaddata[2], w_hssi_gen3_tx_pcs_avmmreaddata[1], w_hssi_gen3_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_rx_pcs = {w_hssi_krfec_rx_pcs_avmmreaddata[7], w_hssi_krfec_rx_pcs_avmmreaddata[6], w_hssi_krfec_rx_pcs_avmmreaddata[5], w_hssi_krfec_rx_pcs_avmmreaddata[4], w_hssi_krfec_rx_pcs_avmmreaddata[3], w_hssi_krfec_rx_pcs_avmmreaddata[2], w_hssi_krfec_rx_pcs_avmmreaddata[1], w_hssi_krfec_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_tx_pcs = {w_hssi_krfec_tx_pcs_avmmreaddata[7], w_hssi_krfec_tx_pcs_avmmreaddata[6], w_hssi_krfec_tx_pcs_avmmreaddata[5], w_hssi_krfec_tx_pcs_avmmreaddata[4], w_hssi_krfec_tx_pcs_avmmreaddata[3], w_hssi_krfec_tx_pcs_avmmreaddata[2], w_hssi_krfec_tx_pcs_avmmreaddata[1], w_hssi_krfec_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen1_2 = {w_hssi_pipe_gen1_2_avmmreaddata[7], w_hssi_pipe_gen1_2_avmmreaddata[6], w_hssi_pipe_gen1_2_avmmreaddata[5], w_hssi_pipe_gen1_2_avmmreaddata[4], w_hssi_pipe_gen1_2_avmmreaddata[3], w_hssi_pipe_gen1_2_avmmreaddata[2], w_hssi_pipe_gen1_2_avmmreaddata[1], w_hssi_pipe_gen1_2_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen3 = {w_hssi_pipe_gen3_avmmreaddata[7], w_hssi_pipe_gen3_avmmreaddata[6], w_hssi_pipe_gen3_avmmreaddata[5], w_hssi_pipe_gen3_avmmreaddata[4], w_hssi_pipe_gen3_avmmreaddata[3], w_hssi_pipe_gen3_avmmreaddata[2], w_hssi_pipe_gen3_avmmreaddata[1], w_hssi_pipe_gen3_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pcs_pma_interface = {w_hssi_rx_pcs_pma_interface_avmmreaddata[7], w_hssi_rx_pcs_pma_interface_avmmreaddata[6], w_hssi_rx_pcs_pma_interface_avmmreaddata[5], w_hssi_rx_pcs_pma_interface_avmmreaddata[4], w_hssi_rx_pcs_pma_interface_avmmreaddata[3], w_hssi_rx_pcs_pma_interface_avmmreaddata[2], w_hssi_rx_pcs_pma_interface_avmmreaddata[1], w_hssi_rx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pld_pcs_interface = {w_hssi_rx_pld_pcs_interface_avmmreaddata[7], w_hssi_rx_pld_pcs_interface_avmmreaddata[6], w_hssi_rx_pld_pcs_interface_avmmreaddata[5], w_hssi_rx_pld_pcs_interface_avmmreaddata[4], w_hssi_rx_pld_pcs_interface_avmmreaddata[3], w_hssi_rx_pld_pcs_interface_avmmreaddata[2], w_hssi_rx_pld_pcs_interface_avmmreaddata[1], w_hssi_rx_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pcs_pma_interface = {w_hssi_tx_pcs_pma_interface_avmmreaddata[7], w_hssi_tx_pcs_pma_interface_avmmreaddata[6], w_hssi_tx_pcs_pma_interface_avmmreaddata[5], w_hssi_tx_pcs_pma_interface_avmmreaddata[4], w_hssi_tx_pcs_pma_interface_avmmreaddata[3], w_hssi_tx_pcs_pma_interface_avmmreaddata[2], w_hssi_tx_pcs_pma_interface_avmmreaddata[1], w_hssi_tx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pld_pcs_interface = {w_hssi_tx_pld_pcs_interface_avmmreaddata[7], w_hssi_tx_pld_pcs_interface_avmmreaddata[6], w_hssi_tx_pld_pcs_interface_avmmreaddata[5], w_hssi_tx_pld_pcs_interface_avmmreaddata[4], w_hssi_tx_pld_pcs_interface_avmmreaddata[3], w_hssi_tx_pld_pcs_interface_avmmreaddata[2], w_hssi_tx_pld_pcs_interface_avmmreaddata[1], w_hssi_tx_pld_pcs_interface_avmmreaddata[0]};
		assign out_blockselect_hssi_10g_rx_pcs = w_hssi_10g_rx_pcs_blockselect;
		assign out_blockselect_hssi_10g_tx_pcs = w_hssi_10g_tx_pcs_blockselect;
		assign out_blockselect_hssi_8g_rx_pcs = w_hssi_8g_rx_pcs_blockselect;
		assign out_blockselect_hssi_8g_tx_pcs = w_hssi_8g_tx_pcs_blockselect;
		assign out_blockselect_hssi_common_pcs_pma_interface = w_hssi_common_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_common_pld_pcs_interface = w_hssi_common_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_fifo_rx_pcs = w_hssi_fifo_rx_pcs_blockselect;
		assign out_blockselect_hssi_fifo_tx_pcs = w_hssi_fifo_tx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_rx_pcs = w_hssi_gen3_rx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_tx_pcs = w_hssi_gen3_tx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_rx_pcs = w_hssi_krfec_rx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_tx_pcs = w_hssi_krfec_tx_pcs_blockselect;
		assign out_blockselect_hssi_pipe_gen1_2 = w_hssi_pipe_gen1_2_blockselect;
		assign out_blockselect_hssi_pipe_gen3 = w_hssi_pipe_gen3_blockselect;
		assign out_blockselect_hssi_rx_pcs_pma_interface = w_hssi_rx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_rx_pld_pcs_interface = w_hssi_rx_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_tx_pcs_pma_interface = w_hssi_tx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_tx_pld_pcs_interface = w_hssi_tx_pld_pcs_interface_blockselect;
		assign out_bond_pcs10g_out_bot = {w_hssi_10g_tx_pcs_distdwn_out_rden, w_hssi_10g_tx_pcs_distdwn_out_wren, w_hssi_10g_tx_pcs_distdwn_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs10g_out_top = {w_hssi_10g_tx_pcs_distup_out_rden, w_hssi_10g_tx_pcs_distup_out_wren, w_hssi_10g_tx_pcs_distup_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs8g_out_bot = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down, w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_down, w_hssi_8g_tx_pcs_wr_enable_out_chnl_down, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_down, w_hssi_8g_rx_pcs_wr_enable_out_chnl_down, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[0]};
		assign out_bond_pcs8g_out_top = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up, w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_up, w_hssi_8g_tx_pcs_wr_enable_out_chnl_up, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_up, w_hssi_8g_rx_pcs_wr_enable_out_chnl_up, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[0]};
		assign out_bond_pmaif_out_bot = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[0]};
		assign out_bond_pmaif_out_top = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[0]};
		assign out_hip_clk_out = {w_hssi_common_pld_pcs_interface_hip_cmn_clk[1], w_hssi_common_pld_pcs_interface_hip_cmn_clk[0], w_hssi_tx_pld_pcs_interface_hip_tx_clk};
		assign out_hip_ctrl_out = {w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[4], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[3], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[2], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[1], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[0], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[0]};
		assign out_hip_iocsr_rdy = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
		assign out_hip_iocsr_rdy_dly = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
		assign out_hip_nfrzdrv = w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
		assign out_hip_npor = w_hssi_common_pld_pcs_interface_hip_npor;
		assign out_hip_rx_data = {w_hssi_rx_pld_pcs_interface_hip_rx_data[50], w_hssi_rx_pld_pcs_interface_hip_rx_data[49], w_hssi_rx_pld_pcs_interface_hip_rx_data[48], w_hssi_rx_pld_pcs_interface_hip_rx_data[47], w_hssi_rx_pld_pcs_interface_hip_rx_data[46], w_hssi_rx_pld_pcs_interface_hip_rx_data[45], w_hssi_rx_pld_pcs_interface_hip_rx_data[44], w_hssi_rx_pld_pcs_interface_hip_rx_data[43], w_hssi_rx_pld_pcs_interface_hip_rx_data[42], w_hssi_rx_pld_pcs_interface_hip_rx_data[41], w_hssi_rx_pld_pcs_interface_hip_rx_data[40], w_hssi_rx_pld_pcs_interface_hip_rx_data[39], w_hssi_rx_pld_pcs_interface_hip_rx_data[38], w_hssi_rx_pld_pcs_interface_hip_rx_data[37], w_hssi_rx_pld_pcs_interface_hip_rx_data[36], w_hssi_rx_pld_pcs_interface_hip_rx_data[35], w_hssi_rx_pld_pcs_interface_hip_rx_data[34], w_hssi_rx_pld_pcs_interface_hip_rx_data[33], w_hssi_rx_pld_pcs_interface_hip_rx_data[32], w_hssi_rx_pld_pcs_interface_hip_rx_data[31], w_hssi_rx_pld_pcs_interface_hip_rx_data[30], w_hssi_rx_pld_pcs_interface_hip_rx_data[29], w_hssi_rx_pld_pcs_interface_hip_rx_data[28], w_hssi_rx_pld_pcs_interface_hip_rx_data[27], w_hssi_rx_pld_pcs_interface_hip_rx_data[26], w_hssi_rx_pld_pcs_interface_hip_rx_data[25], w_hssi_rx_pld_pcs_interface_hip_rx_data[24], w_hssi_rx_pld_pcs_interface_hip_rx_data[23], w_hssi_rx_pld_pcs_interface_hip_rx_data[22], w_hssi_rx_pld_pcs_interface_hip_rx_data[21], w_hssi_rx_pld_pcs_interface_hip_rx_data[20], w_hssi_rx_pld_pcs_interface_hip_rx_data[19], w_hssi_rx_pld_pcs_interface_hip_rx_data[18], w_hssi_rx_pld_pcs_interface_hip_rx_data[17], w_hssi_rx_pld_pcs_interface_hip_rx_data[16], w_hssi_rx_pld_pcs_interface_hip_rx_data[15], w_hssi_rx_pld_pcs_interface_hip_rx_data[14], w_hssi_rx_pld_pcs_interface_hip_rx_data[13], w_hssi_rx_pld_pcs_interface_hip_rx_data[12], w_hssi_rx_pld_pcs_interface_hip_rx_data[11], w_hssi_rx_pld_pcs_interface_hip_rx_data[10], w_hssi_rx_pld_pcs_interface_hip_rx_data[9], w_hssi_rx_pld_pcs_interface_hip_rx_data[8], w_hssi_rx_pld_pcs_interface_hip_rx_data[7], w_hssi_rx_pld_pcs_interface_hip_rx_data[6], w_hssi_rx_pld_pcs_interface_hip_rx_data[5], w_hssi_rx_pld_pcs_interface_hip_rx_data[4], w_hssi_rx_pld_pcs_interface_hip_rx_data[3], w_hssi_rx_pld_pcs_interface_hip_rx_data[2], w_hssi_rx_pld_pcs_interface_hip_rx_data[1], w_hssi_rx_pld_pcs_interface_hip_rx_data[0]};
		assign out_hip_usermode = w_hssi_common_pld_pcs_interface_hip_usermode;
		assign out_pld_10g_krfec_rx_blk_lock = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
		assign out_pld_10g_krfec_rx_diag_data_status = {w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1], w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[0]};
		assign out_pld_10g_krfec_rx_frame = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
		assign out_pld_10g_krfec_tx_frame = w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
		assign out_pld_10g_rx_align_val = w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
		assign out_pld_10g_rx_crc32_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
		assign out_pld_10g_rx_data_valid = w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
		assign out_pld_10g_rx_empty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
		assign out_pld_10g_rx_fifo_del = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
		assign out_pld_10g_rx_fifo_insert = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
		assign out_pld_10g_rx_fifo_num = {w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[3], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[2], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[1], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[0]};
		assign out_pld_10g_rx_frame_lock = w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
		assign out_pld_10g_rx_hi_ber = w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
		assign out_pld_10g_rx_oflw_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
		assign out_pld_10g_rx_pempty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
		assign out_pld_10g_rx_pfull = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
		assign out_pld_10g_tx_burst_en_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
		assign out_pld_10g_tx_empty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
		assign out_pld_10g_tx_fifo_num = {w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[2], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[1], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[0]};
		assign out_pld_10g_tx_full = w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
		assign out_pld_10g_tx_pempty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
		assign out_pld_10g_tx_pfull = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
		assign out_pld_10g_tx_wordslip_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
		assign out_pld_8g_a1a2_k1k2_flag = {w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[2], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[1], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[0]};
		assign out_pld_8g_empty_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
		assign out_pld_8g_empty_rx = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
		assign out_pld_8g_empty_tx = w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
		assign out_pld_8g_full_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
		assign out_pld_8g_full_rx = w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
		assign out_pld_8g_full_tx = w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
		assign out_pld_8g_rxelecidle = w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
		assign out_pld_8g_signal_detect_out = w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
		assign out_pld_8g_wa_boundary = {w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0]};
		assign out_pld_krfec_tx_alignment = w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
		assign out_pld_pcs_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
		assign out_pld_pcs_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
		assign out_pld_pma_adapt_done = w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
		assign out_pld_pma_clkdiv_rx_user = w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
		assign out_pld_pma_clkdiv_tx_user = w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
		assign out_pld_pma_clklow = w_hssi_common_pld_pcs_interface_pld_pma_clklow;
		assign out_pld_pma_fref = w_hssi_common_pld_pcs_interface_pld_pma_fref;
		assign out_pld_pma_hclk = w_hssi_common_pld_pcs_interface_pld_pma_hclk;
		assign out_pld_pma_pcie_sw_done = {w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1], w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[0]};
		assign out_pld_pma_pfdmode_lock = w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
		assign out_pld_pma_reserved_in = {w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[3], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[2], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[1], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[0]};
		assign out_pld_pma_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
		assign out_pld_pma_rx_detect_valid = w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
		assign out_pld_pma_rx_found = w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
		assign out_pld_pma_rxpll_lock = w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
		assign out_pld_pma_signal_ok = w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
		assign out_pld_pma_testbus = {w_hssi_common_pld_pcs_interface_pld_pma_testbus[7], w_hssi_common_pld_pcs_interface_pld_pma_testbus[6], w_hssi_common_pld_pcs_interface_pld_pma_testbus[5], w_hssi_common_pld_pcs_interface_pld_pma_testbus[4], w_hssi_common_pld_pcs_interface_pld_pma_testbus[3], w_hssi_common_pld_pcs_interface_pld_pma_testbus[2], w_hssi_common_pld_pcs_interface_pld_pma_testbus[1], w_hssi_common_pld_pcs_interface_pld_pma_testbus[0]};
		assign out_pld_pma_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
		assign out_pld_pmaif_mask_tx_pll = w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
		assign out_pld_reserved_out = {w_hssi_common_pld_pcs_interface_pld_reserved_out[9], w_hssi_common_pld_pcs_interface_pld_reserved_out[8], w_hssi_common_pld_pcs_interface_pld_reserved_out[7], w_hssi_common_pld_pcs_interface_pld_reserved_out[6], w_hssi_common_pld_pcs_interface_pld_reserved_out[5], w_hssi_common_pld_pcs_interface_pld_reserved_out[4], w_hssi_common_pld_pcs_interface_pld_reserved_out[3], w_hssi_common_pld_pcs_interface_pld_reserved_out[2], w_hssi_common_pld_pcs_interface_pld_reserved_out[1], w_hssi_common_pld_pcs_interface_pld_reserved_out[0]};
		assign out_pld_rx_control = {w_hssi_rx_pld_pcs_interface_pld_rx_control[19], w_hssi_rx_pld_pcs_interface_pld_rx_control[18], w_hssi_rx_pld_pcs_interface_pld_rx_control[17], w_hssi_rx_pld_pcs_interface_pld_rx_control[16], w_hssi_rx_pld_pcs_interface_pld_rx_control[15], w_hssi_rx_pld_pcs_interface_pld_rx_control[14], w_hssi_rx_pld_pcs_interface_pld_rx_control[13], w_hssi_rx_pld_pcs_interface_pld_rx_control[12], w_hssi_rx_pld_pcs_interface_pld_rx_control[11], w_hssi_rx_pld_pcs_interface_pld_rx_control[10], w_hssi_rx_pld_pcs_interface_pld_rx_control[9], w_hssi_rx_pld_pcs_interface_pld_rx_control[8], w_hssi_rx_pld_pcs_interface_pld_rx_control[7], w_hssi_rx_pld_pcs_interface_pld_rx_control[6], w_hssi_rx_pld_pcs_interface_pld_rx_control[5], w_hssi_rx_pld_pcs_interface_pld_rx_control[4], w_hssi_rx_pld_pcs_interface_pld_rx_control[3], w_hssi_rx_pld_pcs_interface_pld_rx_control[2], w_hssi_rx_pld_pcs_interface_pld_rx_control[1], w_hssi_rx_pld_pcs_interface_pld_rx_control[0]};
		assign out_pld_rx_data = {w_hssi_rx_pld_pcs_interface_pld_rx_data[127], w_hssi_rx_pld_pcs_interface_pld_rx_data[126], w_hssi_rx_pld_pcs_interface_pld_rx_data[125], w_hssi_rx_pld_pcs_interface_pld_rx_data[124], w_hssi_rx_pld_pcs_interface_pld_rx_data[123], w_hssi_rx_pld_pcs_interface_pld_rx_data[122], w_hssi_rx_pld_pcs_interface_pld_rx_data[121], w_hssi_rx_pld_pcs_interface_pld_rx_data[120], w_hssi_rx_pld_pcs_interface_pld_rx_data[119], w_hssi_rx_pld_pcs_interface_pld_rx_data[118], w_hssi_rx_pld_pcs_interface_pld_rx_data[117], w_hssi_rx_pld_pcs_interface_pld_rx_data[116], w_hssi_rx_pld_pcs_interface_pld_rx_data[115], w_hssi_rx_pld_pcs_interface_pld_rx_data[114], w_hssi_rx_pld_pcs_interface_pld_rx_data[113], w_hssi_rx_pld_pcs_interface_pld_rx_data[112], w_hssi_rx_pld_pcs_interface_pld_rx_data[111], w_hssi_rx_pld_pcs_interface_pld_rx_data[110], w_hssi_rx_pld_pcs_interface_pld_rx_data[109], w_hssi_rx_pld_pcs_interface_pld_rx_data[108], w_hssi_rx_pld_pcs_interface_pld_rx_data[107], w_hssi_rx_pld_pcs_interface_pld_rx_data[106], w_hssi_rx_pld_pcs_interface_pld_rx_data[105], w_hssi_rx_pld_pcs_interface_pld_rx_data[104], w_hssi_rx_pld_pcs_interface_pld_rx_data[103], w_hssi_rx_pld_pcs_interface_pld_rx_data[102], w_hssi_rx_pld_pcs_interface_pld_rx_data[101], w_hssi_rx_pld_pcs_interface_pld_rx_data[100], w_hssi_rx_pld_pcs_interface_pld_rx_data[99], w_hssi_rx_pld_pcs_interface_pld_rx_data[98], w_hssi_rx_pld_pcs_interface_pld_rx_data[97], w_hssi_rx_pld_pcs_interface_pld_rx_data[96], w_hssi_rx_pld_pcs_interface_pld_rx_data[95], w_hssi_rx_pld_pcs_interface_pld_rx_data[94], w_hssi_rx_pld_pcs_interface_pld_rx_data[93], w_hssi_rx_pld_pcs_interface_pld_rx_data[92], w_hssi_rx_pld_pcs_interface_pld_rx_data[91], w_hssi_rx_pld_pcs_interface_pld_rx_data[90], w_hssi_rx_pld_pcs_interface_pld_rx_data[89], w_hssi_rx_pld_pcs_interface_pld_rx_data[88], w_hssi_rx_pld_pcs_interface_pld_rx_data[87], w_hssi_rx_pld_pcs_interface_pld_rx_data[86], w_hssi_rx_pld_pcs_interface_pld_rx_data[85], w_hssi_rx_pld_pcs_interface_pld_rx_data[84], w_hssi_rx_pld_pcs_interface_pld_rx_data[83], w_hssi_rx_pld_pcs_interface_pld_rx_data[82], w_hssi_rx_pld_pcs_interface_pld_rx_data[81], w_hssi_rx_pld_pcs_interface_pld_rx_data[80], w_hssi_rx_pld_pcs_interface_pld_rx_data[79], w_hssi_rx_pld_pcs_interface_pld_rx_data[78], w_hssi_rx_pld_pcs_interface_pld_rx_data[77], w_hssi_rx_pld_pcs_interface_pld_rx_data[76], w_hssi_rx_pld_pcs_interface_pld_rx_data[75], w_hssi_rx_pld_pcs_interface_pld_rx_data[74], w_hssi_rx_pld_pcs_interface_pld_rx_data[73], w_hssi_rx_pld_pcs_interface_pld_rx_data[72], w_hssi_rx_pld_pcs_interface_pld_rx_data[71], w_hssi_rx_pld_pcs_interface_pld_rx_data[70], w_hssi_rx_pld_pcs_interface_pld_rx_data[69], w_hssi_rx_pld_pcs_interface_pld_rx_data[68], w_hssi_rx_pld_pcs_interface_pld_rx_data[67], w_hssi_rx_pld_pcs_interface_pld_rx_data[66], w_hssi_rx_pld_pcs_interface_pld_rx_data[65], w_hssi_rx_pld_pcs_interface_pld_rx_data[64], w_hssi_rx_pld_pcs_interface_pld_rx_data[63], w_hssi_rx_pld_pcs_interface_pld_rx_data[62], w_hssi_rx_pld_pcs_interface_pld_rx_data[61], w_hssi_rx_pld_pcs_interface_pld_rx_data[60], w_hssi_rx_pld_pcs_interface_pld_rx_data[59], w_hssi_rx_pld_pcs_interface_pld_rx_data[58], w_hssi_rx_pld_pcs_interface_pld_rx_data[57], w_hssi_rx_pld_pcs_interface_pld_rx_data[56], w_hssi_rx_pld_pcs_interface_pld_rx_data[55], w_hssi_rx_pld_pcs_interface_pld_rx_data[54], w_hssi_rx_pld_pcs_interface_pld_rx_data[53], w_hssi_rx_pld_pcs_interface_pld_rx_data[52], w_hssi_rx_pld_pcs_interface_pld_rx_data[51], w_hssi_rx_pld_pcs_interface_pld_rx_data[50], w_hssi_rx_pld_pcs_interface_pld_rx_data[49], w_hssi_rx_pld_pcs_interface_pld_rx_data[48], w_hssi_rx_pld_pcs_interface_pld_rx_data[47], w_hssi_rx_pld_pcs_interface_pld_rx_data[46], w_hssi_rx_pld_pcs_interface_pld_rx_data[45], w_hssi_rx_pld_pcs_interface_pld_rx_data[44], w_hssi_rx_pld_pcs_interface_pld_rx_data[43], w_hssi_rx_pld_pcs_interface_pld_rx_data[42], w_hssi_rx_pld_pcs_interface_pld_rx_data[41], w_hssi_rx_pld_pcs_interface_pld_rx_data[40], w_hssi_rx_pld_pcs_interface_pld_rx_data[39], w_hssi_rx_pld_pcs_interface_pld_rx_data[38], w_hssi_rx_pld_pcs_interface_pld_rx_data[37], w_hssi_rx_pld_pcs_interface_pld_rx_data[36], w_hssi_rx_pld_pcs_interface_pld_rx_data[35], w_hssi_rx_pld_pcs_interface_pld_rx_data[34], w_hssi_rx_pld_pcs_interface_pld_rx_data[33], w_hssi_rx_pld_pcs_interface_pld_rx_data[32], w_hssi_rx_pld_pcs_interface_pld_rx_data[31], w_hssi_rx_pld_pcs_interface_pld_rx_data[30], w_hssi_rx_pld_pcs_interface_pld_rx_data[29], w_hssi_rx_pld_pcs_interface_pld_rx_data[28], w_hssi_rx_pld_pcs_interface_pld_rx_data[27], w_hssi_rx_pld_pcs_interface_pld_rx_data[26], w_hssi_rx_pld_pcs_interface_pld_rx_data[25], w_hssi_rx_pld_pcs_interface_pld_rx_data[24], w_hssi_rx_pld_pcs_interface_pld_rx_data[23], w_hssi_rx_pld_pcs_interface_pld_rx_data[22], w_hssi_rx_pld_pcs_interface_pld_rx_data[21], w_hssi_rx_pld_pcs_interface_pld_rx_data[20], w_hssi_rx_pld_pcs_interface_pld_rx_data[19], w_hssi_rx_pld_pcs_interface_pld_rx_data[18], w_hssi_rx_pld_pcs_interface_pld_rx_data[17], w_hssi_rx_pld_pcs_interface_pld_rx_data[16], w_hssi_rx_pld_pcs_interface_pld_rx_data[15], w_hssi_rx_pld_pcs_interface_pld_rx_data[14], w_hssi_rx_pld_pcs_interface_pld_rx_data[13], w_hssi_rx_pld_pcs_interface_pld_rx_data[12], w_hssi_rx_pld_pcs_interface_pld_rx_data[11], w_hssi_rx_pld_pcs_interface_pld_rx_data[10], w_hssi_rx_pld_pcs_interface_pld_rx_data[9], w_hssi_rx_pld_pcs_interface_pld_rx_data[8], w_hssi_rx_pld_pcs_interface_pld_rx_data[7], w_hssi_rx_pld_pcs_interface_pld_rx_data[6], w_hssi_rx_pld_pcs_interface_pld_rx_data[5], w_hssi_rx_pld_pcs_interface_pld_rx_data[4], w_hssi_rx_pld_pcs_interface_pld_rx_data[3], w_hssi_rx_pld_pcs_interface_pld_rx_data[2], w_hssi_rx_pld_pcs_interface_pld_rx_data[1], w_hssi_rx_pld_pcs_interface_pld_rx_data[0]};
		assign out_pld_rx_prbs_done = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
		assign out_pld_rx_prbs_err = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
		assign out_pld_test_data = {w_hssi_common_pld_pcs_interface_pld_test_data[19], w_hssi_common_pld_pcs_interface_pld_test_data[18], w_hssi_common_pld_pcs_interface_pld_test_data[17], w_hssi_common_pld_pcs_interface_pld_test_data[16], w_hssi_common_pld_pcs_interface_pld_test_data[15], w_hssi_common_pld_pcs_interface_pld_test_data[14], w_hssi_common_pld_pcs_interface_pld_test_data[13], w_hssi_common_pld_pcs_interface_pld_test_data[12], w_hssi_common_pld_pcs_interface_pld_test_data[11], w_hssi_common_pld_pcs_interface_pld_test_data[10], w_hssi_common_pld_pcs_interface_pld_test_data[9], w_hssi_common_pld_pcs_interface_pld_test_data[8], w_hssi_common_pld_pcs_interface_pld_test_data[7], w_hssi_common_pld_pcs_interface_pld_test_data[6], w_hssi_common_pld_pcs_interface_pld_test_data[5], w_hssi_common_pld_pcs_interface_pld_test_data[4], w_hssi_common_pld_pcs_interface_pld_test_data[3], w_hssi_common_pld_pcs_interface_pld_test_data[2], w_hssi_common_pld_pcs_interface_pld_test_data[1], w_hssi_common_pld_pcs_interface_pld_test_data[0]};
		assign out_pld_uhsif_lock = w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
		assign out_pld_uhsif_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
		assign out_pma_adapt_start = w_hssi_common_pcs_pma_interface_pma_adapt_start;
		assign out_pma_atpg_los_en_n = w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
		assign out_pma_csr_test_dis = w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
		assign out_pma_current_coeff = {w_hssi_common_pcs_pma_interface_pma_current_coeff[17], w_hssi_common_pcs_pma_interface_pma_current_coeff[16], w_hssi_common_pcs_pma_interface_pma_current_coeff[15], w_hssi_common_pcs_pma_interface_pma_current_coeff[14], w_hssi_common_pcs_pma_interface_pma_current_coeff[13], w_hssi_common_pcs_pma_interface_pma_current_coeff[12], w_hssi_common_pcs_pma_interface_pma_current_coeff[11], w_hssi_common_pcs_pma_interface_pma_current_coeff[10], w_hssi_common_pcs_pma_interface_pma_current_coeff[9], w_hssi_common_pcs_pma_interface_pma_current_coeff[8], w_hssi_common_pcs_pma_interface_pma_current_coeff[7], w_hssi_common_pcs_pma_interface_pma_current_coeff[6], w_hssi_common_pcs_pma_interface_pma_current_coeff[5], w_hssi_common_pcs_pma_interface_pma_current_coeff[4], w_hssi_common_pcs_pma_interface_pma_current_coeff[3], w_hssi_common_pcs_pma_interface_pma_current_coeff[2], w_hssi_common_pcs_pma_interface_pma_current_coeff[1], w_hssi_common_pcs_pma_interface_pma_current_coeff[0]};
		assign out_pma_current_rxpreset = {w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[1], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[0]};
		assign out_pma_early_eios = w_hssi_common_pcs_pma_interface_pma_early_eios;
		assign out_pma_eye_monitor = {w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0]};
		assign out_pma_interface_select = {w_hssi_common_pcs_pma_interface_pma_interface_select[1], w_hssi_common_pcs_pma_interface_pma_interface_select[0]};
		assign out_pma_ltd_b = w_hssi_common_pcs_pma_interface_pma_ltd_b;
		assign out_pma_ltr = w_hssi_common_pcs_pma_interface_pma_ltr;
		assign out_pma_nfrzdrv = w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
		assign out_pma_nrpi_freeze = w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
		assign out_pma_pcie_switch = {w_hssi_common_pcs_pma_interface_pma_pcie_switch[1], w_hssi_common_pcs_pma_interface_pma_pcie_switch[0]};
		assign out_pma_ppm_lock = w_hssi_common_pcs_pma_interface_pma_ppm_lock;
		assign out_pma_reserved_out = {w_hssi_common_pcs_pma_interface_pma_reserved_out[4], w_hssi_common_pcs_pma_interface_pma_reserved_out[3], w_hssi_common_pcs_pma_interface_pma_reserved_out[2], w_hssi_common_pcs_pma_interface_pma_reserved_out[1], w_hssi_common_pcs_pma_interface_pma_reserved_out[0]};
		assign out_pma_rs_lpbk_b = w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
		assign out_pma_rx_clkslip = w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
		assign out_pma_rx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
		assign out_pma_rxpma_rstb = w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
		assign out_pma_scan_mode_n = w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
		assign out_pma_scan_shift_n = w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
		assign out_pma_tx_bitslip = w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
		assign out_pma_tx_bonding_rstb = w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
		assign out_pma_tx_elec_idle = w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
		assign out_pma_tx_pma_data = {w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0]};
		assign out_pma_tx_qpi_pulldn = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
		assign out_pma_tx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
		assign out_pma_tx_txdetectrx = w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
		assign out_pma_txpma_rstb = w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	endgenerate
endmodule
module twentynm_pcs_rev_20nm5es2
	#(
	//PARAM_LIST_START
		parameter xcvr_native_mode = "mode_duplex",  // mode_duplex, mode_rx_only, mode_tx_only
		
		// parameters for twentynm_hssi_10g_rx_pcs
		parameter hssi_10g_rx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_align_del = "align_del_en", // align_del_dis|align_del_en
		parameter hssi_10g_rx_pcs_ber_bit_err_total_cnt = "bit_err_total_cnt_10g", // bit_err_total_cnt_10g
		parameter hssi_10g_rx_pcs_ber_clken = "ber_clk_dis", // ber_clk_dis|ber_clk_en
		parameter hssi_10g_rx_pcs_ber_xus_timer_window = 21'b100110001001010,
		parameter hssi_10g_rx_pcs_bitslip_mode = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_rx_pcs_blksync_bitslip_type = "bitslip_comb", // bitslip_comb|bitslip_reg
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_cnt = 3'b1,
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_type = "bitslip_match", // bitslip_match|bitslip_cnt
		parameter hssi_10g_rx_pcs_blksync_bypass = "blksync_bypass_dis", // blksync_bypass_dis|blksync_bypass_en
		parameter hssi_10g_rx_pcs_blksync_clken = "blksync_clk_dis", // blksync_clk_dis|blksync_clk_en
		parameter hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt = "enum_invalid_sh_cnt_10g", // enum_invalid_sh_cnt_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock = "knum_sh_cnt_postlock_10g", // knum_sh_cnt_postlock_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock = "knum_sh_cnt_prelock_10g", // knum_sh_cnt_prelock_10g
		parameter hssi_10g_rx_pcs_blksync_pipeln = "blksync_pipeln_dis", // blksync_pipeln_dis|blksync_pipeln_en
		parameter hssi_10g_rx_pcs_clr_errblk_cnt_en = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_control_del = "control_del_all", // control_del_all|control_del_none
		parameter hssi_10g_rx_pcs_crcchk_bypass = "crcchk_bypass_dis", // crcchk_bypass_dis|crcchk_bypass_en
		parameter hssi_10g_rx_pcs_crcchk_clken = "crcchk_clk_dis", // crcchk_clk_dis|crcchk_clk_en
		parameter hssi_10g_rx_pcs_crcchk_inv = "crcchk_inv_dis", // crcchk_inv_dis|crcchk_inv_en
		parameter hssi_10g_rx_pcs_crcchk_pipeln = "crcchk_pipeln_dis", // crcchk_pipeln_dis|crcchk_pipeln_en
		parameter hssi_10g_rx_pcs_crcflag_pipeln = "crcflag_pipeln_dis", // crcflag_pipeln_dis|crcflag_pipeln_en
		parameter hssi_10g_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_rx_pcs_dec64b66b_clken = "dec64b66b_clk_dis", // dec64b66b_clk_dis|dec64b66b_clk_en
		parameter hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass = "dec_64b66b_rxsm_bypass_dis", // dec_64b66b_rxsm_bypass_dis|dec_64b66b_rxsm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_bypass = "descrm_bypass_en", // descrm_bypass_dis|descrm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_clken = "descrm_clk_dis", // descrm_clk_dis|descrm_clk_en
		parameter hssi_10g_rx_pcs_descrm_mode = "async", // async|sync
		parameter hssi_10g_rx_pcs_descrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_dft_clk_out_sel = "rx_master_clk", // rx_master_clk|rx_gbexp_clk|rx_blksync_clk|rx_descrm_clk|rx_frmsync_clk|rx_64b66bdec_clk|rx_ber_clk|rx_rand_clk|rx_crcchk_clk|rx_wrfifo_clk|rx_rdfifo_clk|rx_fec_clk
		parameter hssi_10g_rx_pcs_dis_signal_ok = "dis_signal_ok_dis", // dis_signal_ok_dis|dis_signal_ok_en
		parameter hssi_10g_rx_pcs_dispchk_bypass = "dispchk_bypass_dis", // dispchk_bypass_dis|dispchk_bypass_en
		parameter hssi_10g_rx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_rx_pcs_fast_path = "fast_path_dis", // fast_path_dis|fast_path_en
		parameter hssi_10g_rx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_rx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_rx_pcs_fifo_double_read = "fifo_double_read_dis", // fifo_double_read_dis|fifo_double_read_en
		parameter hssi_10g_rx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_rx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_rx_pcs_force_align = "force_align_dis", // force_align_dis|force_align_en
		parameter hssi_10g_rx_pcs_frmsync_bypass = "frmsync_bypass_dis", // frmsync_bypass_dis|frmsync_bypass_en
		parameter hssi_10g_rx_pcs_frmsync_clken = "frmsync_clk_dis", // frmsync_clk_dis|frmsync_clk_en
		parameter hssi_10g_rx_pcs_frmsync_enum_scrm = "enum_scrm_default", // enum_scrm_default
		parameter hssi_10g_rx_pcs_frmsync_enum_sync = "enum_sync_default", // enum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_flag_type = "all_framing_words", // all_framing_words|location_only
		parameter hssi_10g_rx_pcs_frmsync_knum_sync = "knum_sync_default", // knum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_mfrm_length = 16'b100000000000,
		parameter hssi_10g_rx_pcs_frmsync_pipeln = "frmsync_pipeln_dis", // frmsync_pipeln_dis|frmsync_pipeln_en
		parameter hssi_10g_rx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_rx_pcs_gb_rx_idwidth = "width_32", // width_40|width_32|width_64
		parameter hssi_10g_rx_pcs_gb_rx_odwidth = "width_66", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_rx_pcs_gbexp_clken = "gbexp_clk_dis", // gbexp_clk_dis|gbexp_clk_en
		parameter hssi_10g_rx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_10g_rx_pcs_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_rx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_rx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_rx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_rx_pcs_pld_if_type = "fifo", // fifo|reg
		parameter hssi_10g_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_rx_pcs_rand_clken = "rand_clk_dis", // rand_clk_dis|rand_clk_en
		parameter hssi_10g_rx_pcs_rd_clk_sel = "rd_rx_pma_clk", // rd_rx_pld_clk|rd_rx_pma_clk|rd_refclk_dig
		parameter hssi_10g_rx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_rx_pcs_rx_fifo_write_ctrl = "blklock_stops", // blklock_stops|blklock_ignore
		parameter hssi_10g_rx_pcs_rx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_rx_pcs_rx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_rx_pcs_rx_signal_ok_sel = "synchronized_ver", // synchronized_ver|nonsync_ver
		parameter hssi_10g_rx_pcs_rx_sm_bypass = "rx_sm_bypass_dis", // rx_sm_bypass_dis|rx_sm_bypass_en
		parameter hssi_10g_rx_pcs_rx_sm_hiber = "rx_sm_hiber_en", // rx_sm_hiber_en|rx_sm_hiber_dis
		parameter hssi_10g_rx_pcs_rx_sm_pipeln = "rx_sm_pipeln_dis", // rx_sm_pipeln_dis|rx_sm_pipeln_en
		parameter hssi_10g_rx_pcs_rx_testbus_sel = "crc32_chk_testbus1", // crc32_chk_testbus1|crc32_chk_testbus2|frame_sync_testbus1|frame_sync_testbus2|dec64b66b_testbus|rxsm_testbus|ber_testbus|blksync_testbus1|blksync_testbus2|gearbox_exp_testbus|random_ver_testbus|descramble_testbus|blank_testbus|rx_fifo_testbus1|rx_fifo_testbus2
		parameter hssi_10g_rx_pcs_rx_true_b2b = "b2b", // single|b2b
		parameter hssi_10g_rx_pcs_rxfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_rx_pcs_rxfifo_full = "full_default", // full_default
		parameter hssi_10g_rx_pcs_rxfifo_mode = "phase_comp", // register_mode|clk_comp_10g|generic_interlaken|generic_basic|phase_comp|phase_comp_dv
		parameter hssi_10g_rx_pcs_rxfifo_pempty = 5'b10,
		parameter hssi_10g_rx_pcs_rxfifo_pfull = 5'b10111,
		parameter hssi_10g_rx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_rx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_rx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_10g_tx_pcs
		parameter hssi_10g_tx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_bitslip_en = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_10g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_10g_tx_pcs_comp_cnt = 8'b0,
		parameter hssi_10g_tx_pcs_compin_sel = "compin_master", // compin_master|compin_slave_top|compin_slave_bot|compin_default
		parameter hssi_10g_tx_pcs_crcgen_bypass = "crcgen_bypass_dis", // crcgen_bypass_dis|crcgen_bypass_en
		parameter hssi_10g_tx_pcs_crcgen_clken = "crcgen_clk_dis", // crcgen_clk_dis|crcgen_clk_en
		parameter hssi_10g_tx_pcs_crcgen_err = "crcgen_err_dis", // crcgen_err_dis|crcgen_err_en
		parameter hssi_10g_tx_pcs_crcgen_inv = "crcgen_inv_dis", // crcgen_inv_dis|crcgen_inv_en
		parameter hssi_10g_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_tx_pcs_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_10g_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_tx_pcs_dft_clk_out_sel = "tx_master_clk", // tx_master_clk|tx_rdfifo_clk|tx_frmgen_clk|tx_crcgen_clk|tx_64b66benc_txsm_clk|tx_scrm_clk|tx_dispgen_clk|tx_gbred_clk|tx_wrfifo_clk|tx_fec_clk
		parameter hssi_10g_tx_pcs_dispgen_bypass = "dispgen_bypass_dis", // dispgen_bypass_dis|dispgen_bypass_en
		parameter hssi_10g_tx_pcs_dispgen_clken = "dispgen_clk_dis", // dispgen_clk_dis|dispgen_clk_en
		parameter hssi_10g_tx_pcs_dispgen_err = "dispgen_err_dis", // dispgen_err_dis|dispgen_err_en
		parameter hssi_10g_tx_pcs_dispgen_pipeln = "dispgen_pipeln_dis", // dispgen_pipeln_dis|dispgen_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_bypass_pipeln = "distdwn_bypass_pipeln_dis", // distdwn_bypass_pipeln_dis|distdwn_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_master = "distdwn_master_en", // distdwn_master_en|distdwn_master_dis
		parameter hssi_10g_tx_pcs_distup_bypass_pipeln = "distup_bypass_pipeln_dis", // distup_bypass_pipeln_dis|distup_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distup_master = "distup_master_en", // distup_master_en|distup_master_dis
		parameter hssi_10g_tx_pcs_dv_bond = "dv_bond_dis", // dv_bond_en|dv_bond_dis
		parameter hssi_10g_tx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_tx_pcs_enc64b66b_txsm_clken = "enc64b66b_txsm_clk_dis", // enc64b66b_txsm_clk_dis|enc64b66b_txsm_clk_en
		parameter hssi_10g_tx_pcs_enc_64b66b_txsm_bypass = "enc_64b66b_txsm_bypass_dis", // enc_64b66b_txsm_bypass_dis|enc_64b66b_txsm_bypass_en
		parameter hssi_10g_tx_pcs_fastpath = "fastpath_dis", // fastpath_dis|fastpath_en
		parameter hssi_10g_tx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_tx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_tx_pcs_fifo_double_write = "fifo_double_write_dis", // fifo_double_write_dis|fifo_double_write_en
		parameter hssi_10g_tx_pcs_fifo_reg_fast = "fifo_reg_fast_dis", // fifo_reg_fast_dis|fifo_reg_fast_en
		parameter hssi_10g_tx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_tx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_tx_pcs_frmgen_burst = "frmgen_burst_dis", // frmgen_burst_dis|frmgen_burst_en
		parameter hssi_10g_tx_pcs_frmgen_bypass = "frmgen_bypass_dis", // frmgen_bypass_dis|frmgen_bypass_en
		parameter hssi_10g_tx_pcs_frmgen_clken = "frmgen_clk_dis", // frmgen_clk_dis|frmgen_clk_en
		parameter hssi_10g_tx_pcs_frmgen_mfrm_length = 16'b100000000000,
		parameter hssi_10g_tx_pcs_frmgen_pipeln = "frmgen_pipeln_dis", // frmgen_pipeln_dis|frmgen_pipeln_en
		parameter hssi_10g_tx_pcs_frmgen_pyld_ins = "frmgen_pyld_ins_dis", // frmgen_pyld_ins_dis|frmgen_pyld_ins_en
		parameter hssi_10g_tx_pcs_frmgen_wordslip = "frmgen_wordslip_dis", // frmgen_wordslip_dis|frmgen_wordslip_en
		parameter hssi_10g_tx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_tx_pcs_gb_pipeln_bypass = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_gb_tx_idwidth = "width_50", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_tx_pcs_gb_tx_odwidth = "width_32", // width_32|width_40|width_64
		parameter hssi_10g_tx_pcs_gbred_clken = "gbred_clk_dis", // gbred_clk_dis|gbred_clk_en
		parameter hssi_10g_tx_pcs_indv = "indv_en", // indv_en|indv_dis
		parameter hssi_10g_tx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_tx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_tx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_tx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del6|phcomp_rd_del5|phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_tx_pcs_pld_if_type = "fifo", // fifo|reg|fastreg
		parameter hssi_10g_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_tx_pcs_pseudo_random = "all_0", // two_lf|all_0
		parameter hssi_10g_tx_pcs_pseudo_seed_a = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_pseudo_seed_b = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_random_disp = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_tx_pcs_scrm_bypass = "scrm_bypass_dis", // scrm_bypass_dis|scrm_bypass_en
		parameter hssi_10g_tx_pcs_scrm_clken = "scrm_clk_dis", // scrm_clk_dis|scrm_clk_en
		parameter hssi_10g_tx_pcs_scrm_mode = "async", // async|sync
		parameter hssi_10g_tx_pcs_scrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_sh_err = "sh_err_dis", // sh_err_dis|sh_err_en
		parameter hssi_10g_tx_pcs_sop_mark = "sop_mark_dis", // sop_mark_en|sop_mark_dis
		parameter hssi_10g_tx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_tx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_tx_pcs_tx_scrm_err = "scrm_err_dis", // scrm_err_dis|scrm_err_en
		parameter hssi_10g_tx_pcs_tx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_tx_pcs_tx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_tx_pcs_tx_sm_bypass = "tx_sm_bypass_dis", // tx_sm_bypass_dis|tx_sm_bypass_en
		parameter hssi_10g_tx_pcs_tx_sm_pipeln = "tx_sm_pipeln_dis", // tx_sm_pipeln_dis|tx_sm_pipeln_en
		parameter hssi_10g_tx_pcs_tx_testbus_sel = "crc32_gen_testbus1", // crc32_gen_testbus1|crc32_gen_testbus2|disp_gen_testbus1|disp_gen_testbus2|frame_gen_testbus1|frame_gen_testbus2|enc64b66b_testbus|txsm_testbus|tx_cp_bond_testbus|gearbox_red_testbus|scramble_testbus|blank_testbus|tx_fifo_testbus1|tx_fifo_testbus2
		parameter hssi_10g_tx_pcs_txfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_tx_pcs_txfifo_full = "full_default", // full_default
		parameter hssi_10g_tx_pcs_txfifo_mode = "phase_comp", // register_mode|interlaken_generic|basic_generic|phase_comp
		parameter hssi_10g_tx_pcs_txfifo_pempty = 4'b10,
		parameter hssi_10g_tx_pcs_txfifo_pfull = 4'b1011,
		parameter hssi_10g_tx_pcs_wr_clk_sel = "wr_tx_pma_clk", // wr_tx_pld_clk|wr_tx_pma_clk|wr_refclk_dig
		parameter hssi_10g_tx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_8g_rx_pcs
		parameter hssi_8g_rx_pcs_auto_error_replacement = "dis_err_replace", // dis_err_replace|en_err_replace
		parameter hssi_8g_rx_pcs_auto_speed_nego = "dis_asn", // dis_asn|en_asn_g2_freq_scal
		parameter hssi_8g_rx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_rx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_rx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_rx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_rx_pcs_byte_deserializer = "dis_bds", // dis_bds|en_bds_by_2|en_bds_by_4|en_bds_by_2_det
		parameter hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask = "dis_rxvalid_mask", // dis_rxvalid_mask|en_rxvalid_mask
		parameter hssi_8g_rx_pcs_clkcmp_pattern_n = 20'b0,
		parameter hssi_8g_rx_pcs_clkcmp_pattern_p = 20'b0,
		parameter hssi_8g_rx_pcs_clock_gate_bds_dec_asn = "dis_bds_dec_asn_clk_gating", // dis_bds_dec_asn_clk_gating|en_bds_dec_asn_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_cdr_eidle = "dis_cdr_eidle_clk_gating", // dis_cdr_eidle_clk_gating|en_cdr_eidle_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk = "dis_dw_pc_wrclk_gating", // dis_dw_pc_wrclk_gating|en_dw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_rd = "dis_dw_rm_rdclk_gating", // dis_dw_rm_rdclk_gating|en_dw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_wr = "dis_dw_rm_wrclk_gating", // dis_dw_rm_wrclk_gating|en_dw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_wa = "dis_dw_wa_clk_gating", // dis_dw_wa_clk_gating|en_dw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_pc_rdclk = "dis_pc_rdclk_gating", // dis_pc_rdclk_gating|en_pc_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk = "dis_sw_pc_wrclk_gating", // dis_sw_pc_wrclk_gating|en_sw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_rd = "dis_sw_rm_rdclk_gating", // dis_sw_rm_rdclk_gating|en_sw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_wr = "dis_sw_rm_wrclk_gating", // dis_sw_rm_wrclk_gating|en_sw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_wa = "dis_sw_wa_clk_gating", // dis_sw_wa_clk_gating|en_sw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_observation_in_pld_core = "internal_sw_wa_clk", // internal_sw_wa_clk|internal_dw_wa_clk|internal_cdr_eidle_clk|internal_sm_rm_wr_clk|internal_dw_rm_wr_clk|internal_clk_2_b|internal_sw_rm_rd_clk|internal_dw_rm_rd_clk|internal_sw_rx_wr_clk|internal_dw_rx_wr_clk|internal_rx_rd_clk|internal_rx_pma_clk_gen3|internal_rx_rcvd_clk_gen3
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_rx_pcs_eidle_entry_eios = "dis_eidle_eios", // dis_eidle_eios|en_eidle_eios
		parameter hssi_8g_rx_pcs_eidle_entry_iei = "dis_eidle_iei", // dis_eidle_iei|en_eidle_iei
		parameter hssi_8g_rx_pcs_eidle_entry_sd = "dis_eidle_sd", // dis_eidle_sd|en_eidle_sd
		parameter hssi_8g_rx_pcs_eightb_tenb_decoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_rx_pcs_err_flags_sel = "err_flags_wa", // err_flags_wa|err_flags_8b10b
		parameter hssi_8g_rx_pcs_fixed_pat_det = "dis_fixed_patdet", // dis_fixed_patdet|en_fixed_patdet
		parameter hssi_8g_rx_pcs_fixed_pat_num = 4'b1111,
		parameter hssi_8g_rx_pcs_force_signal_detect = "en_force_signal_detect", // en_force_signal_detect|dis_force_signal_detect
		parameter hssi_8g_rx_pcs_gen3_clk_en = "disable_clk", // disable_clk|enable_clk
		parameter hssi_8g_rx_pcs_gen3_rx_clk_sel = "rcvd_clk", // en_dig_clk1_8g|rcvd_clk
		parameter hssi_8g_rx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // en_dig_clk2_8g|tx_pma_clk
		parameter hssi_8g_rx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_rx_pcs_ibm_invalid_code = "dis_ibm_invalid_code", // dis_ibm_invalid_code|en_ibm_invalid_code
		parameter hssi_8g_rx_pcs_invalid_code_flag_only = "dis_invalid_code_only", // dis_invalid_code_only|en_invalid_code_only
		parameter hssi_8g_rx_pcs_pad_or_edb_error_replace = "replace_edb", // replace_edb|replace_edb_dynamic|replace_pad
		parameter hssi_8g_rx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_rx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_rx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_rx_pcs_pipe_if_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_8g_rx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_rx_pcs_polinv_8b10b_dec = "dis_polinv_8b10b_dec", // dis_polinv_8b10b_dec|en_polinv_8b10b_dec
		parameter hssi_8g_rx_pcs_prot_mode = "gige", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic_rm_enable|basic_rm_disable|disabled_prot_mode
		parameter hssi_8g_rx_pcs_rate_match = "dis_rm", // dis_rm|gige_rm|pipe_rm|pipe_rm_0ppm|sw_basic_rm|dw_basic_rm
		parameter hssi_8g_rx_pcs_rate_match_del_thres = "dis_rm_del_thres", // dis_rm_del_thres|gige_rm_del_thres|pipe_rm_del_thres|pipe_rm_0ppm_del_thres|sw_basic_rm_del_thres|dw_basic_rm_del_thres
		parameter hssi_8g_rx_pcs_rate_match_empty_thres = "dis_rm_empty_thres", // dis_rm_empty_thres|gige_rm_empty_thres|pipe_rm_empty_thres|pipe_rm_0ppm_empty_thres|sw_basic_rm_empty_thres|dw_basic_rm_empty_thres
		parameter hssi_8g_rx_pcs_rate_match_full_thres = "dis_rm_full_thres", // dis_rm_full_thres|gige_rm_full_thres|pipe_rm_full_thres|pipe_rm_0ppm_full_thres|sw_basic_rm_full_thres|dw_basic_rm_full_thres
		parameter hssi_8g_rx_pcs_rate_match_ins_thres = "dis_rm_ins_thres", // dis_rm_ins_thres|gige_rm_ins_thres|pipe_rm_ins_thres|pipe_rm_0ppm_ins_thres|sw_basic_rm_ins_thres|dw_basic_rm_ins_thres
		parameter hssi_8g_rx_pcs_rate_match_start_thres = "dis_rm_start_thres", // dis_rm_start_thres|gige_rm_start_thres|pipe_rm_start_thres|pipe_rm_0ppm_start_thres|sw_basic_rm_start_thres|dw_basic_rm_start_thres
		parameter hssi_8g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_rx_pcs_rx_clk2 = "rcvd_clk_clk2", // rcvd_clk_clk2|tx_pma_clock_clk2|refclk_dig2_clk2
		parameter hssi_8g_rx_pcs_rx_clk_free_running = "en_rx_clk_free_run", // dis_rx_clk_free_run|en_rx_clk_free_run
		parameter hssi_8g_rx_pcs_rx_pcs_urst = "en_rx_pcs_urst", // dis_rx_pcs_urst|en_rx_pcs_urst
		parameter hssi_8g_rx_pcs_rx_rcvd_clk = "rcvd_clk_rcvd_clk", // rcvd_clk_rcvd_clk|tx_pma_clock_rcvd_clk
		parameter hssi_8g_rx_pcs_rx_rd_clk = "pld_rx_clk", // pld_rx_clk|rx_clk
		parameter hssi_8g_rx_pcs_rx_refclk = "dis_refclk_sel", // dis_refclk_sel|en_refclk_sel
		parameter hssi_8g_rx_pcs_rx_wr_clk = "rx_clk2_div_1_2_4", // rx_clk2_div_1_2_4|txfifo_rd_clk
		parameter hssi_8g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_rx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_rx_pcs_sync_sm_idle_eios = "dis_syncsm_idle", // dis_syncsm_idle|en_syncsm_idle
		parameter hssi_8g_rx_pcs_test_bus_sel = "tx_testbus", // tx_testbus|tx_ctrl_plane_testbus|wa_testbus|rm_testbus|rx_ctrl_testbus|pcie_ctrl_testbus|rx_ctrl_plane_testbus
		parameter hssi_8g_rx_pcs_tx_rx_parallel_loopback = "dis_plpbk", // dis_plpbk|en_plpbk
		parameter hssi_8g_rx_pcs_wa_boundary_lock_ctrl = "bit_slip", // bit_slip|sync_sm|deterministic_latency|auto_align_pld_ctrl
		parameter hssi_8g_rx_pcs_wa_clk_slip_spacing = 10'b10000,
		parameter hssi_8g_rx_pcs_wa_det_latency_sync_status_beh = "assert_sync_status_non_imm", // assert_sync_status_imm|assert_sync_status_non_imm|dont_care_assert_sync
		parameter hssi_8g_rx_pcs_wa_disp_err_flag = "dis_disp_err_flag", // dis_disp_err_flag|en_disp_err_flag
		parameter hssi_8g_rx_pcs_wa_kchar = "dis_kchar", // dis_kchar|en_kchar
		parameter hssi_8g_rx_pcs_wa_pd = "wa_pd_10", // wa_pd_7|wa_pd_10|wa_pd_20|wa_pd_40|wa_pd_8_sw|wa_pd_8_dw|wa_pd_16_sw|wa_pd_16_dw|wa_pd_32
		parameter hssi_8g_rx_pcs_wa_pd_data = 40'b0,
		parameter hssi_8g_rx_pcs_wa_pd_polarity = "dis_pd_both_pol", // dis_pd_both_pol|en_pd_both_pol|dont_care_both_pol
		parameter hssi_8g_rx_pcs_wa_pld_controlled = "dis_pld_ctrl", // dis_pld_ctrl|pld_ctrl_sw|rising_edge_sensitive_dw|level_sensitive_dw
		parameter hssi_8g_rx_pcs_wa_renumber_data = 6'b0,
		parameter hssi_8g_rx_pcs_wa_rgnumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rknumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rosnumber_data = 2'b0,
		parameter hssi_8g_rx_pcs_wa_rvnumber_data = 13'b0,
		parameter hssi_8g_rx_pcs_wa_sync_sm_ctrl = "gige_sync_sm", // gige_sync_sm|pipe_sync_sm|sw_basic_sync_sm|dw_basic_sync_sm|fibre_channel_sync_sm
		parameter hssi_8g_rx_pcs_wait_cnt = 12'b0,
		
		// parameters for twentynm_hssi_8g_tx_pcs
		parameter hssi_8g_tx_pcs_auto_speed_nego_gen2 = "dis_asn_g2", // dis_asn_g2|en_asn_g2_freq_scal
		parameter hssi_8g_tx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_tx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_tx_pcs_byte_serializer = "dis_bs", // dis_bs|en_bs_by_2|en_bs_by_4
		parameter hssi_8g_tx_pcs_clock_gate_bs_enc = "dis_bs_enc_clk_gating", // dis_bs_enc_clk_gating|en_bs_enc_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_dw_fifowr = "dis_dw_fifowr_clk_gating", // dis_dw_fifowr_clk_gating|en_dw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_fiford = "dis_fiford_clk_gating", // dis_fiford_clk_gating|en_fiford_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_sw_fifowr = "dis_sw_fifowr_clk_gating", // dis_sw_fifowr_clk_gating|en_sw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_observation_in_pld_core = "internal_refclk_b", // internal_refclk_b|internal_fifo_rd_clk|internal_sw_fifo_wr_clk|internal_dw_fifo_wr_clk|internal_tx_clk_out_gen3|internal_pipe_tx_clk_out_gen3
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_tx_pcs_data_selection_8b10b_encoder_input = "normal_data_path", // normal_data_path|gige_idle_conversion
		parameter hssi_8g_tx_pcs_dynamic_clk_switch = "dis_dyn_clk_switch", // dis_dyn_clk_switch|en_dyn_clk_switch
		parameter hssi_8g_tx_pcs_eightb_tenb_disp_ctrl = "dis_disp_ctrl", // dis_disp_ctrl|en_disp_ctrl|en_ib_disp_ctrl
		parameter hssi_8g_tx_pcs_eightb_tenb_encoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_tx_pcs_force_echar = "dis_force_echar", // dis_force_echar|en_force_echar
		parameter hssi_8g_tx_pcs_force_kchar = "dis_force_kchar", // dis_force_kchar|en_force_kchar
		parameter hssi_8g_tx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // dis_tx_clk|tx_pma_clk
		parameter hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel = "func_clk", // dis_tx_pipe_clk|func_clk
		parameter hssi_8g_tx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_tx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_tx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_tx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_tx_pcs_phfifo_write_clk_sel = "pld_tx_clk", // pld_tx_clk|tx_clk
		parameter hssi_8g_tx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_tx_pcs_prot_mode = "basic", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic|disabled_prot_mode
		parameter hssi_8g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_tx_pcs_refclk_b_clk_sel = "tx_pma_clock", // tx_pma_clock|refclk_dig
		parameter hssi_8g_tx_pcs_revloop_back_rm = "dis_rev_loopback_rx_rm", // dis_rev_loopback_rx_rm|en_rev_loopback_rx_rm
		parameter hssi_8g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_tx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_tx_pcs_tx_bitslip = "dis_tx_bitslip", // dis_tx_bitslip|en_tx_bitslip
		parameter hssi_8g_tx_pcs_tx_compliance_controlled_disparity = "dis_txcompliance", // dis_txcompliance|en_txcompliance_pipe2p0|en_txcompliance_pipe3p0
		parameter hssi_8g_tx_pcs_tx_fast_pld_reg = "dis_tx_fast_pld_reg", // dis_tx_fast_pld_reg|en_tx_fast_pld_reg
		parameter hssi_8g_tx_pcs_txclk_freerun = "dis_freerun_tx", // dis_freerun_tx|en_freerun_tx
		parameter hssi_8g_tx_pcs_txpcs_urst = "en_txpcs_urst", // dis_txpcs_urst|en_txpcs_urst
		
		// parameters for twentynm_hssi_common_pcs_pma_interface
		parameter hssi_common_pcs_pma_interface_asn_clk_enable = "false", // false|true
		parameter hssi_common_pcs_pma_interface_asn_enable = "dis_asn", // dis_asn|en_asn
		parameter hssi_common_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|pcie_gen3
		parameter hssi_common_pcs_pma_interface_bypass_early_eios = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pcie_switch = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_ltr = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_sw_done = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_ppm_lock = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_txdetectrx = "false", // false|true
		parameter hssi_common_pcs_pma_interface_cdr_control = "en_cdr_ctrl", // dis_cdr_ctrl|en_cdr_ctrl
		parameter hssi_common_pcs_pma_interface_cid_enable = "en_cid_mode", // dis_cid_mode|en_cid_mode
		parameter hssi_common_pcs_pma_interface_cp_cons_sel = "cp_cons_default", // cp_cons_master|cp_cons_slave_abv|cp_cons_slave_blw|cp_cons_default
		parameter hssi_common_pcs_pma_interface_cp_dwn_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_cp_up_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_blw|ctrl_slave_abv
		parameter hssi_common_pcs_pma_interface_data_mask_count = 16'b100111000100,
		parameter hssi_common_pcs_pma_interface_data_mask_count_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_dft_observation_clock_selection = "dft_clk_obsrv_tx0", // dft_clk_obsrv_tx0|dft_clk_obsrv_tx1|dft_clk_obsrv_tx2|dft_clk_obsrv_tx3|dft_clk_obsrv_tx4|dft_clk_obsrv_rx|dft_clk_obsrv_hclk|dft_clk_obsrv_fref|dft_clk_obsrv_clklow|dft_clk_obsrv_asn0|dft_clk_obsrv_asn1
		parameter hssi_common_pcs_pma_interface_early_eios_counter = 8'b110010,
		parameter hssi_common_pcs_pma_interface_force_freqdet = "force_freqdet_dis", // force_freqdet_dis|force1_freqdet_en|force0_freqdet_en
		parameter hssi_common_pcs_pma_interface_free_run_clk_enable = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ignore_sigdet_g23 = "false", // false|true
		parameter hssi_common_pcs_pma_interface_pc_en_counter = 7'b110111,
		parameter hssi_common_pcs_pma_interface_pc_rst_counter = 5'b10111,
		parameter hssi_common_pcs_pma_interface_pcie_hip_mode = "hip_disable", // hip_enable|hip_disable
		parameter hssi_common_pcs_pma_interface_ph_fifo_reg_mode = "phfifo_reg_mode_dis", // phfifo_reg_mode_dis|phfifo_reg_mode_en
		parameter hssi_common_pcs_pma_interface_phfifo_flush_wait = 6'b100100,
		parameter hssi_common_pcs_pma_interface_pipe_if_g3pcs = "pipe_if_8gpcs", // pipe_if_g3pcs|pipe_if_8gpcs
		parameter hssi_common_pcs_pma_interface_pma_done_counter = 18'b101010101110011000,
		parameter hssi_common_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_common_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_common_pcs_pma_interface_ppm_cnt_rst = "ppm_cnt_rst_dis", // ppm_cnt_rst_dis|ppm_cnt_rst_en
		parameter hssi_common_pcs_pma_interface_ppm_deassert_early = "deassert_early_dis", // deassert_early_dis|deassert_early_en
		parameter hssi_common_pcs_pma_interface_ppm_det_buckets = "ppm_100_bucket", // disable_prot|ppm_300_bucket|ppm_100_bucket|ppm_300_100_bucket
		parameter hssi_common_pcs_pma_interface_ppm_gen1_2_cnt = "cnt_32k", // cnt_32k|cnt_64k
		parameter hssi_common_pcs_pma_interface_ppm_post_eidle_delay = "cnt_200_cycles", // cnt_200_cycles|cnt_400_cycles
		parameter hssi_common_pcs_pma_interface_ppmsel = "ppmsel_300", // ppmsel_disable|ppmsel_5000|ppmsel_2500|ppmsel_1000|ppmsel_500|ppmsel_300|ppmsel_250|ppmsel_200|ppmsel_125|ppmsel_100|ppmsel_62p5|ppm_other
		parameter hssi_common_pcs_pma_interface_prot_mode = "disable_prot_mode", // disable_prot_mode|pipe_g12|pipe_g3|other_protocols
		parameter hssi_common_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_common_pcs_pma_interface_rxvalid_mask = "rxvalid_mask_en", // rxvalid_mask_dis|rxvalid_mask_en
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter = 12'b100111000100,
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_sim_mode = "disable", // disable|enable
		parameter hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en = "true", // false|true
		parameter hssi_common_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_common_pcs_pma_interface_testout_sel = "ppm_det_test", // ppm_det_test|asn_test|pma_pll_test|rxpmaif_test|prbs_gen_test|prbs_ver_test|uhsif_1_test|uhsif_2_test|uhsif_3_test
		parameter hssi_common_pcs_pma_interface_wait_clk_on_off_timer = 4'b100,
		parameter hssi_common_pcs_pma_interface_wait_pipe_synchronizing = 5'b10111,
		parameter hssi_common_pcs_pma_interface_wait_send_syncp_fbkp = 11'b11111010,
		
		// parameters for twentynm_hssi_common_pld_pcs_interface
		parameter hssi_common_pld_pcs_interface_dft_clk_out_en = "dft_clk_out_disable", // dft_clk_out_disable|dft_clk_out_enable
		parameter hssi_common_pld_pcs_interface_dft_clk_out_sel = "teng_rx_dft_clk", // teng_rx_dft_clk|teng_tx_dft_clk|eightg_rx_dft_clk|eightg_tx_dft_clk|pmaif_dft_clk
		parameter hssi_common_pld_pcs_interface_hrdrstctrl_en = "hrst_dis", // hrst_dis|hrst_en
		parameter hssi_common_pld_pcs_interface_pcs_testbus_block_sel = "eightg", // eightg|g3pcs|teng|krfec|pma_if
		parameter hssi_common_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_fifo_rx_pcs
		parameter hssi_fifo_rx_pcs_double_read_mode = "double_read_dis", // double_read_en|double_read_dis
		parameter hssi_fifo_rx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_fifo_tx_pcs
		parameter hssi_fifo_tx_pcs_double_write_mode = "double_write_dis", // double_write_en|double_write_dis
		parameter hssi_fifo_tx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_gen3_rx_pcs
		parameter hssi_gen3_rx_pcs_block_sync = "enable_block_sync", // bypass_block_sync|enable_block_sync
		parameter hssi_gen3_rx_pcs_block_sync_sm = "enable_blk_sync_sm", // disable_blk_sync_sm|enable_blk_sync_sm
		parameter hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn = "enable", // disable|enable
		parameter hssi_gen3_rx_pcs_lpbk_force = "lpbk_frce_dis", // lpbk_frce_dis|lpbk_frce_en
		parameter hssi_gen3_rx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_rx_pcs_rate_match_fifo = "enable_rm_fifo_600ppm", // bypass_rm_fifo|enable_rm_fifo_600ppm|enable_rm_fifo_0ppm
		parameter hssi_gen3_rx_pcs_rate_match_fifo_latency = "regular_latency", // regular_latency|low_latency
		parameter hssi_gen3_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_gen3_rx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_b4gb_par_lpbk = "b4gb_par_lpbk_dis", // b4gb_par_lpbk_dis|b4gb_par_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_force_balign = "en_force_balign", // en_force_balign|dis_force_balign
		parameter hssi_gen3_rx_pcs_rx_ins_del_one_skip = "ins_del_one_skip_en", // ins_del_one_skip_dis|ins_del_one_skip_en
		parameter hssi_gen3_rx_pcs_rx_num_fixed_pat = 4'b1000,
		parameter hssi_gen3_rx_pcs_rx_test_out_sel = "rx_test_out0", // rx_test_out0|rx_test_out1
		parameter hssi_gen3_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_gen3_tx_pcs
		parameter hssi_gen3_tx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_tx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_gen3_tx_pcs_tx_bitslip = 5'b0,
		parameter hssi_gen3_tx_pcs_tx_gbox_byp = "bypass_gbox", // bypass_gbox|enable_gbox
		
		// parameters for twentynm_hssi_krfec_rx_pcs
		parameter hssi_krfec_rx_pcs_blksync_cor_en = "detect", // detect|correct
		parameter hssi_krfec_rx_pcs_bypass_gb = "bypass_dis", // bypass_dis|bypass_en
		parameter hssi_krfec_rx_pcs_clr_ctrl = "both_enabled", // both_enabled|corr_cnt_only|uncorr_cnt_only
		parameter hssi_krfec_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_rx_pcs_dv_start = "with_blklock", // with_blksync|with_blklock
		parameter hssi_krfec_rx_pcs_err_mark_type = "err_mark_10g", // err_mark_10g|err_mark_40g
		parameter hssi_krfec_rx_pcs_error_marking_en = "err_mark_dis", // err_mark_dis|err_mark_en
		parameter hssi_krfec_rx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_krfec_rx_pcs_parity_invalid_enum = 8'b1000,
		parameter hssi_krfec_rx_pcs_parity_valid_num = 4'b100,
		parameter hssi_krfec_rx_pcs_pipeln_blksync = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_descrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errcorrect = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_ind = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_lfsr = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_loc = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_pat = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_gearbox = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_syndrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_trans_dec = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_rx_pcs_receive_order = "receive_lsb", // receive_lsb|receive_msb
		parameter hssi_krfec_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_krfec_rx_pcs_rx_testbus_sel = "overall", // overall|fast_search|fast_search_cntrs|blksync|blksync_cntrs|decoder_master_sm|decoder_master_sm_cntrs|syndrm_sm|syndrm1|syndrm2|errtrap_sm|errtrap_ind1|errtrap_ind2|errtrap_ind3|errtrap_ind4|errtrap_ind5|errtrap_loc|errtrap_pat1|errtrap_pat2|errtrap_pat3|errtrap_pat4|decoder_rd_sm|gb_and_trans
		parameter hssi_krfec_rx_pcs_signal_ok_en = "sig_ok_dis", // sig_ok_dis|sig_ok_en
		parameter hssi_krfec_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_krfec_tx_pcs
		parameter hssi_krfec_tx_pcs_burst_err = "burst_err_dis", // burst_err_dis|burst_err_en
		parameter hssi_krfec_tx_pcs_burst_err_len = "burst_err_len1", // burst_err_len1|burst_err_len2|burst_err_len3|burst_err_len4|burst_err_len5|burst_err_len6|burst_err_len7|burst_err_len8|burst_err_len9|burst_err_len10|burst_err_len11|burst_err_len12|burst_err_len13|burst_err_len14|burst_err_len15|burst_err_len16
		parameter hssi_krfec_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_tx_pcs_enc_frame_query = "enc_query_dis", // enc_query_dis|enc_query_en
		parameter hssi_krfec_tx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_encoder = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_scrambler = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_krfec_tx_pcs_transcode_err = "trans_err_dis", // trans_err_dis|trans_err_en
		parameter hssi_krfec_tx_pcs_transmit_order = "transmit_lsb", // transmit_lsb|transmit_msb
		parameter hssi_krfec_tx_pcs_tx_testbus_sel = "overall", // overall|encoder1|encoder2|scramble1|scramble2|scramble3|gearbox
		
		// parameters for twentynm_hssi_pipe_gen1_2
		parameter hssi_pipe_gen1_2_elec_idle_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_error_replace_pad = "replace_edb", // replace_edb|replace_pad
		parameter hssi_pipe_gen1_2_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_pipe_gen1_2_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen1_2_phystatus_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_phystatus_rst_toggle = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen1_2_pipe_byte_de_serializer_en = "dont_care_bds", // dis_bds|en_bds_by_2|dont_care_bds
		parameter hssi_pipe_gen1_2_prot_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|basic|disabled_prot_mode
		parameter hssi_pipe_gen1_2_reconfig_settings = "{}", // 
		parameter hssi_pipe_gen1_2_rx_pipe_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_pipe_gen1_2_rxdetect_bypass = "dis_rxdetect_bypass", // dis_rxdetect_bypass|en_rxdetect_bypass
		parameter hssi_pipe_gen1_2_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen1_2_tx_pipe_enable = "dis_pipe_tx", // dis_pipe_tx|en_pipe_tx|en_pipe3_tx
		parameter hssi_pipe_gen1_2_txswing = "dis_txswing", // dis_txswing|en_txswing
		
		// parameters for twentynm_hssi_pipe_gen3
		parameter hssi_pipe_gen3_bypass_rx_detection_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_rx_preset = 3'b0,
		parameter hssi_pipe_gen3_bypass_rx_preset_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_tx_coefficent = 18'b0,
		parameter hssi_pipe_gen3_bypass_tx_coefficent_enable = "false", // false|true
		parameter hssi_pipe_gen3_elecidle_delay_g3 = 3'b110,
		parameter hssi_pipe_gen3_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen3_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|disable_pcs
		parameter hssi_pipe_gen3_phy_status_delay_g12 = 3'b101,
		parameter hssi_pipe_gen3_phy_status_delay_g3 = 3'b101,
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g12 = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g3 = "dis_phystatus_rst_toggle_g3", // dis_phystatus_rst_toggle_g3|en_phystatus_rst_toggle_g3
		parameter hssi_pipe_gen3_rate_match_pad_insertion = "dis_rm_fifo_pad_ins", // dis_rm_fifo_pad_ins|en_rm_fifo_pad_ins
		parameter hssi_pipe_gen3_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen3_test_out_sel = "disable_test_out", // tx_test_out|rx_test_out|pipe_test_out1|pipe_test_out2|pipe_test_out3|pipe_ctrl_test_out|disable_test_out
		
		// parameters for twentynm_hssi_rx_pcs_pma_interface
		parameter hssi_rx_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|ten_g_pcs|direct_pld
		parameter hssi_rx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pcs_pma_interface_clkslip_sel = "pld", // pld|slip_eight_g_pcs
		parameter hssi_rx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pcs_pma_interface_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_rx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_rx_pcs_pma_interface_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_rx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_rx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_rx_pcs_pma_interface_prbs_ver = "prbs_off", // prbs_off|prbs_31|prbs_15|prbs_23|prbs_9|prbs_7
		parameter hssi_rx_pcs_pma_interface_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion = "rx_dyn_polinv_dis", // rx_dyn_polinv_dis|rx_dyn_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_lpbk_en = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok = "unforce_sig_ok", // unforce_sig_ok|force_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mask = "prbsmask128", // prbsmask128|prbsmask256|prbsmask512|prbsmask1024
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mode = "teng_mode", // teng_mode|eightg_mode
		parameter hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel = "sel_sig_det", // sel_sig_det|sel_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_static_polarity_inversion = "rx_stat_polinv_dis", // rx_stat_polinv_dis|rx_stat_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en = "uhsif_lpbk_dis", // uhsif_lpbk_dis|uhsif_lpbk_en
		parameter hssi_rx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_rx_pld_pcs_interface
		parameter hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx = "enable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx = "pma_64b_rx", // pma_32b_rx|pma_40b_rx|pma_64b_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_baser_mode_rx|interlaken_mode_rx|sfis_mode_rx|teng_sdi_mode_rx|basic_mode_rx|test_prp_mode_rx|test_prp_krfec_mode_rx|teng_1588_mode_rx|teng_baser_krfec_mode_rx|teng_1588_krfec_mode_rx|basic_krfec_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx = "disabled_prot_mode_rx", // pipe_g1_rx|pipe_g2_rx|pipe_g3_rx|cpri_rx|cpri_rx_tx_rx|gige_rx|gige_1588_rx|basic_rm_enable_rx|basic_rm_disable_rx|disabled_prot_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcie_g1_capable_rx|pcie_g2_capable_rx|pcie_g3_capable_rx|gige_rx|teng_baser_rx|teng_basekr_krfec_rx|fortyg_basekr_krfec_rx|cpri_8b10b_rx|interlaken_rx|sfis_rx|teng_sdi_rx|gige_1588_rx|teng_1588_baser_rx|teng_1588_basekr_krfec_rx|basic_8gpcs_rm_enable_rx|basic_8gpcs_rm_disable_rx|basic_10gpcs_rx|basic_10gpcs_krfec_rx|pcs_direct_rx|prp_rx|prp_krfec_rx|prbs_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx = "teng_mode_rx", // teng_mode_rx|non_teng_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_basekr_mode_rx|fortyg_basekr_mode_rx|teng_1588_basekr_mode_rx|basic_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|eightg_and_g3_pld_fifo_mode_rx|eightg_and_g3_reg_mode_rx|eightg_and_g3_reg_mode_hip_rx|teng_pld_fifo_mode_rx|teng_reg_mode_rx|teng_and_krfec_pld_fifo_mode_rx|teng_and_krfec_reg_mode_rx|pcs_direct_reg_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_block_sel = "pcs_direct", // eightg|teng|pcs_direct
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_rx_clk|pma_rx_clk_user
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_sel = "pld_rx_clk", // pld_rx_clk|pcs_rx_clk
		parameter hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en = "hip_rx_enable", // hip_rx_enable|hip_rx_disable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_rx_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_tx_pcs_pma_interface
		parameter hssi_tx_pcs_pma_interface_bypass_pma_txelecidle = "false", // false|true
		parameter hssi_tx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pcs_pma_interface_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx = "other_prot_mode", // pipe_g12|pipe_g3|other_prot_mode
		parameter hssi_tx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_tx_pcs_pma_interface_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_tx_pcs_pma_interface_pmagate_en = "pmagate_dis", // pmagate_dis|pmagate_en
		parameter hssi_tx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_tx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_tx_pcs_pma_interface_prbs_gen_pat = "prbs_gen_dis", // prbs_gen_dis|prbs_31|prbs_23|prbs_15|prbs_9|prbs_7
		parameter hssi_tx_pcs_pma_interface_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_tx_pcs_pma_interface_sq_wave_num = "sq_wave_4", // sq_wave_1|sq_wave_4|sq_wave_8|sq_wave_6|sq_wave_default
		parameter hssi_tx_pcs_pma_interface_sqwgen_clken = "sqwgen_clk_dis", // sqwgen_clk_dis|sqwgen_clk_en
		parameter hssi_tx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion = "tx_dyn_polinv_dis", // tx_dyn_polinv_dis|tx_dyn_polinv_en
		parameter hssi_tx_pcs_pma_interface_tx_pma_data_sel = "pld_dir", // pld_dir|pcie_gen3|eight_g_pcs|ten_g_pcs|prbs_pat|sq_wave_pat|block_sel_default|registered_uhsif_dat|directed_uhsif_dat
		parameter hssi_tx_pcs_pma_interface_tx_static_polarity_inversion = "tx_stat_polinv_dis", // tx_stat_polinv_dis|tx_stat_polinv_en
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock = "uhsif_filt_stepsz_b4lock_4", // uhsif_filt_stepsz_b4lock_2|uhsif_filt_stepsz_b4lock_4|uhsif_filt_stepsz_b4lock_6|uhsif_filt_stepsz_b4lock_8
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value = 4'b1011,
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock = "uhsif_filt_cntthr_b4lock_16", // uhsif_filt_cntthr_b4lock_8|uhsif_filt_cntthr_b4lock_16|uhsif_filt_cntthr_b4lock_24|uhsif_filt_cntthr_b4lock_32
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period = "uhsif_dcn_test_period_4", // uhsif_dcn_test_period_4|uhsif_dcn_test_period_8|uhsif_dcn_test_period_12|uhsif_dcn_test_period_16
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable = "uhsif_dcn_test_mode_disable", // uhsif_dcn_test_mode_enable|uhsif_dcn_test_mode_disable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh = "uhsif_dzt_cnt_thr_4", // uhsif_dzt_cnt_thr_2|uhsif_dzt_cnt_thr_4|uhsif_dzt_cnt_thr_6|uhsif_dzt_cnt_thr_8
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable = "uhsif_dzt_enable", // uhsif_dzt_disable|uhsif_dzt_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window = "uhsif_dzt_obr_win_32", // uhsif_dzt_obr_win_16|uhsif_dzt_obr_win_32|uhsif_dzt_obr_win_48|uhsif_dzt_obr_win_64
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size = "uhsif_dzt_skipsz_8", // uhsif_dzt_skipsz_4|uhsif_dzt_skipsz_8|uhsif_dzt_skipsz_12|uhsif_dzt_skipsz_16
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel = "uhsif_index_internal", // uhsif_index_internal|uhsif_index_cram
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin = "uhsif_dcn_margin_4", // uhsif_dcn_margin_2|uhsif_dcn_margin_3|uhsif_dcn_margin_4|uhsif_dcn_margin_5
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value = 8'b10000000,
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control = "uhsif_dft_dz_det_val_0", // uhsif_dft_dz_det_val_0|uhsif_dft_dz_det_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control = "uhsif_dft_up_val_0", // uhsif_dft_up_val_0|uhsif_dft_up_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_enable = "uhsif_disable", // uhsif_disable|uhsif_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock = "uhsif_lkd_segsz_aflock_2048", // uhsif_lkd_segsz_aflock_512|uhsif_lkd_segsz_aflock_1024|uhsif_lkd_segsz_aflock_2048|uhsif_lkd_segsz_aflock_4096
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock = "uhsif_lkd_segsz_b4lock_32", // uhsif_lkd_segsz_b4lock_16|uhsif_lkd_segsz_b4lock_32|uhsif_lkd_segsz_b4lock_64|uhsif_lkd_segsz_b4lock_128
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value = 4'b11,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value = 4'b11,
		
		// parameters for twentynm_hssi_tx_pld_pcs_interface
		parameter hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx = "enable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx = "pma_64b_tx", // pma_32b_tx|pma_40b_tx|pma_64b_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_baser_mode_tx|interlaken_mode_tx|sfis_mode_tx|teng_sdi_mode_tx|basic_mode_tx|test_prp_mode_tx|test_prp_krfec_mode_tx|teng_1588_mode_tx|teng_baser_krfec_mode_tx|teng_1588_krfec_mode_tx|basic_krfec_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx = "disabled_prot_mode_tx", // pipe_g1_tx|pipe_g2_tx|pipe_g3_tx|cpri_tx|cpri_rx_tx_tx|gige_tx|gige_1588_tx|basic_tx|disabled_prot_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcie_g1_capable_tx|pcie_g2_capable_tx|pcie_g3_capable_tx|gige_tx|teng_baser_tx|teng_basekr_krfec_tx|fortyg_basekr_krfec_tx|cpri_8b10b_tx|interlaken_tx|sfis_tx|teng_sdi_tx|gige_1588_tx|teng_1588_baser_tx|teng_1588_basekr_krfec_tx|basic_8gpcs_tx|basic_10gpcs_tx|basic_10gpcs_krfec_tx|pcs_direct_tx|uhsif_tx|prp_tx|prp_krfec_tx|prbs_tx|sqwave_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx = "teng_mode_tx", // teng_mode_tx|non_teng_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_basekr_mode_tx|fortyg_basekr_mode_tx|teng_1588_basekr_mode_tx|basic_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|eightg_and_g3_pld_fifo_mode_tx|eightg_and_g3_reg_mode_tx|eightg_and_g3_reg_mode_hip_tx|eightg_and_g3_fastreg_mode_tx|teng_pld_fifo_mode_tx|teng_reg_mode_tx|teng_fastreg_mode_tx|teng_and_krfec_pld_fifo_mode_tx|teng_and_krfec_reg_mode_tx|teng_and_krfec_fastreg_mode_tx|pcs_direct_fastreg_mode_tx|uhsif_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_tx_clk|pma_tx_clk_user
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_source = "teng", // eightg|teng|pma_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_data_source = "hip_disable", // hip_disable|hip_enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en = "delay1_clk_disable", // delay1_clk_enable|delay1_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel = "pld_tx_clk", // pld_tx_clk|pcs_tx_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl = "delay1_path0", // delay1_path0|delay1_path1|delay1_path2|delay1_path3|delay1_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel = "one_ff_delay", // one_ff_delay|two_ff_delay
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en = "delay2_clk_disable", // delay2_clk_enable|delay2_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl = "delay2_path0", // delay2_path0|delay2_path1|delay2_path2|delay2_path3|delay2_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_tx_pld_pcs_interface_reconfig_settings = "{}" // 
	//PARAM_LIST_END
	)
	(
	//PORT_LIST_START
		input wire	[8:0]	in_avmmaddress,
		input wire		in_avmmclk,
		input wire		in_avmmread,
		input wire		in_avmmrstn,
		input wire		in_avmmwrite,
		input wire	[7:0]	in_avmmwritedata,
		input wire	[4:0]	in_bond_pcs10g_in_bot,
		input wire	[4:0]	in_bond_pcs10g_in_top,
		input wire	[12:0]	in_bond_pcs8g_in_bot,
		input wire	[12:0]	in_bond_pcs8g_in_top,
		input wire	[11:0]	in_bond_pmaif_in_bot,
		input wire	[11:0]	in_bond_pmaif_in_top,
		input wire	[63:0]	in_hip_tx_data,
		input wire		in_iocsr_clk,
		input wire	[5:0]	in_iocsr_config,
		input wire		in_iocsr_rdy,
		input wire		in_iocsr_rdy_dly,
		input wire		in_pld_10g_krfec_rx_clr_errblk_cnt,
		input wire		in_pld_10g_krfec_rx_pld_rst_n,
		input wire		in_pld_10g_krfec_tx_pld_rst_n,
		input wire		in_pld_10g_rx_align_clr,
		input wire		in_pld_10g_rx_clr_ber_count,
		input wire		in_pld_10g_rx_rd_en,
		input wire	[6:0]	in_pld_10g_tx_bitslip,
		input wire		in_pld_10g_tx_burst_en,
		input wire		in_pld_10g_tx_data_valid,
		input wire	[1:0]	in_pld_10g_tx_diag_status,
		input wire		in_pld_10g_tx_wordslip,
		input wire		in_pld_8g_a1a2_size,
		input wire		in_pld_8g_bitloc_rev_en,
		input wire		in_pld_8g_byte_rev_en,
		input wire	[2:0]	in_pld_8g_eidleinfersel,
		input wire		in_pld_8g_encdt,
		input wire		in_pld_8g_g3_rx_pld_rst_n,
		input wire		in_pld_8g_g3_tx_pld_rst_n,
		input wire		in_pld_8g_rddisable_tx,
		input wire		in_pld_8g_rdenable_rx,
		input wire		in_pld_8g_refclk_dig2,
		input wire		in_pld_8g_rxpolarity,
		input wire	[4:0]	in_pld_8g_tx_boundary_sel,
		input wire		in_pld_8g_wrdisable_rx,
		input wire		in_pld_8g_wrenable_tx,
		input wire		in_pld_atpg_los_en_n,
		input wire		in_pld_bitslip,
		input wire	[17:0]	in_pld_g3_current_coeff,
		input wire	[2:0]	in_pld_g3_current_rxpreset,
		input wire		in_pld_ltr,
		input wire		in_pld_mem_krfec_atpg_rst_n,
		input wire		in_pld_partial_reconfig,
		input wire		in_pld_pcs_refclk_dig,
		input wire		in_pld_pma_adapt_start,
		input wire		in_pld_pma_csr_test_dis,
		input wire		in_pld_pma_early_eios,
		input wire	[5:0]	in_pld_pma_eye_monitor,
		input wire		in_pld_pma_ltd_b,
		input wire		in_pld_pma_nrpi_freeze,
		input wire	[1:0]	in_pld_pma_pcie_switch,
		input wire		in_pld_pma_ppm_lock,
		input wire	[4:0]	in_pld_pma_reserved_out,
		input wire		in_pld_pma_rs_lpbk_b,
		input wire		in_pld_pma_rx_qpi_pullup,
		input wire		in_pld_pma_rxpma_rstb,
		input wire		in_pld_pma_tx_bitslip,
		input wire		in_pld_pma_tx_bonding_rstb,
		input wire		in_pld_pma_tx_qpi_pulldn,
		input wire		in_pld_pma_tx_qpi_pullup,
		input wire		in_pld_pma_txdetectrx,
		input wire		in_pld_pma_txpma_rstb,
		input wire		in_pld_pmaif_rx_pld_rst_n,
		input wire		in_pld_pmaif_rxclkslip,
		input wire		in_pld_pmaif_tx_pld_rst_n,
		input wire		in_pld_polinv_rx,
		input wire		in_pld_polinv_tx,
		input wire	[1:0]	in_pld_rate,
		input wire	[9:0]	in_pld_reserved_in,
		input wire		in_pld_rx_clk,
		input wire		in_pld_rx_prbs_err_clr,
		input wire		in_pld_scan_mode_n,
		input wire		in_pld_scan_shift_n,
		input wire		in_pld_syncsm_en,
		input wire		in_pld_tx_clk,
		input wire	[17:0]	in_pld_tx_control,
		input wire	[127:0]	in_pld_tx_data,
		input wire		in_pld_txelecidle,
		input wire		in_pld_uhsif_tx_clk,
		input wire		in_pma_adapt_done,
		input wire		in_pma_clklow,
		input wire		in_pma_fref,
		input wire		in_pma_hclk,
		input wire	[1:0]	in_pma_pcie_sw_done,
		input wire		in_pma_pfdmode_lock,
		input wire	[4:0]	in_pma_reserved_in,
		input wire		in_pma_rx_clkdiv_user,
		input wire		in_pma_rx_detect_valid,
		input wire		in_pma_rx_found,
		input wire		in_pma_rx_pma_clk,
		input wire	[63:0]	in_pma_rx_pma_data,
		input wire		in_pma_rx_signal_ok,
		input wire		in_pma_rxpll_lock,
		input wire		in_pma_signal_det,
		input wire	[7:0]	in_pma_testbus,
		input wire		in_pma_tx_clkdiv_user,
		input wire		in_pma_tx_pma_clk,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen1_2,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen3,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pld_pcs_interface,
		output wire		out_blockselect_hssi_10g_rx_pcs,
		output wire		out_blockselect_hssi_10g_tx_pcs,
		output wire		out_blockselect_hssi_8g_rx_pcs,
		output wire		out_blockselect_hssi_8g_tx_pcs,
		output wire		out_blockselect_hssi_common_pcs_pma_interface,
		output wire		out_blockselect_hssi_common_pld_pcs_interface,
		output wire		out_blockselect_hssi_fifo_rx_pcs,
		output wire		out_blockselect_hssi_fifo_tx_pcs,
		output wire		out_blockselect_hssi_gen3_rx_pcs,
		output wire		out_blockselect_hssi_gen3_tx_pcs,
		output wire		out_blockselect_hssi_krfec_rx_pcs,
		output wire		out_blockselect_hssi_krfec_tx_pcs,
		output wire		out_blockselect_hssi_pipe_gen1_2,
		output wire		out_blockselect_hssi_pipe_gen3,
		output wire		out_blockselect_hssi_rx_pcs_pma_interface,
		output wire		out_blockselect_hssi_rx_pld_pcs_interface,
		output wire		out_blockselect_hssi_tx_pcs_pma_interface,
		output wire		out_blockselect_hssi_tx_pld_pcs_interface,
		output wire	[4:0]	out_bond_pcs10g_out_bot,
		output wire	[4:0]	out_bond_pcs10g_out_top,
		output wire	[12:0]	out_bond_pcs8g_out_bot,
		output wire	[12:0]	out_bond_pcs8g_out_top,
		output wire	[11:0]	out_bond_pmaif_out_bot,
		output wire	[11:0]	out_bond_pmaif_out_top,
		output wire	[2:0]	out_hip_clk_out,
		output wire	[7:0]	out_hip_ctrl_out,
		output wire		out_hip_iocsr_rdy,
		output wire		out_hip_iocsr_rdy_dly,
		output wire		out_hip_nfrzdrv,
		output wire		out_hip_npor,
		output wire	[50:0]	out_hip_rx_data,
		output wire		out_hip_usermode,
		output wire		out_pld_10g_krfec_rx_blk_lock,
		output wire	[1:0]	out_pld_10g_krfec_rx_diag_data_status,
		output wire		out_pld_10g_krfec_rx_frame,
		output wire		out_pld_10g_krfec_tx_frame,
		output wire		out_pld_10g_rx_align_val,
		output wire		out_pld_10g_rx_crc32_err,
		output wire		out_pld_10g_rx_data_valid,
		output wire		out_pld_10g_rx_empty,
		output wire		out_pld_10g_rx_fifo_del,
		output wire		out_pld_10g_rx_fifo_insert,
		output wire	[4:0]	out_pld_10g_rx_fifo_num,
		output wire		out_pld_10g_rx_frame_lock,
		output wire		out_pld_10g_rx_hi_ber,
		output wire		out_pld_10g_rx_oflw_err,
		output wire		out_pld_10g_rx_pempty,
		output wire		out_pld_10g_rx_pfull,
		output wire		out_pld_10g_tx_burst_en_exe,
		output wire		out_pld_10g_tx_empty,
		output wire	[3:0]	out_pld_10g_tx_fifo_num,
		output wire		out_pld_10g_tx_full,
		output wire		out_pld_10g_tx_pempty,
		output wire		out_pld_10g_tx_pfull,
		output wire		out_pld_10g_tx_wordslip_exe,
		output wire	[3:0]	out_pld_8g_a1a2_k1k2_flag,
		output wire		out_pld_8g_empty_rmf,
		output wire		out_pld_8g_empty_rx,
		output wire		out_pld_8g_empty_tx,
		output wire		out_pld_8g_full_rmf,
		output wire		out_pld_8g_full_rx,
		output wire		out_pld_8g_full_tx,
		output wire		out_pld_8g_rxelecidle,
		output wire		out_pld_8g_signal_detect_out,
		output wire	[4:0]	out_pld_8g_wa_boundary,
		output wire		out_pld_krfec_tx_alignment,
		output wire		out_pld_pcs_rx_clk_out,
		output wire		out_pld_pcs_tx_clk_out,
		output wire		out_pld_pma_adapt_done,
		output wire		out_pld_pma_clkdiv_rx_user,
		output wire		out_pld_pma_clkdiv_tx_user,
		output wire		out_pld_pma_clklow,
		output wire		out_pld_pma_fref,
		output wire		out_pld_pma_hclk,
		output wire	[1:0]	out_pld_pma_pcie_sw_done,
		output wire		out_pld_pma_pfdmode_lock,
		output wire	[4:0]	out_pld_pma_reserved_in,
		output wire		out_pld_pma_rx_clk_out,
		output wire		out_pld_pma_rx_detect_valid,
		output wire		out_pld_pma_rx_found,
		output wire		out_pld_pma_rxpll_lock,
		output wire		out_pld_pma_signal_ok,
		output wire	[7:0]	out_pld_pma_testbus,
		output wire		out_pld_pma_tx_clk_out,
		output wire		out_pld_pmaif_mask_tx_pll,
		output wire	[9:0]	out_pld_reserved_out,
		output wire	[19:0]	out_pld_rx_control,
		output wire	[127:0]	out_pld_rx_data,
		output wire		out_pld_rx_prbs_done,
		output wire		out_pld_rx_prbs_err,
		output wire	[19:0]	out_pld_test_data,
		output wire		out_pld_uhsif_lock,
		output wire		out_pld_uhsif_tx_clk_out,
		output wire		out_pma_adapt_start,
		output wire		out_pma_atpg_los_en_n,
		output wire		out_pma_csr_test_dis,
		output wire	[17:0]	out_pma_current_coeff,
		output wire	[2:0]	out_pma_current_rxpreset,
		output wire		out_pma_early_eios,
		output wire	[5:0]	out_pma_eye_monitor,
		output wire	[1:0]	out_pma_interface_select,
		output wire		out_pma_ltd_b,
		output wire		out_pma_ltr,
		output wire		out_pma_nfrzdrv,
		output wire		out_pma_nrpi_freeze,
		output wire	[1:0]	out_pma_pcie_switch,
		output wire		out_pma_ppm_lock,
		output wire	[4:0]	out_pma_reserved_out,
		output wire		out_pma_rs_lpbk_b,
		output wire		out_pma_rx_clkslip,
		output wire		out_pma_rx_qpi_pullup,
		output wire		out_pma_rxpma_rstb,
		output wire		out_pma_scan_mode_n,
		output wire		out_pma_scan_shift_n,
		output wire		out_pma_tx_bitslip,
		output wire		out_pma_tx_bonding_rstb,
		output wire		out_pma_tx_elec_idle,
		output wire	[63:0]	out_pma_tx_pma_data,
		output wire		out_pma_tx_qpi_pulldn,
		output wire		out_pma_tx_qpi_pullup,
		output wire		out_pma_tx_txdetectrx,
		output wire		out_pma_txpma_rstb
	//PORT_LIST_END
	);
	//wire declarations
	
	// wires for module twentynm_hssi_fifo_tx_pcs
	wire	[7:0]	w_hssi_fifo_tx_pcs_avmmreaddata;
	wire		w_hssi_fifo_tx_pcs_blockselect;
	wire	[72:0]	w_hssi_fifo_tx_pcs_data_out_10g;
	wire	[63:0]	w_hssi_fifo_tx_pcs_data_out_8g_phase_comp;
	
	// wires for module twentynm_hssi_gen3_rx_pcs
	wire	[7:0]	w_hssi_gen3_rx_pcs_avmmreaddata;
	wire		w_hssi_gen3_rx_pcs_blk_algnd_int;
	wire		w_hssi_gen3_rx_pcs_blk_start;
	wire		w_hssi_gen3_rx_pcs_blockselect;
	wire		w_hssi_gen3_rx_pcs_clkcomp_delete_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_insert_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_overfl_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_undfl_int;
	wire	[31:0]	w_hssi_gen3_rx_pcs_data_out;
	wire		w_hssi_gen3_rx_pcs_data_valid;
	wire		w_hssi_gen3_rx_pcs_ei_det_int;
	wire		w_hssi_gen3_rx_pcs_ei_partial_det_int;
	wire		w_hssi_gen3_rx_pcs_err_decode_int;
	wire		w_hssi_gen3_rx_pcs_i_det_int;
	wire		w_hssi_gen3_rx_pcs_lpbk_blk_start;
	wire	[33:0]	w_hssi_gen3_rx_pcs_lpbk_data;
	wire		w_hssi_gen3_rx_pcs_lpbk_data_valid;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk;
	wire	[39:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n;
	wire		w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int;
	wire	[19:0]	w_hssi_gen3_rx_pcs_rx_test_out;
	wire	[1:0]	w_hssi_gen3_rx_pcs_sync_hdr;
	
	// wires for module twentynm_hssi_krfec_tx_pcs
	wire	[7:0]	w_hssi_krfec_tx_pcs_avmmreaddata;
	wire		w_hssi_krfec_tx_pcs_blockselect;
	wire		w_hssi_krfec_tx_pcs_tx_alignment;
	wire	[63:0]	w_hssi_krfec_tx_pcs_tx_data_out;
	wire		w_hssi_krfec_tx_pcs_tx_frame;
	wire	[19:0]	w_hssi_krfec_tx_pcs_tx_test_data;
	
	// wires for module twentynm_hssi_krfec_rx_pcs
	wire	[7:0]	w_hssi_krfec_rx_pcs_avmmreaddata;
	wire		w_hssi_krfec_rx_pcs_blockselect;
	wire		w_hssi_krfec_rx_pcs_rx_block_lock;
	wire	[9:0]	w_hssi_krfec_rx_pcs_rx_control_out;
	wire	[63:0]	w_hssi_krfec_rx_pcs_rx_data_out;
	wire	[1:0]	w_hssi_krfec_rx_pcs_rx_data_status;
	wire		w_hssi_krfec_rx_pcs_rx_data_valid_out;
	wire		w_hssi_krfec_rx_pcs_rx_frame;
	wire		w_hssi_krfec_rx_pcs_rx_signal_ok_out;
	
	// wires for module twentynm_hssi_rx_pld_pcs_interface
	wire	[7:0]	w_hssi_rx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_rx_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_hip_rx_ctrl;
	wire	[50:0]	w_hssi_rx_pld_pcs_interface_hip_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
	wire	[3:0]	w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary;
	wire		w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_pld_rx_control;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_pld_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
	
	// wires for module twentynm_hssi_common_pld_pcs_interface
	wire	[7:0]	w_hssi_common_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_common_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_hip_cmn_clk;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_hip_cmn_ctrl;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
	wire		w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_hip_npor;
	wire		w_hssi_common_pld_pcs_interface_hip_usermode;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n;
	wire	[17:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel;
	wire		w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_clklow;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_fref;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_hclk;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_pld_pma_reserved_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
	wire	[7:0]	w_hssi_common_pld_pcs_interface_pld_pma_testbus;
	wire		w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
	wire	[9:0]	w_hssi_common_pld_pcs_interface_pld_reserved_out;
	wire	[19:0]	w_hssi_common_pld_pcs_interface_pld_test_data;
	wire		w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
	wire		w_hssi_common_pld_pcs_interface_scan_mode_n;
	
	// wires for module twentynm_hssi_10g_rx_pcs
	wire	[7:0]	w_hssi_10g_rx_pcs_avmmreaddata;
	wire		w_hssi_10g_rx_pcs_blockselect;
	wire		w_hssi_10g_rx_pcs_rx_align_val;
	wire		w_hssi_10g_rx_pcs_rx_blk_lock;
	wire		w_hssi_10g_rx_pcs_rx_clk_out;
	wire		w_hssi_10g_rx_pcs_rx_clk_out_pld_if;
	wire	[19:0]	w_hssi_10g_rx_pcs_rx_control;
	wire		w_hssi_10g_rx_pcs_rx_crc32_err;
	wire	[127:0]	w_hssi_10g_rx_pcs_rx_data;
	wire		w_hssi_10g_rx_pcs_rx_data_valid;
	wire		w_hssi_10g_rx_pcs_rx_dft_clk_out;
	wire	[1:0]	w_hssi_10g_rx_pcs_rx_diag_status;
	wire		w_hssi_10g_rx_pcs_rx_empty;
	wire		w_hssi_10g_rx_pcs_rx_fec_clk;
	wire		w_hssi_10g_rx_pcs_rx_fifo_del;
	wire		w_hssi_10g_rx_pcs_rx_fifo_insert;
	wire	[4:0]	w_hssi_10g_rx_pcs_rx_fifo_num;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_clk;
	wire	[73:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_data;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_en;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_ptr;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_frame_lock;
	wire		w_hssi_10g_rx_pcs_rx_hi_ber;
	wire		w_hssi_10g_rx_pcs_rx_master_clk;
	wire		w_hssi_10g_rx_pcs_rx_master_clk_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_oflw_err;
	wire		w_hssi_10g_rx_pcs_rx_pempty;
	wire		w_hssi_10g_rx_pcs_rx_pfull;
	wire		w_hssi_10g_rx_pcs_rx_random_err;
	wire		w_hssi_10g_rx_pcs_rx_rx_frame;
	
	// wires for module twentynm_hssi_tx_pld_pcs_interface
	wire	[7:0]	w_hssi_tx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_tx_pld_pcs_interface_blockselect;
	wire		w_hssi_tx_pld_pcs_interface_hip_tx_clk;
	wire	[6:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en;
	wire	[17:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control;
	wire	[8:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg;
	wire	[127:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start;
	wire	[4:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle;
	wire	[2:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
	wire		w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
	
	// wires for module twentynm_hssi_tx_pcs_pma_interface
	wire	[7:0]	w_hssi_tx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_tx_pcs_pma_interface_blockselect;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out;
	wire	[4:0]	w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk;
	wire		w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_pma_tx_pma_data;
	wire		w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_1;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_2;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_3;
	
	// wires for module twentynm_hssi_rx_pcs_pma_interface
	wire	[7:0]	w_hssi_rx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_rx_pcs_pma_interface_blockselect;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni;
	wire	[31:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok;
	wire		w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk;
	wire	[5:0]	w_hssi_rx_pcs_pma_interface_pma_eye_monitor;
	wire		w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
	wire		w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test;
	
	// wires for module twentynm_hssi_10g_tx_pcs
	wire	[7:0]	w_hssi_10g_tx_pcs_avmmreaddata;
	wire		w_hssi_10g_tx_pcs_blockselect;
	wire		w_hssi_10g_tx_pcs_distdwn_out_dv;
	wire		w_hssi_10g_tx_pcs_distdwn_out_rden;
	wire		w_hssi_10g_tx_pcs_distdwn_out_wren;
	wire		w_hssi_10g_tx_pcs_distup_out_dv;
	wire		w_hssi_10g_tx_pcs_distup_out_rden;
	wire		w_hssi_10g_tx_pcs_distup_out_wren;
	wire		w_hssi_10g_tx_pcs_tx_burst_en_exe;
	wire		w_hssi_10g_tx_pcs_tx_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pma_if;
	wire	[8:0]	w_hssi_10g_tx_pcs_tx_control_out_krfec;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_data_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_data_valid_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_dft_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_empty;
	wire		w_hssi_10g_tx_pcs_tx_fec_clk;
	wire	[3:0]	w_hssi_10g_tx_pcs_tx_fifo_num;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_rd_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_clk;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_en;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_frame;
	wire		w_hssi_10g_tx_pcs_tx_full;
	wire		w_hssi_10g_tx_pcs_tx_master_clk;
	wire		w_hssi_10g_tx_pcs_tx_master_clk_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_pempty;
	wire		w_hssi_10g_tx_pcs_tx_pfull;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_data;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_gating_val;
	wire	[19:0]	w_hssi_10g_tx_pcs_tx_test_data;
	wire		w_hssi_10g_tx_pcs_tx_wordslip_exe;
	
	// wires for module twentynm_hssi_8g_tx_pcs
	wire	[7:0]	w_hssi_8g_tx_pcs_avmmreaddata;
	wire		w_hssi_8g_tx_pcs_blockselect;
	wire		w_hssi_8g_tx_pcs_clk_out;
	wire		w_hssi_8g_tx_pcs_clk_out_gen3;
	wire	[19:0]	w_hssi_8g_tx_pcs_dataout;
	wire		w_hssi_8g_tx_pcs_dyn_clk_switch_n;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn;
	wire		w_hssi_8g_tx_pcs_g3_tx_pma_rstn;
	wire	[2:0]	w_hssi_8g_tx_pcs_non_gray_eidleinfersel;
	wire		w_hssi_8g_tx_pcs_ph_fifo_overflow;
	wire		w_hssi_8g_tx_pcs_ph_fifo_underflow;
	wire		w_hssi_8g_tx_pcs_phfifo_txdeemph;
	wire	[2:0]	w_hssi_8g_tx_pcs_phfifo_txmargin;
	wire		w_hssi_8g_tx_pcs_phfifo_txswing;
	wire		w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out;
	wire	[1:0]	w_hssi_8g_tx_pcs_pipe_power_down_out;
	wire		w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3;
	wire		w_hssi_8g_tx_pcs_pmaif_asn_rstn;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_refclk_b;
	wire		w_hssi_8g_tx_pcs_refclk_b_reset;
	wire		w_hssi_8g_tx_pcs_rxpolarity_int;
	wire		w_hssi_8g_tx_pcs_soft_reset_wclk1_n;
	wire		w_hssi_8g_tx_pcs_sw_fifo_wr_clk;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_blk_start_out;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_ctrlplane_testbus;
	wire	[31:0]	w_hssi_8g_tx_pcs_tx_data_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_data_valid_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_datak_out;
	wire		w_hssi_8g_tx_pcs_tx_detect_rxloopback_int;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_tx_pipe_clk;
	wire		w_hssi_8g_tx_pcs_tx_pipe_electidle;
	wire		w_hssi_8g_tx_pcs_tx_pipe_soft_reset;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_sync_hdr_out;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_testbus;
	wire		w_hssi_8g_tx_pcs_txcompliance_out;
	wire		w_hssi_8g_tx_pcs_txelecidle_out;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk;
	wire	[63:0]	w_hssi_8g_tx_pcs_wr_data_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_en_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo;
	
	// wires for module twentynm_hssi_pipe_gen3
	wire	[7:0]	w_hssi_pipe_gen3_avmmreaddata;
	wire		w_hssi_pipe_gen3_blockselect;
	wire		w_hssi_pipe_gen3_gen3_clk_sel;
	wire		w_hssi_pipe_gen3_pcs_rst;
	wire		w_hssi_pipe_gen3_phystatus;
	wire	[17:0]	w_hssi_pipe_gen3_pma_current_coeff;
	wire	[2:0]	w_hssi_pipe_gen3_pma_current_rxpreset;
	wire		w_hssi_pipe_gen3_pma_tx_elec_idle;
	wire		w_hssi_pipe_gen3_pma_txdetectrx;
	wire		w_hssi_pipe_gen3_rev_lpbk_8gpcs_out;
	wire		w_hssi_pipe_gen3_rev_lpbk_int;
	wire	[3:0]	w_hssi_pipe_gen3_rx_blk_start;
	wire	[1:0]	w_hssi_pipe_gen3_rx_sync_hdr;
	wire	[63:0]	w_hssi_pipe_gen3_rxd_8gpcs_out;
	wire	[3:0]	w_hssi_pipe_gen3_rxdataskip;
	wire		w_hssi_pipe_gen3_rxelecidle;
	wire		w_hssi_pipe_gen3_rxpolarity_8gpcs_out;
	wire		w_hssi_pipe_gen3_rxpolarity_int;
	wire	[2:0]	w_hssi_pipe_gen3_rxstatus;
	wire		w_hssi_pipe_gen3_rxvalid;
	wire		w_hssi_pipe_gen3_shutdown_clk;
	wire	[19:0]	w_hssi_pipe_gen3_test_out;
	wire		w_hssi_pipe_gen3_tx_blk_start_int;
	wire	[1:0]	w_hssi_pipe_gen3_tx_sync_hdr_int;
	wire	[31:0]	w_hssi_pipe_gen3_txdata_int;
	wire	[3:0]	w_hssi_pipe_gen3_txdatak_int;
	wire		w_hssi_pipe_gen3_txdataskip_int;
	
	// wires for module twentynm_hssi_pipe_gen1_2
	wire	[7:0]	w_hssi_pipe_gen1_2_avmmreaddata;
	wire		w_hssi_pipe_gen1_2_blockselect;
	wire	[17:0]	w_hssi_pipe_gen1_2_current_coeff;
	wire		w_hssi_pipe_gen1_2_phystatus;
	wire		w_hssi_pipe_gen1_2_polarity_inversion_rx;
	wire		w_hssi_pipe_gen1_2_rev_loopbk;
	wire		w_hssi_pipe_gen1_2_rxelecidle;
	wire		w_hssi_pipe_gen1_2_rxelectricalidle_out;
	wire	[2:0]	w_hssi_pipe_gen1_2_rxstatus;
	wire		w_hssi_pipe_gen1_2_rxvalid;
	wire		w_hssi_pipe_gen1_2_tx_elec_idle_out;
	wire		w_hssi_pipe_gen1_2_txdetectrx;
	
	// wires for module twentynm_hssi_gen3_tx_pcs
	wire	[7:0]	w_hssi_gen3_tx_pcs_avmmreaddata;
	wire		w_hssi_gen3_tx_pcs_blockselect;
	wire	[31:0]	w_hssi_gen3_tx_pcs_data_out;
	wire	[35:0]	w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out;
	wire	[31:0]	w_hssi_gen3_tx_pcs_par_lpbk_out;
	wire	[19:0]	w_hssi_gen3_tx_pcs_tx_test_out;
	
	// wires for module twentynm_hssi_8g_rx_pcs
	wire	[3:0]	w_hssi_8g_rx_pcs_a1a2k1k2flag;
	wire	[7:0]	w_hssi_8g_rx_pcs_avmmreaddata;
	wire		w_hssi_8g_rx_pcs_blockselect;
	wire	[19:0]	w_hssi_8g_rx_pcs_chnl_test_bus_out;
	wire		w_hssi_8g_rx_pcs_clock_to_pld;
	wire	[63:0]	w_hssi_8g_rx_pcs_dataout;
	wire		w_hssi_8g_rx_pcs_dis_pc_byte;
	wire		w_hssi_8g_rx_pcs_eidle_detected;
	wire	[2:0]	w_hssi_8g_rx_pcs_eios_det_cdr_ctrl;
	wire		w_hssi_8g_rx_pcs_g3_rx_pma_rstn;
	wire		w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn;
	wire		w_hssi_8g_rx_pcs_gen2ngen1;
	wire	[19:0]	w_hssi_8g_rx_pcs_parallel_rev_loopback;
	wire		w_hssi_8g_rx_pcs_pc_fifo_empty;
	wire		w_hssi_8g_rx_pcs_pcfifofull;
	wire		w_hssi_8g_rx_pcs_phystatus;
	wire	[63:0]	w_hssi_8g_rx_pcs_pipe_data;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_up;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo;
	wire	[7:0]	w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rm_fifo_empty;
	wire		w_hssi_8g_rx_pcs_rm_fifo_full;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_blk_start;
	wire		w_hssi_8g_rx_pcs_rx_clk_out_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clkslip;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_data_valid;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rx_pipe_clk;
	wire		w_hssi_8g_rx_pcs_rx_pipe_soft_reset;
	wire		w_hssi_8g_rx_pcs_rx_pma_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_sync_hdr;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_up;
	wire	[2:0]	w_hssi_8g_rx_pcs_rxstatus;
	wire		w_hssi_8g_rx_pcs_rxvalid;
	wire		w_hssi_8g_rx_pcs_signal_detect_out;
	wire	[4:0]	w_hssi_8g_rx_pcs_word_align_boundary;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk;
	wire	[79:0]	w_hssi_8g_rx_pcs_wr_data_rx_phfifo;
	wire	[31:0]	w_hssi_8g_rx_pcs_wr_data_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo;
	
	// wires for module twentynm_hssi_fifo_rx_pcs
	wire	[7:0]	w_hssi_fifo_rx_pcs_avmmreaddata;
	wire		w_hssi_fifo_rx_pcs_blockselect;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out2_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out_8g_clock_comp;
	wire	[79:0]	w_hssi_fifo_rx_pcs_data_out_8g_phase_comp;
	wire	[39:0]	w_hssi_fifo_rx_pcs_data_out_gen3;
	
	// wires for module twentynm_hssi_common_pcs_pma_interface
	wire	[7:0]	w_hssi_common_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_common_pcs_pma_interface_blockselect;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in;
	wire	[19:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out;
	wire	[7:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus;
	wire		w_hssi_common_pcs_pma_interface_pma_adapt_start;
	wire		w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
	wire		w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
	wire	[17:0]	w_hssi_common_pcs_pma_interface_pma_current_coeff;
	wire	[2:0]	w_hssi_common_pcs_pma_interface_pma_current_rxpreset;
	wire		w_hssi_common_pcs_pma_interface_pma_early_eios;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_interface_select;
	wire		w_hssi_common_pcs_pma_interface_pma_ltd_b;
	wire		w_hssi_common_pcs_pma_interface_pma_ltr;
	wire		w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
	wire		w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_pcie_switch;
	wire		w_hssi_common_pcs_pma_interface_pma_ppm_lock;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_pma_reserved_out;
	wire		w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
	wire		w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up;
	
	
	generate
		
		//module instantiations
		
		// instantiating twentynm_hssi_10g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_rx_pcs
			twentynm_hssi_10g_rx_pcs #(
				.advanced_user_mode(hssi_10g_rx_pcs_advanced_user_mode),
				.align_del(hssi_10g_rx_pcs_align_del),
				.ber_bit_err_total_cnt(hssi_10g_rx_pcs_ber_bit_err_total_cnt),
				.ber_clken(hssi_10g_rx_pcs_ber_clken),
				.ber_xus_timer_window(hssi_10g_rx_pcs_ber_xus_timer_window),
				.bitslip_mode(hssi_10g_rx_pcs_bitslip_mode),
				.blksync_bitslip_type(hssi_10g_rx_pcs_blksync_bitslip_type),
				.blksync_bitslip_wait_cnt(hssi_10g_rx_pcs_blksync_bitslip_wait_cnt),
				.blksync_bitslip_wait_type(hssi_10g_rx_pcs_blksync_bitslip_wait_type),
				.blksync_bypass(hssi_10g_rx_pcs_blksync_bypass),
				.blksync_clken(hssi_10g_rx_pcs_blksync_clken),
				.blksync_enum_invalid_sh_cnt(hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt),
				.blksync_knum_sh_cnt_postlock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock),
				.blksync_knum_sh_cnt_prelock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock),
				.blksync_pipeln(hssi_10g_rx_pcs_blksync_pipeln),
				.clr_errblk_cnt_en(hssi_10g_rx_pcs_clr_errblk_cnt_en),
				.control_del(hssi_10g_rx_pcs_control_del),
				.crcchk_bypass(hssi_10g_rx_pcs_crcchk_bypass),
				.crcchk_clken(hssi_10g_rx_pcs_crcchk_clken),
				.crcchk_inv(hssi_10g_rx_pcs_crcchk_inv),
				.crcchk_pipeln(hssi_10g_rx_pcs_crcchk_pipeln),
				.crcflag_pipeln(hssi_10g_rx_pcs_crcflag_pipeln),
				.ctrl_bit_reverse(hssi_10g_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_10g_rx_pcs_data_bit_reverse),
				.dec64b66b_clken(hssi_10g_rx_pcs_dec64b66b_clken),
				.dec_64b66b_rxsm_bypass(hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass),
				.descrm_bypass(hssi_10g_rx_pcs_descrm_bypass),
				.descrm_clken(hssi_10g_rx_pcs_descrm_clken),
				.descrm_mode(hssi_10g_rx_pcs_descrm_mode),
				.descrm_pipeln(hssi_10g_rx_pcs_descrm_pipeln),
				.dft_clk_out_sel(hssi_10g_rx_pcs_dft_clk_out_sel),
				.dis_signal_ok(hssi_10g_rx_pcs_dis_signal_ok),
				.dispchk_bypass(hssi_10g_rx_pcs_dispchk_bypass),
				.empty_flag_type(hssi_10g_rx_pcs_empty_flag_type),
				.fast_path(hssi_10g_rx_pcs_fast_path),
				.fec_clken(hssi_10g_rx_pcs_fec_clken),
				.fec_enable(hssi_10g_rx_pcs_fec_enable),
				.fifo_double_read(hssi_10g_rx_pcs_fifo_double_read),
				.fifo_stop_rd(hssi_10g_rx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_rx_pcs_fifo_stop_wr),
				.force_align(hssi_10g_rx_pcs_force_align),
				.frmsync_bypass(hssi_10g_rx_pcs_frmsync_bypass),
				.frmsync_clken(hssi_10g_rx_pcs_frmsync_clken),
				.frmsync_enum_scrm(hssi_10g_rx_pcs_frmsync_enum_scrm),
				.frmsync_enum_sync(hssi_10g_rx_pcs_frmsync_enum_sync),
				.frmsync_flag_type(hssi_10g_rx_pcs_frmsync_flag_type),
				.frmsync_knum_sync(hssi_10g_rx_pcs_frmsync_knum_sync),
				.frmsync_mfrm_length(hssi_10g_rx_pcs_frmsync_mfrm_length),
				.frmsync_pipeln(hssi_10g_rx_pcs_frmsync_pipeln),
				.full_flag_type(hssi_10g_rx_pcs_full_flag_type),
				.gb_rx_idwidth(hssi_10g_rx_pcs_gb_rx_idwidth),
				.gb_rx_odwidth(hssi_10g_rx_pcs_gb_rx_odwidth),
				.gbexp_clken(hssi_10g_rx_pcs_gbexp_clken),
				.low_latency_en(hssi_10g_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_10g_rx_pcs_lpbk_mode),
				.master_clk_sel(hssi_10g_rx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_rx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_rx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_rx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_rx_pcs_pld_if_type),
				.prot_mode(hssi_10g_rx_pcs_prot_mode),
				.rand_clken(hssi_10g_rx_pcs_rand_clken),
				.rd_clk_sel(hssi_10g_rx_pcs_rd_clk_sel),
				.rdfifo_clken(hssi_10g_rx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_rx_pcs_reconfig_settings),
				.rx_fifo_write_ctrl(hssi_10g_rx_pcs_rx_fifo_write_ctrl),
				.rx_scrm_width(hssi_10g_rx_pcs_rx_scrm_width),
				.rx_sh_location(hssi_10g_rx_pcs_rx_sh_location),
				.rx_signal_ok_sel(hssi_10g_rx_pcs_rx_signal_ok_sel),
				.rx_sm_bypass(hssi_10g_rx_pcs_rx_sm_bypass),
				.rx_sm_hiber(hssi_10g_rx_pcs_rx_sm_hiber),
				.rx_sm_pipeln(hssi_10g_rx_pcs_rx_sm_pipeln),
				.rx_testbus_sel(hssi_10g_rx_pcs_rx_testbus_sel),
				.rx_true_b2b(hssi_10g_rx_pcs_rx_true_b2b),
				.rxfifo_empty(hssi_10g_rx_pcs_rxfifo_empty),
				.rxfifo_full(hssi_10g_rx_pcs_rxfifo_full),
				.rxfifo_mode(hssi_10g_rx_pcs_rxfifo_mode),
				.rxfifo_pempty(hssi_10g_rx_pcs_rxfifo_pempty),
				.rxfifo_pfull(hssi_10g_rx_pcs_rxfifo_pfull),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.stretch_num_stages(hssi_10g_rx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_rx_pcs_sup_mode),
				.test_mode(hssi_10g_rx_pcs_test_mode),
				.wrfifo_clken(hssi_10g_rx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_rx_pcs_blockselect),
				.rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.rx_control(w_hssi_10g_rx_pcs_rx_control),
				.rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.rx_data(w_hssi_10g_rx_pcs_rx_data),
				.rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.rx_diag_status(w_hssi_10g_rx_pcs_rx_diag_status),
				.rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.rx_fec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.rx_fifo_num(w_hssi_10g_rx_pcs_rx_fifo_num),
				.rx_fifo_rd_ptr(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr),
				.rx_fifo_rd_ptr2(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2),
				.rx_fifo_wr_clk(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.rx_fifo_wr_data(w_hssi_10g_rx_pcs_rx_fifo_wr_data),
				.rx_fifo_wr_en(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.rx_fifo_wr_ptr(w_hssi_10g_rx_pcs_rx_fifo_wr_ptr),
				.rx_fifo_wr_rst_n(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.rx_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_rx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_rx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.rx_control_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0]}),
				.rx_control_in_krfec({w_hssi_krfec_rx_pcs_rx_control_out[9], w_hssi_krfec_rx_pcs_rx_control_out[8], w_hssi_krfec_rx_pcs_rx_control_out[7], w_hssi_krfec_rx_pcs_rx_control_out[6], w_hssi_krfec_rx_pcs_rx_control_out[5], w_hssi_krfec_rx_pcs_rx_control_out[4], w_hssi_krfec_rx_pcs_rx_control_out[3], w_hssi_krfec_rx_pcs_rx_control_out[2], w_hssi_krfec_rx_pcs_rx_control_out[1], w_hssi_krfec_rx_pcs_rx_control_out[0]}),
				.rx_data_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0]}),
				.rx_data_in_krfec({w_hssi_krfec_rx_pcs_rx_data_out[63], w_hssi_krfec_rx_pcs_rx_data_out[62], w_hssi_krfec_rx_pcs_rx_data_out[61], w_hssi_krfec_rx_pcs_rx_data_out[60], w_hssi_krfec_rx_pcs_rx_data_out[59], w_hssi_krfec_rx_pcs_rx_data_out[58], w_hssi_krfec_rx_pcs_rx_data_out[57], w_hssi_krfec_rx_pcs_rx_data_out[56], w_hssi_krfec_rx_pcs_rx_data_out[55], w_hssi_krfec_rx_pcs_rx_data_out[54], w_hssi_krfec_rx_pcs_rx_data_out[53], w_hssi_krfec_rx_pcs_rx_data_out[52], w_hssi_krfec_rx_pcs_rx_data_out[51], w_hssi_krfec_rx_pcs_rx_data_out[50], w_hssi_krfec_rx_pcs_rx_data_out[49], w_hssi_krfec_rx_pcs_rx_data_out[48], w_hssi_krfec_rx_pcs_rx_data_out[47], w_hssi_krfec_rx_pcs_rx_data_out[46], w_hssi_krfec_rx_pcs_rx_data_out[45], w_hssi_krfec_rx_pcs_rx_data_out[44], w_hssi_krfec_rx_pcs_rx_data_out[43], w_hssi_krfec_rx_pcs_rx_data_out[42], w_hssi_krfec_rx_pcs_rx_data_out[41], w_hssi_krfec_rx_pcs_rx_data_out[40], w_hssi_krfec_rx_pcs_rx_data_out[39], w_hssi_krfec_rx_pcs_rx_data_out[38], w_hssi_krfec_rx_pcs_rx_data_out[37], w_hssi_krfec_rx_pcs_rx_data_out[36], w_hssi_krfec_rx_pcs_rx_data_out[35], w_hssi_krfec_rx_pcs_rx_data_out[34], w_hssi_krfec_rx_pcs_rx_data_out[33], w_hssi_krfec_rx_pcs_rx_data_out[32], w_hssi_krfec_rx_pcs_rx_data_out[31], w_hssi_krfec_rx_pcs_rx_data_out[30], w_hssi_krfec_rx_pcs_rx_data_out[29], w_hssi_krfec_rx_pcs_rx_data_out[28], w_hssi_krfec_rx_pcs_rx_data_out[27], w_hssi_krfec_rx_pcs_rx_data_out[26], w_hssi_krfec_rx_pcs_rx_data_out[25], w_hssi_krfec_rx_pcs_rx_data_out[24], w_hssi_krfec_rx_pcs_rx_data_out[23], w_hssi_krfec_rx_pcs_rx_data_out[22], w_hssi_krfec_rx_pcs_rx_data_out[21], w_hssi_krfec_rx_pcs_rx_data_out[20], w_hssi_krfec_rx_pcs_rx_data_out[19], w_hssi_krfec_rx_pcs_rx_data_out[18], w_hssi_krfec_rx_pcs_rx_data_out[17], w_hssi_krfec_rx_pcs_rx_data_out[16], w_hssi_krfec_rx_pcs_rx_data_out[15], w_hssi_krfec_rx_pcs_rx_data_out[14], w_hssi_krfec_rx_pcs_rx_data_out[13], w_hssi_krfec_rx_pcs_rx_data_out[12], w_hssi_krfec_rx_pcs_rx_data_out[11], w_hssi_krfec_rx_pcs_rx_data_out[10], w_hssi_krfec_rx_pcs_rx_data_out[9], w_hssi_krfec_rx_pcs_rx_data_out[8], w_hssi_krfec_rx_pcs_rx_data_out[7], w_hssi_krfec_rx_pcs_rx_data_out[6], w_hssi_krfec_rx_pcs_rx_data_out[5], w_hssi_krfec_rx_pcs_rx_data_out[4], w_hssi_krfec_rx_pcs_rx_data_out[3], w_hssi_krfec_rx_pcs_rx_data_out[2], w_hssi_krfec_rx_pcs_rx_data_out[1], w_hssi_krfec_rx_pcs_rx_data_out[0]}),
				.rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.rx_data_valid_in_krfec(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_10g[73], w_hssi_fifo_rx_pcs_data_out_10g[72], w_hssi_fifo_rx_pcs_data_out_10g[71], w_hssi_fifo_rx_pcs_data_out_10g[70], w_hssi_fifo_rx_pcs_data_out_10g[69], w_hssi_fifo_rx_pcs_data_out_10g[68], w_hssi_fifo_rx_pcs_data_out_10g[67], w_hssi_fifo_rx_pcs_data_out_10g[66], w_hssi_fifo_rx_pcs_data_out_10g[65], w_hssi_fifo_rx_pcs_data_out_10g[64], w_hssi_fifo_rx_pcs_data_out_10g[63], w_hssi_fifo_rx_pcs_data_out_10g[62], w_hssi_fifo_rx_pcs_data_out_10g[61], w_hssi_fifo_rx_pcs_data_out_10g[60], w_hssi_fifo_rx_pcs_data_out_10g[59], w_hssi_fifo_rx_pcs_data_out_10g[58], w_hssi_fifo_rx_pcs_data_out_10g[57], w_hssi_fifo_rx_pcs_data_out_10g[56], w_hssi_fifo_rx_pcs_data_out_10g[55], w_hssi_fifo_rx_pcs_data_out_10g[54], w_hssi_fifo_rx_pcs_data_out_10g[53], w_hssi_fifo_rx_pcs_data_out_10g[52], w_hssi_fifo_rx_pcs_data_out_10g[51], w_hssi_fifo_rx_pcs_data_out_10g[50], w_hssi_fifo_rx_pcs_data_out_10g[49], w_hssi_fifo_rx_pcs_data_out_10g[48], w_hssi_fifo_rx_pcs_data_out_10g[47], w_hssi_fifo_rx_pcs_data_out_10g[46], w_hssi_fifo_rx_pcs_data_out_10g[45], w_hssi_fifo_rx_pcs_data_out_10g[44], w_hssi_fifo_rx_pcs_data_out_10g[43], w_hssi_fifo_rx_pcs_data_out_10g[42], w_hssi_fifo_rx_pcs_data_out_10g[41], w_hssi_fifo_rx_pcs_data_out_10g[40], w_hssi_fifo_rx_pcs_data_out_10g[39], w_hssi_fifo_rx_pcs_data_out_10g[38], w_hssi_fifo_rx_pcs_data_out_10g[37], w_hssi_fifo_rx_pcs_data_out_10g[36], w_hssi_fifo_rx_pcs_data_out_10g[35], w_hssi_fifo_rx_pcs_data_out_10g[34], w_hssi_fifo_rx_pcs_data_out_10g[33], w_hssi_fifo_rx_pcs_data_out_10g[32], w_hssi_fifo_rx_pcs_data_out_10g[31], w_hssi_fifo_rx_pcs_data_out_10g[30], w_hssi_fifo_rx_pcs_data_out_10g[29], w_hssi_fifo_rx_pcs_data_out_10g[28], w_hssi_fifo_rx_pcs_data_out_10g[27], w_hssi_fifo_rx_pcs_data_out_10g[26], w_hssi_fifo_rx_pcs_data_out_10g[25], w_hssi_fifo_rx_pcs_data_out_10g[24], w_hssi_fifo_rx_pcs_data_out_10g[23], w_hssi_fifo_rx_pcs_data_out_10g[22], w_hssi_fifo_rx_pcs_data_out_10g[21], w_hssi_fifo_rx_pcs_data_out_10g[20], w_hssi_fifo_rx_pcs_data_out_10g[19], w_hssi_fifo_rx_pcs_data_out_10g[18], w_hssi_fifo_rx_pcs_data_out_10g[17], w_hssi_fifo_rx_pcs_data_out_10g[16], w_hssi_fifo_rx_pcs_data_out_10g[15], w_hssi_fifo_rx_pcs_data_out_10g[14], w_hssi_fifo_rx_pcs_data_out_10g[13], w_hssi_fifo_rx_pcs_data_out_10g[12], w_hssi_fifo_rx_pcs_data_out_10g[11], w_hssi_fifo_rx_pcs_data_out_10g[10], w_hssi_fifo_rx_pcs_data_out_10g[9], w_hssi_fifo_rx_pcs_data_out_10g[8], w_hssi_fifo_rx_pcs_data_out_10g[7], w_hssi_fifo_rx_pcs_data_out_10g[6], w_hssi_fifo_rx_pcs_data_out_10g[5], w_hssi_fifo_rx_pcs_data_out_10g[4], w_hssi_fifo_rx_pcs_data_out_10g[3], w_hssi_fifo_rx_pcs_data_out_10g[2], w_hssi_fifo_rx_pcs_data_out_10g[1], w_hssi_fifo_rx_pcs_data_out_10g[0]}),
				.rx_fifo_rd_data_dw({w_hssi_fifo_rx_pcs_data_out2_10g[73], w_hssi_fifo_rx_pcs_data_out2_10g[72], w_hssi_fifo_rx_pcs_data_out2_10g[71], w_hssi_fifo_rx_pcs_data_out2_10g[70], w_hssi_fifo_rx_pcs_data_out2_10g[69], w_hssi_fifo_rx_pcs_data_out2_10g[68], w_hssi_fifo_rx_pcs_data_out2_10g[67], w_hssi_fifo_rx_pcs_data_out2_10g[66], w_hssi_fifo_rx_pcs_data_out2_10g[65], w_hssi_fifo_rx_pcs_data_out2_10g[64], w_hssi_fifo_rx_pcs_data_out2_10g[63], w_hssi_fifo_rx_pcs_data_out2_10g[62], w_hssi_fifo_rx_pcs_data_out2_10g[61], w_hssi_fifo_rx_pcs_data_out2_10g[60], w_hssi_fifo_rx_pcs_data_out2_10g[59], w_hssi_fifo_rx_pcs_data_out2_10g[58], w_hssi_fifo_rx_pcs_data_out2_10g[57], w_hssi_fifo_rx_pcs_data_out2_10g[56], w_hssi_fifo_rx_pcs_data_out2_10g[55], w_hssi_fifo_rx_pcs_data_out2_10g[54], w_hssi_fifo_rx_pcs_data_out2_10g[53], w_hssi_fifo_rx_pcs_data_out2_10g[52], w_hssi_fifo_rx_pcs_data_out2_10g[51], w_hssi_fifo_rx_pcs_data_out2_10g[50], w_hssi_fifo_rx_pcs_data_out2_10g[49], w_hssi_fifo_rx_pcs_data_out2_10g[48], w_hssi_fifo_rx_pcs_data_out2_10g[47], w_hssi_fifo_rx_pcs_data_out2_10g[46], w_hssi_fifo_rx_pcs_data_out2_10g[45], w_hssi_fifo_rx_pcs_data_out2_10g[44], w_hssi_fifo_rx_pcs_data_out2_10g[43], w_hssi_fifo_rx_pcs_data_out2_10g[42], w_hssi_fifo_rx_pcs_data_out2_10g[41], w_hssi_fifo_rx_pcs_data_out2_10g[40], w_hssi_fifo_rx_pcs_data_out2_10g[39], w_hssi_fifo_rx_pcs_data_out2_10g[38], w_hssi_fifo_rx_pcs_data_out2_10g[37], w_hssi_fifo_rx_pcs_data_out2_10g[36], w_hssi_fifo_rx_pcs_data_out2_10g[35], w_hssi_fifo_rx_pcs_data_out2_10g[34], w_hssi_fifo_rx_pcs_data_out2_10g[33], w_hssi_fifo_rx_pcs_data_out2_10g[32], w_hssi_fifo_rx_pcs_data_out2_10g[31], w_hssi_fifo_rx_pcs_data_out2_10g[30], w_hssi_fifo_rx_pcs_data_out2_10g[29], w_hssi_fifo_rx_pcs_data_out2_10g[28], w_hssi_fifo_rx_pcs_data_out2_10g[27], w_hssi_fifo_rx_pcs_data_out2_10g[26], w_hssi_fifo_rx_pcs_data_out2_10g[25], w_hssi_fifo_rx_pcs_data_out2_10g[24], w_hssi_fifo_rx_pcs_data_out2_10g[23], w_hssi_fifo_rx_pcs_data_out2_10g[22], w_hssi_fifo_rx_pcs_data_out2_10g[21], w_hssi_fifo_rx_pcs_data_out2_10g[20], w_hssi_fifo_rx_pcs_data_out2_10g[19], w_hssi_fifo_rx_pcs_data_out2_10g[18], w_hssi_fifo_rx_pcs_data_out2_10g[17], w_hssi_fifo_rx_pcs_data_out2_10g[16], w_hssi_fifo_rx_pcs_data_out2_10g[15], w_hssi_fifo_rx_pcs_data_out2_10g[14], w_hssi_fifo_rx_pcs_data_out2_10g[13], w_hssi_fifo_rx_pcs_data_out2_10g[12], w_hssi_fifo_rx_pcs_data_out2_10g[11], w_hssi_fifo_rx_pcs_data_out2_10g[10], w_hssi_fifo_rx_pcs_data_out2_10g[9], w_hssi_fifo_rx_pcs_data_out2_10g[8], w_hssi_fifo_rx_pcs_data_out2_10g[7], w_hssi_fifo_rx_pcs_data_out2_10g[6], w_hssi_fifo_rx_pcs_data_out2_10g[5], w_hssi_fifo_rx_pcs_data_out2_10g[4], w_hssi_fifo_rx_pcs_data_out2_10g[3], w_hssi_fifo_rx_pcs_data_out2_10g[2], w_hssi_fifo_rx_pcs_data_out2_10g[1], w_hssi_fifo_rx_pcs_data_out2_10g[0]}),
				.rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.rx_pma_data({w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0]}),
				.rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.signal_ok_krfec(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_10g_reg(),
				.pld_10g_krfec_rx_blk_lock_10g_txclk_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_txclk_reg(),
				.pld_10g_krfec_rx_frame_10g_reg(),
				.pld_10g_krfec_rx_frame_10g_txclk_reg(),
				.pld_10g_krfec_rx_pld_rst_n_fifo(),
				.pld_10g_krfec_rx_pld_rst_n_reg(),
				.pld_10g_krfec_rx_pld_rst_n_txclk_reg(),
				.pld_10g_rx_align_clr_fifo(),
				.pld_10g_rx_align_clr_reg(),
				.pld_10g_rx_align_clr_txclk_reg(),
				.pld_10g_rx_align_val_fifo(),
				.pld_10g_rx_align_val_reg(),
				.pld_10g_rx_align_val_txclk_reg(),
				.pld_10g_rx_clr_ber_count_reg(),
				.pld_10g_rx_clr_ber_count_txclk_reg(),
				.pld_10g_rx_crc32_err_reg(),
				.pld_10g_rx_crc32_err_txclk_reg(),
				.pld_10g_rx_data_valid_10g_reg(),
				.pld_10g_rx_data_valid_fifo(),
				.pld_10g_rx_data_valid_pcsdirect_reg(),
				.pld_10g_rx_data_valid_txclk_reg(),
				.pld_10g_rx_empty_fifo(),
				.pld_10g_rx_fifo_del_reg(),
				.pld_10g_rx_fifo_del_txclk_reg(),
				.pld_10g_rx_fifo_insert_fifo(),
				.pld_10g_rx_fifo_num_reg(),
				.pld_10g_rx_fifo_num_txclk_reg(),
				.pld_10g_rx_frame_lock_reg(),
				.pld_10g_rx_frame_lock_txclk_reg(),
				.pld_10g_rx_hi_ber_reg(),
				.pld_10g_rx_hi_ber_txclk_reg(),
				.pld_10g_rx_oflw_err_reg(),
				.pld_10g_rx_oflw_err_txclk_reg(),
				.pld_10g_rx_pempty_fifo(),
				.pld_10g_rx_pfull_reg(),
				.pld_10g_rx_pfull_txclk_reg(),
				.pld_10g_rx_rd_en_fifo(),
				.pld_pcs_rx_clk_out_10g_txclk_wire(),
				.pld_pcs_rx_clk_out_10g_wire(),
				.pld_rx_control_10g_reg(),
				.pld_rx_control_10g_txclk_reg(),
				.pld_rx_data_10g_reg(),
				.pld_rx_data_10g_txclk_reg(),
				.pld_rx_prbs_err_10g_txclk_reg(),
				.pld_rx_prbs_err_clr_10g_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_10g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_align_val = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_blk_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_control[19:0] = 20'b0;
				assign w_hssi_10g_rx_pcs_rx_crc32_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_data[127:0] = 128'b0;
				assign w_hssi_10g_rx_pcs_rx_data_valid = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_dft_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_diag_status[1:0] = 2'b0;
				assign w_hssi_10g_rx_pcs_rx_empty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fec_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_del = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_insert = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_data[73:0] = 74'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_frame_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_hi_ber = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_oflw_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pempty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pfull = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_random_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_rx_frame = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_10g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_tx_pcs
			twentynm_hssi_10g_tx_pcs #(
				.advanced_user_mode(hssi_10g_tx_pcs_advanced_user_mode),
				.bitslip_en(hssi_10g_tx_pcs_bitslip_en),
				.bonding_dft_en(hssi_10g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_10g_tx_pcs_bonding_dft_val),
				.comp_cnt(hssi_10g_tx_pcs_comp_cnt),
				.compin_sel(hssi_10g_tx_pcs_compin_sel),
				.crcgen_bypass(hssi_10g_tx_pcs_crcgen_bypass),
				.crcgen_clken(hssi_10g_tx_pcs_crcgen_clken),
				.crcgen_err(hssi_10g_tx_pcs_crcgen_err),
				.crcgen_inv(hssi_10g_tx_pcs_crcgen_inv),
				.ctrl_bit_reverse(hssi_10g_tx_pcs_ctrl_bit_reverse),
				.ctrl_plane_bonding(hssi_10g_tx_pcs_ctrl_plane_bonding),
				.data_bit_reverse(hssi_10g_tx_pcs_data_bit_reverse),
				.dft_clk_out_sel(hssi_10g_tx_pcs_dft_clk_out_sel),
				.dispgen_bypass(hssi_10g_tx_pcs_dispgen_bypass),
				.dispgen_clken(hssi_10g_tx_pcs_dispgen_clken),
				.dispgen_err(hssi_10g_tx_pcs_dispgen_err),
				.dispgen_pipeln(hssi_10g_tx_pcs_dispgen_pipeln),
				.distdwn_bypass_pipeln(hssi_10g_tx_pcs_distdwn_bypass_pipeln),
				.distdwn_master(hssi_10g_tx_pcs_distdwn_master),
				.distup_bypass_pipeln(hssi_10g_tx_pcs_distup_bypass_pipeln),
				.distup_master(hssi_10g_tx_pcs_distup_master),
				.dv_bond(hssi_10g_tx_pcs_dv_bond),
				.empty_flag_type(hssi_10g_tx_pcs_empty_flag_type),
				.enc64b66b_txsm_clken(hssi_10g_tx_pcs_enc64b66b_txsm_clken),
				.enc_64b66b_txsm_bypass(hssi_10g_tx_pcs_enc_64b66b_txsm_bypass),
				.fastpath(hssi_10g_tx_pcs_fastpath),
				.fec_clken(hssi_10g_tx_pcs_fec_clken),
				.fec_enable(hssi_10g_tx_pcs_fec_enable),
				.fifo_double_write(hssi_10g_tx_pcs_fifo_double_write),
				.fifo_reg_fast(hssi_10g_tx_pcs_fifo_reg_fast),
				.fifo_stop_rd(hssi_10g_tx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_tx_pcs_fifo_stop_wr),
				.frmgen_burst(hssi_10g_tx_pcs_frmgen_burst),
				.frmgen_bypass(hssi_10g_tx_pcs_frmgen_bypass),
				.frmgen_clken(hssi_10g_tx_pcs_frmgen_clken),
				.frmgen_mfrm_length(hssi_10g_tx_pcs_frmgen_mfrm_length),
				.frmgen_pipeln(hssi_10g_tx_pcs_frmgen_pipeln),
				.frmgen_pyld_ins(hssi_10g_tx_pcs_frmgen_pyld_ins),
				.frmgen_wordslip(hssi_10g_tx_pcs_frmgen_wordslip),
				.full_flag_type(hssi_10g_tx_pcs_full_flag_type),
				.gb_pipeln_bypass(hssi_10g_tx_pcs_gb_pipeln_bypass),
				.gb_tx_idwidth(hssi_10g_tx_pcs_gb_tx_idwidth),
				.gb_tx_odwidth(hssi_10g_tx_pcs_gb_tx_odwidth),
				.gbred_clken(hssi_10g_tx_pcs_gbred_clken),
				.indv(hssi_10g_tx_pcs_indv),
				.low_latency_en(hssi_10g_tx_pcs_low_latency_en),
				.master_clk_sel(hssi_10g_tx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_tx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_tx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_tx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_tx_pcs_pld_if_type),
				.prot_mode(hssi_10g_tx_pcs_prot_mode),
				.pseudo_random(hssi_10g_tx_pcs_pseudo_random),
				.pseudo_seed_a(hssi_10g_tx_pcs_pseudo_seed_a),
				.pseudo_seed_b(hssi_10g_tx_pcs_pseudo_seed_b),
				.random_disp(hssi_10g_tx_pcs_random_disp),
				.rdfifo_clken(hssi_10g_tx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_tx_pcs_reconfig_settings),
				.scrm_bypass(hssi_10g_tx_pcs_scrm_bypass),
				.scrm_clken(hssi_10g_tx_pcs_scrm_clken),
				.scrm_mode(hssi_10g_tx_pcs_scrm_mode),
				.scrm_pipeln(hssi_10g_tx_pcs_scrm_pipeln),
				.sh_err(hssi_10g_tx_pcs_sh_err),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sop_mark(hssi_10g_tx_pcs_sop_mark),
				.stretch_num_stages(hssi_10g_tx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_tx_pcs_sup_mode),
				.test_mode(hssi_10g_tx_pcs_test_mode),
				.tx_scrm_err(hssi_10g_tx_pcs_tx_scrm_err),
				.tx_scrm_width(hssi_10g_tx_pcs_tx_scrm_width),
				.tx_sh_location(hssi_10g_tx_pcs_tx_sh_location),
				.tx_sm_bypass(hssi_10g_tx_pcs_tx_sm_bypass),
				.tx_sm_pipeln(hssi_10g_tx_pcs_tx_sm_pipeln),
				.tx_testbus_sel(hssi_10g_tx_pcs_tx_testbus_sel),
				.txfifo_empty(hssi_10g_tx_pcs_txfifo_empty),
				.txfifo_full(hssi_10g_tx_pcs_txfifo_full),
				.txfifo_mode(hssi_10g_tx_pcs_txfifo_mode),
				.txfifo_pempty(hssi_10g_tx_pcs_txfifo_pempty),
				.txfifo_pfull(hssi_10g_tx_pcs_txfifo_pfull),
				.wr_clk_sel(hssi_10g_tx_pcs_wr_clk_sel),
				.wrfifo_clken(hssi_10g_tx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_tx_pcs_blockselect),
				.distdwn_out_dv(w_hssi_10g_tx_pcs_distdwn_out_dv),
				.distdwn_out_rden(w_hssi_10g_tx_pcs_distdwn_out_rden),
				.distdwn_out_wren(w_hssi_10g_tx_pcs_distdwn_out_wren),
				.distup_out_dv(w_hssi_10g_tx_pcs_distup_out_dv),
				.distup_out_rden(w_hssi_10g_tx_pcs_distup_out_rden),
				.distup_out_wren(w_hssi_10g_tx_pcs_distup_out_wren),
				.tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pma_if(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.tx_control_out_krfec(w_hssi_10g_tx_pcs_tx_control_out_krfec),
				.tx_data_out_krfec(w_hssi_10g_tx_pcs_tx_data_out_krfec),
				.tx_data_valid_out_krfec(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.tx_fec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_fifo_num(w_hssi_10g_tx_pcs_tx_fifo_num),
				.tx_fifo_rd_ptr(w_hssi_10g_tx_pcs_tx_fifo_rd_ptr),
				.tx_fifo_wr_clk(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.tx_fifo_wr_data(w_hssi_10g_tx_pcs_tx_fifo_wr_data),
				.tx_fifo_wr_data_dw(w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw),
				.tx_fifo_wr_en(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.tx_fifo_wr_ptr(w_hssi_10g_tx_pcs_tx_fifo_wr_ptr),
				.tx_fifo_wr_rst_n(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.tx_full(w_hssi_10g_tx_pcs_tx_full),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				.tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.tx_pma_data(w_hssi_10g_tx_pcs_tx_pma_data),
				.tx_pma_gating_val(w_hssi_10g_tx_pcs_tx_pma_gating_val),
				.tx_test_data(w_hssi_10g_tx_pcs_tx_test_data),
				.tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.distdwn_in_dv(in_bond_pcs10g_in_bot[2]),
				.distdwn_in_rden(in_bond_pcs10g_in_bot[4]),
				.distdwn_in_wren(in_bond_pcs10g_in_bot[3]),
				.distup_in_dv(in_bond_pcs10g_in_top[2]),
				.distup_in_rden(in_bond_pcs10g_in_top[4]),
				.distup_in_wren(in_bond_pcs10g_in_top[3]),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_tx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_tx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.tx_bitslip({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0]}),
				.tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.tx_control({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0]}),
				.tx_control_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0]}),
				.tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0]}),
				.tx_data_in_krfec({w_hssi_krfec_tx_pcs_tx_data_out[63], w_hssi_krfec_tx_pcs_tx_data_out[62], w_hssi_krfec_tx_pcs_tx_data_out[61], w_hssi_krfec_tx_pcs_tx_data_out[60], w_hssi_krfec_tx_pcs_tx_data_out[59], w_hssi_krfec_tx_pcs_tx_data_out[58], w_hssi_krfec_tx_pcs_tx_data_out[57], w_hssi_krfec_tx_pcs_tx_data_out[56], w_hssi_krfec_tx_pcs_tx_data_out[55], w_hssi_krfec_tx_pcs_tx_data_out[54], w_hssi_krfec_tx_pcs_tx_data_out[53], w_hssi_krfec_tx_pcs_tx_data_out[52], w_hssi_krfec_tx_pcs_tx_data_out[51], w_hssi_krfec_tx_pcs_tx_data_out[50], w_hssi_krfec_tx_pcs_tx_data_out[49], w_hssi_krfec_tx_pcs_tx_data_out[48], w_hssi_krfec_tx_pcs_tx_data_out[47], w_hssi_krfec_tx_pcs_tx_data_out[46], w_hssi_krfec_tx_pcs_tx_data_out[45], w_hssi_krfec_tx_pcs_tx_data_out[44], w_hssi_krfec_tx_pcs_tx_data_out[43], w_hssi_krfec_tx_pcs_tx_data_out[42], w_hssi_krfec_tx_pcs_tx_data_out[41], w_hssi_krfec_tx_pcs_tx_data_out[40], w_hssi_krfec_tx_pcs_tx_data_out[39], w_hssi_krfec_tx_pcs_tx_data_out[38], w_hssi_krfec_tx_pcs_tx_data_out[37], w_hssi_krfec_tx_pcs_tx_data_out[36], w_hssi_krfec_tx_pcs_tx_data_out[35], w_hssi_krfec_tx_pcs_tx_data_out[34], w_hssi_krfec_tx_pcs_tx_data_out[33], w_hssi_krfec_tx_pcs_tx_data_out[32], w_hssi_krfec_tx_pcs_tx_data_out[31], w_hssi_krfec_tx_pcs_tx_data_out[30], w_hssi_krfec_tx_pcs_tx_data_out[29], w_hssi_krfec_tx_pcs_tx_data_out[28], w_hssi_krfec_tx_pcs_tx_data_out[27], w_hssi_krfec_tx_pcs_tx_data_out[26], w_hssi_krfec_tx_pcs_tx_data_out[25], w_hssi_krfec_tx_pcs_tx_data_out[24], w_hssi_krfec_tx_pcs_tx_data_out[23], w_hssi_krfec_tx_pcs_tx_data_out[22], w_hssi_krfec_tx_pcs_tx_data_out[21], w_hssi_krfec_tx_pcs_tx_data_out[20], w_hssi_krfec_tx_pcs_tx_data_out[19], w_hssi_krfec_tx_pcs_tx_data_out[18], w_hssi_krfec_tx_pcs_tx_data_out[17], w_hssi_krfec_tx_pcs_tx_data_out[16], w_hssi_krfec_tx_pcs_tx_data_out[15], w_hssi_krfec_tx_pcs_tx_data_out[14], w_hssi_krfec_tx_pcs_tx_data_out[13], w_hssi_krfec_tx_pcs_tx_data_out[12], w_hssi_krfec_tx_pcs_tx_data_out[11], w_hssi_krfec_tx_pcs_tx_data_out[10], w_hssi_krfec_tx_pcs_tx_data_out[9], w_hssi_krfec_tx_pcs_tx_data_out[8], w_hssi_krfec_tx_pcs_tx_data_out[7], w_hssi_krfec_tx_pcs_tx_data_out[6], w_hssi_krfec_tx_pcs_tx_data_out[5], w_hssi_krfec_tx_pcs_tx_data_out[4], w_hssi_krfec_tx_pcs_tx_data_out[3], w_hssi_krfec_tx_pcs_tx_data_out[2], w_hssi_krfec_tx_pcs_tx_data_out[1], w_hssi_krfec_tx_pcs_tx_data_out[0]}),
				.tx_data_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0]}),
				.tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.tx_diag_status({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0]}),
				.tx_fifo_rd_data({w_hssi_fifo_tx_pcs_data_out_10g[72], w_hssi_fifo_tx_pcs_data_out_10g[71], w_hssi_fifo_tx_pcs_data_out_10g[70], w_hssi_fifo_tx_pcs_data_out_10g[69], w_hssi_fifo_tx_pcs_data_out_10g[68], w_hssi_fifo_tx_pcs_data_out_10g[67], w_hssi_fifo_tx_pcs_data_out_10g[66], w_hssi_fifo_tx_pcs_data_out_10g[65], w_hssi_fifo_tx_pcs_data_out_10g[64], w_hssi_fifo_tx_pcs_data_out_10g[63], w_hssi_fifo_tx_pcs_data_out_10g[62], w_hssi_fifo_tx_pcs_data_out_10g[61], w_hssi_fifo_tx_pcs_data_out_10g[60], w_hssi_fifo_tx_pcs_data_out_10g[59], w_hssi_fifo_tx_pcs_data_out_10g[58], w_hssi_fifo_tx_pcs_data_out_10g[57], w_hssi_fifo_tx_pcs_data_out_10g[56], w_hssi_fifo_tx_pcs_data_out_10g[55], w_hssi_fifo_tx_pcs_data_out_10g[54], w_hssi_fifo_tx_pcs_data_out_10g[53], w_hssi_fifo_tx_pcs_data_out_10g[52], w_hssi_fifo_tx_pcs_data_out_10g[51], w_hssi_fifo_tx_pcs_data_out_10g[50], w_hssi_fifo_tx_pcs_data_out_10g[49], w_hssi_fifo_tx_pcs_data_out_10g[48], w_hssi_fifo_tx_pcs_data_out_10g[47], w_hssi_fifo_tx_pcs_data_out_10g[46], w_hssi_fifo_tx_pcs_data_out_10g[45], w_hssi_fifo_tx_pcs_data_out_10g[44], w_hssi_fifo_tx_pcs_data_out_10g[43], w_hssi_fifo_tx_pcs_data_out_10g[42], w_hssi_fifo_tx_pcs_data_out_10g[41], w_hssi_fifo_tx_pcs_data_out_10g[40], w_hssi_fifo_tx_pcs_data_out_10g[39], w_hssi_fifo_tx_pcs_data_out_10g[38], w_hssi_fifo_tx_pcs_data_out_10g[37], w_hssi_fifo_tx_pcs_data_out_10g[36], w_hssi_fifo_tx_pcs_data_out_10g[35], w_hssi_fifo_tx_pcs_data_out_10g[34], w_hssi_fifo_tx_pcs_data_out_10g[33], w_hssi_fifo_tx_pcs_data_out_10g[32], w_hssi_fifo_tx_pcs_data_out_10g[31], w_hssi_fifo_tx_pcs_data_out_10g[30], w_hssi_fifo_tx_pcs_data_out_10g[29], w_hssi_fifo_tx_pcs_data_out_10g[28], w_hssi_fifo_tx_pcs_data_out_10g[27], w_hssi_fifo_tx_pcs_data_out_10g[26], w_hssi_fifo_tx_pcs_data_out_10g[25], w_hssi_fifo_tx_pcs_data_out_10g[24], w_hssi_fifo_tx_pcs_data_out_10g[23], w_hssi_fifo_tx_pcs_data_out_10g[22], w_hssi_fifo_tx_pcs_data_out_10g[21], w_hssi_fifo_tx_pcs_data_out_10g[20], w_hssi_fifo_tx_pcs_data_out_10g[19], w_hssi_fifo_tx_pcs_data_out_10g[18], w_hssi_fifo_tx_pcs_data_out_10g[17], w_hssi_fifo_tx_pcs_data_out_10g[16], w_hssi_fifo_tx_pcs_data_out_10g[15], w_hssi_fifo_tx_pcs_data_out_10g[14], w_hssi_fifo_tx_pcs_data_out_10g[13], w_hssi_fifo_tx_pcs_data_out_10g[12], w_hssi_fifo_tx_pcs_data_out_10g[11], w_hssi_fifo_tx_pcs_data_out_10g[10], w_hssi_fifo_tx_pcs_data_out_10g[9], w_hssi_fifo_tx_pcs_data_out_10g[8], w_hssi_fifo_tx_pcs_data_out_10g[7], w_hssi_fifo_tx_pcs_data_out_10g[6], w_hssi_fifo_tx_pcs_data_out_10g[5], w_hssi_fifo_tx_pcs_data_out_10g[4], w_hssi_fifo_tx_pcs_data_out_10g[3], w_hssi_fifo_tx_pcs_data_out_10g[2], w_hssi_fifo_tx_pcs_data_out_10g[1], w_hssi_fifo_tx_pcs_data_out_10g[0]}),
				.tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_10g_reg(),
				.pld_10g_krfec_tx_pld_rst_n_fifo(),
				.pld_10g_krfec_tx_pld_rst_n_reg(),
				.pld_10g_tx_bitslip_reg(),
				.pld_10g_tx_burst_en_exe_reg(),
				.pld_10g_tx_data_valid_10g_reg(),
				.pld_10g_tx_data_valid_fifo(),
				.pld_10g_tx_data_valid_reg(),
				.pld_10g_tx_diag_status_reg(),
				.pld_10g_tx_empty_reg(),
				.pld_10g_tx_fifo_num_reg(),
				.pld_10g_tx_full_fifo(),
				.pld_10g_tx_full_reg(),
				.pld_10g_tx_pempty_reg(),
				.pld_10g_tx_pfull_fifo(),
				.pld_10g_tx_wordslip_exe_reg(),
				.pld_10g_tx_wordslip_reg(),
				.pld_pcs_tx_clk_out_10g_wire(),
				.pld_tx_burst_en_reg(),
				.pld_tx_control_lo_10g_reg(),
				.pld_tx_data_10g_fifo(),
				.pld_tx_data_lo_10g_reg()
			);
		end // if generate
		else begin
				assign w_hssi_10g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_burst_en_exe = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pma_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_control_out_krfec[8:0] = 9'b0;
				assign w_hssi_10g_tx_pcs_tx_data_out_krfec[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_data_valid_out_krfec = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_dft_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_empty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fec_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_full = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_pempty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pfull = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_gating_val[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_test_data[19:0] = 20'b0;
				assign w_hssi_10g_tx_pcs_tx_wordslip_exe = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_rx_pcs
			twentynm_hssi_8g_rx_pcs #(
				.auto_error_replacement(hssi_8g_rx_pcs_auto_error_replacement),
				.auto_speed_nego(hssi_8g_rx_pcs_auto_speed_nego),
				.bit_reversal(hssi_8g_rx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_rx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_rx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_rx_pcs_bypass_pipeline_reg),
				.byte_deserializer(hssi_8g_rx_pcs_byte_deserializer),
				.cdr_ctrl_rxvalid_mask(hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask),
				.clkcmp_pattern_n(hssi_8g_rx_pcs_clkcmp_pattern_n),
				.clkcmp_pattern_p(hssi_8g_rx_pcs_clkcmp_pattern_p),
				.clock_gate_bds_dec_asn(hssi_8g_rx_pcs_clock_gate_bds_dec_asn),
				.clock_gate_cdr_eidle(hssi_8g_rx_pcs_clock_gate_cdr_eidle),
				.clock_gate_dw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk),
				.clock_gate_dw_rm_rd(hssi_8g_rx_pcs_clock_gate_dw_rm_rd),
				.clock_gate_dw_rm_wr(hssi_8g_rx_pcs_clock_gate_dw_rm_wr),
				.clock_gate_dw_wa(hssi_8g_rx_pcs_clock_gate_dw_wa),
				.clock_gate_pc_rdclk(hssi_8g_rx_pcs_clock_gate_pc_rdclk),
				.clock_gate_sw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk),
				.clock_gate_sw_rm_rd(hssi_8g_rx_pcs_clock_gate_sw_rm_rd),
				.clock_gate_sw_rm_wr(hssi_8g_rx_pcs_clock_gate_sw_rm_wr),
				.clock_gate_sw_wa(hssi_8g_rx_pcs_clock_gate_sw_wa),
				.clock_observation_in_pld_core(hssi_8g_rx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_rx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_rx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_rx_pcs_ctrl_plane_bonding_distribution),
				.eidle_entry_eios(hssi_8g_rx_pcs_eidle_entry_eios),
				.eidle_entry_iei(hssi_8g_rx_pcs_eidle_entry_iei),
				.eidle_entry_sd(hssi_8g_rx_pcs_eidle_entry_sd),
				.eightb_tenb_decoder(hssi_8g_rx_pcs_eightb_tenb_decoder),
				.err_flags_sel(hssi_8g_rx_pcs_err_flags_sel),
				.fixed_pat_det(hssi_8g_rx_pcs_fixed_pat_det),
				.fixed_pat_num(hssi_8g_rx_pcs_fixed_pat_num),
				.force_signal_detect(hssi_8g_rx_pcs_force_signal_detect),
				.gen3_clk_en(hssi_8g_rx_pcs_gen3_clk_en),
				.gen3_rx_clk_sel(hssi_8g_rx_pcs_gen3_rx_clk_sel),
				.gen3_tx_clk_sel(hssi_8g_rx_pcs_gen3_tx_clk_sel),
				.hip_mode(hssi_8g_rx_pcs_hip_mode),
				.ibm_invalid_code(hssi_8g_rx_pcs_ibm_invalid_code),
				.invalid_code_flag_only(hssi_8g_rx_pcs_invalid_code_flag_only),
				.pad_or_edb_error_replace(hssi_8g_rx_pcs_pad_or_edb_error_replace),
				.pcs_bypass(hssi_8g_rx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_rx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_rx_pcs_phase_compensation_fifo),
				.pipe_if_enable(hssi_8g_rx_pcs_pipe_if_enable),
				.pma_dw(hssi_8g_rx_pcs_pma_dw),
				.polinv_8b10b_dec(hssi_8g_rx_pcs_polinv_8b10b_dec),
				.prot_mode(hssi_8g_rx_pcs_prot_mode),
				.rate_match(hssi_8g_rx_pcs_rate_match),
				.rate_match_del_thres(hssi_8g_rx_pcs_rate_match_del_thres),
				.rate_match_empty_thres(hssi_8g_rx_pcs_rate_match_empty_thres),
				.rate_match_full_thres(hssi_8g_rx_pcs_rate_match_full_thres),
				.rate_match_ins_thres(hssi_8g_rx_pcs_rate_match_ins_thres),
				.rate_match_start_thres(hssi_8g_rx_pcs_rate_match_start_thres),
				.reconfig_settings(hssi_8g_rx_pcs_reconfig_settings),
				.rx_clk2(hssi_8g_rx_pcs_rx_clk2),
				.rx_clk_free_running(hssi_8g_rx_pcs_rx_clk_free_running),
				.rx_pcs_urst(hssi_8g_rx_pcs_rx_pcs_urst),
				.rx_rcvd_clk(hssi_8g_rx_pcs_rx_rcvd_clk),
				.rx_rd_clk(hssi_8g_rx_pcs_rx_rd_clk),
				.rx_refclk(hssi_8g_rx_pcs_rx_refclk),
				.rx_wr_clk(hssi_8g_rx_pcs_rx_wr_clk),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_rx_pcs_sup_mode),
				.symbol_swap(hssi_8g_rx_pcs_symbol_swap),
				.sync_sm_idle_eios(hssi_8g_rx_pcs_sync_sm_idle_eios),
				.test_bus_sel(hssi_8g_rx_pcs_test_bus_sel),
				.tx_rx_parallel_loopback(hssi_8g_rx_pcs_tx_rx_parallel_loopback),
				.wa_boundary_lock_ctrl(hssi_8g_rx_pcs_wa_boundary_lock_ctrl),
				.wa_clk_slip_spacing(hssi_8g_rx_pcs_wa_clk_slip_spacing),
				.wa_det_latency_sync_status_beh(hssi_8g_rx_pcs_wa_det_latency_sync_status_beh),
				.wa_disp_err_flag(hssi_8g_rx_pcs_wa_disp_err_flag),
				.wa_kchar(hssi_8g_rx_pcs_wa_kchar),
				.wa_pd(hssi_8g_rx_pcs_wa_pd),
				.wa_pd_data(hssi_8g_rx_pcs_wa_pd_data),
				.wa_pd_polarity(hssi_8g_rx_pcs_wa_pd_polarity),
				.wa_pld_controlled(hssi_8g_rx_pcs_wa_pld_controlled),
				.wa_renumber_data(hssi_8g_rx_pcs_wa_renumber_data),
				.wa_rgnumber_data(hssi_8g_rx_pcs_wa_rgnumber_data),
				.wa_rknumber_data(hssi_8g_rx_pcs_wa_rknumber_data),
				.wa_rosnumber_data(hssi_8g_rx_pcs_wa_rosnumber_data),
				.wa_rvnumber_data(hssi_8g_rx_pcs_wa_rvnumber_data),
				.wa_sync_sm_ctrl(hssi_8g_rx_pcs_wa_sync_sm_ctrl),
				.wait_cnt(hssi_8g_rx_pcs_wait_cnt)
			) inst_twentynm_hssi_8g_rx_pcs (
				// OUTPUTS
				.a1a2k1k2flag(w_hssi_8g_rx_pcs_a1a2k1k2flag),
				.avmmreaddata(w_hssi_8g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_rx_pcs_blockselect),
				.chnl_test_bus_out(w_hssi_8g_rx_pcs_chnl_test_bus_out),
				.clock_to_pld(w_hssi_8g_rx_pcs_clock_to_pld),
				.dataout(w_hssi_8g_rx_pcs_dataout),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidle_detected(w_hssi_8g_rx_pcs_eidle_detected),
				.eios_det_cdr_ctrl(w_hssi_8g_rx_pcs_eios_det_cdr_ctrl),
				.g3_rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.g3_rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.gen2ngen1(w_hssi_8g_rx_pcs_gen2ngen1),
				.parallel_rev_loopback(w_hssi_8g_rx_pcs_parallel_rev_loopback),
				.pc_fifo_empty(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.pcfifofull(w_hssi_8g_rx_pcs_pcfifofull),
				.phystatus(w_hssi_8g_rx_pcs_phystatus),
				.pipe_data(w_hssi_8g_rx_pcs_pipe_data),
				.rd_enable_out_chnl_down(w_hssi_8g_rx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_rx_pcs_rd_enable_out_chnl_up),
				.rd_ptr1_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo),
				.rd_ptr2_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo),
				.rd_ptr_rx_phfifo(w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.reset_pc_ptrs_out_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down),
				.reset_pc_ptrs_out_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up),
				.rm_fifo_empty(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.rm_fifo_full(w_hssi_8g_rx_pcs_rm_fifo_full),
				.rx_blk_start(w_hssi_8g_rx_pcs_rx_blk_start),
				.rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.rx_data_valid(w_hssi_8g_rx_pcs_rx_data_valid),
				.rx_div_sync_out_chnl_down(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down),
				.rx_div_sync_out_chnl_up(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up),
				.rx_pipe_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.rx_pipe_soft_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rx_pma_clk_gen3(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_rcvd_clk_gen3(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_rstn_sync2wrfifo_8g(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.rx_sync_hdr(w_hssi_8g_rx_pcs_rx_sync_hdr),
				.rx_we_out_chnl_down(w_hssi_8g_rx_pcs_rx_we_out_chnl_down),
				.rx_we_out_chnl_up(w_hssi_8g_rx_pcs_rx_we_out_chnl_up),
				.rxstatus(w_hssi_8g_rx_pcs_rxstatus),
				.rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.word_align_boundary(w_hssi_8g_rx_pcs_word_align_boundary),
				.wr_clk_rx_phfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_rx_phfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_rx_rmfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_rx_rmfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_data_rx_phfifo(w_hssi_8g_rx_pcs_wr_data_rx_phfifo),
				.wr_data_rx_rmfifo(w_hssi_8g_rx_pcs_wr_data_rx_rmfifo),
				.wr_en_rx_phfifo(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_rx_rmfifo(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_rx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_rx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_rx_phfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo),
				.wr_ptr_rx_rmfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo),
				.wr_rst_n_rx_phfifo(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_rx_rmfifo(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				// INPUTS
				.a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bit_reversal_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.datain({w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0]}),
				.disable_pc_fifo_byte_serdes(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4]),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.eidleinfersel({w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0]}),
				.eios_detected_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.enable_comma_detect(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.gen3_clk_sel(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.hrd_rst(1'b0),
				.inferred_rxvalid_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.pc_fifo_rd_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.pc_fifo_wrdisable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.phystatus_int(w_hssi_pipe_gen1_2_phystatus),
				.phystatus_pcs_gen3(w_hssi_pipe_gen3_phystatus),
				.pipe_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.polarity_inversion(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.rd_data1_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0]}),
				.rd_data2_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0]}),
				.rd_data_rx_phfifo({w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[3]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[3]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.reset_pc_ptrs_asn(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5]),
				.reset_pc_ptrs_in_chnl_down(in_bond_pcs8g_in_bot[12]),
				.reset_pc_ptrs_in_chnl_up(in_bond_pcs8g_in_top[12]),
				.reset_ppm_cntrs_pcs_pma(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7]),
				.rm_fifo_read_enable(1'b0),
				.rm_fifo_write_enable(1'b0),
				.rx_blk_start_pcs_gen3({w_hssi_pipe_gen3_rx_blk_start[3], w_hssi_pipe_gen3_rx_blk_start[2], w_hssi_pipe_gen3_rx_blk_start[1], w_hssi_pipe_gen3_rx_blk_start[0]}),
				.rx_data_pcs_gen3({w_hssi_pipe_gen3_rxd_8gpcs_out[63], w_hssi_pipe_gen3_rxd_8gpcs_out[62], w_hssi_pipe_gen3_rxd_8gpcs_out[61], w_hssi_pipe_gen3_rxd_8gpcs_out[60], w_hssi_pipe_gen3_rxd_8gpcs_out[59], w_hssi_pipe_gen3_rxd_8gpcs_out[58], w_hssi_pipe_gen3_rxd_8gpcs_out[57], w_hssi_pipe_gen3_rxd_8gpcs_out[56], w_hssi_pipe_gen3_rxd_8gpcs_out[55], w_hssi_pipe_gen3_rxd_8gpcs_out[54], w_hssi_pipe_gen3_rxd_8gpcs_out[53], w_hssi_pipe_gen3_rxd_8gpcs_out[52], w_hssi_pipe_gen3_rxd_8gpcs_out[51], w_hssi_pipe_gen3_rxd_8gpcs_out[50], w_hssi_pipe_gen3_rxd_8gpcs_out[49], w_hssi_pipe_gen3_rxd_8gpcs_out[48], w_hssi_pipe_gen3_rxd_8gpcs_out[47], w_hssi_pipe_gen3_rxd_8gpcs_out[46], w_hssi_pipe_gen3_rxd_8gpcs_out[45], w_hssi_pipe_gen3_rxd_8gpcs_out[44], w_hssi_pipe_gen3_rxd_8gpcs_out[43], w_hssi_pipe_gen3_rxd_8gpcs_out[42], w_hssi_pipe_gen3_rxd_8gpcs_out[41], w_hssi_pipe_gen3_rxd_8gpcs_out[40], w_hssi_pipe_gen3_rxd_8gpcs_out[39], w_hssi_pipe_gen3_rxd_8gpcs_out[38], w_hssi_pipe_gen3_rxd_8gpcs_out[37], w_hssi_pipe_gen3_rxd_8gpcs_out[36], w_hssi_pipe_gen3_rxd_8gpcs_out[35], w_hssi_pipe_gen3_rxd_8gpcs_out[34], w_hssi_pipe_gen3_rxd_8gpcs_out[33], w_hssi_pipe_gen3_rxd_8gpcs_out[32], w_hssi_pipe_gen3_rxd_8gpcs_out[31], w_hssi_pipe_gen3_rxd_8gpcs_out[30], w_hssi_pipe_gen3_rxd_8gpcs_out[29], w_hssi_pipe_gen3_rxd_8gpcs_out[28], w_hssi_pipe_gen3_rxd_8gpcs_out[27], w_hssi_pipe_gen3_rxd_8gpcs_out[26], w_hssi_pipe_gen3_rxd_8gpcs_out[25], w_hssi_pipe_gen3_rxd_8gpcs_out[24], w_hssi_pipe_gen3_rxd_8gpcs_out[23], w_hssi_pipe_gen3_rxd_8gpcs_out[22], w_hssi_pipe_gen3_rxd_8gpcs_out[21], w_hssi_pipe_gen3_rxd_8gpcs_out[20], w_hssi_pipe_gen3_rxd_8gpcs_out[19], w_hssi_pipe_gen3_rxd_8gpcs_out[18], w_hssi_pipe_gen3_rxd_8gpcs_out[17], w_hssi_pipe_gen3_rxd_8gpcs_out[16], w_hssi_pipe_gen3_rxd_8gpcs_out[15], w_hssi_pipe_gen3_rxd_8gpcs_out[14], w_hssi_pipe_gen3_rxd_8gpcs_out[13], w_hssi_pipe_gen3_rxd_8gpcs_out[12], w_hssi_pipe_gen3_rxd_8gpcs_out[11], w_hssi_pipe_gen3_rxd_8gpcs_out[10], w_hssi_pipe_gen3_rxd_8gpcs_out[9], w_hssi_pipe_gen3_rxd_8gpcs_out[8], w_hssi_pipe_gen3_rxd_8gpcs_out[7], w_hssi_pipe_gen3_rxd_8gpcs_out[6], w_hssi_pipe_gen3_rxd_8gpcs_out[5], w_hssi_pipe_gen3_rxd_8gpcs_out[4], w_hssi_pipe_gen3_rxd_8gpcs_out[3], w_hssi_pipe_gen3_rxd_8gpcs_out[2], w_hssi_pipe_gen3_rxd_8gpcs_out[1], w_hssi_pipe_gen3_rxd_8gpcs_out[0]}),
				.rx_data_valid_pcs_gen3({w_hssi_pipe_gen3_rxdataskip[3], w_hssi_pipe_gen3_rxdataskip[2], w_hssi_pipe_gen3_rxdataskip[1], w_hssi_pipe_gen3_rxdataskip[0]}),
				.rx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[1], in_bond_pcs8g_in_bot[0]}),
				.rx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[1], in_bond_pcs8g_in_top[0]}),
				.rx_pcs_rst(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.rx_sync_hdr_pcs_gen3({w_hssi_pipe_gen3_rx_sync_hdr[1], w_hssi_pipe_gen3_rx_sync_hdr[0]}),
				.rx_we_in_chnl_down({in_bond_pcs8g_in_bot[5], in_bond_pcs8g_in_bot[4]}),
				.rx_we_in_chnl_up({in_bond_pcs8g_in_top[5], in_bond_pcs8g_in_top[4]}),
				.rxstatus_int({w_hssi_pipe_gen1_2_rxstatus[2], w_hssi_pipe_gen1_2_rxstatus[1], w_hssi_pipe_gen1_2_rxstatus[0]}),
				.rxstatus_pcs_gen3({w_hssi_pipe_gen3_rxstatus[2], w_hssi_pipe_gen3_rxstatus[1], w_hssi_pipe_gen3_rxstatus[0]}),
				.rxvalid_int(w_hssi_pipe_gen1_2_rxvalid),
				.rxvalid_pcs_gen3(w_hssi_pipe_gen3_rxvalid),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.sig_det_from_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_ctrlplane_testbus({w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0]}),
				.tx_div_sync({w_hssi_8g_tx_pcs_tx_div_sync[1], w_hssi_8g_tx_pcs_tx_div_sync[0]}),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.tx_testbus({w_hssi_8g_tx_pcs_tx_testbus[19], w_hssi_8g_tx_pcs_tx_testbus[18], w_hssi_8g_tx_pcs_tx_testbus[17], w_hssi_8g_tx_pcs_tx_testbus[16], w_hssi_8g_tx_pcs_tx_testbus[15], w_hssi_8g_tx_pcs_tx_testbus[14], w_hssi_8g_tx_pcs_tx_testbus[13], w_hssi_8g_tx_pcs_tx_testbus[12], w_hssi_8g_tx_pcs_tx_testbus[11], w_hssi_8g_tx_pcs_tx_testbus[10], w_hssi_8g_tx_pcs_tx_testbus[9], w_hssi_8g_tx_pcs_tx_testbus[8], w_hssi_8g_tx_pcs_tx_testbus[7], w_hssi_8g_tx_pcs_tx_testbus[6], w_hssi_8g_tx_pcs_tx_testbus[5], w_hssi_8g_tx_pcs_tx_testbus[4], w_hssi_8g_tx_pcs_tx_testbus[3], w_hssi_8g_tx_pcs_tx_testbus[2], w_hssi_8g_tx_pcs_tx_testbus[1], w_hssi_8g_tx_pcs_tx_testbus[0]}),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[2]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[2]),
				
				// UNUSED
				.byte_deserializer_pcs_clk_div_by_2_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_wire(),
				.byte_deserializer_pcs_clk_div_by_2_wire(),
				.byte_deserializer_pcs_clk_div_by_4_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_2_reg(),
				.byte_deserializer_pld_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_4_txclk_reg(),
				.pld_8g_a1a2_k1k2_flag_reg(),
				.pld_8g_a1a2_k1k2_flag_txclk_reg(),
				.pld_8g_a1a2_size_reg(),
				.pld_8g_a1a2_size_txclk_reg(),
				.pld_8g_bitloc_rev_en_reg(),
				.pld_8g_bitloc_rev_en_txclk_reg(),
				.pld_8g_byte_rev_en_reg(),
				.pld_8g_byte_rev_en_txclk_reg(),
				.pld_8g_elecidle_reg(),
				.pld_8g_empty_rmf_lowlatency_reg(),
				.pld_8g_empty_rmf_lowlatency_txclk_reg(),
				.pld_8g_empty_rmf_reg(),
				.pld_8g_empty_rmf_txclk_reg(),
				.pld_8g_empty_rx_fifo(),
				.pld_8g_empty_rx_reg(),
				.pld_8g_empty_rx_txclk_reg(),
				.pld_8g_encdt_reg(),
				.pld_8g_encdt_txclk_reg(),
				.pld_8g_full_rmf_reg(),
				.pld_8g_full_rmf_txclk_reg(),
				.pld_8g_full_rx_fifo(),
				.pld_8g_full_rx_reg(),
				.pld_8g_full_rx_txclk_reg(),
				.pld_8g_g3_rx_pld_rst_n_reg(),
				.pld_8g_g3_rx_pld_rst_n_txclk_reg(),
				.pld_8g_rxelecidle_txclk_reg(),
				.pld_8g_rxpolarity_reg(),
				.pld_8g_rxpolarity_txclk_reg(),
				.pld_8g_wa_boundary_reg(),
				.pld_8g_wrdisable_rx_reg(),
				.pld_8g_wrdisable_rx_txclk_reg(),
				.pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_rx_clk_out_8g_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_wire(),
				.pld_rx_control_8g_reg(),
				.pld_rx_control_8g_txclk_reg(),
				.pld_rx_data_8g_reg(),
				.pld_rx_data_8g_txclk_reg(),
				.pld_syncsm_en_reg(),
				.pld_syncsm_en_txclk_reg(),
				.rm_fifo_partial_empty(),
				.rm_fifo_partial_full(),
				.sta_rx_clk2_by2_1(),
				.sta_rx_clk2_by2_1_out(),
				.sta_rx_clk2_by2_2(),
				.sta_rx_clk2_by2_2_out(),
				.sta_rx_clk2_by4_1(),
				.sta_rx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_rx_pcs_a1a2k1k2flag[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_rx_pcs_chnl_test_bus_out[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_clock_to_pld = 1'b0;
				assign w_hssi_8g_rx_pcs_dataout[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_dis_pc_byte = 1'b0;
				assign w_hssi_8g_rx_pcs_eidle_detected = 1'b0;
				assign w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_pma_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_gen2ngen1 = 1'b0;
				assign w_hssi_8g_rx_pcs_parallel_rev_loopback[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_pc_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_pcfifofull = 1'b0;
				assign w_hssi_8g_rx_pcs_phystatus = 1'b0;
				assign w_hssi_8g_rx_pcs_pipe_data[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_full = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clkslip = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_data_valid[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pma_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rxstatus[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_rxvalid = 1'b0;
				assign w_hssi_8g_rx_pcs_signal_detect_out = 1'b0;
				assign w_hssi_8g_rx_pcs_word_align_boundary[4:0] = 5'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79:0] = 80'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31:0] = 32'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_rmfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_tx_pcs
			twentynm_hssi_8g_tx_pcs #(
				.auto_speed_nego_gen2(hssi_8g_tx_pcs_auto_speed_nego_gen2),
				.bit_reversal(hssi_8g_tx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_tx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_tx_pcs_bypass_pipeline_reg),
				.byte_serializer(hssi_8g_tx_pcs_byte_serializer),
				.clock_gate_bs_enc(hssi_8g_tx_pcs_clock_gate_bs_enc),
				.clock_gate_dw_fifowr(hssi_8g_tx_pcs_clock_gate_dw_fifowr),
				.clock_gate_fiford(hssi_8g_tx_pcs_clock_gate_fiford),
				.clock_gate_sw_fifowr(hssi_8g_tx_pcs_clock_gate_sw_fifowr),
				.clock_observation_in_pld_core(hssi_8g_tx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_tx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_tx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_tx_pcs_ctrl_plane_bonding_distribution),
				.data_selection_8b10b_encoder_input(hssi_8g_tx_pcs_data_selection_8b10b_encoder_input),
				.dynamic_clk_switch(hssi_8g_tx_pcs_dynamic_clk_switch),
				.eightb_tenb_disp_ctrl(hssi_8g_tx_pcs_eightb_tenb_disp_ctrl),
				.eightb_tenb_encoder(hssi_8g_tx_pcs_eightb_tenb_encoder),
				.force_echar(hssi_8g_tx_pcs_force_echar),
				.force_kchar(hssi_8g_tx_pcs_force_kchar),
				.gen3_tx_clk_sel(hssi_8g_tx_pcs_gen3_tx_clk_sel),
				.gen3_tx_pipe_clk_sel(hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel),
				.hip_mode(hssi_8g_tx_pcs_hip_mode),
				.pcs_bypass(hssi_8g_tx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_tx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_tx_pcs_phase_compensation_fifo),
				.phfifo_write_clk_sel(hssi_8g_tx_pcs_phfifo_write_clk_sel),
				.pma_dw(hssi_8g_tx_pcs_pma_dw),
				.prot_mode(hssi_8g_tx_pcs_prot_mode),
				.reconfig_settings(hssi_8g_tx_pcs_reconfig_settings),
				.refclk_b_clk_sel(hssi_8g_tx_pcs_refclk_b_clk_sel),
				.revloop_back_rm(hssi_8g_tx_pcs_revloop_back_rm),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_tx_pcs_sup_mode),
				.symbol_swap(hssi_8g_tx_pcs_symbol_swap),
				.tx_bitslip(hssi_8g_tx_pcs_tx_bitslip),
				.tx_compliance_controlled_disparity(hssi_8g_tx_pcs_tx_compliance_controlled_disparity),
				.tx_fast_pld_reg(hssi_8g_tx_pcs_tx_fast_pld_reg),
				.txclk_freerun(hssi_8g_tx_pcs_txclk_freerun),
				.txpcs_urst(hssi_8g_tx_pcs_txpcs_urst)
			) inst_twentynm_hssi_8g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_8g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_tx_pcs_blockselect),
				.clk_out(w_hssi_8g_tx_pcs_clk_out),
				.clk_out_gen3(w_hssi_8g_tx_pcs_clk_out_gen3),
				.dataout(w_hssi_8g_tx_pcs_dataout),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.fifo_select_out_chnl_down(w_hssi_8g_tx_pcs_fifo_select_out_chnl_down),
				.fifo_select_out_chnl_up(w_hssi_8g_tx_pcs_fifo_select_out_chnl_up),
				.g3_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.g3_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
				.non_gray_eidleinfersel(w_hssi_8g_tx_pcs_non_gray_eidleinfersel),
				.ph_fifo_overflow(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.ph_fifo_underflow(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.phfifo_txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.phfifo_txmargin(w_hssi_8g_tx_pcs_phfifo_txmargin),
				.phfifo_txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				.pipe_en_rev_parallel_lpbk_out(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.pipe_power_down_out(w_hssi_8g_tx_pcs_pipe_power_down_out),
				.pipe_tx_clk_out_gen3(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pmaif_asn_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.rd_enable_out_chnl_down(w_hssi_8g_tx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_tx_pcs_rd_enable_out_chnl_up),
				.rd_ptr_tx_phfifo(w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rxpolarity_int(w_hssi_8g_tx_pcs_rxpolarity_int),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.tx_blk_start_out(w_hssi_8g_tx_pcs_tx_blk_start_out),
				.tx_clk_out_8g_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.tx_ctrlplane_testbus(w_hssi_8g_tx_pcs_tx_ctrlplane_testbus),
				.tx_data_out(w_hssi_8g_tx_pcs_tx_data_out),
				.tx_data_valid_out(w_hssi_8g_tx_pcs_tx_data_valid_out),
				.tx_datak_out(w_hssi_8g_tx_pcs_tx_datak_out),
				.tx_detect_rxloopback_int(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.tx_div_sync(w_hssi_8g_tx_pcs_tx_div_sync),
				.tx_div_sync_out_chnl_down(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down),
				.tx_div_sync_out_chnl_up(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up),
				.tx_pipe_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.tx_pipe_electidle(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_soft_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.tx_sync_hdr_out(w_hssi_8g_tx_pcs_tx_sync_hdr_out),
				.tx_testbus(w_hssi_8g_tx_pcs_tx_testbus),
				.txcompliance_out(w_hssi_8g_tx_pcs_txcompliance_out),
				.txelecidle_out(w_hssi_8g_tx_pcs_txelecidle_out),
				.wr_clk_tx_phfifo_dw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_tx_phfifo_sw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_data_tx_phfifo(w_hssi_8g_tx_pcs_wr_data_tx_phfifo),
				.wr_en_tx_phfifo(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_tx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_tx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_tx_phfifo(w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo),
				.wr_rst_n_tx_phfifo(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bitslip_boundary_select({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0]}),
				.clk_sel_gen3(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.coreclk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.datain({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.detectrxloopin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidleinfersel({w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0]}),
				.en_rev_parallel_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.fifo_select_in_chnl_down({in_bond_pcs8g_in_bot[11], in_bond_pcs8g_in_bot[10]}),
				.fifo_select_in_chnl_up({in_bond_pcs8g_in_top[11], in_bond_pcs8g_in_top[10]}),
				.hrdrst(1'b0),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.ph_fifo_rd_disable(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.pipe_en_rev_parallel_lpbk_in(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.pipe_tx_deemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.pipe_tx_margin({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0]}),
				.powerdn({w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0]}),
				.rate_switch(w_hssi_8g_rx_pcs_gen2ngen1),
				.rd_data_tx_phfifo({w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[9]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[9]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.rev_parallel_lpbk_data({w_hssi_8g_rx_pcs_parallel_rev_loopback[19], w_hssi_8g_rx_pcs_parallel_rev_loopback[18], w_hssi_8g_rx_pcs_parallel_rev_loopback[17], w_hssi_8g_rx_pcs_parallel_rev_loopback[16], w_hssi_8g_rx_pcs_parallel_rev_loopback[15], w_hssi_8g_rx_pcs_parallel_rev_loopback[14], w_hssi_8g_rx_pcs_parallel_rev_loopback[13], w_hssi_8g_rx_pcs_parallel_rev_loopback[12], w_hssi_8g_rx_pcs_parallel_rev_loopback[11], w_hssi_8g_rx_pcs_parallel_rev_loopback[10], w_hssi_8g_rx_pcs_parallel_rev_loopback[9], w_hssi_8g_rx_pcs_parallel_rev_loopback[8], w_hssi_8g_rx_pcs_parallel_rev_loopback[7], w_hssi_8g_rx_pcs_parallel_rev_loopback[6], w_hssi_8g_rx_pcs_parallel_rev_loopback[5], w_hssi_8g_rx_pcs_parallel_rev_loopback[4], w_hssi_8g_rx_pcs_parallel_rev_loopback[3], w_hssi_8g_rx_pcs_parallel_rev_loopback[2], w_hssi_8g_rx_pcs_parallel_rev_loopback[1], w_hssi_8g_rx_pcs_parallel_rev_loopback[0]}),
				.rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.tx_blk_start({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0]}),
				.tx_data_valid({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0]}),
				.tx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[7], in_bond_pcs8g_in_bot[6]}),
				.tx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[7], in_bond_pcs8g_in_top[6]}),
				.tx_pcs_reset(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.tx_sync_hdr({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0]}),
				.txd_fast_reg({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0]}),
				.txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[8]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[8]),
				.wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				
				// UNUSED
				.byte_serializer_pcs_clk_div_by_2_reg(),
				.byte_serializer_pcs_clk_div_by_2_wire(),
				.byte_serializer_pcs_clk_div_by_4_reg(),
				.byte_serializer_pld_clk_div_by_2_reg(),
				.byte_serializer_pld_clk_div_by_4_reg(),
				.pld_8g_empty_tx_fifo(),
				.pld_8g_empty_tx_reg(),
				.pld_8g_full_tx_fifo(),
				.pld_8g_full_tx_reg(),
				.pld_8g_g3_tx_pld_rst_n_reg(),
				.pld_8g_rddisable_tx_reg(),
				.pld_8g_tx_boundary_sel_reg(),
				.pld_pcs_tx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_tx_clk_out_8g_wire(),
				.pld_tx_data_8g_fifo(),
				.pld_tx_data_lo_8g_reg(),
				.sta_tx_clk2_by2_1(),
				.sta_tx_clk2_by2_1_out(),
				.sta_tx_clk2_by4_1(),
				.sta_tx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_dataout[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_dyn_clk_switch_n = 1'b1;		// Override default tieoff
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_g3_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_overflow = 1'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_underflow = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txdeemph = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txmargin[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txswing = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_power_down_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_pmaif_asn_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_refclk_b = 1'b0;
				assign w_hssi_8g_tx_pcs_refclk_b_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_rxpolarity_int = 1'b0;
				assign w_hssi_8g_tx_pcs_soft_reset_wclk1_n = 1'b0;
				assign w_hssi_8g_tx_pcs_sw_fifo_wr_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_blk_start_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_tx_data_out[31:0] = 32'b0;
				assign w_hssi_8g_tx_pcs_tx_data_valid_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_datak_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_detect_rxloopback_int = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_electidle = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_sync_hdr_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_txcompliance_out = 1'b0;
				assign w_hssi_8g_tx_pcs_txelecidle_out = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63:0] = 64'b0;
				assign w_hssi_8g_tx_pcs_wr_en_tx_phfifo = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pcs_pma_interface
			twentynm_hssi_common_pcs_pma_interface #(
				.asn_clk_enable(hssi_common_pcs_pma_interface_asn_clk_enable),
				.asn_enable(hssi_common_pcs_pma_interface_asn_enable),
				.block_sel(hssi_common_pcs_pma_interface_block_sel),
				.bypass_early_eios(hssi_common_pcs_pma_interface_bypass_early_eios),
				.bypass_pcie_switch(hssi_common_pcs_pma_interface_bypass_pcie_switch),
				.bypass_pma_ltr(hssi_common_pcs_pma_interface_bypass_pma_ltr),
				.bypass_pma_sw_done(hssi_common_pcs_pma_interface_bypass_pma_sw_done),
				.bypass_ppm_lock(hssi_common_pcs_pma_interface_bypass_ppm_lock),
				.bypass_send_syncp_fbkp(hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp),
				.bypass_txdetectrx(hssi_common_pcs_pma_interface_bypass_txdetectrx),
				.cdr_control(hssi_common_pcs_pma_interface_cdr_control),
				.cid_enable(hssi_common_pcs_pma_interface_cid_enable),
				.cp_cons_sel(hssi_common_pcs_pma_interface_cp_cons_sel),
				.cp_dwn_mstr(hssi_common_pcs_pma_interface_cp_dwn_mstr),
				.cp_up_mstr(hssi_common_pcs_pma_interface_cp_up_mstr),
				.ctrl_plane_bonding(hssi_common_pcs_pma_interface_ctrl_plane_bonding),
				.data_mask_count(hssi_common_pcs_pma_interface_data_mask_count),
				.data_mask_count_multi(hssi_common_pcs_pma_interface_data_mask_count_multi),
				.dft_observation_clock_selection(hssi_common_pcs_pma_interface_dft_observation_clock_selection),
				.early_eios_counter(hssi_common_pcs_pma_interface_early_eios_counter),
				.force_freqdet(hssi_common_pcs_pma_interface_force_freqdet),
				.free_run_clk_enable(hssi_common_pcs_pma_interface_free_run_clk_enable),
				.ignore_sigdet_g23(hssi_common_pcs_pma_interface_ignore_sigdet_g23),
				.pc_en_counter(hssi_common_pcs_pma_interface_pc_en_counter),
				.pc_rst_counter(hssi_common_pcs_pma_interface_pc_rst_counter),
				.pcie_hip_mode(hssi_common_pcs_pma_interface_pcie_hip_mode),
				.ph_fifo_reg_mode(hssi_common_pcs_pma_interface_ph_fifo_reg_mode),
				.phfifo_flush_wait(hssi_common_pcs_pma_interface_phfifo_flush_wait),
				.pipe_if_g3pcs(hssi_common_pcs_pma_interface_pipe_if_g3pcs),
				.pma_done_counter(hssi_common_pcs_pma_interface_pma_done_counter),
				.pma_if_dft_en(hssi_common_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_common_pcs_pma_interface_pma_if_dft_val),
				.ppm_cnt_rst(hssi_common_pcs_pma_interface_ppm_cnt_rst),
				.ppm_deassert_early(hssi_common_pcs_pma_interface_ppm_deassert_early),
				.ppm_det_buckets(hssi_common_pcs_pma_interface_ppm_det_buckets),
				.ppm_gen1_2_cnt(hssi_common_pcs_pma_interface_ppm_gen1_2_cnt),
				.ppm_post_eidle_delay(hssi_common_pcs_pma_interface_ppm_post_eidle_delay),
				.ppmsel(hssi_common_pcs_pma_interface_ppmsel),
				.prot_mode(hssi_common_pcs_pma_interface_prot_mode),
				.reconfig_settings(hssi_common_pcs_pma_interface_reconfig_settings),
				.rxvalid_mask(hssi_common_pcs_pma_interface_rxvalid_mask),
				.sigdet_wait_counter(hssi_common_pcs_pma_interface_sigdet_wait_counter),
				.sigdet_wait_counter_multi(hssi_common_pcs_pma_interface_sigdet_wait_counter_multi),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sim_mode(hssi_common_pcs_pma_interface_sim_mode),
				.spd_chg_rst_wait_cnt_en(hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en),
				.sup_mode(hssi_common_pcs_pma_interface_sup_mode),
				.testout_sel(hssi_common_pcs_pma_interface_testout_sel),
				.wait_clk_on_off_timer(hssi_common_pcs_pma_interface_wait_clk_on_off_timer),
				.wait_pipe_synchronizing(hssi_common_pcs_pma_interface_wait_pipe_synchronizing),
				.wait_send_syncp_fbkp(hssi_common_pcs_pma_interface_wait_send_syncp_fbkp)
			) inst_twentynm_hssi_common_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_common_pcs_pma_interface_blockselect),
				.int_pmaif_8g_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in),
				.int_pmaif_8g_eios_detected(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.int_pmaif_8g_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.int_pmaif_8g_power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.int_pmaif_g3_pcs_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in),
				.int_pmaif_pldif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pmaif_pldif_pcie_sw_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done),
				.int_pmaif_pldif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pmaif_pldif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pmaif_pldif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pmaif_pldif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pmaif_pldif_pma_reserved_in(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in),
				.int_pmaif_pldif_test_out(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out),
				.int_pmaif_pldif_testbus(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus),
				.pma_adapt_start(w_hssi_common_pcs_pma_interface_pma_adapt_start),
				.pma_atpg_los_en_n(w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n),
				.pma_csr_test_dis(w_hssi_common_pcs_pma_interface_pma_csr_test_dis),
				.pma_current_coeff(w_hssi_common_pcs_pma_interface_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_common_pcs_pma_interface_pma_current_rxpreset),
				.pma_early_eios(w_hssi_common_pcs_pma_interface_pma_early_eios),
				.pma_interface_select(w_hssi_common_pcs_pma_interface_pma_interface_select),
				.pma_ltd_b(w_hssi_common_pcs_pma_interface_pma_ltd_b),
				.pma_ltr(w_hssi_common_pcs_pma_interface_pma_ltr),
				.pma_nfrzdrv(w_hssi_common_pcs_pma_interface_pma_nfrzdrv),
				.pma_nrpi_freeze(w_hssi_common_pcs_pma_interface_pma_nrpi_freeze),
				.pma_pcie_switch(w_hssi_common_pcs_pma_interface_pma_pcie_switch),
				.pma_ppm_lock(w_hssi_common_pcs_pma_interface_pma_ppm_lock),
				.pma_reserved_out(w_hssi_common_pcs_pma_interface_pma_reserved_out),
				.pma_rs_lpbk_b(w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b),
				.pma_rx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup),
				.pma_scan_mode_n(w_hssi_common_pcs_pma_interface_pma_scan_mode_n),
				.pma_scan_shift_n(w_hssi_common_pcs_pma_interface_pma_scan_shift_n),
				.pma_tx_bitslip(w_hssi_common_pcs_pma_interface_pma_tx_bitslip),
				.pma_tx_bonding_rstb(w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb),
				.pma_tx_qpi_pulldn(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn),
				.pma_tx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup),
				.pma_tx_txdetectrx(w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx),
				.pmaif_bundling_out_down(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down),
				.pmaif_bundling_out_up(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_8g_current_coeff({w_hssi_pipe_gen1_2_current_coeff[17], w_hssi_pipe_gen1_2_current_coeff[16], w_hssi_pipe_gen1_2_current_coeff[15], w_hssi_pipe_gen1_2_current_coeff[14], w_hssi_pipe_gen1_2_current_coeff[13], w_hssi_pipe_gen1_2_current_coeff[12], w_hssi_pipe_gen1_2_current_coeff[11], w_hssi_pipe_gen1_2_current_coeff[10], w_hssi_pipe_gen1_2_current_coeff[9], w_hssi_pipe_gen1_2_current_coeff[8], w_hssi_pipe_gen1_2_current_coeff[7], w_hssi_pipe_gen1_2_current_coeff[6], w_hssi_pipe_gen1_2_current_coeff[5], w_hssi_pipe_gen1_2_current_coeff[4], w_hssi_pipe_gen1_2_current_coeff[3], w_hssi_pipe_gen1_2_current_coeff[2], w_hssi_pipe_gen1_2_current_coeff[1], w_hssi_pipe_gen1_2_current_coeff[0]}),
				.int_pmaif_8g_eios_det({w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0]}),
				.int_pmaif_8g_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.int_pmaif_8g_rev_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.int_pmaif_8g_tx_clk_out_gen3(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.int_pmaif_8g_txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				.int_pmaif_g3_eios_det({w_hssi_gen3_rx_pcs_ei_det_int, w_hssi_gen3_rx_pcs_ei_partial_det_int, w_hssi_gen3_rx_pcs_i_det_int}),
				.int_pmaif_g3_pma_current_coeff({w_hssi_pipe_gen3_pma_current_coeff[17], w_hssi_pipe_gen3_pma_current_coeff[16], w_hssi_pipe_gen3_pma_current_coeff[15], w_hssi_pipe_gen3_pma_current_coeff[14], w_hssi_pipe_gen3_pma_current_coeff[13], w_hssi_pipe_gen3_pma_current_coeff[12], w_hssi_pipe_gen3_pma_current_coeff[11], w_hssi_pipe_gen3_pma_current_coeff[10], w_hssi_pipe_gen3_pma_current_coeff[9], w_hssi_pipe_gen3_pma_current_coeff[8], w_hssi_pipe_gen3_pma_current_coeff[7], w_hssi_pipe_gen3_pma_current_coeff[6], w_hssi_pipe_gen3_pma_current_coeff[5], w_hssi_pipe_gen3_pma_current_coeff[4], w_hssi_pipe_gen3_pma_current_coeff[3], w_hssi_pipe_gen3_pma_current_coeff[2], w_hssi_pipe_gen3_pma_current_coeff[1], w_hssi_pipe_gen3_pma_current_coeff[0]}),
				.int_pmaif_g3_pma_current_rxpreset({w_hssi_pipe_gen3_pma_current_rxpreset[2], w_hssi_pipe_gen3_pma_current_rxpreset[1], w_hssi_pipe_gen3_pma_current_rxpreset[0]}),
				.int_pmaif_g3_pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.int_pmaif_g3_rev_lpbk(w_hssi_pipe_gen3_rev_lpbk_int),
				.int_pmaif_pldif_8g_tx_pld_rstn(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pmaif_pldif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pmaif_pldif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pmaif_pldif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pmaif_pldif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pmaif_pldif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pmaif_pldif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pmaif_pldif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pmaif_pldif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pmaif_pldif_pcie_switch({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0]}),
				.int_pmaif_pldif_pma_reserved_out({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0]}),
				.int_pmaif_pldif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pmaif_pldif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pmaif_pldif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pmaif_pldif_rate({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0]}),
				.int_pmaif_pldif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pmaif_pldif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pmaif_pldif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.int_pmaif_pldif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pmaif_pldif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pmaif_pldif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pmaif_pldif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pmaif_pldif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pmaif_pldif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.int_tx_dft_obsrv_clk({w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0]}),
				.iocsr_clk(in_iocsr_clk),
				.iocsr_config({in_iocsr_config[5], in_iocsr_config[4], in_iocsr_config[3], in_iocsr_config[2], in_iocsr_config[1], in_iocsr_config[0]}),
				.iocsr_rdy(in_iocsr_rdy),
				.iocsr_rdy_dly(in_iocsr_rdy_dly),
				.pma_adapt_done(in_pma_adapt_done),
				.pma_clklow(in_pma_clklow),
				.pma_fref(in_pma_fref),
				.pma_hclk(in_pma_hclk),
				.pma_pcie_sw_done({in_pma_pcie_sw_done[1], in_pma_pcie_sw_done[0]}),
				.pma_pfdmode_lock(in_pma_pfdmode_lock),
				.pma_reserved_in({in_pma_reserved_in[4], in_pma_reserved_in[3], in_pma_reserved_in[2], in_pma_reserved_in[1], in_pma_reserved_in[0]}),
				.pma_signal_det(in_pma_signal_det),
				.pma_testbus({in_pma_testbus[7], in_pma_testbus[6], in_pma_testbus[5], in_pma_testbus[4], in_pma_testbus[3], in_pma_testbus[2], in_pma_testbus[1], in_pma_testbus[0]}),
				.pmaif_bundling_in_down({in_bond_pmaif_in_bot[11], in_bond_pmaif_in_bot[10], in_bond_pmaif_in_bot[9], in_bond_pmaif_in_bot[8], in_bond_pmaif_in_bot[7], in_bond_pmaif_in_bot[6], in_bond_pmaif_in_bot[5], in_bond_pmaif_in_bot[4], in_bond_pmaif_in_bot[3], in_bond_pmaif_in_bot[2], in_bond_pmaif_in_bot[1], in_bond_pmaif_in_bot[0]}),
				.pmaif_bundling_in_up({in_bond_pmaif_in_top[11], in_bond_pmaif_in_top[10], in_bond_pmaif_in_top[9], in_bond_pmaif_in_top[8], in_bond_pmaif_in_top[7], in_bond_pmaif_in_top[6], in_bond_pmaif_in_top[5], in_bond_pmaif_in_top[4], in_bond_pmaif_in_top[3], in_bond_pmaif_in_top[2], in_bond_pmaif_in_top[1], in_bond_pmaif_in_top[0]}),
				.rx_pmaif_test_out({w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0]}),
				.rx_prbs_ver_test({w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0]}),
				.tx_prbs_gen_test({w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0]}),
				.uhsif_test_out_1({w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0]}),
				.uhsif_test_out_2({w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0]}),
				.uhsif_test_out_3({w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0]}),
				
				// UNUSED
				.int_pmaif_avmm_iocsr_clk(),
				.int_pmaif_avmm_iocsr_config(),
				.int_pmaif_avmm_iocsr_rdy(),
				.int_pmaif_avmm_iocsr_rdy_dly(),
				.int_pmaif_pldif_interface_select(),
				.pma_tx_pma_syncp(),
				.sta_pma_hclk_by2()
			);
		end // if generate
		else begin
				assign w_hssi_common_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19:0] = 20'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_pma_adapt_start = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_csr_test_dis = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pcs_pma_interface_pma_early_eios = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_interface_select[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltd_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltr = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nfrzdrv = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nrpi_freeze = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ppm_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_tx_bitslip = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx = in_pld_pma_txdetectrx;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11:0] = 12'b0;
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11:0] = 12'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pld_pcs_interface
			twentynm_hssi_common_pld_pcs_interface #(
				.dft_clk_out_en(hssi_common_pld_pcs_interface_dft_clk_out_en),
				.dft_clk_out_sel(hssi_common_pld_pcs_interface_dft_clk_out_sel),
				.hrdrstctrl_en(hssi_common_pld_pcs_interface_hrdrstctrl_en),
				.pcs_testbus_block_sel(hssi_common_pld_pcs_interface_pcs_testbus_block_sel),
				.reconfig_settings(hssi_common_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm5es2" )       //PARAM_HIDE
			) inst_twentynm_hssi_common_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_common_pld_pcs_interface_blockselect),
				.hip_cmn_clk(w_hssi_common_pld_pcs_interface_hip_cmn_clk),
				.hip_cmn_ctrl(w_hssi_common_pld_pcs_interface_hip_cmn_ctrl),
				.hip_iocsr_rdy(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy),
				.hip_iocsr_rdy_dly(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly),
				.hip_nfrzdrv(w_hssi_common_pld_pcs_interface_hip_nfrzdrv),
				.hip_npor(w_hssi_common_pld_pcs_interface_hip_npor),
				.hip_usermode(w_hssi_common_pld_pcs_interface_hip_usermode),
				.int_pldif_10g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.int_pldif_10g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.int_pldif_8g_eidleinfersel(w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel),
				.int_pldif_8g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.int_pldif_8g_refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.int_pldif_8g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.int_pldif_g3_current_coeff(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff),
				.int_pldif_g3_current_rxpreset(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset),
				.int_pldif_krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.int_pldif_krfec_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.int_pldif_krfec_scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				.int_pldif_mem_atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.int_pldif_mem_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.int_pldif_pmaif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pldif_pmaif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pldif_pmaif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pldif_pmaif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pldif_pmaif_eye_monitor(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor),
				.int_pldif_pmaif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pldif_pmaif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pldif_pmaif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pldif_pmaif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pldif_pmaif_pcie_switch(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch),
				.int_pldif_pmaif_pma_reserved_out(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out),
				.int_pldif_pmaif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pldif_pmaif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pldif_pmaif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pldif_pmaif_rate(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate),
				.int_pldif_pmaif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pldif_pmaif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pldif_pmaif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pldif_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_pldif_pmaif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pldif_pmaif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pldif_pmaif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pldif_pmaif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pldif_pmaif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pldif_pmaif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pldif_pmaif_uhsif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.pld_pma_adapt_done(w_hssi_common_pld_pcs_interface_pld_pma_adapt_done),
				.pld_pma_clklow(w_hssi_common_pld_pcs_interface_pld_pma_clklow),
				.pld_pma_fref(w_hssi_common_pld_pcs_interface_pld_pma_fref),
				.pld_pma_hclk(w_hssi_common_pld_pcs_interface_pld_pma_hclk),
				.pld_pma_pcie_sw_done(w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done),
				.pld_pma_pfdmode_lock(w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock),
				.pld_pma_reserved_in(w_hssi_common_pld_pcs_interface_pld_pma_reserved_in),
				.pld_pma_rx_detect_valid(w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid),
				.pld_pma_rx_found(w_hssi_common_pld_pcs_interface_pld_pma_rx_found),
				.pld_pma_rxpll_lock(w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock),
				.pld_pma_testbus(w_hssi_common_pld_pcs_interface_pld_pma_testbus),
				.pld_pmaif_mask_tx_pll(w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll),
				.pld_reserved_out(w_hssi_common_pld_pcs_interface_pld_reserved_out),
				.pld_test_data(w_hssi_common_pld_pcs_interface_pld_test_data),
				.pld_uhsif_lock(w_hssi_common_pld_pcs_interface_pld_uhsif_lock),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.int_pldif_10g_test_data({w_hssi_10g_tx_pcs_tx_test_data[19], w_hssi_10g_tx_pcs_tx_test_data[18], w_hssi_10g_tx_pcs_tx_test_data[17], w_hssi_10g_tx_pcs_tx_test_data[16], w_hssi_10g_tx_pcs_tx_test_data[15], w_hssi_10g_tx_pcs_tx_test_data[14], w_hssi_10g_tx_pcs_tx_test_data[13], w_hssi_10g_tx_pcs_tx_test_data[12], w_hssi_10g_tx_pcs_tx_test_data[11], w_hssi_10g_tx_pcs_tx_test_data[10], w_hssi_10g_tx_pcs_tx_test_data[9], w_hssi_10g_tx_pcs_tx_test_data[8], w_hssi_10g_tx_pcs_tx_test_data[7], w_hssi_10g_tx_pcs_tx_test_data[6], w_hssi_10g_tx_pcs_tx_test_data[5], w_hssi_10g_tx_pcs_tx_test_data[4], w_hssi_10g_tx_pcs_tx_test_data[3], w_hssi_10g_tx_pcs_tx_test_data[2], w_hssi_10g_tx_pcs_tx_test_data[1], w_hssi_10g_tx_pcs_tx_test_data[0]}),
				.int_pldif_10g_tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.int_pldif_8g_chnl_test_bus_out({w_hssi_8g_rx_pcs_chnl_test_bus_out[19], w_hssi_8g_rx_pcs_chnl_test_bus_out[18], w_hssi_8g_rx_pcs_chnl_test_bus_out[17], w_hssi_8g_rx_pcs_chnl_test_bus_out[16], w_hssi_8g_rx_pcs_chnl_test_bus_out[15], w_hssi_8g_rx_pcs_chnl_test_bus_out[14], w_hssi_8g_rx_pcs_chnl_test_bus_out[13], w_hssi_8g_rx_pcs_chnl_test_bus_out[12], w_hssi_8g_rx_pcs_chnl_test_bus_out[11], w_hssi_8g_rx_pcs_chnl_test_bus_out[10], w_hssi_8g_rx_pcs_chnl_test_bus_out[9], w_hssi_8g_rx_pcs_chnl_test_bus_out[8], w_hssi_8g_rx_pcs_chnl_test_bus_out[7], w_hssi_8g_rx_pcs_chnl_test_bus_out[6], w_hssi_8g_rx_pcs_chnl_test_bus_out[5], w_hssi_8g_rx_pcs_chnl_test_bus_out[4], w_hssi_8g_rx_pcs_chnl_test_bus_out[3], w_hssi_8g_rx_pcs_chnl_test_bus_out[2], w_hssi_8g_rx_pcs_chnl_test_bus_out[1], w_hssi_8g_rx_pcs_chnl_test_bus_out[0]}),
				.int_pldif_8g_rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.int_pldif_8g_tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.int_pldif_g3_test_out({w_hssi_pipe_gen3_test_out[19], w_hssi_pipe_gen3_test_out[18], w_hssi_pipe_gen3_test_out[17], w_hssi_pipe_gen3_test_out[16], w_hssi_pipe_gen3_test_out[15], w_hssi_pipe_gen3_test_out[14], w_hssi_pipe_gen3_test_out[13], w_hssi_pipe_gen3_test_out[12], w_hssi_pipe_gen3_test_out[11], w_hssi_pipe_gen3_test_out[10], w_hssi_pipe_gen3_test_out[9], w_hssi_pipe_gen3_test_out[8], w_hssi_pipe_gen3_test_out[7], w_hssi_pipe_gen3_test_out[6], w_hssi_pipe_gen3_test_out[5], w_hssi_pipe_gen3_test_out[4], w_hssi_pipe_gen3_test_out[3], w_hssi_pipe_gen3_test_out[2], w_hssi_pipe_gen3_test_out[1], w_hssi_pipe_gen3_test_out[0]}),
				.int_pldif_krfec_test_data({w_hssi_krfec_tx_pcs_tx_test_data[19], w_hssi_krfec_tx_pcs_tx_test_data[18], w_hssi_krfec_tx_pcs_tx_test_data[17], w_hssi_krfec_tx_pcs_tx_test_data[16], w_hssi_krfec_tx_pcs_tx_test_data[15], w_hssi_krfec_tx_pcs_tx_test_data[14], w_hssi_krfec_tx_pcs_tx_test_data[13], w_hssi_krfec_tx_pcs_tx_test_data[12], w_hssi_krfec_tx_pcs_tx_test_data[11], w_hssi_krfec_tx_pcs_tx_test_data[10], w_hssi_krfec_tx_pcs_tx_test_data[9], w_hssi_krfec_tx_pcs_tx_test_data[8], w_hssi_krfec_tx_pcs_tx_test_data[7], w_hssi_krfec_tx_pcs_tx_test_data[6], w_hssi_krfec_tx_pcs_tx_test_data[5], w_hssi_krfec_tx_pcs_tx_test_data[4], w_hssi_krfec_tx_pcs_tx_test_data[3], w_hssi_krfec_tx_pcs_tx_test_data[2], w_hssi_krfec_tx_pcs_tx_test_data[1], w_hssi_krfec_tx_pcs_tx_test_data[0]}),
				.int_pldif_pmaif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pldif_pmaif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pldif_pmaif_pcie_sw_done({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0]}),
				.int_pldif_pmaif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pldif_pmaif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pldif_pmaif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pldif_pmaif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pldif_pmaif_pma_reserved_in({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0]}),
				.int_pldif_pmaif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pldif_pmaif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_test_out({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0]}),
				.int_pldif_pmaif_testbus({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0]}),
				.int_pldif_pmaif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.pld_8g_eidleinfersel({in_pld_8g_eidleinfersel[2], in_pld_8g_eidleinfersel[1], in_pld_8g_eidleinfersel[0]}),
				.pld_8g_refclk_dig2(in_pld_8g_refclk_dig2),
				.pld_atpg_los_en_n(in_pld_atpg_los_en_n),
				.pld_g3_current_coeff({in_pld_g3_current_coeff[17], in_pld_g3_current_coeff[16], in_pld_g3_current_coeff[15], in_pld_g3_current_coeff[14], in_pld_g3_current_coeff[13], in_pld_g3_current_coeff[12], in_pld_g3_current_coeff[11], in_pld_g3_current_coeff[10], in_pld_g3_current_coeff[9], in_pld_g3_current_coeff[8], in_pld_g3_current_coeff[7], in_pld_g3_current_coeff[6], in_pld_g3_current_coeff[5], in_pld_g3_current_coeff[4], in_pld_g3_current_coeff[3], in_pld_g3_current_coeff[2], in_pld_g3_current_coeff[1], in_pld_g3_current_coeff[0]}),
				.pld_g3_current_rxpreset({in_pld_g3_current_rxpreset[2], in_pld_g3_current_rxpreset[1], in_pld_g3_current_rxpreset[0]}),
				.pld_ltr(in_pld_ltr),
				.pld_mem_krfec_atpg_rst_n(in_pld_mem_krfec_atpg_rst_n),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pcs_refclk_dig(in_pld_pcs_refclk_dig),
				.pld_pma_adapt_start(in_pld_pma_adapt_start),
				.pld_pma_csr_test_dis(in_pld_pma_csr_test_dis),
				.pld_pma_early_eios(in_pld_pma_early_eios),
				.pld_pma_eye_monitor({in_pld_pma_eye_monitor[5], in_pld_pma_eye_monitor[4], in_pld_pma_eye_monitor[3], in_pld_pma_eye_monitor[2], in_pld_pma_eye_monitor[1], in_pld_pma_eye_monitor[0]}),
				.pld_pma_ltd_b(in_pld_pma_ltd_b),
				.pld_pma_nrpi_freeze(in_pld_pma_nrpi_freeze),
				.pld_pma_pcie_switch({in_pld_pma_pcie_switch[1], in_pld_pma_pcie_switch[0]}),
				.pld_pma_ppm_lock(in_pld_pma_ppm_lock),
				.pld_pma_reserved_out({in_pld_pma_reserved_out[4], in_pld_pma_reserved_out[3], in_pld_pma_reserved_out[2], in_pld_pma_reserved_out[1], in_pld_pma_reserved_out[0]}),
				.pld_pma_rs_lpbk_b(in_pld_pma_rs_lpbk_b),
				.pld_pma_rx_qpi_pullup(in_pld_pma_rx_qpi_pullup),
				.pld_pma_tx_bitslip(in_pld_pma_tx_bitslip),
				.pld_pma_tx_bonding_rstb(in_pld_pma_tx_bonding_rstb),
				.pld_pma_tx_qpi_pulldn(in_pld_pma_tx_qpi_pulldn),
				.pld_pma_tx_qpi_pullup(in_pld_pma_tx_qpi_pullup),
				.pld_pma_txdetectrx(in_pld_pma_txdetectrx),
				.pld_rate({in_pld_rate[1], in_pld_rate[0]}),
				.pld_reserved_in({in_pld_reserved_in[9], in_pld_reserved_in[8], in_pld_reserved_in[7], in_pld_reserved_in[6], in_pld_reserved_in[5], in_pld_reserved_in[4], in_pld_reserved_in[3], in_pld_reserved_in[2], in_pld_reserved_in[1], in_pld_reserved_in[0]}),
				.pld_scan_mode_n(in_pld_scan_mode_n),
				.pld_scan_shift_n(in_pld_scan_shift_n),
				
				// UNUSED
				.int_pldif_8g_ltr(),
				.int_pldif_avmm_pld_avmm1_request(),
				.int_pldif_avmm_pld_avmm2_request(),
				.int_pldif_avmm_refclk_dig_en(),
				.int_pldif_g3_scan_mode_n(),
				.pld_8g_eidleinfersel_fifo(),
				.pld_8g_eidleinfersel_reg(),
				.pld_partial_reconfig_fifo(),
				.pld_partial_reconfig_rx_div_by_2_rxclk_wire(),
				.pld_partial_reconfig_rx_div_by_2_txclk_wire(),
				.pld_partial_reconfig_rxclk_reg(),
				.pld_partial_reconfig_tx_div_by_2_wire(),
				.pld_partial_reconfig_txclk_reg(),
				.pld_rate_reg(),
				.pld_test_data_reg()
			);
		end // if generate
		else begin
				assign w_hssi_common_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_clk[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_npor = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_usermode = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2 = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_adapt_done = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_clklow = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_fref = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_hclk = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_found = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_testbus[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_reserved_out[9:0] = 10'b0;
				assign w_hssi_common_pld_pcs_interface_pld_test_data[19:0] = 20'b0;
				assign w_hssi_common_pld_pcs_interface_pld_uhsif_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_scan_mode_n = 1'b1;		// Override default tieoff
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_rx_pcs
			twentynm_hssi_fifo_rx_pcs #(
				.double_read_mode(hssi_fifo_rx_pcs_double_read_mode),
				.prot_mode(hssi_fifo_rx_pcs_prot_mode),
				.silicon_rev( "20nm5es2" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_rx_pcs_blockselect),
				.data_out2_10g(w_hssi_fifo_rx_pcs_data_out2_10g),
				.data_out2_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp),
				.data_out_10g(w_hssi_fifo_rx_pcs_data_out_10g),
				.data_out_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out_8g_clock_comp),
				.data_out_8g_phase_comp(w_hssi_fifo_rx_pcs_data_out_8g_phase_comp),
				.data_out_gen3(w_hssi_fifo_rx_pcs_data_out_gen3),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_data[73], w_hssi_10g_rx_pcs_rx_fifo_wr_data[72], w_hssi_10g_rx_pcs_rx_fifo_wr_data[71], w_hssi_10g_rx_pcs_rx_fifo_wr_data[70], w_hssi_10g_rx_pcs_rx_fifo_wr_data[69], w_hssi_10g_rx_pcs_rx_fifo_wr_data[68], w_hssi_10g_rx_pcs_rx_fifo_wr_data[67], w_hssi_10g_rx_pcs_rx_fifo_wr_data[66], w_hssi_10g_rx_pcs_rx_fifo_wr_data[65], w_hssi_10g_rx_pcs_rx_fifo_wr_data[64], w_hssi_10g_rx_pcs_rx_fifo_wr_data[63], w_hssi_10g_rx_pcs_rx_fifo_wr_data[62], w_hssi_10g_rx_pcs_rx_fifo_wr_data[61], w_hssi_10g_rx_pcs_rx_fifo_wr_data[60], w_hssi_10g_rx_pcs_rx_fifo_wr_data[59], w_hssi_10g_rx_pcs_rx_fifo_wr_data[58], w_hssi_10g_rx_pcs_rx_fifo_wr_data[57], w_hssi_10g_rx_pcs_rx_fifo_wr_data[56], w_hssi_10g_rx_pcs_rx_fifo_wr_data[55], w_hssi_10g_rx_pcs_rx_fifo_wr_data[54], w_hssi_10g_rx_pcs_rx_fifo_wr_data[53], w_hssi_10g_rx_pcs_rx_fifo_wr_data[52], w_hssi_10g_rx_pcs_rx_fifo_wr_data[51], w_hssi_10g_rx_pcs_rx_fifo_wr_data[50], w_hssi_10g_rx_pcs_rx_fifo_wr_data[49], w_hssi_10g_rx_pcs_rx_fifo_wr_data[48], w_hssi_10g_rx_pcs_rx_fifo_wr_data[47], w_hssi_10g_rx_pcs_rx_fifo_wr_data[46], w_hssi_10g_rx_pcs_rx_fifo_wr_data[45], w_hssi_10g_rx_pcs_rx_fifo_wr_data[44], w_hssi_10g_rx_pcs_rx_fifo_wr_data[43], w_hssi_10g_rx_pcs_rx_fifo_wr_data[42], w_hssi_10g_rx_pcs_rx_fifo_wr_data[41], w_hssi_10g_rx_pcs_rx_fifo_wr_data[40], w_hssi_10g_rx_pcs_rx_fifo_wr_data[39], w_hssi_10g_rx_pcs_rx_fifo_wr_data[38], w_hssi_10g_rx_pcs_rx_fifo_wr_data[37], w_hssi_10g_rx_pcs_rx_fifo_wr_data[36], w_hssi_10g_rx_pcs_rx_fifo_wr_data[35], w_hssi_10g_rx_pcs_rx_fifo_wr_data[34], w_hssi_10g_rx_pcs_rx_fifo_wr_data[33], w_hssi_10g_rx_pcs_rx_fifo_wr_data[32], w_hssi_10g_rx_pcs_rx_fifo_wr_data[31], w_hssi_10g_rx_pcs_rx_fifo_wr_data[30], w_hssi_10g_rx_pcs_rx_fifo_wr_data[29], w_hssi_10g_rx_pcs_rx_fifo_wr_data[28], w_hssi_10g_rx_pcs_rx_fifo_wr_data[27], w_hssi_10g_rx_pcs_rx_fifo_wr_data[26], w_hssi_10g_rx_pcs_rx_fifo_wr_data[25], w_hssi_10g_rx_pcs_rx_fifo_wr_data[24], w_hssi_10g_rx_pcs_rx_fifo_wr_data[23], w_hssi_10g_rx_pcs_rx_fifo_wr_data[22], w_hssi_10g_rx_pcs_rx_fifo_wr_data[21], w_hssi_10g_rx_pcs_rx_fifo_wr_data[20], w_hssi_10g_rx_pcs_rx_fifo_wr_data[19], w_hssi_10g_rx_pcs_rx_fifo_wr_data[18], w_hssi_10g_rx_pcs_rx_fifo_wr_data[17], w_hssi_10g_rx_pcs_rx_fifo_wr_data[16], w_hssi_10g_rx_pcs_rx_fifo_wr_data[15], w_hssi_10g_rx_pcs_rx_fifo_wr_data[14], w_hssi_10g_rx_pcs_rx_fifo_wr_data[13], w_hssi_10g_rx_pcs_rx_fifo_wr_data[12], w_hssi_10g_rx_pcs_rx_fifo_wr_data[11], w_hssi_10g_rx_pcs_rx_fifo_wr_data[10], w_hssi_10g_rx_pcs_rx_fifo_wr_data[9], w_hssi_10g_rx_pcs_rx_fifo_wr_data[8], w_hssi_10g_rx_pcs_rx_fifo_wr_data[7], w_hssi_10g_rx_pcs_rx_fifo_wr_data[6], w_hssi_10g_rx_pcs_rx_fifo_wr_data[5], w_hssi_10g_rx_pcs_rx_fifo_wr_data[4], w_hssi_10g_rx_pcs_rx_fifo_wr_data[3], w_hssi_10g_rx_pcs_rx_fifo_wr_data[2], w_hssi_10g_rx_pcs_rx_fifo_wr_data[1], w_hssi_10g_rx_pcs_rx_fifo_wr_data[0]}),
				.data_in_8g_clock_comp({w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0]}),
				.data_in_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr2_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0]}),
				.rd_ptr2_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0]}),
				.rd_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0]}),
				.rd_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.wr_clk_8g_clock_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_8g_clock_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.wr_en_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.wr_en_8g_clock_comp(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_en_8g_phase_comp(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.wr_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0]}),
				.wr_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0]}),
				.wr_rst_n_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.wr_rst_n_8g_clock_comp(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_n_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_rx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79:0] = 80'b0;
				assign w_hssi_fifo_rx_pcs_data_out_gen3[39:0] = 40'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_tx_pcs
			twentynm_hssi_fifo_tx_pcs #(
				.double_write_mode(hssi_fifo_tx_pcs_double_write_mode),
				.prot_mode(hssi_fifo_tx_pcs_prot_mode),
				.silicon_rev( "20nm5es2" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_tx_pcs_blockselect),
				.data_out_10g(w_hssi_fifo_tx_pcs_data_out_10g),
				.data_out_8g_phase_comp(w_hssi_fifo_tx_pcs_data_out_8g_phase_comp),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in2_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0]}),
				.data_in_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_en_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.wr_en_8g_phase_comp(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0]}),
				.wr_rst_n_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_tx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_tx_pcs_data_out_10g[72:0] = 73'b0;
				assign w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63:0] = 64'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_rx_pcs
			twentynm_hssi_gen3_rx_pcs #(
				.block_sync(hssi_gen3_rx_pcs_block_sync),
				.block_sync_sm(hssi_gen3_rx_pcs_block_sync_sm),
				.cdr_ctrl_force_unalgn(hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn),
				.lpbk_force(hssi_gen3_rx_pcs_lpbk_force),
				.mode(hssi_gen3_rx_pcs_mode),
				.rate_match_fifo(hssi_gen3_rx_pcs_rate_match_fifo),
				.rate_match_fifo_latency(hssi_gen3_rx_pcs_rate_match_fifo_latency),
				.reconfig_settings(hssi_gen3_rx_pcs_reconfig_settings),
				.reverse_lpbk(hssi_gen3_rx_pcs_reverse_lpbk),
				.rx_b4gb_par_lpbk(hssi_gen3_rx_pcs_rx_b4gb_par_lpbk),
				.rx_force_balign(hssi_gen3_rx_pcs_rx_force_balign),
				.rx_ins_del_one_skip(hssi_gen3_rx_pcs_rx_ins_del_one_skip),
				.rx_num_fixed_pat(hssi_gen3_rx_pcs_rx_num_fixed_pat),
				.rx_test_out_sel(hssi_gen3_rx_pcs_rx_test_out_sel),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_rx_pcs_sup_mode)
			) inst_twentynm_hssi_gen3_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_rx_pcs_avmmreaddata),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.blk_start(w_hssi_gen3_rx_pcs_blk_start),
				.blockselect(w_hssi_gen3_rx_pcs_blockselect),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.data_out(w_hssi_gen3_rx_pcs_data_out),
				.data_valid(w_hssi_gen3_rx_pcs_data_valid),
				.ei_det_int(w_hssi_gen3_rx_pcs_ei_det_int),
				.ei_partial_det_int(w_hssi_gen3_rx_pcs_ei_partial_det_int),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.i_det_int(w_hssi_gen3_rx_pcs_i_det_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data(w_hssi_gen3_rx_pcs_lpbk_data),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.mem_rx_fifo_rd_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr),
				.mem_rx_fifo_wr_clk(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.mem_rx_fifo_wr_data(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data),
				.mem_rx_fifo_wr_en(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.mem_rx_fifo_wr_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr),
				.mem_rx_fifo_wr_rst_n(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_test_out(w_hssi_gen3_rx_pcs_rx_test_out),
				.sync_hdr(w_hssi_gen3_rx_pcs_sync_hdr),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0]}),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.mem_rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_gen3[39], w_hssi_fifo_rx_pcs_data_out_gen3[38], w_hssi_fifo_rx_pcs_data_out_gen3[37], w_hssi_fifo_rx_pcs_data_out_gen3[36], w_hssi_fifo_rx_pcs_data_out_gen3[35], w_hssi_fifo_rx_pcs_data_out_gen3[34], w_hssi_fifo_rx_pcs_data_out_gen3[33], w_hssi_fifo_rx_pcs_data_out_gen3[32], w_hssi_fifo_rx_pcs_data_out_gen3[31], w_hssi_fifo_rx_pcs_data_out_gen3[30], w_hssi_fifo_rx_pcs_data_out_gen3[29], w_hssi_fifo_rx_pcs_data_out_gen3[28], w_hssi_fifo_rx_pcs_data_out_gen3[27], w_hssi_fifo_rx_pcs_data_out_gen3[26], w_hssi_fifo_rx_pcs_data_out_gen3[25], w_hssi_fifo_rx_pcs_data_out_gen3[24], w_hssi_fifo_rx_pcs_data_out_gen3[23], w_hssi_fifo_rx_pcs_data_out_gen3[22], w_hssi_fifo_rx_pcs_data_out_gen3[21], w_hssi_fifo_rx_pcs_data_out_gen3[20], w_hssi_fifo_rx_pcs_data_out_gen3[19], w_hssi_fifo_rx_pcs_data_out_gen3[18], w_hssi_fifo_rx_pcs_data_out_gen3[17], w_hssi_fifo_rx_pcs_data_out_gen3[16], w_hssi_fifo_rx_pcs_data_out_gen3[15], w_hssi_fifo_rx_pcs_data_out_gen3[14], w_hssi_fifo_rx_pcs_data_out_gen3[13], w_hssi_fifo_rx_pcs_data_out_gen3[12], w_hssi_fifo_rx_pcs_data_out_gen3[11], w_hssi_fifo_rx_pcs_data_out_gen3[10], w_hssi_fifo_rx_pcs_data_out_gen3[9], w_hssi_fifo_rx_pcs_data_out_gen3[8], w_hssi_fifo_rx_pcs_data_out_gen3[7], w_hssi_fifo_rx_pcs_data_out_gen3[6], w_hssi_fifo_rx_pcs_data_out_gen3[5], w_hssi_fifo_rx_pcs_data_out_gen3[4], w_hssi_fifo_rx_pcs_data_out_gen3[3], w_hssi_fifo_rx_pcs_data_out_gen3[2], w_hssi_fifo_rx_pcs_data_out_gen3[1], w_hssi_fifo_rx_pcs_data_out_gen3[0]}),
				.par_lpbk_b4gb_in({w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0]}),
				.par_lpbk_in({w_hssi_gen3_tx_pcs_par_lpbk_out[31], w_hssi_gen3_tx_pcs_par_lpbk_out[30], w_hssi_gen3_tx_pcs_par_lpbk_out[29], w_hssi_gen3_tx_pcs_par_lpbk_out[28], w_hssi_gen3_tx_pcs_par_lpbk_out[27], w_hssi_gen3_tx_pcs_par_lpbk_out[26], w_hssi_gen3_tx_pcs_par_lpbk_out[25], w_hssi_gen3_tx_pcs_par_lpbk_out[24], w_hssi_gen3_tx_pcs_par_lpbk_out[23], w_hssi_gen3_tx_pcs_par_lpbk_out[22], w_hssi_gen3_tx_pcs_par_lpbk_out[21], w_hssi_gen3_tx_pcs_par_lpbk_out[20], w_hssi_gen3_tx_pcs_par_lpbk_out[19], w_hssi_gen3_tx_pcs_par_lpbk_out[18], w_hssi_gen3_tx_pcs_par_lpbk_out[17], w_hssi_gen3_tx_pcs_par_lpbk_out[16], w_hssi_gen3_tx_pcs_par_lpbk_out[15], w_hssi_gen3_tx_pcs_par_lpbk_out[14], w_hssi_gen3_tx_pcs_par_lpbk_out[13], w_hssi_gen3_tx_pcs_par_lpbk_out[12], w_hssi_gen3_tx_pcs_par_lpbk_out[11], w_hssi_gen3_tx_pcs_par_lpbk_out[10], w_hssi_gen3_tx_pcs_par_lpbk_out[9], w_hssi_gen3_tx_pcs_par_lpbk_out[8], w_hssi_gen3_tx_pcs_par_lpbk_out[7], w_hssi_gen3_tx_pcs_par_lpbk_out[6], w_hssi_gen3_tx_pcs_par_lpbk_out[5], w_hssi_gen3_tx_pcs_par_lpbk_out[4], w_hssi_gen3_tx_pcs_par_lpbk_out[3], w_hssi_gen3_tx_pcs_par_lpbk_out[2], w_hssi_gen3_tx_pcs_par_lpbk_out[1], w_hssi_gen3_tx_pcs_par_lpbk_out[0]}),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.rcvd_clk(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_pma_clk(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.rxpolarity(w_hssi_pipe_gen3_rxpolarity_int),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.sync_sm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.txdatak_in({w_hssi_pipe_gen3_txdatak_int[3], w_hssi_pipe_gen3_txdatak_int[2], w_hssi_pipe_gen3_txdatak_int[1], w_hssi_pipe_gen3_txdatak_int[0]}),
				
				// UNUSED
				.blk_lockd_int(),
				.skp_det_int()
			);
		end // if generate
		else begin
				assign w_hssi_gen3_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_rx_pcs_blk_algnd_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_delete_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_insert_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_overfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_undfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_rx_pcs_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_partial_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_err_decode_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_i_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data[33:0] = 34'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39:0] = 40'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_rx_test_out[19:0] = 20'b0;
				assign w_hssi_gen3_rx_pcs_sync_hdr[1:0] = 2'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_tx_pcs
			twentynm_hssi_gen3_tx_pcs #(
				.mode(hssi_gen3_tx_pcs_mode),
				.reverse_lpbk(hssi_gen3_tx_pcs_reverse_lpbk),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_tx_pcs_sup_mode),
				.tx_bitslip(hssi_gen3_tx_pcs_tx_bitslip),
				.tx_gbox_byp(hssi_gen3_tx_pcs_tx_gbox_byp)
			) inst_twentynm_hssi_gen3_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_gen3_tx_pcs_blockselect),
				.data_out(w_hssi_gen3_tx_pcs_data_out),
				.par_lpbk_b4gb_out(w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out),
				.par_lpbk_out(w_hssi_gen3_tx_pcs_par_lpbk_out),
				.tx_test_out(w_hssi_gen3_tx_pcs_tx_test_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_start_in(w_hssi_pipe_gen3_tx_blk_start_int),
				.data_in({w_hssi_pipe_gen3_txdata_int[31], w_hssi_pipe_gen3_txdata_int[30], w_hssi_pipe_gen3_txdata_int[29], w_hssi_pipe_gen3_txdata_int[28], w_hssi_pipe_gen3_txdata_int[27], w_hssi_pipe_gen3_txdata_int[26], w_hssi_pipe_gen3_txdata_int[25], w_hssi_pipe_gen3_txdata_int[24], w_hssi_pipe_gen3_txdata_int[23], w_hssi_pipe_gen3_txdata_int[22], w_hssi_pipe_gen3_txdata_int[21], w_hssi_pipe_gen3_txdata_int[20], w_hssi_pipe_gen3_txdata_int[19], w_hssi_pipe_gen3_txdata_int[18], w_hssi_pipe_gen3_txdata_int[17], w_hssi_pipe_gen3_txdata_int[16], w_hssi_pipe_gen3_txdata_int[15], w_hssi_pipe_gen3_txdata_int[14], w_hssi_pipe_gen3_txdata_int[13], w_hssi_pipe_gen3_txdata_int[12], w_hssi_pipe_gen3_txdata_int[11], w_hssi_pipe_gen3_txdata_int[10], w_hssi_pipe_gen3_txdata_int[9], w_hssi_pipe_gen3_txdata_int[8], w_hssi_pipe_gen3_txdata_int[7], w_hssi_pipe_gen3_txdata_int[6], w_hssi_pipe_gen3_txdata_int[5], w_hssi_pipe_gen3_txdata_int[4], w_hssi_pipe_gen3_txdata_int[3], w_hssi_pipe_gen3_txdata_int[2], w_hssi_pipe_gen3_txdata_int[1], w_hssi_pipe_gen3_txdata_int[0]}),
				.data_valid(w_hssi_pipe_gen3_txdataskip_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data_in({w_hssi_gen3_rx_pcs_lpbk_data[33], w_hssi_gen3_rx_pcs_lpbk_data[32], w_hssi_gen3_rx_pcs_lpbk_data[31], w_hssi_gen3_rx_pcs_lpbk_data[30], w_hssi_gen3_rx_pcs_lpbk_data[29], w_hssi_gen3_rx_pcs_lpbk_data[28], w_hssi_gen3_rx_pcs_lpbk_data[27], w_hssi_gen3_rx_pcs_lpbk_data[26], w_hssi_gen3_rx_pcs_lpbk_data[25], w_hssi_gen3_rx_pcs_lpbk_data[24], w_hssi_gen3_rx_pcs_lpbk_data[23], w_hssi_gen3_rx_pcs_lpbk_data[22], w_hssi_gen3_rx_pcs_lpbk_data[21], w_hssi_gen3_rx_pcs_lpbk_data[20], w_hssi_gen3_rx_pcs_lpbk_data[19], w_hssi_gen3_rx_pcs_lpbk_data[18], w_hssi_gen3_rx_pcs_lpbk_data[17], w_hssi_gen3_rx_pcs_lpbk_data[16], w_hssi_gen3_rx_pcs_lpbk_data[15], w_hssi_gen3_rx_pcs_lpbk_data[14], w_hssi_gen3_rx_pcs_lpbk_data[13], w_hssi_gen3_rx_pcs_lpbk_data[12], w_hssi_gen3_rx_pcs_lpbk_data[11], w_hssi_gen3_rx_pcs_lpbk_data[10], w_hssi_gen3_rx_pcs_lpbk_data[9], w_hssi_gen3_rx_pcs_lpbk_data[8], w_hssi_gen3_rx_pcs_lpbk_data[7], w_hssi_gen3_rx_pcs_lpbk_data[6], w_hssi_gen3_rx_pcs_lpbk_data[5], w_hssi_gen3_rx_pcs_lpbk_data[4], w_hssi_gen3_rx_pcs_lpbk_data[3], w_hssi_gen3_rx_pcs_lpbk_data[2], w_hssi_gen3_rx_pcs_lpbk_data[1], w_hssi_gen3_rx_pcs_lpbk_data[0]}),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.sync_in({w_hssi_pipe_gen3_tx_sync_hdr_int[1], w_hssi_pipe_gen3_tx_sync_hdr_int[0]}),
				.tx_pma_clk(w_hssi_8g_tx_pcs_clk_out_gen3),
				.tx_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn)
			);
		end // if generate
		else begin
				assign w_hssi_gen3_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_tx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_tx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35:0] = 36'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_tx_test_out[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_rx_pcs
			twentynm_hssi_krfec_rx_pcs #(
				.blksync_cor_en(hssi_krfec_rx_pcs_blksync_cor_en),
				.bypass_gb(hssi_krfec_rx_pcs_bypass_gb),
				.clr_ctrl(hssi_krfec_rx_pcs_clr_ctrl),
				.ctrl_bit_reverse(hssi_krfec_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_rx_pcs_data_bit_reverse),
				.dv_start(hssi_krfec_rx_pcs_dv_start),
				.err_mark_type(hssi_krfec_rx_pcs_err_mark_type),
				.error_marking_en(hssi_krfec_rx_pcs_error_marking_en),
				.low_latency_en(hssi_krfec_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_krfec_rx_pcs_lpbk_mode),
				.parity_invalid_enum(hssi_krfec_rx_pcs_parity_invalid_enum),
				.parity_valid_num(hssi_krfec_rx_pcs_parity_valid_num),
				.pipeln_blksync(hssi_krfec_rx_pcs_pipeln_blksync),
				.pipeln_descrm(hssi_krfec_rx_pcs_pipeln_descrm),
				.pipeln_errcorrect(hssi_krfec_rx_pcs_pipeln_errcorrect),
				.pipeln_errtrap_ind(hssi_krfec_rx_pcs_pipeln_errtrap_ind),
				.pipeln_errtrap_lfsr(hssi_krfec_rx_pcs_pipeln_errtrap_lfsr),
				.pipeln_errtrap_loc(hssi_krfec_rx_pcs_pipeln_errtrap_loc),
				.pipeln_errtrap_pat(hssi_krfec_rx_pcs_pipeln_errtrap_pat),
				.pipeln_gearbox(hssi_krfec_rx_pcs_pipeln_gearbox),
				.pipeln_syndrm(hssi_krfec_rx_pcs_pipeln_syndrm),
				.pipeln_trans_dec(hssi_krfec_rx_pcs_pipeln_trans_dec),
				.prot_mode(hssi_krfec_rx_pcs_prot_mode),
				.receive_order(hssi_krfec_rx_pcs_receive_order),
				.reconfig_settings(hssi_krfec_rx_pcs_reconfig_settings),
				.rx_testbus_sel(hssi_krfec_rx_pcs_rx_testbus_sel),
				.signal_ok_en(hssi_krfec_rx_pcs_signal_ok_en),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_rx_pcs_sup_mode)
			) inst_twentynm_hssi_krfec_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_rx_pcs_blockselect),
				.rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.rx_control_out(w_hssi_krfec_rx_pcs_rx_control_out),
				.rx_data_out(w_hssi_krfec_rx_pcs_rx_data_out),
				.rx_data_status(w_hssi_krfec_rx_pcs_rx_data_status),
				.rx_data_valid_out(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.rx_signal_ok_out(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.rx_data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0]}),
				.rx_krfec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_krfec_reg(),
				.pld_10g_krfec_rx_blk_lock_krfec_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg(),
				.pld_10g_krfec_rx_frame_krfec_reg(),
				.pld_10g_krfec_rx_frame_krfec_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_rx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_block_lock = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_control_out[9:0] = 10'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_status[1:0] = 2'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_valid_out = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_frame = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_signal_ok_out = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_tx_pcs
			twentynm_hssi_krfec_tx_pcs #(
				.burst_err(hssi_krfec_tx_pcs_burst_err),
				.burst_err_len(hssi_krfec_tx_pcs_burst_err_len),
				.ctrl_bit_reverse(hssi_krfec_tx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_tx_pcs_data_bit_reverse),
				.enc_frame_query(hssi_krfec_tx_pcs_enc_frame_query),
				.low_latency_en(hssi_krfec_tx_pcs_low_latency_en),
				.pipeln_encoder(hssi_krfec_tx_pcs_pipeln_encoder),
				.pipeln_scrambler(hssi_krfec_tx_pcs_pipeln_scrambler),
				.prot_mode(hssi_krfec_tx_pcs_prot_mode),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_tx_pcs_sup_mode),
				.transcode_err(hssi_krfec_tx_pcs_transcode_err),
				.transmit_order(hssi_krfec_tx_pcs_transmit_order),
				.tx_testbus_sel(hssi_krfec_tx_pcs_tx_testbus_sel)
			) inst_twentynm_hssi_krfec_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_tx_pcs_blockselect),
				.tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.tx_data_out(w_hssi_krfec_tx_pcs_tx_data_out),
				.tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.tx_test_data(w_hssi_krfec_tx_pcs_tx_test_data),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.tx_control_in({w_hssi_10g_tx_pcs_tx_control_out_krfec[8], w_hssi_10g_tx_pcs_tx_control_out_krfec[7], w_hssi_10g_tx_pcs_tx_control_out_krfec[6], w_hssi_10g_tx_pcs_tx_control_out_krfec[5], w_hssi_10g_tx_pcs_tx_control_out_krfec[4], w_hssi_10g_tx_pcs_tx_control_out_krfec[3], w_hssi_10g_tx_pcs_tx_control_out_krfec[2], w_hssi_10g_tx_pcs_tx_control_out_krfec[1], w_hssi_10g_tx_pcs_tx_control_out_krfec[0]}),
				.tx_data_in({w_hssi_10g_tx_pcs_tx_data_out_krfec[63], w_hssi_10g_tx_pcs_tx_data_out_krfec[62], w_hssi_10g_tx_pcs_tx_data_out_krfec[61], w_hssi_10g_tx_pcs_tx_data_out_krfec[60], w_hssi_10g_tx_pcs_tx_data_out_krfec[59], w_hssi_10g_tx_pcs_tx_data_out_krfec[58], w_hssi_10g_tx_pcs_tx_data_out_krfec[57], w_hssi_10g_tx_pcs_tx_data_out_krfec[56], w_hssi_10g_tx_pcs_tx_data_out_krfec[55], w_hssi_10g_tx_pcs_tx_data_out_krfec[54], w_hssi_10g_tx_pcs_tx_data_out_krfec[53], w_hssi_10g_tx_pcs_tx_data_out_krfec[52], w_hssi_10g_tx_pcs_tx_data_out_krfec[51], w_hssi_10g_tx_pcs_tx_data_out_krfec[50], w_hssi_10g_tx_pcs_tx_data_out_krfec[49], w_hssi_10g_tx_pcs_tx_data_out_krfec[48], w_hssi_10g_tx_pcs_tx_data_out_krfec[47], w_hssi_10g_tx_pcs_tx_data_out_krfec[46], w_hssi_10g_tx_pcs_tx_data_out_krfec[45], w_hssi_10g_tx_pcs_tx_data_out_krfec[44], w_hssi_10g_tx_pcs_tx_data_out_krfec[43], w_hssi_10g_tx_pcs_tx_data_out_krfec[42], w_hssi_10g_tx_pcs_tx_data_out_krfec[41], w_hssi_10g_tx_pcs_tx_data_out_krfec[40], w_hssi_10g_tx_pcs_tx_data_out_krfec[39], w_hssi_10g_tx_pcs_tx_data_out_krfec[38], w_hssi_10g_tx_pcs_tx_data_out_krfec[37], w_hssi_10g_tx_pcs_tx_data_out_krfec[36], w_hssi_10g_tx_pcs_tx_data_out_krfec[35], w_hssi_10g_tx_pcs_tx_data_out_krfec[34], w_hssi_10g_tx_pcs_tx_data_out_krfec[33], w_hssi_10g_tx_pcs_tx_data_out_krfec[32], w_hssi_10g_tx_pcs_tx_data_out_krfec[31], w_hssi_10g_tx_pcs_tx_data_out_krfec[30], w_hssi_10g_tx_pcs_tx_data_out_krfec[29], w_hssi_10g_tx_pcs_tx_data_out_krfec[28], w_hssi_10g_tx_pcs_tx_data_out_krfec[27], w_hssi_10g_tx_pcs_tx_data_out_krfec[26], w_hssi_10g_tx_pcs_tx_data_out_krfec[25], w_hssi_10g_tx_pcs_tx_data_out_krfec[24], w_hssi_10g_tx_pcs_tx_data_out_krfec[23], w_hssi_10g_tx_pcs_tx_data_out_krfec[22], w_hssi_10g_tx_pcs_tx_data_out_krfec[21], w_hssi_10g_tx_pcs_tx_data_out_krfec[20], w_hssi_10g_tx_pcs_tx_data_out_krfec[19], w_hssi_10g_tx_pcs_tx_data_out_krfec[18], w_hssi_10g_tx_pcs_tx_data_out_krfec[17], w_hssi_10g_tx_pcs_tx_data_out_krfec[16], w_hssi_10g_tx_pcs_tx_data_out_krfec[15], w_hssi_10g_tx_pcs_tx_data_out_krfec[14], w_hssi_10g_tx_pcs_tx_data_out_krfec[13], w_hssi_10g_tx_pcs_tx_data_out_krfec[12], w_hssi_10g_tx_pcs_tx_data_out_krfec[11], w_hssi_10g_tx_pcs_tx_data_out_krfec[10], w_hssi_10g_tx_pcs_tx_data_out_krfec[9], w_hssi_10g_tx_pcs_tx_data_out_krfec[8], w_hssi_10g_tx_pcs_tx_data_out_krfec[7], w_hssi_10g_tx_pcs_tx_data_out_krfec[6], w_hssi_10g_tx_pcs_tx_data_out_krfec[5], w_hssi_10g_tx_pcs_tx_data_out_krfec[4], w_hssi_10g_tx_pcs_tx_data_out_krfec[3], w_hssi_10g_tx_pcs_tx_data_out_krfec[2], w_hssi_10g_tx_pcs_tx_data_out_krfec[1], w_hssi_10g_tx_pcs_tx_data_out_krfec[0]}),
				.tx_data_valid_in(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_krfec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_krfec_reg(),
				.pld_krfec_tx_alignment_plddirect_reg(),
				.pld_krfec_tx_alignment_reg()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_tx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_alignment = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_test_data[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen1_2
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen1_2
			twentynm_hssi_pipe_gen1_2 #(
				.elec_idle_delay_val(hssi_pipe_gen1_2_elec_idle_delay_val),
				.error_replace_pad(hssi_pipe_gen1_2_error_replace_pad),
				.hip_mode(hssi_pipe_gen1_2_hip_mode),
				.ind_error_reporting(hssi_pipe_gen1_2_ind_error_reporting),
				.phystatus_delay_val(hssi_pipe_gen1_2_phystatus_delay_val),
				.phystatus_rst_toggle(hssi_pipe_gen1_2_phystatus_rst_toggle),
				.pipe_byte_de_serializer_en(hssi_pipe_gen1_2_pipe_byte_de_serializer_en),
				.prot_mode(hssi_pipe_gen1_2_prot_mode),
				.reconfig_settings(hssi_pipe_gen1_2_reconfig_settings),
				.rx_pipe_enable(hssi_pipe_gen1_2_rx_pipe_enable),
				.rxdetect_bypass(hssi_pipe_gen1_2_rxdetect_bypass),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen1_2_sup_mode),
				.tx_pipe_enable(hssi_pipe_gen1_2_tx_pipe_enable),
				.txswing(hssi_pipe_gen1_2_txswing)
			) inst_twentynm_hssi_pipe_gen1_2 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen1_2_avmmreaddata),
				.blockselect(w_hssi_pipe_gen1_2_blockselect),
				.current_coeff(w_hssi_pipe_gen1_2_current_coeff),
				.phystatus(w_hssi_pipe_gen1_2_phystatus),
				.polarity_inversion_rx(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rev_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.rxelectricalidle_out(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxstatus(w_hssi_pipe_gen1_2_rxstatus),
				.rxvalid(w_hssi_pipe_gen1_2_rxvalid),
				.tx_elec_idle_out(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pipe_rx_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.power_state_transition_done_ena(1'b0),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rev_loopbk_pcs_gen3(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.revloopback(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.rx_pipe_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rxd({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxelectricalidle(w_hssi_8g_rx_pcs_eidle_detected),
				.rxelectricalidle_pcs_gen3(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.rxpolarity_pcs_gen3(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.tx_elec_idle_comp(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.txd_ch({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswingport(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.pld_8g_rxpolarity_pipe3_reg(),
				.rxd_ch(),
				.txd()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen1_2_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen1_2_blockselect = 1'b0;
				assign w_hssi_pipe_gen1_2_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen1_2_phystatus = 1'b0;
				assign w_hssi_pipe_gen1_2_polarity_inversion_rx = 1'b0;
				assign w_hssi_pipe_gen1_2_rev_loopbk = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelectricalidle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen1_2_rxvalid = 1'b0;
				assign w_hssi_pipe_gen1_2_tx_elec_idle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_txdetectrx = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen3
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen3
			twentynm_hssi_pipe_gen3 #(
				.bypass_rx_detection_enable(hssi_pipe_gen3_bypass_rx_detection_enable),
				.bypass_rx_preset(hssi_pipe_gen3_bypass_rx_preset),
				.bypass_rx_preset_enable(hssi_pipe_gen3_bypass_rx_preset_enable),
				.bypass_tx_coefficent(hssi_pipe_gen3_bypass_tx_coefficent),
				.bypass_tx_coefficent_enable(hssi_pipe_gen3_bypass_tx_coefficent_enable),
				.elecidle_delay_g3(hssi_pipe_gen3_elecidle_delay_g3),
				.ind_error_reporting(hssi_pipe_gen3_ind_error_reporting),
				.mode(hssi_pipe_gen3_mode),
				.phy_status_delay_g12(hssi_pipe_gen3_phy_status_delay_g12),
				.phy_status_delay_g3(hssi_pipe_gen3_phy_status_delay_g3),
				.phystatus_rst_toggle_g12(hssi_pipe_gen3_phystatus_rst_toggle_g12),
				.phystatus_rst_toggle_g3(hssi_pipe_gen3_phystatus_rst_toggle_g3),
				.rate_match_pad_insertion(hssi_pipe_gen3_rate_match_pad_insertion),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen3_sup_mode),
				.test_out_sel(hssi_pipe_gen3_test_out_sel)
			) inst_twentynm_hssi_pipe_gen3 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen3_avmmreaddata),
				.blockselect(w_hssi_pipe_gen3_blockselect),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.phystatus(w_hssi_pipe_gen3_phystatus),
				.pma_current_coeff(w_hssi_pipe_gen3_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_pipe_gen3_pma_current_rxpreset),
				.pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.rev_lpbk_8gpcs_out(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.rev_lpbk_int(w_hssi_pipe_gen3_rev_lpbk_int),
				.rx_blk_start(w_hssi_pipe_gen3_rx_blk_start),
				.rx_sync_hdr(w_hssi_pipe_gen3_rx_sync_hdr),
				.rxd_8gpcs_out(w_hssi_pipe_gen3_rxd_8gpcs_out),
				.rxdataskip(w_hssi_pipe_gen3_rxdataskip),
				.rxelecidle(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity_8gpcs_out(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.rxpolarity_int(w_hssi_pipe_gen3_rxpolarity_int),
				.rxstatus(w_hssi_pipe_gen3_rxstatus),
				.rxvalid(w_hssi_pipe_gen3_rxvalid),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.test_out(w_hssi_pipe_gen3_test_out),
				.tx_blk_start_int(w_hssi_pipe_gen3_tx_blk_start_int),
				.tx_sync_hdr_int(w_hssi_pipe_gen3_tx_sync_hdr_int),
				.txdata_int(w_hssi_pipe_gen3_txdata_int),
				.txdatak_int(w_hssi_pipe_gen3_txdatak_int),
				.txdataskip_int(w_hssi_pipe_gen3_txdataskip_int),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.current_coeff({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0]}),
				.current_rxpreset({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0]}),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.pcs_asn_bundling_in({w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0]}),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pipe_tx_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_blk_start_int(w_hssi_gen3_rx_pcs_blk_start),
				.rx_sync_hdr_int({w_hssi_gen3_rx_pcs_sync_hdr[1], w_hssi_gen3_rx_pcs_sync_hdr[0]}),
				.rx_test_out({w_hssi_gen3_rx_pcs_rx_test_out[19], w_hssi_gen3_rx_pcs_rx_test_out[18], w_hssi_gen3_rx_pcs_rx_test_out[17], w_hssi_gen3_rx_pcs_rx_test_out[16], w_hssi_gen3_rx_pcs_rx_test_out[15], w_hssi_gen3_rx_pcs_rx_test_out[14], w_hssi_gen3_rx_pcs_rx_test_out[13], w_hssi_gen3_rx_pcs_rx_test_out[12], w_hssi_gen3_rx_pcs_rx_test_out[11], w_hssi_gen3_rx_pcs_rx_test_out[10], w_hssi_gen3_rx_pcs_rx_test_out[9], w_hssi_gen3_rx_pcs_rx_test_out[8], w_hssi_gen3_rx_pcs_rx_test_out[7], w_hssi_gen3_rx_pcs_rx_test_out[6], w_hssi_gen3_rx_pcs_rx_test_out[5], w_hssi_gen3_rx_pcs_rx_test_out[4], w_hssi_gen3_rx_pcs_rx_test_out[3], w_hssi_gen3_rx_pcs_rx_test_out[2], w_hssi_gen3_rx_pcs_rx_test_out[1], w_hssi_gen3_rx_pcs_rx_test_out[0]}),
				.rxd_8gpcs_in({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxdata_int({w_hssi_gen3_rx_pcs_data_out[31], w_hssi_gen3_rx_pcs_data_out[30], w_hssi_gen3_rx_pcs_data_out[29], w_hssi_gen3_rx_pcs_data_out[28], w_hssi_gen3_rx_pcs_data_out[27], w_hssi_gen3_rx_pcs_data_out[26], w_hssi_gen3_rx_pcs_data_out[25], w_hssi_gen3_rx_pcs_data_out[24], w_hssi_gen3_rx_pcs_data_out[23], w_hssi_gen3_rx_pcs_data_out[22], w_hssi_gen3_rx_pcs_data_out[21], w_hssi_gen3_rx_pcs_data_out[20], w_hssi_gen3_rx_pcs_data_out[19], w_hssi_gen3_rx_pcs_data_out[18], w_hssi_gen3_rx_pcs_data_out[17], w_hssi_gen3_rx_pcs_data_out[16], w_hssi_gen3_rx_pcs_data_out[15], w_hssi_gen3_rx_pcs_data_out[14], w_hssi_gen3_rx_pcs_data_out[13], w_hssi_gen3_rx_pcs_data_out[12], w_hssi_gen3_rx_pcs_data_out[11], w_hssi_gen3_rx_pcs_data_out[10], w_hssi_gen3_rx_pcs_data_out[9], w_hssi_gen3_rx_pcs_data_out[8], w_hssi_gen3_rx_pcs_data_out[7], w_hssi_gen3_rx_pcs_data_out[6], w_hssi_gen3_rx_pcs_data_out[5], w_hssi_gen3_rx_pcs_data_out[4], w_hssi_gen3_rx_pcs_data_out[3], w_hssi_gen3_rx_pcs_data_out[2], w_hssi_gen3_rx_pcs_data_out[1], w_hssi_gen3_rx_pcs_data_out[0]}),
				.rxdatak_int({1'b0, 1'b0, 1'b0, 1'b0}),
				.rxdataskip_int(w_hssi_gen3_rx_pcs_data_valid),
				.rxelecidle_8gpcs_in(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.tx_blk_start(w_hssi_8g_tx_pcs_tx_blk_start_out[0]),
				.tx_sync_hdr({w_hssi_8g_tx_pcs_tx_sync_hdr_out[1], w_hssi_8g_tx_pcs_tx_sync_hdr_out[0]}),
				.tx_test_out({w_hssi_gen3_tx_pcs_tx_test_out[19], w_hssi_gen3_tx_pcs_tx_test_out[18], w_hssi_gen3_tx_pcs_tx_test_out[17], w_hssi_gen3_tx_pcs_tx_test_out[16], w_hssi_gen3_tx_pcs_tx_test_out[15], w_hssi_gen3_tx_pcs_tx_test_out[14], w_hssi_gen3_tx_pcs_tx_test_out[13], w_hssi_gen3_tx_pcs_tx_test_out[12], w_hssi_gen3_tx_pcs_tx_test_out[11], w_hssi_gen3_tx_pcs_tx_test_out[10], w_hssi_gen3_tx_pcs_tx_test_out[9], w_hssi_gen3_tx_pcs_tx_test_out[8], w_hssi_gen3_tx_pcs_tx_test_out[7], w_hssi_gen3_tx_pcs_tx_test_out[6], w_hssi_gen3_tx_pcs_tx_test_out[5], w_hssi_gen3_tx_pcs_tx_test_out[4], w_hssi_gen3_tx_pcs_tx_test_out[3], w_hssi_gen3_tx_pcs_tx_test_out[2], w_hssi_gen3_tx_pcs_tx_test_out[1], w_hssi_gen3_tx_pcs_tx_test_out[0]}),
				.txcompliance(w_hssi_8g_tx_pcs_txcompliance_out),
				.txdata({w_hssi_8g_tx_pcs_tx_data_out[31], w_hssi_8g_tx_pcs_tx_data_out[30], w_hssi_8g_tx_pcs_tx_data_out[29], w_hssi_8g_tx_pcs_tx_data_out[28], w_hssi_8g_tx_pcs_tx_data_out[27], w_hssi_8g_tx_pcs_tx_data_out[26], w_hssi_8g_tx_pcs_tx_data_out[25], w_hssi_8g_tx_pcs_tx_data_out[24], w_hssi_8g_tx_pcs_tx_data_out[23], w_hssi_8g_tx_pcs_tx_data_out[22], w_hssi_8g_tx_pcs_tx_data_out[21], w_hssi_8g_tx_pcs_tx_data_out[20], w_hssi_8g_tx_pcs_tx_data_out[19], w_hssi_8g_tx_pcs_tx_data_out[18], w_hssi_8g_tx_pcs_tx_data_out[17], w_hssi_8g_tx_pcs_tx_data_out[16], w_hssi_8g_tx_pcs_tx_data_out[15], w_hssi_8g_tx_pcs_tx_data_out[14], w_hssi_8g_tx_pcs_tx_data_out[13], w_hssi_8g_tx_pcs_tx_data_out[12], w_hssi_8g_tx_pcs_tx_data_out[11], w_hssi_8g_tx_pcs_tx_data_out[10], w_hssi_8g_tx_pcs_tx_data_out[9], w_hssi_8g_tx_pcs_tx_data_out[8], w_hssi_8g_tx_pcs_tx_data_out[7], w_hssi_8g_tx_pcs_tx_data_out[6], w_hssi_8g_tx_pcs_tx_data_out[5], w_hssi_8g_tx_pcs_tx_data_out[4], w_hssi_8g_tx_pcs_tx_data_out[3], w_hssi_8g_tx_pcs_tx_data_out[2], w_hssi_8g_tx_pcs_tx_data_out[1], w_hssi_8g_tx_pcs_tx_data_out[0]}),
				.txdatak({w_hssi_8g_tx_pcs_tx_datak_out[3], w_hssi_8g_tx_pcs_tx_datak_out[2], w_hssi_8g_tx_pcs_tx_datak_out[1], w_hssi_8g_tx_pcs_tx_datak_out[0]}),
				.txdataskip(w_hssi_8g_tx_pcs_tx_data_valid_out[0]),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_8g_tx_pcs_txelecidle_out),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.dis_pc_byte(),
				.pma_rx_det_pd(),
				.pma_txdeemph(),
				.pma_txmargin(),
				.pma_txswing(),
				.reset_pc_prts()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen3_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen3_blockselect = 1'b0;
				assign w_hssi_pipe_gen3_gen3_clk_sel = 1'b0;
				assign w_hssi_pipe_gen3_pcs_rst = 1'b0;
				assign w_hssi_pipe_gen3_phystatus = 1'b0;
				assign w_hssi_pipe_gen3_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen3_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_pma_tx_elec_idle = 1'b0;
				assign w_hssi_pipe_gen3_pma_txdetectrx = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_int = 1'b0;
				assign w_hssi_pipe_gen3_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_rxd_8gpcs_out[63:0] = 64'b0;
				assign w_hssi_pipe_gen3_rxdataskip[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_int = 1'b0;
				assign w_hssi_pipe_gen3_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_rxvalid = 1'b0;
				assign w_hssi_pipe_gen3_shutdown_clk = 1'b0;
				assign w_hssi_pipe_gen3_test_out[19:0] = 20'b0;
				assign w_hssi_pipe_gen3_tx_blk_start_int = 1'b0;
				assign w_hssi_pipe_gen3_tx_sync_hdr_int[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_txdata_int[31:0] = 32'b0;
				assign w_hssi_pipe_gen3_txdatak_int[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_txdataskip_int = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pcs_pma_interface
			twentynm_hssi_rx_pcs_pma_interface #(
				.block_sel(hssi_rx_pcs_pma_interface_block_sel),
				.channel_operation_mode(hssi_rx_pcs_pma_interface_channel_operation_mode),
				.clkslip_sel(hssi_rx_pcs_pma_interface_clkslip_sel),
				.lpbk_en(hssi_rx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_rx_pcs_pma_interface_master_clk_sel),
				.pldif_datawidth_mode(hssi_rx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_rx(hssi_rx_pcs_pma_interface_pma_dw_rx),
				.pma_if_dft_en(hssi_rx_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_rx_pcs_pma_interface_pma_if_dft_val),
				.prbs9_dwidth(hssi_rx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_rx_pcs_pma_interface_prbs_clken),
				.prbs_ver(hssi_rx_pcs_pma_interface_prbs_ver),
				.prot_mode_rx(hssi_rx_pcs_pma_interface_prot_mode_rx),
				.reconfig_settings(hssi_rx_pcs_pma_interface_reconfig_settings),
				.rx_dyn_polarity_inversion(hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion),
				.rx_lpbk_en(hssi_rx_pcs_pma_interface_rx_lpbk_en),
				.rx_prbs_force_signal_ok(hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok),
				.rx_prbs_mask(hssi_rx_pcs_pma_interface_rx_prbs_mask),
				.rx_prbs_mode(hssi_rx_pcs_pma_interface_rx_prbs_mode),
				.rx_signalok_signaldet_sel(hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel),
				.rx_static_polarity_inversion(hssi_rx_pcs_pma_interface_rx_static_polarity_inversion),
				.rx_uhsif_lpbk_en(hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sup_mode(hssi_rx_pcs_pma_interface_sup_mode)
			) inst_twentynm_hssi_rx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.int_pmaif_10g_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data),
				.int_pmaif_10g_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.int_pmaif_8g_pudi(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi),
				.int_pmaif_8g_rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.int_pmaif_8g_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.int_pmaif_8g_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.int_pmaif_8g_sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.int_pmaif_g3_pma_data_in(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in),
				.int_pmaif_g3_pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.int_pmaif_g3_pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.int_pmaif_g3_pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.int_pmaif_krfec_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data),
				.int_pmaif_krfec_rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.int_pmaif_pldif_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pmaif_pldif_prbs_err_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pmaif_pldif_rx_clkdiv(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pmaif_pldif_rx_clkdiv_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pmaif_pldif_rx_data(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data),
				.int_pmaif_pldif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pmaif_pldif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pmaif_pldif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pmaif_pldif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.pma_eye_monitor(w_hssi_rx_pcs_pma_interface_pma_eye_monitor),
				.pma_rx_clkslip(w_hssi_rx_pcs_pma_interface_pma_rx_clkslip),
				.pma_rxpma_rstb(w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb),
				.rx_pmaif_test_out(w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out),
				.rx_prbs_ver_test(w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.int_pmaif_8g_rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.int_pmaif_pldif_eye_monitor({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0]}),
				.int_pmaif_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pmaif_pldif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pmaif_pldif_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pmaif_pldif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pma_rx_clkdiv_user(in_pma_rx_clkdiv_user),
				.pma_rx_detect_valid(in_pma_rx_detect_valid),
				.pma_rx_found(in_pma_rx_found),
				.pma_rx_pma_clk(in_pma_rx_pma_clk),
				.pma_rx_pma_data({in_pma_rx_pma_data[63], in_pma_rx_pma_data[62], in_pma_rx_pma_data[61], in_pma_rx_pma_data[60], in_pma_rx_pma_data[59], in_pma_rx_pma_data[58], in_pma_rx_pma_data[57], in_pma_rx_pma_data[56], in_pma_rx_pma_data[55], in_pma_rx_pma_data[54], in_pma_rx_pma_data[53], in_pma_rx_pma_data[52], in_pma_rx_pma_data[51], in_pma_rx_pma_data[50], in_pma_rx_pma_data[49], in_pma_rx_pma_data[48], in_pma_rx_pma_data[47], in_pma_rx_pma_data[46], in_pma_rx_pma_data[45], in_pma_rx_pma_data[44], in_pma_rx_pma_data[43], in_pma_rx_pma_data[42], in_pma_rx_pma_data[41], in_pma_rx_pma_data[40], in_pma_rx_pma_data[39], in_pma_rx_pma_data[38], in_pma_rx_pma_data[37], in_pma_rx_pma_data[36], in_pma_rx_pma_data[35], in_pma_rx_pma_data[34], in_pma_rx_pma_data[33], in_pma_rx_pma_data[32], in_pma_rx_pma_data[31], in_pma_rx_pma_data[30], in_pma_rx_pma_data[29], in_pma_rx_pma_data[28], in_pma_rx_pma_data[27], in_pma_rx_pma_data[26], in_pma_rx_pma_data[25], in_pma_rx_pma_data[24], in_pma_rx_pma_data[23], in_pma_rx_pma_data[22], in_pma_rx_pma_data[21], in_pma_rx_pma_data[20], in_pma_rx_pma_data[19], in_pma_rx_pma_data[18], in_pma_rx_pma_data[17], in_pma_rx_pma_data[16], in_pma_rx_pma_data[15], in_pma_rx_pma_data[14], in_pma_rx_pma_data[13], in_pma_rx_pma_data[12], in_pma_rx_pma_data[11], in_pma_rx_pma_data[10], in_pma_rx_pma_data[9], in_pma_rx_pma_data[8], in_pma_rx_pma_data[7], in_pma_rx_pma_data[6], in_pma_rx_pma_data[5], in_pma_rx_pma_data[4], in_pma_rx_pma_data[3], in_pma_rx_pma_data[2], in_pma_rx_pma_data[1], in_pma_rx_pma_data[0]}),
				.pma_rx_signal_ok(in_pma_rx_signal_ok),
				.pma_rxpll_lock(in_pma_rxpll_lock),
				.pma_signal_det(in_pma_signal_det),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.tx_pma_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0]}),
				.tx_pma_uhsif_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0]}),
				
				// UNUSED
				.int_pmaif_g3_rcvd_clk(),
				.prbs_err_lt()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31:0] = 32'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5:0] = 6'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rx_clkslip = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pld_pcs_interface
			twentynm_hssi_rx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx),
				.hd_10g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx),
				.hd_10g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx),
				.hd_10g_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx),
				.hd_10g_lpbk_en(hssi_rx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx),
				.hd_10g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx),
				.hd_10g_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx),
				.hd_10g_test_bus_mode(hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode),
				.hd_8g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx),
				.hd_8g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx),
				.hd_8g_hip_mode(hssi_rx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_rx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx),
				.hd_8g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx),
				.hd_chnl_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_clklow_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz),
				.hd_chnl_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx),
				.hd_chnl_fref_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz),
				.hd_chnl_frequency_rules_en(hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_rx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_rx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx),
				.hd_chnl_lpbk_en(hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx),
				.hd_chnl_pld_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz),
				.hd_chnl_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx),
				.hd_chnl_pma_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz),
				.hd_chnl_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx),
				.hd_chnl_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx),
				.hd_chnl_transparent_pcs_rx(hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx),
				.hd_fifo_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx),
				.hd_fifo_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx),
				.hd_g3_prot_mode(hssi_rx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx),
				.hd_krfec_lpbk_en(hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx),
				.hd_krfec_test_bus_mode(hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode),
				.hd_pldif_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx),
				.hd_pmaif_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_lpbk_en(hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx),
				.hd_pmaif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx),
				.hd_pmaif_sim_mode(hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_rx_block_sel(hssi_rx_pld_pcs_interface_pcs_rx_block_sel),
				.pcs_rx_clk_out_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel),
				.pcs_rx_clk_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_sel),
				.pcs_rx_hip_clk_en(hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en),
				.pcs_rx_output_sel(hssi_rx_pld_pcs_interface_pcs_rx_output_sel),
				.reconfig_settings(hssi_rx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm5es2" )       //PARAM_HIDE
			) inst_twentynm_hssi_rx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pld_pcs_interface_blockselect),
				.hip_rx_ctrl(w_hssi_rx_pld_pcs_interface_hip_rx_ctrl),
				.hip_rx_data(w_hssi_rx_pld_pcs_interface_hip_rx_data),
				.int_pldif_10g_rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.int_pldif_10g_rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.int_pldif_10g_rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.int_pldif_10g_rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.int_pldif_10g_rx_control_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb),
				.int_pldif_10g_rx_data_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb),
				.int_pldif_10g_rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.int_pldif_10g_rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.int_pldif_10g_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.int_pldif_10g_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.int_pldif_10g_rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.int_pldif_8g_a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.int_pldif_8g_bitloc_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.int_pldif_8g_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.int_pldif_8g_byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.int_pldif_8g_encdt(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.int_pldif_8g_pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.int_pldif_8g_rdenable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.int_pldif_8g_rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.int_pldif_8g_rxurstpcs_n(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.int_pldif_8g_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.int_pldif_8g_wrdisable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.int_pldif_g3_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.int_pldif_krfec_rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.int_pldif_pmaif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pldif_pmaif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pldif_pmaif_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pldif_pmaif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pld_10g_krfec_rx_blk_lock(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock),
				.pld_10g_krfec_rx_diag_data_status(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status),
				.pld_10g_krfec_rx_frame(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame),
				.pld_10g_rx_align_val(w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val),
				.pld_10g_rx_crc32_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err),
				.pld_10g_rx_data_valid(w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid),
				.pld_10g_rx_empty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty),
				.pld_10g_rx_fifo_del(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del),
				.pld_10g_rx_fifo_insert(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert),
				.pld_10g_rx_fifo_num(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num),
				.pld_10g_rx_frame_lock(w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock),
				.pld_10g_rx_hi_ber(w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber),
				.pld_10g_rx_oflw_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err),
				.pld_10g_rx_pempty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty),
				.pld_10g_rx_pfull(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull),
				.pld_8g_a1a2_k1k2_flag(w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag),
				.pld_8g_empty_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf),
				.pld_8g_empty_rx(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx),
				.pld_8g_full_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf),
				.pld_8g_full_rx(w_hssi_rx_pld_pcs_interface_pld_8g_full_rx),
				.pld_8g_rxelecidle(w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle),
				.pld_8g_signal_detect_out(w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out),
				.pld_8g_wa_boundary(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary),
				.pld_pcs_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out),
				.pld_pma_clkdiv_rx_user(w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user),
				.pld_pma_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out),
				.pld_pma_signal_ok(w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok),
				.pld_rx_control(w_hssi_rx_pld_pcs_interface_pld_rx_control),
				.pld_rx_data(w_hssi_rx_pld_pcs_interface_pld_rx_data),
				.pld_rx_prbs_done(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done),
				.pld_rx_prbs_err(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.int_pldif_10g_rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.int_pldif_10g_rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.int_pldif_10g_rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_10g_rx_control({w_hssi_10g_rx_pcs_rx_control[19], w_hssi_10g_rx_pcs_rx_control[18], w_hssi_10g_rx_pcs_rx_control[17], w_hssi_10g_rx_pcs_rx_control[16], w_hssi_10g_rx_pcs_rx_control[15], w_hssi_10g_rx_pcs_rx_control[14], w_hssi_10g_rx_pcs_rx_control[13], w_hssi_10g_rx_pcs_rx_control[12], w_hssi_10g_rx_pcs_rx_control[11], w_hssi_10g_rx_pcs_rx_control[10], w_hssi_10g_rx_pcs_rx_control[9], w_hssi_10g_rx_pcs_rx_control[8], w_hssi_10g_rx_pcs_rx_control[7], w_hssi_10g_rx_pcs_rx_control[6], w_hssi_10g_rx_pcs_rx_control[5], w_hssi_10g_rx_pcs_rx_control[4], w_hssi_10g_rx_pcs_rx_control[3], w_hssi_10g_rx_pcs_rx_control[2], w_hssi_10g_rx_pcs_rx_control[1], w_hssi_10g_rx_pcs_rx_control[0]}),
				.int_pldif_10g_rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.int_pldif_10g_rx_data({w_hssi_10g_rx_pcs_rx_data[127], w_hssi_10g_rx_pcs_rx_data[126], w_hssi_10g_rx_pcs_rx_data[125], w_hssi_10g_rx_pcs_rx_data[124], w_hssi_10g_rx_pcs_rx_data[123], w_hssi_10g_rx_pcs_rx_data[122], w_hssi_10g_rx_pcs_rx_data[121], w_hssi_10g_rx_pcs_rx_data[120], w_hssi_10g_rx_pcs_rx_data[119], w_hssi_10g_rx_pcs_rx_data[118], w_hssi_10g_rx_pcs_rx_data[117], w_hssi_10g_rx_pcs_rx_data[116], w_hssi_10g_rx_pcs_rx_data[115], w_hssi_10g_rx_pcs_rx_data[114], w_hssi_10g_rx_pcs_rx_data[113], w_hssi_10g_rx_pcs_rx_data[112], w_hssi_10g_rx_pcs_rx_data[111], w_hssi_10g_rx_pcs_rx_data[110], w_hssi_10g_rx_pcs_rx_data[109], w_hssi_10g_rx_pcs_rx_data[108], w_hssi_10g_rx_pcs_rx_data[107], w_hssi_10g_rx_pcs_rx_data[106], w_hssi_10g_rx_pcs_rx_data[105], w_hssi_10g_rx_pcs_rx_data[104], w_hssi_10g_rx_pcs_rx_data[103], w_hssi_10g_rx_pcs_rx_data[102], w_hssi_10g_rx_pcs_rx_data[101], w_hssi_10g_rx_pcs_rx_data[100], w_hssi_10g_rx_pcs_rx_data[99], w_hssi_10g_rx_pcs_rx_data[98], w_hssi_10g_rx_pcs_rx_data[97], w_hssi_10g_rx_pcs_rx_data[96], w_hssi_10g_rx_pcs_rx_data[95], w_hssi_10g_rx_pcs_rx_data[94], w_hssi_10g_rx_pcs_rx_data[93], w_hssi_10g_rx_pcs_rx_data[92], w_hssi_10g_rx_pcs_rx_data[91], w_hssi_10g_rx_pcs_rx_data[90], w_hssi_10g_rx_pcs_rx_data[89], w_hssi_10g_rx_pcs_rx_data[88], w_hssi_10g_rx_pcs_rx_data[87], w_hssi_10g_rx_pcs_rx_data[86], w_hssi_10g_rx_pcs_rx_data[85], w_hssi_10g_rx_pcs_rx_data[84], w_hssi_10g_rx_pcs_rx_data[83], w_hssi_10g_rx_pcs_rx_data[82], w_hssi_10g_rx_pcs_rx_data[81], w_hssi_10g_rx_pcs_rx_data[80], w_hssi_10g_rx_pcs_rx_data[79], w_hssi_10g_rx_pcs_rx_data[78], w_hssi_10g_rx_pcs_rx_data[77], w_hssi_10g_rx_pcs_rx_data[76], w_hssi_10g_rx_pcs_rx_data[75], w_hssi_10g_rx_pcs_rx_data[74], w_hssi_10g_rx_pcs_rx_data[73], w_hssi_10g_rx_pcs_rx_data[72], w_hssi_10g_rx_pcs_rx_data[71], w_hssi_10g_rx_pcs_rx_data[70], w_hssi_10g_rx_pcs_rx_data[69], w_hssi_10g_rx_pcs_rx_data[68], w_hssi_10g_rx_pcs_rx_data[67], w_hssi_10g_rx_pcs_rx_data[66], w_hssi_10g_rx_pcs_rx_data[65], w_hssi_10g_rx_pcs_rx_data[64], w_hssi_10g_rx_pcs_rx_data[63], w_hssi_10g_rx_pcs_rx_data[62], w_hssi_10g_rx_pcs_rx_data[61], w_hssi_10g_rx_pcs_rx_data[60], w_hssi_10g_rx_pcs_rx_data[59], w_hssi_10g_rx_pcs_rx_data[58], w_hssi_10g_rx_pcs_rx_data[57], w_hssi_10g_rx_pcs_rx_data[56], w_hssi_10g_rx_pcs_rx_data[55], w_hssi_10g_rx_pcs_rx_data[54], w_hssi_10g_rx_pcs_rx_data[53], w_hssi_10g_rx_pcs_rx_data[52], w_hssi_10g_rx_pcs_rx_data[51], w_hssi_10g_rx_pcs_rx_data[50], w_hssi_10g_rx_pcs_rx_data[49], w_hssi_10g_rx_pcs_rx_data[48], w_hssi_10g_rx_pcs_rx_data[47], w_hssi_10g_rx_pcs_rx_data[46], w_hssi_10g_rx_pcs_rx_data[45], w_hssi_10g_rx_pcs_rx_data[44], w_hssi_10g_rx_pcs_rx_data[43], w_hssi_10g_rx_pcs_rx_data[42], w_hssi_10g_rx_pcs_rx_data[41], w_hssi_10g_rx_pcs_rx_data[40], w_hssi_10g_rx_pcs_rx_data[39], w_hssi_10g_rx_pcs_rx_data[38], w_hssi_10g_rx_pcs_rx_data[37], w_hssi_10g_rx_pcs_rx_data[36], w_hssi_10g_rx_pcs_rx_data[35], w_hssi_10g_rx_pcs_rx_data[34], w_hssi_10g_rx_pcs_rx_data[33], w_hssi_10g_rx_pcs_rx_data[32], w_hssi_10g_rx_pcs_rx_data[31], w_hssi_10g_rx_pcs_rx_data[30], w_hssi_10g_rx_pcs_rx_data[29], w_hssi_10g_rx_pcs_rx_data[28], w_hssi_10g_rx_pcs_rx_data[27], w_hssi_10g_rx_pcs_rx_data[26], w_hssi_10g_rx_pcs_rx_data[25], w_hssi_10g_rx_pcs_rx_data[24], w_hssi_10g_rx_pcs_rx_data[23], w_hssi_10g_rx_pcs_rx_data[22], w_hssi_10g_rx_pcs_rx_data[21], w_hssi_10g_rx_pcs_rx_data[20], w_hssi_10g_rx_pcs_rx_data[19], w_hssi_10g_rx_pcs_rx_data[18], w_hssi_10g_rx_pcs_rx_data[17], w_hssi_10g_rx_pcs_rx_data[16], w_hssi_10g_rx_pcs_rx_data[15], w_hssi_10g_rx_pcs_rx_data[14], w_hssi_10g_rx_pcs_rx_data[13], w_hssi_10g_rx_pcs_rx_data[12], w_hssi_10g_rx_pcs_rx_data[11], w_hssi_10g_rx_pcs_rx_data[10], w_hssi_10g_rx_pcs_rx_data[9], w_hssi_10g_rx_pcs_rx_data[8], w_hssi_10g_rx_pcs_rx_data[7], w_hssi_10g_rx_pcs_rx_data[6], w_hssi_10g_rx_pcs_rx_data[5], w_hssi_10g_rx_pcs_rx_data[4], w_hssi_10g_rx_pcs_rx_data[3], w_hssi_10g_rx_pcs_rx_data[2], w_hssi_10g_rx_pcs_rx_data[1], w_hssi_10g_rx_pcs_rx_data[0]}),
				.int_pldif_10g_rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.int_pldif_10g_rx_diag_status({w_hssi_10g_rx_pcs_rx_diag_status[1], w_hssi_10g_rx_pcs_rx_diag_status[0]}),
				.int_pldif_10g_rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.int_pldif_10g_rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.int_pldif_10g_rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.int_pldif_10g_rx_fifo_num({w_hssi_10g_rx_pcs_rx_fifo_num[4], w_hssi_10g_rx_pcs_rx_fifo_num[3], w_hssi_10g_rx_pcs_rx_fifo_num[2], w_hssi_10g_rx_pcs_rx_fifo_num[1], w_hssi_10g_rx_pcs_rx_fifo_num[0]}),
				.int_pldif_10g_rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.int_pldif_10g_rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.int_pldif_10g_rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.int_pldif_10g_rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.int_pldif_10g_rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.int_pldif_10g_rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				.int_pldif_8g_a1a2_k1k2_flag({w_hssi_8g_rx_pcs_a1a2k1k2flag[3], w_hssi_8g_rx_pcs_a1a2k1k2flag[2], w_hssi_8g_rx_pcs_a1a2k1k2flag[1], w_hssi_8g_rx_pcs_a1a2k1k2flag[0]}),
				.int_pldif_8g_empty_rmf(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.int_pldif_8g_empty_rx(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.int_pldif_8g_full_rmf(w_hssi_8g_rx_pcs_rm_fifo_full),
				.int_pldif_8g_full_rx(w_hssi_8g_rx_pcs_pcfifofull),
				.int_pldif_8g_phystatus(w_hssi_8g_rx_pcs_phystatus),
				.int_pldif_8g_rx_blk_start({w_hssi_8g_rx_pcs_rx_blk_start[3], w_hssi_8g_rx_pcs_rx_blk_start[2], w_hssi_8g_rx_pcs_rx_blk_start[1], w_hssi_8g_rx_pcs_rx_blk_start[0]}),
				.int_pldif_8g_rx_clk(w_hssi_8g_rx_pcs_clock_to_pld),
				.int_pldif_8g_rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_8g_rx_data_valid({w_hssi_8g_rx_pcs_rx_data_valid[3], w_hssi_8g_rx_pcs_rx_data_valid[2], w_hssi_8g_rx_pcs_rx_data_valid[1], w_hssi_8g_rx_pcs_rx_data_valid[0]}),
				.int_pldif_8g_rx_rstn_sync2wrfifo(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.int_pldif_8g_rx_sync_hdr({w_hssi_8g_rx_pcs_rx_sync_hdr[1], w_hssi_8g_rx_pcs_rx_sync_hdr[0]}),
				.int_pldif_8g_rxd({w_hssi_8g_rx_pcs_dataout[63], w_hssi_8g_rx_pcs_dataout[62], w_hssi_8g_rx_pcs_dataout[61], w_hssi_8g_rx_pcs_dataout[60], w_hssi_8g_rx_pcs_dataout[59], w_hssi_8g_rx_pcs_dataout[58], w_hssi_8g_rx_pcs_dataout[57], w_hssi_8g_rx_pcs_dataout[56], w_hssi_8g_rx_pcs_dataout[55], w_hssi_8g_rx_pcs_dataout[54], w_hssi_8g_rx_pcs_dataout[53], w_hssi_8g_rx_pcs_dataout[52], w_hssi_8g_rx_pcs_dataout[51], w_hssi_8g_rx_pcs_dataout[50], w_hssi_8g_rx_pcs_dataout[49], w_hssi_8g_rx_pcs_dataout[48], w_hssi_8g_rx_pcs_dataout[47], w_hssi_8g_rx_pcs_dataout[46], w_hssi_8g_rx_pcs_dataout[45], w_hssi_8g_rx_pcs_dataout[44], w_hssi_8g_rx_pcs_dataout[43], w_hssi_8g_rx_pcs_dataout[42], w_hssi_8g_rx_pcs_dataout[41], w_hssi_8g_rx_pcs_dataout[40], w_hssi_8g_rx_pcs_dataout[39], w_hssi_8g_rx_pcs_dataout[38], w_hssi_8g_rx_pcs_dataout[37], w_hssi_8g_rx_pcs_dataout[36], w_hssi_8g_rx_pcs_dataout[35], w_hssi_8g_rx_pcs_dataout[34], w_hssi_8g_rx_pcs_dataout[33], w_hssi_8g_rx_pcs_dataout[32], w_hssi_8g_rx_pcs_dataout[31], w_hssi_8g_rx_pcs_dataout[30], w_hssi_8g_rx_pcs_dataout[29], w_hssi_8g_rx_pcs_dataout[28], w_hssi_8g_rx_pcs_dataout[27], w_hssi_8g_rx_pcs_dataout[26], w_hssi_8g_rx_pcs_dataout[25], w_hssi_8g_rx_pcs_dataout[24], w_hssi_8g_rx_pcs_dataout[23], w_hssi_8g_rx_pcs_dataout[22], w_hssi_8g_rx_pcs_dataout[21], w_hssi_8g_rx_pcs_dataout[20], w_hssi_8g_rx_pcs_dataout[19], w_hssi_8g_rx_pcs_dataout[18], w_hssi_8g_rx_pcs_dataout[17], w_hssi_8g_rx_pcs_dataout[16], w_hssi_8g_rx_pcs_dataout[15], w_hssi_8g_rx_pcs_dataout[14], w_hssi_8g_rx_pcs_dataout[13], w_hssi_8g_rx_pcs_dataout[12], w_hssi_8g_rx_pcs_dataout[11], w_hssi_8g_rx_pcs_dataout[10], w_hssi_8g_rx_pcs_dataout[9], w_hssi_8g_rx_pcs_dataout[8], w_hssi_8g_rx_pcs_dataout[7], w_hssi_8g_rx_pcs_dataout[6], w_hssi_8g_rx_pcs_dataout[5], w_hssi_8g_rx_pcs_dataout[4], w_hssi_8g_rx_pcs_dataout[3], w_hssi_8g_rx_pcs_dataout[2], w_hssi_8g_rx_pcs_dataout[1], w_hssi_8g_rx_pcs_dataout[0]}),
				.int_pldif_8g_rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.int_pldif_8g_rxstatus({w_hssi_8g_rx_pcs_rxstatus[2], w_hssi_8g_rx_pcs_rxstatus[1], w_hssi_8g_rx_pcs_rxstatus[0]}),
				.int_pldif_8g_rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.int_pldif_8g_signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.int_pldif_8g_wa_boundary({w_hssi_8g_rx_pcs_word_align_boundary[4], w_hssi_8g_rx_pcs_word_align_boundary[3], w_hssi_8g_rx_pcs_word_align_boundary[2], w_hssi_8g_rx_pcs_word_align_boundary[1], w_hssi_8g_rx_pcs_word_align_boundary[0]}),
				.int_pldif_krfec_rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.int_pldif_krfec_rx_data_status({w_hssi_krfec_rx_pcs_rx_data_status[1], w_hssi_krfec_rx_pcs_rx_data_status[0]}),
				.int_pldif_krfec_rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.int_pldif_pmaif_clkdiv_rx(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pldif_pmaif_clkdiv_rx_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pldif_pmaif_rx_data({w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0]}),
				.int_pldif_pmaif_rx_prbs_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pldif_pmaif_rx_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.pld_10g_krfec_rx_clr_errblk_cnt(in_pld_10g_krfec_rx_clr_errblk_cnt),
				.pld_10g_krfec_rx_pld_rst_n(in_pld_10g_krfec_rx_pld_rst_n),
				.pld_10g_rx_align_clr(in_pld_10g_rx_align_clr),
				.pld_10g_rx_clr_ber_count(in_pld_10g_rx_clr_ber_count),
				.pld_10g_rx_rd_en(in_pld_10g_rx_rd_en),
				.pld_8g_a1a2_size(in_pld_8g_a1a2_size),
				.pld_8g_bitloc_rev_en(in_pld_8g_bitloc_rev_en),
				.pld_8g_byte_rev_en(in_pld_8g_byte_rev_en),
				.pld_8g_encdt(in_pld_8g_encdt),
				.pld_8g_g3_rx_pld_rst_n(in_pld_8g_g3_rx_pld_rst_n),
				.pld_8g_rdenable_rx(in_pld_8g_rdenable_rx),
				.pld_8g_rxpolarity(in_pld_8g_rxpolarity),
				.pld_8g_wrdisable_rx(in_pld_8g_wrdisable_rx),
				.pld_bitslip(in_pld_bitslip),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_rxpma_rstb(in_pld_pma_rxpma_rstb),
				.pld_pmaif_rx_pld_rst_n(in_pld_pmaif_rx_pld_rst_n),
				.pld_pmaif_rxclkslip(in_pld_pmaif_rxclkslip),
				.pld_polinv_rx(in_pld_polinv_rx),
				.pld_rx_clk(in_pld_rx_clk),
				.pld_rx_prbs_err_clr(in_pld_rx_prbs_err_clr),
				.pld_syncsm_en(in_pld_syncsm_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.int_pldif_pmaif_rx_pld_clk(),
				.pld_8g_wa_boundary_txclk_fastreg(),
				.pld_8g_wa_boundary_txclk_reg(),
				.pld_bitslip_10g_txclk_reg(),
				.pld_bitslip_8g_txclk_reg(),
				.pld_bitslip_rxclk_parallel_loopback_reg(),
				.pld_bitslip_rxclk_reg(),
				.pld_pcs_rx_clk_out_pcsdirect_wire(),
				.pld_pma_rx_clk_out_10g_or_pcsdirect_wire(),
				.pld_pma_rx_clk_out_8g_wire(),
				.pld_pmaif_rx_pld_rst_n_reg(),
				.pld_pmaif_tx_pld_rst_n_txclk_reg(),
				.pld_polinv_rx_reg(),
				.pld_rx_clk_fifo(),
				.pld_rx_control_fifo(),
				.pld_rx_control_pcsdirect_reg(),
				.pld_rx_data_fifo(),
				.pld_rx_data_pcsdirect_reg(),
				.pld_rx_prbs_done_reg(),
				.pld_rx_prbs_done_txclk_reg(),
				.pld_rx_prbs_err_clr_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_clr_reg(),
				.pld_rx_prbs_err_disprbs_reg(),
				.pld_rx_prbs_err_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_reg(),
				.pma_rx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_data[50:0] = 51'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3:0] = 4'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_control[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_data[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pcs_pma_interface
			twentynm_hssi_tx_pcs_pma_interface #(
				.bypass_pma_txelecidle(hssi_tx_pcs_pma_interface_bypass_pma_txelecidle),
				.channel_operation_mode(hssi_tx_pcs_pma_interface_channel_operation_mode),
				.lpbk_en(hssi_tx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_tx_pcs_pma_interface_master_clk_sel),
				.pcie_sub_prot_mode_tx(hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx),
				.pldif_datawidth_mode(hssi_tx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_tx(hssi_tx_pcs_pma_interface_pma_dw_tx),
				.pma_if_dft_en(hssi_tx_pcs_pma_interface_pma_if_dft_en),
				.pmagate_en(hssi_tx_pcs_pma_interface_pmagate_en),
				.prbs9_dwidth(hssi_tx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_tx_pcs_pma_interface_prbs_clken),
				.prbs_gen_pat(hssi_tx_pcs_pma_interface_prbs_gen_pat),
				.prot_mode_tx(hssi_tx_pcs_pma_interface_prot_mode_tx),
				.reconfig_settings(hssi_tx_pcs_pma_interface_reconfig_settings),
				.silicon_rev( "20nm5es2" ),       //PARAM_HIDE
				.sq_wave_num(hssi_tx_pcs_pma_interface_sq_wave_num),
				.sqwgen_clken(hssi_tx_pcs_pma_interface_sqwgen_clken),
				.sup_mode(hssi_tx_pcs_pma_interface_sup_mode),
				.tx_dyn_polarity_inversion(hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion),
				.tx_pma_data_sel(hssi_tx_pcs_pma_interface_tx_pma_data_sel),
				.tx_static_polarity_inversion(hssi_tx_pcs_pma_interface_tx_static_polarity_inversion),
				.uhsif_cnt_step_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock),
				.uhsif_cnt_thresh_filt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value),
				.uhsif_cnt_thresh_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock),
				.uhsif_dcn_test_update_period(hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period),
				.uhsif_dcn_testmode_enable(hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable),
				.uhsif_dead_zone_count_thresh(hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh),
				.uhsif_dead_zone_detection_enable(hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable),
				.uhsif_dead_zone_obser_window(hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window),
				.uhsif_dead_zone_skip_size(hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size),
				.uhsif_delay_cell_index_sel(hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel),
				.uhsif_delay_cell_margin(hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin),
				.uhsif_delay_cell_static_index_value(hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value),
				.uhsif_dft_dead_zone_control(hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control),
				.uhsif_dft_up_filt_control(hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control),
				.uhsif_enable(hssi_tx_pcs_pma_interface_uhsif_enable),
				.uhsif_lock_det_segsz_after_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock),
				.uhsif_lock_det_segsz_before_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock),
				.uhsif_lock_det_thresh_cnt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value),
				.uhsif_lock_det_thresh_cnt_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value),
				.uhsif_lock_det_thresh_diff_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value),
				.uhsif_lock_det_thresh_diff_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value)
			) inst_twentynm_hssi_tx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.int_pmaif_8g_txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.int_pmaif_pldif_tx_clkdiv(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pmaif_pldif_tx_clkdiv_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pmaif_pldif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.int_pmaif_pldif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.int_tx_dft_obsrv_clk(w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk),
				.pma_tx_elec_idle(w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle),
				.pma_tx_pma_data(w_hssi_tx_pcs_pma_interface_pma_tx_pma_data),
				.pma_txpma_rstb(w_hssi_tx_pcs_pma_interface_pma_txpma_rstb),
				.tx_pma_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback),
				.tx_pma_uhsif_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback),
				.tx_prbs_gen_test(w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test),
				.uhsif_test_out_1(w_hssi_tx_pcs_pma_interface_uhsif_test_out_1),
				.uhsif_test_out_2(w_hssi_tx_pcs_pma_interface_uhsif_test_out_2),
				.uhsif_test_out_3(w_hssi_tx_pcs_pma_interface_uhsif_test_out_3),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.int_pmaif_10g_tx_pma_data({w_hssi_10g_tx_pcs_tx_pma_data[63], w_hssi_10g_tx_pcs_tx_pma_data[62], w_hssi_10g_tx_pcs_tx_pma_data[61], w_hssi_10g_tx_pcs_tx_pma_data[60], w_hssi_10g_tx_pcs_tx_pma_data[59], w_hssi_10g_tx_pcs_tx_pma_data[58], w_hssi_10g_tx_pcs_tx_pma_data[57], w_hssi_10g_tx_pcs_tx_pma_data[56], w_hssi_10g_tx_pcs_tx_pma_data[55], w_hssi_10g_tx_pcs_tx_pma_data[54], w_hssi_10g_tx_pcs_tx_pma_data[53], w_hssi_10g_tx_pcs_tx_pma_data[52], w_hssi_10g_tx_pcs_tx_pma_data[51], w_hssi_10g_tx_pcs_tx_pma_data[50], w_hssi_10g_tx_pcs_tx_pma_data[49], w_hssi_10g_tx_pcs_tx_pma_data[48], w_hssi_10g_tx_pcs_tx_pma_data[47], w_hssi_10g_tx_pcs_tx_pma_data[46], w_hssi_10g_tx_pcs_tx_pma_data[45], w_hssi_10g_tx_pcs_tx_pma_data[44], w_hssi_10g_tx_pcs_tx_pma_data[43], w_hssi_10g_tx_pcs_tx_pma_data[42], w_hssi_10g_tx_pcs_tx_pma_data[41], w_hssi_10g_tx_pcs_tx_pma_data[40], w_hssi_10g_tx_pcs_tx_pma_data[39], w_hssi_10g_tx_pcs_tx_pma_data[38], w_hssi_10g_tx_pcs_tx_pma_data[37], w_hssi_10g_tx_pcs_tx_pma_data[36], w_hssi_10g_tx_pcs_tx_pma_data[35], w_hssi_10g_tx_pcs_tx_pma_data[34], w_hssi_10g_tx_pcs_tx_pma_data[33], w_hssi_10g_tx_pcs_tx_pma_data[32], w_hssi_10g_tx_pcs_tx_pma_data[31], w_hssi_10g_tx_pcs_tx_pma_data[30], w_hssi_10g_tx_pcs_tx_pma_data[29], w_hssi_10g_tx_pcs_tx_pma_data[28], w_hssi_10g_tx_pcs_tx_pma_data[27], w_hssi_10g_tx_pcs_tx_pma_data[26], w_hssi_10g_tx_pcs_tx_pma_data[25], w_hssi_10g_tx_pcs_tx_pma_data[24], w_hssi_10g_tx_pcs_tx_pma_data[23], w_hssi_10g_tx_pcs_tx_pma_data[22], w_hssi_10g_tx_pcs_tx_pma_data[21], w_hssi_10g_tx_pcs_tx_pma_data[20], w_hssi_10g_tx_pcs_tx_pma_data[19], w_hssi_10g_tx_pcs_tx_pma_data[18], w_hssi_10g_tx_pcs_tx_pma_data[17], w_hssi_10g_tx_pcs_tx_pma_data[16], w_hssi_10g_tx_pcs_tx_pma_data[15], w_hssi_10g_tx_pcs_tx_pma_data[14], w_hssi_10g_tx_pcs_tx_pma_data[13], w_hssi_10g_tx_pcs_tx_pma_data[12], w_hssi_10g_tx_pcs_tx_pma_data[11], w_hssi_10g_tx_pcs_tx_pma_data[10], w_hssi_10g_tx_pcs_tx_pma_data[9], w_hssi_10g_tx_pcs_tx_pma_data[8], w_hssi_10g_tx_pcs_tx_pma_data[7], w_hssi_10g_tx_pcs_tx_pma_data[6], w_hssi_10g_tx_pcs_tx_pma_data[5], w_hssi_10g_tx_pcs_tx_pma_data[4], w_hssi_10g_tx_pcs_tx_pma_data[3], w_hssi_10g_tx_pcs_tx_pma_data[2], w_hssi_10g_tx_pcs_tx_pma_data[1], w_hssi_10g_tx_pcs_tx_pma_data[0]}),
				.int_pmaif_10g_tx_pma_data_gate_val({w_hssi_10g_tx_pcs_tx_pma_gating_val[63], w_hssi_10g_tx_pcs_tx_pma_gating_val[62], w_hssi_10g_tx_pcs_tx_pma_gating_val[61], w_hssi_10g_tx_pcs_tx_pma_gating_val[60], w_hssi_10g_tx_pcs_tx_pma_gating_val[59], w_hssi_10g_tx_pcs_tx_pma_gating_val[58], w_hssi_10g_tx_pcs_tx_pma_gating_val[57], w_hssi_10g_tx_pcs_tx_pma_gating_val[56], w_hssi_10g_tx_pcs_tx_pma_gating_val[55], w_hssi_10g_tx_pcs_tx_pma_gating_val[54], w_hssi_10g_tx_pcs_tx_pma_gating_val[53], w_hssi_10g_tx_pcs_tx_pma_gating_val[52], w_hssi_10g_tx_pcs_tx_pma_gating_val[51], w_hssi_10g_tx_pcs_tx_pma_gating_val[50], w_hssi_10g_tx_pcs_tx_pma_gating_val[49], w_hssi_10g_tx_pcs_tx_pma_gating_val[48], w_hssi_10g_tx_pcs_tx_pma_gating_val[47], w_hssi_10g_tx_pcs_tx_pma_gating_val[46], w_hssi_10g_tx_pcs_tx_pma_gating_val[45], w_hssi_10g_tx_pcs_tx_pma_gating_val[44], w_hssi_10g_tx_pcs_tx_pma_gating_val[43], w_hssi_10g_tx_pcs_tx_pma_gating_val[42], w_hssi_10g_tx_pcs_tx_pma_gating_val[41], w_hssi_10g_tx_pcs_tx_pma_gating_val[40], w_hssi_10g_tx_pcs_tx_pma_gating_val[39], w_hssi_10g_tx_pcs_tx_pma_gating_val[38], w_hssi_10g_tx_pcs_tx_pma_gating_val[37], w_hssi_10g_tx_pcs_tx_pma_gating_val[36], w_hssi_10g_tx_pcs_tx_pma_gating_val[35], w_hssi_10g_tx_pcs_tx_pma_gating_val[34], w_hssi_10g_tx_pcs_tx_pma_gating_val[33], w_hssi_10g_tx_pcs_tx_pma_gating_val[32], w_hssi_10g_tx_pcs_tx_pma_gating_val[31], w_hssi_10g_tx_pcs_tx_pma_gating_val[30], w_hssi_10g_tx_pcs_tx_pma_gating_val[29], w_hssi_10g_tx_pcs_tx_pma_gating_val[28], w_hssi_10g_tx_pcs_tx_pma_gating_val[27], w_hssi_10g_tx_pcs_tx_pma_gating_val[26], w_hssi_10g_tx_pcs_tx_pma_gating_val[25], w_hssi_10g_tx_pcs_tx_pma_gating_val[24], w_hssi_10g_tx_pcs_tx_pma_gating_val[23], w_hssi_10g_tx_pcs_tx_pma_gating_val[22], w_hssi_10g_tx_pcs_tx_pma_gating_val[21], w_hssi_10g_tx_pcs_tx_pma_gating_val[20], w_hssi_10g_tx_pcs_tx_pma_gating_val[19], w_hssi_10g_tx_pcs_tx_pma_gating_val[18], w_hssi_10g_tx_pcs_tx_pma_gating_val[17], w_hssi_10g_tx_pcs_tx_pma_gating_val[16], w_hssi_10g_tx_pcs_tx_pma_gating_val[15], w_hssi_10g_tx_pcs_tx_pma_gating_val[14], w_hssi_10g_tx_pcs_tx_pma_gating_val[13], w_hssi_10g_tx_pcs_tx_pma_gating_val[12], w_hssi_10g_tx_pcs_tx_pma_gating_val[11], w_hssi_10g_tx_pcs_tx_pma_gating_val[10], w_hssi_10g_tx_pcs_tx_pma_gating_val[9], w_hssi_10g_tx_pcs_tx_pma_gating_val[8], w_hssi_10g_tx_pcs_tx_pma_gating_val[7], w_hssi_10g_tx_pcs_tx_pma_gating_val[6], w_hssi_10g_tx_pcs_tx_pma_gating_val[5], w_hssi_10g_tx_pcs_tx_pma_gating_val[4], w_hssi_10g_tx_pcs_tx_pma_gating_val[3], w_hssi_10g_tx_pcs_tx_pma_gating_val[2], w_hssi_10g_tx_pcs_tx_pma_gating_val[1], w_hssi_10g_tx_pcs_tx_pma_gating_val[0]}),
				.int_pmaif_8g_pudr({w_hssi_8g_tx_pcs_dataout[19], w_hssi_8g_tx_pcs_dataout[18], w_hssi_8g_tx_pcs_dataout[17], w_hssi_8g_tx_pcs_dataout[16], w_hssi_8g_tx_pcs_dataout[15], w_hssi_8g_tx_pcs_dataout[14], w_hssi_8g_tx_pcs_dataout[13], w_hssi_8g_tx_pcs_dataout[12], w_hssi_8g_tx_pcs_dataout[11], w_hssi_8g_tx_pcs_dataout[10], w_hssi_8g_tx_pcs_dataout[9], w_hssi_8g_tx_pcs_dataout[8], w_hssi_8g_tx_pcs_dataout[7], w_hssi_8g_tx_pcs_dataout[6], w_hssi_8g_tx_pcs_dataout[5], w_hssi_8g_tx_pcs_dataout[4], w_hssi_8g_tx_pcs_dataout[3], w_hssi_8g_tx_pcs_dataout[2], w_hssi_8g_tx_pcs_dataout[1], w_hssi_8g_tx_pcs_dataout[0]}),
				.int_pmaif_8g_tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.int_pmaif_8g_tx_elec_idle(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_pma_data_out({w_hssi_gen3_tx_pcs_data_out[31], w_hssi_gen3_tx_pcs_data_out[30], w_hssi_gen3_tx_pcs_data_out[29], w_hssi_gen3_tx_pcs_data_out[28], w_hssi_gen3_tx_pcs_data_out[27], w_hssi_gen3_tx_pcs_data_out[26], w_hssi_gen3_tx_pcs_data_out[25], w_hssi_gen3_tx_pcs_data_out[24], w_hssi_gen3_tx_pcs_data_out[23], w_hssi_gen3_tx_pcs_data_out[22], w_hssi_gen3_tx_pcs_data_out[21], w_hssi_gen3_tx_pcs_data_out[20], w_hssi_gen3_tx_pcs_data_out[19], w_hssi_gen3_tx_pcs_data_out[18], w_hssi_gen3_tx_pcs_data_out[17], w_hssi_gen3_tx_pcs_data_out[16], w_hssi_gen3_tx_pcs_data_out[15], w_hssi_gen3_tx_pcs_data_out[14], w_hssi_gen3_tx_pcs_data_out[13], w_hssi_gen3_tx_pcs_data_out[12], w_hssi_gen3_tx_pcs_data_out[11], w_hssi_gen3_tx_pcs_data_out[10], w_hssi_gen3_tx_pcs_data_out[9], w_hssi_gen3_tx_pcs_data_out[8], w_hssi_gen3_tx_pcs_data_out[7], w_hssi_gen3_tx_pcs_data_out[6], w_hssi_gen3_tx_pcs_data_out[5], w_hssi_gen3_tx_pcs_data_out[4], w_hssi_gen3_tx_pcs_data_out[3], w_hssi_gen3_tx_pcs_data_out[2], w_hssi_gen3_tx_pcs_data_out[1], w_hssi_gen3_tx_pcs_data_out[0]}),
				.int_pmaif_g3_pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.int_pmaif_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pmaif_pldif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pmaif_pldif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0]}),
				.int_pmaif_pldif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pmaif_pldif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.int_pmaif_pldif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pmaif_pldif_uhsif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0]}),
				.pma_tx_clkdiv_user(in_pma_tx_clkdiv_user),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.refclk_dig_uhsif(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.uhsif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.uhsif_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				
				// UNUSED
				.avmm_user_dataout(),
				.write_en(),
				.write_en_ack()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4:0] = 5'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_txpma_rstb = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pld_pcs_interface
			twentynm_hssi_tx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx),
				.hd_10g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx),
				.hd_10g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx),
				.hd_10g_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx),
				.hd_10g_lpbk_en(hssi_tx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx),
				.hd_10g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx),
				.hd_10g_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx),
				.hd_8g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx),
				.hd_8g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx),
				.hd_8g_hip_mode(hssi_tx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_tx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx),
				.hd_8g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx),
				.hd_chnl_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx),
				.hd_chnl_frequency_rules_en(hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_tx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_tx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx),
				.hd_chnl_lpbk_en(hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx),
				.hd_chnl_pld_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz),
				.hd_chnl_pld_uhsif_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz),
				.hd_chnl_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx),
				.hd_chnl_pma_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz),
				.hd_chnl_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx),
				.hd_chnl_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx),
				.hd_fifo_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx),
				.hd_fifo_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx),
				.hd_g3_prot_mode(hssi_tx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx),
				.hd_krfec_lpbk_en(hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx),
				.hd_pldif_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx),
				.hd_pmaif_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_ctrl_plane_bonding(hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding),
				.hd_pmaif_lpbk_en(hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx),
				.hd_pmaif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx),
				.hd_pmaif_sim_mode(hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_tx_clk_out_sel(hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel),
				.pcs_tx_clk_source(hssi_tx_pld_pcs_interface_pcs_tx_clk_source),
				.pcs_tx_data_source(hssi_tx_pld_pcs_interface_pcs_tx_data_source),
				.pcs_tx_delay1_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en),
				.pcs_tx_delay1_clk_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel),
				.pcs_tx_delay1_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl),
				.pcs_tx_delay1_data_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel),
				.pcs_tx_delay2_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en),
				.pcs_tx_delay2_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl),
				.pcs_tx_output_sel(hssi_tx_pld_pcs_interface_pcs_tx_output_sel),
				.reconfig_settings(hssi_tx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm5es2" )       //PARAM_HIDE
			) inst_twentynm_hssi_tx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pld_pcs_interface_blockselect),
				.hip_tx_clk(w_hssi_tx_pld_pcs_interface_hip_tx_clk),
				.int_pldif_10g_tx_bitslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip),
				.int_pldif_10g_tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.int_pldif_10g_tx_control(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control),
				.int_pldif_10g_tx_control_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg),
				.int_pldif_10g_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data),
				.int_pldif_10g_tx_data_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg),
				.int_pldif_10g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.int_pldif_10g_tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.int_pldif_10g_tx_diag_status(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status),
				.int_pldif_10g_tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.int_pldif_10g_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.int_pldif_10g_tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				.int_pldif_8g_pld_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.int_pldif_8g_powerdown(w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown),
				.int_pldif_8g_rddisable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.int_pldif_8g_rev_loopbk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.int_pldif_8g_tx_blk_start(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start),
				.int_pldif_8g_tx_boundary_sel(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel),
				.int_pldif_8g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid),
				.int_pldif_8g_tx_sync_hdr(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr),
				.int_pldif_8g_txd(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd),
				.int_pldif_8g_txd_fast_reg(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg),
				.int_pldif_8g_txdeemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.int_pldif_8g_txdetectrxloopback(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.int_pldif_8g_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.int_pldif_8g_txmargin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin),
				.int_pldif_8g_txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.int_pldif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.int_pldif_8g_wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				.int_pldif_pmaif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pldif_pmaif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pldif_pmaif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data),
				.int_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pldif_pmaif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pldif_pmaif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pldif_pmaif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pldif_pmaif_uhsif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data),
				.pld_10g_krfec_tx_frame(w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame),
				.pld_10g_tx_burst_en_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe),
				.pld_10g_tx_empty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty),
				.pld_10g_tx_fifo_num(w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num),
				.pld_10g_tx_full(w_hssi_tx_pld_pcs_interface_pld_10g_tx_full),
				.pld_10g_tx_pempty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty),
				.pld_10g_tx_pfull(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull),
				.pld_10g_tx_wordslip_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe),
				.pld_8g_empty_tx(w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx),
				.pld_8g_full_tx(w_hssi_tx_pld_pcs_interface_pld_8g_full_tx),
				.pld_krfec_tx_alignment(w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment),
				.pld_pcs_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out),
				.pld_pma_clkdiv_tx_user(w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user),
				.pld_pma_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out),
				.pld_uhsif_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.hip_tx_data({in_hip_tx_data[63], in_hip_tx_data[62], in_hip_tx_data[61], in_hip_tx_data[60], in_hip_tx_data[59], in_hip_tx_data[58], in_hip_tx_data[57], in_hip_tx_data[56], in_hip_tx_data[55], in_hip_tx_data[54], in_hip_tx_data[53], in_hip_tx_data[52], in_hip_tx_data[51], in_hip_tx_data[50], in_hip_tx_data[49], in_hip_tx_data[48], in_hip_tx_data[47], in_hip_tx_data[46], in_hip_tx_data[45], in_hip_tx_data[44], in_hip_tx_data[43], in_hip_tx_data[42], in_hip_tx_data[41], in_hip_tx_data[40], in_hip_tx_data[39], in_hip_tx_data[38], in_hip_tx_data[37], in_hip_tx_data[36], in_hip_tx_data[35], in_hip_tx_data[34], in_hip_tx_data[33], in_hip_tx_data[32], in_hip_tx_data[31], in_hip_tx_data[30], in_hip_tx_data[29], in_hip_tx_data[28], in_hip_tx_data[27], in_hip_tx_data[26], in_hip_tx_data[25], in_hip_tx_data[24], in_hip_tx_data[23], in_hip_tx_data[22], in_hip_tx_data[21], in_hip_tx_data[20], in_hip_tx_data[19], in_hip_tx_data[18], in_hip_tx_data[17], in_hip_tx_data[16], in_hip_tx_data[15], in_hip_tx_data[14], in_hip_tx_data[13], in_hip_tx_data[12], in_hip_tx_data[11], in_hip_tx_data[10], in_hip_tx_data[9], in_hip_tx_data[8], in_hip_tx_data[7], in_hip_tx_data[6], in_hip_tx_data[5], in_hip_tx_data[4], in_hip_tx_data[3], in_hip_tx_data[2], in_hip_tx_data[1], in_hip_tx_data[0]}),
				.int_pldif_10g_tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.int_pldif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.int_pldif_10g_tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_10g_tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.int_pldif_10g_tx_fifo_num({w_hssi_10g_tx_pcs_tx_fifo_num[3], w_hssi_10g_tx_pcs_tx_fifo_num[2], w_hssi_10g_tx_pcs_tx_fifo_num[1], w_hssi_10g_tx_pcs_tx_fifo_num[0]}),
				.int_pldif_10g_tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.int_pldif_10g_tx_full(w_hssi_10g_tx_pcs_tx_full),
				.int_pldif_10g_tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.int_pldif_10g_tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.int_pldif_10g_tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				.int_pldif_8g_empty_tx(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.int_pldif_8g_full_tx(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.int_pldif_8g_tx_clk_out(w_hssi_8g_tx_pcs_clk_out),
				.int_pldif_8g_tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_krfec_tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.int_pldif_krfec_tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.int_pldif_pmaif_clkdiv_tx(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pldif_pmaif_clkdiv_tx_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pldif_pmaif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.pld_10g_krfec_tx_pld_rst_n(in_pld_10g_krfec_tx_pld_rst_n),
				.pld_10g_tx_bitslip({in_pld_10g_tx_bitslip[6], in_pld_10g_tx_bitslip[5], in_pld_10g_tx_bitslip[4], in_pld_10g_tx_bitslip[3], in_pld_10g_tx_bitslip[2], in_pld_10g_tx_bitslip[1], in_pld_10g_tx_bitslip[0]}),
				.pld_10g_tx_burst_en(in_pld_10g_tx_burst_en),
				.pld_10g_tx_data_valid(in_pld_10g_tx_data_valid),
				.pld_10g_tx_diag_status({in_pld_10g_tx_diag_status[1], in_pld_10g_tx_diag_status[0]}),
				.pld_10g_tx_wordslip(in_pld_10g_tx_wordslip),
				.pld_8g_g3_tx_pld_rst_n(in_pld_8g_g3_tx_pld_rst_n),
				.pld_8g_rddisable_tx(in_pld_8g_rddisable_tx),
				.pld_8g_tx_boundary_sel({in_pld_8g_tx_boundary_sel[4], in_pld_8g_tx_boundary_sel[3], in_pld_8g_tx_boundary_sel[2], in_pld_8g_tx_boundary_sel[1], in_pld_8g_tx_boundary_sel[0]}),
				.pld_8g_wrenable_tx(in_pld_8g_wrenable_tx),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_txpma_rstb(in_pld_pma_txpma_rstb),
				.pld_pmaif_tx_pld_rst_n(in_pld_pmaif_tx_pld_rst_n),
				.pld_polinv_tx(in_pld_polinv_tx),
				.pld_tx_clk(in_pld_tx_clk),
				.pld_tx_control({in_pld_tx_control[17], in_pld_tx_control[16], in_pld_tx_control[15], in_pld_tx_control[14], in_pld_tx_control[13], in_pld_tx_control[12], in_pld_tx_control[11], in_pld_tx_control[10], in_pld_tx_control[9], in_pld_tx_control[8], in_pld_tx_control[7], in_pld_tx_control[6], in_pld_tx_control[5], in_pld_tx_control[4], in_pld_tx_control[3], in_pld_tx_control[2], in_pld_tx_control[1], in_pld_tx_control[0]}),
				.pld_tx_data({in_pld_tx_data[127], in_pld_tx_data[126], in_pld_tx_data[125], in_pld_tx_data[124], in_pld_tx_data[123], in_pld_tx_data[122], in_pld_tx_data[121], in_pld_tx_data[120], in_pld_tx_data[119], in_pld_tx_data[118], in_pld_tx_data[117], in_pld_tx_data[116], in_pld_tx_data[115], in_pld_tx_data[114], in_pld_tx_data[113], in_pld_tx_data[112], in_pld_tx_data[111], in_pld_tx_data[110], in_pld_tx_data[109], in_pld_tx_data[108], in_pld_tx_data[107], in_pld_tx_data[106], in_pld_tx_data[105], in_pld_tx_data[104], in_pld_tx_data[103], in_pld_tx_data[102], in_pld_tx_data[101], in_pld_tx_data[100], in_pld_tx_data[99], in_pld_tx_data[98], in_pld_tx_data[97], in_pld_tx_data[96], in_pld_tx_data[95], in_pld_tx_data[94], in_pld_tx_data[93], in_pld_tx_data[92], in_pld_tx_data[91], in_pld_tx_data[90], in_pld_tx_data[89], in_pld_tx_data[88], in_pld_tx_data[87], in_pld_tx_data[86], in_pld_tx_data[85], in_pld_tx_data[84], in_pld_tx_data[83], in_pld_tx_data[82], in_pld_tx_data[81], in_pld_tx_data[80], in_pld_tx_data[79], in_pld_tx_data[78], in_pld_tx_data[77], in_pld_tx_data[76], in_pld_tx_data[75], in_pld_tx_data[74], in_pld_tx_data[73], in_pld_tx_data[72], in_pld_tx_data[71], in_pld_tx_data[70], in_pld_tx_data[69], in_pld_tx_data[68], in_pld_tx_data[67], in_pld_tx_data[66], in_pld_tx_data[65], in_pld_tx_data[64], in_pld_tx_data[63], in_pld_tx_data[62], in_pld_tx_data[61], in_pld_tx_data[60], in_pld_tx_data[59], in_pld_tx_data[58], in_pld_tx_data[57], in_pld_tx_data[56], in_pld_tx_data[55], in_pld_tx_data[54], in_pld_tx_data[53], in_pld_tx_data[52], in_pld_tx_data[51], in_pld_tx_data[50], in_pld_tx_data[49], in_pld_tx_data[48], in_pld_tx_data[47], in_pld_tx_data[46], in_pld_tx_data[45], in_pld_tx_data[44], in_pld_tx_data[43], in_pld_tx_data[42], in_pld_tx_data[41], in_pld_tx_data[40], in_pld_tx_data[39], in_pld_tx_data[38], in_pld_tx_data[37], in_pld_tx_data[36], in_pld_tx_data[35], in_pld_tx_data[34], in_pld_tx_data[33], in_pld_tx_data[32], in_pld_tx_data[31], in_pld_tx_data[30], in_pld_tx_data[29], in_pld_tx_data[28], in_pld_tx_data[27], in_pld_tx_data[26], in_pld_tx_data[25], in_pld_tx_data[24], in_pld_tx_data[23], in_pld_tx_data[22], in_pld_tx_data[21], in_pld_tx_data[20], in_pld_tx_data[19], in_pld_tx_data[18], in_pld_tx_data[17], in_pld_tx_data[16], in_pld_tx_data[15], in_pld_tx_data[14], in_pld_tx_data[13], in_pld_tx_data[12], in_pld_tx_data[11], in_pld_tx_data[10], in_pld_tx_data[9], in_pld_tx_data[8], in_pld_tx_data[7], in_pld_tx_data[6], in_pld_tx_data[5], in_pld_tx_data[4], in_pld_tx_data[3], in_pld_tx_data[2], in_pld_tx_data[1], in_pld_tx_data[0]}),
				.pld_txelecidle(in_pld_txelecidle),
				.pld_uhsif_tx_clk(in_pld_uhsif_tx_clk),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.hip_clk_out_div_by_2_wire(),
				.hip_clk_out_wire(),
				.int_pldif_pmaif_tx_pld_clk(),
				.pld_10g_tx_burst_en_exe_10g_fastreg(),
				.pld_10g_tx_burst_en_exe_plddirect_reg(),
				.pld_10g_tx_data_valid_2ff_delay1_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay3_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg(),
				.pld_10g_tx_data_valid_fastreg(),
				.pld_10g_tx_data_valid_plddirect_fastreg(),
				.pld_pcs_tx_clk_out_pma_wire(),
				.pld_pma_tx_clk_out_wire(),
				.pld_pmaif_tx_pld_rst_n_reg(),
				.pld_polinv_tx_10g_pcsdirect_reg(),
				.pld_polinv_tx_8g_reg(),
				.pld_polinv_tx_pat_reg(),
				.pld_tx_clk_fifo(),
				.pld_tx_control_fifo(),
				.pld_tx_control_hi_10g_reg(),
				.pld_tx_control_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_10g_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_8g_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_control_lo_plddirect_fastreg(),
				.pld_tx_control_lo_plddirect_reg(),
				.pld_tx_data_hi_reg(),
				.pld_tx_data_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_10g_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_8g_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_data_lo_plddirect_fastreg(),
				.pld_tx_data_lo_plddirect_reg(),
				.pld_uhsif_reg(),
				.pma_tx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_hip_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6:0] = 7'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17:0] = 18'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8:0] = 9'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127:0] = 128'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4:0] = 5'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2:0] = 3'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_full = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_full_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out = 1'b0;
		end // if not generate
		
		//output assignments
		assign out_avmmreaddata_hssi_10g_rx_pcs = {w_hssi_10g_rx_pcs_avmmreaddata[7], w_hssi_10g_rx_pcs_avmmreaddata[6], w_hssi_10g_rx_pcs_avmmreaddata[5], w_hssi_10g_rx_pcs_avmmreaddata[4], w_hssi_10g_rx_pcs_avmmreaddata[3], w_hssi_10g_rx_pcs_avmmreaddata[2], w_hssi_10g_rx_pcs_avmmreaddata[1], w_hssi_10g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_10g_tx_pcs = {w_hssi_10g_tx_pcs_avmmreaddata[7], w_hssi_10g_tx_pcs_avmmreaddata[6], w_hssi_10g_tx_pcs_avmmreaddata[5], w_hssi_10g_tx_pcs_avmmreaddata[4], w_hssi_10g_tx_pcs_avmmreaddata[3], w_hssi_10g_tx_pcs_avmmreaddata[2], w_hssi_10g_tx_pcs_avmmreaddata[1], w_hssi_10g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_rx_pcs = {w_hssi_8g_rx_pcs_avmmreaddata[7], w_hssi_8g_rx_pcs_avmmreaddata[6], w_hssi_8g_rx_pcs_avmmreaddata[5], w_hssi_8g_rx_pcs_avmmreaddata[4], w_hssi_8g_rx_pcs_avmmreaddata[3], w_hssi_8g_rx_pcs_avmmreaddata[2], w_hssi_8g_rx_pcs_avmmreaddata[1], w_hssi_8g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_tx_pcs = {w_hssi_8g_tx_pcs_avmmreaddata[7], w_hssi_8g_tx_pcs_avmmreaddata[6], w_hssi_8g_tx_pcs_avmmreaddata[5], w_hssi_8g_tx_pcs_avmmreaddata[4], w_hssi_8g_tx_pcs_avmmreaddata[3], w_hssi_8g_tx_pcs_avmmreaddata[2], w_hssi_8g_tx_pcs_avmmreaddata[1], w_hssi_8g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pcs_pma_interface = {w_hssi_common_pcs_pma_interface_avmmreaddata[7], w_hssi_common_pcs_pma_interface_avmmreaddata[6], w_hssi_common_pcs_pma_interface_avmmreaddata[5], w_hssi_common_pcs_pma_interface_avmmreaddata[4], w_hssi_common_pcs_pma_interface_avmmreaddata[3], w_hssi_common_pcs_pma_interface_avmmreaddata[2], w_hssi_common_pcs_pma_interface_avmmreaddata[1], w_hssi_common_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pld_pcs_interface = {w_hssi_common_pld_pcs_interface_avmmreaddata[7], w_hssi_common_pld_pcs_interface_avmmreaddata[6], w_hssi_common_pld_pcs_interface_avmmreaddata[5], w_hssi_common_pld_pcs_interface_avmmreaddata[4], w_hssi_common_pld_pcs_interface_avmmreaddata[3], w_hssi_common_pld_pcs_interface_avmmreaddata[2], w_hssi_common_pld_pcs_interface_avmmreaddata[1], w_hssi_common_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_rx_pcs = {w_hssi_fifo_rx_pcs_avmmreaddata[7], w_hssi_fifo_rx_pcs_avmmreaddata[6], w_hssi_fifo_rx_pcs_avmmreaddata[5], w_hssi_fifo_rx_pcs_avmmreaddata[4], w_hssi_fifo_rx_pcs_avmmreaddata[3], w_hssi_fifo_rx_pcs_avmmreaddata[2], w_hssi_fifo_rx_pcs_avmmreaddata[1], w_hssi_fifo_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_tx_pcs = {w_hssi_fifo_tx_pcs_avmmreaddata[7], w_hssi_fifo_tx_pcs_avmmreaddata[6], w_hssi_fifo_tx_pcs_avmmreaddata[5], w_hssi_fifo_tx_pcs_avmmreaddata[4], w_hssi_fifo_tx_pcs_avmmreaddata[3], w_hssi_fifo_tx_pcs_avmmreaddata[2], w_hssi_fifo_tx_pcs_avmmreaddata[1], w_hssi_fifo_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_rx_pcs = {w_hssi_gen3_rx_pcs_avmmreaddata[7], w_hssi_gen3_rx_pcs_avmmreaddata[6], w_hssi_gen3_rx_pcs_avmmreaddata[5], w_hssi_gen3_rx_pcs_avmmreaddata[4], w_hssi_gen3_rx_pcs_avmmreaddata[3], w_hssi_gen3_rx_pcs_avmmreaddata[2], w_hssi_gen3_rx_pcs_avmmreaddata[1], w_hssi_gen3_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_tx_pcs = {w_hssi_gen3_tx_pcs_avmmreaddata[7], w_hssi_gen3_tx_pcs_avmmreaddata[6], w_hssi_gen3_tx_pcs_avmmreaddata[5], w_hssi_gen3_tx_pcs_avmmreaddata[4], w_hssi_gen3_tx_pcs_avmmreaddata[3], w_hssi_gen3_tx_pcs_avmmreaddata[2], w_hssi_gen3_tx_pcs_avmmreaddata[1], w_hssi_gen3_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_rx_pcs = {w_hssi_krfec_rx_pcs_avmmreaddata[7], w_hssi_krfec_rx_pcs_avmmreaddata[6], w_hssi_krfec_rx_pcs_avmmreaddata[5], w_hssi_krfec_rx_pcs_avmmreaddata[4], w_hssi_krfec_rx_pcs_avmmreaddata[3], w_hssi_krfec_rx_pcs_avmmreaddata[2], w_hssi_krfec_rx_pcs_avmmreaddata[1], w_hssi_krfec_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_tx_pcs = {w_hssi_krfec_tx_pcs_avmmreaddata[7], w_hssi_krfec_tx_pcs_avmmreaddata[6], w_hssi_krfec_tx_pcs_avmmreaddata[5], w_hssi_krfec_tx_pcs_avmmreaddata[4], w_hssi_krfec_tx_pcs_avmmreaddata[3], w_hssi_krfec_tx_pcs_avmmreaddata[2], w_hssi_krfec_tx_pcs_avmmreaddata[1], w_hssi_krfec_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen1_2 = {w_hssi_pipe_gen1_2_avmmreaddata[7], w_hssi_pipe_gen1_2_avmmreaddata[6], w_hssi_pipe_gen1_2_avmmreaddata[5], w_hssi_pipe_gen1_2_avmmreaddata[4], w_hssi_pipe_gen1_2_avmmreaddata[3], w_hssi_pipe_gen1_2_avmmreaddata[2], w_hssi_pipe_gen1_2_avmmreaddata[1], w_hssi_pipe_gen1_2_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen3 = {w_hssi_pipe_gen3_avmmreaddata[7], w_hssi_pipe_gen3_avmmreaddata[6], w_hssi_pipe_gen3_avmmreaddata[5], w_hssi_pipe_gen3_avmmreaddata[4], w_hssi_pipe_gen3_avmmreaddata[3], w_hssi_pipe_gen3_avmmreaddata[2], w_hssi_pipe_gen3_avmmreaddata[1], w_hssi_pipe_gen3_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pcs_pma_interface = {w_hssi_rx_pcs_pma_interface_avmmreaddata[7], w_hssi_rx_pcs_pma_interface_avmmreaddata[6], w_hssi_rx_pcs_pma_interface_avmmreaddata[5], w_hssi_rx_pcs_pma_interface_avmmreaddata[4], w_hssi_rx_pcs_pma_interface_avmmreaddata[3], w_hssi_rx_pcs_pma_interface_avmmreaddata[2], w_hssi_rx_pcs_pma_interface_avmmreaddata[1], w_hssi_rx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pld_pcs_interface = {w_hssi_rx_pld_pcs_interface_avmmreaddata[7], w_hssi_rx_pld_pcs_interface_avmmreaddata[6], w_hssi_rx_pld_pcs_interface_avmmreaddata[5], w_hssi_rx_pld_pcs_interface_avmmreaddata[4], w_hssi_rx_pld_pcs_interface_avmmreaddata[3], w_hssi_rx_pld_pcs_interface_avmmreaddata[2], w_hssi_rx_pld_pcs_interface_avmmreaddata[1], w_hssi_rx_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pcs_pma_interface = {w_hssi_tx_pcs_pma_interface_avmmreaddata[7], w_hssi_tx_pcs_pma_interface_avmmreaddata[6], w_hssi_tx_pcs_pma_interface_avmmreaddata[5], w_hssi_tx_pcs_pma_interface_avmmreaddata[4], w_hssi_tx_pcs_pma_interface_avmmreaddata[3], w_hssi_tx_pcs_pma_interface_avmmreaddata[2], w_hssi_tx_pcs_pma_interface_avmmreaddata[1], w_hssi_tx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pld_pcs_interface = {w_hssi_tx_pld_pcs_interface_avmmreaddata[7], w_hssi_tx_pld_pcs_interface_avmmreaddata[6], w_hssi_tx_pld_pcs_interface_avmmreaddata[5], w_hssi_tx_pld_pcs_interface_avmmreaddata[4], w_hssi_tx_pld_pcs_interface_avmmreaddata[3], w_hssi_tx_pld_pcs_interface_avmmreaddata[2], w_hssi_tx_pld_pcs_interface_avmmreaddata[1], w_hssi_tx_pld_pcs_interface_avmmreaddata[0]};
		assign out_blockselect_hssi_10g_rx_pcs = w_hssi_10g_rx_pcs_blockselect;
		assign out_blockselect_hssi_10g_tx_pcs = w_hssi_10g_tx_pcs_blockselect;
		assign out_blockselect_hssi_8g_rx_pcs = w_hssi_8g_rx_pcs_blockselect;
		assign out_blockselect_hssi_8g_tx_pcs = w_hssi_8g_tx_pcs_blockselect;
		assign out_blockselect_hssi_common_pcs_pma_interface = w_hssi_common_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_common_pld_pcs_interface = w_hssi_common_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_fifo_rx_pcs = w_hssi_fifo_rx_pcs_blockselect;
		assign out_blockselect_hssi_fifo_tx_pcs = w_hssi_fifo_tx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_rx_pcs = w_hssi_gen3_rx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_tx_pcs = w_hssi_gen3_tx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_rx_pcs = w_hssi_krfec_rx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_tx_pcs = w_hssi_krfec_tx_pcs_blockselect;
		assign out_blockselect_hssi_pipe_gen1_2 = w_hssi_pipe_gen1_2_blockselect;
		assign out_blockselect_hssi_pipe_gen3 = w_hssi_pipe_gen3_blockselect;
		assign out_blockselect_hssi_rx_pcs_pma_interface = w_hssi_rx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_rx_pld_pcs_interface = w_hssi_rx_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_tx_pcs_pma_interface = w_hssi_tx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_tx_pld_pcs_interface = w_hssi_tx_pld_pcs_interface_blockselect;
		assign out_bond_pcs10g_out_bot = {w_hssi_10g_tx_pcs_distdwn_out_rden, w_hssi_10g_tx_pcs_distdwn_out_wren, w_hssi_10g_tx_pcs_distdwn_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs10g_out_top = {w_hssi_10g_tx_pcs_distup_out_rden, w_hssi_10g_tx_pcs_distup_out_wren, w_hssi_10g_tx_pcs_distup_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs8g_out_bot = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down, w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_down, w_hssi_8g_tx_pcs_wr_enable_out_chnl_down, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_down, w_hssi_8g_rx_pcs_wr_enable_out_chnl_down, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[0]};
		assign out_bond_pcs8g_out_top = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up, w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_up, w_hssi_8g_tx_pcs_wr_enable_out_chnl_up, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_up, w_hssi_8g_rx_pcs_wr_enable_out_chnl_up, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[0]};
		assign out_bond_pmaif_out_bot = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[0]};
		assign out_bond_pmaif_out_top = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[0]};
		assign out_hip_clk_out = {w_hssi_common_pld_pcs_interface_hip_cmn_clk[1], w_hssi_common_pld_pcs_interface_hip_cmn_clk[0], w_hssi_tx_pld_pcs_interface_hip_tx_clk};
		assign out_hip_ctrl_out = {w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[4], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[3], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[2], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[1], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[0], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[0]};
		assign out_hip_iocsr_rdy = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
		assign out_hip_iocsr_rdy_dly = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
		assign out_hip_nfrzdrv = w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
		assign out_hip_npor = w_hssi_common_pld_pcs_interface_hip_npor;
		assign out_hip_rx_data = {w_hssi_rx_pld_pcs_interface_hip_rx_data[50], w_hssi_rx_pld_pcs_interface_hip_rx_data[49], w_hssi_rx_pld_pcs_interface_hip_rx_data[48], w_hssi_rx_pld_pcs_interface_hip_rx_data[47], w_hssi_rx_pld_pcs_interface_hip_rx_data[46], w_hssi_rx_pld_pcs_interface_hip_rx_data[45], w_hssi_rx_pld_pcs_interface_hip_rx_data[44], w_hssi_rx_pld_pcs_interface_hip_rx_data[43], w_hssi_rx_pld_pcs_interface_hip_rx_data[42], w_hssi_rx_pld_pcs_interface_hip_rx_data[41], w_hssi_rx_pld_pcs_interface_hip_rx_data[40], w_hssi_rx_pld_pcs_interface_hip_rx_data[39], w_hssi_rx_pld_pcs_interface_hip_rx_data[38], w_hssi_rx_pld_pcs_interface_hip_rx_data[37], w_hssi_rx_pld_pcs_interface_hip_rx_data[36], w_hssi_rx_pld_pcs_interface_hip_rx_data[35], w_hssi_rx_pld_pcs_interface_hip_rx_data[34], w_hssi_rx_pld_pcs_interface_hip_rx_data[33], w_hssi_rx_pld_pcs_interface_hip_rx_data[32], w_hssi_rx_pld_pcs_interface_hip_rx_data[31], w_hssi_rx_pld_pcs_interface_hip_rx_data[30], w_hssi_rx_pld_pcs_interface_hip_rx_data[29], w_hssi_rx_pld_pcs_interface_hip_rx_data[28], w_hssi_rx_pld_pcs_interface_hip_rx_data[27], w_hssi_rx_pld_pcs_interface_hip_rx_data[26], w_hssi_rx_pld_pcs_interface_hip_rx_data[25], w_hssi_rx_pld_pcs_interface_hip_rx_data[24], w_hssi_rx_pld_pcs_interface_hip_rx_data[23], w_hssi_rx_pld_pcs_interface_hip_rx_data[22], w_hssi_rx_pld_pcs_interface_hip_rx_data[21], w_hssi_rx_pld_pcs_interface_hip_rx_data[20], w_hssi_rx_pld_pcs_interface_hip_rx_data[19], w_hssi_rx_pld_pcs_interface_hip_rx_data[18], w_hssi_rx_pld_pcs_interface_hip_rx_data[17], w_hssi_rx_pld_pcs_interface_hip_rx_data[16], w_hssi_rx_pld_pcs_interface_hip_rx_data[15], w_hssi_rx_pld_pcs_interface_hip_rx_data[14], w_hssi_rx_pld_pcs_interface_hip_rx_data[13], w_hssi_rx_pld_pcs_interface_hip_rx_data[12], w_hssi_rx_pld_pcs_interface_hip_rx_data[11], w_hssi_rx_pld_pcs_interface_hip_rx_data[10], w_hssi_rx_pld_pcs_interface_hip_rx_data[9], w_hssi_rx_pld_pcs_interface_hip_rx_data[8], w_hssi_rx_pld_pcs_interface_hip_rx_data[7], w_hssi_rx_pld_pcs_interface_hip_rx_data[6], w_hssi_rx_pld_pcs_interface_hip_rx_data[5], w_hssi_rx_pld_pcs_interface_hip_rx_data[4], w_hssi_rx_pld_pcs_interface_hip_rx_data[3], w_hssi_rx_pld_pcs_interface_hip_rx_data[2], w_hssi_rx_pld_pcs_interface_hip_rx_data[1], w_hssi_rx_pld_pcs_interface_hip_rx_data[0]};
		assign out_hip_usermode = w_hssi_common_pld_pcs_interface_hip_usermode;
		assign out_pld_10g_krfec_rx_blk_lock = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
		assign out_pld_10g_krfec_rx_diag_data_status = {w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1], w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[0]};
		assign out_pld_10g_krfec_rx_frame = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
		assign out_pld_10g_krfec_tx_frame = w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
		assign out_pld_10g_rx_align_val = w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
		assign out_pld_10g_rx_crc32_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
		assign out_pld_10g_rx_data_valid = w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
		assign out_pld_10g_rx_empty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
		assign out_pld_10g_rx_fifo_del = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
		assign out_pld_10g_rx_fifo_insert = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
		assign out_pld_10g_rx_fifo_num = {w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[3], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[2], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[1], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[0]};
		assign out_pld_10g_rx_frame_lock = w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
		assign out_pld_10g_rx_hi_ber = w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
		assign out_pld_10g_rx_oflw_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
		assign out_pld_10g_rx_pempty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
		assign out_pld_10g_rx_pfull = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
		assign out_pld_10g_tx_burst_en_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
		assign out_pld_10g_tx_empty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
		assign out_pld_10g_tx_fifo_num = {w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[2], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[1], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[0]};
		assign out_pld_10g_tx_full = w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
		assign out_pld_10g_tx_pempty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
		assign out_pld_10g_tx_pfull = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
		assign out_pld_10g_tx_wordslip_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
		assign out_pld_8g_a1a2_k1k2_flag = {w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[2], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[1], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[0]};
		assign out_pld_8g_empty_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
		assign out_pld_8g_empty_rx = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
		assign out_pld_8g_empty_tx = w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
		assign out_pld_8g_full_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
		assign out_pld_8g_full_rx = w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
		assign out_pld_8g_full_tx = w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
		assign out_pld_8g_rxelecidle = w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
		assign out_pld_8g_signal_detect_out = w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
		assign out_pld_8g_wa_boundary = {w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0]};
		assign out_pld_krfec_tx_alignment = w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
		assign out_pld_pcs_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
		assign out_pld_pcs_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
		assign out_pld_pma_adapt_done = w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
		assign out_pld_pma_clkdiv_rx_user = w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
		assign out_pld_pma_clkdiv_tx_user = w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
		assign out_pld_pma_clklow = w_hssi_common_pld_pcs_interface_pld_pma_clklow;
		assign out_pld_pma_fref = w_hssi_common_pld_pcs_interface_pld_pma_fref;
		assign out_pld_pma_hclk = w_hssi_common_pld_pcs_interface_pld_pma_hclk;
		assign out_pld_pma_pcie_sw_done = {w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1], w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[0]};
		assign out_pld_pma_pfdmode_lock = w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
		assign out_pld_pma_reserved_in = {w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[3], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[2], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[1], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[0]};
		assign out_pld_pma_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
		assign out_pld_pma_rx_detect_valid = w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
		assign out_pld_pma_rx_found = w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
		assign out_pld_pma_rxpll_lock = w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
		assign out_pld_pma_signal_ok = w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
		assign out_pld_pma_testbus = {w_hssi_common_pld_pcs_interface_pld_pma_testbus[7], w_hssi_common_pld_pcs_interface_pld_pma_testbus[6], w_hssi_common_pld_pcs_interface_pld_pma_testbus[5], w_hssi_common_pld_pcs_interface_pld_pma_testbus[4], w_hssi_common_pld_pcs_interface_pld_pma_testbus[3], w_hssi_common_pld_pcs_interface_pld_pma_testbus[2], w_hssi_common_pld_pcs_interface_pld_pma_testbus[1], w_hssi_common_pld_pcs_interface_pld_pma_testbus[0]};
		assign out_pld_pma_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
		assign out_pld_pmaif_mask_tx_pll = w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
		assign out_pld_reserved_out = {w_hssi_common_pld_pcs_interface_pld_reserved_out[9], w_hssi_common_pld_pcs_interface_pld_reserved_out[8], w_hssi_common_pld_pcs_interface_pld_reserved_out[7], w_hssi_common_pld_pcs_interface_pld_reserved_out[6], w_hssi_common_pld_pcs_interface_pld_reserved_out[5], w_hssi_common_pld_pcs_interface_pld_reserved_out[4], w_hssi_common_pld_pcs_interface_pld_reserved_out[3], w_hssi_common_pld_pcs_interface_pld_reserved_out[2], w_hssi_common_pld_pcs_interface_pld_reserved_out[1], w_hssi_common_pld_pcs_interface_pld_reserved_out[0]};
		assign out_pld_rx_control = {w_hssi_rx_pld_pcs_interface_pld_rx_control[19], w_hssi_rx_pld_pcs_interface_pld_rx_control[18], w_hssi_rx_pld_pcs_interface_pld_rx_control[17], w_hssi_rx_pld_pcs_interface_pld_rx_control[16], w_hssi_rx_pld_pcs_interface_pld_rx_control[15], w_hssi_rx_pld_pcs_interface_pld_rx_control[14], w_hssi_rx_pld_pcs_interface_pld_rx_control[13], w_hssi_rx_pld_pcs_interface_pld_rx_control[12], w_hssi_rx_pld_pcs_interface_pld_rx_control[11], w_hssi_rx_pld_pcs_interface_pld_rx_control[10], w_hssi_rx_pld_pcs_interface_pld_rx_control[9], w_hssi_rx_pld_pcs_interface_pld_rx_control[8], w_hssi_rx_pld_pcs_interface_pld_rx_control[7], w_hssi_rx_pld_pcs_interface_pld_rx_control[6], w_hssi_rx_pld_pcs_interface_pld_rx_control[5], w_hssi_rx_pld_pcs_interface_pld_rx_control[4], w_hssi_rx_pld_pcs_interface_pld_rx_control[3], w_hssi_rx_pld_pcs_interface_pld_rx_control[2], w_hssi_rx_pld_pcs_interface_pld_rx_control[1], w_hssi_rx_pld_pcs_interface_pld_rx_control[0]};
		assign out_pld_rx_data = {w_hssi_rx_pld_pcs_interface_pld_rx_data[127], w_hssi_rx_pld_pcs_interface_pld_rx_data[126], w_hssi_rx_pld_pcs_interface_pld_rx_data[125], w_hssi_rx_pld_pcs_interface_pld_rx_data[124], w_hssi_rx_pld_pcs_interface_pld_rx_data[123], w_hssi_rx_pld_pcs_interface_pld_rx_data[122], w_hssi_rx_pld_pcs_interface_pld_rx_data[121], w_hssi_rx_pld_pcs_interface_pld_rx_data[120], w_hssi_rx_pld_pcs_interface_pld_rx_data[119], w_hssi_rx_pld_pcs_interface_pld_rx_data[118], w_hssi_rx_pld_pcs_interface_pld_rx_data[117], w_hssi_rx_pld_pcs_interface_pld_rx_data[116], w_hssi_rx_pld_pcs_interface_pld_rx_data[115], w_hssi_rx_pld_pcs_interface_pld_rx_data[114], w_hssi_rx_pld_pcs_interface_pld_rx_data[113], w_hssi_rx_pld_pcs_interface_pld_rx_data[112], w_hssi_rx_pld_pcs_interface_pld_rx_data[111], w_hssi_rx_pld_pcs_interface_pld_rx_data[110], w_hssi_rx_pld_pcs_interface_pld_rx_data[109], w_hssi_rx_pld_pcs_interface_pld_rx_data[108], w_hssi_rx_pld_pcs_interface_pld_rx_data[107], w_hssi_rx_pld_pcs_interface_pld_rx_data[106], w_hssi_rx_pld_pcs_interface_pld_rx_data[105], w_hssi_rx_pld_pcs_interface_pld_rx_data[104], w_hssi_rx_pld_pcs_interface_pld_rx_data[103], w_hssi_rx_pld_pcs_interface_pld_rx_data[102], w_hssi_rx_pld_pcs_interface_pld_rx_data[101], w_hssi_rx_pld_pcs_interface_pld_rx_data[100], w_hssi_rx_pld_pcs_interface_pld_rx_data[99], w_hssi_rx_pld_pcs_interface_pld_rx_data[98], w_hssi_rx_pld_pcs_interface_pld_rx_data[97], w_hssi_rx_pld_pcs_interface_pld_rx_data[96], w_hssi_rx_pld_pcs_interface_pld_rx_data[95], w_hssi_rx_pld_pcs_interface_pld_rx_data[94], w_hssi_rx_pld_pcs_interface_pld_rx_data[93], w_hssi_rx_pld_pcs_interface_pld_rx_data[92], w_hssi_rx_pld_pcs_interface_pld_rx_data[91], w_hssi_rx_pld_pcs_interface_pld_rx_data[90], w_hssi_rx_pld_pcs_interface_pld_rx_data[89], w_hssi_rx_pld_pcs_interface_pld_rx_data[88], w_hssi_rx_pld_pcs_interface_pld_rx_data[87], w_hssi_rx_pld_pcs_interface_pld_rx_data[86], w_hssi_rx_pld_pcs_interface_pld_rx_data[85], w_hssi_rx_pld_pcs_interface_pld_rx_data[84], w_hssi_rx_pld_pcs_interface_pld_rx_data[83], w_hssi_rx_pld_pcs_interface_pld_rx_data[82], w_hssi_rx_pld_pcs_interface_pld_rx_data[81], w_hssi_rx_pld_pcs_interface_pld_rx_data[80], w_hssi_rx_pld_pcs_interface_pld_rx_data[79], w_hssi_rx_pld_pcs_interface_pld_rx_data[78], w_hssi_rx_pld_pcs_interface_pld_rx_data[77], w_hssi_rx_pld_pcs_interface_pld_rx_data[76], w_hssi_rx_pld_pcs_interface_pld_rx_data[75], w_hssi_rx_pld_pcs_interface_pld_rx_data[74], w_hssi_rx_pld_pcs_interface_pld_rx_data[73], w_hssi_rx_pld_pcs_interface_pld_rx_data[72], w_hssi_rx_pld_pcs_interface_pld_rx_data[71], w_hssi_rx_pld_pcs_interface_pld_rx_data[70], w_hssi_rx_pld_pcs_interface_pld_rx_data[69], w_hssi_rx_pld_pcs_interface_pld_rx_data[68], w_hssi_rx_pld_pcs_interface_pld_rx_data[67], w_hssi_rx_pld_pcs_interface_pld_rx_data[66], w_hssi_rx_pld_pcs_interface_pld_rx_data[65], w_hssi_rx_pld_pcs_interface_pld_rx_data[64], w_hssi_rx_pld_pcs_interface_pld_rx_data[63], w_hssi_rx_pld_pcs_interface_pld_rx_data[62], w_hssi_rx_pld_pcs_interface_pld_rx_data[61], w_hssi_rx_pld_pcs_interface_pld_rx_data[60], w_hssi_rx_pld_pcs_interface_pld_rx_data[59], w_hssi_rx_pld_pcs_interface_pld_rx_data[58], w_hssi_rx_pld_pcs_interface_pld_rx_data[57], w_hssi_rx_pld_pcs_interface_pld_rx_data[56], w_hssi_rx_pld_pcs_interface_pld_rx_data[55], w_hssi_rx_pld_pcs_interface_pld_rx_data[54], w_hssi_rx_pld_pcs_interface_pld_rx_data[53], w_hssi_rx_pld_pcs_interface_pld_rx_data[52], w_hssi_rx_pld_pcs_interface_pld_rx_data[51], w_hssi_rx_pld_pcs_interface_pld_rx_data[50], w_hssi_rx_pld_pcs_interface_pld_rx_data[49], w_hssi_rx_pld_pcs_interface_pld_rx_data[48], w_hssi_rx_pld_pcs_interface_pld_rx_data[47], w_hssi_rx_pld_pcs_interface_pld_rx_data[46], w_hssi_rx_pld_pcs_interface_pld_rx_data[45], w_hssi_rx_pld_pcs_interface_pld_rx_data[44], w_hssi_rx_pld_pcs_interface_pld_rx_data[43], w_hssi_rx_pld_pcs_interface_pld_rx_data[42], w_hssi_rx_pld_pcs_interface_pld_rx_data[41], w_hssi_rx_pld_pcs_interface_pld_rx_data[40], w_hssi_rx_pld_pcs_interface_pld_rx_data[39], w_hssi_rx_pld_pcs_interface_pld_rx_data[38], w_hssi_rx_pld_pcs_interface_pld_rx_data[37], w_hssi_rx_pld_pcs_interface_pld_rx_data[36], w_hssi_rx_pld_pcs_interface_pld_rx_data[35], w_hssi_rx_pld_pcs_interface_pld_rx_data[34], w_hssi_rx_pld_pcs_interface_pld_rx_data[33], w_hssi_rx_pld_pcs_interface_pld_rx_data[32], w_hssi_rx_pld_pcs_interface_pld_rx_data[31], w_hssi_rx_pld_pcs_interface_pld_rx_data[30], w_hssi_rx_pld_pcs_interface_pld_rx_data[29], w_hssi_rx_pld_pcs_interface_pld_rx_data[28], w_hssi_rx_pld_pcs_interface_pld_rx_data[27], w_hssi_rx_pld_pcs_interface_pld_rx_data[26], w_hssi_rx_pld_pcs_interface_pld_rx_data[25], w_hssi_rx_pld_pcs_interface_pld_rx_data[24], w_hssi_rx_pld_pcs_interface_pld_rx_data[23], w_hssi_rx_pld_pcs_interface_pld_rx_data[22], w_hssi_rx_pld_pcs_interface_pld_rx_data[21], w_hssi_rx_pld_pcs_interface_pld_rx_data[20], w_hssi_rx_pld_pcs_interface_pld_rx_data[19], w_hssi_rx_pld_pcs_interface_pld_rx_data[18], w_hssi_rx_pld_pcs_interface_pld_rx_data[17], w_hssi_rx_pld_pcs_interface_pld_rx_data[16], w_hssi_rx_pld_pcs_interface_pld_rx_data[15], w_hssi_rx_pld_pcs_interface_pld_rx_data[14], w_hssi_rx_pld_pcs_interface_pld_rx_data[13], w_hssi_rx_pld_pcs_interface_pld_rx_data[12], w_hssi_rx_pld_pcs_interface_pld_rx_data[11], w_hssi_rx_pld_pcs_interface_pld_rx_data[10], w_hssi_rx_pld_pcs_interface_pld_rx_data[9], w_hssi_rx_pld_pcs_interface_pld_rx_data[8], w_hssi_rx_pld_pcs_interface_pld_rx_data[7], w_hssi_rx_pld_pcs_interface_pld_rx_data[6], w_hssi_rx_pld_pcs_interface_pld_rx_data[5], w_hssi_rx_pld_pcs_interface_pld_rx_data[4], w_hssi_rx_pld_pcs_interface_pld_rx_data[3], w_hssi_rx_pld_pcs_interface_pld_rx_data[2], w_hssi_rx_pld_pcs_interface_pld_rx_data[1], w_hssi_rx_pld_pcs_interface_pld_rx_data[0]};
		assign out_pld_rx_prbs_done = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
		assign out_pld_rx_prbs_err = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
		assign out_pld_test_data = {w_hssi_common_pld_pcs_interface_pld_test_data[19], w_hssi_common_pld_pcs_interface_pld_test_data[18], w_hssi_common_pld_pcs_interface_pld_test_data[17], w_hssi_common_pld_pcs_interface_pld_test_data[16], w_hssi_common_pld_pcs_interface_pld_test_data[15], w_hssi_common_pld_pcs_interface_pld_test_data[14], w_hssi_common_pld_pcs_interface_pld_test_data[13], w_hssi_common_pld_pcs_interface_pld_test_data[12], w_hssi_common_pld_pcs_interface_pld_test_data[11], w_hssi_common_pld_pcs_interface_pld_test_data[10], w_hssi_common_pld_pcs_interface_pld_test_data[9], w_hssi_common_pld_pcs_interface_pld_test_data[8], w_hssi_common_pld_pcs_interface_pld_test_data[7], w_hssi_common_pld_pcs_interface_pld_test_data[6], w_hssi_common_pld_pcs_interface_pld_test_data[5], w_hssi_common_pld_pcs_interface_pld_test_data[4], w_hssi_common_pld_pcs_interface_pld_test_data[3], w_hssi_common_pld_pcs_interface_pld_test_data[2], w_hssi_common_pld_pcs_interface_pld_test_data[1], w_hssi_common_pld_pcs_interface_pld_test_data[0]};
		assign out_pld_uhsif_lock = w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
		assign out_pld_uhsif_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
		assign out_pma_adapt_start = w_hssi_common_pcs_pma_interface_pma_adapt_start;
		assign out_pma_atpg_los_en_n = w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
		assign out_pma_csr_test_dis = w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
		assign out_pma_current_coeff = {w_hssi_common_pcs_pma_interface_pma_current_coeff[17], w_hssi_common_pcs_pma_interface_pma_current_coeff[16], w_hssi_common_pcs_pma_interface_pma_current_coeff[15], w_hssi_common_pcs_pma_interface_pma_current_coeff[14], w_hssi_common_pcs_pma_interface_pma_current_coeff[13], w_hssi_common_pcs_pma_interface_pma_current_coeff[12], w_hssi_common_pcs_pma_interface_pma_current_coeff[11], w_hssi_common_pcs_pma_interface_pma_current_coeff[10], w_hssi_common_pcs_pma_interface_pma_current_coeff[9], w_hssi_common_pcs_pma_interface_pma_current_coeff[8], w_hssi_common_pcs_pma_interface_pma_current_coeff[7], w_hssi_common_pcs_pma_interface_pma_current_coeff[6], w_hssi_common_pcs_pma_interface_pma_current_coeff[5], w_hssi_common_pcs_pma_interface_pma_current_coeff[4], w_hssi_common_pcs_pma_interface_pma_current_coeff[3], w_hssi_common_pcs_pma_interface_pma_current_coeff[2], w_hssi_common_pcs_pma_interface_pma_current_coeff[1], w_hssi_common_pcs_pma_interface_pma_current_coeff[0]};
		assign out_pma_current_rxpreset = {w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[1], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[0]};
		assign out_pma_early_eios = w_hssi_common_pcs_pma_interface_pma_early_eios;
		assign out_pma_eye_monitor = {w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0]};
		assign out_pma_interface_select = {w_hssi_common_pcs_pma_interface_pma_interface_select[1], w_hssi_common_pcs_pma_interface_pma_interface_select[0]};
		assign out_pma_ltd_b = w_hssi_common_pcs_pma_interface_pma_ltd_b;
		assign out_pma_ltr = w_hssi_common_pcs_pma_interface_pma_ltr;
		assign out_pma_nfrzdrv = w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
		assign out_pma_nrpi_freeze = w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
		assign out_pma_pcie_switch = {w_hssi_common_pcs_pma_interface_pma_pcie_switch[1], w_hssi_common_pcs_pma_interface_pma_pcie_switch[0]};
		assign out_pma_ppm_lock = w_hssi_common_pcs_pma_interface_pma_ppm_lock;
		assign out_pma_reserved_out = {w_hssi_common_pcs_pma_interface_pma_reserved_out[4], w_hssi_common_pcs_pma_interface_pma_reserved_out[3], w_hssi_common_pcs_pma_interface_pma_reserved_out[2], w_hssi_common_pcs_pma_interface_pma_reserved_out[1], w_hssi_common_pcs_pma_interface_pma_reserved_out[0]};
		assign out_pma_rs_lpbk_b = w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
		assign out_pma_rx_clkslip = w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
		assign out_pma_rx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
		assign out_pma_rxpma_rstb = w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
		assign out_pma_scan_mode_n = w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
		assign out_pma_scan_shift_n = w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
		assign out_pma_tx_bitslip = w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
		assign out_pma_tx_bonding_rstb = w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
		assign out_pma_tx_elec_idle = w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
		assign out_pma_tx_pma_data = {w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0]};
		assign out_pma_tx_qpi_pulldn = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
		assign out_pma_tx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
		assign out_pma_tx_txdetectrx = w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
		assign out_pma_txpma_rstb = w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	endgenerate
endmodule
module twentynm_pcs_rev_20nm4es
	#(
	//PARAM_LIST_START
		parameter xcvr_native_mode = "mode_duplex",  // mode_duplex, mode_rx_only, mode_tx_only
		
		// parameters for twentynm_hssi_10g_rx_pcs
		parameter hssi_10g_rx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_align_del = "align_del_en", // align_del_dis|align_del_en
		parameter hssi_10g_rx_pcs_ber_bit_err_total_cnt = "bit_err_total_cnt_10g", // bit_err_total_cnt_10g
		parameter hssi_10g_rx_pcs_ber_clken = "ber_clk_dis", // ber_clk_dis|ber_clk_en
		parameter hssi_10g_rx_pcs_ber_xus_timer_window = 21'b100110001001010,
		parameter hssi_10g_rx_pcs_bitslip_mode = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_rx_pcs_blksync_bitslip_type = "bitslip_comb", // bitslip_comb|bitslip_reg
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_cnt = 3'b1,
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_type = "bitslip_match", // bitslip_match|bitslip_cnt
		parameter hssi_10g_rx_pcs_blksync_bypass = "blksync_bypass_dis", // blksync_bypass_dis|blksync_bypass_en
		parameter hssi_10g_rx_pcs_blksync_clken = "blksync_clk_dis", // blksync_clk_dis|blksync_clk_en
		parameter hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt = "enum_invalid_sh_cnt_10g", // enum_invalid_sh_cnt_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock = "knum_sh_cnt_postlock_10g", // knum_sh_cnt_postlock_10g
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock = "knum_sh_cnt_prelock_10g", // knum_sh_cnt_prelock_10g
		parameter hssi_10g_rx_pcs_blksync_pipeln = "blksync_pipeln_dis", // blksync_pipeln_dis|blksync_pipeln_en
		parameter hssi_10g_rx_pcs_clr_errblk_cnt_en = "disable", // disable|enable
		parameter hssi_10g_rx_pcs_control_del = "control_del_all", // control_del_all|control_del_none
		parameter hssi_10g_rx_pcs_crcchk_bypass = "crcchk_bypass_dis", // crcchk_bypass_dis|crcchk_bypass_en
		parameter hssi_10g_rx_pcs_crcchk_clken = "crcchk_clk_dis", // crcchk_clk_dis|crcchk_clk_en
		parameter hssi_10g_rx_pcs_crcchk_inv = "crcchk_inv_dis", // crcchk_inv_dis|crcchk_inv_en
		parameter hssi_10g_rx_pcs_crcchk_pipeln = "crcchk_pipeln_dis", // crcchk_pipeln_dis|crcchk_pipeln_en
		parameter hssi_10g_rx_pcs_crcflag_pipeln = "crcflag_pipeln_dis", // crcflag_pipeln_dis|crcflag_pipeln_en
		parameter hssi_10g_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_rx_pcs_dec64b66b_clken = "dec64b66b_clk_dis", // dec64b66b_clk_dis|dec64b66b_clk_en
		parameter hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass = "dec_64b66b_rxsm_bypass_dis", // dec_64b66b_rxsm_bypass_dis|dec_64b66b_rxsm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_bypass = "descrm_bypass_en", // descrm_bypass_dis|descrm_bypass_en
		parameter hssi_10g_rx_pcs_descrm_clken = "descrm_clk_dis", // descrm_clk_dis|descrm_clk_en
		parameter hssi_10g_rx_pcs_descrm_mode = "async", // async|sync
		parameter hssi_10g_rx_pcs_descrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_dft_clk_out_sel = "rx_master_clk", // rx_master_clk|rx_gbexp_clk|rx_blksync_clk|rx_descrm_clk|rx_frmsync_clk|rx_64b66bdec_clk|rx_ber_clk|rx_rand_clk|rx_crcchk_clk|rx_wrfifo_clk|rx_rdfifo_clk|rx_fec_clk
		parameter hssi_10g_rx_pcs_dis_signal_ok = "dis_signal_ok_dis", // dis_signal_ok_dis|dis_signal_ok_en
		parameter hssi_10g_rx_pcs_dispchk_bypass = "dispchk_bypass_dis", // dispchk_bypass_dis|dispchk_bypass_en
		parameter hssi_10g_rx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_rx_pcs_fast_path = "fast_path_dis", // fast_path_dis|fast_path_en
		parameter hssi_10g_rx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_rx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_rx_pcs_fifo_double_read = "fifo_double_read_dis", // fifo_double_read_dis|fifo_double_read_en
		parameter hssi_10g_rx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_rx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_rx_pcs_force_align = "force_align_dis", // force_align_dis|force_align_en
		parameter hssi_10g_rx_pcs_frmsync_bypass = "frmsync_bypass_dis", // frmsync_bypass_dis|frmsync_bypass_en
		parameter hssi_10g_rx_pcs_frmsync_clken = "frmsync_clk_dis", // frmsync_clk_dis|frmsync_clk_en
		parameter hssi_10g_rx_pcs_frmsync_enum_scrm = "enum_scrm_default", // enum_scrm_default
		parameter hssi_10g_rx_pcs_frmsync_enum_sync = "enum_sync_default", // enum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_flag_type = "all_framing_words", // all_framing_words|location_only
		parameter hssi_10g_rx_pcs_frmsync_knum_sync = "knum_sync_default", // knum_sync_default
		parameter hssi_10g_rx_pcs_frmsync_mfrm_length = 16'b100000000000,
		parameter hssi_10g_rx_pcs_frmsync_pipeln = "frmsync_pipeln_dis", // frmsync_pipeln_dis|frmsync_pipeln_en
		parameter hssi_10g_rx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_rx_pcs_gb_rx_idwidth = "width_32", // width_40|width_32|width_64
		parameter hssi_10g_rx_pcs_gb_rx_odwidth = "width_66", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_rx_pcs_gbexp_clken = "gbexp_clk_dis", // gbexp_clk_dis|gbexp_clk_en
		parameter hssi_10g_rx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_10g_rx_pcs_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_rx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_rx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_rx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_rx_pcs_pld_if_type = "fifo", // fifo|reg
		parameter hssi_10g_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_rx_pcs_rand_clken = "rand_clk_dis", // rand_clk_dis|rand_clk_en
		parameter hssi_10g_rx_pcs_rd_clk_sel = "rd_rx_pma_clk", // rd_rx_pld_clk|rd_rx_pma_clk|rd_refclk_dig
		parameter hssi_10g_rx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_rx_pcs_rx_fifo_write_ctrl = "blklock_stops", // blklock_stops|blklock_ignore
		parameter hssi_10g_rx_pcs_rx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_rx_pcs_rx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_rx_pcs_rx_signal_ok_sel = "synchronized_ver", // synchronized_ver|nonsync_ver
		parameter hssi_10g_rx_pcs_rx_sm_bypass = "rx_sm_bypass_dis", // rx_sm_bypass_dis|rx_sm_bypass_en
		parameter hssi_10g_rx_pcs_rx_sm_hiber = "rx_sm_hiber_en", // rx_sm_hiber_en|rx_sm_hiber_dis
		parameter hssi_10g_rx_pcs_rx_sm_pipeln = "rx_sm_pipeln_dis", // rx_sm_pipeln_dis|rx_sm_pipeln_en
		parameter hssi_10g_rx_pcs_rx_testbus_sel = "crc32_chk_testbus1", // crc32_chk_testbus1|crc32_chk_testbus2|frame_sync_testbus1|frame_sync_testbus2|dec64b66b_testbus|rxsm_testbus|ber_testbus|blksync_testbus1|blksync_testbus2|gearbox_exp_testbus|random_ver_testbus|descramble_testbus|blank_testbus|rx_fifo_testbus1|rx_fifo_testbus2
		parameter hssi_10g_rx_pcs_rx_true_b2b = "b2b", // single|b2b
		parameter hssi_10g_rx_pcs_rxfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_rx_pcs_rxfifo_full = "full_default", // full_default
		parameter hssi_10g_rx_pcs_rxfifo_mode = "phase_comp", // register_mode|clk_comp_10g|generic_interlaken|generic_basic|phase_comp|phase_comp_dv
		parameter hssi_10g_rx_pcs_rxfifo_pempty = 5'b10,
		parameter hssi_10g_rx_pcs_rxfifo_pfull = 5'b10111,
		parameter hssi_10g_rx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_rx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_rx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_10g_tx_pcs
		parameter hssi_10g_tx_pcs_advanced_user_mode = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_bitslip_en = "bitslip_dis", // bitslip_dis|bitslip_en
		parameter hssi_10g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_10g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_10g_tx_pcs_comp_cnt = 8'b0,
		parameter hssi_10g_tx_pcs_compin_sel = "compin_master", // compin_master|compin_slave_top|compin_slave_bot|compin_default
		parameter hssi_10g_tx_pcs_crcgen_bypass = "crcgen_bypass_dis", // crcgen_bypass_dis|crcgen_bypass_en
		parameter hssi_10g_tx_pcs_crcgen_clken = "crcgen_clk_dis", // crcgen_clk_dis|crcgen_clk_en
		parameter hssi_10g_tx_pcs_crcgen_err = "crcgen_err_dis", // crcgen_err_dis|crcgen_err_en
		parameter hssi_10g_tx_pcs_crcgen_inv = "crcgen_inv_dis", // crcgen_inv_dis|crcgen_inv_en
		parameter hssi_10g_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_10g_tx_pcs_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_10g_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_10g_tx_pcs_dft_clk_out_sel = "tx_master_clk", // tx_master_clk|tx_rdfifo_clk|tx_frmgen_clk|tx_crcgen_clk|tx_64b66benc_txsm_clk|tx_scrm_clk|tx_dispgen_clk|tx_gbred_clk|tx_wrfifo_clk|tx_fec_clk
		parameter hssi_10g_tx_pcs_dispgen_bypass = "dispgen_bypass_dis", // dispgen_bypass_dis|dispgen_bypass_en
		parameter hssi_10g_tx_pcs_dispgen_clken = "dispgen_clk_dis", // dispgen_clk_dis|dispgen_clk_en
		parameter hssi_10g_tx_pcs_dispgen_err = "dispgen_err_dis", // dispgen_err_dis|dispgen_err_en
		parameter hssi_10g_tx_pcs_dispgen_pipeln = "dispgen_pipeln_dis", // dispgen_pipeln_dis|dispgen_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_bypass_pipeln = "distdwn_bypass_pipeln_dis", // distdwn_bypass_pipeln_dis|distdwn_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distdwn_master = "distdwn_master_en", // distdwn_master_en|distdwn_master_dis
		parameter hssi_10g_tx_pcs_distup_bypass_pipeln = "distup_bypass_pipeln_dis", // distup_bypass_pipeln_dis|distup_bypass_pipeln_en
		parameter hssi_10g_tx_pcs_distup_master = "distup_master_en", // distup_master_en|distup_master_dis
		parameter hssi_10g_tx_pcs_dv_bond = "dv_bond_dis", // dv_bond_en|dv_bond_dis
		parameter hssi_10g_tx_pcs_empty_flag_type = "empty_rd_side", // empty_rd_side|empty_wr_side
		parameter hssi_10g_tx_pcs_enc64b66b_txsm_clken = "enc64b66b_txsm_clk_dis", // enc64b66b_txsm_clk_dis|enc64b66b_txsm_clk_en
		parameter hssi_10g_tx_pcs_enc_64b66b_txsm_bypass = "enc_64b66b_txsm_bypass_dis", // enc_64b66b_txsm_bypass_dis|enc_64b66b_txsm_bypass_en
		parameter hssi_10g_tx_pcs_fastpath = "fastpath_dis", // fastpath_dis|fastpath_en
		parameter hssi_10g_tx_pcs_fec_clken = "fec_clk_dis", // fec_clk_dis|fec_clk_en
		parameter hssi_10g_tx_pcs_fec_enable = "fec_dis", // fec_en|fec_dis
		parameter hssi_10g_tx_pcs_fifo_double_write = "fifo_double_write_dis", // fifo_double_write_dis|fifo_double_write_en
		parameter hssi_10g_tx_pcs_fifo_reg_fast = "fifo_reg_fast_dis", // fifo_reg_fast_dis|fifo_reg_fast_en
		parameter hssi_10g_tx_pcs_fifo_stop_rd = "n_rd_empty", // rd_empty|n_rd_empty
		parameter hssi_10g_tx_pcs_fifo_stop_wr = "n_wr_full", // wr_full|n_wr_full
		parameter hssi_10g_tx_pcs_frmgen_burst = "frmgen_burst_dis", // frmgen_burst_dis|frmgen_burst_en
		parameter hssi_10g_tx_pcs_frmgen_bypass = "frmgen_bypass_dis", // frmgen_bypass_dis|frmgen_bypass_en
		parameter hssi_10g_tx_pcs_frmgen_clken = "frmgen_clk_dis", // frmgen_clk_dis|frmgen_clk_en
		parameter hssi_10g_tx_pcs_frmgen_mfrm_length = 16'b100000000000,
		parameter hssi_10g_tx_pcs_frmgen_pipeln = "frmgen_pipeln_dis", // frmgen_pipeln_dis|frmgen_pipeln_en
		parameter hssi_10g_tx_pcs_frmgen_pyld_ins = "frmgen_pyld_ins_dis", // frmgen_pyld_ins_dis|frmgen_pyld_ins_en
		parameter hssi_10g_tx_pcs_frmgen_wordslip = "frmgen_wordslip_dis", // frmgen_wordslip_dis|frmgen_wordslip_en
		parameter hssi_10g_tx_pcs_full_flag_type = "full_wr_side", // full_rd_side|full_wr_side
		parameter hssi_10g_tx_pcs_gb_pipeln_bypass = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_gb_tx_idwidth = "width_50", // width_32|width_40|width_50|width_67|width_64|width_66
		parameter hssi_10g_tx_pcs_gb_tx_odwidth = "width_32", // width_32|width_40|width_64
		parameter hssi_10g_tx_pcs_gbred_clken = "gbred_clk_dis", // gbred_clk_dis|gbred_clk_en
		parameter hssi_10g_tx_pcs_indv = "indv_en", // indv_en|indv_dis
		parameter hssi_10g_tx_pcs_low_latency_en = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_10g_tx_pcs_pempty_flag_type = "pempty_rd_side", // pempty_rd_side|pempty_wr_side
		parameter hssi_10g_tx_pcs_pfull_flag_type = "pfull_wr_side", // pfull_rd_side|pfull_wr_side
		parameter hssi_10g_tx_pcs_phcomp_rd_del = "phcomp_rd_del2", // phcomp_rd_del6|phcomp_rd_del5|phcomp_rd_del4|phcomp_rd_del3|phcomp_rd_del2
		parameter hssi_10g_tx_pcs_pld_if_type = "fifo", // fifo|reg|fastreg
		parameter hssi_10g_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_baser_mode|interlaken_mode|sfis_mode|teng_sdi_mode|basic_mode|test_prp_mode|test_prp_krfec_mode|teng_1588_mode|teng_baser_krfec_mode|teng_1588_krfec_mode|basic_krfec_mode
		parameter hssi_10g_tx_pcs_pseudo_random = "all_0", // two_lf|all_0
		parameter hssi_10g_tx_pcs_pseudo_seed_a = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_pseudo_seed_b = 58'b1111111111111111111111111111111111111111111111111111111111,
		parameter hssi_10g_tx_pcs_random_disp = "disable", // disable|enable
		parameter hssi_10g_tx_pcs_rdfifo_clken = "rdfifo_clk_dis", // rdfifo_clk_dis|rdfifo_clk_en
		parameter hssi_10g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_10g_tx_pcs_scrm_bypass = "scrm_bypass_dis", // scrm_bypass_dis|scrm_bypass_en
		parameter hssi_10g_tx_pcs_scrm_clken = "scrm_clk_dis", // scrm_clk_dis|scrm_clk_en
		parameter hssi_10g_tx_pcs_scrm_mode = "async", // async|sync
		parameter hssi_10g_tx_pcs_scrm_pipeln = "enable", // disable|enable
		parameter hssi_10g_tx_pcs_sh_err = "sh_err_dis", // sh_err_dis|sh_err_en
		parameter hssi_10g_tx_pcs_sop_mark = "sop_mark_dis", // sop_mark_en|sop_mark_dis
		parameter hssi_10g_tx_pcs_stretch_num_stages = "zero_stage", // zero_stage|one_stage|two_stage|three_stage
		parameter hssi_10g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_10g_tx_pcs_test_mode = "test_off", // test_off|pseudo_random
		parameter hssi_10g_tx_pcs_tx_scrm_err = "scrm_err_dis", // scrm_err_dis|scrm_err_en
		parameter hssi_10g_tx_pcs_tx_scrm_width = "bit64", // bit64|bit66|bit67
		parameter hssi_10g_tx_pcs_tx_sh_location = "lsb", // lsb|msb
		parameter hssi_10g_tx_pcs_tx_sm_bypass = "tx_sm_bypass_dis", // tx_sm_bypass_dis|tx_sm_bypass_en
		parameter hssi_10g_tx_pcs_tx_sm_pipeln = "tx_sm_pipeln_dis", // tx_sm_pipeln_dis|tx_sm_pipeln_en
		parameter hssi_10g_tx_pcs_tx_testbus_sel = "crc32_gen_testbus1", // crc32_gen_testbus1|crc32_gen_testbus2|disp_gen_testbus1|disp_gen_testbus2|frame_gen_testbus1|frame_gen_testbus2|enc64b66b_testbus|txsm_testbus|tx_cp_bond_testbus|gearbox_red_testbus|scramble_testbus|blank_testbus|tx_fifo_testbus1|tx_fifo_testbus2
		parameter hssi_10g_tx_pcs_txfifo_empty = "empty_default", // empty_default
		parameter hssi_10g_tx_pcs_txfifo_full = "full_default", // full_default
		parameter hssi_10g_tx_pcs_txfifo_mode = "phase_comp", // register_mode|interlaken_generic|basic_generic|phase_comp
		parameter hssi_10g_tx_pcs_txfifo_pempty = 4'b10,
		parameter hssi_10g_tx_pcs_txfifo_pfull = 4'b1011,
		parameter hssi_10g_tx_pcs_wr_clk_sel = "wr_tx_pma_clk", // wr_tx_pld_clk|wr_tx_pma_clk|wr_refclk_dig
		parameter hssi_10g_tx_pcs_wrfifo_clken = "wrfifo_clk_dis", // wrfifo_clk_dis|wrfifo_clk_en
		
		// parameters for twentynm_hssi_8g_rx_pcs
		parameter hssi_8g_rx_pcs_auto_error_replacement = "dis_err_replace", // dis_err_replace|en_err_replace
		parameter hssi_8g_rx_pcs_auto_speed_nego = "dis_asn", // dis_asn|en_asn_g2_freq_scal
		parameter hssi_8g_rx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_rx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_rx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_rx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_rx_pcs_byte_deserializer = "dis_bds", // dis_bds|en_bds_by_2|en_bds_by_4|en_bds_by_2_det
		parameter hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask = "dis_rxvalid_mask", // dis_rxvalid_mask|en_rxvalid_mask
		parameter hssi_8g_rx_pcs_clkcmp_pattern_n = 20'b0,
		parameter hssi_8g_rx_pcs_clkcmp_pattern_p = 20'b0,
		parameter hssi_8g_rx_pcs_clock_gate_bds_dec_asn = "dis_bds_dec_asn_clk_gating", // dis_bds_dec_asn_clk_gating|en_bds_dec_asn_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_cdr_eidle = "dis_cdr_eidle_clk_gating", // dis_cdr_eidle_clk_gating|en_cdr_eidle_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk = "dis_dw_pc_wrclk_gating", // dis_dw_pc_wrclk_gating|en_dw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_rd = "dis_dw_rm_rdclk_gating", // dis_dw_rm_rdclk_gating|en_dw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_wr = "dis_dw_rm_wrclk_gating", // dis_dw_rm_wrclk_gating|en_dw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_dw_wa = "dis_dw_wa_clk_gating", // dis_dw_wa_clk_gating|en_dw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_gate_pc_rdclk = "dis_pc_rdclk_gating", // dis_pc_rdclk_gating|en_pc_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk = "dis_sw_pc_wrclk_gating", // dis_sw_pc_wrclk_gating|en_sw_pc_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_rd = "dis_sw_rm_rdclk_gating", // dis_sw_rm_rdclk_gating|en_sw_rm_rdclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_wr = "dis_sw_rm_wrclk_gating", // dis_sw_rm_wrclk_gating|en_sw_rm_wrclk_gating
		parameter hssi_8g_rx_pcs_clock_gate_sw_wa = "dis_sw_wa_clk_gating", // dis_sw_wa_clk_gating|en_sw_wa_clk_gating
		parameter hssi_8g_rx_pcs_clock_observation_in_pld_core = "internal_sw_wa_clk", // internal_sw_wa_clk|internal_dw_wa_clk|internal_cdr_eidle_clk|internal_sm_rm_wr_clk|internal_dw_rm_wr_clk|internal_clk_2_b|internal_sw_rm_rd_clk|internal_dw_rm_rd_clk|internal_sw_rx_wr_clk|internal_dw_rx_wr_clk|internal_rx_rd_clk|internal_rx_pma_clk_gen3|internal_rx_rcvd_clk_gen3
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_rx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_rx_pcs_eidle_entry_eios = "dis_eidle_eios", // dis_eidle_eios|en_eidle_eios
		parameter hssi_8g_rx_pcs_eidle_entry_iei = "dis_eidle_iei", // dis_eidle_iei|en_eidle_iei
		parameter hssi_8g_rx_pcs_eidle_entry_sd = "dis_eidle_sd", // dis_eidle_sd|en_eidle_sd
		parameter hssi_8g_rx_pcs_eightb_tenb_decoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_rx_pcs_err_flags_sel = "err_flags_wa", // err_flags_wa|err_flags_8b10b
		parameter hssi_8g_rx_pcs_fixed_pat_det = "dis_fixed_patdet", // dis_fixed_patdet|en_fixed_patdet
		parameter hssi_8g_rx_pcs_fixed_pat_num = 4'b1111,
		parameter hssi_8g_rx_pcs_force_signal_detect = "en_force_signal_detect", // en_force_signal_detect|dis_force_signal_detect
		parameter hssi_8g_rx_pcs_gen3_clk_en = "disable_clk", // disable_clk|enable_clk
		parameter hssi_8g_rx_pcs_gen3_rx_clk_sel = "rcvd_clk", // en_dig_clk1_8g|rcvd_clk
		parameter hssi_8g_rx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // en_dig_clk2_8g|tx_pma_clk
		parameter hssi_8g_rx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_rx_pcs_ibm_invalid_code = "dis_ibm_invalid_code", // dis_ibm_invalid_code|en_ibm_invalid_code
		parameter hssi_8g_rx_pcs_invalid_code_flag_only = "dis_invalid_code_only", // dis_invalid_code_only|en_invalid_code_only
		parameter hssi_8g_rx_pcs_pad_or_edb_error_replace = "replace_edb", // replace_edb|replace_edb_dynamic|replace_pad
		parameter hssi_8g_rx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_rx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_rx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_rx_pcs_pipe_if_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_8g_rx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_rx_pcs_polinv_8b10b_dec = "dis_polinv_8b10b_dec", // dis_polinv_8b10b_dec|en_polinv_8b10b_dec
		parameter hssi_8g_rx_pcs_prot_mode = "gige", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic_rm_enable|basic_rm_disable|disabled_prot_mode
		parameter hssi_8g_rx_pcs_rate_match = "dis_rm", // dis_rm|gige_rm|pipe_rm|pipe_rm_0ppm|sw_basic_rm|dw_basic_rm
		parameter hssi_8g_rx_pcs_rate_match_del_thres = "dis_rm_del_thres", // dis_rm_del_thres|gige_rm_del_thres|pipe_rm_del_thres|pipe_rm_0ppm_del_thres|sw_basic_rm_del_thres|dw_basic_rm_del_thres
		parameter hssi_8g_rx_pcs_rate_match_empty_thres = "dis_rm_empty_thres", // dis_rm_empty_thres|gige_rm_empty_thres|pipe_rm_empty_thres|pipe_rm_0ppm_empty_thres|sw_basic_rm_empty_thres|dw_basic_rm_empty_thres
		parameter hssi_8g_rx_pcs_rate_match_full_thres = "dis_rm_full_thres", // dis_rm_full_thres|gige_rm_full_thres|pipe_rm_full_thres|pipe_rm_0ppm_full_thres|sw_basic_rm_full_thres|dw_basic_rm_full_thres
		parameter hssi_8g_rx_pcs_rate_match_ins_thres = "dis_rm_ins_thres", // dis_rm_ins_thres|gige_rm_ins_thres|pipe_rm_ins_thres|pipe_rm_0ppm_ins_thres|sw_basic_rm_ins_thres|dw_basic_rm_ins_thres
		parameter hssi_8g_rx_pcs_rate_match_start_thres = "dis_rm_start_thres", // dis_rm_start_thres|gige_rm_start_thres|pipe_rm_start_thres|pipe_rm_0ppm_start_thres|sw_basic_rm_start_thres|dw_basic_rm_start_thres
		parameter hssi_8g_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_rx_pcs_rx_clk2 = "rcvd_clk_clk2", // rcvd_clk_clk2|tx_pma_clock_clk2|refclk_dig2_clk2
		parameter hssi_8g_rx_pcs_rx_clk_free_running = "en_rx_clk_free_run", // dis_rx_clk_free_run|en_rx_clk_free_run
		parameter hssi_8g_rx_pcs_rx_pcs_urst = "en_rx_pcs_urst", // dis_rx_pcs_urst|en_rx_pcs_urst
		parameter hssi_8g_rx_pcs_rx_rcvd_clk = "rcvd_clk_rcvd_clk", // rcvd_clk_rcvd_clk|tx_pma_clock_rcvd_clk
		parameter hssi_8g_rx_pcs_rx_rd_clk = "pld_rx_clk", // pld_rx_clk|rx_clk
		parameter hssi_8g_rx_pcs_rx_refclk = "dis_refclk_sel", // dis_refclk_sel|en_refclk_sel
		parameter hssi_8g_rx_pcs_rx_wr_clk = "rx_clk2_div_1_2_4", // rx_clk2_div_1_2_4|txfifo_rd_clk
		parameter hssi_8g_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_rx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_rx_pcs_sync_sm_idle_eios = "dis_syncsm_idle", // dis_syncsm_idle|en_syncsm_idle
		parameter hssi_8g_rx_pcs_test_bus_sel = "tx_testbus", // tx_testbus|tx_ctrl_plane_testbus|wa_testbus|rm_testbus|rx_ctrl_testbus|pcie_ctrl_testbus|rx_ctrl_plane_testbus
		parameter hssi_8g_rx_pcs_tx_rx_parallel_loopback = "dis_plpbk", // dis_plpbk|en_plpbk
		parameter hssi_8g_rx_pcs_wa_boundary_lock_ctrl = "bit_slip", // bit_slip|sync_sm|deterministic_latency|auto_align_pld_ctrl
		parameter hssi_8g_rx_pcs_wa_clk_slip_spacing = 10'b10000,
		parameter hssi_8g_rx_pcs_wa_det_latency_sync_status_beh = "assert_sync_status_non_imm", // assert_sync_status_imm|assert_sync_status_non_imm|dont_care_assert_sync
		parameter hssi_8g_rx_pcs_wa_disp_err_flag = "dis_disp_err_flag", // dis_disp_err_flag|en_disp_err_flag
		parameter hssi_8g_rx_pcs_wa_kchar = "dis_kchar", // dis_kchar|en_kchar
		parameter hssi_8g_rx_pcs_wa_pd = "wa_pd_10", // wa_pd_7|wa_pd_10|wa_pd_20|wa_pd_40|wa_pd_8_sw|wa_pd_8_dw|wa_pd_16_sw|wa_pd_16_dw|wa_pd_32
		parameter hssi_8g_rx_pcs_wa_pd_data = 40'b0,
		parameter hssi_8g_rx_pcs_wa_pd_polarity = "dis_pd_both_pol", // dis_pd_both_pol|en_pd_both_pol|dont_care_both_pol
		parameter hssi_8g_rx_pcs_wa_pld_controlled = "dis_pld_ctrl", // dis_pld_ctrl|pld_ctrl_sw|rising_edge_sensitive_dw|level_sensitive_dw
		parameter hssi_8g_rx_pcs_wa_renumber_data = 6'b0,
		parameter hssi_8g_rx_pcs_wa_rgnumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rknumber_data = 8'b0,
		parameter hssi_8g_rx_pcs_wa_rosnumber_data = 2'b0,
		parameter hssi_8g_rx_pcs_wa_rvnumber_data = 13'b0,
		parameter hssi_8g_rx_pcs_wa_sync_sm_ctrl = "gige_sync_sm", // gige_sync_sm|pipe_sync_sm|sw_basic_sync_sm|dw_basic_sync_sm|fibre_channel_sync_sm
		parameter hssi_8g_rx_pcs_wait_cnt = 12'b0,
		
		// parameters for twentynm_hssi_8g_tx_pcs
		parameter hssi_8g_tx_pcs_auto_speed_nego_gen2 = "dis_asn_g2", // dis_asn_g2|en_asn_g2_freq_scal
		parameter hssi_8g_tx_pcs_bit_reversal = "dis_bit_reversal", // dis_bit_reversal|en_bit_reversal
		parameter hssi_8g_tx_pcs_bonding_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_8g_tx_pcs_bonding_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_8g_tx_pcs_bypass_pipeline_reg = "dis_bypass_pipeline", // dis_bypass_pipeline|en_bypass_pipeline
		parameter hssi_8g_tx_pcs_byte_serializer = "dis_bs", // dis_bs|en_bs_by_2|en_bs_by_4
		parameter hssi_8g_tx_pcs_clock_gate_bs_enc = "dis_bs_enc_clk_gating", // dis_bs_enc_clk_gating|en_bs_enc_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_dw_fifowr = "dis_dw_fifowr_clk_gating", // dis_dw_fifowr_clk_gating|en_dw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_fiford = "dis_fiford_clk_gating", // dis_fiford_clk_gating|en_fiford_clk_gating
		parameter hssi_8g_tx_pcs_clock_gate_sw_fifowr = "dis_sw_fifowr_clk_gating", // dis_sw_fifowr_clk_gating|en_sw_fifowr_clk_gating
		parameter hssi_8g_tx_pcs_clock_observation_in_pld_core = "internal_refclk_b", // internal_refclk_b|internal_fifo_rd_clk|internal_sw_fifo_wr_clk|internal_dw_fifo_wr_clk|internal_tx_clk_out_gen3|internal_pipe_tx_clk_out_gen3
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_compensation = "dis_compensation", // dis_compensation|en_compensation
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_consumption = "individual", // individual|bundled_master|bundled_slave_below|bundled_slave_above
		parameter hssi_8g_tx_pcs_ctrl_plane_bonding_distribution = "not_master_chnl_distr", // not_master_chnl_distr|master_chnl_distr
		parameter hssi_8g_tx_pcs_data_selection_8b10b_encoder_input = "normal_data_path", // normal_data_path|gige_idle_conversion
		parameter hssi_8g_tx_pcs_dynamic_clk_switch = "dis_dyn_clk_switch", // dis_dyn_clk_switch|en_dyn_clk_switch
		parameter hssi_8g_tx_pcs_eightb_tenb_disp_ctrl = "dis_disp_ctrl", // dis_disp_ctrl|en_disp_ctrl|en_ib_disp_ctrl
		parameter hssi_8g_tx_pcs_eightb_tenb_encoder = "dis_8b10b", // dis_8b10b|en_8b10b_ibm|en_8b10b_sgx
		parameter hssi_8g_tx_pcs_force_echar = "dis_force_echar", // dis_force_echar|en_force_echar
		parameter hssi_8g_tx_pcs_force_kchar = "dis_force_kchar", // dis_force_kchar|en_force_kchar
		parameter hssi_8g_tx_pcs_gen3_tx_clk_sel = "tx_pma_clk", // dis_tx_clk|tx_pma_clk
		parameter hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel = "func_clk", // dis_tx_pipe_clk|func_clk
		parameter hssi_8g_tx_pcs_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_8g_tx_pcs_pcs_bypass = "dis_pcs_bypass", // dis_pcs_bypass|en_pcs_bypass
		parameter hssi_8g_tx_pcs_phase_comp_rdptr = "enable_rdptr", // disable_rdptr|enable_rdptr
		parameter hssi_8g_tx_pcs_phase_compensation_fifo = "low_latency", // low_latency|normal_latency|register_fifo|pld_ctrl_low_latency|pld_ctrl_normal_latency
		parameter hssi_8g_tx_pcs_phfifo_write_clk_sel = "pld_tx_clk", // pld_tx_clk|tx_clk
		parameter hssi_8g_tx_pcs_pma_dw = "eight_bit", // eight_bit|ten_bit|sixteen_bit|twenty_bit
		parameter hssi_8g_tx_pcs_prot_mode = "basic", // pipe_g1|pipe_g2|pipe_g3|cpri|cpri_rx_tx|gige|gige_1588|basic|disabled_prot_mode
		parameter hssi_8g_tx_pcs_reconfig_settings = "{}", // 
		parameter hssi_8g_tx_pcs_refclk_b_clk_sel = "tx_pma_clock", // tx_pma_clock|refclk_dig
		parameter hssi_8g_tx_pcs_revloop_back_rm = "dis_rev_loopback_rx_rm", // dis_rev_loopback_rx_rm|en_rev_loopback_rx_rm
		parameter hssi_8g_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_8g_tx_pcs_symbol_swap = "dis_symbol_swap", // dis_symbol_swap|en_symbol_swap
		parameter hssi_8g_tx_pcs_tx_bitslip = "dis_tx_bitslip", // dis_tx_bitslip|en_tx_bitslip
		parameter hssi_8g_tx_pcs_tx_compliance_controlled_disparity = "dis_txcompliance", // dis_txcompliance|en_txcompliance_pipe2p0|en_txcompliance_pipe3p0
		parameter hssi_8g_tx_pcs_tx_fast_pld_reg = "dis_tx_fast_pld_reg", // dis_tx_fast_pld_reg|en_tx_fast_pld_reg
		parameter hssi_8g_tx_pcs_txclk_freerun = "dis_freerun_tx", // dis_freerun_tx|en_freerun_tx
		parameter hssi_8g_tx_pcs_txpcs_urst = "en_txpcs_urst", // dis_txpcs_urst|en_txpcs_urst
		
		// parameters for twentynm_hssi_common_pcs_pma_interface
		parameter hssi_common_pcs_pma_interface_asn_clk_enable = "false", // false|true
		parameter hssi_common_pcs_pma_interface_asn_enable = "dis_asn", // dis_asn|en_asn
		parameter hssi_common_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|pcie_gen3
		parameter hssi_common_pcs_pma_interface_bypass_early_eios = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pcie_switch = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_ltr = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_pma_sw_done = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_ppm_lock = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp = "false", // false|true
		parameter hssi_common_pcs_pma_interface_bypass_txdetectrx = "false", // false|true
		parameter hssi_common_pcs_pma_interface_cdr_control = "en_cdr_ctrl", // dis_cdr_ctrl|en_cdr_ctrl
		parameter hssi_common_pcs_pma_interface_cid_enable = "en_cid_mode", // dis_cid_mode|en_cid_mode
		parameter hssi_common_pcs_pma_interface_cp_cons_sel = "cp_cons_default", // cp_cons_master|cp_cons_slave_abv|cp_cons_slave_blw|cp_cons_default
		parameter hssi_common_pcs_pma_interface_cp_dwn_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_cp_up_mstr = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_blw|ctrl_slave_abv
		parameter hssi_common_pcs_pma_interface_data_mask_count = 16'b100111000100,
		parameter hssi_common_pcs_pma_interface_data_mask_count_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_dft_observation_clock_selection = "dft_clk_obsrv_tx0", // dft_clk_obsrv_tx0|dft_clk_obsrv_tx1|dft_clk_obsrv_tx2|dft_clk_obsrv_tx3|dft_clk_obsrv_tx4|dft_clk_obsrv_rx|dft_clk_obsrv_hclk|dft_clk_obsrv_fref|dft_clk_obsrv_clklow|dft_clk_obsrv_asn0|dft_clk_obsrv_asn1
		parameter hssi_common_pcs_pma_interface_early_eios_counter = 8'b110010,
		parameter hssi_common_pcs_pma_interface_force_freqdet = "force_freqdet_dis", // force_freqdet_dis|force1_freqdet_en|force0_freqdet_en
		parameter hssi_common_pcs_pma_interface_free_run_clk_enable = "true", // false|true
		parameter hssi_common_pcs_pma_interface_ignore_sigdet_g23 = "false", // false|true
		parameter hssi_common_pcs_pma_interface_pc_en_counter = 7'b110111,
		parameter hssi_common_pcs_pma_interface_pc_rst_counter = 5'b10111,
		parameter hssi_common_pcs_pma_interface_pcie_hip_mode = "hip_disable", // hip_enable|hip_disable
		parameter hssi_common_pcs_pma_interface_ph_fifo_reg_mode = "phfifo_reg_mode_dis", // phfifo_reg_mode_dis|phfifo_reg_mode_en
		parameter hssi_common_pcs_pma_interface_phfifo_flush_wait = 6'b100100,
		parameter hssi_common_pcs_pma_interface_pipe_if_g3pcs = "pipe_if_8gpcs", // pipe_if_g3pcs|pipe_if_8gpcs
		parameter hssi_common_pcs_pma_interface_pma_done_counter = 18'b101010101110011000,
		parameter hssi_common_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_common_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_common_pcs_pma_interface_ppm_cnt_rst = "ppm_cnt_rst_dis", // ppm_cnt_rst_dis|ppm_cnt_rst_en
		parameter hssi_common_pcs_pma_interface_ppm_deassert_early = "deassert_early_dis", // deassert_early_dis|deassert_early_en
		parameter hssi_common_pcs_pma_interface_ppm_det_buckets = "ppm_100_bucket", // disable_prot|ppm_300_bucket|ppm_100_bucket|ppm_300_100_bucket
		parameter hssi_common_pcs_pma_interface_ppm_gen1_2_cnt = "cnt_32k", // cnt_32k|cnt_64k
		parameter hssi_common_pcs_pma_interface_ppm_post_eidle_delay = "cnt_200_cycles", // cnt_200_cycles|cnt_400_cycles
		parameter hssi_common_pcs_pma_interface_ppmsel = "ppmsel_300", // ppmsel_disable|ppmsel_5000|ppmsel_2500|ppmsel_1000|ppmsel_500|ppmsel_300|ppmsel_250|ppmsel_200|ppmsel_125|ppmsel_100|ppmsel_62p5|ppm_other
		parameter hssi_common_pcs_pma_interface_prot_mode = "disable_prot_mode", // disable_prot_mode|pipe_g12|pipe_g3|other_protocols
		parameter hssi_common_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_common_pcs_pma_interface_rxvalid_mask = "rxvalid_mask_en", // rxvalid_mask_dis|rxvalid_mask_en
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter = 12'b100111000100,
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter_multi = 3'b1,
		parameter hssi_common_pcs_pma_interface_sim_mode = "disable", // disable|enable
		parameter hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en = "true", // false|true
		parameter hssi_common_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_common_pcs_pma_interface_testout_sel = "ppm_det_test", // ppm_det_test|asn_test|pma_pll_test|rxpmaif_test|prbs_gen_test|prbs_ver_test|uhsif_1_test|uhsif_2_test|uhsif_3_test
		parameter hssi_common_pcs_pma_interface_wait_clk_on_off_timer = 4'b100,
		parameter hssi_common_pcs_pma_interface_wait_pipe_synchronizing = 5'b10111,
		parameter hssi_common_pcs_pma_interface_wait_send_syncp_fbkp = 11'b11111010,
		
		// parameters for twentynm_hssi_common_pld_pcs_interface
		parameter hssi_common_pld_pcs_interface_dft_clk_out_en = "dft_clk_out_disable", // dft_clk_out_disable|dft_clk_out_enable
		parameter hssi_common_pld_pcs_interface_dft_clk_out_sel = "teng_rx_dft_clk", // teng_rx_dft_clk|teng_tx_dft_clk|eightg_rx_dft_clk|eightg_tx_dft_clk|pmaif_dft_clk
		parameter hssi_common_pld_pcs_interface_hrdrstctrl_en = "hrst_dis", // hrst_dis|hrst_en
		parameter hssi_common_pld_pcs_interface_pcs_testbus_block_sel = "eightg", // eightg|g3pcs|teng|krfec|pma_if
		parameter hssi_common_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_fifo_rx_pcs
		parameter hssi_fifo_rx_pcs_double_read_mode = "double_read_dis", // double_read_en|double_read_dis
		parameter hssi_fifo_rx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_fifo_tx_pcs
		parameter hssi_fifo_tx_pcs_double_write_mode = "double_write_dis", // double_write_en|double_write_dis
		parameter hssi_fifo_tx_pcs_prot_mode = "teng_mode", // teng_mode|non_teng_mode
		
		// parameters for twentynm_hssi_gen3_rx_pcs
		parameter hssi_gen3_rx_pcs_block_sync = "enable_block_sync", // bypass_block_sync|enable_block_sync
		parameter hssi_gen3_rx_pcs_block_sync_sm = "enable_blk_sync_sm", // disable_blk_sync_sm|enable_blk_sync_sm
		parameter hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn = "enable", // disable|enable
		parameter hssi_gen3_rx_pcs_lpbk_force = "lpbk_frce_dis", // lpbk_frce_dis|lpbk_frce_en
		parameter hssi_gen3_rx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_rx_pcs_rate_match_fifo = "enable_rm_fifo_600ppm", // bypass_rm_fifo|enable_rm_fifo_600ppm|enable_rm_fifo_0ppm
		parameter hssi_gen3_rx_pcs_rate_match_fifo_latency = "regular_latency", // regular_latency|low_latency
		parameter hssi_gen3_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_gen3_rx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_b4gb_par_lpbk = "b4gb_par_lpbk_dis", // b4gb_par_lpbk_dis|b4gb_par_lpbk_en
		parameter hssi_gen3_rx_pcs_rx_force_balign = "en_force_balign", // en_force_balign|dis_force_balign
		parameter hssi_gen3_rx_pcs_rx_ins_del_one_skip = "ins_del_one_skip_en", // ins_del_one_skip_dis|ins_del_one_skip_en
		parameter hssi_gen3_rx_pcs_rx_num_fixed_pat = 4'b1000,
		parameter hssi_gen3_rx_pcs_rx_test_out_sel = "rx_test_out0", // rx_test_out0|rx_test_out1
		parameter hssi_gen3_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_gen3_tx_pcs
		parameter hssi_gen3_tx_pcs_mode = "gen3_func", // gen3_func|disable_pcs
		parameter hssi_gen3_tx_pcs_reverse_lpbk = "rev_lpbk_en", // rev_lpbk_dis|rev_lpbk_en
		parameter hssi_gen3_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_gen3_tx_pcs_tx_bitslip = 5'b0,
		parameter hssi_gen3_tx_pcs_tx_gbox_byp = "bypass_gbox", // bypass_gbox|enable_gbox
		
		// parameters for twentynm_hssi_krfec_rx_pcs
		parameter hssi_krfec_rx_pcs_blksync_cor_en = "detect", // detect|correct
		parameter hssi_krfec_rx_pcs_bypass_gb = "bypass_dis", // bypass_dis|bypass_en
		parameter hssi_krfec_rx_pcs_clr_ctrl = "both_enabled", // both_enabled|corr_cnt_only|uncorr_cnt_only
		parameter hssi_krfec_rx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_rx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_rx_pcs_dv_start = "with_blklock", // with_blksync|with_blklock
		parameter hssi_krfec_rx_pcs_err_mark_type = "err_mark_10g", // err_mark_10g|err_mark_40g
		parameter hssi_krfec_rx_pcs_error_marking_en = "err_mark_dis", // err_mark_dis|err_mark_en
		parameter hssi_krfec_rx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_rx_pcs_lpbk_mode = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_krfec_rx_pcs_parity_invalid_enum = 8'b1000,
		parameter hssi_krfec_rx_pcs_parity_valid_num = 4'b100,
		parameter hssi_krfec_rx_pcs_pipeln_blksync = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_descrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errcorrect = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_ind = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_lfsr = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_loc = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_pat = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_gearbox = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_syndrm = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_pipeln_trans_dec = "enable", // disable|enable
		parameter hssi_krfec_rx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_rx_pcs_receive_order = "receive_lsb", // receive_lsb|receive_msb
		parameter hssi_krfec_rx_pcs_reconfig_settings = "{}", // 
		parameter hssi_krfec_rx_pcs_rx_testbus_sel = "overall", // overall|fast_search|fast_search_cntrs|blksync|blksync_cntrs|decoder_master_sm|decoder_master_sm_cntrs|syndrm_sm|syndrm1|syndrm2|errtrap_sm|errtrap_ind1|errtrap_ind2|errtrap_ind3|errtrap_ind4|errtrap_ind5|errtrap_loc|errtrap_pat1|errtrap_pat2|errtrap_pat3|errtrap_pat4|decoder_rd_sm|gb_and_trans
		parameter hssi_krfec_rx_pcs_signal_ok_en = "sig_ok_dis", // sig_ok_dis|sig_ok_en
		parameter hssi_krfec_rx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_krfec_tx_pcs
		parameter hssi_krfec_tx_pcs_burst_err = "burst_err_dis", // burst_err_dis|burst_err_en
		parameter hssi_krfec_tx_pcs_burst_err_len = "burst_err_len1", // burst_err_len1|burst_err_len2|burst_err_len3|burst_err_len4|burst_err_len5|burst_err_len6|burst_err_len7|burst_err_len8|burst_err_len9|burst_err_len10|burst_err_len11|burst_err_len12|burst_err_len13|burst_err_len14|burst_err_len15|burst_err_len16
		parameter hssi_krfec_tx_pcs_ctrl_bit_reverse = "ctrl_bit_reverse_dis", // ctrl_bit_reverse_dis|ctrl_bit_reverse_en
		parameter hssi_krfec_tx_pcs_data_bit_reverse = "data_bit_reverse_dis", // data_bit_reverse_dis|data_bit_reverse_en
		parameter hssi_krfec_tx_pcs_enc_frame_query = "enc_query_dis", // enc_query_dis|enc_query_en
		parameter hssi_krfec_tx_pcs_low_latency_en = "disable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_encoder = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_pipeln_scrambler = "enable", // disable|enable
		parameter hssi_krfec_tx_pcs_prot_mode = "disable_mode", // disable_mode|teng_basekr_mode|fortyg_basekr_mode|teng_1588_basekr_mode|basic_mode
		parameter hssi_krfec_tx_pcs_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_krfec_tx_pcs_transcode_err = "trans_err_dis", // trans_err_dis|trans_err_en
		parameter hssi_krfec_tx_pcs_transmit_order = "transmit_lsb", // transmit_lsb|transmit_msb
		parameter hssi_krfec_tx_pcs_tx_testbus_sel = "overall", // overall|encoder1|encoder2|scramble1|scramble2|scramble3|gearbox
		
		// parameters for twentynm_hssi_pipe_gen1_2
		parameter hssi_pipe_gen1_2_elec_idle_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_error_replace_pad = "replace_edb", // replace_edb|replace_pad
		parameter hssi_pipe_gen1_2_hip_mode = "dis_hip", // dis_hip|en_hip
		parameter hssi_pipe_gen1_2_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen1_2_phystatus_delay_val = 3'b0,
		parameter hssi_pipe_gen1_2_phystatus_rst_toggle = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen1_2_pipe_byte_de_serializer_en = "dont_care_bds", // dis_bds|en_bds_by_2|dont_care_bds
		parameter hssi_pipe_gen1_2_prot_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|basic|disabled_prot_mode
		parameter hssi_pipe_gen1_2_reconfig_settings = "{}", // 
		parameter hssi_pipe_gen1_2_rx_pipe_enable = "dis_pipe_rx", // dis_pipe_rx|en_pipe_rx|en_pipe3_rx
		parameter hssi_pipe_gen1_2_rxdetect_bypass = "dis_rxdetect_bypass", // dis_rxdetect_bypass|en_rxdetect_bypass
		parameter hssi_pipe_gen1_2_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen1_2_tx_pipe_enable = "dis_pipe_tx", // dis_pipe_tx|en_pipe_tx|en_pipe3_tx
		parameter hssi_pipe_gen1_2_txswing = "dis_txswing", // dis_txswing|en_txswing
		
		// parameters for twentynm_hssi_pipe_gen3
		parameter hssi_pipe_gen3_bypass_rx_detection_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_rx_preset = 3'b0,
		parameter hssi_pipe_gen3_bypass_rx_preset_enable = "false", // false|true
		parameter hssi_pipe_gen3_bypass_tx_coefficent = 18'b0,
		parameter hssi_pipe_gen3_bypass_tx_coefficent_enable = "false", // false|true
		parameter hssi_pipe_gen3_elecidle_delay_g3 = 3'b110,
		parameter hssi_pipe_gen3_ind_error_reporting = "dis_ind_error_reporting", // dis_ind_error_reporting|en_ind_error_reporting
		parameter hssi_pipe_gen3_mode = "pipe_g1", // pipe_g1|pipe_g2|pipe_g3|disable_pcs
		parameter hssi_pipe_gen3_phy_status_delay_g12 = 3'b101,
		parameter hssi_pipe_gen3_phy_status_delay_g3 = 3'b101,
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g12 = "dis_phystatus_rst_toggle", // dis_phystatus_rst_toggle|en_phystatus_rst_toggle
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g3 = "dis_phystatus_rst_toggle_g3", // dis_phystatus_rst_toggle_g3|en_phystatus_rst_toggle_g3
		parameter hssi_pipe_gen3_rate_match_pad_insertion = "dis_rm_fifo_pad_ins", // dis_rm_fifo_pad_ins|en_rm_fifo_pad_ins
		parameter hssi_pipe_gen3_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_pipe_gen3_test_out_sel = "disable_test_out", // tx_test_out|rx_test_out|pipe_test_out1|pipe_test_out2|pipe_test_out3|pipe_ctrl_test_out|disable_test_out
		
		// parameters for twentynm_hssi_rx_pcs_pma_interface
		parameter hssi_rx_pcs_pma_interface_block_sel = "eight_g_pcs", // eight_g_pcs|ten_g_pcs|direct_pld
		parameter hssi_rx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pcs_pma_interface_clkslip_sel = "pld", // pld|slip_eight_g_pcs
		parameter hssi_rx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pcs_pma_interface_master_clk_sel = "master_rx_pma_clk", // master_rx_pma_clk|master_tx_pma_clk|master_refclk_dig
		parameter hssi_rx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_rx_pcs_pma_interface_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_val = "dft_0", // dft_0|dft_1
		parameter hssi_rx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_rx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_rx_pcs_pma_interface_prbs_ver = "prbs_off", // prbs_off|prbs_31|prbs_15|prbs_23|prbs_9|prbs_7
		parameter hssi_rx_pcs_pma_interface_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion = "rx_dyn_polinv_dis", // rx_dyn_polinv_dis|rx_dyn_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_lpbk_en = "lpbk_dis", // lpbk_dis|lpbk_en
		parameter hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok = "unforce_sig_ok", // unforce_sig_ok|force_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mask = "prbsmask128", // prbsmask128|prbsmask256|prbsmask512|prbsmask1024
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mode = "teng_mode", // teng_mode|eightg_mode
		parameter hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel = "sel_sig_det", // sel_sig_det|sel_sig_ok
		parameter hssi_rx_pcs_pma_interface_rx_static_polarity_inversion = "rx_stat_polinv_dis", // rx_stat_polinv_dis|rx_stat_polinv_en
		parameter hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en = "uhsif_lpbk_dis", // uhsif_lpbk_dis|uhsif_lpbk_en
		parameter hssi_rx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		
		// parameters for twentynm_hssi_rx_pld_pcs_interface
		parameter hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx = "enable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx = "pma_64b_rx", // pma_32b_rx|pma_40b_rx|pma_64b_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_baser_mode_rx|interlaken_mode_rx|sfis_mode_rx|teng_sdi_mode_rx|basic_mode_rx|test_prp_mode_rx|test_prp_krfec_mode_rx|teng_1588_mode_rx|teng_baser_krfec_mode_rx|teng_1588_krfec_mode_rx|basic_krfec_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx
		parameter hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx = "disabled_prot_mode_rx", // pipe_g1_rx|pipe_g2_rx|pipe_g3_rx|cpri_rx|cpri_rx_tx_rx|gige_rx|gige_1588_rx|basic_rm_enable_rx|basic_rm_disable_rx|disabled_prot_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx = "individual_rx", // individual_rx|ctrl_master_rx|ctrl_slave_abv_rx|ctrl_slave_blw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx = "fifo_rx", // fifo_rx|reg_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz = 30'b0,
		parameter hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcie_g1_capable_rx|pcie_g2_capable_rx|pcie_g3_capable_rx|gige_rx|teng_baser_rx|teng_basekr_krfec_rx|fortyg_basekr_krfec_rx|cpri_8b10b_rx|interlaken_rx|sfis_rx|teng_sdi_rx|gige_1588_rx|teng_1588_baser_rx|teng_1588_basekr_krfec_rx|basic_8gpcs_rm_enable_rx|basic_8gpcs_rm_disable_rx|basic_10gpcs_rx|basic_10gpcs_krfec_rx|pcs_direct_rx|prp_rx|prp_krfec_rx|prbs_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx = "teng_mode_rx", // teng_mode_rx|non_teng_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx = "single_rx", // single_rx|double_rx
		parameter hssi_rx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|teng_basekr_mode_rx|fortyg_basekr_mode_rx|teng_1588_basekr_mode_rx|basic_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode = "tx", // tx|rx
		parameter hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|eightg_and_g3_pld_fifo_mode_rx|eightg_and_g3_reg_mode_rx|eightg_and_g3_reg_mode_hip_rx|teng_pld_fifo_mode_rx|teng_reg_mode_rx|teng_and_krfec_pld_fifo_mode_rx|teng_and_krfec_reg_mode_rx|pcs_direct_reg_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx = "pma_8b_rx", // pma_8b_rx|pma_10b_rx|pma_16b_rx|pma_20b_rx|pma_32b_rx|pma_40b_rx|pma_64b_rx|pcie_g3_dyn_dw_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx = "disabled_prot_mode_rx", // disabled_prot_mode_rx|pcs_direct_mode_rx|eightg_only_pld_mode_rx|eightg_pcie_g12_pld_mode_rx|eightg_g3_pcie_g3_pld_mode_rx|eightg_pcie_g12_hip_mode_rx|eightg_g3_pcie_g3_hip_mode_rx|teng_krfec_mode_rx|eightg_basic_mode_rx|teng_basic_mode_rx|teng_sfis_sdi_mode_rx|prbs_mode_rx
		parameter hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_block_sel = "pcs_direct", // eightg|teng|pcs_direct
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_rx_clk|pma_rx_clk_user
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_sel = "pld_rx_clk", // pld_rx_clk|pcs_rx_clk
		parameter hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en = "hip_rx_enable", // hip_rx_enable|hip_rx_disable
		parameter hssi_rx_pld_pcs_interface_pcs_rx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_rx_pld_pcs_interface_reconfig_settings = "{}", // 
		
		// parameters for twentynm_hssi_tx_pcs_pma_interface
		parameter hssi_tx_pcs_pma_interface_bypass_pma_txelecidle = "false", // false|true
		parameter hssi_tx_pcs_pma_interface_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pcs_pma_interface_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pcs_pma_interface_master_clk_sel = "master_tx_pma_clk", // master_tx_pma_clk|master_refclk_dig
		parameter hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx = "other_prot_mode", // pipe_g12|pipe_g3|other_prot_mode
		parameter hssi_tx_pcs_pma_interface_pldif_datawidth_mode = "pldif_data_10bit", // pldif_data_10bit|pldif_data_8bit
		parameter hssi_tx_pcs_pma_interface_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pcs_pma_interface_pma_if_dft_en = "dft_dis", // dft_dis|dft_en
		parameter hssi_tx_pcs_pma_interface_pmagate_en = "pmagate_dis", // pmagate_dis|pmagate_en
		parameter hssi_tx_pcs_pma_interface_prbs9_dwidth = "prbs9_64b", // prbs9_64b|prbs9_10b
		parameter hssi_tx_pcs_pma_interface_prbs_clken = "prbs_clk_dis", // prbs_clk_dis|prbs_clk_en
		parameter hssi_tx_pcs_pma_interface_prbs_gen_pat = "prbs_gen_dis", // prbs_gen_dis|prbs_31|prbs_23|prbs_15|prbs_9|prbs_7
		parameter hssi_tx_pcs_pma_interface_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pcs_pma_interface_reconfig_settings = "{}", // 
		parameter hssi_tx_pcs_pma_interface_sq_wave_num = "sq_wave_4", // sq_wave_1|sq_wave_4|sq_wave_8|sq_wave_6|sq_wave_default
		parameter hssi_tx_pcs_pma_interface_sqwgen_clken = "sqwgen_clk_dis", // sqwgen_clk_dis|sqwgen_clk_en
		parameter hssi_tx_pcs_pma_interface_sup_mode = "user_mode", // user_mode|engineering_mode
		parameter hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion = "tx_dyn_polinv_dis", // tx_dyn_polinv_dis|tx_dyn_polinv_en
		parameter hssi_tx_pcs_pma_interface_tx_pma_data_sel = "pld_dir", // pld_dir|pcie_gen3|eight_g_pcs|ten_g_pcs|prbs_pat|sq_wave_pat|block_sel_default|registered_uhsif_dat|directed_uhsif_dat
		parameter hssi_tx_pcs_pma_interface_tx_static_polarity_inversion = "tx_stat_polinv_dis", // tx_stat_polinv_dis|tx_stat_polinv_en
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock = "uhsif_filt_stepsz_b4lock_4", // uhsif_filt_stepsz_b4lock_2|uhsif_filt_stepsz_b4lock_4|uhsif_filt_stepsz_b4lock_6|uhsif_filt_stepsz_b4lock_8
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value = 4'b1011,
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock = "uhsif_filt_cntthr_b4lock_16", // uhsif_filt_cntthr_b4lock_8|uhsif_filt_cntthr_b4lock_16|uhsif_filt_cntthr_b4lock_24|uhsif_filt_cntthr_b4lock_32
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period = "uhsif_dcn_test_period_4", // uhsif_dcn_test_period_4|uhsif_dcn_test_period_8|uhsif_dcn_test_period_12|uhsif_dcn_test_period_16
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable = "uhsif_dcn_test_mode_disable", // uhsif_dcn_test_mode_enable|uhsif_dcn_test_mode_disable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh = "uhsif_dzt_cnt_thr_4", // uhsif_dzt_cnt_thr_2|uhsif_dzt_cnt_thr_4|uhsif_dzt_cnt_thr_6|uhsif_dzt_cnt_thr_8
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable = "uhsif_dzt_enable", // uhsif_dzt_disable|uhsif_dzt_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window = "uhsif_dzt_obr_win_32", // uhsif_dzt_obr_win_16|uhsif_dzt_obr_win_32|uhsif_dzt_obr_win_48|uhsif_dzt_obr_win_64
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size = "uhsif_dzt_skipsz_8", // uhsif_dzt_skipsz_4|uhsif_dzt_skipsz_8|uhsif_dzt_skipsz_12|uhsif_dzt_skipsz_16
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel = "uhsif_index_internal", // uhsif_index_internal|uhsif_index_cram
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin = "uhsif_dcn_margin_4", // uhsif_dcn_margin_2|uhsif_dcn_margin_3|uhsif_dcn_margin_4|uhsif_dcn_margin_5
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value = 8'b10000000,
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control = "uhsif_dft_dz_det_val_0", // uhsif_dft_dz_det_val_0|uhsif_dft_dz_det_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control = "uhsif_dft_up_val_0", // uhsif_dft_up_val_0|uhsif_dft_up_val_1
		parameter hssi_tx_pcs_pma_interface_uhsif_enable = "uhsif_disable", // uhsif_disable|uhsif_enable
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock = "uhsif_lkd_segsz_aflock_2048", // uhsif_lkd_segsz_aflock_512|uhsif_lkd_segsz_aflock_1024|uhsif_lkd_segsz_aflock_2048|uhsif_lkd_segsz_aflock_4096
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock = "uhsif_lkd_segsz_b4lock_32", // uhsif_lkd_segsz_b4lock_16|uhsif_lkd_segsz_b4lock_32|uhsif_lkd_segsz_b4lock_64|uhsif_lkd_segsz_b4lock_128
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value = 4'b1000,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value = 4'b11,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value = 4'b11,
		
		// parameters for twentynm_hssi_tx_pld_pcs_interface
		parameter hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx = "enable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx = "pma_64b_tx", // pma_32b_tx|pma_40b_tx|pma_64b_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_baser_mode_tx|interlaken_mode_tx|sfis_mode_tx|teng_sdi_mode_tx|basic_mode_tx|test_prp_mode_tx|test_prp_krfec_mode_tx|teng_1588_mode_tx|teng_baser_krfec_mode_tx|teng_1588_krfec_mode_tx|basic_krfec_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_hip_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx
		parameter hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx = "disabled_prot_mode_tx", // pipe_g1_tx|pipe_g2_tx|pipe_g3_tx|cpri_tx|cpri_rx_tx_tx|gige_tx|gige_1588_tx|basic_tx|disabled_prot_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx = "individual_tx", // individual_tx|ctrl_master_tx|ctrl_slave_abv_tx|ctrl_slave_blw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_func_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hip_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx = "fifo_tx", // fifo_tx|reg_tx|fastreg_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz = 30'b0,
		parameter hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcie_g1_capable_tx|pcie_g2_capable_tx|pcie_g3_capable_tx|gige_tx|teng_baser_tx|teng_basekr_krfec_tx|fortyg_basekr_krfec_tx|cpri_8b10b_tx|interlaken_tx|sfis_tx|teng_sdi_tx|gige_1588_tx|teng_1588_baser_tx|teng_1588_basekr_krfec_tx|basic_8gpcs_tx|basic_10gpcs_tx|basic_10gpcs_krfec_tx|pcs_direct_tx|uhsif_tx|prp_tx|prp_krfec_tx|prbs_tx|sqwave_tx
		parameter hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx = "teng_mode_tx", // teng_mode_tx|non_teng_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx = "single_tx", // single_tx|double_tx
		parameter hssi_tx_pld_pcs_interface_hd_g3_prot_mode = "disabled_prot_mode", // pipe_g1|pipe_g2|pipe_g3|disabled_prot_mode
		parameter hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|teng_basekr_mode_tx|fortyg_basekr_mode_tx|teng_1588_basekr_mode_tx|basic_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|eightg_and_g3_pld_fifo_mode_tx|eightg_and_g3_reg_mode_tx|eightg_and_g3_reg_mode_hip_tx|eightg_and_g3_fastreg_mode_tx|teng_pld_fifo_mode_tx|teng_reg_mode_tx|teng_fastreg_mode_tx|teng_and_krfec_pld_fifo_mode_tx|teng_and_krfec_reg_mode_tx|teng_and_krfec_fastreg_mode_tx|pcs_direct_fastreg_mode_tx|uhsif_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled", // tx_rx_pair_enabled|tx_rx_independent
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding = "individual", // individual|ctrl_master|ctrl_slave_abv|ctrl_slave_blw
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx = "pma_8b_tx", // pma_8b_tx|pma_10b_tx|pma_16b_tx|pma_20b_tx|pma_32b_tx|pma_40b_tx|pma_64b_tx|pcie_g3_dyn_dw_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx = "disabled_prot_mode_tx", // disabled_prot_mode_tx|pcs_direct_mode_tx|uhsif_reg_mode_tx|uhsif_direct_mode_tx|eightg_only_pld_mode_tx|eightg_pcie_g12_pld_mode_tx|eightg_g3_pcie_g3_pld_mode_tx|eightg_pcie_g12_hip_mode_tx|eightg_g3_pcie_g3_hip_mode_tx|teng_krfec_mode_tx|eightg_basic_mode_tx|teng_basic_mode_tx|teng_sfis_sdi_mode_tx|prbs_mode_tx|sqwave_mode_tx
		parameter hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode = "disable", // disable|enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel = "teng_clk_out", // eightg_clk_out|teng_clk_out|pma_tx_clk|pma_tx_clk_user
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_source = "teng", // eightg|teng|pma_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_data_source = "hip_disable", // hip_disable|hip_enable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en = "delay1_clk_disable", // delay1_clk_enable|delay1_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel = "pld_tx_clk", // pld_tx_clk|pcs_tx_clk
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl = "delay1_path0", // delay1_path0|delay1_path1|delay1_path2|delay1_path3|delay1_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel = "one_ff_delay", // one_ff_delay|two_ff_delay
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en = "delay2_clk_disable", // delay2_clk_enable|delay2_clk_disable
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl = "delay2_path0", // delay2_path0|delay2_path1|delay2_path2|delay2_path3|delay2_path4
		parameter hssi_tx_pld_pcs_interface_pcs_tx_output_sel = "teng_output", // krfec_output|teng_output
		parameter hssi_tx_pld_pcs_interface_reconfig_settings = "{}" // 
	//PARAM_LIST_END
	)
	(
	//PORT_LIST_START
		input wire	[8:0]	in_avmmaddress,
		input wire		in_avmmclk,
		input wire		in_avmmread,
		input wire		in_avmmrstn,
		input wire		in_avmmwrite,
		input wire	[7:0]	in_avmmwritedata,
		input wire	[4:0]	in_bond_pcs10g_in_bot,
		input wire	[4:0]	in_bond_pcs10g_in_top,
		input wire	[12:0]	in_bond_pcs8g_in_bot,
		input wire	[12:0]	in_bond_pcs8g_in_top,
		input wire	[11:0]	in_bond_pmaif_in_bot,
		input wire	[11:0]	in_bond_pmaif_in_top,
		input wire	[63:0]	in_hip_tx_data,
		input wire		in_iocsr_clk,
		input wire	[5:0]	in_iocsr_config,
		input wire		in_iocsr_rdy,
		input wire		in_iocsr_rdy_dly,
		input wire		in_pld_10g_krfec_rx_clr_errblk_cnt,
		input wire		in_pld_10g_krfec_rx_pld_rst_n,
		input wire		in_pld_10g_krfec_tx_pld_rst_n,
		input wire		in_pld_10g_rx_align_clr,
		input wire		in_pld_10g_rx_clr_ber_count,
		input wire		in_pld_10g_rx_rd_en,
		input wire	[6:0]	in_pld_10g_tx_bitslip,
		input wire		in_pld_10g_tx_burst_en,
		input wire		in_pld_10g_tx_data_valid,
		input wire	[1:0]	in_pld_10g_tx_diag_status,
		input wire		in_pld_10g_tx_wordslip,
		input wire		in_pld_8g_a1a2_size,
		input wire		in_pld_8g_bitloc_rev_en,
		input wire		in_pld_8g_byte_rev_en,
		input wire	[2:0]	in_pld_8g_eidleinfersel,
		input wire		in_pld_8g_encdt,
		input wire		in_pld_8g_g3_rx_pld_rst_n,
		input wire		in_pld_8g_g3_tx_pld_rst_n,
		input wire		in_pld_8g_rddisable_tx,
		input wire		in_pld_8g_rdenable_rx,
		input wire		in_pld_8g_refclk_dig2,
		input wire		in_pld_8g_rxpolarity,
		input wire	[4:0]	in_pld_8g_tx_boundary_sel,
		input wire		in_pld_8g_wrdisable_rx,
		input wire		in_pld_8g_wrenable_tx,
		input wire		in_pld_atpg_los_en_n,
		input wire		in_pld_bitslip,
		input wire	[17:0]	in_pld_g3_current_coeff,
		input wire	[2:0]	in_pld_g3_current_rxpreset,
		input wire		in_pld_ltr,
		input wire		in_pld_mem_krfec_atpg_rst_n,
		input wire		in_pld_partial_reconfig,
		input wire		in_pld_pcs_refclk_dig,
		input wire		in_pld_pma_adapt_start,
		input wire		in_pld_pma_csr_test_dis,
		input wire		in_pld_pma_early_eios,
		input wire	[5:0]	in_pld_pma_eye_monitor,
		input wire		in_pld_pma_ltd_b,
		input wire		in_pld_pma_nrpi_freeze,
		input wire	[1:0]	in_pld_pma_pcie_switch,
		input wire		in_pld_pma_ppm_lock,
		input wire	[4:0]	in_pld_pma_reserved_out,
		input wire		in_pld_pma_rs_lpbk_b,
		input wire		in_pld_pma_rx_qpi_pullup,
		input wire		in_pld_pma_rxpma_rstb,
		input wire		in_pld_pma_tx_bitslip,
		input wire		in_pld_pma_tx_bonding_rstb,
		input wire		in_pld_pma_tx_qpi_pulldn,
		input wire		in_pld_pma_tx_qpi_pullup,
		input wire		in_pld_pma_txdetectrx,
		input wire		in_pld_pma_txpma_rstb,
		input wire		in_pld_pmaif_rx_pld_rst_n,
		input wire		in_pld_pmaif_rxclkslip,
		input wire		in_pld_pmaif_tx_pld_rst_n,
		input wire		in_pld_polinv_rx,
		input wire		in_pld_polinv_tx,
		input wire	[1:0]	in_pld_rate,
		input wire	[9:0]	in_pld_reserved_in,
		input wire		in_pld_rx_clk,
		input wire		in_pld_rx_prbs_err_clr,
		input wire		in_pld_scan_mode_n,
		input wire		in_pld_scan_shift_n,
		input wire		in_pld_syncsm_en,
		input wire		in_pld_tx_clk,
		input wire	[17:0]	in_pld_tx_control,
		input wire	[127:0]	in_pld_tx_data,
		input wire		in_pld_txelecidle,
		input wire		in_pld_uhsif_tx_clk,
		input wire		in_pma_adapt_done,
		input wire		in_pma_clklow,
		input wire		in_pma_fref,
		input wire		in_pma_hclk,
		input wire	[1:0]	in_pma_pcie_sw_done,
		input wire		in_pma_pfdmode_lock,
		input wire	[4:0]	in_pma_reserved_in,
		input wire		in_pma_rx_clkdiv_user,
		input wire		in_pma_rx_detect_valid,
		input wire		in_pma_rx_found,
		input wire		in_pma_rx_pma_clk,
		input wire	[63:0]	in_pma_rx_pma_data,
		input wire		in_pma_rx_signal_ok,
		input wire		in_pma_rxpll_lock,
		input wire		in_pma_signal_det,
		input wire	[7:0]	in_pma_testbus,
		input wire		in_pma_tx_clkdiv_user,
		input wire		in_pma_tx_pma_clk,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_10g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_8g_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_common_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_fifo_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_gen3_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_rx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_krfec_tx_pcs,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen1_2,
		output wire	[7:0]	out_avmmreaddata_hssi_pipe_gen3,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_rx_pld_pcs_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pcs_pma_interface,
		output wire	[7:0]	out_avmmreaddata_hssi_tx_pld_pcs_interface,
		output wire		out_blockselect_hssi_10g_rx_pcs,
		output wire		out_blockselect_hssi_10g_tx_pcs,
		output wire		out_blockselect_hssi_8g_rx_pcs,
		output wire		out_blockselect_hssi_8g_tx_pcs,
		output wire		out_blockselect_hssi_common_pcs_pma_interface,
		output wire		out_blockselect_hssi_common_pld_pcs_interface,
		output wire		out_blockselect_hssi_fifo_rx_pcs,
		output wire		out_blockselect_hssi_fifo_tx_pcs,
		output wire		out_blockselect_hssi_gen3_rx_pcs,
		output wire		out_blockselect_hssi_gen3_tx_pcs,
		output wire		out_blockselect_hssi_krfec_rx_pcs,
		output wire		out_blockselect_hssi_krfec_tx_pcs,
		output wire		out_blockselect_hssi_pipe_gen1_2,
		output wire		out_blockselect_hssi_pipe_gen3,
		output wire		out_blockselect_hssi_rx_pcs_pma_interface,
		output wire		out_blockselect_hssi_rx_pld_pcs_interface,
		output wire		out_blockselect_hssi_tx_pcs_pma_interface,
		output wire		out_blockselect_hssi_tx_pld_pcs_interface,
		output wire	[4:0]	out_bond_pcs10g_out_bot,
		output wire	[4:0]	out_bond_pcs10g_out_top,
		output wire	[12:0]	out_bond_pcs8g_out_bot,
		output wire	[12:0]	out_bond_pcs8g_out_top,
		output wire	[11:0]	out_bond_pmaif_out_bot,
		output wire	[11:0]	out_bond_pmaif_out_top,
		output wire	[2:0]	out_hip_clk_out,
		output wire	[7:0]	out_hip_ctrl_out,
		output wire		out_hip_iocsr_rdy,
		output wire		out_hip_iocsr_rdy_dly,
		output wire		out_hip_nfrzdrv,
		output wire		out_hip_npor,
		output wire	[50:0]	out_hip_rx_data,
		output wire		out_hip_usermode,
		output wire		out_pld_10g_krfec_rx_blk_lock,
		output wire	[1:0]	out_pld_10g_krfec_rx_diag_data_status,
		output wire		out_pld_10g_krfec_rx_frame,
		output wire		out_pld_10g_krfec_tx_frame,
		output wire		out_pld_10g_rx_align_val,
		output wire		out_pld_10g_rx_crc32_err,
		output wire		out_pld_10g_rx_data_valid,
		output wire		out_pld_10g_rx_empty,
		output wire		out_pld_10g_rx_fifo_del,
		output wire		out_pld_10g_rx_fifo_insert,
		output wire	[4:0]	out_pld_10g_rx_fifo_num,
		output wire		out_pld_10g_rx_frame_lock,
		output wire		out_pld_10g_rx_hi_ber,
		output wire		out_pld_10g_rx_oflw_err,
		output wire		out_pld_10g_rx_pempty,
		output wire		out_pld_10g_rx_pfull,
		output wire		out_pld_10g_tx_burst_en_exe,
		output wire		out_pld_10g_tx_empty,
		output wire	[3:0]	out_pld_10g_tx_fifo_num,
		output wire		out_pld_10g_tx_full,
		output wire		out_pld_10g_tx_pempty,
		output wire		out_pld_10g_tx_pfull,
		output wire		out_pld_10g_tx_wordslip_exe,
		output wire	[3:0]	out_pld_8g_a1a2_k1k2_flag,
		output wire		out_pld_8g_empty_rmf,
		output wire		out_pld_8g_empty_rx,
		output wire		out_pld_8g_empty_tx,
		output wire		out_pld_8g_full_rmf,
		output wire		out_pld_8g_full_rx,
		output wire		out_pld_8g_full_tx,
		output wire		out_pld_8g_rxelecidle,
		output wire		out_pld_8g_signal_detect_out,
		output wire	[4:0]	out_pld_8g_wa_boundary,
		output wire		out_pld_krfec_tx_alignment,
		output wire		out_pld_pcs_rx_clk_out,
		output wire		out_pld_pcs_tx_clk_out,
		output wire		out_pld_pma_adapt_done,
		output wire		out_pld_pma_clkdiv_rx_user,
		output wire		out_pld_pma_clkdiv_tx_user,
		output wire		out_pld_pma_clklow,
		output wire		out_pld_pma_fref,
		output wire		out_pld_pma_hclk,
		output wire	[1:0]	out_pld_pma_pcie_sw_done,
		output wire		out_pld_pma_pfdmode_lock,
		output wire	[4:0]	out_pld_pma_reserved_in,
		output wire		out_pld_pma_rx_clk_out,
		output wire		out_pld_pma_rx_detect_valid,
		output wire		out_pld_pma_rx_found,
		output wire		out_pld_pma_rxpll_lock,
		output wire		out_pld_pma_signal_ok,
		output wire	[7:0]	out_pld_pma_testbus,
		output wire		out_pld_pma_tx_clk_out,
		output wire		out_pld_pmaif_mask_tx_pll,
		output wire	[9:0]	out_pld_reserved_out,
		output wire	[19:0]	out_pld_rx_control,
		output wire	[127:0]	out_pld_rx_data,
		output wire		out_pld_rx_prbs_done,
		output wire		out_pld_rx_prbs_err,
		output wire	[19:0]	out_pld_test_data,
		output wire		out_pld_uhsif_lock,
		output wire		out_pld_uhsif_tx_clk_out,
		output wire		out_pma_adapt_start,
		output wire		out_pma_atpg_los_en_n,
		output wire		out_pma_csr_test_dis,
		output wire	[17:0]	out_pma_current_coeff,
		output wire	[2:0]	out_pma_current_rxpreset,
		output wire		out_pma_early_eios,
		output wire	[5:0]	out_pma_eye_monitor,
		output wire	[1:0]	out_pma_interface_select,
		output wire		out_pma_ltd_b,
		output wire		out_pma_ltr,
		output wire		out_pma_nfrzdrv,
		output wire		out_pma_nrpi_freeze,
		output wire	[1:0]	out_pma_pcie_switch,
		output wire		out_pma_ppm_lock,
		output wire	[4:0]	out_pma_reserved_out,
		output wire		out_pma_rs_lpbk_b,
		output wire		out_pma_rx_clkslip,
		output wire		out_pma_rx_qpi_pullup,
		output wire		out_pma_rxpma_rstb,
		output wire		out_pma_scan_mode_n,
		output wire		out_pma_scan_shift_n,
		output wire		out_pma_tx_bitslip,
		output wire		out_pma_tx_bonding_rstb,
		output wire		out_pma_tx_elec_idle,
		output wire	[63:0]	out_pma_tx_pma_data,
		output wire		out_pma_tx_qpi_pulldn,
		output wire		out_pma_tx_qpi_pullup,
		output wire		out_pma_tx_txdetectrx,
		output wire		out_pma_txpma_rstb
	//PORT_LIST_END
	);
	//wire declarations
	
	// wires for module twentynm_hssi_fifo_tx_pcs
	wire	[7:0]	w_hssi_fifo_tx_pcs_avmmreaddata;
	wire		w_hssi_fifo_tx_pcs_blockselect;
	wire	[72:0]	w_hssi_fifo_tx_pcs_data_out_10g;
	wire	[63:0]	w_hssi_fifo_tx_pcs_data_out_8g_phase_comp;
	
	// wires for module twentynm_hssi_gen3_rx_pcs
	wire	[7:0]	w_hssi_gen3_rx_pcs_avmmreaddata;
	wire		w_hssi_gen3_rx_pcs_blk_algnd_int;
	wire		w_hssi_gen3_rx_pcs_blk_start;
	wire		w_hssi_gen3_rx_pcs_blockselect;
	wire		w_hssi_gen3_rx_pcs_clkcomp_delete_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_insert_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_overfl_int;
	wire		w_hssi_gen3_rx_pcs_clkcomp_undfl_int;
	wire	[31:0]	w_hssi_gen3_rx_pcs_data_out;
	wire		w_hssi_gen3_rx_pcs_data_valid;
	wire		w_hssi_gen3_rx_pcs_ei_det_int;
	wire		w_hssi_gen3_rx_pcs_ei_partial_det_int;
	wire		w_hssi_gen3_rx_pcs_err_decode_int;
	wire		w_hssi_gen3_rx_pcs_i_det_int;
	wire		w_hssi_gen3_rx_pcs_lpbk_blk_start;
	wire	[33:0]	w_hssi_gen3_rx_pcs_lpbk_data;
	wire		w_hssi_gen3_rx_pcs_lpbk_data_valid;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk;
	wire	[39:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en;
	wire	[15:0]	w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr;
	wire		w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n;
	wire		w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int;
	wire	[19:0]	w_hssi_gen3_rx_pcs_rx_test_out;
	wire	[1:0]	w_hssi_gen3_rx_pcs_sync_hdr;
	
	// wires for module twentynm_hssi_krfec_tx_pcs
	wire	[7:0]	w_hssi_krfec_tx_pcs_avmmreaddata;
	wire		w_hssi_krfec_tx_pcs_blockselect;
	wire		w_hssi_krfec_tx_pcs_tx_alignment;
	wire	[63:0]	w_hssi_krfec_tx_pcs_tx_data_out;
	wire		w_hssi_krfec_tx_pcs_tx_frame;
	wire	[19:0]	w_hssi_krfec_tx_pcs_tx_test_data;
	
	// wires for module twentynm_hssi_krfec_rx_pcs
	wire	[7:0]	w_hssi_krfec_rx_pcs_avmmreaddata;
	wire		w_hssi_krfec_rx_pcs_blockselect;
	wire		w_hssi_krfec_rx_pcs_rx_block_lock;
	wire	[9:0]	w_hssi_krfec_rx_pcs_rx_control_out;
	wire	[63:0]	w_hssi_krfec_rx_pcs_rx_data_out;
	wire	[1:0]	w_hssi_krfec_rx_pcs_rx_data_status;
	wire		w_hssi_krfec_rx_pcs_rx_data_valid_out;
	wire		w_hssi_krfec_rx_pcs_rx_frame;
	wire		w_hssi_krfec_rx_pcs_rx_signal_ok_out;
	
	// wires for module twentynm_hssi_rx_pld_pcs_interface
	wire	[7:0]	w_hssi_rx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_rx_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_hip_rx_ctrl;
	wire	[50:0]	w_hssi_rx_pld_pcs_interface_hip_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr;
	wire		w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
	wire	[1:0]	w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
	wire		w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
	wire	[3:0]	w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
	wire		w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
	wire	[4:0]	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary;
	wire		w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
	wire		w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
	wire	[19:0]	w_hssi_rx_pld_pcs_interface_pld_rx_control;
	wire	[127:0]	w_hssi_rx_pld_pcs_interface_pld_rx_data;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
	wire		w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
	
	// wires for module twentynm_hssi_common_pld_pcs_interface
	wire	[7:0]	w_hssi_common_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_common_pld_pcs_interface_blockselect;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_hip_cmn_clk;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_hip_cmn_ctrl;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
	wire		w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
	wire		w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_hip_npor;
	wire		w_hssi_common_pld_pcs_interface_hip_usermode;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n;
	wire	[17:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff;
	wire	[2:0]	w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios;
	wire	[5:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig;
	wire		w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel;
	wire		w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_clklow;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_fref;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_hclk;
	wire	[1:0]	w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
	wire	[4:0]	w_hssi_common_pld_pcs_interface_pld_pma_reserved_in;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
	wire		w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
	wire	[7:0]	w_hssi_common_pld_pcs_interface_pld_pma_testbus;
	wire		w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
	wire	[9:0]	w_hssi_common_pld_pcs_interface_pld_reserved_out;
	wire	[19:0]	w_hssi_common_pld_pcs_interface_pld_test_data;
	wire		w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
	wire		w_hssi_common_pld_pcs_interface_scan_mode_n;
	
	// wires for module twentynm_hssi_10g_rx_pcs
	wire	[7:0]	w_hssi_10g_rx_pcs_avmmreaddata;
	wire		w_hssi_10g_rx_pcs_blockselect;
	wire		w_hssi_10g_rx_pcs_rx_align_val;
	wire		w_hssi_10g_rx_pcs_rx_blk_lock;
	wire		w_hssi_10g_rx_pcs_rx_clk_out;
	wire		w_hssi_10g_rx_pcs_rx_clk_out_pld_if;
	wire	[19:0]	w_hssi_10g_rx_pcs_rx_control;
	wire		w_hssi_10g_rx_pcs_rx_crc32_err;
	wire	[127:0]	w_hssi_10g_rx_pcs_rx_data;
	wire		w_hssi_10g_rx_pcs_rx_data_valid;
	wire		w_hssi_10g_rx_pcs_rx_dft_clk_out;
	wire	[1:0]	w_hssi_10g_rx_pcs_rx_diag_status;
	wire		w_hssi_10g_rx_pcs_rx_empty;
	wire		w_hssi_10g_rx_pcs_rx_fec_clk;
	wire		w_hssi_10g_rx_pcs_rx_fifo_del;
	wire		w_hssi_10g_rx_pcs_rx_fifo_insert;
	wire	[4:0]	w_hssi_10g_rx_pcs_rx_fifo_num;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_clk;
	wire	[73:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_data;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_en;
	wire	[31:0]	w_hssi_10g_rx_pcs_rx_fifo_wr_ptr;
	wire		w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_frame_lock;
	wire		w_hssi_10g_rx_pcs_rx_hi_ber;
	wire		w_hssi_10g_rx_pcs_rx_master_clk;
	wire		w_hssi_10g_rx_pcs_rx_master_clk_rst_n;
	wire		w_hssi_10g_rx_pcs_rx_oflw_err;
	wire		w_hssi_10g_rx_pcs_rx_pempty;
	wire		w_hssi_10g_rx_pcs_rx_pfull;
	wire		w_hssi_10g_rx_pcs_rx_random_err;
	wire		w_hssi_10g_rx_pcs_rx_rx_frame;
	
	// wires for module twentynm_hssi_tx_pld_pcs_interface
	wire	[7:0]	w_hssi_tx_pld_pcs_interface_avmmreaddata;
	wire		w_hssi_tx_pld_pcs_interface_blockselect;
	wire		w_hssi_tx_pld_pcs_interface_hip_tx_clk;
	wire	[6:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en;
	wire	[17:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control;
	wire	[8:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg;
	wire	[127:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start;
	wire	[4:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid;
	wire	[1:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd;
	wire	[43:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle;
	wire	[2:0]	w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb;
	wire		w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk;
	wire	[63:0]	w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
	wire	[3:0]	w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
	wire		w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
	wire		w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
	wire		w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
	wire		w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
	wire		w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
	
	// wires for module twentynm_hssi_tx_pcs_pma_interface
	wire	[7:0]	w_hssi_tx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_tx_pcs_pma_interface_blockselect;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out;
	wire		w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out;
	wire	[4:0]	w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk;
	wire		w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_pma_tx_pma_data;
	wire		w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback;
	wire	[63:0]	w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_1;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_2;
	wire	[19:0]	w_hssi_tx_pcs_pma_interface_uhsif_test_out_3;
	
	// wires for module twentynm_hssi_rx_pcs_pma_interface
	wire	[7:0]	w_hssi_rx_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_rx_pcs_pma_interface_blockselect;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni;
	wire	[31:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user;
	wire	[63:0]	w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock;
	wire		w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok;
	wire		w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk;
	wire	[5:0]	w_hssi_rx_pcs_pma_interface_pma_eye_monitor;
	wire		w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
	wire		w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out;
	wire	[19:0]	w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test;
	
	// wires for module twentynm_hssi_10g_tx_pcs
	wire	[7:0]	w_hssi_10g_tx_pcs_avmmreaddata;
	wire		w_hssi_10g_tx_pcs_blockselect;
	wire		w_hssi_10g_tx_pcs_distdwn_out_dv;
	wire		w_hssi_10g_tx_pcs_distdwn_out_rden;
	wire		w_hssi_10g_tx_pcs_distdwn_out_wren;
	wire		w_hssi_10g_tx_pcs_distup_out_dv;
	wire		w_hssi_10g_tx_pcs_distup_out_rden;
	wire		w_hssi_10g_tx_pcs_distup_out_wren;
	wire		w_hssi_10g_tx_pcs_tx_burst_en_exe;
	wire		w_hssi_10g_tx_pcs_tx_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_10g_tx_pcs_tx_clk_out_pma_if;
	wire	[8:0]	w_hssi_10g_tx_pcs_tx_control_out_krfec;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_data_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_data_valid_out_krfec;
	wire		w_hssi_10g_tx_pcs_tx_dft_clk_out;
	wire		w_hssi_10g_tx_pcs_tx_empty;
	wire		w_hssi_10g_tx_pcs_tx_fec_clk;
	wire	[3:0]	w_hssi_10g_tx_pcs_tx_fifo_num;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_rd_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_clk;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data;
	wire	[72:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_en;
	wire	[15:0]	w_hssi_10g_tx_pcs_tx_fifo_wr_ptr;
	wire		w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_frame;
	wire		w_hssi_10g_tx_pcs_tx_full;
	wire		w_hssi_10g_tx_pcs_tx_master_clk;
	wire		w_hssi_10g_tx_pcs_tx_master_clk_rst_n;
	wire		w_hssi_10g_tx_pcs_tx_pempty;
	wire		w_hssi_10g_tx_pcs_tx_pfull;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_data;
	wire	[63:0]	w_hssi_10g_tx_pcs_tx_pma_gating_val;
	wire	[19:0]	w_hssi_10g_tx_pcs_tx_test_data;
	wire		w_hssi_10g_tx_pcs_tx_wordslip_exe;
	
	// wires for module twentynm_hssi_8g_tx_pcs
	wire	[7:0]	w_hssi_8g_tx_pcs_avmmreaddata;
	wire		w_hssi_8g_tx_pcs_blockselect;
	wire		w_hssi_8g_tx_pcs_clk_out;
	wire		w_hssi_8g_tx_pcs_clk_out_gen3;
	wire	[19:0]	w_hssi_8g_tx_pcs_dataout;
	wire		w_hssi_8g_tx_pcs_dyn_clk_switch_n;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_fifo_select_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn;
	wire		w_hssi_8g_tx_pcs_g3_tx_pma_rstn;
	wire	[2:0]	w_hssi_8g_tx_pcs_non_gray_eidleinfersel;
	wire		w_hssi_8g_tx_pcs_ph_fifo_overflow;
	wire		w_hssi_8g_tx_pcs_ph_fifo_underflow;
	wire		w_hssi_8g_tx_pcs_phfifo_txdeemph;
	wire	[2:0]	w_hssi_8g_tx_pcs_phfifo_txmargin;
	wire		w_hssi_8g_tx_pcs_phfifo_txswing;
	wire		w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out;
	wire	[1:0]	w_hssi_8g_tx_pcs_pipe_power_down_out;
	wire		w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3;
	wire		w_hssi_8g_tx_pcs_pmaif_asn_rstn;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_rd_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_refclk_b;
	wire		w_hssi_8g_tx_pcs_refclk_b_reset;
	wire		w_hssi_8g_tx_pcs_rxpolarity_int;
	wire		w_hssi_8g_tx_pcs_soft_reset_wclk1_n;
	wire		w_hssi_8g_tx_pcs_sw_fifo_wr_clk;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_blk_start_out;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pld_if;
	wire		w_hssi_8g_tx_pcs_tx_clk_out_pmaif;
	wire		w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_ctrlplane_testbus;
	wire	[31:0]	w_hssi_8g_tx_pcs_tx_data_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_data_valid_out;
	wire	[3:0]	w_hssi_8g_tx_pcs_tx_datak_out;
	wire		w_hssi_8g_tx_pcs_tx_detect_rxloopback_int;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up;
	wire		w_hssi_8g_tx_pcs_tx_pipe_clk;
	wire		w_hssi_8g_tx_pcs_tx_pipe_electidle;
	wire		w_hssi_8g_tx_pcs_tx_pipe_soft_reset;
	wire	[1:0]	w_hssi_8g_tx_pcs_tx_sync_hdr_out;
	wire	[19:0]	w_hssi_8g_tx_pcs_tx_testbus;
	wire		w_hssi_8g_tx_pcs_txcompliance_out;
	wire		w_hssi_8g_tx_pcs_txelecidle_out;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk;
	wire		w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk;
	wire	[63:0]	w_hssi_8g_tx_pcs_wr_data_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_en_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_tx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo;
	wire		w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo;
	
	// wires for module twentynm_hssi_pipe_gen3
	wire	[7:0]	w_hssi_pipe_gen3_avmmreaddata;
	wire		w_hssi_pipe_gen3_blockselect;
	wire		w_hssi_pipe_gen3_gen3_clk_sel;
	wire		w_hssi_pipe_gen3_pcs_rst;
	wire		w_hssi_pipe_gen3_phystatus;
	wire	[17:0]	w_hssi_pipe_gen3_pma_current_coeff;
	wire	[2:0]	w_hssi_pipe_gen3_pma_current_rxpreset;
	wire		w_hssi_pipe_gen3_pma_tx_elec_idle;
	wire		w_hssi_pipe_gen3_pma_txdetectrx;
	wire		w_hssi_pipe_gen3_rev_lpbk_8gpcs_out;
	wire		w_hssi_pipe_gen3_rev_lpbk_int;
	wire	[3:0]	w_hssi_pipe_gen3_rx_blk_start;
	wire	[1:0]	w_hssi_pipe_gen3_rx_sync_hdr;
	wire	[63:0]	w_hssi_pipe_gen3_rxd_8gpcs_out;
	wire	[3:0]	w_hssi_pipe_gen3_rxdataskip;
	wire		w_hssi_pipe_gen3_rxelecidle;
	wire		w_hssi_pipe_gen3_rxpolarity_8gpcs_out;
	wire		w_hssi_pipe_gen3_rxpolarity_int;
	wire	[2:0]	w_hssi_pipe_gen3_rxstatus;
	wire		w_hssi_pipe_gen3_rxvalid;
	wire		w_hssi_pipe_gen3_shutdown_clk;
	wire	[19:0]	w_hssi_pipe_gen3_test_out;
	wire		w_hssi_pipe_gen3_tx_blk_start_int;
	wire	[1:0]	w_hssi_pipe_gen3_tx_sync_hdr_int;
	wire	[31:0]	w_hssi_pipe_gen3_txdata_int;
	wire	[3:0]	w_hssi_pipe_gen3_txdatak_int;
	wire		w_hssi_pipe_gen3_txdataskip_int;
	
	// wires for module twentynm_hssi_pipe_gen1_2
	wire	[7:0]	w_hssi_pipe_gen1_2_avmmreaddata;
	wire		w_hssi_pipe_gen1_2_blockselect;
	wire	[17:0]	w_hssi_pipe_gen1_2_current_coeff;
	wire		w_hssi_pipe_gen1_2_phystatus;
	wire		w_hssi_pipe_gen1_2_polarity_inversion_rx;
	wire		w_hssi_pipe_gen1_2_rev_loopbk;
	wire		w_hssi_pipe_gen1_2_rxelecidle;
	wire		w_hssi_pipe_gen1_2_rxelectricalidle_out;
	wire	[2:0]	w_hssi_pipe_gen1_2_rxstatus;
	wire		w_hssi_pipe_gen1_2_rxvalid;
	wire		w_hssi_pipe_gen1_2_tx_elec_idle_out;
	wire		w_hssi_pipe_gen1_2_txdetectrx;
	
	// wires for module twentynm_hssi_gen3_tx_pcs
	wire	[7:0]	w_hssi_gen3_tx_pcs_avmmreaddata;
	wire		w_hssi_gen3_tx_pcs_blockselect;
	wire	[31:0]	w_hssi_gen3_tx_pcs_data_out;
	wire	[35:0]	w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out;
	wire	[31:0]	w_hssi_gen3_tx_pcs_par_lpbk_out;
	wire	[19:0]	w_hssi_gen3_tx_pcs_tx_test_out;
	
	// wires for module twentynm_hssi_8g_rx_pcs
	wire	[3:0]	w_hssi_8g_rx_pcs_a1a2k1k2flag;
	wire	[7:0]	w_hssi_8g_rx_pcs_avmmreaddata;
	wire		w_hssi_8g_rx_pcs_blockselect;
	wire	[19:0]	w_hssi_8g_rx_pcs_chnl_test_bus_out;
	wire		w_hssi_8g_rx_pcs_clock_to_pld;
	wire	[63:0]	w_hssi_8g_rx_pcs_dataout;
	wire		w_hssi_8g_rx_pcs_dis_pc_byte;
	wire		w_hssi_8g_rx_pcs_eidle_detected;
	wire	[2:0]	w_hssi_8g_rx_pcs_eios_det_cdr_ctrl;
	wire		w_hssi_8g_rx_pcs_g3_rx_pma_rstn;
	wire		w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn;
	wire		w_hssi_8g_rx_pcs_gen2ngen1;
	wire	[19:0]	w_hssi_8g_rx_pcs_parallel_rev_loopback;
	wire		w_hssi_8g_rx_pcs_pc_fifo_empty;
	wire		w_hssi_8g_rx_pcs_pcfifofull;
	wire		w_hssi_8g_rx_pcs_phystatus;
	wire	[63:0]	w_hssi_8g_rx_pcs_pipe_data;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_rd_enable_out_chnl_up;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo;
	wire	[7:0]	w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rm_fifo_empty;
	wire		w_hssi_8g_rx_pcs_rm_fifo_full;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_blk_start;
	wire		w_hssi_8g_rx_pcs_rx_clk_out_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if;
	wire		w_hssi_8g_rx_pcs_rx_clkslip;
	wire	[3:0]	w_hssi_8g_rx_pcs_rx_data_valid;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up;
	wire		w_hssi_8g_rx_pcs_rx_pipe_clk;
	wire		w_hssi_8g_rx_pcs_rx_pipe_soft_reset;
	wire		w_hssi_8g_rx_pcs_rx_pma_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3;
	wire		w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_sync_hdr;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_down;
	wire	[1:0]	w_hssi_8g_rx_pcs_rx_we_out_chnl_up;
	wire	[2:0]	w_hssi_8g_rx_pcs_rxstatus;
	wire		w_hssi_8g_rx_pcs_rxvalid;
	wire		w_hssi_8g_rx_pcs_signal_detect_out;
	wire	[4:0]	w_hssi_8g_rx_pcs_word_align_boundary;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk;
	wire		w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk;
	wire	[79:0]	w_hssi_8g_rx_pcs_wr_data_rx_phfifo;
	wire	[31:0]	w_hssi_8g_rx_pcs_wr_data_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_en_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_down;
	wire		w_hssi_8g_rx_pcs_wr_enable_out_chnl_up;
	wire	[7:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo;
	wire	[19:0]	w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo;
	wire		w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo;
	
	// wires for module twentynm_hssi_fifo_rx_pcs
	wire	[7:0]	w_hssi_fifo_rx_pcs_avmmreaddata;
	wire		w_hssi_fifo_rx_pcs_blockselect;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out2_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp;
	wire	[73:0]	w_hssi_fifo_rx_pcs_data_out_10g;
	wire	[31:0]	w_hssi_fifo_rx_pcs_data_out_8g_clock_comp;
	wire	[79:0]	w_hssi_fifo_rx_pcs_data_out_8g_phase_comp;
	wire	[39:0]	w_hssi_fifo_rx_pcs_data_out_gen3;
	
	// wires for module twentynm_hssi_common_pcs_pma_interface
	wire	[7:0]	w_hssi_common_pcs_pma_interface_avmmreaddata;
	wire		w_hssi_common_pcs_pma_interface_blockselect;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid;
	wire	[8:0]	w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref;
	wire		w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in;
	wire	[19:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out;
	wire	[7:0]	w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus;
	wire		w_hssi_common_pcs_pma_interface_pma_adapt_start;
	wire		w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
	wire		w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
	wire	[17:0]	w_hssi_common_pcs_pma_interface_pma_current_coeff;
	wire	[2:0]	w_hssi_common_pcs_pma_interface_pma_current_rxpreset;
	wire		w_hssi_common_pcs_pma_interface_pma_early_eios;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_interface_select;
	wire		w_hssi_common_pcs_pma_interface_pma_ltd_b;
	wire		w_hssi_common_pcs_pma_interface_pma_ltr;
	wire		w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
	wire		w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
	wire	[1:0]	w_hssi_common_pcs_pma_interface_pma_pcie_switch;
	wire		w_hssi_common_pcs_pma_interface_pma_ppm_lock;
	wire	[4:0]	w_hssi_common_pcs_pma_interface_pma_reserved_out;
	wire		w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
	wire		w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
	wire		w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
	wire		w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down;
	wire	[11:0]	w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up;
	
	
	generate
		
		//module instantiations
		
		// instantiating twentynm_hssi_10g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_rx_pcs
			twentynm_hssi_10g_rx_pcs #(
				.advanced_user_mode(hssi_10g_rx_pcs_advanced_user_mode),
				.align_del(hssi_10g_rx_pcs_align_del),
				.ber_bit_err_total_cnt(hssi_10g_rx_pcs_ber_bit_err_total_cnt),
				.ber_clken(hssi_10g_rx_pcs_ber_clken),
				.ber_xus_timer_window(hssi_10g_rx_pcs_ber_xus_timer_window),
				.bitslip_mode(hssi_10g_rx_pcs_bitslip_mode),
				.blksync_bitslip_type(hssi_10g_rx_pcs_blksync_bitslip_type),
				.blksync_bitslip_wait_cnt(hssi_10g_rx_pcs_blksync_bitslip_wait_cnt),
				.blksync_bitslip_wait_type(hssi_10g_rx_pcs_blksync_bitslip_wait_type),
				.blksync_bypass(hssi_10g_rx_pcs_blksync_bypass),
				.blksync_clken(hssi_10g_rx_pcs_blksync_clken),
				.blksync_enum_invalid_sh_cnt(hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt),
				.blksync_knum_sh_cnt_postlock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock),
				.blksync_knum_sh_cnt_prelock(hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock),
				.blksync_pipeln(hssi_10g_rx_pcs_blksync_pipeln),
				.clr_errblk_cnt_en(hssi_10g_rx_pcs_clr_errblk_cnt_en),
				.control_del(hssi_10g_rx_pcs_control_del),
				.crcchk_bypass(hssi_10g_rx_pcs_crcchk_bypass),
				.crcchk_clken(hssi_10g_rx_pcs_crcchk_clken),
				.crcchk_inv(hssi_10g_rx_pcs_crcchk_inv),
				.crcchk_pipeln(hssi_10g_rx_pcs_crcchk_pipeln),
				.crcflag_pipeln(hssi_10g_rx_pcs_crcflag_pipeln),
				.ctrl_bit_reverse(hssi_10g_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_10g_rx_pcs_data_bit_reverse),
				.dec64b66b_clken(hssi_10g_rx_pcs_dec64b66b_clken),
				.dec_64b66b_rxsm_bypass(hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass),
				.descrm_bypass(hssi_10g_rx_pcs_descrm_bypass),
				.descrm_clken(hssi_10g_rx_pcs_descrm_clken),
				.descrm_mode(hssi_10g_rx_pcs_descrm_mode),
				.descrm_pipeln(hssi_10g_rx_pcs_descrm_pipeln),
				.dft_clk_out_sel(hssi_10g_rx_pcs_dft_clk_out_sel),
				.dis_signal_ok(hssi_10g_rx_pcs_dis_signal_ok),
				.dispchk_bypass(hssi_10g_rx_pcs_dispchk_bypass),
				.empty_flag_type(hssi_10g_rx_pcs_empty_flag_type),
				.fast_path(hssi_10g_rx_pcs_fast_path),
				.fec_clken(hssi_10g_rx_pcs_fec_clken),
				.fec_enable(hssi_10g_rx_pcs_fec_enable),
				.fifo_double_read(hssi_10g_rx_pcs_fifo_double_read),
				.fifo_stop_rd(hssi_10g_rx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_rx_pcs_fifo_stop_wr),
				.force_align(hssi_10g_rx_pcs_force_align),
				.frmsync_bypass(hssi_10g_rx_pcs_frmsync_bypass),
				.frmsync_clken(hssi_10g_rx_pcs_frmsync_clken),
				.frmsync_enum_scrm(hssi_10g_rx_pcs_frmsync_enum_scrm),
				.frmsync_enum_sync(hssi_10g_rx_pcs_frmsync_enum_sync),
				.frmsync_flag_type(hssi_10g_rx_pcs_frmsync_flag_type),
				.frmsync_knum_sync(hssi_10g_rx_pcs_frmsync_knum_sync),
				.frmsync_mfrm_length(hssi_10g_rx_pcs_frmsync_mfrm_length),
				.frmsync_pipeln(hssi_10g_rx_pcs_frmsync_pipeln),
				.full_flag_type(hssi_10g_rx_pcs_full_flag_type),
				.gb_rx_idwidth(hssi_10g_rx_pcs_gb_rx_idwidth),
				.gb_rx_odwidth(hssi_10g_rx_pcs_gb_rx_odwidth),
				.gbexp_clken(hssi_10g_rx_pcs_gbexp_clken),
				.low_latency_en(hssi_10g_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_10g_rx_pcs_lpbk_mode),
				.master_clk_sel(hssi_10g_rx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_rx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_rx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_rx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_rx_pcs_pld_if_type),
				.prot_mode(hssi_10g_rx_pcs_prot_mode),
				.rand_clken(hssi_10g_rx_pcs_rand_clken),
				.rd_clk_sel(hssi_10g_rx_pcs_rd_clk_sel),
				.rdfifo_clken(hssi_10g_rx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_rx_pcs_reconfig_settings),
				.rx_fifo_write_ctrl(hssi_10g_rx_pcs_rx_fifo_write_ctrl),
				.rx_scrm_width(hssi_10g_rx_pcs_rx_scrm_width),
				.rx_sh_location(hssi_10g_rx_pcs_rx_sh_location),
				.rx_signal_ok_sel(hssi_10g_rx_pcs_rx_signal_ok_sel),
				.rx_sm_bypass(hssi_10g_rx_pcs_rx_sm_bypass),
				.rx_sm_hiber(hssi_10g_rx_pcs_rx_sm_hiber),
				.rx_sm_pipeln(hssi_10g_rx_pcs_rx_sm_pipeln),
				.rx_testbus_sel(hssi_10g_rx_pcs_rx_testbus_sel),
				.rx_true_b2b(hssi_10g_rx_pcs_rx_true_b2b),
				.rxfifo_empty(hssi_10g_rx_pcs_rxfifo_empty),
				.rxfifo_full(hssi_10g_rx_pcs_rxfifo_full),
				.rxfifo_mode(hssi_10g_rx_pcs_rxfifo_mode),
				.rxfifo_pempty(hssi_10g_rx_pcs_rxfifo_pempty),
				.rxfifo_pfull(hssi_10g_rx_pcs_rxfifo_pfull),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.stretch_num_stages(hssi_10g_rx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_rx_pcs_sup_mode),
				.test_mode(hssi_10g_rx_pcs_test_mode),
				.wrfifo_clken(hssi_10g_rx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_rx_pcs_blockselect),
				.rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.rx_control(w_hssi_10g_rx_pcs_rx_control),
				.rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.rx_data(w_hssi_10g_rx_pcs_rx_data),
				.rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.rx_diag_status(w_hssi_10g_rx_pcs_rx_diag_status),
				.rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.rx_fec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.rx_fifo_num(w_hssi_10g_rx_pcs_rx_fifo_num),
				.rx_fifo_rd_ptr(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr),
				.rx_fifo_rd_ptr2(w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2),
				.rx_fifo_wr_clk(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.rx_fifo_wr_data(w_hssi_10g_rx_pcs_rx_fifo_wr_data),
				.rx_fifo_wr_en(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.rx_fifo_wr_ptr(w_hssi_10g_rx_pcs_rx_fifo_wr_ptr),
				.rx_fifo_wr_rst_n(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.rx_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_rx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_rx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_rx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.rx_control_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0]}),
				.rx_control_in_krfec({w_hssi_krfec_rx_pcs_rx_control_out[9], w_hssi_krfec_rx_pcs_rx_control_out[8], w_hssi_krfec_rx_pcs_rx_control_out[7], w_hssi_krfec_rx_pcs_rx_control_out[6], w_hssi_krfec_rx_pcs_rx_control_out[5], w_hssi_krfec_rx_pcs_rx_control_out[4], w_hssi_krfec_rx_pcs_rx_control_out[3], w_hssi_krfec_rx_pcs_rx_control_out[2], w_hssi_krfec_rx_pcs_rx_control_out[1], w_hssi_krfec_rx_pcs_rx_control_out[0]}),
				.rx_data_fb({w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1], w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0]}),
				.rx_data_in_krfec({w_hssi_krfec_rx_pcs_rx_data_out[63], w_hssi_krfec_rx_pcs_rx_data_out[62], w_hssi_krfec_rx_pcs_rx_data_out[61], w_hssi_krfec_rx_pcs_rx_data_out[60], w_hssi_krfec_rx_pcs_rx_data_out[59], w_hssi_krfec_rx_pcs_rx_data_out[58], w_hssi_krfec_rx_pcs_rx_data_out[57], w_hssi_krfec_rx_pcs_rx_data_out[56], w_hssi_krfec_rx_pcs_rx_data_out[55], w_hssi_krfec_rx_pcs_rx_data_out[54], w_hssi_krfec_rx_pcs_rx_data_out[53], w_hssi_krfec_rx_pcs_rx_data_out[52], w_hssi_krfec_rx_pcs_rx_data_out[51], w_hssi_krfec_rx_pcs_rx_data_out[50], w_hssi_krfec_rx_pcs_rx_data_out[49], w_hssi_krfec_rx_pcs_rx_data_out[48], w_hssi_krfec_rx_pcs_rx_data_out[47], w_hssi_krfec_rx_pcs_rx_data_out[46], w_hssi_krfec_rx_pcs_rx_data_out[45], w_hssi_krfec_rx_pcs_rx_data_out[44], w_hssi_krfec_rx_pcs_rx_data_out[43], w_hssi_krfec_rx_pcs_rx_data_out[42], w_hssi_krfec_rx_pcs_rx_data_out[41], w_hssi_krfec_rx_pcs_rx_data_out[40], w_hssi_krfec_rx_pcs_rx_data_out[39], w_hssi_krfec_rx_pcs_rx_data_out[38], w_hssi_krfec_rx_pcs_rx_data_out[37], w_hssi_krfec_rx_pcs_rx_data_out[36], w_hssi_krfec_rx_pcs_rx_data_out[35], w_hssi_krfec_rx_pcs_rx_data_out[34], w_hssi_krfec_rx_pcs_rx_data_out[33], w_hssi_krfec_rx_pcs_rx_data_out[32], w_hssi_krfec_rx_pcs_rx_data_out[31], w_hssi_krfec_rx_pcs_rx_data_out[30], w_hssi_krfec_rx_pcs_rx_data_out[29], w_hssi_krfec_rx_pcs_rx_data_out[28], w_hssi_krfec_rx_pcs_rx_data_out[27], w_hssi_krfec_rx_pcs_rx_data_out[26], w_hssi_krfec_rx_pcs_rx_data_out[25], w_hssi_krfec_rx_pcs_rx_data_out[24], w_hssi_krfec_rx_pcs_rx_data_out[23], w_hssi_krfec_rx_pcs_rx_data_out[22], w_hssi_krfec_rx_pcs_rx_data_out[21], w_hssi_krfec_rx_pcs_rx_data_out[20], w_hssi_krfec_rx_pcs_rx_data_out[19], w_hssi_krfec_rx_pcs_rx_data_out[18], w_hssi_krfec_rx_pcs_rx_data_out[17], w_hssi_krfec_rx_pcs_rx_data_out[16], w_hssi_krfec_rx_pcs_rx_data_out[15], w_hssi_krfec_rx_pcs_rx_data_out[14], w_hssi_krfec_rx_pcs_rx_data_out[13], w_hssi_krfec_rx_pcs_rx_data_out[12], w_hssi_krfec_rx_pcs_rx_data_out[11], w_hssi_krfec_rx_pcs_rx_data_out[10], w_hssi_krfec_rx_pcs_rx_data_out[9], w_hssi_krfec_rx_pcs_rx_data_out[8], w_hssi_krfec_rx_pcs_rx_data_out[7], w_hssi_krfec_rx_pcs_rx_data_out[6], w_hssi_krfec_rx_pcs_rx_data_out[5], w_hssi_krfec_rx_pcs_rx_data_out[4], w_hssi_krfec_rx_pcs_rx_data_out[3], w_hssi_krfec_rx_pcs_rx_data_out[2], w_hssi_krfec_rx_pcs_rx_data_out[1], w_hssi_krfec_rx_pcs_rx_data_out[0]}),
				.rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.rx_data_valid_in_krfec(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_10g[73], w_hssi_fifo_rx_pcs_data_out_10g[72], w_hssi_fifo_rx_pcs_data_out_10g[71], w_hssi_fifo_rx_pcs_data_out_10g[70], w_hssi_fifo_rx_pcs_data_out_10g[69], w_hssi_fifo_rx_pcs_data_out_10g[68], w_hssi_fifo_rx_pcs_data_out_10g[67], w_hssi_fifo_rx_pcs_data_out_10g[66], w_hssi_fifo_rx_pcs_data_out_10g[65], w_hssi_fifo_rx_pcs_data_out_10g[64], w_hssi_fifo_rx_pcs_data_out_10g[63], w_hssi_fifo_rx_pcs_data_out_10g[62], w_hssi_fifo_rx_pcs_data_out_10g[61], w_hssi_fifo_rx_pcs_data_out_10g[60], w_hssi_fifo_rx_pcs_data_out_10g[59], w_hssi_fifo_rx_pcs_data_out_10g[58], w_hssi_fifo_rx_pcs_data_out_10g[57], w_hssi_fifo_rx_pcs_data_out_10g[56], w_hssi_fifo_rx_pcs_data_out_10g[55], w_hssi_fifo_rx_pcs_data_out_10g[54], w_hssi_fifo_rx_pcs_data_out_10g[53], w_hssi_fifo_rx_pcs_data_out_10g[52], w_hssi_fifo_rx_pcs_data_out_10g[51], w_hssi_fifo_rx_pcs_data_out_10g[50], w_hssi_fifo_rx_pcs_data_out_10g[49], w_hssi_fifo_rx_pcs_data_out_10g[48], w_hssi_fifo_rx_pcs_data_out_10g[47], w_hssi_fifo_rx_pcs_data_out_10g[46], w_hssi_fifo_rx_pcs_data_out_10g[45], w_hssi_fifo_rx_pcs_data_out_10g[44], w_hssi_fifo_rx_pcs_data_out_10g[43], w_hssi_fifo_rx_pcs_data_out_10g[42], w_hssi_fifo_rx_pcs_data_out_10g[41], w_hssi_fifo_rx_pcs_data_out_10g[40], w_hssi_fifo_rx_pcs_data_out_10g[39], w_hssi_fifo_rx_pcs_data_out_10g[38], w_hssi_fifo_rx_pcs_data_out_10g[37], w_hssi_fifo_rx_pcs_data_out_10g[36], w_hssi_fifo_rx_pcs_data_out_10g[35], w_hssi_fifo_rx_pcs_data_out_10g[34], w_hssi_fifo_rx_pcs_data_out_10g[33], w_hssi_fifo_rx_pcs_data_out_10g[32], w_hssi_fifo_rx_pcs_data_out_10g[31], w_hssi_fifo_rx_pcs_data_out_10g[30], w_hssi_fifo_rx_pcs_data_out_10g[29], w_hssi_fifo_rx_pcs_data_out_10g[28], w_hssi_fifo_rx_pcs_data_out_10g[27], w_hssi_fifo_rx_pcs_data_out_10g[26], w_hssi_fifo_rx_pcs_data_out_10g[25], w_hssi_fifo_rx_pcs_data_out_10g[24], w_hssi_fifo_rx_pcs_data_out_10g[23], w_hssi_fifo_rx_pcs_data_out_10g[22], w_hssi_fifo_rx_pcs_data_out_10g[21], w_hssi_fifo_rx_pcs_data_out_10g[20], w_hssi_fifo_rx_pcs_data_out_10g[19], w_hssi_fifo_rx_pcs_data_out_10g[18], w_hssi_fifo_rx_pcs_data_out_10g[17], w_hssi_fifo_rx_pcs_data_out_10g[16], w_hssi_fifo_rx_pcs_data_out_10g[15], w_hssi_fifo_rx_pcs_data_out_10g[14], w_hssi_fifo_rx_pcs_data_out_10g[13], w_hssi_fifo_rx_pcs_data_out_10g[12], w_hssi_fifo_rx_pcs_data_out_10g[11], w_hssi_fifo_rx_pcs_data_out_10g[10], w_hssi_fifo_rx_pcs_data_out_10g[9], w_hssi_fifo_rx_pcs_data_out_10g[8], w_hssi_fifo_rx_pcs_data_out_10g[7], w_hssi_fifo_rx_pcs_data_out_10g[6], w_hssi_fifo_rx_pcs_data_out_10g[5], w_hssi_fifo_rx_pcs_data_out_10g[4], w_hssi_fifo_rx_pcs_data_out_10g[3], w_hssi_fifo_rx_pcs_data_out_10g[2], w_hssi_fifo_rx_pcs_data_out_10g[1], w_hssi_fifo_rx_pcs_data_out_10g[0]}),
				.rx_fifo_rd_data_dw({w_hssi_fifo_rx_pcs_data_out2_10g[73], w_hssi_fifo_rx_pcs_data_out2_10g[72], w_hssi_fifo_rx_pcs_data_out2_10g[71], w_hssi_fifo_rx_pcs_data_out2_10g[70], w_hssi_fifo_rx_pcs_data_out2_10g[69], w_hssi_fifo_rx_pcs_data_out2_10g[68], w_hssi_fifo_rx_pcs_data_out2_10g[67], w_hssi_fifo_rx_pcs_data_out2_10g[66], w_hssi_fifo_rx_pcs_data_out2_10g[65], w_hssi_fifo_rx_pcs_data_out2_10g[64], w_hssi_fifo_rx_pcs_data_out2_10g[63], w_hssi_fifo_rx_pcs_data_out2_10g[62], w_hssi_fifo_rx_pcs_data_out2_10g[61], w_hssi_fifo_rx_pcs_data_out2_10g[60], w_hssi_fifo_rx_pcs_data_out2_10g[59], w_hssi_fifo_rx_pcs_data_out2_10g[58], w_hssi_fifo_rx_pcs_data_out2_10g[57], w_hssi_fifo_rx_pcs_data_out2_10g[56], w_hssi_fifo_rx_pcs_data_out2_10g[55], w_hssi_fifo_rx_pcs_data_out2_10g[54], w_hssi_fifo_rx_pcs_data_out2_10g[53], w_hssi_fifo_rx_pcs_data_out2_10g[52], w_hssi_fifo_rx_pcs_data_out2_10g[51], w_hssi_fifo_rx_pcs_data_out2_10g[50], w_hssi_fifo_rx_pcs_data_out2_10g[49], w_hssi_fifo_rx_pcs_data_out2_10g[48], w_hssi_fifo_rx_pcs_data_out2_10g[47], w_hssi_fifo_rx_pcs_data_out2_10g[46], w_hssi_fifo_rx_pcs_data_out2_10g[45], w_hssi_fifo_rx_pcs_data_out2_10g[44], w_hssi_fifo_rx_pcs_data_out2_10g[43], w_hssi_fifo_rx_pcs_data_out2_10g[42], w_hssi_fifo_rx_pcs_data_out2_10g[41], w_hssi_fifo_rx_pcs_data_out2_10g[40], w_hssi_fifo_rx_pcs_data_out2_10g[39], w_hssi_fifo_rx_pcs_data_out2_10g[38], w_hssi_fifo_rx_pcs_data_out2_10g[37], w_hssi_fifo_rx_pcs_data_out2_10g[36], w_hssi_fifo_rx_pcs_data_out2_10g[35], w_hssi_fifo_rx_pcs_data_out2_10g[34], w_hssi_fifo_rx_pcs_data_out2_10g[33], w_hssi_fifo_rx_pcs_data_out2_10g[32], w_hssi_fifo_rx_pcs_data_out2_10g[31], w_hssi_fifo_rx_pcs_data_out2_10g[30], w_hssi_fifo_rx_pcs_data_out2_10g[29], w_hssi_fifo_rx_pcs_data_out2_10g[28], w_hssi_fifo_rx_pcs_data_out2_10g[27], w_hssi_fifo_rx_pcs_data_out2_10g[26], w_hssi_fifo_rx_pcs_data_out2_10g[25], w_hssi_fifo_rx_pcs_data_out2_10g[24], w_hssi_fifo_rx_pcs_data_out2_10g[23], w_hssi_fifo_rx_pcs_data_out2_10g[22], w_hssi_fifo_rx_pcs_data_out2_10g[21], w_hssi_fifo_rx_pcs_data_out2_10g[20], w_hssi_fifo_rx_pcs_data_out2_10g[19], w_hssi_fifo_rx_pcs_data_out2_10g[18], w_hssi_fifo_rx_pcs_data_out2_10g[17], w_hssi_fifo_rx_pcs_data_out2_10g[16], w_hssi_fifo_rx_pcs_data_out2_10g[15], w_hssi_fifo_rx_pcs_data_out2_10g[14], w_hssi_fifo_rx_pcs_data_out2_10g[13], w_hssi_fifo_rx_pcs_data_out2_10g[12], w_hssi_fifo_rx_pcs_data_out2_10g[11], w_hssi_fifo_rx_pcs_data_out2_10g[10], w_hssi_fifo_rx_pcs_data_out2_10g[9], w_hssi_fifo_rx_pcs_data_out2_10g[8], w_hssi_fifo_rx_pcs_data_out2_10g[7], w_hssi_fifo_rx_pcs_data_out2_10g[6], w_hssi_fifo_rx_pcs_data_out2_10g[5], w_hssi_fifo_rx_pcs_data_out2_10g[4], w_hssi_fifo_rx_pcs_data_out2_10g[3], w_hssi_fifo_rx_pcs_data_out2_10g[2], w_hssi_fifo_rx_pcs_data_out2_10g[1], w_hssi_fifo_rx_pcs_data_out2_10g[0]}),
				.rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.rx_pma_data({w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0]}),
				.rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.signal_ok_krfec(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_10g_reg(),
				.pld_10g_krfec_rx_blk_lock_10g_txclk_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_reg(),
				.pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_reg(),
				.pld_10g_krfec_rx_diag_data_status_10g_txclk_reg(),
				.pld_10g_krfec_rx_frame_10g_reg(),
				.pld_10g_krfec_rx_frame_10g_txclk_reg(),
				.pld_10g_krfec_rx_pld_rst_n_fifo(),
				.pld_10g_krfec_rx_pld_rst_n_reg(),
				.pld_10g_krfec_rx_pld_rst_n_txclk_reg(),
				.pld_10g_rx_align_clr_fifo(),
				.pld_10g_rx_align_clr_reg(),
				.pld_10g_rx_align_clr_txclk_reg(),
				.pld_10g_rx_align_val_fifo(),
				.pld_10g_rx_align_val_reg(),
				.pld_10g_rx_align_val_txclk_reg(),
				.pld_10g_rx_clr_ber_count_reg(),
				.pld_10g_rx_clr_ber_count_txclk_reg(),
				.pld_10g_rx_crc32_err_reg(),
				.pld_10g_rx_crc32_err_txclk_reg(),
				.pld_10g_rx_data_valid_10g_reg(),
				.pld_10g_rx_data_valid_fifo(),
				.pld_10g_rx_data_valid_pcsdirect_reg(),
				.pld_10g_rx_data_valid_txclk_reg(),
				.pld_10g_rx_empty_fifo(),
				.pld_10g_rx_fifo_del_reg(),
				.pld_10g_rx_fifo_del_txclk_reg(),
				.pld_10g_rx_fifo_insert_fifo(),
				.pld_10g_rx_fifo_num_reg(),
				.pld_10g_rx_fifo_num_txclk_reg(),
				.pld_10g_rx_frame_lock_reg(),
				.pld_10g_rx_frame_lock_txclk_reg(),
				.pld_10g_rx_hi_ber_reg(),
				.pld_10g_rx_hi_ber_txclk_reg(),
				.pld_10g_rx_oflw_err_reg(),
				.pld_10g_rx_oflw_err_txclk_reg(),
				.pld_10g_rx_pempty_fifo(),
				.pld_10g_rx_pfull_reg(),
				.pld_10g_rx_pfull_txclk_reg(),
				.pld_10g_rx_rd_en_fifo(),
				.pld_pcs_rx_clk_out_10g_txclk_wire(),
				.pld_pcs_rx_clk_out_10g_wire(),
				.pld_rx_control_10g_reg(),
				.pld_rx_control_10g_txclk_reg(),
				.pld_rx_data_10g_reg(),
				.pld_rx_data_10g_txclk_reg(),
				.pld_rx_prbs_err_10g_txclk_reg(),
				.pld_rx_prbs_err_clr_10g_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_10g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_align_val = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_blk_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_control[19:0] = 20'b0;
				assign w_hssi_10g_rx_pcs_rx_crc32_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_data[127:0] = 128'b0;
				assign w_hssi_10g_rx_pcs_rx_data_valid = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_dft_clk_out = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_diag_status[1:0] = 2'b0;
				assign w_hssi_10g_rx_pcs_rx_empty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fec_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_del = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_insert = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_data[73:0] = 74'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31:0] = 32'b0;
				assign w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_frame_lock = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_hi_ber = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_rx_pcs_rx_oflw_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pempty = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_pfull = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_random_err = 1'b0;
				assign w_hssi_10g_rx_pcs_rx_rx_frame = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_10g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_10g_tx_pcs
			twentynm_hssi_10g_tx_pcs #(
				.advanced_user_mode(hssi_10g_tx_pcs_advanced_user_mode),
				.bitslip_en(hssi_10g_tx_pcs_bitslip_en),
				.bonding_dft_en(hssi_10g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_10g_tx_pcs_bonding_dft_val),
				.comp_cnt(hssi_10g_tx_pcs_comp_cnt),
				.compin_sel(hssi_10g_tx_pcs_compin_sel),
				.crcgen_bypass(hssi_10g_tx_pcs_crcgen_bypass),
				.crcgen_clken(hssi_10g_tx_pcs_crcgen_clken),
				.crcgen_err(hssi_10g_tx_pcs_crcgen_err),
				.crcgen_inv(hssi_10g_tx_pcs_crcgen_inv),
				.ctrl_bit_reverse(hssi_10g_tx_pcs_ctrl_bit_reverse),
				.ctrl_plane_bonding(hssi_10g_tx_pcs_ctrl_plane_bonding),
				.data_bit_reverse(hssi_10g_tx_pcs_data_bit_reverse),
				.dft_clk_out_sel(hssi_10g_tx_pcs_dft_clk_out_sel),
				.dispgen_bypass(hssi_10g_tx_pcs_dispgen_bypass),
				.dispgen_clken(hssi_10g_tx_pcs_dispgen_clken),
				.dispgen_err(hssi_10g_tx_pcs_dispgen_err),
				.dispgen_pipeln(hssi_10g_tx_pcs_dispgen_pipeln),
				.distdwn_bypass_pipeln(hssi_10g_tx_pcs_distdwn_bypass_pipeln),
				.distdwn_master(hssi_10g_tx_pcs_distdwn_master),
				.distup_bypass_pipeln(hssi_10g_tx_pcs_distup_bypass_pipeln),
				.distup_master(hssi_10g_tx_pcs_distup_master),
				.dv_bond(hssi_10g_tx_pcs_dv_bond),
				.empty_flag_type(hssi_10g_tx_pcs_empty_flag_type),
				.enc64b66b_txsm_clken(hssi_10g_tx_pcs_enc64b66b_txsm_clken),
				.enc_64b66b_txsm_bypass(hssi_10g_tx_pcs_enc_64b66b_txsm_bypass),
				.fastpath(hssi_10g_tx_pcs_fastpath),
				.fec_clken(hssi_10g_tx_pcs_fec_clken),
				.fec_enable(hssi_10g_tx_pcs_fec_enable),
				.fifo_double_write(hssi_10g_tx_pcs_fifo_double_write),
				.fifo_reg_fast(hssi_10g_tx_pcs_fifo_reg_fast),
				.fifo_stop_rd(hssi_10g_tx_pcs_fifo_stop_rd),
				.fifo_stop_wr(hssi_10g_tx_pcs_fifo_stop_wr),
				.frmgen_burst(hssi_10g_tx_pcs_frmgen_burst),
				.frmgen_bypass(hssi_10g_tx_pcs_frmgen_bypass),
				.frmgen_clken(hssi_10g_tx_pcs_frmgen_clken),
				.frmgen_mfrm_length(hssi_10g_tx_pcs_frmgen_mfrm_length),
				.frmgen_pipeln(hssi_10g_tx_pcs_frmgen_pipeln),
				.frmgen_pyld_ins(hssi_10g_tx_pcs_frmgen_pyld_ins),
				.frmgen_wordslip(hssi_10g_tx_pcs_frmgen_wordslip),
				.full_flag_type(hssi_10g_tx_pcs_full_flag_type),
				.gb_pipeln_bypass(hssi_10g_tx_pcs_gb_pipeln_bypass),
				.gb_tx_idwidth(hssi_10g_tx_pcs_gb_tx_idwidth),
				.gb_tx_odwidth(hssi_10g_tx_pcs_gb_tx_odwidth),
				.gbred_clken(hssi_10g_tx_pcs_gbred_clken),
				.indv(hssi_10g_tx_pcs_indv),
				.low_latency_en(hssi_10g_tx_pcs_low_latency_en),
				.master_clk_sel(hssi_10g_tx_pcs_master_clk_sel),
				.pempty_flag_type(hssi_10g_tx_pcs_pempty_flag_type),
				.pfull_flag_type(hssi_10g_tx_pcs_pfull_flag_type),
				.phcomp_rd_del(hssi_10g_tx_pcs_phcomp_rd_del),
				.pld_if_type(hssi_10g_tx_pcs_pld_if_type),
				.prot_mode(hssi_10g_tx_pcs_prot_mode),
				.pseudo_random(hssi_10g_tx_pcs_pseudo_random),
				.pseudo_seed_a(hssi_10g_tx_pcs_pseudo_seed_a),
				.pseudo_seed_b(hssi_10g_tx_pcs_pseudo_seed_b),
				.random_disp(hssi_10g_tx_pcs_random_disp),
				.rdfifo_clken(hssi_10g_tx_pcs_rdfifo_clken),
				.reconfig_settings(hssi_10g_tx_pcs_reconfig_settings),
				.scrm_bypass(hssi_10g_tx_pcs_scrm_bypass),
				.scrm_clken(hssi_10g_tx_pcs_scrm_clken),
				.scrm_mode(hssi_10g_tx_pcs_scrm_mode),
				.scrm_pipeln(hssi_10g_tx_pcs_scrm_pipeln),
				.sh_err(hssi_10g_tx_pcs_sh_err),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sop_mark(hssi_10g_tx_pcs_sop_mark),
				.stretch_num_stages(hssi_10g_tx_pcs_stretch_num_stages),
				.sup_mode(hssi_10g_tx_pcs_sup_mode),
				.test_mode(hssi_10g_tx_pcs_test_mode),
				.tx_scrm_err(hssi_10g_tx_pcs_tx_scrm_err),
				.tx_scrm_width(hssi_10g_tx_pcs_tx_scrm_width),
				.tx_sh_location(hssi_10g_tx_pcs_tx_sh_location),
				.tx_sm_bypass(hssi_10g_tx_pcs_tx_sm_bypass),
				.tx_sm_pipeln(hssi_10g_tx_pcs_tx_sm_pipeln),
				.tx_testbus_sel(hssi_10g_tx_pcs_tx_testbus_sel),
				.txfifo_empty(hssi_10g_tx_pcs_txfifo_empty),
				.txfifo_full(hssi_10g_tx_pcs_txfifo_full),
				.txfifo_mode(hssi_10g_tx_pcs_txfifo_mode),
				.txfifo_pempty(hssi_10g_tx_pcs_txfifo_pempty),
				.txfifo_pfull(hssi_10g_tx_pcs_txfifo_pfull),
				.wr_clk_sel(hssi_10g_tx_pcs_wr_clk_sel),
				.wrfifo_clken(hssi_10g_tx_pcs_wrfifo_clken)
			) inst_twentynm_hssi_10g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_10g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_10g_tx_pcs_blockselect),
				.distdwn_out_dv(w_hssi_10g_tx_pcs_distdwn_out_dv),
				.distdwn_out_rden(w_hssi_10g_tx_pcs_distdwn_out_rden),
				.distdwn_out_wren(w_hssi_10g_tx_pcs_distdwn_out_wren),
				.distup_out_dv(w_hssi_10g_tx_pcs_distup_out_dv),
				.distup_out_rden(w_hssi_10g_tx_pcs_distup_out_rden),
				.distup_out_wren(w_hssi_10g_tx_pcs_distup_out_wren),
				.tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pma_if(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.tx_control_out_krfec(w_hssi_10g_tx_pcs_tx_control_out_krfec),
				.tx_data_out_krfec(w_hssi_10g_tx_pcs_tx_data_out_krfec),
				.tx_data_valid_out_krfec(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.tx_fec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_fifo_num(w_hssi_10g_tx_pcs_tx_fifo_num),
				.tx_fifo_rd_ptr(w_hssi_10g_tx_pcs_tx_fifo_rd_ptr),
				.tx_fifo_wr_clk(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.tx_fifo_wr_data(w_hssi_10g_tx_pcs_tx_fifo_wr_data),
				.tx_fifo_wr_data_dw(w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw),
				.tx_fifo_wr_en(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.tx_fifo_wr_ptr(w_hssi_10g_tx_pcs_tx_fifo_wr_ptr),
				.tx_fifo_wr_rst_n(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.tx_full(w_hssi_10g_tx_pcs_tx_full),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				.tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.tx_pma_data(w_hssi_10g_tx_pcs_tx_pma_data),
				.tx_pma_gating_val(w_hssi_10g_tx_pcs_tx_pma_gating_val),
				.tx_test_data(w_hssi_10g_tx_pcs_tx_test_data),
				.tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.distdwn_in_dv(in_bond_pcs10g_in_bot[2]),
				.distdwn_in_rden(in_bond_pcs10g_in_bot[4]),
				.distdwn_in_wren(in_bond_pcs10g_in_bot[3]),
				.distup_in_dv(in_bond_pcs10g_in_top[2]),
				.distup_in_rden(in_bond_pcs10g_in_top[4]),
				.distup_in_wren(in_bond_pcs10g_in_top[3]),
				.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.r_tx_diag_word({1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_scrm_word({1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
				.r_tx_skip_word({1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}),
				.r_tx_sync_word({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0}),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.tx_bitslip({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0]}),
				.tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.tx_control({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0]}),
				.tx_control_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0]}),
				.tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0]}),
				.tx_data_in_krfec({w_hssi_krfec_tx_pcs_tx_data_out[63], w_hssi_krfec_tx_pcs_tx_data_out[62], w_hssi_krfec_tx_pcs_tx_data_out[61], w_hssi_krfec_tx_pcs_tx_data_out[60], w_hssi_krfec_tx_pcs_tx_data_out[59], w_hssi_krfec_tx_pcs_tx_data_out[58], w_hssi_krfec_tx_pcs_tx_data_out[57], w_hssi_krfec_tx_pcs_tx_data_out[56], w_hssi_krfec_tx_pcs_tx_data_out[55], w_hssi_krfec_tx_pcs_tx_data_out[54], w_hssi_krfec_tx_pcs_tx_data_out[53], w_hssi_krfec_tx_pcs_tx_data_out[52], w_hssi_krfec_tx_pcs_tx_data_out[51], w_hssi_krfec_tx_pcs_tx_data_out[50], w_hssi_krfec_tx_pcs_tx_data_out[49], w_hssi_krfec_tx_pcs_tx_data_out[48], w_hssi_krfec_tx_pcs_tx_data_out[47], w_hssi_krfec_tx_pcs_tx_data_out[46], w_hssi_krfec_tx_pcs_tx_data_out[45], w_hssi_krfec_tx_pcs_tx_data_out[44], w_hssi_krfec_tx_pcs_tx_data_out[43], w_hssi_krfec_tx_pcs_tx_data_out[42], w_hssi_krfec_tx_pcs_tx_data_out[41], w_hssi_krfec_tx_pcs_tx_data_out[40], w_hssi_krfec_tx_pcs_tx_data_out[39], w_hssi_krfec_tx_pcs_tx_data_out[38], w_hssi_krfec_tx_pcs_tx_data_out[37], w_hssi_krfec_tx_pcs_tx_data_out[36], w_hssi_krfec_tx_pcs_tx_data_out[35], w_hssi_krfec_tx_pcs_tx_data_out[34], w_hssi_krfec_tx_pcs_tx_data_out[33], w_hssi_krfec_tx_pcs_tx_data_out[32], w_hssi_krfec_tx_pcs_tx_data_out[31], w_hssi_krfec_tx_pcs_tx_data_out[30], w_hssi_krfec_tx_pcs_tx_data_out[29], w_hssi_krfec_tx_pcs_tx_data_out[28], w_hssi_krfec_tx_pcs_tx_data_out[27], w_hssi_krfec_tx_pcs_tx_data_out[26], w_hssi_krfec_tx_pcs_tx_data_out[25], w_hssi_krfec_tx_pcs_tx_data_out[24], w_hssi_krfec_tx_pcs_tx_data_out[23], w_hssi_krfec_tx_pcs_tx_data_out[22], w_hssi_krfec_tx_pcs_tx_data_out[21], w_hssi_krfec_tx_pcs_tx_data_out[20], w_hssi_krfec_tx_pcs_tx_data_out[19], w_hssi_krfec_tx_pcs_tx_data_out[18], w_hssi_krfec_tx_pcs_tx_data_out[17], w_hssi_krfec_tx_pcs_tx_data_out[16], w_hssi_krfec_tx_pcs_tx_data_out[15], w_hssi_krfec_tx_pcs_tx_data_out[14], w_hssi_krfec_tx_pcs_tx_data_out[13], w_hssi_krfec_tx_pcs_tx_data_out[12], w_hssi_krfec_tx_pcs_tx_data_out[11], w_hssi_krfec_tx_pcs_tx_data_out[10], w_hssi_krfec_tx_pcs_tx_data_out[9], w_hssi_krfec_tx_pcs_tx_data_out[8], w_hssi_krfec_tx_pcs_tx_data_out[7], w_hssi_krfec_tx_pcs_tx_data_out[6], w_hssi_krfec_tx_pcs_tx_data_out[5], w_hssi_krfec_tx_pcs_tx_data_out[4], w_hssi_krfec_tx_pcs_tx_data_out[3], w_hssi_krfec_tx_pcs_tx_data_out[2], w_hssi_krfec_tx_pcs_tx_data_out[1], w_hssi_krfec_tx_pcs_tx_data_out[0]}),
				.tx_data_reg({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0]}),
				.tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.tx_diag_status({w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1], w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0]}),
				.tx_fifo_rd_data({w_hssi_fifo_tx_pcs_data_out_10g[72], w_hssi_fifo_tx_pcs_data_out_10g[71], w_hssi_fifo_tx_pcs_data_out_10g[70], w_hssi_fifo_tx_pcs_data_out_10g[69], w_hssi_fifo_tx_pcs_data_out_10g[68], w_hssi_fifo_tx_pcs_data_out_10g[67], w_hssi_fifo_tx_pcs_data_out_10g[66], w_hssi_fifo_tx_pcs_data_out_10g[65], w_hssi_fifo_tx_pcs_data_out_10g[64], w_hssi_fifo_tx_pcs_data_out_10g[63], w_hssi_fifo_tx_pcs_data_out_10g[62], w_hssi_fifo_tx_pcs_data_out_10g[61], w_hssi_fifo_tx_pcs_data_out_10g[60], w_hssi_fifo_tx_pcs_data_out_10g[59], w_hssi_fifo_tx_pcs_data_out_10g[58], w_hssi_fifo_tx_pcs_data_out_10g[57], w_hssi_fifo_tx_pcs_data_out_10g[56], w_hssi_fifo_tx_pcs_data_out_10g[55], w_hssi_fifo_tx_pcs_data_out_10g[54], w_hssi_fifo_tx_pcs_data_out_10g[53], w_hssi_fifo_tx_pcs_data_out_10g[52], w_hssi_fifo_tx_pcs_data_out_10g[51], w_hssi_fifo_tx_pcs_data_out_10g[50], w_hssi_fifo_tx_pcs_data_out_10g[49], w_hssi_fifo_tx_pcs_data_out_10g[48], w_hssi_fifo_tx_pcs_data_out_10g[47], w_hssi_fifo_tx_pcs_data_out_10g[46], w_hssi_fifo_tx_pcs_data_out_10g[45], w_hssi_fifo_tx_pcs_data_out_10g[44], w_hssi_fifo_tx_pcs_data_out_10g[43], w_hssi_fifo_tx_pcs_data_out_10g[42], w_hssi_fifo_tx_pcs_data_out_10g[41], w_hssi_fifo_tx_pcs_data_out_10g[40], w_hssi_fifo_tx_pcs_data_out_10g[39], w_hssi_fifo_tx_pcs_data_out_10g[38], w_hssi_fifo_tx_pcs_data_out_10g[37], w_hssi_fifo_tx_pcs_data_out_10g[36], w_hssi_fifo_tx_pcs_data_out_10g[35], w_hssi_fifo_tx_pcs_data_out_10g[34], w_hssi_fifo_tx_pcs_data_out_10g[33], w_hssi_fifo_tx_pcs_data_out_10g[32], w_hssi_fifo_tx_pcs_data_out_10g[31], w_hssi_fifo_tx_pcs_data_out_10g[30], w_hssi_fifo_tx_pcs_data_out_10g[29], w_hssi_fifo_tx_pcs_data_out_10g[28], w_hssi_fifo_tx_pcs_data_out_10g[27], w_hssi_fifo_tx_pcs_data_out_10g[26], w_hssi_fifo_tx_pcs_data_out_10g[25], w_hssi_fifo_tx_pcs_data_out_10g[24], w_hssi_fifo_tx_pcs_data_out_10g[23], w_hssi_fifo_tx_pcs_data_out_10g[22], w_hssi_fifo_tx_pcs_data_out_10g[21], w_hssi_fifo_tx_pcs_data_out_10g[20], w_hssi_fifo_tx_pcs_data_out_10g[19], w_hssi_fifo_tx_pcs_data_out_10g[18], w_hssi_fifo_tx_pcs_data_out_10g[17], w_hssi_fifo_tx_pcs_data_out_10g[16], w_hssi_fifo_tx_pcs_data_out_10g[15], w_hssi_fifo_tx_pcs_data_out_10g[14], w_hssi_fifo_tx_pcs_data_out_10g[13], w_hssi_fifo_tx_pcs_data_out_10g[12], w_hssi_fifo_tx_pcs_data_out_10g[11], w_hssi_fifo_tx_pcs_data_out_10g[10], w_hssi_fifo_tx_pcs_data_out_10g[9], w_hssi_fifo_tx_pcs_data_out_10g[8], w_hssi_fifo_tx_pcs_data_out_10g[7], w_hssi_fifo_tx_pcs_data_out_10g[6], w_hssi_fifo_tx_pcs_data_out_10g[5], w_hssi_fifo_tx_pcs_data_out_10g[4], w_hssi_fifo_tx_pcs_data_out_10g[3], w_hssi_fifo_tx_pcs_data_out_10g[2], w_hssi_fifo_tx_pcs_data_out_10g[1], w_hssi_fifo_tx_pcs_data_out_10g[0]}),
				.tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_10g_reg(),
				.pld_10g_krfec_tx_pld_rst_n_fifo(),
				.pld_10g_krfec_tx_pld_rst_n_reg(),
				.pld_10g_tx_bitslip_reg(),
				.pld_10g_tx_burst_en_exe_reg(),
				.pld_10g_tx_data_valid_10g_reg(),
				.pld_10g_tx_data_valid_fifo(),
				.pld_10g_tx_data_valid_reg(),
				.pld_10g_tx_diag_status_reg(),
				.pld_10g_tx_empty_reg(),
				.pld_10g_tx_fifo_num_reg(),
				.pld_10g_tx_full_fifo(),
				.pld_10g_tx_full_reg(),
				.pld_10g_tx_pempty_reg(),
				.pld_10g_tx_pfull_fifo(),
				.pld_10g_tx_wordslip_exe_reg(),
				.pld_10g_tx_wordslip_reg(),
				.pld_pcs_tx_clk_out_10g_wire(),
				.pld_tx_burst_en_reg(),
				.pld_tx_control_lo_10g_reg(),
				.pld_tx_data_10g_fifo(),
				.pld_tx_data_lo_10g_reg()
			);
		end // if generate
		else begin
				assign w_hssi_10g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_10g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distdwn_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_dv = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_rden = 1'b0;
				assign w_hssi_10g_tx_pcs_distup_out_wren = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_burst_en_exe = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_clk_out_pma_if = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_control_out_krfec[8:0] = 9'b0;
				assign w_hssi_10g_tx_pcs_tx_data_out_krfec[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_data_valid_out_krfec = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_dft_clk_out = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_empty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fec_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72:0] = 73'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_en = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_full = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_master_clk_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_10g_tx_pcs_tx_pempty = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pfull = 1'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_pma_gating_val[63:0] = 64'b0;
				assign w_hssi_10g_tx_pcs_tx_test_data[19:0] = 20'b0;
				assign w_hssi_10g_tx_pcs_tx_wordslip_exe = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_rx_pcs
			twentynm_hssi_8g_rx_pcs #(
				.auto_error_replacement(hssi_8g_rx_pcs_auto_error_replacement),
				.auto_speed_nego(hssi_8g_rx_pcs_auto_speed_nego),
				.bit_reversal(hssi_8g_rx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_rx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_rx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_rx_pcs_bypass_pipeline_reg),
				.byte_deserializer(hssi_8g_rx_pcs_byte_deserializer),
				.cdr_ctrl_rxvalid_mask(hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask),
				.clkcmp_pattern_n(hssi_8g_rx_pcs_clkcmp_pattern_n),
				.clkcmp_pattern_p(hssi_8g_rx_pcs_clkcmp_pattern_p),
				.clock_gate_bds_dec_asn(hssi_8g_rx_pcs_clock_gate_bds_dec_asn),
				.clock_gate_cdr_eidle(hssi_8g_rx_pcs_clock_gate_cdr_eidle),
				.clock_gate_dw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk),
				.clock_gate_dw_rm_rd(hssi_8g_rx_pcs_clock_gate_dw_rm_rd),
				.clock_gate_dw_rm_wr(hssi_8g_rx_pcs_clock_gate_dw_rm_wr),
				.clock_gate_dw_wa(hssi_8g_rx_pcs_clock_gate_dw_wa),
				.clock_gate_pc_rdclk(hssi_8g_rx_pcs_clock_gate_pc_rdclk),
				.clock_gate_sw_pc_wrclk(hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk),
				.clock_gate_sw_rm_rd(hssi_8g_rx_pcs_clock_gate_sw_rm_rd),
				.clock_gate_sw_rm_wr(hssi_8g_rx_pcs_clock_gate_sw_rm_wr),
				.clock_gate_sw_wa(hssi_8g_rx_pcs_clock_gate_sw_wa),
				.clock_observation_in_pld_core(hssi_8g_rx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_rx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_rx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_rx_pcs_ctrl_plane_bonding_distribution),
				.eidle_entry_eios(hssi_8g_rx_pcs_eidle_entry_eios),
				.eidle_entry_iei(hssi_8g_rx_pcs_eidle_entry_iei),
				.eidle_entry_sd(hssi_8g_rx_pcs_eidle_entry_sd),
				.eightb_tenb_decoder(hssi_8g_rx_pcs_eightb_tenb_decoder),
				.err_flags_sel(hssi_8g_rx_pcs_err_flags_sel),
				.fixed_pat_det(hssi_8g_rx_pcs_fixed_pat_det),
				.fixed_pat_num(hssi_8g_rx_pcs_fixed_pat_num),
				.force_signal_detect(hssi_8g_rx_pcs_force_signal_detect),
				.gen3_clk_en(hssi_8g_rx_pcs_gen3_clk_en),
				.gen3_rx_clk_sel(hssi_8g_rx_pcs_gen3_rx_clk_sel),
				.gen3_tx_clk_sel(hssi_8g_rx_pcs_gen3_tx_clk_sel),
				.hip_mode(hssi_8g_rx_pcs_hip_mode),
				.ibm_invalid_code(hssi_8g_rx_pcs_ibm_invalid_code),
				.invalid_code_flag_only(hssi_8g_rx_pcs_invalid_code_flag_only),
				.pad_or_edb_error_replace(hssi_8g_rx_pcs_pad_or_edb_error_replace),
				.pcs_bypass(hssi_8g_rx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_rx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_rx_pcs_phase_compensation_fifo),
				.pipe_if_enable(hssi_8g_rx_pcs_pipe_if_enable),
				.pma_dw(hssi_8g_rx_pcs_pma_dw),
				.polinv_8b10b_dec(hssi_8g_rx_pcs_polinv_8b10b_dec),
				.prot_mode(hssi_8g_rx_pcs_prot_mode),
				.rate_match(hssi_8g_rx_pcs_rate_match),
				.rate_match_del_thres(hssi_8g_rx_pcs_rate_match_del_thres),
				.rate_match_empty_thres(hssi_8g_rx_pcs_rate_match_empty_thres),
				.rate_match_full_thres(hssi_8g_rx_pcs_rate_match_full_thres),
				.rate_match_ins_thres(hssi_8g_rx_pcs_rate_match_ins_thres),
				.rate_match_start_thres(hssi_8g_rx_pcs_rate_match_start_thres),
				.reconfig_settings(hssi_8g_rx_pcs_reconfig_settings),
				.rx_clk2(hssi_8g_rx_pcs_rx_clk2),
				.rx_clk_free_running(hssi_8g_rx_pcs_rx_clk_free_running),
				.rx_pcs_urst(hssi_8g_rx_pcs_rx_pcs_urst),
				.rx_rcvd_clk(hssi_8g_rx_pcs_rx_rcvd_clk),
				.rx_rd_clk(hssi_8g_rx_pcs_rx_rd_clk),
				.rx_refclk(hssi_8g_rx_pcs_rx_refclk),
				.rx_wr_clk(hssi_8g_rx_pcs_rx_wr_clk),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_rx_pcs_sup_mode),
				.symbol_swap(hssi_8g_rx_pcs_symbol_swap),
				.sync_sm_idle_eios(hssi_8g_rx_pcs_sync_sm_idle_eios),
				.test_bus_sel(hssi_8g_rx_pcs_test_bus_sel),
				.tx_rx_parallel_loopback(hssi_8g_rx_pcs_tx_rx_parallel_loopback),
				.wa_boundary_lock_ctrl(hssi_8g_rx_pcs_wa_boundary_lock_ctrl),
				.wa_clk_slip_spacing(hssi_8g_rx_pcs_wa_clk_slip_spacing),
				.wa_det_latency_sync_status_beh(hssi_8g_rx_pcs_wa_det_latency_sync_status_beh),
				.wa_disp_err_flag(hssi_8g_rx_pcs_wa_disp_err_flag),
				.wa_kchar(hssi_8g_rx_pcs_wa_kchar),
				.wa_pd(hssi_8g_rx_pcs_wa_pd),
				.wa_pd_data(hssi_8g_rx_pcs_wa_pd_data),
				.wa_pd_polarity(hssi_8g_rx_pcs_wa_pd_polarity),
				.wa_pld_controlled(hssi_8g_rx_pcs_wa_pld_controlled),
				.wa_renumber_data(hssi_8g_rx_pcs_wa_renumber_data),
				.wa_rgnumber_data(hssi_8g_rx_pcs_wa_rgnumber_data),
				.wa_rknumber_data(hssi_8g_rx_pcs_wa_rknumber_data),
				.wa_rosnumber_data(hssi_8g_rx_pcs_wa_rosnumber_data),
				.wa_rvnumber_data(hssi_8g_rx_pcs_wa_rvnumber_data),
				.wa_sync_sm_ctrl(hssi_8g_rx_pcs_wa_sync_sm_ctrl),
				.wait_cnt(hssi_8g_rx_pcs_wait_cnt)
			) inst_twentynm_hssi_8g_rx_pcs (
				// OUTPUTS
				.a1a2k1k2flag(w_hssi_8g_rx_pcs_a1a2k1k2flag),
				.avmmreaddata(w_hssi_8g_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_rx_pcs_blockselect),
				.chnl_test_bus_out(w_hssi_8g_rx_pcs_chnl_test_bus_out),
				.clock_to_pld(w_hssi_8g_rx_pcs_clock_to_pld),
				.dataout(w_hssi_8g_rx_pcs_dataout),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidle_detected(w_hssi_8g_rx_pcs_eidle_detected),
				.eios_det_cdr_ctrl(w_hssi_8g_rx_pcs_eios_det_cdr_ctrl),
				.g3_rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.g3_rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.gen2ngen1(w_hssi_8g_rx_pcs_gen2ngen1),
				.parallel_rev_loopback(w_hssi_8g_rx_pcs_parallel_rev_loopback),
				.pc_fifo_empty(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.pcfifofull(w_hssi_8g_rx_pcs_pcfifofull),
				.phystatus(w_hssi_8g_rx_pcs_phystatus),
				.pipe_data(w_hssi_8g_rx_pcs_pipe_data),
				.rd_enable_out_chnl_down(w_hssi_8g_rx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_rx_pcs_rd_enable_out_chnl_up),
				.rd_ptr1_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo),
				.rd_ptr2_rx_rmfifo(w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo),
				.rd_ptr_rx_phfifo(w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.reset_pc_ptrs_out_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down),
				.reset_pc_ptrs_out_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up),
				.rm_fifo_empty(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.rm_fifo_full(w_hssi_8g_rx_pcs_rm_fifo_full),
				.rx_blk_start(w_hssi_8g_rx_pcs_rx_blk_start),
				.rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.rx_data_valid(w_hssi_8g_rx_pcs_rx_data_valid),
				.rx_div_sync_out_chnl_down(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down),
				.rx_div_sync_out_chnl_up(w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up),
				.rx_pipe_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.rx_pipe_soft_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rx_pma_clk_gen3(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_rcvd_clk_gen3(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_rstn_sync2wrfifo_8g(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.rx_sync_hdr(w_hssi_8g_rx_pcs_rx_sync_hdr),
				.rx_we_out_chnl_down(w_hssi_8g_rx_pcs_rx_we_out_chnl_down),
				.rx_we_out_chnl_up(w_hssi_8g_rx_pcs_rx_we_out_chnl_up),
				.rxstatus(w_hssi_8g_rx_pcs_rxstatus),
				.rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.word_align_boundary(w_hssi_8g_rx_pcs_word_align_boundary),
				.wr_clk_rx_phfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_rx_phfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_rx_rmfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_rx_rmfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_data_rx_phfifo(w_hssi_8g_rx_pcs_wr_data_rx_phfifo),
				.wr_data_rx_rmfifo(w_hssi_8g_rx_pcs_wr_data_rx_rmfifo),
				.wr_en_rx_phfifo(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_rx_rmfifo(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_rx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_rx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_rx_phfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo),
				.wr_ptr_rx_rmfifo(w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo),
				.wr_rst_n_rx_phfifo(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_rx_rmfifo(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				// INPUTS
				.a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bit_reversal_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.datain({w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1], w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0]}),
				.disable_pc_fifo_byte_serdes(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4]),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.eidleinfersel({w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1], w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0]}),
				.eios_detected_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.enable_comma_detect(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.gen3_clk_sel(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.hrd_rst(1'b0),
				.inferred_rxvalid_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.pc_fifo_rd_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.pc_fifo_wrdisable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.phystatus_int(w_hssi_pipe_gen1_2_phystatus),
				.phystatus_pcs_gen3(w_hssi_pipe_gen3_phystatus),
				.pipe_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.polarity_inversion(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.rd_data1_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0]}),
				.rd_data2_rx_rmfifo({w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1], w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0]}),
				.rd_data_rx_phfifo({w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[3]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[3]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.reset_pc_ptrs_asn(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5]),
				.reset_pc_ptrs_in_chnl_down(in_bond_pcs8g_in_bot[12]),
				.reset_pc_ptrs_in_chnl_up(in_bond_pcs8g_in_top[12]),
				.reset_ppm_cntrs_pcs_pma(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7]),
				.rm_fifo_read_enable(1'b0),
				.rm_fifo_write_enable(1'b0),
				.rx_blk_start_pcs_gen3({w_hssi_pipe_gen3_rx_blk_start[3], w_hssi_pipe_gen3_rx_blk_start[2], w_hssi_pipe_gen3_rx_blk_start[1], w_hssi_pipe_gen3_rx_blk_start[0]}),
				.rx_data_pcs_gen3({w_hssi_pipe_gen3_rxd_8gpcs_out[63], w_hssi_pipe_gen3_rxd_8gpcs_out[62], w_hssi_pipe_gen3_rxd_8gpcs_out[61], w_hssi_pipe_gen3_rxd_8gpcs_out[60], w_hssi_pipe_gen3_rxd_8gpcs_out[59], w_hssi_pipe_gen3_rxd_8gpcs_out[58], w_hssi_pipe_gen3_rxd_8gpcs_out[57], w_hssi_pipe_gen3_rxd_8gpcs_out[56], w_hssi_pipe_gen3_rxd_8gpcs_out[55], w_hssi_pipe_gen3_rxd_8gpcs_out[54], w_hssi_pipe_gen3_rxd_8gpcs_out[53], w_hssi_pipe_gen3_rxd_8gpcs_out[52], w_hssi_pipe_gen3_rxd_8gpcs_out[51], w_hssi_pipe_gen3_rxd_8gpcs_out[50], w_hssi_pipe_gen3_rxd_8gpcs_out[49], w_hssi_pipe_gen3_rxd_8gpcs_out[48], w_hssi_pipe_gen3_rxd_8gpcs_out[47], w_hssi_pipe_gen3_rxd_8gpcs_out[46], w_hssi_pipe_gen3_rxd_8gpcs_out[45], w_hssi_pipe_gen3_rxd_8gpcs_out[44], w_hssi_pipe_gen3_rxd_8gpcs_out[43], w_hssi_pipe_gen3_rxd_8gpcs_out[42], w_hssi_pipe_gen3_rxd_8gpcs_out[41], w_hssi_pipe_gen3_rxd_8gpcs_out[40], w_hssi_pipe_gen3_rxd_8gpcs_out[39], w_hssi_pipe_gen3_rxd_8gpcs_out[38], w_hssi_pipe_gen3_rxd_8gpcs_out[37], w_hssi_pipe_gen3_rxd_8gpcs_out[36], w_hssi_pipe_gen3_rxd_8gpcs_out[35], w_hssi_pipe_gen3_rxd_8gpcs_out[34], w_hssi_pipe_gen3_rxd_8gpcs_out[33], w_hssi_pipe_gen3_rxd_8gpcs_out[32], w_hssi_pipe_gen3_rxd_8gpcs_out[31], w_hssi_pipe_gen3_rxd_8gpcs_out[30], w_hssi_pipe_gen3_rxd_8gpcs_out[29], w_hssi_pipe_gen3_rxd_8gpcs_out[28], w_hssi_pipe_gen3_rxd_8gpcs_out[27], w_hssi_pipe_gen3_rxd_8gpcs_out[26], w_hssi_pipe_gen3_rxd_8gpcs_out[25], w_hssi_pipe_gen3_rxd_8gpcs_out[24], w_hssi_pipe_gen3_rxd_8gpcs_out[23], w_hssi_pipe_gen3_rxd_8gpcs_out[22], w_hssi_pipe_gen3_rxd_8gpcs_out[21], w_hssi_pipe_gen3_rxd_8gpcs_out[20], w_hssi_pipe_gen3_rxd_8gpcs_out[19], w_hssi_pipe_gen3_rxd_8gpcs_out[18], w_hssi_pipe_gen3_rxd_8gpcs_out[17], w_hssi_pipe_gen3_rxd_8gpcs_out[16], w_hssi_pipe_gen3_rxd_8gpcs_out[15], w_hssi_pipe_gen3_rxd_8gpcs_out[14], w_hssi_pipe_gen3_rxd_8gpcs_out[13], w_hssi_pipe_gen3_rxd_8gpcs_out[12], w_hssi_pipe_gen3_rxd_8gpcs_out[11], w_hssi_pipe_gen3_rxd_8gpcs_out[10], w_hssi_pipe_gen3_rxd_8gpcs_out[9], w_hssi_pipe_gen3_rxd_8gpcs_out[8], w_hssi_pipe_gen3_rxd_8gpcs_out[7], w_hssi_pipe_gen3_rxd_8gpcs_out[6], w_hssi_pipe_gen3_rxd_8gpcs_out[5], w_hssi_pipe_gen3_rxd_8gpcs_out[4], w_hssi_pipe_gen3_rxd_8gpcs_out[3], w_hssi_pipe_gen3_rxd_8gpcs_out[2], w_hssi_pipe_gen3_rxd_8gpcs_out[1], w_hssi_pipe_gen3_rxd_8gpcs_out[0]}),
				.rx_data_valid_pcs_gen3({w_hssi_pipe_gen3_rxdataskip[3], w_hssi_pipe_gen3_rxdataskip[2], w_hssi_pipe_gen3_rxdataskip[1], w_hssi_pipe_gen3_rxdataskip[0]}),
				.rx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[1], in_bond_pcs8g_in_bot[0]}),
				.rx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[1], in_bond_pcs8g_in_top[0]}),
				.rx_pcs_rst(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.rx_sync_hdr_pcs_gen3({w_hssi_pipe_gen3_rx_sync_hdr[1], w_hssi_pipe_gen3_rx_sync_hdr[0]}),
				.rx_we_in_chnl_down({in_bond_pcs8g_in_bot[5], in_bond_pcs8g_in_bot[4]}),
				.rx_we_in_chnl_up({in_bond_pcs8g_in_top[5], in_bond_pcs8g_in_top[4]}),
				.rxstatus_int({w_hssi_pipe_gen1_2_rxstatus[2], w_hssi_pipe_gen1_2_rxstatus[1], w_hssi_pipe_gen1_2_rxstatus[0]}),
				.rxstatus_pcs_gen3({w_hssi_pipe_gen3_rxstatus[2], w_hssi_pipe_gen3_rxstatus[1], w_hssi_pipe_gen3_rxstatus[0]}),
				.rxvalid_int(w_hssi_pipe_gen1_2_rxvalid),
				.rxvalid_pcs_gen3(w_hssi_pipe_gen3_rxvalid),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.sig_det_from_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_ctrlplane_testbus({w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1], w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0]}),
				.tx_div_sync({w_hssi_8g_tx_pcs_tx_div_sync[1], w_hssi_8g_tx_pcs_tx_div_sync[0]}),
				.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.tx_testbus({w_hssi_8g_tx_pcs_tx_testbus[19], w_hssi_8g_tx_pcs_tx_testbus[18], w_hssi_8g_tx_pcs_tx_testbus[17], w_hssi_8g_tx_pcs_tx_testbus[16], w_hssi_8g_tx_pcs_tx_testbus[15], w_hssi_8g_tx_pcs_tx_testbus[14], w_hssi_8g_tx_pcs_tx_testbus[13], w_hssi_8g_tx_pcs_tx_testbus[12], w_hssi_8g_tx_pcs_tx_testbus[11], w_hssi_8g_tx_pcs_tx_testbus[10], w_hssi_8g_tx_pcs_tx_testbus[9], w_hssi_8g_tx_pcs_tx_testbus[8], w_hssi_8g_tx_pcs_tx_testbus[7], w_hssi_8g_tx_pcs_tx_testbus[6], w_hssi_8g_tx_pcs_tx_testbus[5], w_hssi_8g_tx_pcs_tx_testbus[4], w_hssi_8g_tx_pcs_tx_testbus[3], w_hssi_8g_tx_pcs_tx_testbus[2], w_hssi_8g_tx_pcs_tx_testbus[1], w_hssi_8g_tx_pcs_tx_testbus[0]}),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[2]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[2]),
				
				// UNUSED
				.byte_deserializer_pcs_clk_div_by_2_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pcs_clk_div_by_2_txclk_wire(),
				.byte_deserializer_pcs_clk_div_by_2_wire(),
				.byte_deserializer_pcs_clk_div_by_4_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_2_reg(),
				.byte_deserializer_pld_clk_div_by_2_txclk_reg(),
				.byte_deserializer_pld_clk_div_by_4_txclk_reg(),
				.pld_8g_a1a2_k1k2_flag_reg(),
				.pld_8g_a1a2_k1k2_flag_txclk_reg(),
				.pld_8g_a1a2_size_reg(),
				.pld_8g_a1a2_size_txclk_reg(),
				.pld_8g_bitloc_rev_en_reg(),
				.pld_8g_bitloc_rev_en_txclk_reg(),
				.pld_8g_byte_rev_en_reg(),
				.pld_8g_byte_rev_en_txclk_reg(),
				.pld_8g_elecidle_reg(),
				.pld_8g_empty_rmf_lowlatency_reg(),
				.pld_8g_empty_rmf_lowlatency_txclk_reg(),
				.pld_8g_empty_rmf_reg(),
				.pld_8g_empty_rmf_txclk_reg(),
				.pld_8g_empty_rx_fifo(),
				.pld_8g_empty_rx_reg(),
				.pld_8g_empty_rx_txclk_reg(),
				.pld_8g_encdt_reg(),
				.pld_8g_encdt_txclk_reg(),
				.pld_8g_full_rmf_reg(),
				.pld_8g_full_rmf_txclk_reg(),
				.pld_8g_full_rx_fifo(),
				.pld_8g_full_rx_reg(),
				.pld_8g_full_rx_txclk_reg(),
				.pld_8g_g3_rx_pld_rst_n_reg(),
				.pld_8g_g3_rx_pld_rst_n_txclk_reg(),
				.pld_8g_rxelecidle_txclk_reg(),
				.pld_8g_rxpolarity_reg(),
				.pld_8g_rxpolarity_txclk_reg(),
				.pld_8g_wa_boundary_reg(),
				.pld_8g_wrdisable_rx_reg(),
				.pld_8g_wrdisable_rx_txclk_reg(),
				.pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_rx_clk_out_8g_txclk_wire(),
				.pld_pcs_rx_clk_out_8g_wire(),
				.pld_rx_control_8g_reg(),
				.pld_rx_control_8g_txclk_reg(),
				.pld_rx_data_8g_reg(),
				.pld_rx_data_8g_txclk_reg(),
				.pld_syncsm_en_reg(),
				.pld_syncsm_en_txclk_reg(),
				.rm_fifo_partial_empty(),
				.rm_fifo_partial_full(),
				.sta_rx_clk2_by2_1(),
				.sta_rx_clk2_by2_1_out(),
				.sta_rx_clk2_by2_2(),
				.sta_rx_clk2_by2_2_out(),
				.sta_rx_clk2_by4_1(),
				.sta_rx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_rx_pcs_a1a2k1k2flag[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_rx_pcs_chnl_test_bus_out[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_clock_to_pld = 1'b0;
				assign w_hssi_8g_rx_pcs_dataout[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_dis_pc_byte = 1'b0;
				assign w_hssi_8g_rx_pcs_eidle_detected = 1'b0;
				assign w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_pma_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn = 1'b0;
				assign w_hssi_8g_rx_pcs_gen2ngen1 = 1'b0;
				assign w_hssi_8g_rx_pcs_parallel_rev_loopback[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_pc_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_pcfifofull = 1'b0;
				assign w_hssi_8g_rx_pcs_phystatus = 1'b0;
				assign w_hssi_8g_rx_pcs_pipe_data[63:0] = 64'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_empty = 1'b0;
				assign w_hssi_8g_rx_pcs_rm_fifo_full = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_clkslip = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_data_valid[3:0] = 4'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_pma_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3 = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g = 1'b0;
				assign w_hssi_8g_rx_pcs_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_rx_pcs_rxstatus[2:0] = 3'b0;
				assign w_hssi_8g_rx_pcs_rxvalid = 1'b0;
				assign w_hssi_8g_rx_pcs_signal_detect_out = 1'b0;
				assign w_hssi_8g_rx_pcs_word_align_boundary[4:0] = 5'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79:0] = 80'b0;
				assign w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31:0] = 32'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_en_rx_rmfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19:0] = 20'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo = 1'b0;
				assign w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_8g_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_8g_tx_pcs
			twentynm_hssi_8g_tx_pcs #(
				.auto_speed_nego_gen2(hssi_8g_tx_pcs_auto_speed_nego_gen2),
				.bit_reversal(hssi_8g_tx_pcs_bit_reversal),
				.bonding_dft_en(hssi_8g_tx_pcs_bonding_dft_en),
				.bonding_dft_val(hssi_8g_tx_pcs_bonding_dft_val),
				.bypass_pipeline_reg(hssi_8g_tx_pcs_bypass_pipeline_reg),
				.byte_serializer(hssi_8g_tx_pcs_byte_serializer),
				.clock_gate_bs_enc(hssi_8g_tx_pcs_clock_gate_bs_enc),
				.clock_gate_dw_fifowr(hssi_8g_tx_pcs_clock_gate_dw_fifowr),
				.clock_gate_fiford(hssi_8g_tx_pcs_clock_gate_fiford),
				.clock_gate_sw_fifowr(hssi_8g_tx_pcs_clock_gate_sw_fifowr),
				.clock_observation_in_pld_core(hssi_8g_tx_pcs_clock_observation_in_pld_core),
				.ctrl_plane_bonding_compensation(hssi_8g_tx_pcs_ctrl_plane_bonding_compensation),
				.ctrl_plane_bonding_consumption(hssi_8g_tx_pcs_ctrl_plane_bonding_consumption),
				.ctrl_plane_bonding_distribution(hssi_8g_tx_pcs_ctrl_plane_bonding_distribution),
				.data_selection_8b10b_encoder_input(hssi_8g_tx_pcs_data_selection_8b10b_encoder_input),
				.dynamic_clk_switch(hssi_8g_tx_pcs_dynamic_clk_switch),
				.eightb_tenb_disp_ctrl(hssi_8g_tx_pcs_eightb_tenb_disp_ctrl),
				.eightb_tenb_encoder(hssi_8g_tx_pcs_eightb_tenb_encoder),
				.force_echar(hssi_8g_tx_pcs_force_echar),
				.force_kchar(hssi_8g_tx_pcs_force_kchar),
				.gen3_tx_clk_sel(hssi_8g_tx_pcs_gen3_tx_clk_sel),
				.gen3_tx_pipe_clk_sel(hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel),
				.hip_mode(hssi_8g_tx_pcs_hip_mode),
				.pcs_bypass(hssi_8g_tx_pcs_pcs_bypass),
				.phase_comp_rdptr(hssi_8g_tx_pcs_phase_comp_rdptr),
				.phase_compensation_fifo(hssi_8g_tx_pcs_phase_compensation_fifo),
				.phfifo_write_clk_sel(hssi_8g_tx_pcs_phfifo_write_clk_sel),
				.pma_dw(hssi_8g_tx_pcs_pma_dw),
				.prot_mode(hssi_8g_tx_pcs_prot_mode),
				.reconfig_settings(hssi_8g_tx_pcs_reconfig_settings),
				.refclk_b_clk_sel(hssi_8g_tx_pcs_refclk_b_clk_sel),
				.revloop_back_rm(hssi_8g_tx_pcs_revloop_back_rm),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sup_mode(hssi_8g_tx_pcs_sup_mode),
				.symbol_swap(hssi_8g_tx_pcs_symbol_swap),
				.tx_bitslip(hssi_8g_tx_pcs_tx_bitslip),
				.tx_compliance_controlled_disparity(hssi_8g_tx_pcs_tx_compliance_controlled_disparity),
				.tx_fast_pld_reg(hssi_8g_tx_pcs_tx_fast_pld_reg),
				.txclk_freerun(hssi_8g_tx_pcs_txclk_freerun),
				.txpcs_urst(hssi_8g_tx_pcs_txpcs_urst)
			) inst_twentynm_hssi_8g_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_8g_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_8g_tx_pcs_blockselect),
				.clk_out(w_hssi_8g_tx_pcs_clk_out),
				.clk_out_gen3(w_hssi_8g_tx_pcs_clk_out_gen3),
				.dataout(w_hssi_8g_tx_pcs_dataout),
				.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
				.fifo_select_out_chnl_down(w_hssi_8g_tx_pcs_fifo_select_out_chnl_down),
				.fifo_select_out_chnl_up(w_hssi_8g_tx_pcs_fifo_select_out_chnl_up),
				.g3_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.g3_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
				.non_gray_eidleinfersel(w_hssi_8g_tx_pcs_non_gray_eidleinfersel),
				.ph_fifo_overflow(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.ph_fifo_underflow(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.phfifo_txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.phfifo_txmargin(w_hssi_8g_tx_pcs_phfifo_txmargin),
				.phfifo_txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				.pipe_en_rev_parallel_lpbk_out(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.pipe_power_down_out(w_hssi_8g_tx_pcs_pipe_power_down_out),
				.pipe_tx_clk_out_gen3(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pmaif_asn_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.rd_enable_out_chnl_down(w_hssi_8g_tx_pcs_rd_enable_out_chnl_down),
				.rd_enable_out_chnl_up(w_hssi_8g_tx_pcs_rd_enable_out_chnl_up),
				.rd_ptr_tx_phfifo(w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rxpolarity_int(w_hssi_8g_tx_pcs_rxpolarity_int),
				.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
				.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
				.tx_blk_start_out(w_hssi_8g_tx_pcs_tx_blk_start_out),
				.tx_clk_out_8g_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.tx_clk_out_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.tx_ctrlplane_testbus(w_hssi_8g_tx_pcs_tx_ctrlplane_testbus),
				.tx_data_out(w_hssi_8g_tx_pcs_tx_data_out),
				.tx_data_valid_out(w_hssi_8g_tx_pcs_tx_data_valid_out),
				.tx_datak_out(w_hssi_8g_tx_pcs_tx_datak_out),
				.tx_detect_rxloopback_int(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.tx_div_sync(w_hssi_8g_tx_pcs_tx_div_sync),
				.tx_div_sync_out_chnl_down(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down),
				.tx_div_sync_out_chnl_up(w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up),
				.tx_pipe_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.tx_pipe_electidle(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_soft_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.tx_sync_hdr_out(w_hssi_8g_tx_pcs_tx_sync_hdr_out),
				.tx_testbus(w_hssi_8g_tx_pcs_tx_testbus),
				.txcompliance_out(w_hssi_8g_tx_pcs_txcompliance_out),
				.txelecidle_out(w_hssi_8g_tx_pcs_txelecidle_out),
				.wr_clk_tx_phfifo_dw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_tx_phfifo_sw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_data_tx_phfifo(w_hssi_8g_tx_pcs_wr_data_tx_phfifo),
				.wr_en_tx_phfifo(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_enable_out_chnl_down(w_hssi_8g_tx_pcs_wr_enable_out_chnl_down),
				.wr_enable_out_chnl_up(w_hssi_8g_tx_pcs_wr_enable_out_chnl_up),
				.wr_ptr_tx_phfifo(w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo),
				.wr_rst_n_tx_phfifo(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.bitslip_boundary_select({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0]}),
				.clk_sel_gen3(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]),
				.coreclk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.datain({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.detectrxloopin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
				.eidleinfersel({w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1], w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0]}),
				.en_rev_parallel_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.fifo_select_in_chnl_down({in_bond_pcs8g_in_bot[11], in_bond_pcs8g_in_bot[10]}),
				.fifo_select_in_chnl_up({in_bond_pcs8g_in_top[11], in_bond_pcs8g_in_top[10]}),
				.hrdrst(1'b0),
				.pcs_rst(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]),
				.ph_fifo_rd_disable(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.pipe_en_rev_parallel_lpbk_in(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.pipe_tx_deemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.pipe_tx_margin({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0]}),
				.powerdn({w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0]}),
				.rate_switch(w_hssi_8g_rx_pcs_gen2ngen1),
				.rd_data_tx_phfifo({w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1], w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0]}),
				.rd_enable_in_chnl_down(in_bond_pcs8g_in_bot[9]),
				.rd_enable_in_chnl_up(in_bond_pcs8g_in_top[9]),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
				.reset_pc_ptrs_in_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
				.reset_pc_ptrs_in_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
				.rev_parallel_lpbk_data({w_hssi_8g_rx_pcs_parallel_rev_loopback[19], w_hssi_8g_rx_pcs_parallel_rev_loopback[18], w_hssi_8g_rx_pcs_parallel_rev_loopback[17], w_hssi_8g_rx_pcs_parallel_rev_loopback[16], w_hssi_8g_rx_pcs_parallel_rev_loopback[15], w_hssi_8g_rx_pcs_parallel_rev_loopback[14], w_hssi_8g_rx_pcs_parallel_rev_loopback[13], w_hssi_8g_rx_pcs_parallel_rev_loopback[12], w_hssi_8g_rx_pcs_parallel_rev_loopback[11], w_hssi_8g_rx_pcs_parallel_rev_loopback[10], w_hssi_8g_rx_pcs_parallel_rev_loopback[9], w_hssi_8g_rx_pcs_parallel_rev_loopback[8], w_hssi_8g_rx_pcs_parallel_rev_loopback[7], w_hssi_8g_rx_pcs_parallel_rev_loopback[6], w_hssi_8g_rx_pcs_parallel_rev_loopback[5], w_hssi_8g_rx_pcs_parallel_rev_loopback[4], w_hssi_8g_rx_pcs_parallel_rev_loopback[3], w_hssi_8g_rx_pcs_parallel_rev_loopback[2], w_hssi_8g_rx_pcs_parallel_rev_loopback[1], w_hssi_8g_rx_pcs_parallel_rev_loopback[0]}),
				.rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.tx_blk_start({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0]}),
				.tx_data_valid({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0]}),
				.tx_div_sync_in_chnl_down({in_bond_pcs8g_in_bot[7], in_bond_pcs8g_in_bot[6]}),
				.tx_div_sync_in_chnl_up({in_bond_pcs8g_in_top[7], in_bond_pcs8g_in_top[6]}),
				.tx_pcs_reset(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.tx_sync_hdr({w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0]}),
				.txd_fast_reg({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0]}),
				.txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.wr_enable_in_chnl_down(in_bond_pcs8g_in_bot[8]),
				.wr_enable_in_chnl_up(in_bond_pcs8g_in_top[8]),
				.wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				
				// UNUSED
				.byte_serializer_pcs_clk_div_by_2_reg(),
				.byte_serializer_pcs_clk_div_by_2_wire(),
				.byte_serializer_pcs_clk_div_by_4_reg(),
				.byte_serializer_pld_clk_div_by_2_reg(),
				.byte_serializer_pld_clk_div_by_4_reg(),
				.pld_8g_empty_tx_fifo(),
				.pld_8g_empty_tx_reg(),
				.pld_8g_full_tx_fifo(),
				.pld_8g_full_tx_reg(),
				.pld_8g_g3_tx_pld_rst_n_reg(),
				.pld_8g_rddisable_tx_reg(),
				.pld_8g_tx_boundary_sel_reg(),
				.pld_pcs_tx_clk_out_8g_div_by_2_wire(),
				.pld_pcs_tx_clk_out_8g_wire(),
				.pld_tx_data_8g_fifo(),
				.pld_tx_data_lo_8g_reg(),
				.sta_tx_clk2_by2_1(),
				.sta_tx_clk2_by2_1_out(),
				.sta_tx_clk2_by4_1(),
				.sta_tx_clk2_by4_1_out()
			);
		end // if generate
		else begin
				assign w_hssi_8g_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_blockselect = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_dataout[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_dyn_clk_switch_n = 1'b1;		// Override default tieoff
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_g3_tx_pma_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_overflow = 1'b0;
				assign w_hssi_8g_tx_pcs_ph_fifo_underflow = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txdeemph = 1'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txmargin[2:0] = 3'b0;
				assign w_hssi_8g_tx_pcs_phfifo_txswing = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out = 1'b0;
				assign w_hssi_8g_tx_pcs_pipe_power_down_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3 = 1'b0;
				assign w_hssi_8g_tx_pcs_pmaif_asn_rstn = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_refclk_b = 1'b0;
				assign w_hssi_8g_tx_pcs_refclk_b_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_rxpolarity_int = 1'b0;
				assign w_hssi_8g_tx_pcs_soft_reset_wclk1_n = 1'b0;
				assign w_hssi_8g_tx_pcs_sw_fifo_wr_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_blk_start_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_out_pmaif = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_tx_data_out[31:0] = 32'b0;
				assign w_hssi_8g_tx_pcs_tx_data_valid_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_datak_out[3:0] = 4'b0;
				assign w_hssi_8g_tx_pcs_tx_detect_rxloopback_int = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_electidle = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_pipe_soft_reset = 1'b0;
				assign w_hssi_8g_tx_pcs_tx_sync_hdr_out[1:0] = 2'b0;
				assign w_hssi_8g_tx_pcs_tx_testbus[19:0] = 20'b0;
				assign w_hssi_8g_tx_pcs_txcompliance_out = 1'b0;
				assign w_hssi_8g_tx_pcs_txelecidle_out = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63:0] = 64'b0;
				assign w_hssi_8g_tx_pcs_wr_en_tx_phfifo = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_down = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_enable_out_chnl_up = 1'b0;
				assign w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7:0] = 8'b0;
				assign w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pcs_pma_interface
			twentynm_hssi_common_pcs_pma_interface #(
				.asn_clk_enable(hssi_common_pcs_pma_interface_asn_clk_enable),
				.asn_enable(hssi_common_pcs_pma_interface_asn_enable),
				.block_sel(hssi_common_pcs_pma_interface_block_sel),
				.bypass_early_eios(hssi_common_pcs_pma_interface_bypass_early_eios),
				.bypass_pcie_switch(hssi_common_pcs_pma_interface_bypass_pcie_switch),
				.bypass_pma_ltr(hssi_common_pcs_pma_interface_bypass_pma_ltr),
				.bypass_pma_sw_done(hssi_common_pcs_pma_interface_bypass_pma_sw_done),
				.bypass_ppm_lock(hssi_common_pcs_pma_interface_bypass_ppm_lock),
				.bypass_send_syncp_fbkp(hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp),
				.bypass_txdetectrx(hssi_common_pcs_pma_interface_bypass_txdetectrx),
				.cdr_control(hssi_common_pcs_pma_interface_cdr_control),
				.cid_enable(hssi_common_pcs_pma_interface_cid_enable),
				.cp_cons_sel(hssi_common_pcs_pma_interface_cp_cons_sel),
				.cp_dwn_mstr(hssi_common_pcs_pma_interface_cp_dwn_mstr),
				.cp_up_mstr(hssi_common_pcs_pma_interface_cp_up_mstr),
				.ctrl_plane_bonding(hssi_common_pcs_pma_interface_ctrl_plane_bonding),
				.data_mask_count(hssi_common_pcs_pma_interface_data_mask_count),
				.data_mask_count_multi(hssi_common_pcs_pma_interface_data_mask_count_multi),
				.dft_observation_clock_selection(hssi_common_pcs_pma_interface_dft_observation_clock_selection),
				.early_eios_counter(hssi_common_pcs_pma_interface_early_eios_counter),
				.force_freqdet(hssi_common_pcs_pma_interface_force_freqdet),
				.free_run_clk_enable(hssi_common_pcs_pma_interface_free_run_clk_enable),
				.ignore_sigdet_g23(hssi_common_pcs_pma_interface_ignore_sigdet_g23),
				.pc_en_counter(hssi_common_pcs_pma_interface_pc_en_counter),
				.pc_rst_counter(hssi_common_pcs_pma_interface_pc_rst_counter),
				.pcie_hip_mode(hssi_common_pcs_pma_interface_pcie_hip_mode),
				.ph_fifo_reg_mode(hssi_common_pcs_pma_interface_ph_fifo_reg_mode),
				.phfifo_flush_wait(hssi_common_pcs_pma_interface_phfifo_flush_wait),
				.pipe_if_g3pcs(hssi_common_pcs_pma_interface_pipe_if_g3pcs),
				.pma_done_counter(hssi_common_pcs_pma_interface_pma_done_counter),
				.pma_if_dft_en(hssi_common_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_common_pcs_pma_interface_pma_if_dft_val),
				.ppm_cnt_rst(hssi_common_pcs_pma_interface_ppm_cnt_rst),
				.ppm_deassert_early(hssi_common_pcs_pma_interface_ppm_deassert_early),
				.ppm_det_buckets(hssi_common_pcs_pma_interface_ppm_det_buckets),
				.ppm_gen1_2_cnt(hssi_common_pcs_pma_interface_ppm_gen1_2_cnt),
				.ppm_post_eidle_delay(hssi_common_pcs_pma_interface_ppm_post_eidle_delay),
				.ppmsel(hssi_common_pcs_pma_interface_ppmsel),
				.prot_mode(hssi_common_pcs_pma_interface_prot_mode),
				.reconfig_settings(hssi_common_pcs_pma_interface_reconfig_settings),
				.rxvalid_mask(hssi_common_pcs_pma_interface_rxvalid_mask),
				.sigdet_wait_counter(hssi_common_pcs_pma_interface_sigdet_wait_counter),
				.sigdet_wait_counter_multi(hssi_common_pcs_pma_interface_sigdet_wait_counter_multi),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sim_mode(hssi_common_pcs_pma_interface_sim_mode),
				.spd_chg_rst_wait_cnt_en(hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en),
				.sup_mode(hssi_common_pcs_pma_interface_sup_mode),
				.testout_sel(hssi_common_pcs_pma_interface_testout_sel),
				.wait_clk_on_off_timer(hssi_common_pcs_pma_interface_wait_clk_on_off_timer),
				.wait_pipe_synchronizing(hssi_common_pcs_pma_interface_wait_pipe_synchronizing),
				.wait_send_syncp_fbkp(hssi_common_pcs_pma_interface_wait_send_syncp_fbkp)
			) inst_twentynm_hssi_common_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_common_pcs_pma_interface_blockselect),
				.int_pmaif_8g_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in),
				.int_pmaif_8g_eios_detected(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
				.int_pmaif_8g_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
				.int_pmaif_8g_power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.int_pmaif_g3_pcs_asn_bundling_in(w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in),
				.int_pmaif_pldif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pmaif_pldif_pcie_sw_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done),
				.int_pmaif_pldif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pmaif_pldif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pmaif_pldif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pmaif_pldif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pmaif_pldif_pma_reserved_in(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in),
				.int_pmaif_pldif_test_out(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out),
				.int_pmaif_pldif_testbus(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus),
				.pma_adapt_start(w_hssi_common_pcs_pma_interface_pma_adapt_start),
				.pma_atpg_los_en_n(w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n),
				.pma_csr_test_dis(w_hssi_common_pcs_pma_interface_pma_csr_test_dis),
				.pma_current_coeff(w_hssi_common_pcs_pma_interface_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_common_pcs_pma_interface_pma_current_rxpreset),
				.pma_early_eios(w_hssi_common_pcs_pma_interface_pma_early_eios),
				.pma_interface_select(w_hssi_common_pcs_pma_interface_pma_interface_select),
				.pma_ltd_b(w_hssi_common_pcs_pma_interface_pma_ltd_b),
				.pma_ltr(w_hssi_common_pcs_pma_interface_pma_ltr),
				.pma_nfrzdrv(w_hssi_common_pcs_pma_interface_pma_nfrzdrv),
				.pma_nrpi_freeze(w_hssi_common_pcs_pma_interface_pma_nrpi_freeze),
				.pma_pcie_switch(w_hssi_common_pcs_pma_interface_pma_pcie_switch),
				.pma_ppm_lock(w_hssi_common_pcs_pma_interface_pma_ppm_lock),
				.pma_reserved_out(w_hssi_common_pcs_pma_interface_pma_reserved_out),
				.pma_rs_lpbk_b(w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b),
				.pma_rx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup),
				.pma_scan_mode_n(w_hssi_common_pcs_pma_interface_pma_scan_mode_n),
				.pma_scan_shift_n(w_hssi_common_pcs_pma_interface_pma_scan_shift_n),
				.pma_tx_bitslip(w_hssi_common_pcs_pma_interface_pma_tx_bitslip),
				.pma_tx_bonding_rstb(w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb),
				.pma_tx_qpi_pulldn(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn),
				.pma_tx_qpi_pullup(w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup),
				.pma_tx_txdetectrx(w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx),
				.pmaif_bundling_out_down(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down),
				.pmaif_bundling_out_up(w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_8g_current_coeff({w_hssi_pipe_gen1_2_current_coeff[17], w_hssi_pipe_gen1_2_current_coeff[16], w_hssi_pipe_gen1_2_current_coeff[15], w_hssi_pipe_gen1_2_current_coeff[14], w_hssi_pipe_gen1_2_current_coeff[13], w_hssi_pipe_gen1_2_current_coeff[12], w_hssi_pipe_gen1_2_current_coeff[11], w_hssi_pipe_gen1_2_current_coeff[10], w_hssi_pipe_gen1_2_current_coeff[9], w_hssi_pipe_gen1_2_current_coeff[8], w_hssi_pipe_gen1_2_current_coeff[7], w_hssi_pipe_gen1_2_current_coeff[6], w_hssi_pipe_gen1_2_current_coeff[5], w_hssi_pipe_gen1_2_current_coeff[4], w_hssi_pipe_gen1_2_current_coeff[3], w_hssi_pipe_gen1_2_current_coeff[2], w_hssi_pipe_gen1_2_current_coeff[1], w_hssi_pipe_gen1_2_current_coeff[0]}),
				.int_pmaif_8g_eios_det({w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1], w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0]}),
				.int_pmaif_8g_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
				.int_pmaif_8g_rev_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.int_pmaif_8g_tx_clk_out_gen3(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
				.int_pmaif_8g_txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				.int_pmaif_g3_eios_det({w_hssi_gen3_rx_pcs_ei_det_int, w_hssi_gen3_rx_pcs_ei_partial_det_int, w_hssi_gen3_rx_pcs_i_det_int}),
				.int_pmaif_g3_pma_current_coeff({w_hssi_pipe_gen3_pma_current_coeff[17], w_hssi_pipe_gen3_pma_current_coeff[16], w_hssi_pipe_gen3_pma_current_coeff[15], w_hssi_pipe_gen3_pma_current_coeff[14], w_hssi_pipe_gen3_pma_current_coeff[13], w_hssi_pipe_gen3_pma_current_coeff[12], w_hssi_pipe_gen3_pma_current_coeff[11], w_hssi_pipe_gen3_pma_current_coeff[10], w_hssi_pipe_gen3_pma_current_coeff[9], w_hssi_pipe_gen3_pma_current_coeff[8], w_hssi_pipe_gen3_pma_current_coeff[7], w_hssi_pipe_gen3_pma_current_coeff[6], w_hssi_pipe_gen3_pma_current_coeff[5], w_hssi_pipe_gen3_pma_current_coeff[4], w_hssi_pipe_gen3_pma_current_coeff[3], w_hssi_pipe_gen3_pma_current_coeff[2], w_hssi_pipe_gen3_pma_current_coeff[1], w_hssi_pipe_gen3_pma_current_coeff[0]}),
				.int_pmaif_g3_pma_current_rxpreset({w_hssi_pipe_gen3_pma_current_rxpreset[2], w_hssi_pipe_gen3_pma_current_rxpreset[1], w_hssi_pipe_gen3_pma_current_rxpreset[0]}),
				.int_pmaif_g3_pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.int_pmaif_g3_rev_lpbk(w_hssi_pipe_gen3_rev_lpbk_int),
				.int_pmaif_pldif_8g_tx_pld_rstn(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pmaif_pldif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pmaif_pldif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pmaif_pldif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pmaif_pldif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pmaif_pldif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pmaif_pldif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pmaif_pldif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pmaif_pldif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pmaif_pldif_pcie_switch({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0]}),
				.int_pmaif_pldif_pma_reserved_out({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0]}),
				.int_pmaif_pldif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pmaif_pldif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pmaif_pldif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pmaif_pldif_rate({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0]}),
				.int_pmaif_pldif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pmaif_pldif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pmaif_pldif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.int_pmaif_pldif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pmaif_pldif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pmaif_pldif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pmaif_pldif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pmaif_pldif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pmaif_pldif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.int_tx_dft_obsrv_clk({w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1], w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0]}),
				.iocsr_clk(in_iocsr_clk),
				.iocsr_config({in_iocsr_config[5], in_iocsr_config[4], in_iocsr_config[3], in_iocsr_config[2], in_iocsr_config[1], in_iocsr_config[0]}),
				.iocsr_rdy(in_iocsr_rdy),
				.iocsr_rdy_dly(in_iocsr_rdy_dly),
				.pma_adapt_done(in_pma_adapt_done),
				.pma_clklow(in_pma_clklow),
				.pma_fref(in_pma_fref),
				.pma_hclk(in_pma_hclk),
				.pma_pcie_sw_done({in_pma_pcie_sw_done[1], in_pma_pcie_sw_done[0]}),
				.pma_pfdmode_lock(in_pma_pfdmode_lock),
				.pma_reserved_in({in_pma_reserved_in[4], in_pma_reserved_in[3], in_pma_reserved_in[2], in_pma_reserved_in[1], in_pma_reserved_in[0]}),
				.pma_signal_det(in_pma_signal_det),
				.pma_testbus({in_pma_testbus[7], in_pma_testbus[6], in_pma_testbus[5], in_pma_testbus[4], in_pma_testbus[3], in_pma_testbus[2], in_pma_testbus[1], in_pma_testbus[0]}),
				.pmaif_bundling_in_down({in_bond_pmaif_in_bot[11], in_bond_pmaif_in_bot[10], in_bond_pmaif_in_bot[9], in_bond_pmaif_in_bot[8], in_bond_pmaif_in_bot[7], in_bond_pmaif_in_bot[6], in_bond_pmaif_in_bot[5], in_bond_pmaif_in_bot[4], in_bond_pmaif_in_bot[3], in_bond_pmaif_in_bot[2], in_bond_pmaif_in_bot[1], in_bond_pmaif_in_bot[0]}),
				.pmaif_bundling_in_up({in_bond_pmaif_in_top[11], in_bond_pmaif_in_top[10], in_bond_pmaif_in_top[9], in_bond_pmaif_in_top[8], in_bond_pmaif_in_top[7], in_bond_pmaif_in_top[6], in_bond_pmaif_in_top[5], in_bond_pmaif_in_top[4], in_bond_pmaif_in_top[3], in_bond_pmaif_in_top[2], in_bond_pmaif_in_top[1], in_bond_pmaif_in_top[0]}),
				.rx_pmaif_test_out({w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1], w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0]}),
				.rx_prbs_ver_test({w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1], w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0]}),
				.tx_prbs_gen_test({w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1], w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0]}),
				.uhsif_test_out_1({w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0]}),
				.uhsif_test_out_2({w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0]}),
				.uhsif_test_out_3({w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1], w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0]}),
				
				// UNUSED
				.int_pmaif_avmm_iocsr_clk(),
				.int_pmaif_avmm_iocsr_config(),
				.int_pmaif_avmm_iocsr_rdy(),
				.int_pmaif_avmm_iocsr_rdy_dly(),
				.int_pmaif_pldif_interface_select(),
				.pma_tx_pma_syncp(),
				.sta_pma_hclk_by2()
			);
		end // if generate
		else begin
				assign w_hssi_common_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8:0] = 9'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk = 1'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19:0] = 20'b0;
				assign w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7:0] = 8'b0;
				assign w_hssi_common_pcs_pma_interface_pma_adapt_start = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_csr_test_dis = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pcs_pma_interface_pma_early_eios = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_interface_select[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltd_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ltr = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nfrzdrv = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_nrpi_freeze = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pcs_pma_interface_pma_ppm_lock = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pma_tx_bitslip = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx = in_pld_pma_txdetectrx;		// Override default tieoff
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11:0] = 12'b0;
				assign w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11:0] = 12'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_common_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_common_pld_pcs_interface
			twentynm_hssi_common_pld_pcs_interface #(
				.dft_clk_out_en(hssi_common_pld_pcs_interface_dft_clk_out_en),
				.dft_clk_out_sel(hssi_common_pld_pcs_interface_dft_clk_out_sel),
				.hrdrstctrl_en(hssi_common_pld_pcs_interface_hrdrstctrl_en),
				.pcs_testbus_block_sel(hssi_common_pld_pcs_interface_pcs_testbus_block_sel),
				.reconfig_settings(hssi_common_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm4es" )       //PARAM_HIDE
			) inst_twentynm_hssi_common_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_common_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_common_pld_pcs_interface_blockselect),
				.hip_cmn_clk(w_hssi_common_pld_pcs_interface_hip_cmn_clk),
				.hip_cmn_ctrl(w_hssi_common_pld_pcs_interface_hip_cmn_ctrl),
				.hip_iocsr_rdy(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy),
				.hip_iocsr_rdy_dly(w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly),
				.hip_nfrzdrv(w_hssi_common_pld_pcs_interface_hip_nfrzdrv),
				.hip_npor(w_hssi_common_pld_pcs_interface_hip_npor),
				.hip_usermode(w_hssi_common_pld_pcs_interface_hip_usermode),
				.int_pldif_10g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
				.int_pldif_10g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
				.int_pldif_8g_eidleinfersel(w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel),
				.int_pldif_8g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
				.int_pldif_8g_refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
				.int_pldif_8g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
				.int_pldif_g3_current_coeff(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff),
				.int_pldif_g3_current_rxpreset(w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset),
				.int_pldif_krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
				.int_pldif_krfec_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.int_pldif_krfec_scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				.int_pldif_mem_atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.int_pldif_mem_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.int_pldif_pmaif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
				.int_pldif_pmaif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
				.int_pldif_pmaif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
				.int_pldif_pmaif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
				.int_pldif_pmaif_eye_monitor(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor),
				.int_pldif_pmaif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
				.int_pldif_pmaif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
				.int_pldif_pmaif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
				.int_pldif_pmaif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
				.int_pldif_pmaif_pcie_switch(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch),
				.int_pldif_pmaif_pma_reserved_out(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out),
				.int_pldif_pmaif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.int_pldif_pmaif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				.int_pldif_pmaif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
				.int_pldif_pmaif_rate(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate),
				.int_pldif_pmaif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.int_pldif_pmaif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
				.int_pldif_pmaif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
				.int_pldif_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.int_pldif_pmaif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
				.int_pldif_pmaif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
				.int_pldif_pmaif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
				.int_pldif_pmaif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
				.int_pldif_pmaif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
				.int_pldif_pmaif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
				.int_pldif_pmaif_uhsif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.pld_pma_adapt_done(w_hssi_common_pld_pcs_interface_pld_pma_adapt_done),
				.pld_pma_clklow(w_hssi_common_pld_pcs_interface_pld_pma_clklow),
				.pld_pma_fref(w_hssi_common_pld_pcs_interface_pld_pma_fref),
				.pld_pma_hclk(w_hssi_common_pld_pcs_interface_pld_pma_hclk),
				.pld_pma_pcie_sw_done(w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done),
				.pld_pma_pfdmode_lock(w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock),
				.pld_pma_reserved_in(w_hssi_common_pld_pcs_interface_pld_pma_reserved_in),
				.pld_pma_rx_detect_valid(w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid),
				.pld_pma_rx_found(w_hssi_common_pld_pcs_interface_pld_pma_rx_found),
				.pld_pma_rxpll_lock(w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock),
				.pld_pma_testbus(w_hssi_common_pld_pcs_interface_pld_pma_testbus),
				.pld_pmaif_mask_tx_pll(w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll),
				.pld_reserved_out(w_hssi_common_pld_pcs_interface_pld_reserved_out),
				.pld_test_data(w_hssi_common_pld_pcs_interface_pld_test_data),
				.pld_uhsif_lock(w_hssi_common_pld_pcs_interface_pld_uhsif_lock),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
				.int_pldif_10g_test_data({w_hssi_10g_tx_pcs_tx_test_data[19], w_hssi_10g_tx_pcs_tx_test_data[18], w_hssi_10g_tx_pcs_tx_test_data[17], w_hssi_10g_tx_pcs_tx_test_data[16], w_hssi_10g_tx_pcs_tx_test_data[15], w_hssi_10g_tx_pcs_tx_test_data[14], w_hssi_10g_tx_pcs_tx_test_data[13], w_hssi_10g_tx_pcs_tx_test_data[12], w_hssi_10g_tx_pcs_tx_test_data[11], w_hssi_10g_tx_pcs_tx_test_data[10], w_hssi_10g_tx_pcs_tx_test_data[9], w_hssi_10g_tx_pcs_tx_test_data[8], w_hssi_10g_tx_pcs_tx_test_data[7], w_hssi_10g_tx_pcs_tx_test_data[6], w_hssi_10g_tx_pcs_tx_test_data[5], w_hssi_10g_tx_pcs_tx_test_data[4], w_hssi_10g_tx_pcs_tx_test_data[3], w_hssi_10g_tx_pcs_tx_test_data[2], w_hssi_10g_tx_pcs_tx_test_data[1], w_hssi_10g_tx_pcs_tx_test_data[0]}),
				.int_pldif_10g_tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
				.int_pldif_8g_chnl_test_bus_out({w_hssi_8g_rx_pcs_chnl_test_bus_out[19], w_hssi_8g_rx_pcs_chnl_test_bus_out[18], w_hssi_8g_rx_pcs_chnl_test_bus_out[17], w_hssi_8g_rx_pcs_chnl_test_bus_out[16], w_hssi_8g_rx_pcs_chnl_test_bus_out[15], w_hssi_8g_rx_pcs_chnl_test_bus_out[14], w_hssi_8g_rx_pcs_chnl_test_bus_out[13], w_hssi_8g_rx_pcs_chnl_test_bus_out[12], w_hssi_8g_rx_pcs_chnl_test_bus_out[11], w_hssi_8g_rx_pcs_chnl_test_bus_out[10], w_hssi_8g_rx_pcs_chnl_test_bus_out[9], w_hssi_8g_rx_pcs_chnl_test_bus_out[8], w_hssi_8g_rx_pcs_chnl_test_bus_out[7], w_hssi_8g_rx_pcs_chnl_test_bus_out[6], w_hssi_8g_rx_pcs_chnl_test_bus_out[5], w_hssi_8g_rx_pcs_chnl_test_bus_out[4], w_hssi_8g_rx_pcs_chnl_test_bus_out[3], w_hssi_8g_rx_pcs_chnl_test_bus_out[2], w_hssi_8g_rx_pcs_chnl_test_bus_out[1], w_hssi_8g_rx_pcs_chnl_test_bus_out[0]}),
				.int_pldif_8g_rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
				.int_pldif_8g_tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
				.int_pldif_g3_test_out({w_hssi_pipe_gen3_test_out[19], w_hssi_pipe_gen3_test_out[18], w_hssi_pipe_gen3_test_out[17], w_hssi_pipe_gen3_test_out[16], w_hssi_pipe_gen3_test_out[15], w_hssi_pipe_gen3_test_out[14], w_hssi_pipe_gen3_test_out[13], w_hssi_pipe_gen3_test_out[12], w_hssi_pipe_gen3_test_out[11], w_hssi_pipe_gen3_test_out[10], w_hssi_pipe_gen3_test_out[9], w_hssi_pipe_gen3_test_out[8], w_hssi_pipe_gen3_test_out[7], w_hssi_pipe_gen3_test_out[6], w_hssi_pipe_gen3_test_out[5], w_hssi_pipe_gen3_test_out[4], w_hssi_pipe_gen3_test_out[3], w_hssi_pipe_gen3_test_out[2], w_hssi_pipe_gen3_test_out[1], w_hssi_pipe_gen3_test_out[0]}),
				.int_pldif_krfec_test_data({w_hssi_krfec_tx_pcs_tx_test_data[19], w_hssi_krfec_tx_pcs_tx_test_data[18], w_hssi_krfec_tx_pcs_tx_test_data[17], w_hssi_krfec_tx_pcs_tx_test_data[16], w_hssi_krfec_tx_pcs_tx_test_data[15], w_hssi_krfec_tx_pcs_tx_test_data[14], w_hssi_krfec_tx_pcs_tx_test_data[13], w_hssi_krfec_tx_pcs_tx_test_data[12], w_hssi_krfec_tx_pcs_tx_test_data[11], w_hssi_krfec_tx_pcs_tx_test_data[10], w_hssi_krfec_tx_pcs_tx_test_data[9], w_hssi_krfec_tx_pcs_tx_test_data[8], w_hssi_krfec_tx_pcs_tx_test_data[7], w_hssi_krfec_tx_pcs_tx_test_data[6], w_hssi_krfec_tx_pcs_tx_test_data[5], w_hssi_krfec_tx_pcs_tx_test_data[4], w_hssi_krfec_tx_pcs_tx_test_data[3], w_hssi_krfec_tx_pcs_tx_test_data[2], w_hssi_krfec_tx_pcs_tx_test_data[1], w_hssi_krfec_tx_pcs_tx_test_data[0]}),
				.int_pldif_pmaif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
				.int_pldif_pmaif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
				.int_pldif_pmaif_pcie_sw_done({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0]}),
				.int_pldif_pmaif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
				.int_pldif_pmaif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
				.int_pldif_pmaif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
				.int_pldif_pmaif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
				.int_pldif_pmaif_pma_reserved_in({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0]}),
				.int_pldif_pmaif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pldif_pmaif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_test_out({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0]}),
				.int_pldif_pmaif_testbus({w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1], w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0]}),
				.int_pldif_pmaif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.pld_8g_eidleinfersel({in_pld_8g_eidleinfersel[2], in_pld_8g_eidleinfersel[1], in_pld_8g_eidleinfersel[0]}),
				.pld_8g_refclk_dig2(in_pld_8g_refclk_dig2),
				.pld_atpg_los_en_n(in_pld_atpg_los_en_n),
				.pld_g3_current_coeff({in_pld_g3_current_coeff[17], in_pld_g3_current_coeff[16], in_pld_g3_current_coeff[15], in_pld_g3_current_coeff[14], in_pld_g3_current_coeff[13], in_pld_g3_current_coeff[12], in_pld_g3_current_coeff[11], in_pld_g3_current_coeff[10], in_pld_g3_current_coeff[9], in_pld_g3_current_coeff[8], in_pld_g3_current_coeff[7], in_pld_g3_current_coeff[6], in_pld_g3_current_coeff[5], in_pld_g3_current_coeff[4], in_pld_g3_current_coeff[3], in_pld_g3_current_coeff[2], in_pld_g3_current_coeff[1], in_pld_g3_current_coeff[0]}),
				.pld_g3_current_rxpreset({in_pld_g3_current_rxpreset[2], in_pld_g3_current_rxpreset[1], in_pld_g3_current_rxpreset[0]}),
				.pld_ltr(in_pld_ltr),
				.pld_mem_krfec_atpg_rst_n(in_pld_mem_krfec_atpg_rst_n),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pcs_refclk_dig(in_pld_pcs_refclk_dig),
				.pld_pma_adapt_start(in_pld_pma_adapt_start),
				.pld_pma_csr_test_dis(in_pld_pma_csr_test_dis),
				.pld_pma_early_eios(in_pld_pma_early_eios),
				.pld_pma_eye_monitor({in_pld_pma_eye_monitor[5], in_pld_pma_eye_monitor[4], in_pld_pma_eye_monitor[3], in_pld_pma_eye_monitor[2], in_pld_pma_eye_monitor[1], in_pld_pma_eye_monitor[0]}),
				.pld_pma_ltd_b(in_pld_pma_ltd_b),
				.pld_pma_nrpi_freeze(in_pld_pma_nrpi_freeze),
				.pld_pma_pcie_switch({in_pld_pma_pcie_switch[1], in_pld_pma_pcie_switch[0]}),
				.pld_pma_ppm_lock(in_pld_pma_ppm_lock),
				.pld_pma_reserved_out({in_pld_pma_reserved_out[4], in_pld_pma_reserved_out[3], in_pld_pma_reserved_out[2], in_pld_pma_reserved_out[1], in_pld_pma_reserved_out[0]}),
				.pld_pma_rs_lpbk_b(in_pld_pma_rs_lpbk_b),
				.pld_pma_rx_qpi_pullup(in_pld_pma_rx_qpi_pullup),
				.pld_pma_tx_bitslip(in_pld_pma_tx_bitslip),
				.pld_pma_tx_bonding_rstb(in_pld_pma_tx_bonding_rstb),
				.pld_pma_tx_qpi_pulldn(in_pld_pma_tx_qpi_pulldn),
				.pld_pma_tx_qpi_pullup(in_pld_pma_tx_qpi_pullup),
				.pld_pma_txdetectrx(in_pld_pma_txdetectrx),
				.pld_rate({in_pld_rate[1], in_pld_rate[0]}),
				.pld_reserved_in({in_pld_reserved_in[9], in_pld_reserved_in[8], in_pld_reserved_in[7], in_pld_reserved_in[6], in_pld_reserved_in[5], in_pld_reserved_in[4], in_pld_reserved_in[3], in_pld_reserved_in[2], in_pld_reserved_in[1], in_pld_reserved_in[0]}),
				.pld_scan_mode_n(in_pld_scan_mode_n),
				.pld_scan_shift_n(in_pld_scan_shift_n),
				
				// UNUSED
				.int_pldif_8g_ltr(),
				.int_pldif_avmm_pld_avmm1_request(),
				.int_pldif_avmm_pld_avmm2_request(),
				.int_pldif_avmm_refclk_dig_en(),
				.int_pldif_g3_scan_mode_n(),
				.pld_8g_eidleinfersel_fifo(),
				.pld_8g_eidleinfersel_reg(),
				.pld_partial_reconfig_fifo(),
				.pld_partial_reconfig_rx_div_by_2_rxclk_wire(),
				.pld_partial_reconfig_rx_div_by_2_txclk_wire(),
				.pld_partial_reconfig_rxclk_reg(),
				.pld_partial_reconfig_tx_div_by_2_wire(),
				.pld_partial_reconfig_txclk_reg(),
				.pld_rate_reg(),
				.pld_test_data_reg()
			);
		end // if generate
		else begin
				assign w_hssi_common_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_clk[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_npor = 1'b0;
				assign w_hssi_common_pld_pcs_interface_hip_usermode = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2 = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17:0] = 18'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5:0] = 6'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n = 1'b1;		// Override default tieoff
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel = 1'b0;
				assign w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_adapt_done = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_clklow = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_fref = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_hclk = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1:0] = 2'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4:0] = 5'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rx_found = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pma_testbus[7:0] = 8'b0;
				assign w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll = 1'b0;
				assign w_hssi_common_pld_pcs_interface_pld_reserved_out[9:0] = 10'b0;
				assign w_hssi_common_pld_pcs_interface_pld_test_data[19:0] = 20'b0;
				assign w_hssi_common_pld_pcs_interface_pld_uhsif_lock = 1'b0;
				assign w_hssi_common_pld_pcs_interface_scan_mode_n = 1'b1;		// Override default tieoff
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_rx_pcs
			twentynm_hssi_fifo_rx_pcs #(
				.double_read_mode(hssi_fifo_rx_pcs_double_read_mode),
				.prot_mode(hssi_fifo_rx_pcs_prot_mode),
				.silicon_rev( "20nm4es" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_rx_pcs_blockselect),
				.data_out2_10g(w_hssi_fifo_rx_pcs_data_out2_10g),
				.data_out2_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp),
				.data_out_10g(w_hssi_fifo_rx_pcs_data_out_10g),
				.data_out_8g_clock_comp(w_hssi_fifo_rx_pcs_data_out_8g_clock_comp),
				.data_out_8g_phase_comp(w_hssi_fifo_rx_pcs_data_out_8g_phase_comp),
				.data_out_gen3(w_hssi_fifo_rx_pcs_data_out_gen3),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_data[73], w_hssi_10g_rx_pcs_rx_fifo_wr_data[72], w_hssi_10g_rx_pcs_rx_fifo_wr_data[71], w_hssi_10g_rx_pcs_rx_fifo_wr_data[70], w_hssi_10g_rx_pcs_rx_fifo_wr_data[69], w_hssi_10g_rx_pcs_rx_fifo_wr_data[68], w_hssi_10g_rx_pcs_rx_fifo_wr_data[67], w_hssi_10g_rx_pcs_rx_fifo_wr_data[66], w_hssi_10g_rx_pcs_rx_fifo_wr_data[65], w_hssi_10g_rx_pcs_rx_fifo_wr_data[64], w_hssi_10g_rx_pcs_rx_fifo_wr_data[63], w_hssi_10g_rx_pcs_rx_fifo_wr_data[62], w_hssi_10g_rx_pcs_rx_fifo_wr_data[61], w_hssi_10g_rx_pcs_rx_fifo_wr_data[60], w_hssi_10g_rx_pcs_rx_fifo_wr_data[59], w_hssi_10g_rx_pcs_rx_fifo_wr_data[58], w_hssi_10g_rx_pcs_rx_fifo_wr_data[57], w_hssi_10g_rx_pcs_rx_fifo_wr_data[56], w_hssi_10g_rx_pcs_rx_fifo_wr_data[55], w_hssi_10g_rx_pcs_rx_fifo_wr_data[54], w_hssi_10g_rx_pcs_rx_fifo_wr_data[53], w_hssi_10g_rx_pcs_rx_fifo_wr_data[52], w_hssi_10g_rx_pcs_rx_fifo_wr_data[51], w_hssi_10g_rx_pcs_rx_fifo_wr_data[50], w_hssi_10g_rx_pcs_rx_fifo_wr_data[49], w_hssi_10g_rx_pcs_rx_fifo_wr_data[48], w_hssi_10g_rx_pcs_rx_fifo_wr_data[47], w_hssi_10g_rx_pcs_rx_fifo_wr_data[46], w_hssi_10g_rx_pcs_rx_fifo_wr_data[45], w_hssi_10g_rx_pcs_rx_fifo_wr_data[44], w_hssi_10g_rx_pcs_rx_fifo_wr_data[43], w_hssi_10g_rx_pcs_rx_fifo_wr_data[42], w_hssi_10g_rx_pcs_rx_fifo_wr_data[41], w_hssi_10g_rx_pcs_rx_fifo_wr_data[40], w_hssi_10g_rx_pcs_rx_fifo_wr_data[39], w_hssi_10g_rx_pcs_rx_fifo_wr_data[38], w_hssi_10g_rx_pcs_rx_fifo_wr_data[37], w_hssi_10g_rx_pcs_rx_fifo_wr_data[36], w_hssi_10g_rx_pcs_rx_fifo_wr_data[35], w_hssi_10g_rx_pcs_rx_fifo_wr_data[34], w_hssi_10g_rx_pcs_rx_fifo_wr_data[33], w_hssi_10g_rx_pcs_rx_fifo_wr_data[32], w_hssi_10g_rx_pcs_rx_fifo_wr_data[31], w_hssi_10g_rx_pcs_rx_fifo_wr_data[30], w_hssi_10g_rx_pcs_rx_fifo_wr_data[29], w_hssi_10g_rx_pcs_rx_fifo_wr_data[28], w_hssi_10g_rx_pcs_rx_fifo_wr_data[27], w_hssi_10g_rx_pcs_rx_fifo_wr_data[26], w_hssi_10g_rx_pcs_rx_fifo_wr_data[25], w_hssi_10g_rx_pcs_rx_fifo_wr_data[24], w_hssi_10g_rx_pcs_rx_fifo_wr_data[23], w_hssi_10g_rx_pcs_rx_fifo_wr_data[22], w_hssi_10g_rx_pcs_rx_fifo_wr_data[21], w_hssi_10g_rx_pcs_rx_fifo_wr_data[20], w_hssi_10g_rx_pcs_rx_fifo_wr_data[19], w_hssi_10g_rx_pcs_rx_fifo_wr_data[18], w_hssi_10g_rx_pcs_rx_fifo_wr_data[17], w_hssi_10g_rx_pcs_rx_fifo_wr_data[16], w_hssi_10g_rx_pcs_rx_fifo_wr_data[15], w_hssi_10g_rx_pcs_rx_fifo_wr_data[14], w_hssi_10g_rx_pcs_rx_fifo_wr_data[13], w_hssi_10g_rx_pcs_rx_fifo_wr_data[12], w_hssi_10g_rx_pcs_rx_fifo_wr_data[11], w_hssi_10g_rx_pcs_rx_fifo_wr_data[10], w_hssi_10g_rx_pcs_rx_fifo_wr_data[9], w_hssi_10g_rx_pcs_rx_fifo_wr_data[8], w_hssi_10g_rx_pcs_rx_fifo_wr_data[7], w_hssi_10g_rx_pcs_rx_fifo_wr_data[6], w_hssi_10g_rx_pcs_rx_fifo_wr_data[5], w_hssi_10g_rx_pcs_rx_fifo_wr_data[4], w_hssi_10g_rx_pcs_rx_fifo_wr_data[3], w_hssi_10g_rx_pcs_rx_fifo_wr_data[2], w_hssi_10g_rx_pcs_rx_fifo_wr_data[1], w_hssi_10g_rx_pcs_rx_fifo_wr_data[0]}),
				.data_in_8g_clock_comp({w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0]}),
				.data_in_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr2_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0]}),
				.rd_ptr2_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0]}),
				.rd_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1], w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0]}),
				.rd_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
				.wr_clk_8g_clock_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
				.wr_clk_8g_clock_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
				.wr_clk_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.wr_en_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
				.wr_en_8g_clock_comp(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
				.wr_en_8g_phase_comp(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
				.wr_en_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.wr_ptr_10g({w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1], w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_clock_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1], w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0]}),
				.wr_ptr_gen3({w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1], w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0]}),
				.wr_rst_n_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
				.wr_rst_n_8g_clock_comp(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
				.wr_rst_n_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_rx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_10g[73:0] = 74'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31:0] = 32'b0;
				assign w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79:0] = 80'b0;
				assign w_hssi_fifo_rx_pcs_data_out_gen3[39:0] = 40'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_fifo_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_fifo_tx_pcs
			twentynm_hssi_fifo_tx_pcs #(
				.double_write_mode(hssi_fifo_tx_pcs_double_write_mode),
				.prot_mode(hssi_fifo_tx_pcs_prot_mode),
				.silicon_rev( "20nm4es" )       //PARAM_HIDE
			) inst_twentynm_hssi_fifo_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_fifo_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_fifo_tx_pcs_blockselect),
				.data_out_10g(w_hssi_fifo_tx_pcs_data_out_10g),
				.data_out_8g_phase_comp(w_hssi_fifo_tx_pcs_data_out_8g_phase_comp),
				// INPUTS
				.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in2_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0]}),
				.data_in_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_data[72], w_hssi_10g_tx_pcs_tx_fifo_wr_data[71], w_hssi_10g_tx_pcs_tx_fifo_wr_data[70], w_hssi_10g_tx_pcs_tx_fifo_wr_data[69], w_hssi_10g_tx_pcs_tx_fifo_wr_data[68], w_hssi_10g_tx_pcs_tx_fifo_wr_data[67], w_hssi_10g_tx_pcs_tx_fifo_wr_data[66], w_hssi_10g_tx_pcs_tx_fifo_wr_data[65], w_hssi_10g_tx_pcs_tx_fifo_wr_data[64], w_hssi_10g_tx_pcs_tx_fifo_wr_data[63], w_hssi_10g_tx_pcs_tx_fifo_wr_data[62], w_hssi_10g_tx_pcs_tx_fifo_wr_data[61], w_hssi_10g_tx_pcs_tx_fifo_wr_data[60], w_hssi_10g_tx_pcs_tx_fifo_wr_data[59], w_hssi_10g_tx_pcs_tx_fifo_wr_data[58], w_hssi_10g_tx_pcs_tx_fifo_wr_data[57], w_hssi_10g_tx_pcs_tx_fifo_wr_data[56], w_hssi_10g_tx_pcs_tx_fifo_wr_data[55], w_hssi_10g_tx_pcs_tx_fifo_wr_data[54], w_hssi_10g_tx_pcs_tx_fifo_wr_data[53], w_hssi_10g_tx_pcs_tx_fifo_wr_data[52], w_hssi_10g_tx_pcs_tx_fifo_wr_data[51], w_hssi_10g_tx_pcs_tx_fifo_wr_data[50], w_hssi_10g_tx_pcs_tx_fifo_wr_data[49], w_hssi_10g_tx_pcs_tx_fifo_wr_data[48], w_hssi_10g_tx_pcs_tx_fifo_wr_data[47], w_hssi_10g_tx_pcs_tx_fifo_wr_data[46], w_hssi_10g_tx_pcs_tx_fifo_wr_data[45], w_hssi_10g_tx_pcs_tx_fifo_wr_data[44], w_hssi_10g_tx_pcs_tx_fifo_wr_data[43], w_hssi_10g_tx_pcs_tx_fifo_wr_data[42], w_hssi_10g_tx_pcs_tx_fifo_wr_data[41], w_hssi_10g_tx_pcs_tx_fifo_wr_data[40], w_hssi_10g_tx_pcs_tx_fifo_wr_data[39], w_hssi_10g_tx_pcs_tx_fifo_wr_data[38], w_hssi_10g_tx_pcs_tx_fifo_wr_data[37], w_hssi_10g_tx_pcs_tx_fifo_wr_data[36], w_hssi_10g_tx_pcs_tx_fifo_wr_data[35], w_hssi_10g_tx_pcs_tx_fifo_wr_data[34], w_hssi_10g_tx_pcs_tx_fifo_wr_data[33], w_hssi_10g_tx_pcs_tx_fifo_wr_data[32], w_hssi_10g_tx_pcs_tx_fifo_wr_data[31], w_hssi_10g_tx_pcs_tx_fifo_wr_data[30], w_hssi_10g_tx_pcs_tx_fifo_wr_data[29], w_hssi_10g_tx_pcs_tx_fifo_wr_data[28], w_hssi_10g_tx_pcs_tx_fifo_wr_data[27], w_hssi_10g_tx_pcs_tx_fifo_wr_data[26], w_hssi_10g_tx_pcs_tx_fifo_wr_data[25], w_hssi_10g_tx_pcs_tx_fifo_wr_data[24], w_hssi_10g_tx_pcs_tx_fifo_wr_data[23], w_hssi_10g_tx_pcs_tx_fifo_wr_data[22], w_hssi_10g_tx_pcs_tx_fifo_wr_data[21], w_hssi_10g_tx_pcs_tx_fifo_wr_data[20], w_hssi_10g_tx_pcs_tx_fifo_wr_data[19], w_hssi_10g_tx_pcs_tx_fifo_wr_data[18], w_hssi_10g_tx_pcs_tx_fifo_wr_data[17], w_hssi_10g_tx_pcs_tx_fifo_wr_data[16], w_hssi_10g_tx_pcs_tx_fifo_wr_data[15], w_hssi_10g_tx_pcs_tx_fifo_wr_data[14], w_hssi_10g_tx_pcs_tx_fifo_wr_data[13], w_hssi_10g_tx_pcs_tx_fifo_wr_data[12], w_hssi_10g_tx_pcs_tx_fifo_wr_data[11], w_hssi_10g_tx_pcs_tx_fifo_wr_data[10], w_hssi_10g_tx_pcs_tx_fifo_wr_data[9], w_hssi_10g_tx_pcs_tx_fifo_wr_data[8], w_hssi_10g_tx_pcs_tx_fifo_wr_data[7], w_hssi_10g_tx_pcs_tx_fifo_wr_data[6], w_hssi_10g_tx_pcs_tx_fifo_wr_data[5], w_hssi_10g_tx_pcs_tx_fifo_wr_data[4], w_hssi_10g_tx_pcs_tx_fifo_wr_data[3], w_hssi_10g_tx_pcs_tx_fifo_wr_data[2], w_hssi_10g_tx_pcs_tx_fifo_wr_data[1], w_hssi_10g_tx_pcs_tx_fifo_wr_data[0]}),
				.data_in_8g_phase_comp({w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0]}),
				.hard_reset_n(1'b0),
				.rd_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0]}),
				.rd_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0]}),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
				.wr_clk_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
				.wr_clk_8g_phase_comp_dw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
				.wr_clk_8g_phase_comp_sw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
				.wr_en_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
				.wr_en_8g_phase_comp(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
				.wr_ptr_10g({w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1], w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0]}),
				.wr_ptr_8g_phase_comp({w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1], w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0]}),
				.wr_rst_n_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
				.wr_rst_n_8g_phase_comp(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo)
			);
		end // if generate
		else begin
				assign w_hssi_fifo_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_fifo_tx_pcs_blockselect = 1'b0;
				assign w_hssi_fifo_tx_pcs_data_out_10g[72:0] = 73'b0;
				assign w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63:0] = 64'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_rx_pcs
			twentynm_hssi_gen3_rx_pcs #(
				.block_sync(hssi_gen3_rx_pcs_block_sync),
				.block_sync_sm(hssi_gen3_rx_pcs_block_sync_sm),
				.cdr_ctrl_force_unalgn(hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn),
				.lpbk_force(hssi_gen3_rx_pcs_lpbk_force),
				.mode(hssi_gen3_rx_pcs_mode),
				.rate_match_fifo(hssi_gen3_rx_pcs_rate_match_fifo),
				.rate_match_fifo_latency(hssi_gen3_rx_pcs_rate_match_fifo_latency),
				.reconfig_settings(hssi_gen3_rx_pcs_reconfig_settings),
				.reverse_lpbk(hssi_gen3_rx_pcs_reverse_lpbk),
				.rx_b4gb_par_lpbk(hssi_gen3_rx_pcs_rx_b4gb_par_lpbk),
				.rx_force_balign(hssi_gen3_rx_pcs_rx_force_balign),
				.rx_ins_del_one_skip(hssi_gen3_rx_pcs_rx_ins_del_one_skip),
				.rx_num_fixed_pat(hssi_gen3_rx_pcs_rx_num_fixed_pat),
				.rx_test_out_sel(hssi_gen3_rx_pcs_rx_test_out_sel),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_rx_pcs_sup_mode)
			) inst_twentynm_hssi_gen3_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_rx_pcs_avmmreaddata),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.blk_start(w_hssi_gen3_rx_pcs_blk_start),
				.blockselect(w_hssi_gen3_rx_pcs_blockselect),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.data_out(w_hssi_gen3_rx_pcs_data_out),
				.data_valid(w_hssi_gen3_rx_pcs_data_valid),
				.ei_det_int(w_hssi_gen3_rx_pcs_ei_det_int),
				.ei_partial_det_int(w_hssi_gen3_rx_pcs_ei_partial_det_int),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.i_det_int(w_hssi_gen3_rx_pcs_i_det_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data(w_hssi_gen3_rx_pcs_lpbk_data),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.mem_rx_fifo_rd_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr),
				.mem_rx_fifo_wr_clk(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
				.mem_rx_fifo_wr_data(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data),
				.mem_rx_fifo_wr_en(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
				.mem_rx_fifo_wr_ptr(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr),
				.mem_rx_fifo_wr_rst_n(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_test_out(w_hssi_gen3_rx_pcs_rx_test_out),
				.sync_hdr(w_hssi_gen3_rx_pcs_sync_hdr),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1], w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0]}),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.mem_rx_fifo_rd_data({w_hssi_fifo_rx_pcs_data_out_gen3[39], w_hssi_fifo_rx_pcs_data_out_gen3[38], w_hssi_fifo_rx_pcs_data_out_gen3[37], w_hssi_fifo_rx_pcs_data_out_gen3[36], w_hssi_fifo_rx_pcs_data_out_gen3[35], w_hssi_fifo_rx_pcs_data_out_gen3[34], w_hssi_fifo_rx_pcs_data_out_gen3[33], w_hssi_fifo_rx_pcs_data_out_gen3[32], w_hssi_fifo_rx_pcs_data_out_gen3[31], w_hssi_fifo_rx_pcs_data_out_gen3[30], w_hssi_fifo_rx_pcs_data_out_gen3[29], w_hssi_fifo_rx_pcs_data_out_gen3[28], w_hssi_fifo_rx_pcs_data_out_gen3[27], w_hssi_fifo_rx_pcs_data_out_gen3[26], w_hssi_fifo_rx_pcs_data_out_gen3[25], w_hssi_fifo_rx_pcs_data_out_gen3[24], w_hssi_fifo_rx_pcs_data_out_gen3[23], w_hssi_fifo_rx_pcs_data_out_gen3[22], w_hssi_fifo_rx_pcs_data_out_gen3[21], w_hssi_fifo_rx_pcs_data_out_gen3[20], w_hssi_fifo_rx_pcs_data_out_gen3[19], w_hssi_fifo_rx_pcs_data_out_gen3[18], w_hssi_fifo_rx_pcs_data_out_gen3[17], w_hssi_fifo_rx_pcs_data_out_gen3[16], w_hssi_fifo_rx_pcs_data_out_gen3[15], w_hssi_fifo_rx_pcs_data_out_gen3[14], w_hssi_fifo_rx_pcs_data_out_gen3[13], w_hssi_fifo_rx_pcs_data_out_gen3[12], w_hssi_fifo_rx_pcs_data_out_gen3[11], w_hssi_fifo_rx_pcs_data_out_gen3[10], w_hssi_fifo_rx_pcs_data_out_gen3[9], w_hssi_fifo_rx_pcs_data_out_gen3[8], w_hssi_fifo_rx_pcs_data_out_gen3[7], w_hssi_fifo_rx_pcs_data_out_gen3[6], w_hssi_fifo_rx_pcs_data_out_gen3[5], w_hssi_fifo_rx_pcs_data_out_gen3[4], w_hssi_fifo_rx_pcs_data_out_gen3[3], w_hssi_fifo_rx_pcs_data_out_gen3[2], w_hssi_fifo_rx_pcs_data_out_gen3[1], w_hssi_fifo_rx_pcs_data_out_gen3[0]}),
				.par_lpbk_b4gb_in({w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1], w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0]}),
				.par_lpbk_in({w_hssi_gen3_tx_pcs_par_lpbk_out[31], w_hssi_gen3_tx_pcs_par_lpbk_out[30], w_hssi_gen3_tx_pcs_par_lpbk_out[29], w_hssi_gen3_tx_pcs_par_lpbk_out[28], w_hssi_gen3_tx_pcs_par_lpbk_out[27], w_hssi_gen3_tx_pcs_par_lpbk_out[26], w_hssi_gen3_tx_pcs_par_lpbk_out[25], w_hssi_gen3_tx_pcs_par_lpbk_out[24], w_hssi_gen3_tx_pcs_par_lpbk_out[23], w_hssi_gen3_tx_pcs_par_lpbk_out[22], w_hssi_gen3_tx_pcs_par_lpbk_out[21], w_hssi_gen3_tx_pcs_par_lpbk_out[20], w_hssi_gen3_tx_pcs_par_lpbk_out[19], w_hssi_gen3_tx_pcs_par_lpbk_out[18], w_hssi_gen3_tx_pcs_par_lpbk_out[17], w_hssi_gen3_tx_pcs_par_lpbk_out[16], w_hssi_gen3_tx_pcs_par_lpbk_out[15], w_hssi_gen3_tx_pcs_par_lpbk_out[14], w_hssi_gen3_tx_pcs_par_lpbk_out[13], w_hssi_gen3_tx_pcs_par_lpbk_out[12], w_hssi_gen3_tx_pcs_par_lpbk_out[11], w_hssi_gen3_tx_pcs_par_lpbk_out[10], w_hssi_gen3_tx_pcs_par_lpbk_out[9], w_hssi_gen3_tx_pcs_par_lpbk_out[8], w_hssi_gen3_tx_pcs_par_lpbk_out[7], w_hssi_gen3_tx_pcs_par_lpbk_out[6], w_hssi_gen3_tx_pcs_par_lpbk_out[5], w_hssi_gen3_tx_pcs_par_lpbk_out[4], w_hssi_gen3_tx_pcs_par_lpbk_out[3], w_hssi_gen3_tx_pcs_par_lpbk_out[2], w_hssi_gen3_tx_pcs_par_lpbk_out[1], w_hssi_gen3_tx_pcs_par_lpbk_out[0]}),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.rcvd_clk(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
				.rx_pma_clk(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
				.rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
				.rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
				.rxpolarity(w_hssi_pipe_gen3_rxpolarity_int),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.sync_sm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.txdatak_in({w_hssi_pipe_gen3_txdatak_int[3], w_hssi_pipe_gen3_txdatak_int[2], w_hssi_pipe_gen3_txdatak_int[1], w_hssi_pipe_gen3_txdatak_int[0]}),
				
				// UNUSED
				.blk_lockd_int(),
				.skp_det_int()
			);
		end // if generate
		else begin
				assign w_hssi_gen3_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_rx_pcs_blk_algnd_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_delete_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_insert_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_overfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_clkcomp_undfl_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_rx_pcs_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_ei_partial_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_err_decode_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_i_det_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_blk_start = 1'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data[33:0] = 34'b0;
				assign w_hssi_gen3_rx_pcs_lpbk_data_valid = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39:0] = 40'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en = 1'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15:0] = 16'b0;
				assign w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int = 1'b0;
				assign w_hssi_gen3_rx_pcs_rx_test_out[19:0] = 20'b0;
				assign w_hssi_gen3_rx_pcs_sync_hdr[1:0] = 2'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_gen3_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_gen3_tx_pcs
			twentynm_hssi_gen3_tx_pcs #(
				.mode(hssi_gen3_tx_pcs_mode),
				.reverse_lpbk(hssi_gen3_tx_pcs_reverse_lpbk),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sup_mode(hssi_gen3_tx_pcs_sup_mode),
				.tx_bitslip(hssi_gen3_tx_pcs_tx_bitslip),
				.tx_gbox_byp(hssi_gen3_tx_pcs_tx_gbox_byp)
			) inst_twentynm_hssi_gen3_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_gen3_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_gen3_tx_pcs_blockselect),
				.data_out(w_hssi_gen3_tx_pcs_data_out),
				.par_lpbk_b4gb_out(w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out),
				.par_lpbk_out(w_hssi_gen3_tx_pcs_par_lpbk_out),
				.tx_test_out(w_hssi_gen3_tx_pcs_tx_test_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_start_in(w_hssi_pipe_gen3_tx_blk_start_int),
				.data_in({w_hssi_pipe_gen3_txdata_int[31], w_hssi_pipe_gen3_txdata_int[30], w_hssi_pipe_gen3_txdata_int[29], w_hssi_pipe_gen3_txdata_int[28], w_hssi_pipe_gen3_txdata_int[27], w_hssi_pipe_gen3_txdata_int[26], w_hssi_pipe_gen3_txdata_int[25], w_hssi_pipe_gen3_txdata_int[24], w_hssi_pipe_gen3_txdata_int[23], w_hssi_pipe_gen3_txdata_int[22], w_hssi_pipe_gen3_txdata_int[21], w_hssi_pipe_gen3_txdata_int[20], w_hssi_pipe_gen3_txdata_int[19], w_hssi_pipe_gen3_txdata_int[18], w_hssi_pipe_gen3_txdata_int[17], w_hssi_pipe_gen3_txdata_int[16], w_hssi_pipe_gen3_txdata_int[15], w_hssi_pipe_gen3_txdata_int[14], w_hssi_pipe_gen3_txdata_int[13], w_hssi_pipe_gen3_txdata_int[12], w_hssi_pipe_gen3_txdata_int[11], w_hssi_pipe_gen3_txdata_int[10], w_hssi_pipe_gen3_txdata_int[9], w_hssi_pipe_gen3_txdata_int[8], w_hssi_pipe_gen3_txdata_int[7], w_hssi_pipe_gen3_txdata_int[6], w_hssi_pipe_gen3_txdata_int[5], w_hssi_pipe_gen3_txdata_int[4], w_hssi_pipe_gen3_txdata_int[3], w_hssi_pipe_gen3_txdata_int[2], w_hssi_pipe_gen3_txdata_int[1], w_hssi_pipe_gen3_txdata_int[0]}),
				.data_valid(w_hssi_pipe_gen3_txdataskip_int),
				.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
				.lpbk_data_in({w_hssi_gen3_rx_pcs_lpbk_data[33], w_hssi_gen3_rx_pcs_lpbk_data[32], w_hssi_gen3_rx_pcs_lpbk_data[31], w_hssi_gen3_rx_pcs_lpbk_data[30], w_hssi_gen3_rx_pcs_lpbk_data[29], w_hssi_gen3_rx_pcs_lpbk_data[28], w_hssi_gen3_rx_pcs_lpbk_data[27], w_hssi_gen3_rx_pcs_lpbk_data[26], w_hssi_gen3_rx_pcs_lpbk_data[25], w_hssi_gen3_rx_pcs_lpbk_data[24], w_hssi_gen3_rx_pcs_lpbk_data[23], w_hssi_gen3_rx_pcs_lpbk_data[22], w_hssi_gen3_rx_pcs_lpbk_data[21], w_hssi_gen3_rx_pcs_lpbk_data[20], w_hssi_gen3_rx_pcs_lpbk_data[19], w_hssi_gen3_rx_pcs_lpbk_data[18], w_hssi_gen3_rx_pcs_lpbk_data[17], w_hssi_gen3_rx_pcs_lpbk_data[16], w_hssi_gen3_rx_pcs_lpbk_data[15], w_hssi_gen3_rx_pcs_lpbk_data[14], w_hssi_gen3_rx_pcs_lpbk_data[13], w_hssi_gen3_rx_pcs_lpbk_data[12], w_hssi_gen3_rx_pcs_lpbk_data[11], w_hssi_gen3_rx_pcs_lpbk_data[10], w_hssi_gen3_rx_pcs_lpbk_data[9], w_hssi_gen3_rx_pcs_lpbk_data[8], w_hssi_gen3_rx_pcs_lpbk_data[7], w_hssi_gen3_rx_pcs_lpbk_data[6], w_hssi_gen3_rx_pcs_lpbk_data[5], w_hssi_gen3_rx_pcs_lpbk_data[4], w_hssi_gen3_rx_pcs_lpbk_data[3], w_hssi_gen3_rx_pcs_lpbk_data[2], w_hssi_gen3_rx_pcs_lpbk_data[1], w_hssi_gen3_rx_pcs_lpbk_data[0]}),
				.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
				.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
				.sync_in({w_hssi_pipe_gen3_tx_sync_hdr_int[1], w_hssi_pipe_gen3_tx_sync_hdr_int[0]}),
				.tx_pma_clk(w_hssi_8g_tx_pcs_clk_out_gen3),
				.tx_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn)
			);
		end // if generate
		else begin
				assign w_hssi_gen3_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_gen3_tx_pcs_blockselect = 1'b0;
				assign w_hssi_gen3_tx_pcs_data_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35:0] = 36'b0;
				assign w_hssi_gen3_tx_pcs_par_lpbk_out[31:0] = 32'b0;
				assign w_hssi_gen3_tx_pcs_tx_test_out[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_rx_pcs
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_rx_pcs
			twentynm_hssi_krfec_rx_pcs #(
				.blksync_cor_en(hssi_krfec_rx_pcs_blksync_cor_en),
				.bypass_gb(hssi_krfec_rx_pcs_bypass_gb),
				.clr_ctrl(hssi_krfec_rx_pcs_clr_ctrl),
				.ctrl_bit_reverse(hssi_krfec_rx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_rx_pcs_data_bit_reverse),
				.dv_start(hssi_krfec_rx_pcs_dv_start),
				.err_mark_type(hssi_krfec_rx_pcs_err_mark_type),
				.error_marking_en(hssi_krfec_rx_pcs_error_marking_en),
				.low_latency_en(hssi_krfec_rx_pcs_low_latency_en),
				.lpbk_mode(hssi_krfec_rx_pcs_lpbk_mode),
				.parity_invalid_enum(hssi_krfec_rx_pcs_parity_invalid_enum),
				.parity_valid_num(hssi_krfec_rx_pcs_parity_valid_num),
				.pipeln_blksync(hssi_krfec_rx_pcs_pipeln_blksync),
				.pipeln_descrm(hssi_krfec_rx_pcs_pipeln_descrm),
				.pipeln_errcorrect(hssi_krfec_rx_pcs_pipeln_errcorrect),
				.pipeln_errtrap_ind(hssi_krfec_rx_pcs_pipeln_errtrap_ind),
				.pipeln_errtrap_lfsr(hssi_krfec_rx_pcs_pipeln_errtrap_lfsr),
				.pipeln_errtrap_loc(hssi_krfec_rx_pcs_pipeln_errtrap_loc),
				.pipeln_errtrap_pat(hssi_krfec_rx_pcs_pipeln_errtrap_pat),
				.pipeln_gearbox(hssi_krfec_rx_pcs_pipeln_gearbox),
				.pipeln_syndrm(hssi_krfec_rx_pcs_pipeln_syndrm),
				.pipeln_trans_dec(hssi_krfec_rx_pcs_pipeln_trans_dec),
				.prot_mode(hssi_krfec_rx_pcs_prot_mode),
				.receive_order(hssi_krfec_rx_pcs_receive_order),
				.reconfig_settings(hssi_krfec_rx_pcs_reconfig_settings),
				.rx_testbus_sel(hssi_krfec_rx_pcs_rx_testbus_sel),
				.signal_ok_en(hssi_krfec_rx_pcs_signal_ok_en),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_rx_pcs_sup_mode)
			) inst_twentynm_hssi_krfec_rx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_rx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_rx_pcs_blockselect),
				.rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.rx_control_out(w_hssi_krfec_rx_pcs_rx_control_out),
				.rx_data_out(w_hssi_krfec_rx_pcs_rx_data_out),
				.rx_data_status(w_hssi_krfec_rx_pcs_rx_data_status),
				.rx_data_valid_out(w_hssi_krfec_rx_pcs_rx_data_valid_out),
				.rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.rx_signal_ok_out(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.rx_data_in({w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0]}),
				.rx_krfec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
				.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
				.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
				.rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
				.scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
				
				// UNUSED
				.pld_10g_krfec_rx_blk_lock_krfec_reg(),
				.pld_10g_krfec_rx_blk_lock_krfec_txclk_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_reg(),
				.pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg(),
				.pld_10g_krfec_rx_frame_krfec_reg(),
				.pld_10g_krfec_rx_frame_krfec_txclk_reg(),
				.rx_test_data()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_rx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_rx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_block_lock = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_control_out[9:0] = 10'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_status[1:0] = 2'b0;
				assign w_hssi_krfec_rx_pcs_rx_data_valid_out = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_frame = 1'b0;
				assign w_hssi_krfec_rx_pcs_rx_signal_ok_out = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_krfec_tx_pcs
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_krfec_tx_pcs
			twentynm_hssi_krfec_tx_pcs #(
				.burst_err(hssi_krfec_tx_pcs_burst_err),
				.burst_err_len(hssi_krfec_tx_pcs_burst_err_len),
				.ctrl_bit_reverse(hssi_krfec_tx_pcs_ctrl_bit_reverse),
				.data_bit_reverse(hssi_krfec_tx_pcs_data_bit_reverse),
				.enc_frame_query(hssi_krfec_tx_pcs_enc_frame_query),
				.low_latency_en(hssi_krfec_tx_pcs_low_latency_en),
				.pipeln_encoder(hssi_krfec_tx_pcs_pipeln_encoder),
				.pipeln_scrambler(hssi_krfec_tx_pcs_pipeln_scrambler),
				.prot_mode(hssi_krfec_tx_pcs_prot_mode),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sup_mode(hssi_krfec_tx_pcs_sup_mode),
				.transcode_err(hssi_krfec_tx_pcs_transcode_err),
				.transmit_order(hssi_krfec_tx_pcs_transmit_order),
				.tx_testbus_sel(hssi_krfec_tx_pcs_tx_testbus_sel)
			) inst_twentynm_hssi_krfec_tx_pcs (
				// OUTPUTS
				.avmmreaddata(w_hssi_krfec_tx_pcs_avmmreaddata),
				.blockselect(w_hssi_krfec_tx_pcs_blockselect),
				.tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.tx_data_out(w_hssi_krfec_tx_pcs_tx_data_out),
				.tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.tx_test_data(w_hssi_krfec_tx_pcs_tx_test_data),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.tx_control_in({w_hssi_10g_tx_pcs_tx_control_out_krfec[8], w_hssi_10g_tx_pcs_tx_control_out_krfec[7], w_hssi_10g_tx_pcs_tx_control_out_krfec[6], w_hssi_10g_tx_pcs_tx_control_out_krfec[5], w_hssi_10g_tx_pcs_tx_control_out_krfec[4], w_hssi_10g_tx_pcs_tx_control_out_krfec[3], w_hssi_10g_tx_pcs_tx_control_out_krfec[2], w_hssi_10g_tx_pcs_tx_control_out_krfec[1], w_hssi_10g_tx_pcs_tx_control_out_krfec[0]}),
				.tx_data_in({w_hssi_10g_tx_pcs_tx_data_out_krfec[63], w_hssi_10g_tx_pcs_tx_data_out_krfec[62], w_hssi_10g_tx_pcs_tx_data_out_krfec[61], w_hssi_10g_tx_pcs_tx_data_out_krfec[60], w_hssi_10g_tx_pcs_tx_data_out_krfec[59], w_hssi_10g_tx_pcs_tx_data_out_krfec[58], w_hssi_10g_tx_pcs_tx_data_out_krfec[57], w_hssi_10g_tx_pcs_tx_data_out_krfec[56], w_hssi_10g_tx_pcs_tx_data_out_krfec[55], w_hssi_10g_tx_pcs_tx_data_out_krfec[54], w_hssi_10g_tx_pcs_tx_data_out_krfec[53], w_hssi_10g_tx_pcs_tx_data_out_krfec[52], w_hssi_10g_tx_pcs_tx_data_out_krfec[51], w_hssi_10g_tx_pcs_tx_data_out_krfec[50], w_hssi_10g_tx_pcs_tx_data_out_krfec[49], w_hssi_10g_tx_pcs_tx_data_out_krfec[48], w_hssi_10g_tx_pcs_tx_data_out_krfec[47], w_hssi_10g_tx_pcs_tx_data_out_krfec[46], w_hssi_10g_tx_pcs_tx_data_out_krfec[45], w_hssi_10g_tx_pcs_tx_data_out_krfec[44], w_hssi_10g_tx_pcs_tx_data_out_krfec[43], w_hssi_10g_tx_pcs_tx_data_out_krfec[42], w_hssi_10g_tx_pcs_tx_data_out_krfec[41], w_hssi_10g_tx_pcs_tx_data_out_krfec[40], w_hssi_10g_tx_pcs_tx_data_out_krfec[39], w_hssi_10g_tx_pcs_tx_data_out_krfec[38], w_hssi_10g_tx_pcs_tx_data_out_krfec[37], w_hssi_10g_tx_pcs_tx_data_out_krfec[36], w_hssi_10g_tx_pcs_tx_data_out_krfec[35], w_hssi_10g_tx_pcs_tx_data_out_krfec[34], w_hssi_10g_tx_pcs_tx_data_out_krfec[33], w_hssi_10g_tx_pcs_tx_data_out_krfec[32], w_hssi_10g_tx_pcs_tx_data_out_krfec[31], w_hssi_10g_tx_pcs_tx_data_out_krfec[30], w_hssi_10g_tx_pcs_tx_data_out_krfec[29], w_hssi_10g_tx_pcs_tx_data_out_krfec[28], w_hssi_10g_tx_pcs_tx_data_out_krfec[27], w_hssi_10g_tx_pcs_tx_data_out_krfec[26], w_hssi_10g_tx_pcs_tx_data_out_krfec[25], w_hssi_10g_tx_pcs_tx_data_out_krfec[24], w_hssi_10g_tx_pcs_tx_data_out_krfec[23], w_hssi_10g_tx_pcs_tx_data_out_krfec[22], w_hssi_10g_tx_pcs_tx_data_out_krfec[21], w_hssi_10g_tx_pcs_tx_data_out_krfec[20], w_hssi_10g_tx_pcs_tx_data_out_krfec[19], w_hssi_10g_tx_pcs_tx_data_out_krfec[18], w_hssi_10g_tx_pcs_tx_data_out_krfec[17], w_hssi_10g_tx_pcs_tx_data_out_krfec[16], w_hssi_10g_tx_pcs_tx_data_out_krfec[15], w_hssi_10g_tx_pcs_tx_data_out_krfec[14], w_hssi_10g_tx_pcs_tx_data_out_krfec[13], w_hssi_10g_tx_pcs_tx_data_out_krfec[12], w_hssi_10g_tx_pcs_tx_data_out_krfec[11], w_hssi_10g_tx_pcs_tx_data_out_krfec[10], w_hssi_10g_tx_pcs_tx_data_out_krfec[9], w_hssi_10g_tx_pcs_tx_data_out_krfec[8], w_hssi_10g_tx_pcs_tx_data_out_krfec[7], w_hssi_10g_tx_pcs_tx_data_out_krfec[6], w_hssi_10g_tx_pcs_tx_data_out_krfec[5], w_hssi_10g_tx_pcs_tx_data_out_krfec[4], w_hssi_10g_tx_pcs_tx_data_out_krfec[3], w_hssi_10g_tx_pcs_tx_data_out_krfec[2], w_hssi_10g_tx_pcs_tx_data_out_krfec[1], w_hssi_10g_tx_pcs_tx_data_out_krfec[0]}),
				.tx_data_valid_in(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
				.tx_krfec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
				.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
				.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
				
				// UNUSED
				.pld_10g_krfec_tx_frame_krfec_reg(),
				.pld_krfec_tx_alignment_plddirect_reg(),
				.pld_krfec_tx_alignment_reg()
			);
		end // if generate
		else begin
				assign w_hssi_krfec_tx_pcs_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_krfec_tx_pcs_blockselect = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_alignment = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_data_out[63:0] = 64'b0;
				assign w_hssi_krfec_tx_pcs_tx_frame = 1'b0;
				assign w_hssi_krfec_tx_pcs_tx_test_data[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen1_2
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen1_2
			twentynm_hssi_pipe_gen1_2 #(
				.elec_idle_delay_val(hssi_pipe_gen1_2_elec_idle_delay_val),
				.error_replace_pad(hssi_pipe_gen1_2_error_replace_pad),
				.hip_mode(hssi_pipe_gen1_2_hip_mode),
				.ind_error_reporting(hssi_pipe_gen1_2_ind_error_reporting),
				.phystatus_delay_val(hssi_pipe_gen1_2_phystatus_delay_val),
				.phystatus_rst_toggle(hssi_pipe_gen1_2_phystatus_rst_toggle),
				.pipe_byte_de_serializer_en(hssi_pipe_gen1_2_pipe_byte_de_serializer_en),
				.prot_mode(hssi_pipe_gen1_2_prot_mode),
				.reconfig_settings(hssi_pipe_gen1_2_reconfig_settings),
				.rx_pipe_enable(hssi_pipe_gen1_2_rx_pipe_enable),
				.rxdetect_bypass(hssi_pipe_gen1_2_rxdetect_bypass),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen1_2_sup_mode),
				.tx_pipe_enable(hssi_pipe_gen1_2_tx_pipe_enable),
				.txswing(hssi_pipe_gen1_2_txswing)
			) inst_twentynm_hssi_pipe_gen1_2 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen1_2_avmmreaddata),
				.blockselect(w_hssi_pipe_gen1_2_blockselect),
				.current_coeff(w_hssi_pipe_gen1_2_current_coeff),
				.phystatus(w_hssi_pipe_gen1_2_phystatus),
				.polarity_inversion_rx(w_hssi_pipe_gen1_2_polarity_inversion_rx),
				.rev_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
				.rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.rxelectricalidle_out(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxstatus(w_hssi_pipe_gen1_2_rxstatus),
				.rxvalid(w_hssi_pipe_gen1_2_rxvalid),
				.tx_elec_idle_out(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.pcie_switch(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]),
				.pipe_rx_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
				.power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
				.power_state_transition_done_ena(1'b0),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
				.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
				.rev_loopbk_pcs_gen3(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.revloopback(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
				.rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.rx_pipe_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
				.rxd({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxelectricalidle(w_hssi_8g_rx_pcs_eidle_detected),
				.rxelectricalidle_pcs_gen3(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.rxpolarity_pcs_gen3(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.speed_change(w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]),
				.tx_elec_idle_comp(w_hssi_8g_tx_pcs_tx_pipe_electidle),
				.tx_pipe_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
				.txd_ch({w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1], w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]}),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswingport(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.pld_8g_rxpolarity_pipe3_reg(),
				.rxd_ch(),
				.txd()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen1_2_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen1_2_blockselect = 1'b0;
				assign w_hssi_pipe_gen1_2_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen1_2_phystatus = 1'b0;
				assign w_hssi_pipe_gen1_2_polarity_inversion_rx = 1'b0;
				assign w_hssi_pipe_gen1_2_rev_loopbk = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen1_2_rxelectricalidle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen1_2_rxvalid = 1'b0;
				assign w_hssi_pipe_gen1_2_tx_elec_idle_out = 1'b0;
				assign w_hssi_pipe_gen1_2_txdetectrx = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_pipe_gen3
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_pipe_gen3
			twentynm_hssi_pipe_gen3 #(
				.bypass_rx_detection_enable(hssi_pipe_gen3_bypass_rx_detection_enable),
				.bypass_rx_preset(hssi_pipe_gen3_bypass_rx_preset),
				.bypass_rx_preset_enable(hssi_pipe_gen3_bypass_rx_preset_enable),
				.bypass_tx_coefficent(hssi_pipe_gen3_bypass_tx_coefficent),
				.bypass_tx_coefficent_enable(hssi_pipe_gen3_bypass_tx_coefficent_enable),
				.elecidle_delay_g3(hssi_pipe_gen3_elecidle_delay_g3),
				.ind_error_reporting(hssi_pipe_gen3_ind_error_reporting),
				.mode(hssi_pipe_gen3_mode),
				.phy_status_delay_g12(hssi_pipe_gen3_phy_status_delay_g12),
				.phy_status_delay_g3(hssi_pipe_gen3_phy_status_delay_g3),
				.phystatus_rst_toggle_g12(hssi_pipe_gen3_phystatus_rst_toggle_g12),
				.phystatus_rst_toggle_g3(hssi_pipe_gen3_phystatus_rst_toggle_g3),
				.rate_match_pad_insertion(hssi_pipe_gen3_rate_match_pad_insertion),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sup_mode(hssi_pipe_gen3_sup_mode),
				.test_out_sel(hssi_pipe_gen3_test_out_sel)
			) inst_twentynm_hssi_pipe_gen3 (
				// OUTPUTS
				.avmmreaddata(w_hssi_pipe_gen3_avmmreaddata),
				.blockselect(w_hssi_pipe_gen3_blockselect),
				.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
				.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
				.phystatus(w_hssi_pipe_gen3_phystatus),
				.pma_current_coeff(w_hssi_pipe_gen3_pma_current_coeff),
				.pma_current_rxpreset(w_hssi_pipe_gen3_pma_current_rxpreset),
				.pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
				.rev_lpbk_8gpcs_out(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
				.rev_lpbk_int(w_hssi_pipe_gen3_rev_lpbk_int),
				.rx_blk_start(w_hssi_pipe_gen3_rx_blk_start),
				.rx_sync_hdr(w_hssi_pipe_gen3_rx_sync_hdr),
				.rxd_8gpcs_out(w_hssi_pipe_gen3_rxd_8gpcs_out),
				.rxdataskip(w_hssi_pipe_gen3_rxdataskip),
				.rxelecidle(w_hssi_pipe_gen3_rxelecidle),
				.rxpolarity_8gpcs_out(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
				.rxpolarity_int(w_hssi_pipe_gen3_rxpolarity_int),
				.rxstatus(w_hssi_pipe_gen3_rxstatus),
				.rxvalid(w_hssi_pipe_gen3_rxvalid),
				.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
				.test_out(w_hssi_pipe_gen3_test_out),
				.tx_blk_start_int(w_hssi_pipe_gen3_tx_blk_start_int),
				.tx_sync_hdr_int(w_hssi_pipe_gen3_tx_sync_hdr_int),
				.txdata_int(w_hssi_pipe_gen3_txdata_int),
				.txdatak_int(w_hssi_pipe_gen3_txdatak_int),
				.txdataskip_int(w_hssi_pipe_gen3_txdataskip_int),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
				.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
				.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
				.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
				.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
				.current_coeff({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0]}),
				.current_rxpreset({w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1], w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0]}),
				.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
				.pcs_asn_bundling_in({w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1], w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0]}),
				.pipe_tx_clk(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
				.pipe_tx_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
				.pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.powerdown({w_hssi_8g_tx_pcs_pipe_power_down_out[1], w_hssi_8g_tx_pcs_pipe_power_down_out[0]}),
				.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
				.rx_blk_start_int(w_hssi_gen3_rx_pcs_blk_start),
				.rx_sync_hdr_int({w_hssi_gen3_rx_pcs_sync_hdr[1], w_hssi_gen3_rx_pcs_sync_hdr[0]}),
				.rx_test_out({w_hssi_gen3_rx_pcs_rx_test_out[19], w_hssi_gen3_rx_pcs_rx_test_out[18], w_hssi_gen3_rx_pcs_rx_test_out[17], w_hssi_gen3_rx_pcs_rx_test_out[16], w_hssi_gen3_rx_pcs_rx_test_out[15], w_hssi_gen3_rx_pcs_rx_test_out[14], w_hssi_gen3_rx_pcs_rx_test_out[13], w_hssi_gen3_rx_pcs_rx_test_out[12], w_hssi_gen3_rx_pcs_rx_test_out[11], w_hssi_gen3_rx_pcs_rx_test_out[10], w_hssi_gen3_rx_pcs_rx_test_out[9], w_hssi_gen3_rx_pcs_rx_test_out[8], w_hssi_gen3_rx_pcs_rx_test_out[7], w_hssi_gen3_rx_pcs_rx_test_out[6], w_hssi_gen3_rx_pcs_rx_test_out[5], w_hssi_gen3_rx_pcs_rx_test_out[4], w_hssi_gen3_rx_pcs_rx_test_out[3], w_hssi_gen3_rx_pcs_rx_test_out[2], w_hssi_gen3_rx_pcs_rx_test_out[1], w_hssi_gen3_rx_pcs_rx_test_out[0]}),
				.rxd_8gpcs_in({w_hssi_8g_rx_pcs_pipe_data[63], w_hssi_8g_rx_pcs_pipe_data[62], w_hssi_8g_rx_pcs_pipe_data[61], w_hssi_8g_rx_pcs_pipe_data[60], w_hssi_8g_rx_pcs_pipe_data[59], w_hssi_8g_rx_pcs_pipe_data[58], w_hssi_8g_rx_pcs_pipe_data[57], w_hssi_8g_rx_pcs_pipe_data[56], w_hssi_8g_rx_pcs_pipe_data[55], w_hssi_8g_rx_pcs_pipe_data[54], w_hssi_8g_rx_pcs_pipe_data[53], w_hssi_8g_rx_pcs_pipe_data[52], w_hssi_8g_rx_pcs_pipe_data[51], w_hssi_8g_rx_pcs_pipe_data[50], w_hssi_8g_rx_pcs_pipe_data[49], w_hssi_8g_rx_pcs_pipe_data[48], w_hssi_8g_rx_pcs_pipe_data[47], w_hssi_8g_rx_pcs_pipe_data[46], w_hssi_8g_rx_pcs_pipe_data[45], w_hssi_8g_rx_pcs_pipe_data[44], w_hssi_8g_rx_pcs_pipe_data[43], w_hssi_8g_rx_pcs_pipe_data[42], w_hssi_8g_rx_pcs_pipe_data[41], w_hssi_8g_rx_pcs_pipe_data[40], w_hssi_8g_rx_pcs_pipe_data[39], w_hssi_8g_rx_pcs_pipe_data[38], w_hssi_8g_rx_pcs_pipe_data[37], w_hssi_8g_rx_pcs_pipe_data[36], w_hssi_8g_rx_pcs_pipe_data[35], w_hssi_8g_rx_pcs_pipe_data[34], w_hssi_8g_rx_pcs_pipe_data[33], w_hssi_8g_rx_pcs_pipe_data[32], w_hssi_8g_rx_pcs_pipe_data[31], w_hssi_8g_rx_pcs_pipe_data[30], w_hssi_8g_rx_pcs_pipe_data[29], w_hssi_8g_rx_pcs_pipe_data[28], w_hssi_8g_rx_pcs_pipe_data[27], w_hssi_8g_rx_pcs_pipe_data[26], w_hssi_8g_rx_pcs_pipe_data[25], w_hssi_8g_rx_pcs_pipe_data[24], w_hssi_8g_rx_pcs_pipe_data[23], w_hssi_8g_rx_pcs_pipe_data[22], w_hssi_8g_rx_pcs_pipe_data[21], w_hssi_8g_rx_pcs_pipe_data[20], w_hssi_8g_rx_pcs_pipe_data[19], w_hssi_8g_rx_pcs_pipe_data[18], w_hssi_8g_rx_pcs_pipe_data[17], w_hssi_8g_rx_pcs_pipe_data[16], w_hssi_8g_rx_pcs_pipe_data[15], w_hssi_8g_rx_pcs_pipe_data[14], w_hssi_8g_rx_pcs_pipe_data[13], w_hssi_8g_rx_pcs_pipe_data[12], w_hssi_8g_rx_pcs_pipe_data[11], w_hssi_8g_rx_pcs_pipe_data[10], w_hssi_8g_rx_pcs_pipe_data[9], w_hssi_8g_rx_pcs_pipe_data[8], w_hssi_8g_rx_pcs_pipe_data[7], w_hssi_8g_rx_pcs_pipe_data[6], w_hssi_8g_rx_pcs_pipe_data[5], w_hssi_8g_rx_pcs_pipe_data[4], w_hssi_8g_rx_pcs_pipe_data[3], w_hssi_8g_rx_pcs_pipe_data[2], w_hssi_8g_rx_pcs_pipe_data[1], w_hssi_8g_rx_pcs_pipe_data[0]}),
				.rxdata_int({w_hssi_gen3_rx_pcs_data_out[31], w_hssi_gen3_rx_pcs_data_out[30], w_hssi_gen3_rx_pcs_data_out[29], w_hssi_gen3_rx_pcs_data_out[28], w_hssi_gen3_rx_pcs_data_out[27], w_hssi_gen3_rx_pcs_data_out[26], w_hssi_gen3_rx_pcs_data_out[25], w_hssi_gen3_rx_pcs_data_out[24], w_hssi_gen3_rx_pcs_data_out[23], w_hssi_gen3_rx_pcs_data_out[22], w_hssi_gen3_rx_pcs_data_out[21], w_hssi_gen3_rx_pcs_data_out[20], w_hssi_gen3_rx_pcs_data_out[19], w_hssi_gen3_rx_pcs_data_out[18], w_hssi_gen3_rx_pcs_data_out[17], w_hssi_gen3_rx_pcs_data_out[16], w_hssi_gen3_rx_pcs_data_out[15], w_hssi_gen3_rx_pcs_data_out[14], w_hssi_gen3_rx_pcs_data_out[13], w_hssi_gen3_rx_pcs_data_out[12], w_hssi_gen3_rx_pcs_data_out[11], w_hssi_gen3_rx_pcs_data_out[10], w_hssi_gen3_rx_pcs_data_out[9], w_hssi_gen3_rx_pcs_data_out[8], w_hssi_gen3_rx_pcs_data_out[7], w_hssi_gen3_rx_pcs_data_out[6], w_hssi_gen3_rx_pcs_data_out[5], w_hssi_gen3_rx_pcs_data_out[4], w_hssi_gen3_rx_pcs_data_out[3], w_hssi_gen3_rx_pcs_data_out[2], w_hssi_gen3_rx_pcs_data_out[1], w_hssi_gen3_rx_pcs_data_out[0]}),
				.rxdatak_int({1'b0, 1'b0, 1'b0, 1'b0}),
				.rxdataskip_int(w_hssi_gen3_rx_pcs_data_valid),
				.rxelecidle_8gpcs_in(w_hssi_pipe_gen1_2_rxelectricalidle_out),
				.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
				.tx_blk_start(w_hssi_8g_tx_pcs_tx_blk_start_out[0]),
				.tx_sync_hdr({w_hssi_8g_tx_pcs_tx_sync_hdr_out[1], w_hssi_8g_tx_pcs_tx_sync_hdr_out[0]}),
				.tx_test_out({w_hssi_gen3_tx_pcs_tx_test_out[19], w_hssi_gen3_tx_pcs_tx_test_out[18], w_hssi_gen3_tx_pcs_tx_test_out[17], w_hssi_gen3_tx_pcs_tx_test_out[16], w_hssi_gen3_tx_pcs_tx_test_out[15], w_hssi_gen3_tx_pcs_tx_test_out[14], w_hssi_gen3_tx_pcs_tx_test_out[13], w_hssi_gen3_tx_pcs_tx_test_out[12], w_hssi_gen3_tx_pcs_tx_test_out[11], w_hssi_gen3_tx_pcs_tx_test_out[10], w_hssi_gen3_tx_pcs_tx_test_out[9], w_hssi_gen3_tx_pcs_tx_test_out[8], w_hssi_gen3_tx_pcs_tx_test_out[7], w_hssi_gen3_tx_pcs_tx_test_out[6], w_hssi_gen3_tx_pcs_tx_test_out[5], w_hssi_gen3_tx_pcs_tx_test_out[4], w_hssi_gen3_tx_pcs_tx_test_out[3], w_hssi_gen3_tx_pcs_tx_test_out[2], w_hssi_gen3_tx_pcs_tx_test_out[1], w_hssi_gen3_tx_pcs_tx_test_out[0]}),
				.txcompliance(w_hssi_8g_tx_pcs_txcompliance_out),
				.txdata({w_hssi_8g_tx_pcs_tx_data_out[31], w_hssi_8g_tx_pcs_tx_data_out[30], w_hssi_8g_tx_pcs_tx_data_out[29], w_hssi_8g_tx_pcs_tx_data_out[28], w_hssi_8g_tx_pcs_tx_data_out[27], w_hssi_8g_tx_pcs_tx_data_out[26], w_hssi_8g_tx_pcs_tx_data_out[25], w_hssi_8g_tx_pcs_tx_data_out[24], w_hssi_8g_tx_pcs_tx_data_out[23], w_hssi_8g_tx_pcs_tx_data_out[22], w_hssi_8g_tx_pcs_tx_data_out[21], w_hssi_8g_tx_pcs_tx_data_out[20], w_hssi_8g_tx_pcs_tx_data_out[19], w_hssi_8g_tx_pcs_tx_data_out[18], w_hssi_8g_tx_pcs_tx_data_out[17], w_hssi_8g_tx_pcs_tx_data_out[16], w_hssi_8g_tx_pcs_tx_data_out[15], w_hssi_8g_tx_pcs_tx_data_out[14], w_hssi_8g_tx_pcs_tx_data_out[13], w_hssi_8g_tx_pcs_tx_data_out[12], w_hssi_8g_tx_pcs_tx_data_out[11], w_hssi_8g_tx_pcs_tx_data_out[10], w_hssi_8g_tx_pcs_tx_data_out[9], w_hssi_8g_tx_pcs_tx_data_out[8], w_hssi_8g_tx_pcs_tx_data_out[7], w_hssi_8g_tx_pcs_tx_data_out[6], w_hssi_8g_tx_pcs_tx_data_out[5], w_hssi_8g_tx_pcs_tx_data_out[4], w_hssi_8g_tx_pcs_tx_data_out[3], w_hssi_8g_tx_pcs_tx_data_out[2], w_hssi_8g_tx_pcs_tx_data_out[1], w_hssi_8g_tx_pcs_tx_data_out[0]}),
				.txdatak({w_hssi_8g_tx_pcs_tx_datak_out[3], w_hssi_8g_tx_pcs_tx_datak_out[2], w_hssi_8g_tx_pcs_tx_datak_out[1], w_hssi_8g_tx_pcs_tx_datak_out[0]}),
				.txdataskip(w_hssi_8g_tx_pcs_tx_data_valid_out[0]),
				.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
				.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
				.txelecidle(w_hssi_8g_tx_pcs_txelecidle_out),
				.txmargin({w_hssi_8g_tx_pcs_phfifo_txmargin[2], w_hssi_8g_tx_pcs_phfifo_txmargin[1], w_hssi_8g_tx_pcs_phfifo_txmargin[0]}),
				.txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
				
				// UNUSED
				.dis_pc_byte(),
				.pma_rx_det_pd(),
				.pma_txdeemph(),
				.pma_txmargin(),
				.pma_txswing(),
				.reset_pc_prts()
			);
		end // if generate
		else begin
				assign w_hssi_pipe_gen3_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_pipe_gen3_blockselect = 1'b0;
				assign w_hssi_pipe_gen3_gen3_clk_sel = 1'b0;
				assign w_hssi_pipe_gen3_pcs_rst = 1'b0;
				assign w_hssi_pipe_gen3_phystatus = 1'b0;
				assign w_hssi_pipe_gen3_pma_current_coeff[17:0] = 18'b0;
				assign w_hssi_pipe_gen3_pma_current_rxpreset[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_pma_tx_elec_idle = 1'b0;
				assign w_hssi_pipe_gen3_pma_txdetectrx = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rev_lpbk_int = 1'b0;
				assign w_hssi_pipe_gen3_rx_blk_start[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_rxd_8gpcs_out[63:0] = 64'b0;
				assign w_hssi_pipe_gen3_rxdataskip[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_rxelecidle = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_8gpcs_out = 1'b0;
				assign w_hssi_pipe_gen3_rxpolarity_int = 1'b0;
				assign w_hssi_pipe_gen3_rxstatus[2:0] = 3'b0;
				assign w_hssi_pipe_gen3_rxvalid = 1'b0;
				assign w_hssi_pipe_gen3_shutdown_clk = 1'b0;
				assign w_hssi_pipe_gen3_test_out[19:0] = 20'b0;
				assign w_hssi_pipe_gen3_tx_blk_start_int = 1'b0;
				assign w_hssi_pipe_gen3_tx_sync_hdr_int[1:0] = 2'b0;
				assign w_hssi_pipe_gen3_txdata_int[31:0] = 32'b0;
				assign w_hssi_pipe_gen3_txdatak_int[3:0] = 4'b0;
				assign w_hssi_pipe_gen3_txdataskip_int = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pcs_pma_interface
			twentynm_hssi_rx_pcs_pma_interface #(
				.block_sel(hssi_rx_pcs_pma_interface_block_sel),
				.channel_operation_mode(hssi_rx_pcs_pma_interface_channel_operation_mode),
				.clkslip_sel(hssi_rx_pcs_pma_interface_clkslip_sel),
				.lpbk_en(hssi_rx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_rx_pcs_pma_interface_master_clk_sel),
				.pldif_datawidth_mode(hssi_rx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_rx(hssi_rx_pcs_pma_interface_pma_dw_rx),
				.pma_if_dft_en(hssi_rx_pcs_pma_interface_pma_if_dft_en),
				.pma_if_dft_val(hssi_rx_pcs_pma_interface_pma_if_dft_val),
				.prbs9_dwidth(hssi_rx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_rx_pcs_pma_interface_prbs_clken),
				.prbs_ver(hssi_rx_pcs_pma_interface_prbs_ver),
				.prot_mode_rx(hssi_rx_pcs_pma_interface_prot_mode_rx),
				.reconfig_settings(hssi_rx_pcs_pma_interface_reconfig_settings),
				.rx_dyn_polarity_inversion(hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion),
				.rx_lpbk_en(hssi_rx_pcs_pma_interface_rx_lpbk_en),
				.rx_prbs_force_signal_ok(hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok),
				.rx_prbs_mask(hssi_rx_pcs_pma_interface_rx_prbs_mask),
				.rx_prbs_mode(hssi_rx_pcs_pma_interface_rx_prbs_mode),
				.rx_signalok_signaldet_sel(hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel),
				.rx_static_polarity_inversion(hssi_rx_pcs_pma_interface_rx_static_polarity_inversion),
				.rx_uhsif_lpbk_en(hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sup_mode(hssi_rx_pcs_pma_interface_sup_mode)
			) inst_twentynm_hssi_rx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
				.int_pmaif_10g_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data),
				.int_pmaif_10g_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
				.int_pmaif_8g_pudi(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi),
				.int_pmaif_8g_rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
				.int_pmaif_8g_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
				.int_pmaif_8g_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
				.int_pmaif_8g_sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
				.int_pmaif_g3_pma_data_in(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in),
				.int_pmaif_g3_pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
				.int_pmaif_g3_pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
				.int_pmaif_g3_pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
				.int_pmaif_krfec_rx_pma_data(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data),
				.int_pmaif_krfec_rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
				.int_pmaif_pldif_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pmaif_pldif_prbs_err_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pmaif_pldif_rx_clkdiv(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pmaif_pldif_rx_clkdiv_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pmaif_pldif_rx_data(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data),
				.int_pmaif_pldif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
				.int_pmaif_pldif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
				.int_pmaif_pldif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pmaif_pldif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
				.pma_eye_monitor(w_hssi_rx_pcs_pma_interface_pma_eye_monitor),
				.pma_rx_clkslip(w_hssi_rx_pcs_pma_interface_pma_rx_clkslip),
				.pma_rxpma_rstb(w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb),
				.rx_pmaif_test_out(w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out),
				.rx_prbs_ver_test(w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_random_err(w_hssi_10g_rx_pcs_rx_random_err),
				.int_pmaif_8g_rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
				.int_pmaif_pldif_eye_monitor({w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1], w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0]}),
				.int_pmaif_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pmaif_pldif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pmaif_pldif_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pmaif_pldif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pma_rx_clkdiv_user(in_pma_rx_clkdiv_user),
				.pma_rx_detect_valid(in_pma_rx_detect_valid),
				.pma_rx_found(in_pma_rx_found),
				.pma_rx_pma_clk(in_pma_rx_pma_clk),
				.pma_rx_pma_data({in_pma_rx_pma_data[63], in_pma_rx_pma_data[62], in_pma_rx_pma_data[61], in_pma_rx_pma_data[60], in_pma_rx_pma_data[59], in_pma_rx_pma_data[58], in_pma_rx_pma_data[57], in_pma_rx_pma_data[56], in_pma_rx_pma_data[55], in_pma_rx_pma_data[54], in_pma_rx_pma_data[53], in_pma_rx_pma_data[52], in_pma_rx_pma_data[51], in_pma_rx_pma_data[50], in_pma_rx_pma_data[49], in_pma_rx_pma_data[48], in_pma_rx_pma_data[47], in_pma_rx_pma_data[46], in_pma_rx_pma_data[45], in_pma_rx_pma_data[44], in_pma_rx_pma_data[43], in_pma_rx_pma_data[42], in_pma_rx_pma_data[41], in_pma_rx_pma_data[40], in_pma_rx_pma_data[39], in_pma_rx_pma_data[38], in_pma_rx_pma_data[37], in_pma_rx_pma_data[36], in_pma_rx_pma_data[35], in_pma_rx_pma_data[34], in_pma_rx_pma_data[33], in_pma_rx_pma_data[32], in_pma_rx_pma_data[31], in_pma_rx_pma_data[30], in_pma_rx_pma_data[29], in_pma_rx_pma_data[28], in_pma_rx_pma_data[27], in_pma_rx_pma_data[26], in_pma_rx_pma_data[25], in_pma_rx_pma_data[24], in_pma_rx_pma_data[23], in_pma_rx_pma_data[22], in_pma_rx_pma_data[21], in_pma_rx_pma_data[20], in_pma_rx_pma_data[19], in_pma_rx_pma_data[18], in_pma_rx_pma_data[17], in_pma_rx_pma_data[16], in_pma_rx_pma_data[15], in_pma_rx_pma_data[14], in_pma_rx_pma_data[13], in_pma_rx_pma_data[12], in_pma_rx_pma_data[11], in_pma_rx_pma_data[10], in_pma_rx_pma_data[9], in_pma_rx_pma_data[8], in_pma_rx_pma_data[7], in_pma_rx_pma_data[6], in_pma_rx_pma_data[5], in_pma_rx_pma_data[4], in_pma_rx_pma_data[3], in_pma_rx_pma_data[2], in_pma_rx_pma_data[1], in_pma_rx_pma_data[0]}),
				.pma_rx_signal_ok(in_pma_rx_signal_ok),
				.pma_rxpll_lock(in_pma_rxpll_lock),
				.pma_signal_det(in_pma_signal_det),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.tx_pma_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0]}),
				.tx_pma_uhsif_data_loopback({w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1], w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0]}),
				
				// UNUSED
				.int_pmaif_g3_rcvd_clk(),
				.prbs_err_lt()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31:0] = 32'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63:0] = 64'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5:0] = 6'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rx_clkslip = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19:0] = 20'b0;
				assign w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_rx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_rx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_rx_pld_pcs_interface
			twentynm_hssi_rx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx),
				.hd_10g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_rx),
				.hd_10g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx),
				.hd_10g_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx),
				.hd_10g_lpbk_en(hssi_rx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx),
				.hd_10g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx),
				.hd_10g_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx),
				.hd_10g_test_bus_mode(hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode),
				.hd_8g_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_rx),
				.hd_8g_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx),
				.hd_8g_hip_mode(hssi_rx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_rx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx),
				.hd_8g_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx),
				.hd_chnl_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_clklow_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz),
				.hd_chnl_ctrl_plane_bonding_rx(hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx),
				.hd_chnl_fref_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz),
				.hd_chnl_frequency_rules_en(hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_rx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_rx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx),
				.hd_chnl_lpbk_en(hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx),
				.hd_chnl_pld_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz),
				.hd_chnl_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx),
				.hd_chnl_pma_rx_clk_hz(hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz),
				.hd_chnl_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx),
				.hd_chnl_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx),
				.hd_chnl_transparent_pcs_rx(hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx),
				.hd_fifo_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx),
				.hd_fifo_shared_fifo_width_rx(hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx),
				.hd_g3_prot_mode(hssi_rx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_rx(hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx),
				.hd_krfec_lpbk_en(hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx),
				.hd_krfec_test_bus_mode(hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode),
				.hd_pldif_hrdrstctl_en(hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx),
				.hd_pmaif_channel_operation_mode(hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_lpbk_en(hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_rx(hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx),
				.hd_pmaif_prot_mode_rx(hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx),
				.hd_pmaif_sim_mode(hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_rx_block_sel(hssi_rx_pld_pcs_interface_pcs_rx_block_sel),
				.pcs_rx_clk_out_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel),
				.pcs_rx_clk_sel(hssi_rx_pld_pcs_interface_pcs_rx_clk_sel),
				.pcs_rx_hip_clk_en(hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en),
				.pcs_rx_output_sel(hssi_rx_pld_pcs_interface_pcs_rx_output_sel),
				.reconfig_settings(hssi_rx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm4es" )       //PARAM_HIDE
			) inst_twentynm_hssi_rx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_rx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_rx_pld_pcs_interface_blockselect),
				.hip_rx_ctrl(w_hssi_rx_pld_pcs_interface_hip_rx_ctrl),
				.hip_rx_data(w_hssi_rx_pld_pcs_interface_hip_rx_data),
				.int_pldif_10g_rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
				.int_pldif_10g_rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
				.int_pldif_10g_rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
				.int_pldif_10g_rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
				.int_pldif_10g_rx_control_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb),
				.int_pldif_10g_rx_data_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb),
				.int_pldif_10g_rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
				.int_pldif_10g_rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
				.int_pldif_10g_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
				.int_pldif_10g_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
				.int_pldif_10g_rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
				.int_pldif_8g_a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
				.int_pldif_8g_bitloc_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
				.int_pldif_8g_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
				.int_pldif_8g_byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
				.int_pldif_8g_encdt(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
				.int_pldif_8g_pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
				.int_pldif_8g_rdenable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
				.int_pldif_8g_rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
				.int_pldif_8g_rxurstpcs_n(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
				.int_pldif_8g_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
				.int_pldif_8g_wrdisable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
				.int_pldif_g3_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
				.int_pldif_krfec_rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
				.int_pldif_pmaif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
				.int_pldif_pmaif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
				.int_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
				.int_pldif_pmaif_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
				.int_pldif_pmaif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
				.pld_10g_krfec_rx_blk_lock(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock),
				.pld_10g_krfec_rx_diag_data_status(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status),
				.pld_10g_krfec_rx_frame(w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame),
				.pld_10g_rx_align_val(w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val),
				.pld_10g_rx_crc32_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err),
				.pld_10g_rx_data_valid(w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid),
				.pld_10g_rx_empty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty),
				.pld_10g_rx_fifo_del(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del),
				.pld_10g_rx_fifo_insert(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert),
				.pld_10g_rx_fifo_num(w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num),
				.pld_10g_rx_frame_lock(w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock),
				.pld_10g_rx_hi_ber(w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber),
				.pld_10g_rx_oflw_err(w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err),
				.pld_10g_rx_pempty(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty),
				.pld_10g_rx_pfull(w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull),
				.pld_8g_a1a2_k1k2_flag(w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag),
				.pld_8g_empty_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf),
				.pld_8g_empty_rx(w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx),
				.pld_8g_full_rmf(w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf),
				.pld_8g_full_rx(w_hssi_rx_pld_pcs_interface_pld_8g_full_rx),
				.pld_8g_rxelecidle(w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle),
				.pld_8g_signal_detect_out(w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out),
				.pld_8g_wa_boundary(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary),
				.pld_pcs_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out),
				.pld_pma_clkdiv_rx_user(w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user),
				.pld_pma_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out),
				.pld_pma_signal_ok(w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok),
				.pld_rx_control(w_hssi_rx_pld_pcs_interface_pld_rx_control),
				.pld_rx_data(w_hssi_rx_pld_pcs_interface_pld_rx_data),
				.pld_rx_prbs_done(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done),
				.pld_rx_prbs_err(w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pldif_10g_rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
				.int_pldif_10g_rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
				.int_pldif_10g_rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
				.int_pldif_10g_rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_10g_rx_control({w_hssi_10g_rx_pcs_rx_control[19], w_hssi_10g_rx_pcs_rx_control[18], w_hssi_10g_rx_pcs_rx_control[17], w_hssi_10g_rx_pcs_rx_control[16], w_hssi_10g_rx_pcs_rx_control[15], w_hssi_10g_rx_pcs_rx_control[14], w_hssi_10g_rx_pcs_rx_control[13], w_hssi_10g_rx_pcs_rx_control[12], w_hssi_10g_rx_pcs_rx_control[11], w_hssi_10g_rx_pcs_rx_control[10], w_hssi_10g_rx_pcs_rx_control[9], w_hssi_10g_rx_pcs_rx_control[8], w_hssi_10g_rx_pcs_rx_control[7], w_hssi_10g_rx_pcs_rx_control[6], w_hssi_10g_rx_pcs_rx_control[5], w_hssi_10g_rx_pcs_rx_control[4], w_hssi_10g_rx_pcs_rx_control[3], w_hssi_10g_rx_pcs_rx_control[2], w_hssi_10g_rx_pcs_rx_control[1], w_hssi_10g_rx_pcs_rx_control[0]}),
				.int_pldif_10g_rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
				.int_pldif_10g_rx_data({w_hssi_10g_rx_pcs_rx_data[127], w_hssi_10g_rx_pcs_rx_data[126], w_hssi_10g_rx_pcs_rx_data[125], w_hssi_10g_rx_pcs_rx_data[124], w_hssi_10g_rx_pcs_rx_data[123], w_hssi_10g_rx_pcs_rx_data[122], w_hssi_10g_rx_pcs_rx_data[121], w_hssi_10g_rx_pcs_rx_data[120], w_hssi_10g_rx_pcs_rx_data[119], w_hssi_10g_rx_pcs_rx_data[118], w_hssi_10g_rx_pcs_rx_data[117], w_hssi_10g_rx_pcs_rx_data[116], w_hssi_10g_rx_pcs_rx_data[115], w_hssi_10g_rx_pcs_rx_data[114], w_hssi_10g_rx_pcs_rx_data[113], w_hssi_10g_rx_pcs_rx_data[112], w_hssi_10g_rx_pcs_rx_data[111], w_hssi_10g_rx_pcs_rx_data[110], w_hssi_10g_rx_pcs_rx_data[109], w_hssi_10g_rx_pcs_rx_data[108], w_hssi_10g_rx_pcs_rx_data[107], w_hssi_10g_rx_pcs_rx_data[106], w_hssi_10g_rx_pcs_rx_data[105], w_hssi_10g_rx_pcs_rx_data[104], w_hssi_10g_rx_pcs_rx_data[103], w_hssi_10g_rx_pcs_rx_data[102], w_hssi_10g_rx_pcs_rx_data[101], w_hssi_10g_rx_pcs_rx_data[100], w_hssi_10g_rx_pcs_rx_data[99], w_hssi_10g_rx_pcs_rx_data[98], w_hssi_10g_rx_pcs_rx_data[97], w_hssi_10g_rx_pcs_rx_data[96], w_hssi_10g_rx_pcs_rx_data[95], w_hssi_10g_rx_pcs_rx_data[94], w_hssi_10g_rx_pcs_rx_data[93], w_hssi_10g_rx_pcs_rx_data[92], w_hssi_10g_rx_pcs_rx_data[91], w_hssi_10g_rx_pcs_rx_data[90], w_hssi_10g_rx_pcs_rx_data[89], w_hssi_10g_rx_pcs_rx_data[88], w_hssi_10g_rx_pcs_rx_data[87], w_hssi_10g_rx_pcs_rx_data[86], w_hssi_10g_rx_pcs_rx_data[85], w_hssi_10g_rx_pcs_rx_data[84], w_hssi_10g_rx_pcs_rx_data[83], w_hssi_10g_rx_pcs_rx_data[82], w_hssi_10g_rx_pcs_rx_data[81], w_hssi_10g_rx_pcs_rx_data[80], w_hssi_10g_rx_pcs_rx_data[79], w_hssi_10g_rx_pcs_rx_data[78], w_hssi_10g_rx_pcs_rx_data[77], w_hssi_10g_rx_pcs_rx_data[76], w_hssi_10g_rx_pcs_rx_data[75], w_hssi_10g_rx_pcs_rx_data[74], w_hssi_10g_rx_pcs_rx_data[73], w_hssi_10g_rx_pcs_rx_data[72], w_hssi_10g_rx_pcs_rx_data[71], w_hssi_10g_rx_pcs_rx_data[70], w_hssi_10g_rx_pcs_rx_data[69], w_hssi_10g_rx_pcs_rx_data[68], w_hssi_10g_rx_pcs_rx_data[67], w_hssi_10g_rx_pcs_rx_data[66], w_hssi_10g_rx_pcs_rx_data[65], w_hssi_10g_rx_pcs_rx_data[64], w_hssi_10g_rx_pcs_rx_data[63], w_hssi_10g_rx_pcs_rx_data[62], w_hssi_10g_rx_pcs_rx_data[61], w_hssi_10g_rx_pcs_rx_data[60], w_hssi_10g_rx_pcs_rx_data[59], w_hssi_10g_rx_pcs_rx_data[58], w_hssi_10g_rx_pcs_rx_data[57], w_hssi_10g_rx_pcs_rx_data[56], w_hssi_10g_rx_pcs_rx_data[55], w_hssi_10g_rx_pcs_rx_data[54], w_hssi_10g_rx_pcs_rx_data[53], w_hssi_10g_rx_pcs_rx_data[52], w_hssi_10g_rx_pcs_rx_data[51], w_hssi_10g_rx_pcs_rx_data[50], w_hssi_10g_rx_pcs_rx_data[49], w_hssi_10g_rx_pcs_rx_data[48], w_hssi_10g_rx_pcs_rx_data[47], w_hssi_10g_rx_pcs_rx_data[46], w_hssi_10g_rx_pcs_rx_data[45], w_hssi_10g_rx_pcs_rx_data[44], w_hssi_10g_rx_pcs_rx_data[43], w_hssi_10g_rx_pcs_rx_data[42], w_hssi_10g_rx_pcs_rx_data[41], w_hssi_10g_rx_pcs_rx_data[40], w_hssi_10g_rx_pcs_rx_data[39], w_hssi_10g_rx_pcs_rx_data[38], w_hssi_10g_rx_pcs_rx_data[37], w_hssi_10g_rx_pcs_rx_data[36], w_hssi_10g_rx_pcs_rx_data[35], w_hssi_10g_rx_pcs_rx_data[34], w_hssi_10g_rx_pcs_rx_data[33], w_hssi_10g_rx_pcs_rx_data[32], w_hssi_10g_rx_pcs_rx_data[31], w_hssi_10g_rx_pcs_rx_data[30], w_hssi_10g_rx_pcs_rx_data[29], w_hssi_10g_rx_pcs_rx_data[28], w_hssi_10g_rx_pcs_rx_data[27], w_hssi_10g_rx_pcs_rx_data[26], w_hssi_10g_rx_pcs_rx_data[25], w_hssi_10g_rx_pcs_rx_data[24], w_hssi_10g_rx_pcs_rx_data[23], w_hssi_10g_rx_pcs_rx_data[22], w_hssi_10g_rx_pcs_rx_data[21], w_hssi_10g_rx_pcs_rx_data[20], w_hssi_10g_rx_pcs_rx_data[19], w_hssi_10g_rx_pcs_rx_data[18], w_hssi_10g_rx_pcs_rx_data[17], w_hssi_10g_rx_pcs_rx_data[16], w_hssi_10g_rx_pcs_rx_data[15], w_hssi_10g_rx_pcs_rx_data[14], w_hssi_10g_rx_pcs_rx_data[13], w_hssi_10g_rx_pcs_rx_data[12], w_hssi_10g_rx_pcs_rx_data[11], w_hssi_10g_rx_pcs_rx_data[10], w_hssi_10g_rx_pcs_rx_data[9], w_hssi_10g_rx_pcs_rx_data[8], w_hssi_10g_rx_pcs_rx_data[7], w_hssi_10g_rx_pcs_rx_data[6], w_hssi_10g_rx_pcs_rx_data[5], w_hssi_10g_rx_pcs_rx_data[4], w_hssi_10g_rx_pcs_rx_data[3], w_hssi_10g_rx_pcs_rx_data[2], w_hssi_10g_rx_pcs_rx_data[1], w_hssi_10g_rx_pcs_rx_data[0]}),
				.int_pldif_10g_rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
				.int_pldif_10g_rx_diag_status({w_hssi_10g_rx_pcs_rx_diag_status[1], w_hssi_10g_rx_pcs_rx_diag_status[0]}),
				.int_pldif_10g_rx_empty(w_hssi_10g_rx_pcs_rx_empty),
				.int_pldif_10g_rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
				.int_pldif_10g_rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
				.int_pldif_10g_rx_fifo_num({w_hssi_10g_rx_pcs_rx_fifo_num[4], w_hssi_10g_rx_pcs_rx_fifo_num[3], w_hssi_10g_rx_pcs_rx_fifo_num[2], w_hssi_10g_rx_pcs_rx_fifo_num[1], w_hssi_10g_rx_pcs_rx_fifo_num[0]}),
				.int_pldif_10g_rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
				.int_pldif_10g_rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
				.int_pldif_10g_rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
				.int_pldif_10g_rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
				.int_pldif_10g_rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
				.int_pldif_10g_rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
				.int_pldif_8g_a1a2_k1k2_flag({w_hssi_8g_rx_pcs_a1a2k1k2flag[3], w_hssi_8g_rx_pcs_a1a2k1k2flag[2], w_hssi_8g_rx_pcs_a1a2k1k2flag[1], w_hssi_8g_rx_pcs_a1a2k1k2flag[0]}),
				.int_pldif_8g_empty_rmf(w_hssi_8g_rx_pcs_rm_fifo_empty),
				.int_pldif_8g_empty_rx(w_hssi_8g_rx_pcs_pc_fifo_empty),
				.int_pldif_8g_full_rmf(w_hssi_8g_rx_pcs_rm_fifo_full),
				.int_pldif_8g_full_rx(w_hssi_8g_rx_pcs_pcfifofull),
				.int_pldif_8g_phystatus(w_hssi_8g_rx_pcs_phystatus),
				.int_pldif_8g_rx_blk_start({w_hssi_8g_rx_pcs_rx_blk_start[3], w_hssi_8g_rx_pcs_rx_blk_start[2], w_hssi_8g_rx_pcs_rx_blk_start[1], w_hssi_8g_rx_pcs_rx_blk_start[0]}),
				.int_pldif_8g_rx_clk(w_hssi_8g_rx_pcs_clock_to_pld),
				.int_pldif_8g_rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
				.int_pldif_8g_rx_data_valid({w_hssi_8g_rx_pcs_rx_data_valid[3], w_hssi_8g_rx_pcs_rx_data_valid[2], w_hssi_8g_rx_pcs_rx_data_valid[1], w_hssi_8g_rx_pcs_rx_data_valid[0]}),
				.int_pldif_8g_rx_rstn_sync2wrfifo(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
				.int_pldif_8g_rx_sync_hdr({w_hssi_8g_rx_pcs_rx_sync_hdr[1], w_hssi_8g_rx_pcs_rx_sync_hdr[0]}),
				.int_pldif_8g_rxd({w_hssi_8g_rx_pcs_dataout[63], w_hssi_8g_rx_pcs_dataout[62], w_hssi_8g_rx_pcs_dataout[61], w_hssi_8g_rx_pcs_dataout[60], w_hssi_8g_rx_pcs_dataout[59], w_hssi_8g_rx_pcs_dataout[58], w_hssi_8g_rx_pcs_dataout[57], w_hssi_8g_rx_pcs_dataout[56], w_hssi_8g_rx_pcs_dataout[55], w_hssi_8g_rx_pcs_dataout[54], w_hssi_8g_rx_pcs_dataout[53], w_hssi_8g_rx_pcs_dataout[52], w_hssi_8g_rx_pcs_dataout[51], w_hssi_8g_rx_pcs_dataout[50], w_hssi_8g_rx_pcs_dataout[49], w_hssi_8g_rx_pcs_dataout[48], w_hssi_8g_rx_pcs_dataout[47], w_hssi_8g_rx_pcs_dataout[46], w_hssi_8g_rx_pcs_dataout[45], w_hssi_8g_rx_pcs_dataout[44], w_hssi_8g_rx_pcs_dataout[43], w_hssi_8g_rx_pcs_dataout[42], w_hssi_8g_rx_pcs_dataout[41], w_hssi_8g_rx_pcs_dataout[40], w_hssi_8g_rx_pcs_dataout[39], w_hssi_8g_rx_pcs_dataout[38], w_hssi_8g_rx_pcs_dataout[37], w_hssi_8g_rx_pcs_dataout[36], w_hssi_8g_rx_pcs_dataout[35], w_hssi_8g_rx_pcs_dataout[34], w_hssi_8g_rx_pcs_dataout[33], w_hssi_8g_rx_pcs_dataout[32], w_hssi_8g_rx_pcs_dataout[31], w_hssi_8g_rx_pcs_dataout[30], w_hssi_8g_rx_pcs_dataout[29], w_hssi_8g_rx_pcs_dataout[28], w_hssi_8g_rx_pcs_dataout[27], w_hssi_8g_rx_pcs_dataout[26], w_hssi_8g_rx_pcs_dataout[25], w_hssi_8g_rx_pcs_dataout[24], w_hssi_8g_rx_pcs_dataout[23], w_hssi_8g_rx_pcs_dataout[22], w_hssi_8g_rx_pcs_dataout[21], w_hssi_8g_rx_pcs_dataout[20], w_hssi_8g_rx_pcs_dataout[19], w_hssi_8g_rx_pcs_dataout[18], w_hssi_8g_rx_pcs_dataout[17], w_hssi_8g_rx_pcs_dataout[16], w_hssi_8g_rx_pcs_dataout[15], w_hssi_8g_rx_pcs_dataout[14], w_hssi_8g_rx_pcs_dataout[13], w_hssi_8g_rx_pcs_dataout[12], w_hssi_8g_rx_pcs_dataout[11], w_hssi_8g_rx_pcs_dataout[10], w_hssi_8g_rx_pcs_dataout[9], w_hssi_8g_rx_pcs_dataout[8], w_hssi_8g_rx_pcs_dataout[7], w_hssi_8g_rx_pcs_dataout[6], w_hssi_8g_rx_pcs_dataout[5], w_hssi_8g_rx_pcs_dataout[4], w_hssi_8g_rx_pcs_dataout[3], w_hssi_8g_rx_pcs_dataout[2], w_hssi_8g_rx_pcs_dataout[1], w_hssi_8g_rx_pcs_dataout[0]}),
				.int_pldif_8g_rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
				.int_pldif_8g_rxstatus({w_hssi_8g_rx_pcs_rxstatus[2], w_hssi_8g_rx_pcs_rxstatus[1], w_hssi_8g_rx_pcs_rxstatus[0]}),
				.int_pldif_8g_rxvalid(w_hssi_8g_rx_pcs_rxvalid),
				.int_pldif_8g_signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
				.int_pldif_8g_wa_boundary({w_hssi_8g_rx_pcs_word_align_boundary[4], w_hssi_8g_rx_pcs_word_align_boundary[3], w_hssi_8g_rx_pcs_word_align_boundary[2], w_hssi_8g_rx_pcs_word_align_boundary[1], w_hssi_8g_rx_pcs_word_align_boundary[0]}),
				.int_pldif_krfec_rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
				.int_pldif_krfec_rx_data_status({w_hssi_krfec_rx_pcs_rx_data_status[1], w_hssi_krfec_rx_pcs_rx_data_status[0]}),
				.int_pldif_krfec_rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
				.int_pldif_pmaif_clkdiv_rx(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
				.int_pldif_pmaif_clkdiv_rx_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
				.int_pldif_pmaif_rx_data({w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1], w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0]}),
				.int_pldif_pmaif_rx_prbs_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
				.int_pldif_pmaif_rx_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
				.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
				.int_pldif_pmaif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
				.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
				.pld_10g_krfec_rx_clr_errblk_cnt(in_pld_10g_krfec_rx_clr_errblk_cnt),
				.pld_10g_krfec_rx_pld_rst_n(in_pld_10g_krfec_rx_pld_rst_n),
				.pld_10g_rx_align_clr(in_pld_10g_rx_align_clr),
				.pld_10g_rx_clr_ber_count(in_pld_10g_rx_clr_ber_count),
				.pld_10g_rx_rd_en(in_pld_10g_rx_rd_en),
				.pld_8g_a1a2_size(in_pld_8g_a1a2_size),
				.pld_8g_bitloc_rev_en(in_pld_8g_bitloc_rev_en),
				.pld_8g_byte_rev_en(in_pld_8g_byte_rev_en),
				.pld_8g_encdt(in_pld_8g_encdt),
				.pld_8g_g3_rx_pld_rst_n(in_pld_8g_g3_rx_pld_rst_n),
				.pld_8g_rdenable_rx(in_pld_8g_rdenable_rx),
				.pld_8g_rxpolarity(in_pld_8g_rxpolarity),
				.pld_8g_wrdisable_rx(in_pld_8g_wrdisable_rx),
				.pld_bitslip(in_pld_bitslip),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_rxpma_rstb(in_pld_pma_rxpma_rstb),
				.pld_pmaif_rx_pld_rst_n(in_pld_pmaif_rx_pld_rst_n),
				.pld_pmaif_rxclkslip(in_pld_pmaif_rxclkslip),
				.pld_polinv_rx(in_pld_polinv_rx),
				.pld_rx_clk(in_pld_rx_clk),
				.pld_rx_prbs_err_clr(in_pld_rx_prbs_err_clr),
				.pld_syncsm_en(in_pld_syncsm_en),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.int_pldif_pmaif_rx_pld_clk(),
				.pld_8g_wa_boundary_txclk_fastreg(),
				.pld_8g_wa_boundary_txclk_reg(),
				.pld_bitslip_10g_txclk_reg(),
				.pld_bitslip_8g_txclk_reg(),
				.pld_bitslip_rxclk_parallel_loopback_reg(),
				.pld_bitslip_rxclk_reg(),
				.pld_pcs_rx_clk_out_pcsdirect_wire(),
				.pld_pma_rx_clk_out_10g_or_pcsdirect_wire(),
				.pld_pma_rx_clk_out_8g_wire(),
				.pld_pmaif_rx_pld_rst_n_reg(),
				.pld_pmaif_tx_pld_rst_n_txclk_reg(),
				.pld_polinv_rx_reg(),
				.pld_rx_clk_fifo(),
				.pld_rx_control_fifo(),
				.pld_rx_control_pcsdirect_reg(),
				.pld_rx_data_fifo(),
				.pld_rx_data_pcsdirect_reg(),
				.pld_rx_prbs_done_reg(),
				.pld_rx_prbs_done_txclk_reg(),
				.pld_rx_prbs_err_clr_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_clr_reg(),
				.pld_rx_prbs_err_disprbs_reg(),
				.pld_rx_prbs_err_pcsdirect_txclk_reg(),
				.pld_rx_prbs_err_reg(),
				.pma_rx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_rx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_rx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_hip_rx_data[50:0] = 51'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1:0] = 2'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3:0] = 4'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_full_rx = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4:0] = 5'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_control[19:0] = 20'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_data[127:0] = 128'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done = 1'b0;
				assign w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err = 1'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pcs_pma_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pcs_pma_interface
			twentynm_hssi_tx_pcs_pma_interface #(
				.bypass_pma_txelecidle(hssi_tx_pcs_pma_interface_bypass_pma_txelecidle),
				.channel_operation_mode(hssi_tx_pcs_pma_interface_channel_operation_mode),
				.lpbk_en(hssi_tx_pcs_pma_interface_lpbk_en),
				.master_clk_sel(hssi_tx_pcs_pma_interface_master_clk_sel),
				.pcie_sub_prot_mode_tx(hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx),
				.pldif_datawidth_mode(hssi_tx_pcs_pma_interface_pldif_datawidth_mode),
				.pma_dw_tx(hssi_tx_pcs_pma_interface_pma_dw_tx),
				.pma_if_dft_en(hssi_tx_pcs_pma_interface_pma_if_dft_en),
				.pmagate_en(hssi_tx_pcs_pma_interface_pmagate_en),
				.prbs9_dwidth(hssi_tx_pcs_pma_interface_prbs9_dwidth),
				.prbs_clken(hssi_tx_pcs_pma_interface_prbs_clken),
				.prbs_gen_pat(hssi_tx_pcs_pma_interface_prbs_gen_pat),
				.prot_mode_tx(hssi_tx_pcs_pma_interface_prot_mode_tx),
				.reconfig_settings(hssi_tx_pcs_pma_interface_reconfig_settings),
				.silicon_rev( "20nm4es" ),       //PARAM_HIDE
				.sq_wave_num(hssi_tx_pcs_pma_interface_sq_wave_num),
				.sqwgen_clken(hssi_tx_pcs_pma_interface_sqwgen_clken),
				.sup_mode(hssi_tx_pcs_pma_interface_sup_mode),
				.tx_dyn_polarity_inversion(hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion),
				.tx_pma_data_sel(hssi_tx_pcs_pma_interface_tx_pma_data_sel),
				.tx_static_polarity_inversion(hssi_tx_pcs_pma_interface_tx_static_polarity_inversion),
				.uhsif_cnt_step_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock),
				.uhsif_cnt_thresh_filt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value),
				.uhsif_cnt_thresh_filt_before_lock(hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock),
				.uhsif_dcn_test_update_period(hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period),
				.uhsif_dcn_testmode_enable(hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable),
				.uhsif_dead_zone_count_thresh(hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh),
				.uhsif_dead_zone_detection_enable(hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable),
				.uhsif_dead_zone_obser_window(hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window),
				.uhsif_dead_zone_skip_size(hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size),
				.uhsif_delay_cell_index_sel(hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel),
				.uhsif_delay_cell_margin(hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin),
				.uhsif_delay_cell_static_index_value(hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value),
				.uhsif_dft_dead_zone_control(hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control),
				.uhsif_dft_up_filt_control(hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control),
				.uhsif_enable(hssi_tx_pcs_pma_interface_uhsif_enable),
				.uhsif_lock_det_segsz_after_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock),
				.uhsif_lock_det_segsz_before_lock(hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock),
				.uhsif_lock_det_thresh_cnt_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value),
				.uhsif_lock_det_thresh_cnt_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value),
				.uhsif_lock_det_thresh_diff_after_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value),
				.uhsif_lock_det_thresh_diff_before_lock_value(hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value)
			) inst_twentynm_hssi_tx_pcs_pma_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pcs_pma_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pcs_pma_interface_blockselect),
				.int_pmaif_10g_tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
				.int_pmaif_8g_txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
				.int_pmaif_pldif_tx_clkdiv(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pmaif_pldif_tx_clkdiv_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pmaif_pldif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
				.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
				.int_pmaif_pldif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.int_tx_dft_obsrv_clk(w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk),
				.pma_tx_elec_idle(w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle),
				.pma_tx_pma_data(w_hssi_tx_pcs_pma_interface_pma_tx_pma_data),
				.pma_txpma_rstb(w_hssi_tx_pcs_pma_interface_pma_txpma_rstb),
				.tx_pma_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback),
				.tx_pma_uhsif_data_loopback(w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback),
				.tx_prbs_gen_test(w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test),
				.uhsif_test_out_1(w_hssi_tx_pcs_pma_interface_uhsif_test_out_1),
				.uhsif_test_out_2(w_hssi_tx_pcs_pma_interface_uhsif_test_out_2),
				.uhsif_test_out_3(w_hssi_tx_pcs_pma_interface_uhsif_test_out_3),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.int_pmaif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
				.int_pmaif_10g_tx_pma_data({w_hssi_10g_tx_pcs_tx_pma_data[63], w_hssi_10g_tx_pcs_tx_pma_data[62], w_hssi_10g_tx_pcs_tx_pma_data[61], w_hssi_10g_tx_pcs_tx_pma_data[60], w_hssi_10g_tx_pcs_tx_pma_data[59], w_hssi_10g_tx_pcs_tx_pma_data[58], w_hssi_10g_tx_pcs_tx_pma_data[57], w_hssi_10g_tx_pcs_tx_pma_data[56], w_hssi_10g_tx_pcs_tx_pma_data[55], w_hssi_10g_tx_pcs_tx_pma_data[54], w_hssi_10g_tx_pcs_tx_pma_data[53], w_hssi_10g_tx_pcs_tx_pma_data[52], w_hssi_10g_tx_pcs_tx_pma_data[51], w_hssi_10g_tx_pcs_tx_pma_data[50], w_hssi_10g_tx_pcs_tx_pma_data[49], w_hssi_10g_tx_pcs_tx_pma_data[48], w_hssi_10g_tx_pcs_tx_pma_data[47], w_hssi_10g_tx_pcs_tx_pma_data[46], w_hssi_10g_tx_pcs_tx_pma_data[45], w_hssi_10g_tx_pcs_tx_pma_data[44], w_hssi_10g_tx_pcs_tx_pma_data[43], w_hssi_10g_tx_pcs_tx_pma_data[42], w_hssi_10g_tx_pcs_tx_pma_data[41], w_hssi_10g_tx_pcs_tx_pma_data[40], w_hssi_10g_tx_pcs_tx_pma_data[39], w_hssi_10g_tx_pcs_tx_pma_data[38], w_hssi_10g_tx_pcs_tx_pma_data[37], w_hssi_10g_tx_pcs_tx_pma_data[36], w_hssi_10g_tx_pcs_tx_pma_data[35], w_hssi_10g_tx_pcs_tx_pma_data[34], w_hssi_10g_tx_pcs_tx_pma_data[33], w_hssi_10g_tx_pcs_tx_pma_data[32], w_hssi_10g_tx_pcs_tx_pma_data[31], w_hssi_10g_tx_pcs_tx_pma_data[30], w_hssi_10g_tx_pcs_tx_pma_data[29], w_hssi_10g_tx_pcs_tx_pma_data[28], w_hssi_10g_tx_pcs_tx_pma_data[27], w_hssi_10g_tx_pcs_tx_pma_data[26], w_hssi_10g_tx_pcs_tx_pma_data[25], w_hssi_10g_tx_pcs_tx_pma_data[24], w_hssi_10g_tx_pcs_tx_pma_data[23], w_hssi_10g_tx_pcs_tx_pma_data[22], w_hssi_10g_tx_pcs_tx_pma_data[21], w_hssi_10g_tx_pcs_tx_pma_data[20], w_hssi_10g_tx_pcs_tx_pma_data[19], w_hssi_10g_tx_pcs_tx_pma_data[18], w_hssi_10g_tx_pcs_tx_pma_data[17], w_hssi_10g_tx_pcs_tx_pma_data[16], w_hssi_10g_tx_pcs_tx_pma_data[15], w_hssi_10g_tx_pcs_tx_pma_data[14], w_hssi_10g_tx_pcs_tx_pma_data[13], w_hssi_10g_tx_pcs_tx_pma_data[12], w_hssi_10g_tx_pcs_tx_pma_data[11], w_hssi_10g_tx_pcs_tx_pma_data[10], w_hssi_10g_tx_pcs_tx_pma_data[9], w_hssi_10g_tx_pcs_tx_pma_data[8], w_hssi_10g_tx_pcs_tx_pma_data[7], w_hssi_10g_tx_pcs_tx_pma_data[6], w_hssi_10g_tx_pcs_tx_pma_data[5], w_hssi_10g_tx_pcs_tx_pma_data[4], w_hssi_10g_tx_pcs_tx_pma_data[3], w_hssi_10g_tx_pcs_tx_pma_data[2], w_hssi_10g_tx_pcs_tx_pma_data[1], w_hssi_10g_tx_pcs_tx_pma_data[0]}),
				.int_pmaif_10g_tx_pma_data_gate_val({w_hssi_10g_tx_pcs_tx_pma_gating_val[63], w_hssi_10g_tx_pcs_tx_pma_gating_val[62], w_hssi_10g_tx_pcs_tx_pma_gating_val[61], w_hssi_10g_tx_pcs_tx_pma_gating_val[60], w_hssi_10g_tx_pcs_tx_pma_gating_val[59], w_hssi_10g_tx_pcs_tx_pma_gating_val[58], w_hssi_10g_tx_pcs_tx_pma_gating_val[57], w_hssi_10g_tx_pcs_tx_pma_gating_val[56], w_hssi_10g_tx_pcs_tx_pma_gating_val[55], w_hssi_10g_tx_pcs_tx_pma_gating_val[54], w_hssi_10g_tx_pcs_tx_pma_gating_val[53], w_hssi_10g_tx_pcs_tx_pma_gating_val[52], w_hssi_10g_tx_pcs_tx_pma_gating_val[51], w_hssi_10g_tx_pcs_tx_pma_gating_val[50], w_hssi_10g_tx_pcs_tx_pma_gating_val[49], w_hssi_10g_tx_pcs_tx_pma_gating_val[48], w_hssi_10g_tx_pcs_tx_pma_gating_val[47], w_hssi_10g_tx_pcs_tx_pma_gating_val[46], w_hssi_10g_tx_pcs_tx_pma_gating_val[45], w_hssi_10g_tx_pcs_tx_pma_gating_val[44], w_hssi_10g_tx_pcs_tx_pma_gating_val[43], w_hssi_10g_tx_pcs_tx_pma_gating_val[42], w_hssi_10g_tx_pcs_tx_pma_gating_val[41], w_hssi_10g_tx_pcs_tx_pma_gating_val[40], w_hssi_10g_tx_pcs_tx_pma_gating_val[39], w_hssi_10g_tx_pcs_tx_pma_gating_val[38], w_hssi_10g_tx_pcs_tx_pma_gating_val[37], w_hssi_10g_tx_pcs_tx_pma_gating_val[36], w_hssi_10g_tx_pcs_tx_pma_gating_val[35], w_hssi_10g_tx_pcs_tx_pma_gating_val[34], w_hssi_10g_tx_pcs_tx_pma_gating_val[33], w_hssi_10g_tx_pcs_tx_pma_gating_val[32], w_hssi_10g_tx_pcs_tx_pma_gating_val[31], w_hssi_10g_tx_pcs_tx_pma_gating_val[30], w_hssi_10g_tx_pcs_tx_pma_gating_val[29], w_hssi_10g_tx_pcs_tx_pma_gating_val[28], w_hssi_10g_tx_pcs_tx_pma_gating_val[27], w_hssi_10g_tx_pcs_tx_pma_gating_val[26], w_hssi_10g_tx_pcs_tx_pma_gating_val[25], w_hssi_10g_tx_pcs_tx_pma_gating_val[24], w_hssi_10g_tx_pcs_tx_pma_gating_val[23], w_hssi_10g_tx_pcs_tx_pma_gating_val[22], w_hssi_10g_tx_pcs_tx_pma_gating_val[21], w_hssi_10g_tx_pcs_tx_pma_gating_val[20], w_hssi_10g_tx_pcs_tx_pma_gating_val[19], w_hssi_10g_tx_pcs_tx_pma_gating_val[18], w_hssi_10g_tx_pcs_tx_pma_gating_val[17], w_hssi_10g_tx_pcs_tx_pma_gating_val[16], w_hssi_10g_tx_pcs_tx_pma_gating_val[15], w_hssi_10g_tx_pcs_tx_pma_gating_val[14], w_hssi_10g_tx_pcs_tx_pma_gating_val[13], w_hssi_10g_tx_pcs_tx_pma_gating_val[12], w_hssi_10g_tx_pcs_tx_pma_gating_val[11], w_hssi_10g_tx_pcs_tx_pma_gating_val[10], w_hssi_10g_tx_pcs_tx_pma_gating_val[9], w_hssi_10g_tx_pcs_tx_pma_gating_val[8], w_hssi_10g_tx_pcs_tx_pma_gating_val[7], w_hssi_10g_tx_pcs_tx_pma_gating_val[6], w_hssi_10g_tx_pcs_tx_pma_gating_val[5], w_hssi_10g_tx_pcs_tx_pma_gating_val[4], w_hssi_10g_tx_pcs_tx_pma_gating_val[3], w_hssi_10g_tx_pcs_tx_pma_gating_val[2], w_hssi_10g_tx_pcs_tx_pma_gating_val[1], w_hssi_10g_tx_pcs_tx_pma_gating_val[0]}),
				.int_pmaif_8g_pudr({w_hssi_8g_tx_pcs_dataout[19], w_hssi_8g_tx_pcs_dataout[18], w_hssi_8g_tx_pcs_dataout[17], w_hssi_8g_tx_pcs_dataout[16], w_hssi_8g_tx_pcs_dataout[15], w_hssi_8g_tx_pcs_dataout[14], w_hssi_8g_tx_pcs_dataout[13], w_hssi_8g_tx_pcs_dataout[12], w_hssi_8g_tx_pcs_dataout[11], w_hssi_8g_tx_pcs_dataout[10], w_hssi_8g_tx_pcs_dataout[9], w_hssi_8g_tx_pcs_dataout[8], w_hssi_8g_tx_pcs_dataout[7], w_hssi_8g_tx_pcs_dataout[6], w_hssi_8g_tx_pcs_dataout[5], w_hssi_8g_tx_pcs_dataout[4], w_hssi_8g_tx_pcs_dataout[3], w_hssi_8g_tx_pcs_dataout[2], w_hssi_8g_tx_pcs_dataout[1], w_hssi_8g_tx_pcs_dataout[0]}),
				.int_pmaif_8g_tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
				.int_pmaif_8g_tx_elec_idle(w_hssi_pipe_gen1_2_tx_elec_idle_out),
				.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
				.int_pmaif_g3_pma_data_out({w_hssi_gen3_tx_pcs_data_out[31], w_hssi_gen3_tx_pcs_data_out[30], w_hssi_gen3_tx_pcs_data_out[29], w_hssi_gen3_tx_pcs_data_out[28], w_hssi_gen3_tx_pcs_data_out[27], w_hssi_gen3_tx_pcs_data_out[26], w_hssi_gen3_tx_pcs_data_out[25], w_hssi_gen3_tx_pcs_data_out[24], w_hssi_gen3_tx_pcs_data_out[23], w_hssi_gen3_tx_pcs_data_out[22], w_hssi_gen3_tx_pcs_data_out[21], w_hssi_gen3_tx_pcs_data_out[20], w_hssi_gen3_tx_pcs_data_out[19], w_hssi_gen3_tx_pcs_data_out[18], w_hssi_gen3_tx_pcs_data_out[17], w_hssi_gen3_tx_pcs_data_out[16], w_hssi_gen3_tx_pcs_data_out[15], w_hssi_gen3_tx_pcs_data_out[14], w_hssi_gen3_tx_pcs_data_out[13], w_hssi_gen3_tx_pcs_data_out[12], w_hssi_gen3_tx_pcs_data_out[11], w_hssi_gen3_tx_pcs_data_out[10], w_hssi_gen3_tx_pcs_data_out[9], w_hssi_gen3_tx_pcs_data_out[8], w_hssi_gen3_tx_pcs_data_out[7], w_hssi_gen3_tx_pcs_data_out[6], w_hssi_gen3_tx_pcs_data_out[5], w_hssi_gen3_tx_pcs_data_out[4], w_hssi_gen3_tx_pcs_data_out[3], w_hssi_gen3_tx_pcs_data_out[2], w_hssi_gen3_tx_pcs_data_out[1], w_hssi_gen3_tx_pcs_data_out[0]}),
				.int_pmaif_g3_pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
				.int_pmaif_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pmaif_pldif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pmaif_pldif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0]}),
				.int_pmaif_pldif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pmaif_pldif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
				.int_pmaif_pldif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pmaif_pldif_uhsif_tx_data({w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1], w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0]}),
				.pma_tx_clkdiv_user(in_pma_tx_clkdiv_user),
				.pma_tx_pma_clk(in_pma_tx_pma_clk),
				.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
				.refclk_dig_uhsif(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
				.uhsif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
				.uhsif_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
				
				// UNUSED
				.avmm_user_dataout(),
				.write_en(),
				.write_en_ack()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pcs_pma_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pcs_pma_interface_blockselect = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4:0] = 5'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_pma_txpma_rstb = 1'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63:0] = 64'b0;
				assign w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19:0] = 20'b0;
				assign w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19:0] = 20'b0;
		end // if not generate
		
		// instantiating twentynm_hssi_tx_pld_pcs_interface
		if ((xcvr_native_mode == "mode_tx_only") || (xcvr_native_mode == "mode_duplex")) begin:gen_twentynm_hssi_tx_pld_pcs_interface
			twentynm_hssi_tx_pld_pcs_interface #(
				.hd_10g_advanced_user_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx),
				.hd_10g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode),
				.hd_10g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_10g_ctrl_plane_bonding_tx),
				.hd_10g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx),
				.hd_10g_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx),
				.hd_10g_lpbk_en(hssi_tx_pld_pcs_interface_hd_10g_lpbk_en),
				.hd_10g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx),
				.hd_10g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx),
				.hd_10g_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx),
				.hd_8g_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode),
				.hd_8g_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_8g_ctrl_plane_bonding_tx),
				.hd_8g_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx),
				.hd_8g_hip_mode(hssi_tx_pld_pcs_interface_hd_8g_hip_mode),
				.hd_8g_lpbk_en(hssi_tx_pld_pcs_interface_hd_8g_lpbk_en),
				.hd_8g_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx),
				.hd_8g_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx),
				.hd_chnl_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode),
				.hd_chnl_ctrl_plane_bonding_tx(hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx),
				.hd_chnl_frequency_rules_en(hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en),
				.hd_chnl_func_mode(hssi_tx_pld_pcs_interface_hd_chnl_func_mode),
				.hd_chnl_hip_en(hssi_tx_pld_pcs_interface_hd_chnl_hip_en),
				.hd_chnl_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en),
				.hd_chnl_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx),
				.hd_chnl_lpbk_en(hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en),
				.hd_chnl_pld_fifo_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx),
				.hd_chnl_pld_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz),
				.hd_chnl_pld_uhsif_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz),
				.hd_chnl_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx),
				.hd_chnl_pma_tx_clk_hz(hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz),
				.hd_chnl_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx),
				.hd_chnl_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx),
				.hd_fifo_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode),
				.hd_fifo_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx),
				.hd_fifo_shared_fifo_width_tx(hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx),
				.hd_g3_prot_mode(hssi_tx_pld_pcs_interface_hd_g3_prot_mode),
				.hd_krfec_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode),
				.hd_krfec_low_latency_en_tx(hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx),
				.hd_krfec_lpbk_en(hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en),
				.hd_krfec_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx),
				.hd_pldif_hrdrstctl_en(hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en),
				.hd_pldif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx),
				.hd_pmaif_channel_operation_mode(hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode),
				.hd_pmaif_ctrl_plane_bonding(hssi_tx_pld_pcs_interface_hd_pmaif_ctrl_plane_bonding),
				.hd_pmaif_lpbk_en(hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en),
				.hd_pmaif_pma_dw_tx(hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx),
				.hd_pmaif_prot_mode_tx(hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx),
				.hd_pmaif_sim_mode(hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode),
				.pcs_tx_clk_out_sel(hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel),
				.pcs_tx_clk_source(hssi_tx_pld_pcs_interface_pcs_tx_clk_source),
				.pcs_tx_data_source(hssi_tx_pld_pcs_interface_pcs_tx_data_source),
				.pcs_tx_delay1_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en),
				.pcs_tx_delay1_clk_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel),
				.pcs_tx_delay1_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl),
				.pcs_tx_delay1_data_sel(hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel),
				.pcs_tx_delay2_clk_en(hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en),
				.pcs_tx_delay2_ctrl(hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl),
				.pcs_tx_output_sel(hssi_tx_pld_pcs_interface_pcs_tx_output_sel),
				.reconfig_settings(hssi_tx_pld_pcs_interface_reconfig_settings),
				.silicon_rev( "20nm4es" )       //PARAM_HIDE
			) inst_twentynm_hssi_tx_pld_pcs_interface (
				// OUTPUTS
				.avmmreaddata(w_hssi_tx_pld_pcs_interface_avmmreaddata),
				.blockselect(w_hssi_tx_pld_pcs_interface_blockselect),
				.hip_tx_clk(w_hssi_tx_pld_pcs_interface_hip_tx_clk),
				.int_pldif_10g_tx_bitslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip),
				.int_pldif_10g_tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
				.int_pldif_10g_tx_control(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control),
				.int_pldif_10g_tx_control_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg),
				.int_pldif_10g_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data),
				.int_pldif_10g_tx_data_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg),
				.int_pldif_10g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
				.int_pldif_10g_tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
				.int_pldif_10g_tx_diag_status(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status),
				.int_pldif_10g_tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
				.int_pldif_10g_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
				.int_pldif_10g_tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
				.int_pldif_8g_pld_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
				.int_pldif_8g_powerdown(w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown),
				.int_pldif_8g_rddisable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
				.int_pldif_8g_rev_loopbk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
				.int_pldif_8g_tx_blk_start(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start),
				.int_pldif_8g_tx_boundary_sel(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel),
				.int_pldif_8g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid),
				.int_pldif_8g_tx_sync_hdr(w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr),
				.int_pldif_8g_txd(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd),
				.int_pldif_8g_txd_fast_reg(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg),
				.int_pldif_8g_txdeemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
				.int_pldif_8g_txdetectrxloopback(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
				.int_pldif_8g_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
				.int_pldif_8g_txmargin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin),
				.int_pldif_8g_txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
				.int_pldif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
				.int_pldif_8g_wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
				.int_pldif_pmaif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
				.int_pldif_pmaif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
				.int_pldif_pmaif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data),
				.int_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
				.int_pldif_pmaif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
				.int_pldif_pmaif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
				.int_pldif_pmaif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
				.int_pldif_pmaif_uhsif_tx_data(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data),
				.pld_10g_krfec_tx_frame(w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame),
				.pld_10g_tx_burst_en_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe),
				.pld_10g_tx_empty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty),
				.pld_10g_tx_fifo_num(w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num),
				.pld_10g_tx_full(w_hssi_tx_pld_pcs_interface_pld_10g_tx_full),
				.pld_10g_tx_pempty(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty),
				.pld_10g_tx_pfull(w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull),
				.pld_10g_tx_wordslip_exe(w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe),
				.pld_8g_empty_tx(w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx),
				.pld_8g_full_tx(w_hssi_tx_pld_pcs_interface_pld_8g_full_tx),
				.pld_krfec_tx_alignment(w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment),
				.pld_pcs_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out),
				.pld_pma_clkdiv_tx_user(w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user),
				.pld_pma_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out),
				.pld_uhsif_tx_clk_out(w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out),
				// INPUTS
				.avmmaddress({in_avmmaddress[8], in_avmmaddress[7], in_avmmaddress[6], in_avmmaddress[5], in_avmmaddress[4], in_avmmaddress[3], in_avmmaddress[2], in_avmmaddress[1], in_avmmaddress[0]}),
				.avmmclk(in_avmmclk),
				.avmmread(in_avmmread),
				.avmmrstn(in_avmmrstn),
				.avmmwrite(in_avmmwrite),
				.avmmwritedata({in_avmmwritedata[7], in_avmmwritedata[6], in_avmmwritedata[5], in_avmmwritedata[4], in_avmmwritedata[3], in_avmmwritedata[2], in_avmmwritedata[1], in_avmmwritedata[0]}),
				.hip_tx_data({in_hip_tx_data[63], in_hip_tx_data[62], in_hip_tx_data[61], in_hip_tx_data[60], in_hip_tx_data[59], in_hip_tx_data[58], in_hip_tx_data[57], in_hip_tx_data[56], in_hip_tx_data[55], in_hip_tx_data[54], in_hip_tx_data[53], in_hip_tx_data[52], in_hip_tx_data[51], in_hip_tx_data[50], in_hip_tx_data[49], in_hip_tx_data[48], in_hip_tx_data[47], in_hip_tx_data[46], in_hip_tx_data[45], in_hip_tx_data[44], in_hip_tx_data[43], in_hip_tx_data[42], in_hip_tx_data[41], in_hip_tx_data[40], in_hip_tx_data[39], in_hip_tx_data[38], in_hip_tx_data[37], in_hip_tx_data[36], in_hip_tx_data[35], in_hip_tx_data[34], in_hip_tx_data[33], in_hip_tx_data[32], in_hip_tx_data[31], in_hip_tx_data[30], in_hip_tx_data[29], in_hip_tx_data[28], in_hip_tx_data[27], in_hip_tx_data[26], in_hip_tx_data[25], in_hip_tx_data[24], in_hip_tx_data[23], in_hip_tx_data[22], in_hip_tx_data[21], in_hip_tx_data[20], in_hip_tx_data[19], in_hip_tx_data[18], in_hip_tx_data[17], in_hip_tx_data[16], in_hip_tx_data[15], in_hip_tx_data[14], in_hip_tx_data[13], in_hip_tx_data[12], in_hip_tx_data[11], in_hip_tx_data[10], in_hip_tx_data[9], in_hip_tx_data[8], in_hip_tx_data[7], in_hip_tx_data[6], in_hip_tx_data[5], in_hip_tx_data[4], in_hip_tx_data[3], in_hip_tx_data[2], in_hip_tx_data[1], in_hip_tx_data[0]}),
				.int_pldif_10g_tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
				.int_pldif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
				.int_pldif_10g_tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_10g_tx_empty(w_hssi_10g_tx_pcs_tx_empty),
				.int_pldif_10g_tx_fifo_num({w_hssi_10g_tx_pcs_tx_fifo_num[3], w_hssi_10g_tx_pcs_tx_fifo_num[2], w_hssi_10g_tx_pcs_tx_fifo_num[1], w_hssi_10g_tx_pcs_tx_fifo_num[0]}),
				.int_pldif_10g_tx_frame(w_hssi_10g_tx_pcs_tx_frame),
				.int_pldif_10g_tx_full(w_hssi_10g_tx_pcs_tx_full),
				.int_pldif_10g_tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
				.int_pldif_10g_tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
				.int_pldif_10g_tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
				.int_pldif_8g_empty_tx(w_hssi_8g_tx_pcs_ph_fifo_underflow),
				.int_pldif_8g_full_tx(w_hssi_8g_tx_pcs_ph_fifo_overflow),
				.int_pldif_8g_tx_clk_out(w_hssi_8g_tx_pcs_clk_out),
				.int_pldif_8g_tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
				.int_pldif_krfec_tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
				.int_pldif_krfec_tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
				.int_pldif_pmaif_clkdiv_tx(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
				.int_pldif_pmaif_clkdiv_tx_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
				.int_pldif_pmaif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
				.pld_10g_krfec_tx_pld_rst_n(in_pld_10g_krfec_tx_pld_rst_n),
				.pld_10g_tx_bitslip({in_pld_10g_tx_bitslip[6], in_pld_10g_tx_bitslip[5], in_pld_10g_tx_bitslip[4], in_pld_10g_tx_bitslip[3], in_pld_10g_tx_bitslip[2], in_pld_10g_tx_bitslip[1], in_pld_10g_tx_bitslip[0]}),
				.pld_10g_tx_burst_en(in_pld_10g_tx_burst_en),
				.pld_10g_tx_data_valid(in_pld_10g_tx_data_valid),
				.pld_10g_tx_diag_status({in_pld_10g_tx_diag_status[1], in_pld_10g_tx_diag_status[0]}),
				.pld_10g_tx_wordslip(in_pld_10g_tx_wordslip),
				.pld_8g_g3_tx_pld_rst_n(in_pld_8g_g3_tx_pld_rst_n),
				.pld_8g_rddisable_tx(in_pld_8g_rddisable_tx),
				.pld_8g_tx_boundary_sel({in_pld_8g_tx_boundary_sel[4], in_pld_8g_tx_boundary_sel[3], in_pld_8g_tx_boundary_sel[2], in_pld_8g_tx_boundary_sel[1], in_pld_8g_tx_boundary_sel[0]}),
				.pld_8g_wrenable_tx(in_pld_8g_wrenable_tx),
				.pld_partial_reconfig(in_pld_partial_reconfig),
				.pld_pma_txpma_rstb(in_pld_pma_txpma_rstb),
				.pld_pmaif_tx_pld_rst_n(in_pld_pmaif_tx_pld_rst_n),
				.pld_polinv_tx(in_pld_polinv_tx),
				.pld_tx_clk(in_pld_tx_clk),
				.pld_tx_control({in_pld_tx_control[17], in_pld_tx_control[16], in_pld_tx_control[15], in_pld_tx_control[14], in_pld_tx_control[13], in_pld_tx_control[12], in_pld_tx_control[11], in_pld_tx_control[10], in_pld_tx_control[9], in_pld_tx_control[8], in_pld_tx_control[7], in_pld_tx_control[6], in_pld_tx_control[5], in_pld_tx_control[4], in_pld_tx_control[3], in_pld_tx_control[2], in_pld_tx_control[1], in_pld_tx_control[0]}),
				.pld_tx_data({in_pld_tx_data[127], in_pld_tx_data[126], in_pld_tx_data[125], in_pld_tx_data[124], in_pld_tx_data[123], in_pld_tx_data[122], in_pld_tx_data[121], in_pld_tx_data[120], in_pld_tx_data[119], in_pld_tx_data[118], in_pld_tx_data[117], in_pld_tx_data[116], in_pld_tx_data[115], in_pld_tx_data[114], in_pld_tx_data[113], in_pld_tx_data[112], in_pld_tx_data[111], in_pld_tx_data[110], in_pld_tx_data[109], in_pld_tx_data[108], in_pld_tx_data[107], in_pld_tx_data[106], in_pld_tx_data[105], in_pld_tx_data[104], in_pld_tx_data[103], in_pld_tx_data[102], in_pld_tx_data[101], in_pld_tx_data[100], in_pld_tx_data[99], in_pld_tx_data[98], in_pld_tx_data[97], in_pld_tx_data[96], in_pld_tx_data[95], in_pld_tx_data[94], in_pld_tx_data[93], in_pld_tx_data[92], in_pld_tx_data[91], in_pld_tx_data[90], in_pld_tx_data[89], in_pld_tx_data[88], in_pld_tx_data[87], in_pld_tx_data[86], in_pld_tx_data[85], in_pld_tx_data[84], in_pld_tx_data[83], in_pld_tx_data[82], in_pld_tx_data[81], in_pld_tx_data[80], in_pld_tx_data[79], in_pld_tx_data[78], in_pld_tx_data[77], in_pld_tx_data[76], in_pld_tx_data[75], in_pld_tx_data[74], in_pld_tx_data[73], in_pld_tx_data[72], in_pld_tx_data[71], in_pld_tx_data[70], in_pld_tx_data[69], in_pld_tx_data[68], in_pld_tx_data[67], in_pld_tx_data[66], in_pld_tx_data[65], in_pld_tx_data[64], in_pld_tx_data[63], in_pld_tx_data[62], in_pld_tx_data[61], in_pld_tx_data[60], in_pld_tx_data[59], in_pld_tx_data[58], in_pld_tx_data[57], in_pld_tx_data[56], in_pld_tx_data[55], in_pld_tx_data[54], in_pld_tx_data[53], in_pld_tx_data[52], in_pld_tx_data[51], in_pld_tx_data[50], in_pld_tx_data[49], in_pld_tx_data[48], in_pld_tx_data[47], in_pld_tx_data[46], in_pld_tx_data[45], in_pld_tx_data[44], in_pld_tx_data[43], in_pld_tx_data[42], in_pld_tx_data[41], in_pld_tx_data[40], in_pld_tx_data[39], in_pld_tx_data[38], in_pld_tx_data[37], in_pld_tx_data[36], in_pld_tx_data[35], in_pld_tx_data[34], in_pld_tx_data[33], in_pld_tx_data[32], in_pld_tx_data[31], in_pld_tx_data[30], in_pld_tx_data[29], in_pld_tx_data[28], in_pld_tx_data[27], in_pld_tx_data[26], in_pld_tx_data[25], in_pld_tx_data[24], in_pld_tx_data[23], in_pld_tx_data[22], in_pld_tx_data[21], in_pld_tx_data[20], in_pld_tx_data[19], in_pld_tx_data[18], in_pld_tx_data[17], in_pld_tx_data[16], in_pld_tx_data[15], in_pld_tx_data[14], in_pld_tx_data[13], in_pld_tx_data[12], in_pld_tx_data[11], in_pld_tx_data[10], in_pld_tx_data[9], in_pld_tx_data[8], in_pld_tx_data[7], in_pld_tx_data[6], in_pld_tx_data[5], in_pld_tx_data[4], in_pld_tx_data[3], in_pld_tx_data[2], in_pld_tx_data[1], in_pld_tx_data[0]}),
				.pld_txelecidle(in_pld_txelecidle),
				.pld_uhsif_tx_clk(in_pld_uhsif_tx_clk),
				.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
				
				// UNUSED
				.hip_clk_out_div_by_2_wire(),
				.hip_clk_out_wire(),
				.int_pldif_pmaif_tx_pld_clk(),
				.pld_10g_tx_burst_en_exe_10g_fastreg(),
				.pld_10g_tx_burst_en_exe_plddirect_reg(),
				.pld_10g_tx_data_valid_2ff_delay1_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay3_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_fastreg(),
				.pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg(),
				.pld_10g_tx_data_valid_fastreg(),
				.pld_10g_tx_data_valid_plddirect_fastreg(),
				.pld_pcs_tx_clk_out_pma_wire(),
				.pld_pma_tx_clk_out_wire(),
				.pld_pmaif_tx_pld_rst_n_reg(),
				.pld_polinv_tx_10g_pcsdirect_reg(),
				.pld_polinv_tx_8g_reg(),
				.pld_polinv_tx_pat_reg(),
				.pld_tx_clk_fifo(),
				.pld_tx_control_fifo(),
				.pld_tx_control_hi_10g_reg(),
				.pld_tx_control_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_10g_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_control_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_control_lo_8g_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_control_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_control_lo_plddirect_fastreg(),
				.pld_tx_control_lo_plddirect_reg(),
				.pld_tx_data_hi_reg(),
				.pld_tx_data_lo_10g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_10g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_10g_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay4_fastreg(),
				.pld_tx_data_lo_8g_2ff_delay6_fastreg(),
				.pld_tx_data_lo_8g_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay1_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay3_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay4_fastreg(),
				.pld_tx_data_lo_plddirect_2ff_delay6_fastreg(),
				.pld_tx_data_lo_plddirect_fastreg(),
				.pld_tx_data_lo_plddirect_reg(),
				.pld_uhsif_reg(),
				.pma_tx_pma_clk_reg()
			);
		end // if generate
		else begin
				assign w_hssi_tx_pld_pcs_interface_avmmreaddata[7:0] = 8'b0;
				assign w_hssi_tx_pld_pcs_interface_blockselect = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_hip_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6:0] = 7'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17:0] = 18'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8:0] = 9'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127:0] = 128'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4:0] = 5'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1:0] = 2'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43:0] = 44'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2:0] = 3'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n = 1'b1;		// Override default tieoff
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63:0] = 64'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3:0] = 4'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_full = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_8g_full_tx = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out = 1'b0;
				assign w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out = 1'b0;
		end // if not generate
		
		//output assignments
		assign out_avmmreaddata_hssi_10g_rx_pcs = {w_hssi_10g_rx_pcs_avmmreaddata[7], w_hssi_10g_rx_pcs_avmmreaddata[6], w_hssi_10g_rx_pcs_avmmreaddata[5], w_hssi_10g_rx_pcs_avmmreaddata[4], w_hssi_10g_rx_pcs_avmmreaddata[3], w_hssi_10g_rx_pcs_avmmreaddata[2], w_hssi_10g_rx_pcs_avmmreaddata[1], w_hssi_10g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_10g_tx_pcs = {w_hssi_10g_tx_pcs_avmmreaddata[7], w_hssi_10g_tx_pcs_avmmreaddata[6], w_hssi_10g_tx_pcs_avmmreaddata[5], w_hssi_10g_tx_pcs_avmmreaddata[4], w_hssi_10g_tx_pcs_avmmreaddata[3], w_hssi_10g_tx_pcs_avmmreaddata[2], w_hssi_10g_tx_pcs_avmmreaddata[1], w_hssi_10g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_rx_pcs = {w_hssi_8g_rx_pcs_avmmreaddata[7], w_hssi_8g_rx_pcs_avmmreaddata[6], w_hssi_8g_rx_pcs_avmmreaddata[5], w_hssi_8g_rx_pcs_avmmreaddata[4], w_hssi_8g_rx_pcs_avmmreaddata[3], w_hssi_8g_rx_pcs_avmmreaddata[2], w_hssi_8g_rx_pcs_avmmreaddata[1], w_hssi_8g_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_8g_tx_pcs = {w_hssi_8g_tx_pcs_avmmreaddata[7], w_hssi_8g_tx_pcs_avmmreaddata[6], w_hssi_8g_tx_pcs_avmmreaddata[5], w_hssi_8g_tx_pcs_avmmreaddata[4], w_hssi_8g_tx_pcs_avmmreaddata[3], w_hssi_8g_tx_pcs_avmmreaddata[2], w_hssi_8g_tx_pcs_avmmreaddata[1], w_hssi_8g_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pcs_pma_interface = {w_hssi_common_pcs_pma_interface_avmmreaddata[7], w_hssi_common_pcs_pma_interface_avmmreaddata[6], w_hssi_common_pcs_pma_interface_avmmreaddata[5], w_hssi_common_pcs_pma_interface_avmmreaddata[4], w_hssi_common_pcs_pma_interface_avmmreaddata[3], w_hssi_common_pcs_pma_interface_avmmreaddata[2], w_hssi_common_pcs_pma_interface_avmmreaddata[1], w_hssi_common_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_common_pld_pcs_interface = {w_hssi_common_pld_pcs_interface_avmmreaddata[7], w_hssi_common_pld_pcs_interface_avmmreaddata[6], w_hssi_common_pld_pcs_interface_avmmreaddata[5], w_hssi_common_pld_pcs_interface_avmmreaddata[4], w_hssi_common_pld_pcs_interface_avmmreaddata[3], w_hssi_common_pld_pcs_interface_avmmreaddata[2], w_hssi_common_pld_pcs_interface_avmmreaddata[1], w_hssi_common_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_rx_pcs = {w_hssi_fifo_rx_pcs_avmmreaddata[7], w_hssi_fifo_rx_pcs_avmmreaddata[6], w_hssi_fifo_rx_pcs_avmmreaddata[5], w_hssi_fifo_rx_pcs_avmmreaddata[4], w_hssi_fifo_rx_pcs_avmmreaddata[3], w_hssi_fifo_rx_pcs_avmmreaddata[2], w_hssi_fifo_rx_pcs_avmmreaddata[1], w_hssi_fifo_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_fifo_tx_pcs = {w_hssi_fifo_tx_pcs_avmmreaddata[7], w_hssi_fifo_tx_pcs_avmmreaddata[6], w_hssi_fifo_tx_pcs_avmmreaddata[5], w_hssi_fifo_tx_pcs_avmmreaddata[4], w_hssi_fifo_tx_pcs_avmmreaddata[3], w_hssi_fifo_tx_pcs_avmmreaddata[2], w_hssi_fifo_tx_pcs_avmmreaddata[1], w_hssi_fifo_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_rx_pcs = {w_hssi_gen3_rx_pcs_avmmreaddata[7], w_hssi_gen3_rx_pcs_avmmreaddata[6], w_hssi_gen3_rx_pcs_avmmreaddata[5], w_hssi_gen3_rx_pcs_avmmreaddata[4], w_hssi_gen3_rx_pcs_avmmreaddata[3], w_hssi_gen3_rx_pcs_avmmreaddata[2], w_hssi_gen3_rx_pcs_avmmreaddata[1], w_hssi_gen3_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_gen3_tx_pcs = {w_hssi_gen3_tx_pcs_avmmreaddata[7], w_hssi_gen3_tx_pcs_avmmreaddata[6], w_hssi_gen3_tx_pcs_avmmreaddata[5], w_hssi_gen3_tx_pcs_avmmreaddata[4], w_hssi_gen3_tx_pcs_avmmreaddata[3], w_hssi_gen3_tx_pcs_avmmreaddata[2], w_hssi_gen3_tx_pcs_avmmreaddata[1], w_hssi_gen3_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_rx_pcs = {w_hssi_krfec_rx_pcs_avmmreaddata[7], w_hssi_krfec_rx_pcs_avmmreaddata[6], w_hssi_krfec_rx_pcs_avmmreaddata[5], w_hssi_krfec_rx_pcs_avmmreaddata[4], w_hssi_krfec_rx_pcs_avmmreaddata[3], w_hssi_krfec_rx_pcs_avmmreaddata[2], w_hssi_krfec_rx_pcs_avmmreaddata[1], w_hssi_krfec_rx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_krfec_tx_pcs = {w_hssi_krfec_tx_pcs_avmmreaddata[7], w_hssi_krfec_tx_pcs_avmmreaddata[6], w_hssi_krfec_tx_pcs_avmmreaddata[5], w_hssi_krfec_tx_pcs_avmmreaddata[4], w_hssi_krfec_tx_pcs_avmmreaddata[3], w_hssi_krfec_tx_pcs_avmmreaddata[2], w_hssi_krfec_tx_pcs_avmmreaddata[1], w_hssi_krfec_tx_pcs_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen1_2 = {w_hssi_pipe_gen1_2_avmmreaddata[7], w_hssi_pipe_gen1_2_avmmreaddata[6], w_hssi_pipe_gen1_2_avmmreaddata[5], w_hssi_pipe_gen1_2_avmmreaddata[4], w_hssi_pipe_gen1_2_avmmreaddata[3], w_hssi_pipe_gen1_2_avmmreaddata[2], w_hssi_pipe_gen1_2_avmmreaddata[1], w_hssi_pipe_gen1_2_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_pipe_gen3 = {w_hssi_pipe_gen3_avmmreaddata[7], w_hssi_pipe_gen3_avmmreaddata[6], w_hssi_pipe_gen3_avmmreaddata[5], w_hssi_pipe_gen3_avmmreaddata[4], w_hssi_pipe_gen3_avmmreaddata[3], w_hssi_pipe_gen3_avmmreaddata[2], w_hssi_pipe_gen3_avmmreaddata[1], w_hssi_pipe_gen3_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pcs_pma_interface = {w_hssi_rx_pcs_pma_interface_avmmreaddata[7], w_hssi_rx_pcs_pma_interface_avmmreaddata[6], w_hssi_rx_pcs_pma_interface_avmmreaddata[5], w_hssi_rx_pcs_pma_interface_avmmreaddata[4], w_hssi_rx_pcs_pma_interface_avmmreaddata[3], w_hssi_rx_pcs_pma_interface_avmmreaddata[2], w_hssi_rx_pcs_pma_interface_avmmreaddata[1], w_hssi_rx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_rx_pld_pcs_interface = {w_hssi_rx_pld_pcs_interface_avmmreaddata[7], w_hssi_rx_pld_pcs_interface_avmmreaddata[6], w_hssi_rx_pld_pcs_interface_avmmreaddata[5], w_hssi_rx_pld_pcs_interface_avmmreaddata[4], w_hssi_rx_pld_pcs_interface_avmmreaddata[3], w_hssi_rx_pld_pcs_interface_avmmreaddata[2], w_hssi_rx_pld_pcs_interface_avmmreaddata[1], w_hssi_rx_pld_pcs_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pcs_pma_interface = {w_hssi_tx_pcs_pma_interface_avmmreaddata[7], w_hssi_tx_pcs_pma_interface_avmmreaddata[6], w_hssi_tx_pcs_pma_interface_avmmreaddata[5], w_hssi_tx_pcs_pma_interface_avmmreaddata[4], w_hssi_tx_pcs_pma_interface_avmmreaddata[3], w_hssi_tx_pcs_pma_interface_avmmreaddata[2], w_hssi_tx_pcs_pma_interface_avmmreaddata[1], w_hssi_tx_pcs_pma_interface_avmmreaddata[0]};
		assign out_avmmreaddata_hssi_tx_pld_pcs_interface = {w_hssi_tx_pld_pcs_interface_avmmreaddata[7], w_hssi_tx_pld_pcs_interface_avmmreaddata[6], w_hssi_tx_pld_pcs_interface_avmmreaddata[5], w_hssi_tx_pld_pcs_interface_avmmreaddata[4], w_hssi_tx_pld_pcs_interface_avmmreaddata[3], w_hssi_tx_pld_pcs_interface_avmmreaddata[2], w_hssi_tx_pld_pcs_interface_avmmreaddata[1], w_hssi_tx_pld_pcs_interface_avmmreaddata[0]};
		assign out_blockselect_hssi_10g_rx_pcs = w_hssi_10g_rx_pcs_blockselect;
		assign out_blockselect_hssi_10g_tx_pcs = w_hssi_10g_tx_pcs_blockselect;
		assign out_blockselect_hssi_8g_rx_pcs = w_hssi_8g_rx_pcs_blockselect;
		assign out_blockselect_hssi_8g_tx_pcs = w_hssi_8g_tx_pcs_blockselect;
		assign out_blockselect_hssi_common_pcs_pma_interface = w_hssi_common_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_common_pld_pcs_interface = w_hssi_common_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_fifo_rx_pcs = w_hssi_fifo_rx_pcs_blockselect;
		assign out_blockselect_hssi_fifo_tx_pcs = w_hssi_fifo_tx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_rx_pcs = w_hssi_gen3_rx_pcs_blockselect;
		assign out_blockselect_hssi_gen3_tx_pcs = w_hssi_gen3_tx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_rx_pcs = w_hssi_krfec_rx_pcs_blockselect;
		assign out_blockselect_hssi_krfec_tx_pcs = w_hssi_krfec_tx_pcs_blockselect;
		assign out_blockselect_hssi_pipe_gen1_2 = w_hssi_pipe_gen1_2_blockselect;
		assign out_blockselect_hssi_pipe_gen3 = w_hssi_pipe_gen3_blockselect;
		assign out_blockselect_hssi_rx_pcs_pma_interface = w_hssi_rx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_rx_pld_pcs_interface = w_hssi_rx_pld_pcs_interface_blockselect;
		assign out_blockselect_hssi_tx_pcs_pma_interface = w_hssi_tx_pcs_pma_interface_blockselect;
		assign out_blockselect_hssi_tx_pld_pcs_interface = w_hssi_tx_pld_pcs_interface_blockselect;
		assign out_bond_pcs10g_out_bot = {w_hssi_10g_tx_pcs_distdwn_out_rden, w_hssi_10g_tx_pcs_distdwn_out_wren, w_hssi_10g_tx_pcs_distdwn_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs10g_out_top = {w_hssi_10g_tx_pcs_distup_out_rden, w_hssi_10g_tx_pcs_distup_out_wren, w_hssi_10g_tx_pcs_distup_out_dv, 1'b0, 1'b0};
		assign out_bond_pcs8g_out_bot = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_down, w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_down[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_down, w_hssi_8g_tx_pcs_wr_enable_out_chnl_down, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_down[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_down[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_down, w_hssi_8g_rx_pcs_wr_enable_out_chnl_down, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_down[0]};
		assign out_bond_pcs8g_out_top = {w_hssi_8g_rx_pcs_reset_pc_ptrs_out_chnl_up, w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[1], w_hssi_8g_tx_pcs_fifo_select_out_chnl_up[0], w_hssi_8g_tx_pcs_rd_enable_out_chnl_up, w_hssi_8g_tx_pcs_wr_enable_out_chnl_up, w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[1], w_hssi_8g_tx_pcs_tx_div_sync_out_chnl_up[0], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_we_out_chnl_up[0], w_hssi_8g_rx_pcs_rd_enable_out_chnl_up, w_hssi_8g_rx_pcs_wr_enable_out_chnl_up, w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[1], w_hssi_8g_rx_pcs_rx_div_sync_out_chnl_up[0]};
		assign out_bond_pmaif_out_bot = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_down[0]};
		assign out_bond_pmaif_out_top = {w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[11], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[10], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[9], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[8], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[7], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[6], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[5], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[4], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[3], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[2], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[1], w_hssi_common_pcs_pma_interface_pmaif_bundling_out_up[0]};
		assign out_hip_clk_out = {w_hssi_common_pld_pcs_interface_hip_cmn_clk[1], w_hssi_common_pld_pcs_interface_hip_cmn_clk[0], w_hssi_tx_pld_pcs_interface_hip_tx_clk};
		assign out_hip_ctrl_out = {w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[5], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[4], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[3], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[2], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[1], w_hssi_common_pld_pcs_interface_hip_cmn_ctrl[0], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[1], w_hssi_rx_pld_pcs_interface_hip_rx_ctrl[0]};
		assign out_hip_iocsr_rdy = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy;
		assign out_hip_iocsr_rdy_dly = w_hssi_common_pld_pcs_interface_hip_iocsr_rdy_dly;
		assign out_hip_nfrzdrv = w_hssi_common_pld_pcs_interface_hip_nfrzdrv;
		assign out_hip_npor = w_hssi_common_pld_pcs_interface_hip_npor;
		assign out_hip_rx_data = {w_hssi_rx_pld_pcs_interface_hip_rx_data[50], w_hssi_rx_pld_pcs_interface_hip_rx_data[49], w_hssi_rx_pld_pcs_interface_hip_rx_data[48], w_hssi_rx_pld_pcs_interface_hip_rx_data[47], w_hssi_rx_pld_pcs_interface_hip_rx_data[46], w_hssi_rx_pld_pcs_interface_hip_rx_data[45], w_hssi_rx_pld_pcs_interface_hip_rx_data[44], w_hssi_rx_pld_pcs_interface_hip_rx_data[43], w_hssi_rx_pld_pcs_interface_hip_rx_data[42], w_hssi_rx_pld_pcs_interface_hip_rx_data[41], w_hssi_rx_pld_pcs_interface_hip_rx_data[40], w_hssi_rx_pld_pcs_interface_hip_rx_data[39], w_hssi_rx_pld_pcs_interface_hip_rx_data[38], w_hssi_rx_pld_pcs_interface_hip_rx_data[37], w_hssi_rx_pld_pcs_interface_hip_rx_data[36], w_hssi_rx_pld_pcs_interface_hip_rx_data[35], w_hssi_rx_pld_pcs_interface_hip_rx_data[34], w_hssi_rx_pld_pcs_interface_hip_rx_data[33], w_hssi_rx_pld_pcs_interface_hip_rx_data[32], w_hssi_rx_pld_pcs_interface_hip_rx_data[31], w_hssi_rx_pld_pcs_interface_hip_rx_data[30], w_hssi_rx_pld_pcs_interface_hip_rx_data[29], w_hssi_rx_pld_pcs_interface_hip_rx_data[28], w_hssi_rx_pld_pcs_interface_hip_rx_data[27], w_hssi_rx_pld_pcs_interface_hip_rx_data[26], w_hssi_rx_pld_pcs_interface_hip_rx_data[25], w_hssi_rx_pld_pcs_interface_hip_rx_data[24], w_hssi_rx_pld_pcs_interface_hip_rx_data[23], w_hssi_rx_pld_pcs_interface_hip_rx_data[22], w_hssi_rx_pld_pcs_interface_hip_rx_data[21], w_hssi_rx_pld_pcs_interface_hip_rx_data[20], w_hssi_rx_pld_pcs_interface_hip_rx_data[19], w_hssi_rx_pld_pcs_interface_hip_rx_data[18], w_hssi_rx_pld_pcs_interface_hip_rx_data[17], w_hssi_rx_pld_pcs_interface_hip_rx_data[16], w_hssi_rx_pld_pcs_interface_hip_rx_data[15], w_hssi_rx_pld_pcs_interface_hip_rx_data[14], w_hssi_rx_pld_pcs_interface_hip_rx_data[13], w_hssi_rx_pld_pcs_interface_hip_rx_data[12], w_hssi_rx_pld_pcs_interface_hip_rx_data[11], w_hssi_rx_pld_pcs_interface_hip_rx_data[10], w_hssi_rx_pld_pcs_interface_hip_rx_data[9], w_hssi_rx_pld_pcs_interface_hip_rx_data[8], w_hssi_rx_pld_pcs_interface_hip_rx_data[7], w_hssi_rx_pld_pcs_interface_hip_rx_data[6], w_hssi_rx_pld_pcs_interface_hip_rx_data[5], w_hssi_rx_pld_pcs_interface_hip_rx_data[4], w_hssi_rx_pld_pcs_interface_hip_rx_data[3], w_hssi_rx_pld_pcs_interface_hip_rx_data[2], w_hssi_rx_pld_pcs_interface_hip_rx_data[1], w_hssi_rx_pld_pcs_interface_hip_rx_data[0]};
		assign out_hip_usermode = w_hssi_common_pld_pcs_interface_hip_usermode;
		assign out_pld_10g_krfec_rx_blk_lock = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_blk_lock;
		assign out_pld_10g_krfec_rx_diag_data_status = {w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[1], w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_diag_data_status[0]};
		assign out_pld_10g_krfec_rx_frame = w_hssi_rx_pld_pcs_interface_pld_10g_krfec_rx_frame;
		assign out_pld_10g_krfec_tx_frame = w_hssi_tx_pld_pcs_interface_pld_10g_krfec_tx_frame;
		assign out_pld_10g_rx_align_val = w_hssi_rx_pld_pcs_interface_pld_10g_rx_align_val;
		assign out_pld_10g_rx_crc32_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_crc32_err;
		assign out_pld_10g_rx_data_valid = w_hssi_rx_pld_pcs_interface_pld_10g_rx_data_valid;
		assign out_pld_10g_rx_empty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_empty;
		assign out_pld_10g_rx_fifo_del = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_del;
		assign out_pld_10g_rx_fifo_insert = w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_insert;
		assign out_pld_10g_rx_fifo_num = {w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[4], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[3], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[2], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[1], w_hssi_rx_pld_pcs_interface_pld_10g_rx_fifo_num[0]};
		assign out_pld_10g_rx_frame_lock = w_hssi_rx_pld_pcs_interface_pld_10g_rx_frame_lock;
		assign out_pld_10g_rx_hi_ber = w_hssi_rx_pld_pcs_interface_pld_10g_rx_hi_ber;
		assign out_pld_10g_rx_oflw_err = w_hssi_rx_pld_pcs_interface_pld_10g_rx_oflw_err;
		assign out_pld_10g_rx_pempty = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pempty;
		assign out_pld_10g_rx_pfull = w_hssi_rx_pld_pcs_interface_pld_10g_rx_pfull;
		assign out_pld_10g_tx_burst_en_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_burst_en_exe;
		assign out_pld_10g_tx_empty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_empty;
		assign out_pld_10g_tx_fifo_num = {w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[3], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[2], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[1], w_hssi_tx_pld_pcs_interface_pld_10g_tx_fifo_num[0]};
		assign out_pld_10g_tx_full = w_hssi_tx_pld_pcs_interface_pld_10g_tx_full;
		assign out_pld_10g_tx_pempty = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pempty;
		assign out_pld_10g_tx_pfull = w_hssi_tx_pld_pcs_interface_pld_10g_tx_pfull;
		assign out_pld_10g_tx_wordslip_exe = w_hssi_tx_pld_pcs_interface_pld_10g_tx_wordslip_exe;
		assign out_pld_8g_a1a2_k1k2_flag = {w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[3], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[2], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[1], w_hssi_rx_pld_pcs_interface_pld_8g_a1a2_k1k2_flag[0]};
		assign out_pld_8g_empty_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rmf;
		assign out_pld_8g_empty_rx = w_hssi_rx_pld_pcs_interface_pld_8g_empty_rx;
		assign out_pld_8g_empty_tx = w_hssi_tx_pld_pcs_interface_pld_8g_empty_tx;
		assign out_pld_8g_full_rmf = w_hssi_rx_pld_pcs_interface_pld_8g_full_rmf;
		assign out_pld_8g_full_rx = w_hssi_rx_pld_pcs_interface_pld_8g_full_rx;
		assign out_pld_8g_full_tx = w_hssi_tx_pld_pcs_interface_pld_8g_full_tx;
		assign out_pld_8g_rxelecidle = w_hssi_rx_pld_pcs_interface_pld_8g_rxelecidle;
		assign out_pld_8g_signal_detect_out = w_hssi_rx_pld_pcs_interface_pld_8g_signal_detect_out;
		assign out_pld_8g_wa_boundary = {w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1], w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0]};
		assign out_pld_krfec_tx_alignment = w_hssi_tx_pld_pcs_interface_pld_krfec_tx_alignment;
		assign out_pld_pcs_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
		assign out_pld_pcs_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out;
		assign out_pld_pma_adapt_done = w_hssi_common_pld_pcs_interface_pld_pma_adapt_done;
		assign out_pld_pma_clkdiv_rx_user = w_hssi_rx_pld_pcs_interface_pld_pma_clkdiv_rx_user;
		assign out_pld_pma_clkdiv_tx_user = w_hssi_tx_pld_pcs_interface_pld_pma_clkdiv_tx_user;
		assign out_pld_pma_clklow = w_hssi_common_pld_pcs_interface_pld_pma_clklow;
		assign out_pld_pma_fref = w_hssi_common_pld_pcs_interface_pld_pma_fref;
		assign out_pld_pma_hclk = w_hssi_common_pld_pcs_interface_pld_pma_hclk;
		assign out_pld_pma_pcie_sw_done = {w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[1], w_hssi_common_pld_pcs_interface_pld_pma_pcie_sw_done[0]};
		assign out_pld_pma_pfdmode_lock = w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
		assign out_pld_pma_reserved_in = {w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[4], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[3], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[2], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[1], w_hssi_common_pld_pcs_interface_pld_pma_reserved_in[0]};
		assign out_pld_pma_rx_clk_out = w_hssi_rx_pld_pcs_interface_pld_pma_rx_clk_out;
		assign out_pld_pma_rx_detect_valid = w_hssi_common_pld_pcs_interface_pld_pma_rx_detect_valid;
		assign out_pld_pma_rx_found = w_hssi_common_pld_pcs_interface_pld_pma_rx_found;
		assign out_pld_pma_rxpll_lock = w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
		assign out_pld_pma_signal_ok = w_hssi_rx_pld_pcs_interface_pld_pma_signal_ok;
		assign out_pld_pma_testbus = {w_hssi_common_pld_pcs_interface_pld_pma_testbus[7], w_hssi_common_pld_pcs_interface_pld_pma_testbus[6], w_hssi_common_pld_pcs_interface_pld_pma_testbus[5], w_hssi_common_pld_pcs_interface_pld_pma_testbus[4], w_hssi_common_pld_pcs_interface_pld_pma_testbus[3], w_hssi_common_pld_pcs_interface_pld_pma_testbus[2], w_hssi_common_pld_pcs_interface_pld_pma_testbus[1], w_hssi_common_pld_pcs_interface_pld_pma_testbus[0]};
		assign out_pld_pma_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_pma_tx_clk_out;
		assign out_pld_pmaif_mask_tx_pll = w_hssi_common_pld_pcs_interface_pld_pmaif_mask_tx_pll;
		assign out_pld_reserved_out = {w_hssi_common_pld_pcs_interface_pld_reserved_out[9], w_hssi_common_pld_pcs_interface_pld_reserved_out[8], w_hssi_common_pld_pcs_interface_pld_reserved_out[7], w_hssi_common_pld_pcs_interface_pld_reserved_out[6], w_hssi_common_pld_pcs_interface_pld_reserved_out[5], w_hssi_common_pld_pcs_interface_pld_reserved_out[4], w_hssi_common_pld_pcs_interface_pld_reserved_out[3], w_hssi_common_pld_pcs_interface_pld_reserved_out[2], w_hssi_common_pld_pcs_interface_pld_reserved_out[1], w_hssi_common_pld_pcs_interface_pld_reserved_out[0]};
		assign out_pld_rx_control = {w_hssi_rx_pld_pcs_interface_pld_rx_control[19], w_hssi_rx_pld_pcs_interface_pld_rx_control[18], w_hssi_rx_pld_pcs_interface_pld_rx_control[17], w_hssi_rx_pld_pcs_interface_pld_rx_control[16], w_hssi_rx_pld_pcs_interface_pld_rx_control[15], w_hssi_rx_pld_pcs_interface_pld_rx_control[14], w_hssi_rx_pld_pcs_interface_pld_rx_control[13], w_hssi_rx_pld_pcs_interface_pld_rx_control[12], w_hssi_rx_pld_pcs_interface_pld_rx_control[11], w_hssi_rx_pld_pcs_interface_pld_rx_control[10], w_hssi_rx_pld_pcs_interface_pld_rx_control[9], w_hssi_rx_pld_pcs_interface_pld_rx_control[8], w_hssi_rx_pld_pcs_interface_pld_rx_control[7], w_hssi_rx_pld_pcs_interface_pld_rx_control[6], w_hssi_rx_pld_pcs_interface_pld_rx_control[5], w_hssi_rx_pld_pcs_interface_pld_rx_control[4], w_hssi_rx_pld_pcs_interface_pld_rx_control[3], w_hssi_rx_pld_pcs_interface_pld_rx_control[2], w_hssi_rx_pld_pcs_interface_pld_rx_control[1], w_hssi_rx_pld_pcs_interface_pld_rx_control[0]};
		assign out_pld_rx_data = {w_hssi_rx_pld_pcs_interface_pld_rx_data[127], w_hssi_rx_pld_pcs_interface_pld_rx_data[126], w_hssi_rx_pld_pcs_interface_pld_rx_data[125], w_hssi_rx_pld_pcs_interface_pld_rx_data[124], w_hssi_rx_pld_pcs_interface_pld_rx_data[123], w_hssi_rx_pld_pcs_interface_pld_rx_data[122], w_hssi_rx_pld_pcs_interface_pld_rx_data[121], w_hssi_rx_pld_pcs_interface_pld_rx_data[120], w_hssi_rx_pld_pcs_interface_pld_rx_data[119], w_hssi_rx_pld_pcs_interface_pld_rx_data[118], w_hssi_rx_pld_pcs_interface_pld_rx_data[117], w_hssi_rx_pld_pcs_interface_pld_rx_data[116], w_hssi_rx_pld_pcs_interface_pld_rx_data[115], w_hssi_rx_pld_pcs_interface_pld_rx_data[114], w_hssi_rx_pld_pcs_interface_pld_rx_data[113], w_hssi_rx_pld_pcs_interface_pld_rx_data[112], w_hssi_rx_pld_pcs_interface_pld_rx_data[111], w_hssi_rx_pld_pcs_interface_pld_rx_data[110], w_hssi_rx_pld_pcs_interface_pld_rx_data[109], w_hssi_rx_pld_pcs_interface_pld_rx_data[108], w_hssi_rx_pld_pcs_interface_pld_rx_data[107], w_hssi_rx_pld_pcs_interface_pld_rx_data[106], w_hssi_rx_pld_pcs_interface_pld_rx_data[105], w_hssi_rx_pld_pcs_interface_pld_rx_data[104], w_hssi_rx_pld_pcs_interface_pld_rx_data[103], w_hssi_rx_pld_pcs_interface_pld_rx_data[102], w_hssi_rx_pld_pcs_interface_pld_rx_data[101], w_hssi_rx_pld_pcs_interface_pld_rx_data[100], w_hssi_rx_pld_pcs_interface_pld_rx_data[99], w_hssi_rx_pld_pcs_interface_pld_rx_data[98], w_hssi_rx_pld_pcs_interface_pld_rx_data[97], w_hssi_rx_pld_pcs_interface_pld_rx_data[96], w_hssi_rx_pld_pcs_interface_pld_rx_data[95], w_hssi_rx_pld_pcs_interface_pld_rx_data[94], w_hssi_rx_pld_pcs_interface_pld_rx_data[93], w_hssi_rx_pld_pcs_interface_pld_rx_data[92], w_hssi_rx_pld_pcs_interface_pld_rx_data[91], w_hssi_rx_pld_pcs_interface_pld_rx_data[90], w_hssi_rx_pld_pcs_interface_pld_rx_data[89], w_hssi_rx_pld_pcs_interface_pld_rx_data[88], w_hssi_rx_pld_pcs_interface_pld_rx_data[87], w_hssi_rx_pld_pcs_interface_pld_rx_data[86], w_hssi_rx_pld_pcs_interface_pld_rx_data[85], w_hssi_rx_pld_pcs_interface_pld_rx_data[84], w_hssi_rx_pld_pcs_interface_pld_rx_data[83], w_hssi_rx_pld_pcs_interface_pld_rx_data[82], w_hssi_rx_pld_pcs_interface_pld_rx_data[81], w_hssi_rx_pld_pcs_interface_pld_rx_data[80], w_hssi_rx_pld_pcs_interface_pld_rx_data[79], w_hssi_rx_pld_pcs_interface_pld_rx_data[78], w_hssi_rx_pld_pcs_interface_pld_rx_data[77], w_hssi_rx_pld_pcs_interface_pld_rx_data[76], w_hssi_rx_pld_pcs_interface_pld_rx_data[75], w_hssi_rx_pld_pcs_interface_pld_rx_data[74], w_hssi_rx_pld_pcs_interface_pld_rx_data[73], w_hssi_rx_pld_pcs_interface_pld_rx_data[72], w_hssi_rx_pld_pcs_interface_pld_rx_data[71], w_hssi_rx_pld_pcs_interface_pld_rx_data[70], w_hssi_rx_pld_pcs_interface_pld_rx_data[69], w_hssi_rx_pld_pcs_interface_pld_rx_data[68], w_hssi_rx_pld_pcs_interface_pld_rx_data[67], w_hssi_rx_pld_pcs_interface_pld_rx_data[66], w_hssi_rx_pld_pcs_interface_pld_rx_data[65], w_hssi_rx_pld_pcs_interface_pld_rx_data[64], w_hssi_rx_pld_pcs_interface_pld_rx_data[63], w_hssi_rx_pld_pcs_interface_pld_rx_data[62], w_hssi_rx_pld_pcs_interface_pld_rx_data[61], w_hssi_rx_pld_pcs_interface_pld_rx_data[60], w_hssi_rx_pld_pcs_interface_pld_rx_data[59], w_hssi_rx_pld_pcs_interface_pld_rx_data[58], w_hssi_rx_pld_pcs_interface_pld_rx_data[57], w_hssi_rx_pld_pcs_interface_pld_rx_data[56], w_hssi_rx_pld_pcs_interface_pld_rx_data[55], w_hssi_rx_pld_pcs_interface_pld_rx_data[54], w_hssi_rx_pld_pcs_interface_pld_rx_data[53], w_hssi_rx_pld_pcs_interface_pld_rx_data[52], w_hssi_rx_pld_pcs_interface_pld_rx_data[51], w_hssi_rx_pld_pcs_interface_pld_rx_data[50], w_hssi_rx_pld_pcs_interface_pld_rx_data[49], w_hssi_rx_pld_pcs_interface_pld_rx_data[48], w_hssi_rx_pld_pcs_interface_pld_rx_data[47], w_hssi_rx_pld_pcs_interface_pld_rx_data[46], w_hssi_rx_pld_pcs_interface_pld_rx_data[45], w_hssi_rx_pld_pcs_interface_pld_rx_data[44], w_hssi_rx_pld_pcs_interface_pld_rx_data[43], w_hssi_rx_pld_pcs_interface_pld_rx_data[42], w_hssi_rx_pld_pcs_interface_pld_rx_data[41], w_hssi_rx_pld_pcs_interface_pld_rx_data[40], w_hssi_rx_pld_pcs_interface_pld_rx_data[39], w_hssi_rx_pld_pcs_interface_pld_rx_data[38], w_hssi_rx_pld_pcs_interface_pld_rx_data[37], w_hssi_rx_pld_pcs_interface_pld_rx_data[36], w_hssi_rx_pld_pcs_interface_pld_rx_data[35], w_hssi_rx_pld_pcs_interface_pld_rx_data[34], w_hssi_rx_pld_pcs_interface_pld_rx_data[33], w_hssi_rx_pld_pcs_interface_pld_rx_data[32], w_hssi_rx_pld_pcs_interface_pld_rx_data[31], w_hssi_rx_pld_pcs_interface_pld_rx_data[30], w_hssi_rx_pld_pcs_interface_pld_rx_data[29], w_hssi_rx_pld_pcs_interface_pld_rx_data[28], w_hssi_rx_pld_pcs_interface_pld_rx_data[27], w_hssi_rx_pld_pcs_interface_pld_rx_data[26], w_hssi_rx_pld_pcs_interface_pld_rx_data[25], w_hssi_rx_pld_pcs_interface_pld_rx_data[24], w_hssi_rx_pld_pcs_interface_pld_rx_data[23], w_hssi_rx_pld_pcs_interface_pld_rx_data[22], w_hssi_rx_pld_pcs_interface_pld_rx_data[21], w_hssi_rx_pld_pcs_interface_pld_rx_data[20], w_hssi_rx_pld_pcs_interface_pld_rx_data[19], w_hssi_rx_pld_pcs_interface_pld_rx_data[18], w_hssi_rx_pld_pcs_interface_pld_rx_data[17], w_hssi_rx_pld_pcs_interface_pld_rx_data[16], w_hssi_rx_pld_pcs_interface_pld_rx_data[15], w_hssi_rx_pld_pcs_interface_pld_rx_data[14], w_hssi_rx_pld_pcs_interface_pld_rx_data[13], w_hssi_rx_pld_pcs_interface_pld_rx_data[12], w_hssi_rx_pld_pcs_interface_pld_rx_data[11], w_hssi_rx_pld_pcs_interface_pld_rx_data[10], w_hssi_rx_pld_pcs_interface_pld_rx_data[9], w_hssi_rx_pld_pcs_interface_pld_rx_data[8], w_hssi_rx_pld_pcs_interface_pld_rx_data[7], w_hssi_rx_pld_pcs_interface_pld_rx_data[6], w_hssi_rx_pld_pcs_interface_pld_rx_data[5], w_hssi_rx_pld_pcs_interface_pld_rx_data[4], w_hssi_rx_pld_pcs_interface_pld_rx_data[3], w_hssi_rx_pld_pcs_interface_pld_rx_data[2], w_hssi_rx_pld_pcs_interface_pld_rx_data[1], w_hssi_rx_pld_pcs_interface_pld_rx_data[0]};
		assign out_pld_rx_prbs_done = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_done;
		assign out_pld_rx_prbs_err = w_hssi_rx_pld_pcs_interface_pld_rx_prbs_err;
		assign out_pld_test_data = {w_hssi_common_pld_pcs_interface_pld_test_data[19], w_hssi_common_pld_pcs_interface_pld_test_data[18], w_hssi_common_pld_pcs_interface_pld_test_data[17], w_hssi_common_pld_pcs_interface_pld_test_data[16], w_hssi_common_pld_pcs_interface_pld_test_data[15], w_hssi_common_pld_pcs_interface_pld_test_data[14], w_hssi_common_pld_pcs_interface_pld_test_data[13], w_hssi_common_pld_pcs_interface_pld_test_data[12], w_hssi_common_pld_pcs_interface_pld_test_data[11], w_hssi_common_pld_pcs_interface_pld_test_data[10], w_hssi_common_pld_pcs_interface_pld_test_data[9], w_hssi_common_pld_pcs_interface_pld_test_data[8], w_hssi_common_pld_pcs_interface_pld_test_data[7], w_hssi_common_pld_pcs_interface_pld_test_data[6], w_hssi_common_pld_pcs_interface_pld_test_data[5], w_hssi_common_pld_pcs_interface_pld_test_data[4], w_hssi_common_pld_pcs_interface_pld_test_data[3], w_hssi_common_pld_pcs_interface_pld_test_data[2], w_hssi_common_pld_pcs_interface_pld_test_data[1], w_hssi_common_pld_pcs_interface_pld_test_data[0]};
		assign out_pld_uhsif_lock = w_hssi_common_pld_pcs_interface_pld_uhsif_lock;
		assign out_pld_uhsif_tx_clk_out = w_hssi_tx_pld_pcs_interface_pld_uhsif_tx_clk_out;
		assign out_pma_adapt_start = w_hssi_common_pcs_pma_interface_pma_adapt_start;
		assign out_pma_atpg_los_en_n = w_hssi_common_pcs_pma_interface_pma_atpg_los_en_n;
		assign out_pma_csr_test_dis = w_hssi_common_pcs_pma_interface_pma_csr_test_dis;
		assign out_pma_current_coeff = {w_hssi_common_pcs_pma_interface_pma_current_coeff[17], w_hssi_common_pcs_pma_interface_pma_current_coeff[16], w_hssi_common_pcs_pma_interface_pma_current_coeff[15], w_hssi_common_pcs_pma_interface_pma_current_coeff[14], w_hssi_common_pcs_pma_interface_pma_current_coeff[13], w_hssi_common_pcs_pma_interface_pma_current_coeff[12], w_hssi_common_pcs_pma_interface_pma_current_coeff[11], w_hssi_common_pcs_pma_interface_pma_current_coeff[10], w_hssi_common_pcs_pma_interface_pma_current_coeff[9], w_hssi_common_pcs_pma_interface_pma_current_coeff[8], w_hssi_common_pcs_pma_interface_pma_current_coeff[7], w_hssi_common_pcs_pma_interface_pma_current_coeff[6], w_hssi_common_pcs_pma_interface_pma_current_coeff[5], w_hssi_common_pcs_pma_interface_pma_current_coeff[4], w_hssi_common_pcs_pma_interface_pma_current_coeff[3], w_hssi_common_pcs_pma_interface_pma_current_coeff[2], w_hssi_common_pcs_pma_interface_pma_current_coeff[1], w_hssi_common_pcs_pma_interface_pma_current_coeff[0]};
		assign out_pma_current_rxpreset = {w_hssi_common_pcs_pma_interface_pma_current_rxpreset[2], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[1], w_hssi_common_pcs_pma_interface_pma_current_rxpreset[0]};
		assign out_pma_early_eios = w_hssi_common_pcs_pma_interface_pma_early_eios;
		assign out_pma_eye_monitor = {w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1], w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0]};
		assign out_pma_interface_select = {w_hssi_common_pcs_pma_interface_pma_interface_select[1], w_hssi_common_pcs_pma_interface_pma_interface_select[0]};
		assign out_pma_ltd_b = w_hssi_common_pcs_pma_interface_pma_ltd_b;
		assign out_pma_ltr = w_hssi_common_pcs_pma_interface_pma_ltr;
		assign out_pma_nfrzdrv = w_hssi_common_pcs_pma_interface_pma_nfrzdrv;
		assign out_pma_nrpi_freeze = w_hssi_common_pcs_pma_interface_pma_nrpi_freeze;
		assign out_pma_pcie_switch = {w_hssi_common_pcs_pma_interface_pma_pcie_switch[1], w_hssi_common_pcs_pma_interface_pma_pcie_switch[0]};
		assign out_pma_ppm_lock = w_hssi_common_pcs_pma_interface_pma_ppm_lock;
		assign out_pma_reserved_out = {w_hssi_common_pcs_pma_interface_pma_reserved_out[4], w_hssi_common_pcs_pma_interface_pma_reserved_out[3], w_hssi_common_pcs_pma_interface_pma_reserved_out[2], w_hssi_common_pcs_pma_interface_pma_reserved_out[1], w_hssi_common_pcs_pma_interface_pma_reserved_out[0]};
		assign out_pma_rs_lpbk_b = w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b;
		assign out_pma_rx_clkslip = w_hssi_rx_pcs_pma_interface_pma_rx_clkslip;
		assign out_pma_rx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup;
		assign out_pma_rxpma_rstb = w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb;
		assign out_pma_scan_mode_n = w_hssi_common_pcs_pma_interface_pma_scan_mode_n;
		assign out_pma_scan_shift_n = w_hssi_common_pcs_pma_interface_pma_scan_shift_n;
		assign out_pma_tx_bitslip = w_hssi_common_pcs_pma_interface_pma_tx_bitslip;
		assign out_pma_tx_bonding_rstb = w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb;
		assign out_pma_tx_elec_idle = w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle;
		assign out_pma_tx_pma_data = {w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1], w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0]};
		assign out_pma_tx_qpi_pulldn = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn;
		assign out_pma_tx_qpi_pullup = w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup;
		assign out_pma_tx_txdetectrx = w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx;
		assign out_pma_txpma_rstb = w_hssi_tx_pcs_pma_interface_pma_txpma_rstb;
	endgenerate
endmodule


 // altera message_on 10036

