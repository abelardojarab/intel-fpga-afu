// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// 19 bit val == const(4e1fb) equality comparator.  Latency 2.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_eqc19h4e1fbt2 #(
    parameter SIM_EMULATE = 1'b0
) (
    input clk,
    input [18:0] din,
    output dout
);

wire [3:0] leaf;

alt_e100s10_eqc5h1bt1 cmp0 (
    .clk(clk),
    .din(din[4:0]),
    .dout(leaf[0])
);
defparam cmp0 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_eqc5h0ft1 cmp1 (
    .clk(clk),
    .din(din[9:5]),
    .dout(leaf[1])
);
defparam cmp1 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_eqc5h18t1 cmp2 (
    .clk(clk),
    .din(din[14:10]),
    .dout(leaf[2])
);
defparam cmp2 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_eqc4h9t1 cmp3 (
    .clk(clk),
    .din(din[18:15]),
    .dout(leaf[3])
);
defparam cmp3 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_and4t1 c4 (
    .clk(clk),
    .din(leaf),
    .dout(dout)
);
defparam c4 .SIM_EMULATE = SIM_EMULATE;

endmodule

