`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C3D51sAwcmM9yWiic2Y/eeV/gMG8oVefZcbBf/GKw/pCNpip+bDsCBGNaUVzc2Co
SHpzH9/KnXbewXEJ5gyrItuktWPpDitHPhUgng6T10zcvDoFFrxLDRrNjAEEpXWZ
GJq4EFBHGi6epxJiKnvEVaXyV3Zr17mdznaYAPqGsEo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4096)
anL30IwMoSnMku5iBbYhOe9rvmSFg9WezmS5ospd/9gK9/LupErkGXLVrUiNCjbt
k3RIXGhc1iAXhwEjt1bEs2pYBTd2imVmTjhBH/qxYWH2m6nkbl46ruWfEaHoZ4rp
2U6vZs6Mw7zaO5KL7V0ea7LzFwW5fC1f1fLpM2PPpwhVZC02cC0oR3wWPgVsf7O9
RhqLzmVJmI0ub1y3K3W8Kd4Hvi5Q1jD9tmB1gWi95+RXiyF17Ev6KcylflI5mPRS
b+JFEjV0Pier+k3Ah3a1xNODWt5DfB1R1iaoy3+ztlzquUiUY0lvU368UJk5z2zu
MGexnq6OOL/ja+wG+7vm2Vk8j6TfNKBWMfk4tj61JkxyECyuULYvv6lvVzpxKg8l
iFPhf7eB+aB9XINIVxhaMW5BucQ048iOO0/J27F0dSVy/DF79rz1KctNMyGEXLxC
aQLn0mDvmYaNudVjTrIqiVLLBGMQzF0PER/0Q9Q5VtYkohcLmFTSJCH/GtrVeww7
iXHHafiJ95W8j61254BuZYszN0k8VOQ7xW3SJpDrAsp9b8Z2Eu6nqVQhGMy6IqxL
KA+8qrOrzWdprs9UuQAd2BBi457+c0/U2JFPFU1uo25vWVqU3UaE8Xp4+AdCSGjf
vXv5yJXB8K4fCU6OOGprm4XNKYzbne/QviOqsm3Qmaw3b2V2BGCSpE87o/KRAd61
QLfPl21uLfmxCPVa0KTQlEX4vt9pY9uPNUPQpAIEKLhhmjThGX9uPzebKzs8H4/h
0YZPa+I5fprELPYxjPE80fKwBbEccJOhAkXZsGXWr3m5UxwSv5UvgP41gC+4sZDK
W0H4xoHGsntTaXH4glupT9eMCCdvA5Jn/nhbaqfGiDPpTgWuppu3WYGUNlGQbWDm
8fC8mbmRspjJNLFBl4dE/m0/cWIlOUODFOh4zYPzRmRNSi7xH4CeTrW3AMiWILsk
fx1Rhy8XqTxjlfTTqwrj5dC8YyM0dizUnHpdyR4TR4za63l5qvNVnJnA7APjAgPe
WfBaI+02b6eqedDXAQmVFCvxUohohhQEfPMn+ihOkeVcVRoDv55XLAKjnF8kH7LB
bc+0W278EkO/CSyucSrK8Ro/SxIaymn+DxcHIW+e7QUXxaWah0t6jIYmxZPEc7pQ
tNVF6ZT6j+6w72a/FuitW0MwC2oanxOB6S6yKbwIoj8p+Ida7pH33nw8WDS1gtub
mDIV7b2DKVGdRHWUOxeillhaqRsLTQb5I6qMAE9tog6r+sMTEVi2qeCJL1vh6097
HoaHI2JvRH1smXcBxYQY0PSOtrqznEyxgVjRbQiy9qDPIjx787lAUJRoauZXOqpo
BsWd2HMTAoa/3k82bFbMUesJs7fAKtZq5dFTY0JHAQlC0wwpMhF6VYH9dmiDGMrH
dElzRd8iXq9EijMPreFFvQaNgsYb4AciNPt338fbDvGIfqRd1SJGsbvisJ8z0wEi
n4dy58x6d4PNmADECWOFHDzki9IvQhFG+WNVIgPW5DGqRxz8otjxBY+9xaye1msy
r8FFeB9JrlaPI2ru3yfcSz8oHOo16vff43WoR4+NqYNB6/G3hkSYlfGoIlAkMZ+F
ZnCTkW6ErOUaL4WOlly88Oq1Z7uFco+EOFiG6jiqiZcQppdEuV7uWMaQAdd7FX6y
KeWfGsqtJ/GTH3FVZFfsQZuIg92KFK0bBnzilk5AUFyk2u1AcbjswK57Ps1+7Vzy
H0QPTMrfJdkLbL5pyAqakeHwJBVwF6nwdFQrhVF9u/GA3bOLzQZIC/Xz3j+8qJUh
hO+JtzQd3VsNH72oV2ApDS6yiEvm1gaK0jSieD9AZqQS98s002ghtUhnErVC3iq1
ho3xHSp44BCKh6JZdisnkHvkdP5kUHEAmBvWORACpRTqOWEfkpe6QaC+gRq635wJ
tTO/og2iSpJVx5exqwnXl7ImpSj/usp04cNu28KNpJWu4Fx57M7arjMro6onMuq/
B2fKGbOi66eb11jl82ZA1xFgdhvtxDY3a4ioWDTsraZCcAEQAheRSg8ooYeB+psV
BKS8CO/hUOCLxFUdz9WMfrk/aAQAj+jssT97doX54fpWO9xgwzsGaYUK+q6RqGAT
/yny5tAUsnWjMtDrlw2sFLMJkdDip3YhPu/d0Kv8DVm0QjFBPWQJTkvbM79yS79L
4EZ1sQixiJ1Jc4xNnPHezkd/1Wb3D3juDiZ9eOCjC+hhY+37yt0tfOLanwOaeHlc
4NLQGibnf20S7C0mEZygi/1I6Mc+2rpaHGINIMzrDaqfapjiWB7b7YxcV2SOQ+AM
PtuHZBNs8HKoAk1m4dFeNCn7FyisKxb27EeWrM1+qRhucA4/Z0jQyJLfbd+6aKAg
dg0sNXXTF1GvW6HsVDbCK7DRzhrcqVMXUDKSEPytJ9NTelexs26KTFL7jxdUjRgI
hOSb84qD1TIn0ntvMxG19jHFHJUtc6ak06zyxtWlCeBBYUzqT3Lg6xBjVb8m2zFF
jp9DuhwDTbMG1hMjIbxCzoRsoOf8DbTpZgbjIWvdiqNbRHX2CrQFl0OvQpuxZM1B
3bgXm734DEPya5NrvoLfsuewtAj0Ii1vF20utkm3szbcLuVmAcmmEoVxv5Ke4j8/
1Dd+gsl7Nse4lbIxrJ8Xm/YZcsQzlrkZ4KXVZnPuGG+rPGtZ/6kEhYtDa9Ruk8FQ
q3FldAlYiWGZrpE17w3NFWVzaF+W/NowONjeTyp6T6EW2oGap25WuxdVmK/JCHjY
YjyC1Ri+y9aZZouVtdz3Z/At2i7xC6ugyOBb29HdDdfsiz5wLFWqe71iFZwX+blA
AhKFj5AonBPJ/OTrv1jPYkwLML9wemjVFqexN1ZxHZAmW0DJ445A4aXnZGyhUwKd
m8bfmy9J9okv0iWEeFL7F9xi9sPsd9zwWbEecVhd4q4qhpEYtGh3ZyyAN38WnZZx
HPX5MiaZQrynuA0lzdkmXzsTpMEd8KVlPsmN22ytUt99fBitu8bI/QXxoNjbi3CO
tyTguZ8ixVhkFd3E38wUhgB40Qzw4aSeuUiS1iMrSLdsXOB7+8eAdBtY/Z69EuRG
Rwr2vQWnXveSnp3rcEnQ+9AtEpvvvvfDnoC4BlruX+vg7ASIrP8A9MtyOEYMG4hZ
8WFV6w0IZw7E3p33zTCD5AIwPliRhhBMcqtGxO3FO9EAPFVf56ZU+N2bMwLZkE1Z
IDADGdg9fK6Y78SZ+3xHDSLaJ1XFsWs+m8RokV69Cm5P9l6iAZ5jkTCcEEAYol+w
S+2ocGwEFmrv2P2SxxCS91w4WiFp16CDkcSNaIm5jP5Ly8mxYLcC3wz0vKEI75oQ
T8POR6RTp0Od//0TNVkd4wFu2MQ/K7+Y2xb+iPidsgFVVh3u+ey955MAO7+rribZ
U7lCmera7CBUivZWu+ugVeqLHaQve/E7m4zW0XRJ7nBC1HCBWZmtNb4fN+u2vfis
4uRxOhQ4CRJaZC0939Wa0IvdWvUTt/PH6ny3kP4gzU3jgn8FZV0yssxm5pXVz/fK
6x6/TNVGhAiBBy3ol5LpAoTOU8MN3ZXFUpHPN9g3EYyZaG3Rs/4GQ/TVVX5AfSTX
B/zy6Fo2b/3OahBsWeuYHNiTHL4jYPwq56cMbKX7e0lEtuQFF0lyqXhFULDUtdI/
JfkafxL1FyRvRr81MILj0Qg4BKhH2OZKiw3rfdRqB8yJqoH/DzmAEd4z1T32FnrK
QFjnNUX4rGr8+QxsCFAO7hb6ESClROdIyIDonEQVqFuCBd+6zLqSzizbkKHoEfpI
DFhHAUaEzo8AVMjziJudBmRXdgF5RaUe3fCTgq6ZEdRnvMylpdfns4GaF4vPnoib
VCrYTl6uKy8H9TVLiukxEAyjg75niy0hT9Ke/q5ChRceJ2cWH96zmwos8Cjah4UJ
Ta1aphJN0yTzIEV92cWTZPsRIzcGVoN8YhjOrhTPtjv64B5aFn8nxbyP8ThR2q9n
Vt3qcpP85NxDn/elqLRf43agip0Wsdr2y6X0XQyJeXWnZoVx8hpHl7kfJFIA7jmL
XHHpVOYOXmfaip1zbnof7JRdEB5Mptkex5eOURdemhlxam3DRZtX6i89fFQZFS0p
p650vSXZcviDOD85oUMSJMIInOi38pxSmoDAoCIFdcNRMZv3zDq2co1jLD/SuZ0I
xologY7xFYZntGR1iyZK79+ARShemb1c68BAEss2qhU8V1BvN+5R7x6xcsFByUq6
0ePO9ScA0PhS7p6QtlXjMDkqXYPEMi9nUQ1w5ka6WkKZ6YucGTcrL6qsDtFxiswV
Y7c+jSf2LFJ9Eaqy7RBH251pNWzRh9wCeoAI9NxRLCZ5x0wfuUJsFN/sFyZwG3US
dfln/R77Uc6yuZS2EnSHBO2RMrEzQlertyIyxC3dVjACvhR4Oi723/5sFc190AgL
2zZ9fzZg0mjCIOciWIF2G1pPug0UaQIzVxuYbXLzzFZpVp0Y1qwC5inm47vhTAGs
25C7mq1ufFL275FfCNLOXtKB3f3gj9PheYhrYM4dva+bExTkb2uDvVp70l0jvXi5
jHcLuqWi83w0JckrRHtZHgpPw8ENWzwwOtmWXZrpIbDfFZVhsb9TOCM9LYITRkvF
ukbq44FRvwSH3X9ZXxsuQV+QNUG2Bm85SXj3gxNBUdvIK/QbHY7ETW13lxk/1B/O
Gz9CzXD/dYREn/IpAYQsWBu7y1M6X+6dkeeDocFypxu+8nxytngPFlhoNm4RbuW5
T/HhfiR1+Ex1zHfJzl3trsWLWLFlbClH4mo341tsh3Mq6TJFQVpjHTUhWgAIAZH+
WbhmVb2Cfnbk4JC6TSt8UgcCZi7ICbj+Quz07nfp2v4dtNE1D7g/wJ4bjN9Qt/eJ
SskEmOWgv4do0yGFrCJeHPEn+SvV4ZgloTzmXXBXg5NGfWIYokOn0Z9B+NNEvfdH
3/wDuAsq8oRFjvqXsWf98T30jNFe1AuhsiMKbJwTs9b6sYaSOuZXPrxvmyuGwWj3
iasH9rvr+Q2S1Y0Uw+zTdsxGyR/E6cs86NriUmRyOGT78K3nO9QjSlg8r0rhnUx3
N2ZUduGjbHvn7AMdzKzd+HhQveuyp1wp/XwJvjPao7vNKtyuOa+RWWdRqb9RoArc
oB7KwLjJU20wbUts1Hcgpzj1VnkWnAzEIMTrrNpr1rqaF6Mepb16bdZ6dmW1AdGY
MmQKYwZlKYMykp+BfQw7OzwQyyVdRTDugKRzWOEbU/NRiJZ3ZcZcQ1IQgzKrHZ1g
JHW2nm/tEeygLivCb75sa+Ue6lSNj8vWwXarWPPF56iKkcncuitonGzpGsQthOoC
0dyUm+LAr9dcM8q2K+XpW1vOSX/QlrhDbF56NZSwuZzBY0UgL/wvPQkLfiv1VE4c
vouO/qdl4L0i1EfHefjea+mJf6VqVAH58o9Lgsns8fU84f76iVc0jvLJ2Ksc4fb0
27CsB6c8sN7kGA+U+5UX7w==
`pragma protect end_protected
