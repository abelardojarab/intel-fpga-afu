`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
le/26fRGZbk96EMJi9ALgr8rPfYqlWLKzCXV2Zq0nHNpLGxfjf4LraZTPhHP4LhL
QjKlVJZjjhiFXJ6c/uS7YCpq2Rkv1oO95qYtGmJOgKSzDCXNpa3RCJArfNHnCVmF
XUvvaAtGunma720EQg6CFDBdiTtG9+Vs4jKJ4gz4ksw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4080), data_block
vGe60qNktEjpLrf789mgY2Ozm9q83IXDn4h14bgCvOkPJtnIkMTRXy960TWZ/6Vp
T/93wT43j7RMF4qmSo/ohBGiSfqT4Cm6AxGLrL3DHY1cZKRyRDsLXCg8PczUrqI1
gcy217b3M27Wk6M4ijGbrQWCqURbCZ95OiEpIHaIyFkx/mHE+ebbQOfaJix8BNLV
FfYhGLlC5TUCJMWX0GBJIchiGcLfMEe6fNlZPIQKEHU6XbxYB3kFyXTBlPpHbbl0
y7Kz09FDacihMZckKqMkDWUo3ZlrFlsm9+VMGFH/2Tv9UVuAkLy9bytiMX9AWbnF
o62wBH2oCvzo6FHb1ldKoX7hBCgUGiS0JIOtgeMPclRTyuaXmXluNvS97DOwo589
TEZ/CyqX4f98bNmnGYSF+89Y2CX891iNgCVkJLoyjuDZln3bdACN3TWE2KtjqRmM
/goyanwgtozuHj+XIrlAsddWXClcmtugKOci6okW2rdFWDPNbjLhovq5IFb75Oe3
s0vlMljIhhTwX6sx4K/x46b2RxNdjjApbulsA3Z3Hchy6eUG/dVjEX6Pb52V6Qjo
Ueu4QPBf+/ZMjlADDTjLdfqmN6QFwrNwn4nYpG5MdTKI//PrjQ3rAxOQCMSPNin7
zQDodORkRA8PIOzHlKfhWPJXG3nnvQR4h4w6Ljk07hHM2nszWo71RYPtFRkpuCLV
W8hxe86YqP4DTWK8rAZj67KEhmUip2DL+UlOT9ng2ecJ8+Eo9GXw5waK+OIrHEej
QjDoyK7xuQzcP3eAOEsUDuUHkPiB5wlYSVO2BgMy8m9VgDRf7bVGlLMRYuPE8pKk
UNF0Kbq+NxmnUXhK+LrOAWjtXLDtWsGsm/XO1NPmoJdMt6LqjM1h8uSTdtLJ59EH
g7YCQzRNCkv95lyRwkCeua1WpfbuKO4GSO6FalCAU/oPZ3JpG9YXAkgqaJ1YgOST
tSJB/STAz4s1jie6YH+wWVWw8gkdQBABj13FLox4qjvwx73xWaUByLOKQb6KlzLw
/qDat8DN0EHNQlql6pPIyy7lyCHbtcZjhx3fvmhVvuRaofi/WRZINGITAB2XTH1Q
UCGlnELess9Xoy8wP36CIhX9+ZNcHPde5mkiF599kKuC/Za6skoDKBbGOn0pdaPG
3czKU4WcZjB6MLxFGjmiDMybgOj9twie2B1VbHxp9Qwq3AZmo5HY8GvmfOJuXNOU
2Dkt0JhutuFiOdHurqZ56y3f5W6A/mIp0Qu3lSQKkU5g2ufmG56hUDiqtv+QCGc1
f31pDB56GNrMmdNevXk40z7AjnNBO8GIVnXUouWzyqSedgbaYi1Em+t+mk36bs85
tnlayqrJuLcxUY1Zmjobt1O4BN3LR9wxHAoRmm6oG+fbu49EtOEuYw387KD75L9B
oQBgJvukQwK/A5godx0qBL6STiBHQv3nR8dlNuKTAfXysoVUYDHjncKRV4bXoOjs
P5TXWa9ppoYzsN0op6gcoN8t+pORmw87zxrtQfiJI7LQ+lwBdWOJqzy02GZVU2+E
V3KvFgFn+bY+JziP3LXNX0nq46jcNl8eB2PrIGNsm5C6GqJKiJvITGNpn0VWhyYF
iQNiZSdd4MJrEmu9/W3vnTXTSOo3l/Yz2rWtL/ANZSAOJES8ql1cvRQCH5GYRkCa
oVdA/wGwg2iFcbsi7wdp1S8tUVRDZqHdXxr1lPEnlRZv5ZrvDky449FQ9iOmvSYg
KaFOMiTaVOFzr1l8PDX6e4/+NoCIVd8o3PI+kmN7a5HRpJ480MBaAz/thiRUtRo7
sdN/fVG+RgTpkb1jtDwiyY9kIccvZ0FHq/oaubuRla5B6VFCP6AxZPlaftvVibt5
+tTztI9Fi7cxXQIjHnZOl7jAmQT4t6Tz+qqn7b7Ff5PXrXutQH4cXjEKh5wZfvIQ
cyoPSuZ2UpeI6dUFOaAemAZ4edJ0glwcNa/EMgdCzK1CON5hParrHf5F1X1PnXXX
XQXMuLZs8S1vc727TM6619uuixQKW644313Zah/MuycSl6oX9p6jeV23UahJnhNG
CTEevsSngpt0fAt+UAiiL+HsEduA85WqhInada3rsw0qQaI9pb44gErKzBR4D1Vm
CQYVBpmTPNCkNXxVFkzJ64R1yWlkQfYQO1eQIx/+1d+t/J/8uDqwlXUzTrXfYuwK
kWv1v71e6krOp5O0jQfu6lDpU+fuNPawcW7n1FcfrIXTPawl2D6HLsl5dcrlo2b3
Yn1t8rz9c7TybDij/j+PIAO71KokLkJP35bREnrXKJUyAFBH2n3s3MJYEad8yt1C
TnhjjZar5x8cfcirxZcZ1mgvjLwQSWknSfsbu+UL19FYJjQP28W7CaW1gOhxzb6V
DZqcAzwk1USmzSAlAr5Io5Kt2JrF8R1nwgMGAJvSHFW928E9BVsjfbt07H4pQSH9
G8utN4hhQqvbmQJtQOkAjPL1rLeg089XvjlyhvtqatMGXRh/s78+g5HH7wTb/Gql
IH/tifSoDGI0qQMIIQLdzmiwOG/SKwGL7YdYckK697H+pkAh4ZbV8cAQ0ElMHX0g
8xvGYa4huPIc4pV372++zBiflA5cwJXO5wkXcuiPi4rSlDguZKQJ5Lfubcre7cxK
ygO7zNE6oTqNhfLRaX3V5vZ9+bMfbWg6o1UPH+FKFF1ChMc907eK/iGnu77wclOX
Bmktl/hVezdCz8QkChoja8+Vk14KsPudXjaRhXVP/ftA6/eo83Fdu0HLK0dDd1Zc
UVe4QESNIPIIedFFMD4cTM5MX6b1e38S0Ebn45NMp6fCT+2Po7ZSufrpxraJyFqs
N2UXceYHx/Y8KxAlgNoahmwsh2ZgaVfZjVJi8DCwaWXKC7PwbLl66DqE1J0OEf8s
l7lQQvPJyUjzRTa20cgyJHyBVo6GUDcngPKhd27cU/rZsW1bApMBe3mOCYlV88gK
1v/yKWHo4FVlmuNWDGoQQbMCjxsea086FVadu1QW8qRd1W6rDigdqeymZn9RCTC3
rLsyofrOcarDpJzExvMTnHJ45zsaJPcTiL932gn2rNFf5s5BBfINjtien/iU/G9Y
W11KnDsnog9ID7soarxwVoD8yJHfQpax465XscFEr3TloqnHUe5cz1aqoIwCUD5S
7xebAc/77Z7Kn/tyAHaDp6i2bhTVVpJfW/gqpNk0lEVjaVPNNG31kG6oxGr5ai82
vr5dDiMN8Hm+5WTLX2IaxYYNCPoq4YhLWpcKHt3S40gCopOMD440iyU5gw1RXDyP
vtUdANNBTt/65t+kEmk3A5ITrtIGiTIkk9aBYoTtU3tLXfIC2LRgaLsO7oChNAa9
BfmIReWJXUcYOwnwm6+974LLhhf9IyRvHkaliSKIADIMkgl2YKBql9CwWfxiJ5S+
YQvSsbKeL7uX8O0rm4V6uB2YvOA0myX/ldUZSABTibhB8CVd960BNR0c1dtj8R6u
Aik+B6WnhK25yvk9R/5LzCltAaUfBnJgX0a1aRLrewdwujofV/ISIlhUBWjALFt8
GOYFajyiyHF60I/JDohklQVgn4Mb0UtahBFoko52+6xveYwlkF4EKj3ciqe/2tx8
k4D4Kh96kUFiF7/tPYROxBG2qIC57pfNfC690Dr1mMo5ARFdaYgtyxgRaVyjbhyJ
sWgJ4VYqW+okO7kFZU0whzInuXIra5ssGa2tQK+THWhMjnd3dI9bDKELSs1lTpWZ
2ooKOwHiHTniB0S3pNzs2ac+R9ZWIFOdj398OOMPRc3/VJ8xMxbI9wUxOnoiWcBw
uce6617BBDzhfzSbSarru01yhukociwTyIthlGyvDH3FMkcAD+VA6ecGHok+fqcg
4m3zjPjDZ0Pawsd9/QikrDDvptp74zGNP/z1/4z6cIsGghTbNj7EDShDhdgcC5QL
AWhDUvo3qD+PhkI/pQY/b0EPNF9t4AyXBAJyeU6Z7FheduXJG7z1TRi9Ss05PDDs
LFNbI9b1iE0aUhnptVg8ZuysESQR69RDj4tMSvChrqzdKrmJ9Xom8AsPbP5RVOF+
P8PW82JujkQtgf7/Z/68QlSBR/wWX2iOv2YFq1EYD+fw/XhH9Q/Y4++4TEwUPGtd
eH0s44UpOFdGAukMUDIq85GdD8TOZlRY2t5rexmAZD7PqVv8VPwStInhGsQnNvwX
73o+jQJhlZ+K31isQcr1aP2Of18HYNJgP1u97H3sJ8dRwJPnkMYfJUT6dh7Z8IL9
emozNSlzAcWqjOKE8vZd7lkTIy4X+TFBrjwNlaO1q9lxV8a59gKNafMgAH0VL6OJ
L+v2fv5ZBzOcvDTdKHWbByuhtMWK5/iBS0+a9H521NX1Rt3lYloHikqt+/qekFYI
JSYIwGl3L4Fdwv/EW/EUBd2wlX1qEkb7GqVKz9+IDq8aCjvFE00qj3gNdpNfbULH
Du0QM7vP+1MGVwzIxZ3p/1J2kuYmpZ9VzdPwcstgGY4tt+QWgM4eEvuiV0v0QtSR
5D7smw2MR8PxQCULeWNQs7xrZGQ2BdT/acZ1a1FFAc6d/LOcjjQgozh/g/BRXwlD
xMwNEAdQBWk9VM2PP3NBQ00oOn7a0vQpn2TAB45Ek1ol+Upe6Az+WkWBeki1Kr5/
lB0a8i+tkn8VTTBAv+ad/S5qDnPwQOJQo3dVP0kSun/bfSy4puDQTrgIZb+/4sL1
NKVQp7aQhw4F0KWNpsI9jpryiLfmz8OYcbyKKbrE5LfVroBiy5lwKxuJIuBZB3MS
1HEHA0BFojnuW3p3Tz+JhFtuDtPZBd1WGJTcw882O0yy4phISayBKtBajil2B8fs
XI9GSxXawmvd1h6ODK7mX+aLCLEIDRerblpScflSm+EwhQC7C57r8glNM+PMkF3H
E6vHlhx3XxpkdqbsZFRAmNtSp+xw1FYYKngO4Z8iA3nh1cp0s5Sc4Zj8xQnbXdtg
NS5XKLpRPP1phIo7aA2bdNr1C7CWs7ioYiCWXYnkT5WMDmfxkPAg4fgqbmWJYH7W
bW8Hho+6igj+Au076OvNut4hMi2gMrN1zJ8iOE8dJLHsXlOj3ehyHy982hyxTZeU
ztAwAd6qTPF0mgMRNuWR3fb3EI0j7Ni9o8Gwd82e0r4TMRKRi+BRQh5JzOpo1wDn
80ngo8BDicTrCU71AM/HQwnL0kHiJiEfeS8SCVVLDi9q+3TxxkD40nhAIgckNPxq
tUvm+CqYV02qE5BAdq1GRXmV8/EybDRy0TJGywHMm28nVadmJvGdJAsqshVs+3Qh
Cw2XDe9K+52zUWJwcBIiGYgTrknzSpZ1qfnJe0qXblIr3Z2/JKiUEqm2GxET+q6n
HqToyhSHBRCSm1bYPm6GpKxkld4xlUixDH7s64UmG738mo8NP2KZEepUsPRKDmeg
prTwCOSptVJo7y4MHlOJv2EogB8IIFXZk3YB9DV/9HBurobmJXXWtwkqfQX+OOwt
`pragma protect end_protected
