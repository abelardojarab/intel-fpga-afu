`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
nUpgGKccmUXt5F5LdQvZbPDh0dBLeriBWSsVmOEaRHvmw280uo6NDbDhdmbsBPOL
McQ7LCfMa3zIEsXMTNg8TPWoZ4/eGHP7CR333FdYdVCy5CewAl6E55GsVHnw2MFa
Kwz6bJL+h9lIQ/pJkFVGV86ILTWpx2w1U89M3W786uQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 28640), data_block
CI/72LAD/yeXazsi0cLTfMGmNIGcx7R6FnyD1knvZC3De5XO73unVyoUKrosjoBV
X41j0b2Rt/rptWdYBjzXLjVFUmNS1pO2l+8W/f0XAbjKSPL93rRAVSlmgusJS332
EWLEtr/kbzuKiVcUyG9B8mFJh/QdHg4/lDT1b1Is5XgZ/CGzgEaNeCFHy7FGXv+l
myf6kqQGpQeqpOuZ031/Y1fQ6+wK2/kHX6cLcVj7RfvQnnxQI5ASIDTlRBrJOrPr
VAlSO4sGrw7sPEoqWXo3x8xSj2mANN1wxvfEozBexgDHR9LQq1SvNBPTfbgrX8+F
lGlIrq15KPOb5v0+TUlvGQNKiabxlG2UuE0LB53ZlHQPVAE+ToFscJI1TlxVGWFM
Tq7+MxtNLIk5tUNgJq4dTkkb5YmfwA/FbRo9M9Eyrx2xqWlqOntzdQ0/7/9+axl3
DFmiIghhPcMxUpIvWhWN4abBHHvvT4ZClvsac+rL2Hlqt2KGCz6TVVQbIDWNYEJv
vOng9rTAFTdKngbvBlppG8RE6G9j1RANUSuhItwZbr9F97xS/VZtmy77mPbN2tji
GnmwqlG+7natOom0nu0KMFrd/+Iry944Fm4fqoI2ZvMmy+pcS79FIsqQjbTZEotU
TxM4iIw0gTzDJwZkp2Ym0MGdxIE1qNxfylMuc40CCE+Az26Ecfd8mDCeNOrihGBI
PlXa5l25+qV0Gwif5iq0OOMRZfAFWwMLqFJB+UkVP7VDOUoQnLHES9fex2utDFBp
Xc8i9cD8EK0WnzkHhF6DzIQE4z0gIHISXUZlZqwnI6dyp4vyeEzB0AK4u/gMqGou
1nT9pt0MZOT7OJjy64ivIbzi5JmAykTRfETmluycTfo0rbAFPBtYsZQWdmq34CUn
uEJltEHGxHjtG4QP/ZSCPmZ7jhygOjjrKs4KejSrqeG/I7N7L8limUvaJmpurffh
Rj9f7TzfLSKWwkzo3c22pCivTPVy2raLYDVrd+b3wKn5Mcq5YEfjhJ1FneMiOYhJ
iOzpSgKAUmqwxzDLdGQan8cnE5KTVeKoXO8uQUyK4FCqxUomIHXAQGD2Hodp+09A
HTvJMcV+LLTJ6omWAPrbttZJsjuLK1QAbvz5bpucXra2NeOsgsge4OCxAzfsG0S8
rIHX9yr86kDvUn2he4/0VwKmCYLaSuXM3uzLeSEx2Gm2t83uAT1yhKMgQBmnFjac
WYt5g9Jjeg7pn5REG0hRUWV5Xvy2n2nol9knF0PMPVrpBpAHu+tpDjhVzNgWkehf
wL/RMjyBiZyk0ntlVfgt8sM0ZB6oDlXm4ECYqY/uqa2bvEJHahPPm2dQXhB+uAZB
4HLxNUD8hIxSxoQX3vWM7b98yaz9vLUBfqEQOSRak21DjgBfaw0cvCnvQQp14wCb
SPWWIvcOsWfRc8gwM0t1rQmNJmhLFSTBlFLox1ya4dvTXi6Qz3Ikoypyt3uGEx2q
lBNPjuETY+k+3Sn+yZbJNYXWLFhH8iDXJQZ4EPx0eook3QAyIJXB9c7d/5o3a0xy
cfoL1FHpMluc7yqai6KiEWy6TtYz458D5lfzHYlbTYZJuoPd5izkskSuz2X7sY/8
e7jNzBRg04KtNq4+tTwcJBpeif7MYlI2PrmiTR6PJc07KASKdtsl54HsRNqTTNf0
ETj/sS8pzQJiLCVxW/VYhltvVB7YSb1Hk8HJsg1SdVl8O0Kfc6yDrsaK9o3jeMbx
BAXNXbGgOK0vh+NhQ/sCgyL3JY/uZ1D5HlVJTB9ZOBeeYq26WZdV/6vIq6qpSpL6
ud9vl61Zs6+iBy+wfvof/DOTS95mOIQg/5PGv115fKiNh6VEpN0kjNSyRNPGubHy
Jh0MOjoRR36HXImxYH0Mi7eYNkQRjQn/LoyhPJnlJrtRwBj9qGZpXLBe4mMAHQp+
VuLHN6RKzy8im1jzG2B1uEb50wdAiCYvkguYltOTKc+Faz4HteXtfo1Yk6vDMxXR
S4JIVWwxo+tvU/bSA7p54DtO1Ytq0OLhtLE7lFq+l4d7/9L39Eddq5qTAYcsAKF3
YCyP1tKYwyEVJLNHGM2o0IMmQOz1ICIW3tdRsAzSwe+P+7tNL9dnIDwqN+NfA5S5
XIp+XK9vFUrex4+/yXfLnbCBsZxQF/cKO41+SvPyKvRViAQuTzNtnSOfNYCzmM6s
KN6pTry0iCSe6DFQIzqFAosPoAJosZJEAgPO9iT8Zt4U6KNe/IRZDCXAqAway+ki
4e+RBv25N+cTMMJKfL0Bd4aWNFuKMtGnXznXkZofczOlvLWrXZCX+GbzMSvJMPMB
fs70zfJ+B3HAg/vRfiT7pGm55Hr0IAyF2Xz3BTMr2nMhwTots48nPUw2yCsOFiVA
0mey1eFR1JhwPnKBzTNavaWf6497G/oqvD1mIgzV+gay0rHh4cYJMKgVI30hio4h
JFJr3CEi569a4vRtMHqiNxRXp5fmIO+ohP4dUykRXGhqgnTm2UOOZmTUEE3rHoCI
g1sBSivzaleUdWzs5lf8UzcKLd2uY25HbAiT6I6wjXUepzdAZylo6aaUnSBSmIII
VACz0/YvtrF0mvRjUBS1tHfxFak2timj+658JqraegZ6YUuKEd6QH96qS6P+h0Ty
DjCaULvn9LFb3NxcULWirXMl5PdTiQ1UKN7SrOXOa7XkMJj9GnVbJ9LOwMhFoiMG
JgAyzkDd8QL+WUskFcddhhEI+Fwfrb42MnuJylnf9k6b0FEAt/rg9HNojPVgFRV0
8q50u+lkpCsXPstVbw0twcW7XkjtU/xzBwx0f+bmIVd1EvTqNVNZRD6ENjqesADL
NH/lr9zt0A1v09VW+L+O77SbL95VFSTdXVt1+jC2Y/9MzXTcBjh6ogCmb1TWRO/r
1RHXgw2jMgYTiTOM43KNjsQjb6sDKi72r8+wpDUVQJmwfvx81X7BhbWA9zqrCyte
odKTQhYcPowQ/kdTYRvEAlnKUyMAwsKC+rDk5w5x5vAl2DosIDqzLXBGcA6KGO1Q
MhZ+0IfqqKzhSKJafxjS8v/+wyYibQgLlipzZpybdQOUnP0VzeeuaoaODvoq4pmy
f5TMRENkEs5Qm8TyzA1J0D3Ug073nPuTM+rQDlbCFebT80XPZsagXGPwtuU3j3hE
X8WfgEbPJj5tDi5R+wjQkRwg049RTSej3589K5pTZNPasX+Em6Ww4v+srqp+YUOO
+mPf8pyEN2r6foplfpU6MekTvHeG7CrrIkkyz7+MU4L4i8Em6TwpminsDbTG86UW
PnCjdkANUGFZaKc8GUHonYTzxmyAzyBUXwIUiXKQsHNF9h6+MX4+fcUNyepXXWt6
NVuuMvRRazttM97L0rLIrw+XC5d72JfK9Tz06R/1JFjj0IHJrL8yZKtKiyO8DkWP
j1DD9jF93vcCZZR9uEnDs/th525o6Wa4oO5zmEljhmYuwpnYBSwfyRqiZsroY20Y
8Czss8TNGcP9TEtP+2uxZF6VT1MIsM6jHNxqjhKEw80PBq8cyVxFKJWJOnH9zdNR
vVkffe+Cjge+RWTpkSWgTdgCWHij0jcR0lxYVNjG5U1CiIl0FiU5gdW0Uo6JETt6
WcOWAKuffLlnwS5EO1RQeWMdAKnEwA8AR5Lm9SVR891X6OVbatxm+B5Q1eQ86RV/
iWIxdguhYWDND6leyrg27wOOZ0J19GZ+DHGTtqj/er1ss5octZwZ4P7YAvRp7+WM
THeLGqUWRVrxGcdUm3IjrqnnTTswpNxlY+4wXW0Q8X9iuFvEw2KA37Pxy9TDyMAm
QlUOd4KP+boIoTZ9FR3JS4/AOCUBtrtvkQclPCTeZu3CLZsXQVsU/qQtE8u/s9k8
IxwbvTmmDURxF++KehD93yBl5OOcASprAMa9gRqKsU4bw8M/27ej+u8bRggORLim
ofl4nQIZcTXXOg1F3A2d7NviQHSS9gD6QXe0TQvLmrEF5/Fx9kGNxhJx3+YIW97+
9o+Q4jthzhtGh/1q6Np3e1979XKQyG3WYWf9+h1WIjdSGZivBNhJe2c80XupYABp
dVvLcKYVng2GB5FzlO/4hKk6vPOEvc7q3kABp8FgGjA6j/XxMso6y7jpVJ3VuN03
JB51VO37V383MAIC/yl338WpWVP1ZWSd+JVNmIyTvcl3T3qIyhMJwUb7WnduiET/
5PqaH556zBPVhMtHbQRKJsr+Muqlac0Oi3Mtk0lHY2hU5HQ7HVg7dVE4wW/rDPwa
WH3R3fhXSFUtKBn8t7YF8vOogtfERC14pbM7xwiiekM9dhgyr820P2gtTiPfgtAH
G0NCydxgFOsQfZ2pgrlH0OTi5F64ZO4gEZI67xxZWsNRjgw50QeELohkHc1Ss47I
SfdhjoP/vZZ/Qw5AkI5K2W9RPRfkZOkI2r/DWutbSnJU2s2JMXWEDLqKrjVT+Go3
TYZH4NZu1qm5WRkApnQ1HnJMH1NdusbF7llOaBIO8So46vqgAUsq6oCR4Nt2ys+U
nohgVhvwla33tQK8gvqOpbGRhGRIS1u+TYf6+O5WYn/Wq2qbPAhVdvJuDfYlFS7/
a1ZMXzQzvbiDexbGDBYyfQntGTHtbK6Tuz9Z6wNxacVxJDoi1NMpL/k/R1ybYpfm
CGFF/wh1lTTZ+JZy6p2xSLWCZ44wHmnJhczGsKPcrRlN9OlMKf9/7TPD7u8ZOYEN
tBXp19IKZ28Uo/+HV1UMbfCN4eEZ/F3IiUISq+a7PHHM+iPA3z3TG0LDHQVLlfCb
rJT3JRL8yv6GY0C7icfr0X7nXKIlcD+4CSQXuvjXHT0UlydzHsv0hb6iDvdH0p2Z
xyyAtTCF3/KVF7NNxARSk5C99PDBJmQzP670uarz0npuloVuS+s0YWxK+qRxPQNF
zxdYjbhzfnfImdsLz2FuNk1uqXlwXDr817ggpzekhiC/DkYT/FeJZ9jbMgpcK5Mp
IM6Q+48+VQ8Jpy0dOITv/5di66d6+Lm7ezqta8q9ok8zLg+f7XHEc61/dE0hLti2
/z0MQfV+XSuv7z8IyWMF9Lt28TZvuDJZPK9fg6iZMd3NNvvT7DH+eyvrudsvJOzv
yKqHFFYgJi5pjSG0FXsXzfCFi8PkLHNcVZ6TuCL6p0M3CPp25FN9iPjDmUGNWOY7
fupXM9gjpLgpm5CLajebopH4hKpo5ULIx1m1oA+Qs3dzADdI6qxi43NPY7itl4fw
RXI7S7lrxVur81BjhmkW42DqNjQ29X+32PzJ3xQODvHgRQqCqPjcwLNXakB6qP5u
yk5svYk2tnP3aZQ2ym2KkN0hD/PRLJTeEnrYMkFgkFGxwxawrVBVQGu1Sdd8+JKN
dYgItqHzy0z9n9XLGDq9xjnaUyNDdB+t4Vqt8RZabxpiRLu7hF/5191EAzo4a9ja
NcC4pI/p9hn4RJC0KQe+FaKS44ewluiY2msJtJXwX4AvDTpXTodJGdSmQ7aQtJWe
Jy6lK8T5hhfjdBzZ9QjqKtBKpSFOoS7+1etB3KMMp4T8IVo9bODEo21n6W0x8S31
G5tIXJR5Q9ZmHWOTbisTeM9PlxJQzAgHGrdpt/ukBi7d4+w/WHXEaayQYOndAn7Y
n+VcRvPyl85LcIHUtuuM5CVBNxLtdF6L90+PWtg+4Pyr3DfP1/uSzu6S5lh63/iD
CsVVIUJqPWde69Pn6ezdx+iIM3hec1cH5Xd4OwCbEZv/pfLZsxAFsLUM/btjHu9S
9UqKw5CVH++bgEnIGY/WwAkMdVvA7JjIBjwYcVmcJ8U5P2vQlXwdj4HMlYKg0ZdI
Edt7kLX3JjGinbnQfZuxsBLF2pXB2gJF7neXIX/g4o+io23MjO10oKj4rccJGAM4
1VnKrujCKmXVRfZdyihpoy+GWs2sTidRNvT9Zh1+VvTvYiKc/+NNM2AIbI5XypHv
+be1P7ya7xRwEOpe8ObdTcfjlxMtyrRvwHOWWVI30lQCmrc1g5rJ5T6fUPSrczCP
gsd0B25Y3/O4a0AbDAaJJVKl/B/gKp9ouECaKUHIlqhBfYFrX4Ps4/r3Lpdf7/zH
asIrJqonNFgUjJsxkRJ9SDUkp4SGoAn5Zz/xGp1v6/8gOINyL5ljC+3RR44tupzN
BXisHFbBW5jYx4+kZSUKor+uTIj1io7kPpXewHG9w0vpF4J6t5n/e4URKJHHaOrd
wRnJbFeXSi06aZqqPbhRH7f3YlnyMCTiDu8btrgIn/NlOf3JRabbIccq8spgOD25
H1fqJx6vjDcETqYAbRk0StMxWzQfhD311cQFqdpjVV8LoEPeTGEXY5RWN0QIqXBT
6Fj7Hxu0opCwrlXCQpsKAm/b0WCJsSeT5Ntr8MnvgVNyxY/Q/vcLVp9Qb7yZWUoX
IQLo3QeNzwNTyAhOkvgLzPs2TEgwogbRiOZwu5OjCnBXfDYPWQg2s3UF+KQYevny
vKE+/BjsOr3kj96ZLIoPlCwGoyxpP1PuJ4jSx0fNSsAQtAhEdhzYhQ+d6GDW94LM
FcEd/PgwFE4d0njy3CDjPWGX485498Z4OZ4QXryQAH7j8vMxNpzu3Z6sUtsRmw2s
rCRwMqPTJmWd77v04sRNB8Q+X3vmFWS3LGpOHEJl8X6HrLZtWTMOkAn1RM8tttas
RLQRqfdoBHVzWzSMoVZFnHXf8QNaskhx8waaUDcnbqPojIavPFgGcPWybJfHJmda
WR6/kQDofzHqJXy3yrEMpDLlTjbm/DqggNnkDcCeizww38Dzq/5ViT3CrElHycot
Sq2fmzXdAhU7t2IL2pu+VZTEVQdBV2sGij0aHVy/Kmf6hImjWKVcKE2qDgtIfJYn
HOk4Bkq3HXDeLjX0/hhS0QHY8qoBQ1VzL2CKGm/DA3PXLPbJVcXnmjjunCMoU+KS
3joAvwCexdWnOadtb4kRkQZK/N5WjwDoIlKPkG/5hV/3vgLy5G2UipMho1aa5v6T
LOmnjelD63qDXqSTLXRqFXgChB2YvX7Ub2u0KhWsaTbmL9sK0ppDkGv053xOO48o
7cvObKU0VtaVPS9FcDzekCGMtfWNKo6ADcHo6eV2+f0gACU2mH/g/mQcn1IxvkGk
XM47WXE/+aECAtkNcTrn3s24XQhh4cB4qqJX2UfLbJW1+6m1XXAcCiNlqdXEuFGU
B32lWAGyUaE63+Yeo+e0tXmCeacLKq81we8iyhOFU7xbK5gQsZ4d19VXThk12Jli
77Fy0sDUbimkDtN2rp6mYuw3i/EFoIFHwIOADd+CqzqTA2SDNEx68A8alMFm5joI
zk/ry8zV7rPj/IA+EiMUx7dbv9UlFDzi20cKpyNrxxNJoZNF99wab1dG/6r7/8dL
EeAHm76EtP0IeQ1+fofVnujrHn2qKIdO/YVAqZIZyo6RlUT21gDKrhqKZuJqwRj/
mb3BFMmd4ygzsJ/hlMI5hI5i7d01wMcjcJwZPFJwJka6yqFXWCCBzapUr+eXDBXI
ZTV8EI+2RNk5UzHEDMDGV81VZ6sEBdE0BiFiGBhrPiF1hGA8hy5fWd+YSx6ktXPY
eQRgF3CsGGADqJPynvPWpJMQC2aeqKYvaSFKmeZAK/BE/h2jy+lE4BbhkUI0utXp
5h+gZ6+iKCrEoccPuar3taqYPW7guryo0F68GhGr33V+jO3LLX2STL/S+jpfojad
j7UscPtnlzsHzhci9Dq9XzRCLCmQhJW0KUvxmYj0R9FMQfZZdSi9mtJwXrLNE8zH
4Ve22d7kaelnHwnbjcFKcyk+gw/Q5s6Dn3Z1j+cAaIp1g1RI72+nb1vQLNUMO5Qu
rPDXkKhYNusOuRka27tAkWCyq+s9OQyhZbgbFAYEGnONCl0Tni4Sroppl74FS7ja
OKj/XI/z5u0kYMpVfAUbAecQk+4gbkWiM7MSDbaOKv1TRl0fEqA0mYGXgxVEqEu3
dycykMJjuqJWtLem8yW9+6UK7XK/Scgf+cd2aGLwuZwrHbOyZloYT+72HIYI4QXM
I+90R8yLQAcIDflYjwAWhbngczW0dOkirw0SI1iGi3uZeIC4h2X+EekVoNYvPR9w
/m/gUD/yNFKFrz4mdmyEg6v4ceHxmN56lhASmZiS00da4aFjoS0eAlivY/RjNI+p
ALEQxa1fTMiEt2IBcF2GyF2xxQ+5Sv9mTUlbW1Ol1C5McOCnhuIV1NaPEfrQ/gck
pZRiblKtj1Ey1kgmI/hc6cx3bGDVe8aaYPyS09GMz+A/S8ExQcj2DjiUvO+wpTM/
9As5CZQRUEP4MCIRxQxND15RNAvEALnRkU3TskKVoUNan7KipitP2ivaPTRe6H6W
TWDH6OT90cis4Q8iqlwzvodPAIqBwpAxxQ/mKCPgzZY5kjUh8UB/hdLhajni1rYC
XKgOGI4WHHQ1/8BbCYYQGon6N3kZTmw4RnEX+RSUkpMzZoskxQvF2ZSvE1uP19LW
/JHvfgPnm5vYZ4V6nmXtBiRcmd5zve5MKBONQ1CrcRyVq4pYkyimdGBUmtecn2BP
DOeeOjvYOZTI4kc4DI83OK9TaH+7Cu7X/9qR0GMCN4K5PbUZGk4TzZMfNidSx3r+
YeKIperz4JZMWaISIW27ydY/pUOpnnYRIFnXSYh9qqo3IljHCM9zIY2k+aU2h6/N
g/B7hwm67GBvP7EplmoRhMe6y6r9cU/grF2eT7rZqlBapsOgz9qkK7qfJuFIiuH7
1AK0xOb6R281xY7Letjy7rpm4Wlgcw/wUzvPm1aCt5DyUkKubTe3T6EAPtZay+aq
ZHc3nBJTv5hxm+PabS+rNJAPw1Uc0A1MSaIonMgSd3MtoiAuwYppLiyYAsrdNEej
TiJjRoAxXhhVmz61rT8K4kCqot/XiHrSQz5oPgy/BEE51bhLlPArnbi5PPJkOQ1U
FhLY+nfqd7wgubjEpB5ERL3NicG9p5S7QGKM/7wrhdcNyPQLn5ceZmwEU4OQoBui
dwHRvLBIJorHrRHxK2jvP0RSUwvJcKr5/lIBKTPHh9lbb0T2e6ikk+szccBgRL+C
5hzG3nRq7LMPKc+QqxwKwgob0I8uTliPLJqe1DU8Oi7EbLhvjyG7VCKtWolB73z/
zJaa6fmowfgSp51Ujrxe6evVIdFnuuUb+sZuNZWtdiKZ4UYxCDd3lq8brE9Dn6Z3
32oqM6YkyyAsCa4T+pzpb/aYNWVMqvoKwMjCBcZXsH/92YFQvqoyIWqDsaUmmWdx
rDKwzCaOPeAQID4Z23D+Wv48Hme9i/k0I2bj/zaaMwklwKT8HziFvjUNRdSa4FtE
jzoXy2vE4aaWiWuNKHzigvVkF0t7FbA+VYIfR3rsiCZsEZvfgtH0GVn3/RlRa8Xp
aWH507+X8wI2CuiH1ZHiEoj3+UySGCoriiowGmfMRku8wvGYDIpM0W/rExmFhvS0
3xIA7avvInBw2URom/rawIq8nPiZ5aNlu2pRF0R+EXr2GJVh0HQkOTJFYIWWsot9
+Up88b0aHhg7xm+yWGr4oaNdS065pm+gfJ/A2rx4Oie9WmPRNC9W7GCNouOoIuAI
6DnaGZU1M/HeO3PChGG6z8PtRo/bgGzDPWQsTTqPBB7BxtXmDcMTZEuqhV+htRFL
36Qx92BWkGyuatfG73G/g/uDQwxNDL2Tf6qzR7eFz0gE0wHQWtZP6skOnT5pX2qZ
YToffTnJBqXMlwIb05b6dUK+EnXhoT4aEbfeCfNDakoUlthTAdtlXv5ia90nmWou
uKzk1ViS/zu2v//++F5gBWhCuz46zBcCXYoKqgA9o2SWGJuMdMAagb8fq2jcOVj2
mOTRcnq22LwLUCZ30HnEZ9kbxf3mgs7EOwkWKxNM9N7k/kB4ZKcGoAJzo8xxr0DV
6Scjl4r7XJbN7rovBwTAuePNE+t1eE7GaRH2z90Et+9a3eTO5sU8qUD8jvji+0pe
BNEPnI4z3LzUmwukuAI6FcO23Akp0NkYb0rEfKTMxaJRdDHwfM4c3v0b3AQeHRpq
evEq/SBN9R0tl5ZcAzxDoTOLP5HMWowQIxJdqJEbUlXmHc2dAGoNPLER3FUZ1dkm
9lCsRCIyVfbZCvjq0YbI6UsdPX2+tG4AsctoCUPBR1/jzOK6LBWIN5PTwq/2AI6E
ttEB6wbpw9YUDqVU0mwJUgIlsNtDsWyODER9xvMYZrLOVPDKY0ixsQyZdaiUZFYy
nbp+1zDrxH+TM93SO7yjwhdSbCHlvnb/toj+mdBP2X2UpxGEoWG1rN1Sd5WYa5YX
jd6OQ9B4Mpha8JIiVrXV5uD8uAq+hR+KeQGhkM1LnCzFjq+n/uWVA8h7AkY9RGFT
4q9EsE9r23cnNFQlI44J8KnKKUtqqIV2oCosQ/jEUpF438l0+aae1R4sQsP8ERXO
dn8CXyfhSj/7JisWTlhx+2830ck1jGEHP26d0EgbY1ZxH3SWxhJ1d1yR6BYqSFry
x13dDkNKD5mMn2kwaAq/YYfVBiqxEwHD3Z8bLnAuys40JYEoA3PiMyRreOHSHDyI
gZZ87TiZB5wI5/TLrcbrBRzSVpwdIWa39tz0jqARi4sz4ruMMo0z9BWTLX/4cmBf
AYssRrGTx9gyZDEhxPj7HMLH1X8etVulW72LJC0haXi5PO2oCXFXGWSOt+90JhU1
oyO0089eBbNvwcRHqbUytzxFoC+JrNwd0Uixv0j8iAwOuTAqdHYEyINDngxPJMhZ
J0KCTrax8dQhvRBWGPGRvxmzQ3jTwhgsnYR2XDqJEApNR9TJqfoV8DIFl2dg09DP
WVW0xDQq+8HdaGg3Vn+01LJs6GqS6Q6k8Zjy9KKTRtuYFWkvhxbnTzKJeVbTYdSC
W+6EK80lUejwCXZ1GgrLEc7gTIv6MgUfM0ZYIJl3JESrkps6ApQtSnQJyq/STDZt
fl/k9NP113G3GzO7mr9QYSYetSzqh49kwD7EacYfjkV9LEFsaK8nbwHc0ZxT3bFW
woBGl4tBu+3hr6ZGdZNB1dP5V9CGw2wtvjFOggDpfXc5UPfsn83qQeB2ga/afnOk
ASJoxa7tSqBZGfH19WE5HrFsZyoQxc4Rtlj1yUXppVRXjv4XaSNoX48k8JJN/5+U
Uj8QH8bvpHVTY28r5xiyBIHQUJ6DSV2qIZnkzJ3yaR12SwnF81ktWR9CI8B2C+27
qn49cJhv5seQafJ/LiLjBzPMxqb2qDPN9PGRgJ1mfDDWFIbyehCXDGObRlZh3GB5
BmcvI4A2dZHcPkdNvW658ORo2SqsYSebZ4ywHyLxAlAcHiWcGF7tyX/96nOlNjjc
gELSM2eWe55/xd+USsfflCXKFAfIWAiF0TOyXEBhh3BwiE/kG2o93Fr8YYuhBN+0
E8WjNIuKThLLthxGpkne76uu+5l82WNGEfHxi8K2pGoyv3fugUXVmi0ZHDUBpMTk
9CRQuR1u+ss7Oi76BIwZzlNVCQ7DJupQjUPkqCxSJjAIKJDnnbat//cfgc8aJdPZ
0zYvyxYSPEvpCTQrjJ62kdT9B4l5jvRejywfoN9GXhRKyhATUmVEyOWWggiITNHz
ftm+ry0nduAZYg+BwDI4XYhOL9AHua/UWR13HU08OroWcnOsfIdUibSG+Xk1y4od
66fkw5cMRk5RFcnPw+XUOEQzyKflUvkTwomzd4e0FhzpkGUFKIKvFTFUJ5QbxpE7
m3OzCls+4yEkpNxDwCW5uKGG0XrolKTIyonIytxzDeCDxEfZ1ZqBNMR/v81qxqsl
tjm5MEQfV3q9do8b7KKjQi8Ox5dI3FhWOuMmuNPdKjY4iF9SGJYfGQwUQYQrTe2o
i4/71BYBpv+0bp7Q8msdViwvgge8MLiMo+Urhac1SVccjJObJVkSIjxqP5pdkMsX
OujoTtdDz0BuIEzl425HYQQ8E/g0UaeDxWIHvG4EQkdVRT4y+ZorqpiW16sN0+L4
300ZdVH0+WITfGEgbRLvrwqlyG5SfI5AgDj80F845QaG6o2VkaBTl8RrmOsx97V9
VxcH5Nl1FDAoXsrCNLEFUD3Y9Hwj0pfVO59CwPnH5PLs2t5cVrGutj1O093FA0Ci
JQbM2BvCGCQ/R15BTk13CMS0lx737GLuISyIlbi8lJjgNd24Lk1AiH4rSxNTa2F5
AG7bFcB4c8M0TlmPAewaqfxoyG7Ydr+YIWxAM7sDwf/NzXgqadHWDhEcr/9wofIo
qozoTFsk6pvSVGP3XbEy+QIfzpgIb4YOAg+ZLWLDTahuST5zbn+P8IcUjkD5ZpfS
L3ZFz75pnvc1iLZLRSegMKv9ElIKIiDjwhjgrBpJeJLrfizIWmcenMSh7u60HD1b
ciD6UNk1qwXUl83FoGe4vo3dRA2gocFHBP2BOhjLHw1WYVsQaBQnebTQ/U7htSBu
yaegJq6KK8jsPH85+LJ2mXT/0QSlsg4+C/TUiHWjtg3Bk5KYRdqUs8pJ544os99L
K9zNd2StSbF8imd05RusbVOfbdGJbIC0Wf3vXDMmv5o6JaokjX9pNlzwJnwVhqag
B1FN3PDY77mAV6s1n9LrO+ULi9iSVwLK+TvEUHgjMm3dG/Ux5RuFr83PhkdaURKn
lNJoab9/gIHPkNPiomfrQFAFqYyQznScuFdBAG86LXA7rG6lahsVA/4AvO8mFOgj
BvltdUBfAbfjvUXvw1Y9QRofkAufWAKjr4tPKG1jNfKZYvhvHeCOHg13jlmL5iC1
HCOF7QdMAF2wdmCo/3KLBn2bPkgDLYmm9mVNXXIQF1hRpf1SZONRCpHpRehSQb8e
hKXodCHyV/BHPW73aMnCapFBlgmuTEQ5EmsBFsfw0w3FpraJKoXJUcqmjNtV70Jo
aYyuszeAPIvYBvNOOtmUmK1X8ZuurOqXsdXmm9OtoONl17F7evd2EQitGxk9ICdm
5myOSjwVcLhjz0TAG/BpRj792cbWN0fxuNbQvqaOuNJgRsXq5EaTWkDwRoXCYwg1
W2T9AuYXqaTiorp9qmJwaJMHm+gxsIIEoY0QZUdsabGRyImE/TiFJ6nhzzZI4JSn
vwXVwMIou5JWS4q+ZHZe+i1YY9ElhI3dfrXJQckrfMd0XU0MKBgFJXA/zLhwALci
Dv7l9DQY5bBHM55UAeuK47gAALJ1T1PmVIWyUhSmATU5vebCS3X9pf6vr9iypIAp
AynyFevZgmMIAfODN6PViuaNcTqgfRiPxKBG3pahPqcbxU8bi0SRwdztO8w2bXK8
WkA8e18dOoeTSUZ2EMd6CEod6tMG+SccHn2dq9uK86NqIIK0ic9HpBy0+joBmjXD
gGd1+CeRn12TC4qySEBK9NFA1n+4LOnOZ+lhc7RSxiVuPwzJBM/Ito2J7dJa90M1
IjFbmUlBp+wqX3CRqAbdWrXV1V7FWMmOKpHihyVwsey9Dxc8/1+UfnAufeGyBpIa
UXQ32HzLzlJoO/EIKRhZbYkCUxbAT+66y5SWWdP7VapeY3OQTESzOABXnHCIgr9R
vv6TcvpxBfMt1GoFoq23vQXSyj5OniOdMn2AjMtA8K6lbTIQCsy69jvJQLX3fjiM
L+JR+6lgBbafkOYIRejm4pvg2tfFOwSgGNk77+o+IZ29zMeMtfw7pd/Hri336ysD
lja7Zy+vvxCHYumn8XiIc9LIxXOd7wKF15Iv/VEsHMcscGfFpURKWwbRqzl+TH7/
0eVWar/lOgt0SScIaa1w5rWmsZczKwEN8pqHRPl4KZkkeayq00e7BS7I95LROdSn
S2gZCksJc9dKdeNSAl+owoeMXxP5Cnx0E+slHPuDq++m21wUZtCY281C93QnS74k
CtdhOR51x/og2X0AdVphiMPY869JcGRe6iOjYGOBXOrgMZNywelfts5Rs/SPasFA
cxXGkLhsXbR/vpg3ZE4fXxULInvDH6DzYWFjjgaNGOdaOY2TomCLk9sH5gnXYkcO
bG+jVoeI43vfvUzcaLmwQr2LQGh7nrwirsRdeMomnfiTup4vUBSIEmrCuK0sJRl/
wUWGJ0o9LRNts6WfUKRPxQSnHcSYWZIDS/Az7GjesvdQto73O0nDYVJDuHp/56g2
k70obfzfMoOlYSl+1/RUW4MoCjTB5Jv86yhoS3BEvTe6I/xiYB/GHGtNS0rjqSad
FQ2LF4IOU9UCtlzMkBv1yG2mJQ7rTF6neNf57PsxOyBINRE3d/4+YZyJEoubIHQK
1TlqeW5SpyKvXVi62Wk8TINu6SPo68JSRcc3RzgP+P/2bchvYtyXltz3QkH9SozP
oc4aBQPOFjkmoAsvLy0QrgyaEgAbFD8glJcVXKaECDkGRnmrDtGD0iHputIb+UdD
Nb5RM6iwHerKD0I+8IOltAvFJR9rhRXQrRyjhJzMmgk8jLCoXtKqD14maqppTzIU
PQojBxCsSk7tgEHrz4Zd3RMuaze/FSY7gDBIUliNJklXHemrGs+UAfL0OpBDKy0m
SUDANZSq4U+Mh5ExnxeDah91hIM0xtIWc0bPBsYyxPx4fd8hnXrFi/uGYzUL8h5v
DvXkBSsusI4rQcs1uNFbIUm9agoSgPTnaCuV/dGUuaWZLze2spTapKKSMAxLFCTq
ncpkvH6uuEjyWybrfJPVsBSUaxaGxZyWQKv4jcXE8if0n/uJ2F0lQUvUjDpWe2u4
z0O6s+6+APrd3Bqfb8KanZ/atvBLcqq7OyYTNfuS65VfDa4nx3Hm18iFTLNPmS0b
a3zwmICHiG8YOwUKDTibuWnH8kF1NnL9gkA93j9FMAqodHGL6cl0S4fV3zlpUkr7
bX4w/mHF/MWgU8XvYbht6zHP5o+LWFw72daQpophn1GXz6hhogI/BQL7+/A4iax5
Wc8aIdSk3XPgnXlTPJFtH+zVlasp551z56QGW2UGilMGroMOfBDCnLnnHkxHjZ7E
VT8jSuwN8v0zeO0nHBArfVn/WeuVGNXpj7KD6CnEypVbwvyIgZemPu932UxJOipN
WIrH6GvVk/p65lxcxExuBp0bdsL2GI+I6/ZyjJ0rPNWjW4CZbOoUI3oW7RblpkH7
yHGKvPkON3w9VCVKxD2LOvXAlvgOe7xRYD4z7KE7Z7szqfqNE4aIoR3tUZk4BOAx
h+QW5Dm2g3+500OLiTJLetCwYD4//X45yPKMl+0AW4chI90CexZgljmPKum9z+Ac
FIqUH4ecPCbhEHauVqUMP4Qh9S+HR4uC8Ns/wFbJumDUcy3JDD25kvM7PtArvhG/
skj3x/IQ990QXK0PBMFP979XKJ6st4BeCFDdeH12kfKZvsRZ92Mqb7jqsFq9YNDs
n7n5qh+4lal+AWgyz/3396DW7IUhv/SoKC60MrREHCp95DQpQi6Jl9zkYDHVUTYN
twNYvOHAcfOxSXrGY9C9eQvqocgv48NXC41hf0yojotI5Zjx2HwIHzMSCfxXKxfO
o2p+tW69dmJoLVKh4E47T3HnQVzaCGYv1zvh/1wpqXgUACiNnNcX5qUBDYngCiJQ
fJM7pegh9t+gc7VNMK1IkwxaXxViO9liQSLJ/58gL+TgD9fmp6nM4R21E0bBaONy
5/WtrqkX2Zjvhljs/+eaeSMpBzq8lFibXXBVF7Aj/C0ixXfy9FlP5/rCnd0MPWbS
fLe7HoKOGv+icI9KtjvpZnW/dqXHC+Wq0IescxwJdFf0NH1JAiyzWp40H/CVERME
GdIblMi5ci0WU49o8sy8/aggBzW9JbeTDaZAVInJhYPGz7sat/ORLatVuIiZQIkr
a6PpnablRhxE8u2uql6SgLfBmnwKuebaxB1dZUjgyT0ImaAP7BPO7mt++DStAPvB
dqvhY97s0FxxXltYmdOm/wTEwRxEUo+aKEO0BNNPc9aUXA0yPtOEmiWX7MyOfDYl
8mC44XmEyoRHq/t43l9OwHaNDRwoZPAkhyNIXFOLVRkILdG/L0S+fMds+Kn1WV+0
giXCoWZFQEXBB4f6Lop413pwI5yzWR+2ZFyMdNRaLod5DDOmIqeeKixVPayyE8Sk
XHJbxJgwxTWJry2JG0XSxK/yaHk+lD9bSEYkIKRpFd+wE0RZs8FhOxgtZL3gxIxE
f/sCkVO8ZHLX4TCsESgktxTY3eWf8gCj+HJxlgybJqNBF6U79ENhWS3YV3lQ00xp
QCH1HG7fRvZcb7KlD/oM42YY+ZK0bKr4YD2nnkSnM2xje/Ek5kI1qbflJjjoZdvv
+3CkhsXfswaFKlWVOobAg4oy5ql1kycv3vT9PqXcJ9qoixUhQQdfBO1igtdGCRTC
ZWD3YwwkCCtxs7hTCc6vPDGIsS9w9Lav3DMEI7bYAzgLg3gDEbf25YaG6MpKj2c2
258R42+MmpgGnPeIAW0KMYENtKFWK6h1f58AV41Je8sV1FuGmatdwGLkg94cV9WL
jdgKx7Oydz9gzJFbuQ1c9ReJczUF9FgHpjfRe7SzzNQPo01nVWcHOh6W7IO4BThE
eIk2Qb/UE72flSg/3AUedHRZ2fAfoWQlEeRjN8NV48YnK9q5O6JR++S38glJYyXw
XfBNb0DWbOlXcbcOhdX6cFmVLGl9AMJYvYm0HpOn17uBaWyASwEAI2ZldNgyFUM+
p+wnAfjva4PRFKrhjoylbdkVLJxTr/X6oi+RhbIcn09EBZzrhxEzCaITEvqjHvUf
HKhXOSHLNfUnD61tEXS8hGISjHRA0McNWytl0zj3wQCasdsxtFqI+ioomI0UYCdd
OVwUIBaPm136W/p0XrOhXERpiHR/Cu7+RFTDYyFXJMOmNOkb5AZZy95WpOplJLFE
F4PlOYUuu2/gRyRr6CV50WPpWoSZnnst3v9N+hPJqtcHWxC4AmAPi1yUnOmk1Jp8
EgZhYvPnG/oDZh4qFVNGhbFbXFyA9xrcqMDzcmBSOaMPsF468aV9+l9RQMsfHsqM
bgFaECSygI2TdUdGjcpLNnFk1xkMWFPk9lYHCOLk/r5FihsXRc0e8TcUWcMwV0Z4
Zo7ro2NP3Hmwmetvvjze821IflQzNCZCbpgyQJXaE7Un2CmvrKYFpVXCeILVttbJ
dwv7gMgovjMZjvBHRaemgqYwDtBhfDvnKEax9AmhMh20Itnt3InWgo4NKkSY2/HK
wI+3afxKNLz2jmosMvpqAo4Bl3b4I+rdRldL//y0KnjNJ04Oe4g0fN/qOSxn3KCz
GB/gFiAuz9LHR4gKz3mF4lAC4TWWBgdq04eD6+lJ0Na3vo9JZo9XW7C0jzpr7oMC
Rs4o9Li73WCNc45Ieb3uhTIvPwYmWTHfnpPIl+dHm2BWS1KJDqZoEZX1uiMy3noU
mVKjSiZLtHMpLLUGt2nAqdphtEhGEI3/bKASg3IetCQFwzmddTDYkZO9KzPFkhtE
+he75KssfIxq0k2R+DlGXrizUQsMOTbYNNRR3VdwqOLNHe8xR4V0vVl4awNxJDUj
scTfvXpZDJjSd9cCwAndxkNw0tv3SUIJ4yCmJ9JrcfTug1LT5AqCn58+1mY2p0hn
B9KruRfZRdNqaflEQhV1cynJDNob2xiENUb2xPPrEqkrtBu+J1UllJGjETqyQ/IV
3CzYyiobvHBjDZDMDvjlMaQSCfhTq1Y20BRFRr34EXdU2EW7g7G2JWb1UqX0RAG6
NPAkwUXU7mM+dm7Jg3ezZH7vhm4W+Bc5fWVSu/PjTvCI5G/QZcgyJhrh1RHKSKsp
j3aQKPtwiV6fyNsP7fGW3sDBIzQvrPVSv7+cr9IYCP+lodBAbLlMGD9laKotf4S7
yq6QumJ5AbGdDJnBC6f5QvDN6W77WGQ5CkFpJSPRxMpIZBH2C7Ndrx8jv0/0bAky
p3x+MPgqIYm8pD6XojrWWD5TepxwZHkmqHBZ/ghw1tpoWwh3a4T4oVEJwjj5J/ac
yjoG+lHIL8Q7Be6C4G/BZ0yOfofhjJiumMkmRLxsyqL967JjI+H7SqdNQzeD5b5z
11u+qHYVA+lrLnEFUF5T00j6mUa/aGWk7bgQJ8dDdFKTk2bh6b0lqxuG2Doc4oNH
6f9w2vGpfa1FGJjoMNi1isnY/gcL5VYCTL3xm1xP8hZpjsMcgW2PyUgeCIgAUoAO
wnMR0YEeHPUTZ0251/FH7XXO/CJC0D+1asKVLAa0DfN2Z7BaO4A24TjKSViG1LtN
eCM+nxu5K5rtLjZgDeGgjt3S7sGYdiPh88TSq3QMGUyMLohuC90LhdbKwGfQnf29
LsZaecoiPjAVVy7hC3ZdtCyhhNrFZ5JQBth/aolrJ5FHG/GZuwxieW1iC6VdMPWo
uk9XXKI3h5ehPZYG3pH0SkPwY3LeP7LoAu77DbW2jOy8jE6qZpBZXj/xqaXGcYtG
vBubB0jlY7yuq9dnigX14hGakgks95HN5dDTqFBesHpRn0kU7MJLjyT+uOoftc36
WibI4n0LTKnZMsNZJRLDMnYGeBesQBhXBajeqVurPC/BIJWel7SbdS1zRPN7Es5t
R0Fk/vi/AXmqiPpQKeHriYpYnvQZOkoshhUvIDTvcE5KSLeBBziMvZ2LzKniZ7Ux
B2J5F+mH/DHchOrxvfMfcYm+NEtXevfQ4VimaPgTQPLUYipRJ5Y3qxgrLDF05j7q
WvzyiuqpmOygRmgKoGlxJYNhuwx7gN6quzjZ13qudWM+bqvOaK4WUPJ24TfUusuB
IZtL1YduwZ6NA7E9Y48vmJivaRo7KGOB74+UeHEJP4HV0YiQZdjZI1Ik4SdPjAaS
v524VwOcUaKwG+VIwRQj7y6iXpeitoSMjIJFkzth8SANrPs5vrqed9NS4jA7KI11
YUgtLPQqc6drW/zudRcxLewDZDq3rAN1tHa1rnsiWF70u4NIgFQyywpuEkVtRP0k
4j6FLLbWSkY3dLLcVJNEmi7rMgwkfg2bNkQEjiz8AlJJ9ZYfHox8MV6lqKs+MSej
QpSOxH7kzzuhnGwFs9Aou58TfC9XVJ773nh6z3zEYqNLU7PnYQiNNp1FALVK0OUx
CAJdfhkzq1ua1JYBeCb6eZLrSvwq1Y2s5QzKpMflja6mvZeD+HmybLrid582WltQ
2E0CPQB7ZUHcWiI0gPQPxRK9G+q7b2Xc7vAV74sVDzIak+dHX7EyfdCQYwJiPC36
1TKQRyKCfiJZWdpHaEDpydC08e+p31FUxS3R8dvGYxwIgKx2hyWDVLPRxx0P/vlY
QrL+2nACofrkg4UNIwQGs3EF9Uwd22OuT8CrTOjoRrQnlsK7aPkiVf7Lo7fyne/j
aL71nQeQQlAvjqI3hRJA4Yg6gjQL3NZ46acEwqNw9tSjFY8jDsWD+3PloHL7sCre
AkY32YJMl7gfhDMwZKqGHorK25XbHLNvO1+/oco+mZGZo46EdUnz0QcsiRUb24/n
WGPX3F3Y96+ly8/TsGRC9T83AHv7ue1fdsqc7hip3mKULga7wmeQGtfkF4Tu+RMc
qRVmEKi3ZPFY0fRfwL3v6epAcrH4skHRxRp87Qt3Z60TtBaClXoD4S/2NSVNEXbs
ZREtVpbPu6i+nR8KwliIgKFQanjvyUAaqXLAplUV1ry/OZH2KmyZM3W09NJRmQCQ
a4iRaTrK0QNn00Y6qjq7Hp89z/7e+dolgwmMTQ07flDRisGwqS5uMhgr6E1xwnnN
gzWPYxkR8Hiq8+P07hDLElETIDQOl/fJPe2mNZNEGUrmByjhLua0uhhQuaO/D6ga
xd9JEnGqHMFq2zxBQy+Y1CGpxiYQ65Ilh3KHe6YKaKtbNSxFmFtrw8+0WDHliVrm
IuSj9zqXLNa5wbwPLTtL3ZHVfeQ6nAOM/rp5uT5NAqLb74n5VKHKPHwA4rpzMGmC
393pCoGkmOTZ8ImX3rOMXERLdJo5cytXdk67C1zXVOhqr5Njq5b00jr0m7yxvmyS
yacDA3Fza+XWU1/Pa0xfgI/KjwcW3YQnIcHhF0Y+FggcvQN1w6PIejF2OxELTsuh
X2Z66uzOdW1Db+eeEBzuOMtgQC9rO+mowBgFM1PERgcnrvfX5GkOM52nGa2Mjk8n
TaJty8ngKU29ONejfdY4gTcoKmWrBAJtVNACzTZxlg3uA4WufkYG8dgniZ9YBFNX
0iDJaNgOGkv0eK/mFbQp1puZnuePCzndZNx23FhuD72694BzLjlwgOVDJNs1txM/
aW3n7hPCbfmBDirJvtXFW+USVXs7VCTvrIv5bRnZRRH2nbE3LIVTn0ikzF4Q9dgf
6kNIB8v9hQCwtTrO2qvm9bAfCI/tgq7HifGKD3WIemGgA27OlRrphjuABWfxn40L
FtWA9sW2Yn190kYBs8iiogsdnC5FalmiqZ7trQ2WqugyIWBYuxWPVkuabucP5eru
FS4+9WLArqT/sVretlihDZp/muTEb7KrQ5SeWQJVkZnOSWcYvVi+WXtyTiOKJWht
JhmWWh9dhODdPukHlZOIQadfYQvlFRl5l8F/bEZwr92b2ULWfRl9fcoCSEtQRbZg
V8Pnaj85NxygQeBLU23ZSRdyRC/jXu746wFRdYPl8Nh683fHK7fXcs/18IUQtfOb
7WyRyz8arsZeBzobKDPA7/zcSxlWX+xsLwfKmAgvUu1UJTFMbeLkfrpOrGa7hF82
N82Mk9Txx0Ml4Tl3Jc2j0coZ+JL078PL7UMCmcaxs/kVok4uc1X1m9REKj4SH4OO
AChvRNqzXfdTSEGquQC9dTzFPWZ6Sfr2vYy3hxtd8P/JxNVa05nYe0tFLTOReCrK
F8+GpbRxx3F2FOya757om+69C/QnsIYhIHEupj2BGvhSBSvvG/lU3EN4jqWnt4zc
HR0/h+h8goWnt49poCeCZmWV8hBLg0WdY1oykubd5GspRNVAxLR45wsWZ4W8ilWL
z737m8QyLsuBZmrNSUtX3hv1ylW/oes9ypyOgB+d257chStYRoVlugOC8DKqkqVI
g4mQkVcS5cHt2Cyybb8m1Hhpd6VLpZCdBqvABGicloGezJch4Tmn1i/W5M7PUKMC
5gAWOLOGaIfDZS7zj42zs5e8ZRerXeIqq8FiVBVazuhJAxJ9G51wJ7vAJtJTETBQ
3Vbu1j+v9/aJIKjPXV7RjGpsaSvWsDRbL1QBxFtCwwaTMwaMbBdf0bd92tzFVteN
OZbGjf//PdN2IRhAgufbeJJCnDqCW/hQXK7zI/B/Q8NLBqAkYDcbZjgxTqvnz4/L
hA5NZmWm4/D7/XckTtK8UM8bm5SkfZEapSx5c6FR12UZ+UV34J10kGZmdnJh7k9J
HQs+LqchbanoFP0Xce9BApNCmqkRM7qbDggMIzLrh7bJ+VGBq5pj9JoN37Sum3LE
MY8lfejSxX+L2iQyJAwG+3X9pAftb7TrLmL+2WNXoe8ODFa/QMwLtQS0qjCGmn2W
FiF9WAz1kc8FkIbmNPYueBbmOBrd9AjninoLnn8QLnmw7uJ7qIXy15k+lh/BKZii
Sj2I62Xjx/Hn4htHnmYIAiN+dXVm8hws9KkfZ4yxAQZ6kmOwW46/sAx9RN3dJHaf
Qjzk0cfNSSzmvJhwXyX3JTJsy093CCdR6yC9WzkXPd0gjcdFsQvCvywvsSFGYnpk
UyyySNjGk36PCwxjPVROePOLOJ/i4SjxhwCv1vc1yd3HobERgFxLDv40mRZHHoLz
uoKdwQJrB5BdcpLc/nLmXVusWv0wk7+76WLPwG+pPuk/k44yMArD5S02B0F5syq2
r//zkC4fa3IOjz9Dn2hjBpjhnvEf+Ejxe2iXdhZYeYEMGDdIbH0GlVf02UJUnGtS
G3bWUxEbD20/zyMYy2burufyM8lm0kxlbkuS3iFi0WM0IZnrRgeeJPrRFEwWKwe+
f3dsDXM3+BtAAXWt0nOk7fLUJh9G8dFrSmXZJrtYBTJFOCxkCBrmnFlJHUX5R7Cv
xb9cBANz3rBJbABD+Ugmy/vAqthP1+4d+B+tIDiYl4WnWdekfL0ldzFglEEcPTEj
7++Pu3u8F3VvTDGtX7PrabMYLnNCj4LQZb+BxWRQnihgQ2d9maEARnEU7sgrtjKM
DcPBASlTXg4R0RhYqozkmFa0hsIywY93j/oGTpQcWRgjBMCeFd4XNsL+5cDDRQxD
g/kvgdl6xY2bmu/q5LaQsvjYV4oB7Gc+PSeeo1+r5eOaZ8uDfyLj9U29BQCY1gvT
dceAYajYpMHxPvxdEEwfvzTJYzv25IeJEtM9oNmtzfhvAVlBS/56M739bxTp7KYW
k1RuU6nZDqiHwRNgHRrv+xN8jf8JBvLOkFy9lagUTlk4dvnYaakY7fo8SOvDYV0U
EutRG5gkFAw6f7vIE8WJdAIPkZ7/w0M8+Erg2NwKXs0Z+vs8Ur6mLeoDR81KYnx0
0PybIq2g7AbCPiEyHmB/ZRtmWVx8qMDGlDsPd991qgGCrKvkY7kVK5BKdIuZxwbb
fCNK1UzhB9uOYWkmxDKFlQKoWY+YS+Lo0o9LYW3ZGDFJ58kk9qyf7hPszFKigVlJ
zLLfp2uJt2t3N7wrAE6qC/jHUFB1tYAE3aEpSbpUJ1pzPRi1nHdjU10Pm/aszdRK
pGPUkds+GHW5JdfyypSRHiOZLi7l5eSeYeP08sHZ1biisJfXPRkAIG7n4ZdEiWOP
Fs0hpn0xNnGNA6NMCYrflS+WPy/S4zDJXEjeHvYoWz/7zslGtTS7j5UKZJTad5Qf
fl9XjMp7poDRW6ShfMWUHi7xmzkT7Xb4tCV1ZS2paEjqkbd/tTcMuoyItH3KTLJL
72EmI67kJNo+3Yfp0aBRbawHTZBW0t5mP7PGacvf+i2rs6TWcndaEMhXYh6L2Fsj
jxK+qgGJBd/XmiTbdiq5yXeCpNNUmPNTrcMTmpO8cnvVXQ295CiUABh8tzj7k3yQ
Pj3F8cJ1PJPt3E87T2xbUzgdZqw2sfAxWa+6pgIozzOEQA5cg3vjH0vPp/ccPi0z
TZlUT3yHDbEHy5x/vnvnfAuQpJBraEO3xyrRrtjSKqQb5HcQ95XLOxMO4INKIJeI
xAzkyOsB7A5AUkVhd6mk5GX0pwEDu/bKBxwfsgkgtu6mjP3w5GjuLbt8NJuA6zdV
+SGBmabi2z6HwC9hMG4cuysLsth4oDDNwg4mxAuuDmOsLB5CB08BflBEXXWWUoKg
p/osmRLFr/b0V0no1gy/ZhVzjRWaGv4MMqOWVBLZbAZtpgQvtsf2VxJ5bkUG9jG+
bSpTrUS673zz7azfjLBjA3B2ExC7wOb/mvJ6ET/i0wWnT2nMD5fGJ045noMS3JQV
9oPfm0KhRH5rxOKOuiyNpnXqQuZiatFzlT/kr2R9LQRjhgmrpSO3JOse21pdRxpL
cgLFEtcccV2jQ5aEMVCNE4avCRvasxkwIsrE8RGPt5/b8zUGrFo31D0oOIPPUB/o
MkaJ1MPwR5fAhzAZCNr8sfmZ8qFSo5XL+ioEtsVlMIMnlyBUn1QurGq0XJ8ir183
YIgnBG7eUMNS23nVcz13p9Kyfb4kmSMcP2c5cSrzvUjHdW3Vc1ZmYBB48+/zCZcV
Q2A7WxSI7YRlOlnumvB7e70tfqRmSul8Nhy2E0qnK7OYuS16Rdbx3mb6DvvXKvua
xYX6nfYO32n6dQbsQBrHIu8PBf1wl4CrbnrLVXCXu0U9MfYADHbfghOwEZlhNYgX
dBXW413lyvXT4sXzgUziw+mclDJAgEUp7XtXz7kdEJ1uZuWMlBOqf0bCqnow8xqT
FAAbHzfX5FRIDJIxg+mp6ZJBifqU23CVtUVQViond66aGlHhfNL1cLhjNEThXsdm
zHwHqoYbuo/Vi6T7t7YdoVBAtLYGvH22Aqy78xTyJP5Gpml4Ah6EDFLqqcSLwu9q
cLKD9znBOgJlb5s6v5rhCGRhivoytnC04i56BR/J7f/b6qH3NvIoCxskk6dX9hwJ
PEkjxdPOTlMIoEHDaExee9DW8mdY8yTwQM4oUH158O9tnQknEXo2my1Qus3FgFr0
JU37VUtXJJwCXRyEhG4PDuA/KfbgGJ01Xh889XvT17YLVQF2Nb4syHx/+JRvFffO
PRh2IlYBdA1cZHU99VDzVsxMgpA6sstPSRP/lTRHVewNR7Bvzy4Gj4LRgSMVECt4
evocFST7PDsYWDz7tKGNGgZPVxI2MCX4ptr7YIVF+bTtlgEV3d96nqwtRq/hXtRx
+Bun1ONrXMaNMOvpzXN0HiEgvJgIMl30PBP2OrkP1GE/8GIRyyzuRdnM1g5VlHKL
qbAK7FieWGs9qvrJnDsdr1WKQ8oNveh2b+WuraZBCKqST4VbLV8ZdPCek8TPU2mF
d/P1VusV8JJDkrDgdbk7kQwg9wzQuts7Vph4HD1q8E884Z3qiTxtONS39HqWQx+i
XOjGwM+Svc3WDTeKR313R8/LimWAig6RJqU9ZDje1jM2iUm3OJXE0Lm1GUpOi8un
MpsOdcVaMStOa+LPH9fqcLgbKq2mcGSwrBUE1qv4W8tmVWjBKtcx8AUlHSyN6rNY
oTt1KyJneJDzcZ/ecuum3eewdV8ENHuMyueNPG6TZFoA11BdG/Wc8mYlgO8Zz/aM
0ylM07Ep4JSO+Xu6r7nVuK3181lDr/INyt56lz3MSOWHUMzDyPQSttiGjk+mb6WA
fr+91nfL5VXYMcKSkgRvilk+Kwi4Yp4oHvBFtfKz3PiEEFbFDSdOQMUVlqbufJpx
9VzPVrU7oy6qlifmo1Skv6uUgdN2kIJU0Xb7KWxNtNMOysv8W5WXvuP2V+wnGE3L
gH5/uJekW54v1Ny5RbteQThqotRhflaL8wqOBb3n0V/+1snPledOZtdHsAJZviZ4
BpMjR1tIOKYFZfKPqzftz60fUFMvs/Trfce5AWo0Yrm7nLwIepQ68mfvQzYgbDFP
YpdYb38b17wWvPQryEfB/bw/DB+xHYNJaiPz09h8luxnkk8o2MIdz+57hrw+tdA0
DG6jSJg81CQbYMUaYuLCatxNglvYxFB7gjaarno/D6p4aHCPjXd3mWOA76ZsKCb3
rlUO9sePpkaNNN+MAujtjGpBNt2y/AEtCCHzMWrK7/O94zeGVwNsOb9UiPDR6wWs
POY3wDnIOizkxKyYu0Z1Ibl18LdoBhu2XM4fsC49RXpNywo5rgMgsddFGTzC6895
Pnu4bYVl5b4upL5b3ZIzqVXtgmz+KxTQaNV/VY39JTKIsgX5VJRa3GHGSFPy3W/E
Y93AVoZyL4Od1qHd/vgVcTMCgkaxP6fKvVesvUtbfe+5CjWS6K/ZV2yvIq/io6D7
cjBFJbNXxkcQqA+3Srf1y8JswCTI6DHYXOC/5i/zwnRFLQboGSSKFhMXchUk3iIU
zs58vfPCwl1AK2hZNuqp55WFBcCZNvByu27dVYP2bJZw/UwwOBSNuCw+pweV4N/j
9sf4XHbFdyvJ6nZchIkclAFJKRUjMXX1VdPe/fkwHALPkinFlzkiAOdNTapQqDTF
51puZRUtR+UQ9FVBfX4Nvwbz9qFfOamOts9K9vKBjZuqSR6RHuzVOPNDozerT2sU
r+jNhWJsCrpLBk7PO1D6JSTaMiF24yBXL6LUELWwSWL85Wyg/HV9zUgGaMJp+sL9
Kf+Ro8NUp1G4MLfFKSXWZVlAwzskwtkWPJExnk1YbTTLTPboKOWNC/0OD/nRm8FI
Td/bwax8a2vLh/KYCuSH89O9oRtYVJWezoP/uLj5xrYjrK2BhgL8+XMH98kbGy2Y
wqVuBg3vtwHy4xBhJ/aqclSRAzdnznRdgk/FyGyE80lUU40LYemxWNC/fj3G8k8h
IQntr9f1DfBv0C6Sgz+jN20FrP22KF24sURbvaZq9road3ZEoIvnzmL9tyy57tPT
bMh6Bcz01lRHV589dmm1HxTPf0VMwxuD8R4CDnNODU8MdxijumlzMqzW1/IqgiQ2
OEcXOxgTadYoQsFeo3LjCQt7PvIimZOUNgbs/wA8zSL6PTlOoxWQxBToL773n6Lg
KdP22C+QcWyi0nyn+e46zkqta2xni0gJTzsV4WZadqR9GKVP6IeB3MCa23tmpU7L
ted5yJgTQLk80aPMiOKNgBfswGG6268UOOTWHPZr7gaWmDF7M9iykUY92hTi2Azf
U7e7+DSudEq/MPivt5QDjwXWirShx9rRDNEY4zZSjAtLWHD2utHh55pa3bPMsqtA
CQHLnS70J0wB1BBdl6pL6J/1X2aAKrjwaMP39i4PlHOUInKm8ymTaYTSg2c3uQQB
9lB8lZBvV2QOL1ECXgNmf7keLLbd5sbNj2V3L3/q2CVHh8Z7V/VqSbTLm2sZ+kNN
fj10/g5qCnzy7rq9r0WA9uwV927Qn8rr4BwQRXRBb+K/1mWZXIUVhsjmCxjPGXro
kT4LZhcuDncdHgrSTuBD6a4/FBDykshd8og2zHs/rs+50pI5IpgJNwPBydz9NAZP
+5s17qyY3INo9WEwQKF1GxEgQrkrtJRQ7HqGbDHCcOwWyM6SLYGA3/TYWl99yRvh
uePAqnKFm6eDInqq71o5eXfQcKrxd/Q8oto6uWr07Ei84iZkThOhqilRjkeruycv
qlQHADLiDBtp0pFTe29SrXHCVzPxQeDfyvSeBStuek2quuZ2seLo0ojek9noDTnm
FZIdJE7bgNFT8kIHNdvktPIX4n229LNbI0WrlB3DcOos4nnUhuPeljLgQqI5nrBr
v5LhB1uljRLkSnqwYvJeQspWSy4ynQB9tr6hUAM/WG3RRoAY76eUxHvBNEws2w1X
eY1Woooq0k+BSMvEPLOgJmfzbkxoGkeDSI19OAQyD9FqQRQKlb0FBdswRH5r/cp6
PRd5vwXRNRObYFyzghlqofLTVJIzMqCKyVCrdVQJXIl4NWxWVPC9UXo20kCGoCAV
PcxfWLvzZFLSCu0Ld3cCwvA8l7ojU30joxGhQkahCl72GBbkbWgN+a0iLaGRgDC8
pR9dpXGpCte85ywxBmcdRlpBNP4wFQi+T/tLBsDzAxfzN+9MruZtEAYLxNS/ey48
asZntzKi223wtLLxrD/zWGxa7K6c0gM2NiSceKWZx578hZD/FavhJT/eoTs3FJf4
6umBEwSmuu8iDA2btvmbn+8OlvvAarC5oqJB7SYLgnipk0ukcpGlGiZBxXDppaTO
duihLtgmLRldv/IcxDDK0T+PHSxFdjPDbVy/mgb0qRUj9lDeBWKthtQACoDlnVcc
LaAS0QRxwOGpHSzIjeh6uXjw3PUKWxkILqkbJd3abguG2ztDBMeafWJKOjK0sSfD
67s5psJjACoD9rBhpAYnpkAytuqf7ihyc+u87z9rKG4oYHrVqoxeNZd7/hPAPt8Y
aJIg1rRlI0MJ+xGBQlvLRzMBq7VasSkUHu7XjoPXhPtLI4wQIzRYIP7c1jeswnog
LoqAJlcaEYE9Dj7I/WYz6ueWbBdXnogQj9zgYstcyX75i2Xb70mgFLTxVJZNRgRN
1mq1n2ujT6tvGZL1qA+b83yupbb7dOkjFrz18m4hBNWBW0wWxC9fg+1GqNqtqaDO
mFDU0OPJWHdWDj0ByyVudSRs8gJJjve6c7kyc9xXcU5B7ATefxf6KjnssVvgd6a+
qrv0US3Gkp3q/VnpRSN8R3eycjSAXG/V2SeH9hEYJV3CqqCxoEiHccXV55naBrDO
zAJxylluNM7t2+LO/wg61KGL785DvNtFrj2j8OtdJqztwEaykfRuY44fyyqVaJaR
QeQ3Sn5RkGeXf5jdjI8loNCMduZV5NJRak8iiGtPUSHVXurVLdYVLe0aeieYWsvU
YWsWboLtFpkCjgC4YT8wm+wrg57pUiWpKHv6vfy7fWHXoWL/3xmsEwxqQ8U41Nwa
gpafFCpBt63KfXZXYbC1p2okf9Fb1kaq1KJ2IqLVgP6CwRoATZKpFfppaVPBVaiv
nqM5pAIlkK/VRjI06FKPedL3hITg91lxwmUXRzo3KIuY81UXRs2vrPEoeA0iEMd0
eXuUVR8A9NAc2w9oN2EgfjgNqht/rSoG9eIhnAAvj9aqns8NUtqtkARO71+TiAuY
4pw3ru6bISXoit2FGoT8mGDoVO8qIOkVZo3MJRLZc5D3MNj6dKrDZAT3gQsx1bHV
O0eb1F18o46NuRCfg47qYmRpKcjp/l7glds9GyQRL1Hmf2PkORmilQfgKyE7hKpl
puwcdi4gj41oy3WfYEyv2xppx6zQdaOI5zHDiP4SDAlJU3kpDW6kSieTCU58fmDt
GVOD2S/y83UIb9vuExIOcKkB2uGeLhhJAkvHG5MCGkkpZmcqYCnic8/zRyeOPk7E
3gc/HmwBiqYbGzjl799JtUrIiqUk9tuZFdP1Wlo60c2myqQlhULgHFRi6s3UjKap
vn2uHQiifCwsCqRbmt980GpGDeQPiQNCdgbnXA+YnKHNu+KH36ZF2me3WHDozsvR
F+nV35M+c0581lC3bFz7Yvv2uL7Y1XFkbB4n+cOeyfMjVQDTwK5r4FQp4kPJYsXT
RMBkiIEUp+1m46MaXlZ68/1eoabhPUU7gZI/an8SbN3tgU+xq2xgXvxM698h47ho
C3WrgtkKUQ8V7gark66YV0gWcQmA7j5yV93MkYeI8ArxAD6BcRqBgT0Hs3gAHtYX
nkj+AcWMcvuIdDbyZu75nyzhXKgaMj9Xn0zWFqJqBJp6MnYWLtzayrjlGz5yDaMk
uk0OluFw+QWOrdpNOa1bfPEbsD1TWnqDOZm3rcehsTTFXMJAYpfO1+d4HWyJvIRf
OiK3sdBZKc6dD4XNq3l0FBX3gJsJxRtk9Gr5cCyVVxIFGp1G6uns81RmvBC4vC9K
5F3AZG05VJ3fsFbEMsgGLr21LDrTKP9BUhnzqeWORv+l+M8C2oKmlmK1wNz2CimR
3fEIwtZOZloKAa/HRiNOlfe04O9twcDfBJe5PiB+kXeMRQZ0w1h8DVN/cjPOWl66
zaBZ7aK5tSD9dKlK5lcCTMUj+cN+sfkjN+tpnCbzfuc5dL8SjkemfsxUFfGgtR9M
HGU1I2PO0nlk5+cOkO5fkOyrIJlzPCBvitlps7AlqFlc2AR2FpbUHDVGATgRluYP
oQxR+R68Bew2HwyFFIun7SiILd5UJD4nB8xbbxCXBr3AD+NP70G7bxYpXJty91xw
hGTwdWwrtH2WQUVP8ZY5+44SwRH8U8p79FH/W9jO1Weu/FxjPtLIyYS7dpO/TPpV
EBBmGeVvC71hO0MDObzqBEqUPho0q3ONLZPnBgl9Bq7tecxHYyihovnXdCFFTQ/W
z7H09RE6everdbUm5RA5iP8FCzNF49VoDMEBVvFrwkht0X6bakwOgUnR7tdAZZV4
Rx+bws35wt4PdRsiKt7DhBD+4CXkJyjq9/TZ5eATUlionksITgH/bbxla+yAq7ot
x749d6ZfXY6/BTzodxM56AgOwH6a6QZbRTiqHadytGLIyzBf0UHYLH3ixyEDOgj2
h2IwBqLclRgwuLTYtOiAO0o9MyIwbUf7u4/DpaWZGHmJuxQu+usNQy2Jlxf+KV+a
NbeDpQJl2B7deJXPx8am90pbZb53F52tWu2f+6h3T0HxTbcLLnvdRz9Y17maj0Az
ppLWdfdW3t6BQ28YFHcNx0zxHFUA06xFE4RVQJkeeG+YmYuoE8TILT7JFoUxARXp
Ybk1uhnA9cfnbwhvfIQRa1Rt3Q+0BDYQQW0BQni2kvxXuuUvw3nclTvrxciOx013
wSBshbUYK+5TZ3jay9SAZM6TSJYQxfUE5xsZ40vAN23gguidaxgR1hre1FVCHR9R
fEDzFYtup9gZGZn+ikyriXdiA/+5BbvrjJr6VBTAtitKeNag44k4pjsfbcuSzmt+
vpEYx2FBWM/Jy79XEKg4SOUMpKLCEcE1SEYdehsp2qLkUTchJhI0JXpdobvwJ6Lt
7pcsjc3+YmsZZ8OYGkGgJtGX8ETWGWCOjkXZXr09d/oES8yk71W00FI+6PltpE1R
yURGRCJzoNVlILbBq0jgUhuEGiFvSHmzIfIQMnOBS32CtFfqCtgT9uQF8S2K8m1r
iqO10OyA3YG8eF4M03WN0vT2AwGoHLwfLoQ1v5nA2mU4uFlM8oEalt7Cqf431QCZ
NXT+EcI141DrloeaNCc5MFdhYxo3X2G+TvWZoHPU4BFW8SjtkIRE01VaR1XGt2qo
bTpr1Gqt3s5vJsGa0LselFKK7+X/0Q05J55MGfEdPZdtbdR0YoR7QDK3IXZQEe4F
UroPlvDvBwSMAIbL+yBT/L37eBK4Rqe87Dib/gPAINIsqyI4CmNbgbQ99CQ7cvbb
TdO4NHU3DXG6/a0txbEWNEZKDzAlLq2/9lfjjMpXkFnnYDdlqzJ8DcYjp0O3OIZh
6DWAtxHmKO7zrr791kC9SfnkASFl/slDjhAkftbVBsrTqyFwOPYNIeUY3dtIGnHk
5PZPqSGvzMZb/OSm3XI7zxpREjr3Fosy8KQKyYGKKMSueSxe4fNLqGTg2cxxMzEF
gThzFrWROWM0ewrkjxkYyiFanyz64IbUWdOS5VMnmVKMHd7PscOM7RQzM+FB5pKl
vl2EA/t5VuEHCjWunl2K0i2f3587izpsn0DZLGe9ktxaZ6gbiUbEZX6Cl10lVNOr
6cLLDWumMw4yLwVYdLskbT6hm12nVJoviISujTee+j1eH4IRnRnjPv3ZNbVeLz8g
a58bAHLO5ruZdEytQkIeT3rsbaWagTuPWBX0vjh8MFECbwu86X1AcBiFZWTRwKda
SYK3rBobJoVnY83ppCGrD8T/kc1MHJItKD8v+hHI+FS8Jmf1VLrMkdJ7VBs4oZE9
RxoWcf0b6GlEmT4PH3j7KTiNtkJO0luqGMEG/T2hLvW4HP6Ov/SKQ614Gv+ax3NO
8OtTY8dttTSbnV2B8JOlJNbLrPoKnOul0eRumi0xN+DF/VuXvWxDoX3LJhQ/Ke9o
Y18qcXLpd7/OAN705Ss6XVtC9jEs+bhDjzgjDs7vssTIVyZp+3GhQvOrf9idaQKd
CZ6RE1TSy+ntTBNajsvFtcEyeC18wsGmbNOfEwTJyIPzq+kDiZKVC+oY/tTBMREC
rsltYEUGUekNjjTId3kmsa03JgqHjJSGBgTk3ThAk+Ubn98woV8sYBAVIvZfYtIv
SxA05CJbQVbhagt9xxmjnIjft0HdUbChLUiPFA1P1CW3i66xBZEcpi9WdH34d4tz
I6ktKmXlEvWZPrJPJs4XtZ93k7LPXag1Q/f3dUeLVKzEZ9tfkr2/UzN6wjq4s0a9
x1PuYKQKXF0raubMovVPJEHIHnWC+cy+CYEPikmnx6JJhQQgO6pvrlMkx7YwEwaJ
7WVFDGsKJJiA+blB/CSp21jVMhILiIyhbeUIJ//g3IIqwN+rtAwRgzaeBSviZFkN
76U281UUzKpJLIO6vvEVfG1fPpn3IIbIxl6Aw+SL2IzeB2oavOj5FJvhqL6zVyVx
sevNKAu820xffVTYdH7Q8ZRutAhAbKlZvYakdtcIEWnTwFFvY4cRNXqiQKSnouvx
L4faM4iIg9VYl6r2inng9ckMQlGfYrdW0KNUKVdr3lJubigfxDiLAteoXdAktDpV
laZzmFZaThk4N3cGcPDMFVT06o77k5q/gbcF9du5oQtOaqiQhT6wroQDx1lUKcyr
hAdzNIy1f7qh5FQQPHKBRgHyvNbj9pWP2hlo9/H8sr3M94KvRh+PygCBytliRhRg
JQ25vIrCP/chjjrR2P/RaN9F2lScfCHmbgjrkUW3Pn0P/mYJNrcNKailSP5KhB1b
6KRLOkVqBu3RiYKnH0BLBxrVqtJCgsXqlSfphjHurw8XyH08smD+mVu4veUXp5Ap
fwFMJ3UB76Jrd81lBeoo36MvVYXHFwRv5irjMAJTsM685o2YZ6UEUNwZiASr7/01
5BCa75H4R/CxlXobeAB3N/5dvjGKMt/UfEGNzp+EAncGRK8vuYH+8b1zAf95JKu8
KyS52QRYxTl8iav6ZvxtgBXv6w4cHr7/Ha+D6N89NcxtwO8o7rSb8laQqw8hDkQ+
WpvrzdMeQxQOToW9Z9F/jl54f5M2vb0XiSRWwo3WmBfX2JcvGCN32Ts5+2VLv2gF
D95FfK1nANaQfRWT3Gp2vG3ulB7BJJyPkFhRbkOI3kSXpK04XpMaaqw+wjpFeU3L
LL6YMq5loxmA7UkkzGA/9BUbWxETlTO0opdyU7F2JBGHJB8yY6v+H9AuGpG+LQam
XyNV+CbIvKJkFdA7VzCTBGfnMBGYhDaeAXpJ4YZxq8+TBASggDmnvVZikjZ1tgiK
mcZdLA+cX8SSbqp2nFwCbNrPhoWeszWOJVih+yq91rl6osPRtkry/PF50Xyth5A/
rsYVyKSiiS0OD1wjLNXCGWc2kg6WHTrAkzDrGLkbdH33qbdcd8tItIYZeDoh7LyO
mZNZ1qvSisp6/CFOHnBL9nglsGJKeL5Ms+DYMlU8Vrf7pbHoK0OBBH4VvlA8wO5c
HQfVFEoNmjHTKXXwHUpdsFLXkCNdCWXW+jmfcPvlzSSqjupWqKrhENQrj+gok7Aw
EFh/YbGCJ9B8RPHUaWiZT6UWMEZa+E6hzbfQv9yQY566D4JsLF6x929yJmvOiYG9
31nTzxSIS5eVgZ4AVyvx5q0LBFqj+Yjj+SmAAE0BaB7J6/EIEzDIsFNr2b7a+bDc
hduTp1kkF8ZhBPibgSxX4PQuXyV8pPxX8MfbyoO+PTyZs+AKQ/aIz4oQkN2D3YhS
Wk5BfAcXzQDOEEP6H12L2XoTt0Igapk6uOfi5m1yL+pRSGnYSJmfzpczIBiL6ApQ
+cHGBLoAoRrN5kXfo2RPT6ZUTZiraea2tEPgTuPJ767I16ZjsJeO1+amihdbJAoZ
vvxWf7PU5WUxMpOvC6bKhkmZCVmG/7jzsCAqIyyoRevo3KNu7qISyYmwlwknO3X7
UK2lNCawIRAqEcQoEbRS5TmGOtVZpZ9D5Edrv41NvpYsJD+aTDxC9hvI99sXS1GI
XDqBV9BHqjZRrbSRysWcqqOrlUdxjT8CmigCinINvVJKzS7XatbTIAlVbTI556Mo
IZlP3IoGrE4ubrZlLN8QTgvNAxwuAGRCQrO1F7SEbCKQTpsu0feIN0RHyhxTICDw
mnO/uuZ4d2Tndd4yepGLs1xDQ5WDsPi/7ICULQ5Pjst5ip3+7+DHAXINQbsRdVPh
azo7SvhxVGRCSUqwwJ+/TsJ/Z7KM1cZCZt5j9L/fQnYyM/6p/B5QLx8EOoKfkVFo
bYmfhqUckxMWK1mkQvn2wf4IY53o4zksVsIugNC8Jdp+DdzcjHkXJKP/4Z7Ewaak
T/+kutHkM/7Oeqs9s/SQ7MP2LE0UDx3ZJPwHKbrtM2drTjDzvC0Y5qehPBG1FvGQ
eiSeF0JojscIHtIeqHjBI/iweNL14IJKQn9pZEYbDJAm+LH8lKp2BvvugJsHUZy0
3YUMHpyUPZ5GUB3gAYhVMK7oVuNN2tbUEOUH8giyXLwoDBQ5y9H4guLF09ctg1Z+
zy6KZer443zF4ZOyXm8EPMxgZnGnSYrsOl4fOPCgIIk8ZXVCSvVDC1iAdZK3a5dz
KaihYWwa1ZJuZTSuW1l1xGI2KUhcBEQIli+biRsdcSXPp5bOnU2AyL+6b+purd9b
+xkBF0FiIejqvH4d6kQTxgrkS1ewZf4JiBI/P27qHiPNVn3/Xf8NAm5nokGraHeX
ASN1PnyOGdZp/v2J7vO+RHuBD7iXeR7TieweLWGcg2kM2nFzUti3ASFOTyp52Dx5
sTJqvkU4ormvUt546IbrQnvldEcAHmBO+wFJDxurnN9r+uXFWZm6m1SzScC/HZWX
4gMTuelJxjrEzShEbATthtgr5SBn8z9s0KLvxVQJAeI2vU7mth2IqCMkEn2V/U1x
mUDfA468Ikkfn0SFB84eFAWX9MTj9Z3oM7mwVrUcfaycZuundNaJU/Ylqpi7YYPf
Cs2EI0u6bv0j8j3KXAAfOMXhQbDvuPiS8FJsPJ0f1KJnsoe3P0jQ+hZd3ZDDfv40
1Uz+KbWHVydKEtaiXLVI+cZQvjHnS/F8P+OLGalKAKZRu/UuUJ9+9VMgU07cnve7
ayWENkKtQ06gRsju+YsbZ3Kwx9dmbDEvbX1voSj8FRjWAtgONdYHq4SlhE1s+Wlz
Lw2BxCw7qve8dzriQpDJ+0sP6AaNIXcPiMm57CwahQr4gajzET31q/aIo9Ny9BWS
BZe47GGfeXH2bdowKR0HfzaD9jd0sWz5SKvqET+KfPmonfLEzDKkCqCY5HU9ju8j
0f2nX65nHIVkhdVzwH5B8qwph2gU/FTWH9cW0E6/sy2LdMAAaaajf3j/kFrAUy0h
2MjRx5FbjhwytTbtInsIKPTvNa/QPueS9Cglau+gxBfL5tVaMZnQuFuKOGpG7iBG
asD7mhdLABqpYC66O6OqqvOEnRlZpacXDrJ57feJA1OQlKfcHFRIQgVmd3azGDyY
QkmRdG7zMtQMSP5Wkyt9L6gZZDSb7AKDq9pYE6QXDuLOLGLrdN9KZmQhZvjfmEI4
Xfr+g3kW5dHz8piQ10C7cgRUMnPQtRNN8SDzfvckYPCS5FS9B4bQhRgJKYd8NUeH
+981X0Phu41fsE27OhPSYFYB12ELDqZDmSDaWsaGpZbEsCygYFuYpEPNhRJIjTPb
i2gOeyC9wV/lA7obVb5X0cJdDeSc8fqC6KAzZ9RExdz78DTMaButv7TZKGWra4LG
V1zx/dk0mpHGU8c4lDX/qkFWh56STyqYogmKyahIAyXMN0SKTiZ1PPkc2cXEPaZc
Z4ar3UraHEdXyqilqES3Boiey4T4RemjbIxVBSVvHN3oYG3F2SACqxYKUWV/EQFh
VciK57zXqVWR1xyLbJM27wNMMPmRwScJWs+H0J8E4dbmx1pzndUByFWsroQK4Biw
+9K37TgZl6kxJF3OSUvjaiKYHcvjMI12H3BqETzM3WLSKOHsfqjla84OMcSBL09l
lAGCTcyxkQMLiniwmJuWfyki1OlDPm36Zj6OeoUszrJeoLpVCA58KVkGK+Qk0kUF
jt4T+TCWbZtJPdXO63d53Y5Mcq7nLuhkI1UD5/+NPjaZQgMSu1bbF9/7Ro5tmJPc
8KAaoODYyiY6Ct2DB+/bRWZBUGosy5CFBmEwhL5tnke2/s0i982c7Ph/+EbObZfh
2EncJABByasM8FDdhuSPxqSJMRtTwqUx3bznawmF0mVbLEHBE3iQxi5qvvc5E5PI
/X3SrAAwzOZjuqLSJ6mTdJDLDqIUcptRl6mm9GRVbODxpEi6jSJCgOoBaJzqLoe1
5k3Ld/4ZvSMBmvE+IVIJ8vViYIbxZETt4VCu/+G31/72VGEynK53JQVwT1IJ7Rzn
aHFwrBMlcotzhS2WIgMlk7xlWk1+dTt1xES+vhgC5aNFsja/GjCu262qEVqNNfTJ
i8UbczrHoleo0NyIjmjeqDZh3jfbvHQXzKqFFO0I/eNRADr0tSHhbKtGC3uwwTXJ
qXwRhFN+AL7HX/qPoF8sRyqNqAm6lQ4k0mmT3n2hQeygvLo1ZpXx/Sd3blSj4WVt
lQ1JUycvsnX+qSjvnr38jqTepgOIvWzWbSLrskNXGFVmUkom6cBF3k3GrXQ61h+8
/FDT6JAtD7LV7723ATcjXB6DjVZR5XR59BVzt5pVlBCZYnr2e148ePWzkPziEse0
e1o+/X6UMc7yQm2Fy4KZopziyNwb0U6slHbj+/udvNHwSmSQsbz6c6KaW8Ur7nvZ
n1OrMYj+0JTIq6RFPrFWNwR0awUYWPcF2hkFS9Ewjy3D/wo5JZBzMV1qa3caIXQR
dMGBsvylcsb6jETZg6C2GxPLBWKiO8btnxk7S7RL1r1fbIqEXPMyZ2sJYHebCS7l
1FLLHWMNCnMRpghKT7IWnvRFSGYNPDNgK3jRl8nz5yXzM7JrxS+2Fn5RuAjrBpRc
VmGreuxKxLYW8ZcC1rauWYMGuSe4lAiJIA54qPkGB/rmR4Q37pcFnb/O+RTv+5f/
Jli0Fg3fqFIUw5hloWHhScSVc7ERYpwuQFAoEvLO87n2tr1wnSNBfAPLL7uisqks
1OfZ+lXf+chVILoe8X5Lae/H+Li/hOEkyTckIWp17uDGQ2b6Zps0DZ+x7XRHk0OU
MQBjCvd1Ex2xTDFzNOMfB0V4W8yxTy0IXcIm1/IMFq7Y4as8MJDq7acebRnUYILQ
qmedu6e+G779Gnq5MRmhIwbKom6/Xy1sFYURVEwVdW2kj4JtiAYq5BOqZJwqrmiF
ck38d4R+jpeCZXtliQjQB+PAlE1KlQa8g/s+lmSbP+pY3Rj8pALeSkX76/bN0IQj
Ioe/H2kN1hl2Sx7Y8XvFH6ji0eRvP06xRgjLh96xUZw4YhJqrWxBcGVHJNPM3X2l
OCfNNhoMd3zMxKN7sQ+0lySJ0xTu+5aV8BaRJTB36VtQYe5pSttj6bEBoPHkBnrc
Oqci8OemcatjYEZPS3dLsc6k7IOLyGfFHSfjPvECDTGEhWWXwdTVMm+yNET2mNAD
o+ZgfN8ViEHPanOddlORDDqry50aE3M3T+PjNM6K0ogFdXSUzve2nEi2FEcwEj5a
5W4zPclCMrB5WbjHq1e36o/DHt1lOQG1MdJKlk2+tJ++SHfjtI/NXFS4fkIkzBQA
uqz79faiiiTwuEe6dnA9mDe0AjJtS7V2aicsl3WFE2ndSWaMEswVzhOOPZWWkFf+
nNqw3gYtpImeDggQ/d2fHOfeHTWJplLDoIr7dcNHNokKQnQzgQN1UStSjWyWY31W
tGuC6/NxLfWaZEXxLqbAko71JJUzFZOJpvqDZ8QX4KLmdmT1B2RgeV7guTUK/Yxh
zapsRY1Ub+cGVJK5HqBXhrowlQ6RaP5QrwmhBiVfWZ0npXndIk7DU3PzRC5V8AIK
vCDu7N1W6sZZngdTvh/2txtR6xGRVLeKw6In6Kx4SPHdKOLVCRIQkIvMlXgfXhPh
sDltBLaNc3OeHAwB62gKW6PBqwjhO9aU+hqICXniOZY5ipHHauzwNfSNcoeA8ouU
MR3hWHbe1+m3mhQAJqu/wEC/O6Tb+cgLweH4f0NMJU7ww6//OXr0pI6TObVmhXhx
o51ycyMscI26T3qOBWGoqtLKSekU1VHtOjABXTOPnuOPakUmhbOBVS5EgH4wiaZ+
051ex8ivD7SP/NdSL/ZSPGAHhRddDrKk5Ypqf5ksIemegsLIA31YzFIA5W6uVOJq
nILJGQ07HieeQ49nxxYts+6MzM9W7ZYKjXB7I0Gtk3nnIMjv5TAjr6g/5/uu0DL/
XVHDrHplhUKcW8pPt+XtZEDycAPOHd5BeNO+uxIjb5UYWyhK6+rdpF1H2atwLGRG
cHWOr9aWhLqxjQTH/4ZrclAcSm37VNr4Aam+juORgkoFr1VJP59iHjp4IGRJe7Ao
EDD4FFPx87eelPVuvl7BK10awWC3cswe0tx3eeiH+CaFpBSbDf4mqLbNrN9m03a9
XqgoY5XawDQmXjNr1mfhOYMfwbns3Re28JR+8KWQae4JpFiQG3U44brSC7lnXtpU
99KNEWeQ+j8Yho0BlelQSdbD2HhnPv/N0ZI6mmVx4gQncNDvrsHbjTO4vNcA1Z91
JwfZ462tJyzprClzWURD6zbseOsQ2dZjMCAqTU/y/GXVOkYnD4ojkTQ1kYPFxM76
NKwERmTw/3K2TflX3OQd0CXU27guBhH4ohupgGsunvmmneIU4HYtil6pCmwZeChh
TUCUc5dN8GuCFBJnCAr95lWloJfAkc7OjzYtmW2homqC2jXgp5kUJiPpuPC9zpbb
zVO+AeXuJjKHLEJVtX4fmwA65cFjkgGtL2RqKAfsoyiptXR2ra/XdN7IAWMSJcFo
RfzwFAovaoMiPtJ/yIv6vhJJPbpQ70NZSPs+u7468MzqzFtYCrU3rsAzmuOzoIyq
9wHVy7Jcr7m4mPw5FYWJdc9HIOY4qcylOHPc4OgbR46YaxSWpN+ile2Nh6O4y1Mn
IF6r9nCwCoYFk4T6CGa1EHIyAsBdCBzddDJtaIk5eblSlu5WaTXmYjMKjzk4MVai
KlG7kwS2TVzB+Z0ZfdGSOg6NevM+aPvXg6YYDlJamnwmWcEAsZma1cE9Omjtk6ko
mPnodsD1yM5qKrnGUqvrF2o6Zseb8+N2KXnC9l0y2UpVQGXv9qUB5vFe7am0Dhbc
1rmv/QX4wFX8ToIt4Thk4n2B+kJgKDrEXpp0PdSgqpBkaXboZ/lQAL1jdNFOotnp
D55RH7K3ymjiTpzp9pwSUSvsVfU8WXuClzg0k7Ex/+L3NtpBtSuGgT+OAk8BU+6T
kmRTBOeESV3uqJJ8pTlLBuZ825Tw5e2Pi+coKEFQzGX2OxwtFK2ScFkQ7Vdzhxw4
Mi5kqbVzuBOOYmv1ggM5Gqzsn8hk2b8QT62WMBLN8j3gVpQlqDCRsL5iM8S8mQfi
sZWNDbTB/Pp2uMC+1F5EsXAHueLQEVIq3tMK9yeuGkw=
`pragma protect end_protected
