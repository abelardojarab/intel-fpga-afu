`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
a5fLRlu3xAt4h9DUqVK34XvlzW3rTpxoPuErggZQVABWYwngjqIUyHPCw3XsNUKp
33KqXDOBmCHQl7KzwIPiWdV4sXosdPtWcaTo2k9Lthr83hy0FhCW9OSNrv1pHDTD
eFTw/GS/6FqUt3krnXP6IYJvZ6hysVS1+IVTwSMm2nw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10528)
yHkEmxeSlozjGWnpUgx6n4QbZJjehMSTGE3cOxNLk/fA4QSj6/QZt8nz2YQk44qD
lSrJ9m5HhDLqA4dg4YabAV/Pc3AKLxiZKCQYXT9H8cSS1wcQx4SJhodV4opDT+8L
kpkBS8azGpLYt87UpEqqnzhYN9WJAqb8t2+lIrw1FJVXwGSb+Qw3Fvrm9w87AEc/
5Hj8qhziQo7Mu3Oao7FdiXRnZ7/NznbRuD7u//rFO5Z5aAKAm5y6q+TT6LoS8T75
FX42ZEUh/Jn9LazSX9Q0DS3tlD/m4vbA8qSSKywTbxgP88OHmZo1RLQDLVNFvf0X
ugAxgZJzJ6EeZbt71AeAykLon8NwTwTNBCfePcz5r10tLGP5bHURr7Pu8z+Rz7vv
itQ43vxZgZoFOZU5gHrGMHhTq0vmEzuMwt4Tr7hOCrwXa1F9J+QnbSZhHZe3ng7M
svuZnku+TMQirFtBgLPitLRKw3zxeu1OsCI+xDFKA3KBkNfCnOLqhy0MkIhPwkw+
/W2DX8q3DNkheFrRCQZStVFWi1UoYcYDNOvWqLqoltyx+iVwYa/sPFo5dUNVlLbI
1/uJ/BaiwRMwMrWhk0cp/n/XN9mpk8i10m70G/E2nsYukWbE4A5ytoN7J53M2RF9
PF+t97kqSi9Dh6rf01l2Io3PpYyylOohv4YeDTkoLfk8tV7kYcYoZPGW+cTnZvc8
EtsOoGt8tnQ906iabNG9GtAfNe59JqzJp1Qj23gWMklYMSQkyCfCE9iDeetcNKQB
6QBKBSvKhA1ATQVXqcxwefUN1o8pLrKquFyd+1PsaVZtr5Gb23HmMuY7BsB1UNyK
3nkzuOxL0zstqsiZg8Rc8uw5sFS0IJoKU7YjWFcoEni8edeHN3jaFjxVxe3ZYqTs
vVge2VYhWmPCLYr4uk5JjaJnt69RZoYbK67q6oyPaOFsX0rai+4SpU1LOfftbWFy
NLRmu+a42YrmF/hcdJu7B40wqCuHYqoga1/gC9PK5oHzumDn4KMCbAeBvZDjol8J
PWdEF1F8OvITEjErIq7bKvWMmFsKHCMvV+JjRrGHJOYXluMGSQ13SCEAi+B2Y/T3
p6mYGrXO8OLSWg60xz+mhGVwRZa8O2koeVs6GI/czIpqxo+5gcsB5wzPp4Rw84XJ
RvXk7gcPHaKcgBQ7ajFtexHHXcnhZ2nthXLGaq2SjhM59RGSXGLPkkxBjsqyqG/q
s6aPcSorcx2JMZfY+GQ3Cn76W1FgLlnqyFSEuLC/faqhUCC+PtXwPxCjjpU1Bih4
kXJKgXU5u5pmn7s4Dali3rs+vePw5ko2gnJNEW9YBTVHKJpZaV2Be2hqjYuqHeY/
Cll+XxqJUqSqtl6aDvWJ8ilXSu60x/A+ei7mUlrgeUmR+6BJ7tUMklMEVu127u52
Q+60ewXrynb9F9hrf/lgYEBfsuDfvRAJSyr71J9dSI9mkhHh+sCyjDqZpQ6mqgDv
a89t/oqJtNGHnYwJUbMyv4pFYMjr63ry3zIGsJ9of+qnyi0FznKDQJbPZWJlTpN0
m2mArREeE0O1XZrmxbuAZI6mv5hptl6RKQP6jtuA3waEPKzCaJq1iQyXGi9s2WqX
P1bhVGhyquvnSr3N9JDmdVLZvKP7CJiJmte2AiubxUK0qDFUhcxOm1PFapJgXL2C
FoNr6GtKHQv7j2mftuIqG56WZ02w4xE2A9ROsrVIw92K2ophuaCTYsLo76Eq5irG
WrwdSbghWx1FBRGaUHMDT7uduT/c1NQ+VfwzowD9biu63j8maMo/P0dBN0eJ9VyJ
eC/sBb7s3V/ye4QzWUvFXMwIdVbue9TdN6zi4TRPPsYwF8AIWs1etICMdJzXqLse
rfy8XdtnnpXSpolcutTQsJyfiszQ+BbLLUOTvLTIeuQLrFFfRy2TruZUiE/RvQgz
ZGp6xFXNtnCgDgJh9gJEE7qqpsfWXaFmlfohlycIt6I0iAynk8XXS7NIAy5Ya8F2
QUuS68SreHVuiUo80TTAzaf46c3U5NvvbXtroDycMcoD/4RuToqqK7SdBLLOV6RM
e7ntzhz62ygh08od6XQWZWnJV9TissPmU4XNT87Tb1qMp2rzVQ7y3vFKXY2mi7XS
PrQ/wW+p8UDt7o/mGCIkXn2aRONljihlRArU+uv3f+V6Qi3VWtyndFSgP5W/lQgl
Pj0tKRKSx/Zr1F3awUNirQ240UL3sEKeHAX3nenKV8TMLFqXh1Uk5cWMgwzVAEhX
b+aVLRv0ShT3PXj7PkSYotqVqcz/Ca5uYQCXDyILbDwBbyf4vozbC11rbQndip48
Ek6KvzbAIW4dMtOwy9vS71LEtWW+O4hZ0hhMKn0KEss2qkUDalkEk9FmsIE+yI8C
VLJuPfT/KoZqS/ZzjZJ5berkDhFFcwn7f8t1+6PutzTsYf9PkpINfIXdaD4NPgji
dJl4hejWD71dXIPGq55DOsKIoYap3A2u8lfxrkLuMeRACzJ0F5812RI3gmTV3ZMq
HQAIjShkeKQxWn9RKYzjuK3Hl4g4GMG0p5bDSDxAZJfHVJSzdnYELqSTR3iN5XrP
f/BmiyNmFSNtM0K1zwpKcdqF0XqK/JLCvyoR4va2ppO1RydPsiNdertrtG2JfcWb
WqyiIAJKHIW56Yum696vyXsBNmG1KYgFLZStujpnOzVui4QBV3BwEF4wdcP1bi4I
jfHI29gFZS+ZlYLjxHWcoGLrkyFHBkO4pTexWsfFC+kZpay4+DaY85gGclUlMU0Y
aSLBZNsEJftljGHMpUA2IytxsWbekQQTNdpFC2VhvhlmYr+pdfX9X8sZxW9Gin5y
cIRFUVcHQof9JYLpNcBkGlPczp0jtTCW5I8KF22YkI/3KKGb4u2HR4oZrtQcNA0y
TJhd+vocSOdb2lVEMxVj9816ONrUiZhRGHbdpECQdGY61SbU3OwL1rjwowQmmqdU
fruMXeqf56+bdLVgpmWiv6Yj8Ar5oIwHqB40UCMxiTBDKEox4sfnE10PrDLxIBIW
BpRINrV+0XuWGooYLcdyh+pejEE81/st3zvH2sb+06Zgi/UPh5Ox8f5AHyI7Z8og
shKyYXVEqYoKe4mBZd2go+wipDfhetP/euWWaWlR/xs8/rn6fcw2aKc94x72XWlU
uuvd39Z0Dmc0IOwBlt03ves41KZRaYr8rHqHbWVI+pZC+zlqGPqqrCopX7V4RSW8
lYI/I2C6BDkmrAWXmO7Z/U0G0ypM8gjbY3kV/LLR3MWvQxT/X33KPbOyeJsFM3Y8
Lh3+Xek1pS0tg6LcYR2ApoTfhfuRDbH1g7MU03USKp18HY6LU8kgWuUFiXModOQM
A2GCyekaCeCZUAASFi8RYyysrSmYoAr8/tbX1WWFEzRTGPyHTuaT/O2/T+o8dxyO
LEzewrnAYY7/gb8vGeDCE8WUkSOYrbYQTjwNeWcW8TN90J5jkS+5rP7I03fqzYum
bzM2mLHmov8/qL8Ixf0yGhgZDl+r0cv39Cvl0Dla+p/p9jj6rbtzzcgswdohag4r
bfUFpIV+32TWKdpHrjpkkqqsQDyNBtH5iPaB8bofUw5i7/X+y0xk9AdVBlSo2ilI
OvK1D6CViYn7iHwwz8l3v9swJaP87N58rqUz1cNvCuqGFY361TDSLzHLSBpVV0a1
c+nrnz9ln6nOBB8/h4ymh8VhalQagkzXIQSHg4VVhMz7Fd1d6D+HoWNVPIudWWMu
EyNWc/wUzT6B6UYz58RNhmJ5BKMBlhPXb2LGEt1efr0EHTRVF+lJ2nowaqNHTqSK
M7lZoeLujhgg8E1aF4fo3AohhnRQ9tdpyz66zHRYGgOu2mNkCRNc9MIIONPxXsd2
veTVSH83oZ7xoM+KMYWASoKe93wMdtj9Z8g1KxEYJEZ7rz6iqg46wcXdgzungSaP
W87BoA4E+CmoQ+U5o9TVqtM5fX3lOaC2qaNS+9yCHwn1l1G3QmWler6ein2HPW4O
REaNMAM/9Low0DbmDsrKWFBOGT+w/qAr+flkyVXwggrRlMjZYwEAouS+LYOjA7sB
yJklFeeJMhcKl2Qy44KwzzoXYh3BbzFsLSbpwGcZ/1zNr5+5ePECNl3itLQ4qjxg
W7jGaqzeTSau7HJX0H7M4I16IReClBEoAHGFjKOkxdFoMrayGNI+ElMdz+HJm2kw
yXGgEka/QwMiAYhigOXzh5Yjl/WUN9d7qliKkd9H00CHLBo6yP6AIWPj/7lYIS2d
/Xy6Zorf8Ie4o5h3lQoxSvsuCt/txC9tAx2hjLqkgEaCc5WQojYm/SSaAK1m0o+y
6BoXJ0FyR1eH2ie4KYiZ+mmJWvcjto9tBFGoAifKiRiy/8f1/4atQmqfppz+lEBC
BZHtGbVsHqvL36+8jhD7/AazuwwlgZXxddeGbtphUX1i6ngCll1ASkR5vNwxm8Dk
fR8DNwCd/+YMrV7sDwAL1LsEjN9oCH7jwK/YU3m3fXV9O0OY5u1oNPEsijFJiXEH
zkIN4/DuT1CILKYwnnrawy/1Saa6xwLN5d60wrSry+vH2I+hC1JjZqWAjjwMHho4
Q9CBVNmNUoMSAH5O9sOj5FUZEJoQ2Isgoz+urDVAICkZEJj81iXvzst+VgJlFY79
ZP+o5bQ4f+3WayeNMm2xSvj2EdXBpxMdBAVJASEGIGNbEb63Qqxr0kas3MqdZLOj
vyOzYBuKH9EisXI1YMZjPFvdg6G2WGiHOSg+Yij8SyvPx10yVcPxJui3EdfGQV1c
LFgNgneD6k9oRI/by7ZxfzndWAUut8CEmZnk36KgT7tlbwaeAmcjJ+5Fu79tgGqP
7wEv1fJYs6gH1rWBDrmJCgVKVR1LWgtnWoKVHtjfAgKOPnid/0ycH/Q5C7VkorJf
Is8ccZk9yykzWSTVUYo88R0OhZ4k9UwgIzv4IcAgE/di8aYAxXCEwyR3SH00wqMY
kkeJvqWXKebB36D3x08wFWioN3PX/4JR9v03mVXMnkLfu0B8IkCEvNQBJgEy2H4l
mwJdTcXIDboa/7XG2vc+ZOSxDh9LvcWR3rt7WGA+hQ79Xm+I7nNi1S/ugahqypgR
8KWM2vvGrx11xurQJ86yjBR/HuIWGKTy8gFmt1W9zuusQ4/hmg3gbQDIM2F3fe/h
1Z81D6KNdeFFJW3oNnKks1CTwPT4qIeC8m6wXyWT03Pb/KbmSndRpJ7Q8dd44j1b
7biufz6DmVR0SPzOxwnXKVVGeFGuI+FBwA2lLGNOGXWPAPKGZeubkgBhNc4P1HPu
+qCxGr4Q81zXt8clqsYKt9puaxnXr5amhLi65y1puWYUtpYDcrMt9+n6ycGuqfvM
HvSKN/pj+XJujyYOFlWH7YlfsM6HJbmaEroQuwur4ZANlWuJIR62TUSWMyER3jN+
cR4lia+t2mKdoZ3MBkpsgJkR4usu5CAbmMHTzNwjh4j+lAqyUUFeZVT/WsYSwyRZ
Ph2IbqOcHV3gVXNwqQj5YRWJpuasAXEaqXcsPtQQd6/B/5tgVsCtzuuFfLPaflUD
z1eNBBCeUIcuTchEBoz3igyp5SpPjhIheVJCkU7bQKGiNRmRnyCTjvvQ/Spn0sy5
LtAwRsf03Tb5I8dMbQOWGtbhPZzVzR0kC0gHR8rByQ778MoIpHPt9XbQzdAGhA3s
d/Qlfg3VI9DJkj/q5I9FEvlEJZjizFmz1q0ENdDDHtZcCgskn+gt6avxQAfqlTId
P3NwSopo3vU4mQyQH96C392mrfaf5tjdU1f5LTgW8sxpwe2ZMf9ks3w1Li+kfWQF
WVPmOfHX0H/GsIA6/dRlUL+RUibwlvl8ApaAsCwrrMJ4iZuB8pNbyKzdS3jO13v1
k5QaLigEoFtSsU8ONnckU5ICFR9MGuFaCIcUnv3DI9vphqamB+HyqgXVkEOH7Hqm
ar7AABwrKvjptQAalXjeSujLAv9lZrPN/zJ/OvbaXAFzdnq3xil+yw9TE731NUDw
PICUkegiO7RxNyJtjI8+zWeZdY6Ihkzc+xnvHq7WwkXgJZAMVsWZbg4Z5YkoVzaR
zsajXV4LBNeRfoH/bGNwpKI/sVCdF5GCLtlgOfWmeTdM24ZAtTxKL0TnOjTVKkwq
yvwYzsc36ARueIGYcTeOF1WEE1s9xSRrNl0apKmCoojtlGOwM+NuY4w486wnRA8j
5skSmjd4PYA1VkvtXUWrGkcDsjwzYRoH0WLCpMOyzVgJQXI64HIr/z4pXzBmbPHK
luuFvuAxg8bSYce0CQsq4arIqKG1n86vcVwz69g/xIlqCDawGQ4Ks6YhkBQZQ8hK
5Aj1xTDT/zbjdbvCd+RyrxV/cjfiVAdYuDjejUJDglXwTJJdnx6bUZrikgnTlXv+
OUnuQfpPN8FmeB+9l/8VzwOVQ27DrY89d1W/ZB2gQq7BPZweKva19ddxEMiaqvsR
+jjGBHAyT12xp8Z45cDYLpSfhuree9UVajlcnOy+0prYnykjoC9b9hFnOi5HwQ6j
KnRnw2VpsdW4ksnb1vQ6ixcA6sxY3+Hw5rZBVu5nJPAd3XsXc8W/zIzZLyZ698uy
D7WO67sTvZBBoN/aPsY3hLIVhA76T/3BBzsa3krCi+Ko1TTYx9JrQgyBbuzBN2mP
C5DPEkiYnu4nEbLQKGRNqJ2hbxbawR4ut83dZDlsmgziryRobH9UFg/BdimmEv/0
JkVO32RMbHEsfERPG1yUHzEn2bh6GmePVA4aamzQ/1mDsoTm7lJ7Zvf1va7JdQPy
RjT6dDwU/ZJv4HoGnjVXUSCH2aFFIXg9jnHUt63BxIUUHW3oadicgFo0+MpTbyA5
rjDiMu3vDEA8bVbF97LNC8eH/Jq5RyzwpPJrX2bD6JaPBY2oN40muDAbn/CRjcAO
KCp7Sm5b4aHWXnYiVschZQTGKRV+kJDdLpbwnJ7cFI1TCHmil5fYI0VLz+kY9SU5
36WKnIyrkHhuMpRL4vVd9doEnJeYVcF6NOBeTcxaLGMx3rhUwLpzPSa6OM8OnMPm
pcDbN054s+hL8FqfMOV0/aN8Ta6oYu48M8B2wahfG2zZJHQEvltNJhK3o8JIKZT3
LjBeKFBRJ606BD3YD1qWzT4T4Gpoj1NS7brAIEnM1A1RfSww20pkK/p5+bZ3ii4K
nzeqBkYLUzwJZvtyqGa9q6ZMSGSJ8Eu86UdPUaXRRP2Nvb2z4opR4ZykyivqBP/f
VGrX0xHjCC4SiZeAAjcsASyDX7E6YwiGRFWRoBULIMOuxvrQA2nljmzMFOar+r1H
gOujrpTBXLl/WNR21VbXwdH5GBZfL7qgEfAuWifpFjA9l/9Y+HrmmDv+gigr0SyF
NyNImyJtaNK+2h8Oi0lskyoQcoyKJ77wJzQPCfH6o8apAKRJfDwuJmUZqDREdDcd
sY2xTRq9EJdc6xYOQ3nJnSKvU6EuMTBNeFCHqYKq5iKuYbI1LQfTQJV0WVgnBmZz
6VO0k9z6eAVZ0cUEIXCtSsIQdDBluXuiOpsnm5+/lN1g0yoFHSvBaPdjr4kiloFM
ZcbcoxH8CZdpWZjRryX9e6tPKJoZc5WuGHKtzdjWUy3SHVFmm/47WhvXpbY4hzKw
UEFGMZ0i+PLqnVOS1JfosEeuKaAuyPoF+SB50FuHx11T/+Hw0ljLKQEBvUKCy+Xj
LRs5adK321aOK0EZH+o3ogwJZplOXNXFXmY65vv31K2FOmVejp5IINKY6njsNliO
o5SuIzH9kLxpCPVpuPt0gltDIouyBOlSB4mmdgXji4ruBEnkyEsMD8GCca7r8twh
HWnFmzWvfnKP7GU5bu/PgtLodIBsP4yKcRaMRRMM5lFFkZuoPOuXnOwiASSsveOP
ILiZW6uFuFFlChqYlolfdIyov9Ql5OCUh6LZSNGhXkjUS9WTv27CUr4wbq3W6bwP
FCRK0xoHWtFsaMgxXtj3fM7vJItYzNU2AjsVfBueshbelPS3ui/iXhVHmnye4f/7
tS53CrrzSgS8d+h31wk9JD+Wm8CvNIoOPFlyJM+UD8JUSx+wbFi1vp5oHu+fpwMA
et1AAXnw4Rfq/qePNcIOqlzUQOYHZ8HiuMPAFnpaAQGs5pFkw1gpEhjnxK27XpUe
mnaMaZUHZxS7ex0RuX+sXXX2EXABmwr7mWBq24z7yvGyGVM82alNHYeLApINiWoG
dsyeTVYVB087qpKHrirG5z76hWWN0LQsK38cz+KDOs+SaZyBns6Yvre5RBoYralU
CHrD2Nzv63a5RlOKZIEgBV5l4J/v0h7Z7OU9NO+qDLpvQDfjjwi/owA/ch/jUTTG
qEI7/WMHMOdy/J/MVk5h5dmBtAmPBT8la1ro89NdG0Jq6r8yDqS2T7D81R1vH5vY
x59O5AU6u4MWjYbNnPTGly8Jqyphx6soUyC/nWPzV0tCwHmni2fdI4rl0ckeibow
TRGTAy7gzSjyAK3FdXn7e7ENZNiPq0WqvulmrTZc8JLrZ3bmci+Ig2wCNxEE/0mt
TC09SyPbkvWcMHSlQqMlghWy3sZiXhgaEJee4XJi+JwJ20knbHqvXl8JCbj3hfqu
PNFbDqlpTYYE/x93ckwUrTAhahYXC2zgZAi9190nPICg7JwRloOfC10Csbbm5CaW
VNDuwfEq9ZkMUNHWTvTUQKGh0uJuxu3x737rDfI+eTRQeV/V+oUsanhdP2Xfs2+F
ZVBisuV7L6AdDVoKFMSyjb1Klg+45rZimomsAZIv9a9d7UGkeCAV4dXobkypojv6
rBn+SZMyIKa2kk4awlxYlSH0BBstuj05sSX99y+ZjEMACf9WHKGt5PdBa0fyGh1G
wAdxyDBD6aG8ilw7Oz8huFm+pZml0mbzlnNmIiK/1/V2j3cWpkmG+ToVZKIwz6PV
Fjp77rHEu2LqG+MngkvNGKyWsvuuQKKwepdTe0LRYDozaj7bmVbyTCwpCdNCDV/H
sAcK6gNbrASz2Mt64NMaDJ/TnyWc5NrEdkD4MXYGHvxUCnOYOemgYA1sss9nhqa2
hrYugxwS8CFEa5t3vVeV9VM6gjgRM1crN9OI9+XcbWG8NPYakvlfHcCM9fkO10tO
p6yGndtCN6rVlHie+Bb31XFwJSXKPWyXYEBDAfEwvBdyu4AhnlUE0G+zZIVDhElb
vyirOmn8uDOpgh5DFUG544vdDTlZT1IfCh2JXnPJaZngZK6r2G+s+i2X9jnspqzq
a3SISL0ZQXp+zDxyQNSYcpWeqq4v+W1lsZ0bmgDSgvn9Ej3132C76AFBUS4wK8uk
Rpdt5a++/sAqDOHZaBvoe/A4Ztf1HhoPDUidVZh15XSSmkVn3uk1QlUC537EgGys
Fhhw3wKIlXq/B2mQisvpObcES7wSK97nwFlsBbbywKaS+Qy3qggsZYXoShw2EJMH
fGuawmgiy9uQSvA8EOJ5upXaZBS78sO4/AI/avowErd2HjCEj0XN8xD8sUnfMwGf
EUWoQO/3qgA6WjaRFY5i7O7fUaHJF2I0KrMnj1JNv+49Gl+Ac+XGcE7cFf1t4ClL
6VqnLdCykqykuvJup1RlZWQtpCjSwHgZX5CnSdxKtVluXNkGq9xrvdcush1meLJg
LqPgF2iS7JDf22XKCFyaziG0Ra4gRGN9EeeSfDh7CYEyC6f9Y4jFJ2UNJjBQ7wAf
rkzUIAEd182jwM1kObFUrhPqgqx8cUg9P6Ktj4/0+9kmP7M4xJYsrN6aE08bIze2
oay8o84MlXaZ/IDdYHMqDGbulNAU+xVrrD+OE3QNOa3s93G6qQq3bAsKQe5AaXlZ
dvFUsK/GkNQCcVZiUhpvulqdG+cY/OO+lF4fdRsSiPpImUdmDNaYvtAfTblXZhY1
pRwJISXFpDHBd9RoUrpW762HfQ0euZcgkvqaU+ZpLcFaHUcBv6R/HDeVjgDFF2lX
PAzXFXv1XVXp6L+dboChogAreGx1YZjGl2nYwov01G2+SFN+8TIJnxZwNrIE3qui
9dTngElM+F/xNixACm7MW2lNqzSCo3/L3SmIlR7IgvyTeotLQ1WumzLwwJXzZ4iW
pgfPYLSo7C3l4bAzbUCcT5oqNOdGoaR9BP6+3+5h7We9BwsUeq2VgrTECYpeROoU
QBKrGCzBKceIn+l2F0QclfVjeG9sdOY/17ACuVncHu9nSJMKx/6ErivhGVBSmEqP
XofVQUDMGQtMbGGhTcTbtjMtCl64VRMaQGJq06ixcs7FGQIpM9U2qckEDmV14dqW
R+kfLXlG7G/UOfxz3o5E6i79cWbojkMVo0rc05tL6uySV1wuLHn19yAIJ4ROiTl5
83ZNpd29/IMedw3E4dJDfUKPbkwF5+QPCyuI0rmqqdtLq9asAX06sPCm1XfzoV4j
4dbc2rX0WgvSTmNnl1ybSJJm67yHOVLgsjf5Lq5VTzg5B+oORUAstq/ZO2ShyWBF
59/KNupW5xKue1h/9xSrD+HI6D1+iuZ1l90sRuMuRsD1BDgDH5XQTIxiPWoSLAGX
Eq88svFmpUa+1vqg5mctJ+DHTSraoo4z/BSyDWv9OSpL837aQnctZOT+wMdaaXjI
voPrcjYKe0QS7azw/LWl84i9v7aTUSdA2hzsXqc2llV+xS3WYj6J0NHXNXBI+ngt
mw8wdPol6E4Va1WuD/QeT9bBdAFKvW/a9gFxM3wpAhFim91T5VKF+qb2KGUb7cZq
9TFTRCBjymADUKuW1+qsuKhRRBnpjEpVDejg9eyUSdzhAOQOyVhce4n26f5REOkm
QKpulVBYeTXXCnfQ44N0Jz9x4jaA9Xt8lBdYrVuQ4Q/RZ6wpf4LwISMr8SGf5FY0
CiaXTRKsECPd5PKZ5OK5Wxm74voKgHenxIA+yKvrrcgOAp7i7Y4dg0Xztc1Y7yD6
ztliEtyp5NJqa1neulVap9J3hweZ/6GIPEW+2EIkY086RQqdu1+8GaRBbAHKaxnq
7T8zz8ulIQTjO4CfWdWTTyHYHwa6mA6LJHRPBKURhEJEJIufc+By9ijX6hRRBmGb
km80wukfB8KOiuOptGf7wRGG8PiEeniaFifxiNtJS4TlHFNa1yPE9tpvLfjGqMP4
6Pd2IhroJoMBeiR8TPFo8ypD30ilZGkof6pJW9vwb2ptHGMyDoG/V3sLPpDvC8qS
gyhh68YUAYIYD86TZ51JCOnr6fiPcctoDK8VmMG923UNJOVu0W4IUzFYGYz0oxy3
qpI0SfPXm8iImy8gazn/okzI/dxfkTi/SmLKAvRK5iEyszkYgeN/WlPD3aAYEQop
q+uLr/nQWmBYTWaGjSGT1J50CJ05VnPQs23qCm2sbRKmqIzAQFfw/6BSy/9nDUKN
lG1KyNoMACFRSycBaXCteqDtD6tCXvYYEZ8YTqjTN2tnWE6RxGtJT9cMfsUNHuXf
oDEVDJWLBDrA4Z7qcMjA3401IIJiQA++N+US2Vy0r9IIVnhe+QlJbzfrR499MW9s
WI8T6NyX1nuvhnuzXhVEHV+umcyDMGWuJgTTpjT9lVHDQ6iVLQbsZ6Q6qSvdvunH
U6wvEt0So344Tavdh6NuHrSi9CEck1UP8C9a2N+9aCPZhNOA0+t0j1mq7Fs/aGkI
Egw740cYx/kenoQlSkpVzT5DA5kp+tRAaBKjIk2efTyr7ZaUWakjZyHB++sXViNf
RAUMgQe3mn8jzeh3w8psgewJG5rPojfGWUgp5am9zJK3Adt3St2ALvY33MGcNd3m
IYvxTsrpFrWLpLYjLRHPoePm8zO9CZyO55EzG+ZMNffVrusNwZTsEzqVHR+Y1aAA
bG7Y4b9hOH3Ryr6lfUkLtJ4IgoXsxf0twLRibRHFjUPCma6hPVE/9VxLc9Hkc+iY
o9K2FaHQWRVeYKejtnTriggHkYyytmxaXkHU+wGTw/3AhBGX5BuuMqgEP6od1vSl
sgcO8O6oha9vlKXjb2Wro/FIpaa+IglDFvXE3/x2HQW5nsmX0sB+Rg84AU+Wd6O5
OsvOvImWVs4wFjcloR0LWkxKT/BRH2prjPXjlR18N4oLfLZVNHG7MYA0ybxPfpaB
Uv+6lKHXhVvHdAdIN9I8gkTiCEQOGeFSIyeOMNAojOLDJVSnNDCf2DgHEjzdZr1+
HBiv9Tdz7TXwfIaviZtRjac2W5i0v24ba2z+9LWE7JWxeU6D15IGWSAldXd4VOA8
jCZkF0b1ZZyeihjY4VBwP2YPbHhFLgHm4XImsn2W8ETVm9clfnmhaAySqoYlmyJ9
4oIBmVTEmjnjGmZca5migJMStz3Z8bJBBxU0mk4OPmXfOpMeOg/pdiIeFs1Idyua
5Bn7er78GJkq5tGWNFYuEVpbzli6lUTsFh4/6L2eAno0CbVvaMPzjpb5SyLR3g5U
Of7CmRXsfrBXKYLXaP5KOfywN6HK8OQvHkct3RbamBPW6S03S38u/QY6S20UqTtP
UWWJnO7ai+7gDu1+RncVvvuJb+pE6DqO4v9m4zYm6G5396o2YTHAkXW6pmeDsXGu
rJGcDhlbMUVJyiajm0d9K93dF16eT+mvbWMdr4pxehWk0oNRziID77VHwHVmYZ2W
EfUdvzX76uKbydyYT/Ll+RWmrtU3It94IC6/3fQbdsGo9xl9jwx1FSFST0SXMeTK
AX/pKDE9RO/+FccEDFTr0LhNz9YrVex8+Y3P4mWUhBpVTjpGX1NVBfMYRbts4cH3
lLkHjxfHJTOEVRzGMCY0CCgISR1whp0sJfPnezMCPUPG22sZJ8yu2nKBaj93mgVL
+yEykbzTAGShMnZ7vaNlmjquudfRlVq4lTj3EG+wUl7MeedIkt4Hbbks3Y86p5H9
pBWW3+FmlUFazkfii0JkU893CMHrTV6g+NYiuBVmUTYxsjrsQozWBAsxkmYPRDZS
aSvJiQvDGlQMfEm1dBlQBAIVGvCTB9iVmWFYx52GloZLm9fed0meGnV3dgxio1mJ
ceVCdNcIZm/z0N3Eozcg20obp8WzRAqHy4/w6U/NoXk6ckmgwWyzzwt/QM7hLtuT
Zc6mXDz8LRG2WTY6kvr8lsA8Xe+9JSBBQghK+vgHAJ/51+LNmuqW/73VXi8nIS3/
NCd6BMND8AQ8yGPcuzNvihr1KOfFMGjHFRWwTDwKmZlRXMAZEIZeLAx7urth0Mdk
+82Py6ZH/5YOxq8qdBTgPFs/mwcaWiV6G7L+0N1PRoeLZigFWV3x9PT8cML3rOml
sOMYFqPUndVuHPipTLM5ue5XUaIy8ePJ+CWnUpDa5CY6ojdm/zzHgrbjovQKRvb3
Max+XkiNxdJGHdWAePPRH9gEa7rn/+J46uJk6Bo5KpypKUYo4hcDoAEGQBDG4x2H
wfhqkOR0oIELFEY3zOelj6ZwK18cD0Ig6WkOFSpdUOb4qzIfZUm5P43fAOHymLBe
Zu79nPAutDzuGwEFtGfajFNvAI3R7Inkvoqmbiac15U8kyH65zbrBPhDEurFjsBq
r23RPlCamVJe1Bb5thViOf/lidLkNbKwvhKMWnreQuBMtjTlaQFxuiOqRf/I0Wfk
RG1O8UOrofdJdc60qUsAo4rOCzCKsucEYqZg+y32HDHu3zf7LOkrrnURiBWsYois
ZH90DX5pWi3J2/p42RwNpe5I2EQ23aiZcwcVcIOeTZ34R6b1IcSnpryrqjPICcQR
sONDAOm87JMN4aZMJyJ66i5L/mRUyilKK0w4LSXc/gpEF8GLQwwLQtwPA50VkIGq
MhikYCxOJWxubEjjdBltVOtjKKJWGonDSHCnlWDy4DaGdEAZKfcl+mlZ3mohNrzc
jYOA6H2GKoWBHiqQQcddlYcQOyyIPEwze8zvE/rm7vpP7ny40dg81N8tQcWbmShC
NulDra0kIatRZ4/i3OjGHQCIGUAOJ9AJJvKwaXjqWnG61+OHX+0W6pM1VrcImpTH
Sds8NeW+STdAGfmYrYeKafiLuoWbWFnDxw3TGMZlZjVA/bzQ+4HodcrrRlYMXN1c
VizOpspNuQvc4u8tYfq5DZQtV1KZ/12LTEPrREiyNFvHdrQDXXpD8c6hxbWX3KZ4
53yPb6bGa+OtZJ0yamnTaQBVXWz+hyYyEpOQWm3oL1sAR3/TjtpO9c9POY+ImYGZ
p/ffEeSMGJhCwL1KelCRBg==
`pragma protect end_protected
