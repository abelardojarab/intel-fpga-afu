// dc_fifo.v

// Generated using ACDS version 18.1 221

`timescale 1 ps / 1 ps
module dc_fifo (
		input  wire [31:0] dc_fifo_0_in_data,               //            dc_fifo_0_in.data
		input  wire        dc_fifo_0_in_valid,              //                        .valid
		output wire        dc_fifo_0_in_ready,              //                        .ready
		input  wire        dc_fifo_0_in_startofpacket,      //                        .startofpacket
		input  wire        dc_fifo_0_in_endofpacket,        //                        .endofpacket
		input  wire [1:0]  dc_fifo_0_in_empty,              //                        .empty
		input  wire [0:0]  dc_fifo_0_in_error,              //                        .error
		input  wire        dc_fifo_0_in_clk_clk,            //        dc_fifo_0_in_clk.clk
		input  wire        dc_fifo_0_in_clk_reset_reset_n,  //  dc_fifo_0_in_clk_reset.reset_n
		output wire [31:0] dc_fifo_0_out_data,              //           dc_fifo_0_out.data
		output wire        dc_fifo_0_out_valid,             //                        .valid
		input  wire        dc_fifo_0_out_ready,             //                        .ready
		output wire        dc_fifo_0_out_startofpacket,     //                        .startofpacket
		output wire        dc_fifo_0_out_endofpacket,       //                        .endofpacket
		output wire [1:0]  dc_fifo_0_out_empty,             //                        .empty
		output wire [0:0]  dc_fifo_0_out_error,             //                        .error
		input  wire        dc_fifo_0_out_clk_clk,           //       dc_fifo_0_out_clk.clk
		input  wire        dc_fifo_0_out_clk_reset_reset_n  // dc_fifo_0_out_clk_reset.reset_n
	);

	dc_fifo_0 dc_fifo_0 (
		.in_data           (dc_fifo_0_in_data),               //   input,  width = 32,            in.data
		.in_valid          (dc_fifo_0_in_valid),              //   input,   width = 1,              .valid
		.in_ready          (dc_fifo_0_in_ready),              //  output,   width = 1,              .ready
		.in_startofpacket  (dc_fifo_0_in_startofpacket),      //   input,   width = 1,              .startofpacket
		.in_endofpacket    (dc_fifo_0_in_endofpacket),        //   input,   width = 1,              .endofpacket
		.in_empty          (dc_fifo_0_in_empty),              //   input,   width = 2,              .empty
		.in_error          (dc_fifo_0_in_error),              //   input,   width = 1,              .error
		.in_clk            (dc_fifo_0_in_clk_clk),            //   input,   width = 1,        in_clk.clk
		.in_reset_n        (dc_fifo_0_in_clk_reset_reset_n),  //   input,   width = 1,  in_clk_reset.reset_n
		.out_data          (dc_fifo_0_out_data),              //  output,  width = 32,           out.data
		.out_valid         (dc_fifo_0_out_valid),             //  output,   width = 1,              .valid
		.out_ready         (dc_fifo_0_out_ready),             //   input,   width = 1,              .ready
		.out_startofpacket (dc_fifo_0_out_startofpacket),     //  output,   width = 1,              .startofpacket
		.out_endofpacket   (dc_fifo_0_out_endofpacket),       //  output,   width = 1,              .endofpacket
		.out_empty         (dc_fifo_0_out_empty),             //  output,   width = 2,              .empty
		.out_error         (dc_fifo_0_out_error),             //  output,   width = 1,              .error
		.out_clk           (dc_fifo_0_out_clk_clk),           //   input,   width = 1,       out_clk.clk
		.out_reset_n       (dc_fifo_0_out_clk_reset_reset_n)  //   input,   width = 1, out_clk_reset.reset_n
	);

endmodule
