`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p7WRdFPMud05xwIVX+2OiE9eFTFjgmHoYaLvBKI60oOG4zHdor3ITbNeBtfk5x1E
XWgvQo0QbAev0NnBS+jzgY8ocLV8GXPj0TDq8nWcwz+GoyBl3hwORDgCStoRROqW
ZQObar50rOU/yNKXW2TEZUaiZ1nMdElv8ndjVlsGXdc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36320)
bzJtaRDclyR9hXNy6fSHZGPnbv6EVrBTmJ66+9upz3MZMpkjIfSxJc8aDacfsFav
9cNxCQCWEN2hzN/+d0WtM33MXlAWuYjaInD0a8tBORmQlGEGdPTkGBHYltsbU/vt
6qmSS3enRXA8OiEdo0NOjArJQpo2XtB9Bnaq6FSgFLZOMWAkj8/G1wJhltPIbqVF
mal89eID0DVP1XEJmBEiBdzlkKaweGzP8isuGU91rq2e6Kw+G3QPq/STWBLG/0Lf
za5jIKk3iFasL+5RIsfG8ZneFRRQG5unSDDKvTWfxH717/o6C7lyNXtKdRcN/axx
pmJUL3968T47RuJ9l5P5Xq3uSuozeQL99C0DL5xblfeE3iy9+ucgjgQSa8h13DzR
MLk9XNEUdA5HovtOwFOkxQ0MtsxSdxFLGV3i+d2Pgh9cMkqvhVv6+glea9Dk2d86
0LaCl1bal77MadDnz/vcC3O2honSWk2yXH78L+GPyKH+AooMFp7RTFCTBdbCZYgE
MsbpEpsH9w8RvqS+cfYKlosH92Y6F2NQxV1376zOEYJza5z042XRTGVascUIXjSr
i/3avit28Ql3HCWHC8DNP8Z/mmQdPb3DWN0o7+IPbwjJNtHqOtkHx5951sVxXDQK
3+rrlom1pjRzT4q6cJ9poPGaxj4XmFm42pPdwYfQp4wXe2itJ03BgF7sz0p3L1Y8
/H7Z0f+Jyamz4oGLjdrrItDb79JfRu062XCYrbuziuJMCxQbbf+HOPdCI6EQXknm
Whkm2f5yHZvrh8EnM7mOxUwtsz14k6iUzLklURExRFUrv8+HVyb1W+vo9EiKxjz6
zDJepQ596ZAmce3wpj2xtZfO8r0lh0QjkEQBFw3p2YowpY+DvN8PGxc1hJ5SCh2z
/C0hsfxNxv5r4GHjkZHQy53931lNzSVZ5zZrI0MZv00rRoEZ4Nnsm9M/P/3kkt+S
GLF8NwZvL3RUxogRfR7URQL4LVWE32ufEShYEEgyZpUEahMKEMo1iHJDd0VP7FeA
Q6tYeprvwdO/7pACsAbFlBKZiq+5zWzB/LxyKw+Pv3YOtIEFnUgVlKNhpE44YhCZ
/xPDxFAOezjd96x+O2gyB1c6Q9V4zAGx342EIVUB7T/6/AjY/MkNdfjz/RWkvswn
MGdHaR0kypmQ6zPTsRoK/bjPf8bYb+FWiOifZls9niO+rV4rnFjaF001J3Kn34k9
jpxKfO5by4Cx83Ig8rwTqLebibMMKEd5e8KFVLkaMzczXHpUBblcpST9YIBT7qJZ
urLRpaI3KRqzJC8n4S7wlZTw9tKROuR7lgBPsYo2nQprRNbh9lj1UhXJr4z07hHK
nxTMRvjtsTRnfqLKw1NzXbZVfg8JPe44OT46FqEJJ580rSUgCHGF5eYMZEK0tAGZ
g0DNBQJlipc57dS0aG3/LNqYTKr48/oAZuXiE5vbY+COEcWDxhcMICWK1KtqIhNg
fQtXusMxBlKNJwWFM1RIy0X6vY2qFi3jQVaYg+GerTtLCKqdFhaWSZf7ssg9Cb6S
4JLdHfJ0jC3S9JeH9sdZ6oM4YrFoxPKjeldZPeCgZ24p0RDzOnQNte+5blZqbeV4
h8rI9onupHn4RK9Gp42UQ+JG4L0BRtEi9xR6WcsOJ2Pq3Ysj3vr+ZZ5zA0JWx2gH
If1z83QO9v60dtXDEJ6r0X639XK636wzQ9taAYmp4y8VFd1SLXVR8MuPXhAXWEdR
xUkSaWIbJrWgDGcz3wOQcggGCzIfmbmGD2wgJqJcnQ6nTRSN3tZI5NitseqZD1Jr
VrRsChrqVI44YXrwjaSmKrTiuCfaOyF3fMr4vSwyHxnDQLaizDQCfRiRS36CIeKA
dLJd/nqXNE95lBTNzW5N/q0hYM5Xip/s4vbsPxso9N6eZ4h0VCGd2h1D6hgUPcMf
APNZT14GC04Vr2KB4OmmFNvggMyGZ/zk12o6yLDrDSJVOqSbZDXgnQBb/fERtFDW
tbC6SxRmM5UzagF7ICnTF2mfSsoKoQaX8sdBYDVD9DvXSWnqBz5YxZ9jlD0KES1H
Qx0ndfhNdnOdoz4vBmLIHcUHjMHrEcC1HcjYPZRAd/uYB/NX+2wOkT6lTzqUPeZv
eKOyeTVAhKWjG3aAvExW3BBKv+ykTXVRH9tmXM+gElkCVHnEtsW75Rm/RUUs/Ygb
4F8lpbcJEGX00/H+zk+apQuug1uy7+BfgXXJbtlPx2WuLVWQ115EEjEhH924SRzh
TZ3xVFQXZvmQAH3R14YnIuVofFzHFstNSgyN56xEnIae+roeNLX+Z8gTX+z2VSXf
GSG88XbdgG6zHUY0/5pvOLVg8CB2blXuPxW7uCstqck3xHRGLqFRDsoMPgJiuT5r
tE8fzTRyppHKew9bxe6uiZ+uneCyQRqARxv4VSXFWaQ9ao7B7HHEwIUwylKY4bdd
gbNsqBjAP7X/e4SnNeN3Nq2r/xAONYk8lcvlhMVIaZm2p67ZWPrrpTV0N3wjFHut
z52aUgv/6rlwLVzICpZNlSlGwQE/aQeLQsgyeLGpyUGHumtKM/0dJdJNRL+X62dj
Q0Yib2CJkUVuOukauL5SUbfDov1mmqdiZemOTBBovXYl8JVBSroC23Z3TOJqN0cP
YykIlopRye90OzjM8lmb8gNXUPYQv0lTMiG5m/VCEFPycr2SQ39NwsrUh2+EN+Bp
Ean6ueVrPMTWqSg1cASRE+OfNSGkXYnNEeilf1PIukgwXz6S0+SH1PrblSsLay1I
U7vFh/8xlUdgYhZenuurymLiuz2lTZVkP9y74XHUNGlguoyc1SehqABcBgbC/GQH
ps0o3TNJ1Lee+M9WFyf0UQJ/k6LJz/kSSKj/JCRjDk6VvjP3T8wG5obuLcTezbMl
jnRIVFLlAohJjcob4vXOW0vw7nZQ4Yc2sB4GE5Qs7qd0j/wqVjfDcuO/c/g7FXAF
UJD8fubzeBqNZrzIsp46b1Mu84RQkZoOaR9jSXC6gSprLsduM3lv91M3E005QwCr
Y27kJREkGnRLXvhra9eSWoaMywW2IgsyiTI1ia+gSB2N3kTIBQGKLWYfBe1e61Ju
AWFPwxIv747cqYAU5hCNQ4G8C3ygRYbH7hBcvpRQcIIg5XJif5nZbkcru9e5Ev4z
mb0/YOCp9vghyb3QtEN5w6KISVjWSxMswj2kxtmhv88QnwxM7Dzdf/phnNR/Dwos
UWXuBd4I/gEjHaOMyorZJ5aiOQoQ4F8jXfzPQiSSsoAPS52Mww/Ftqw71eBMM498
8FEyCJsALX7RH47EJQxz5Vr9ngVxubbcj8O3OXbRJJtrrC168n0S89d6akLT8/yf
M0Yhg4l1eX1RpwjpChadS2yP91mCm0FpesGnITFEfQdzUtelt9zhXwxRf62oN0g2
jwtDC1MJu9mI5LWQVisrv6Gm4KefrQhQjl0ZYAFnHgOgn/fR+QZulgYLZ4OdJy8U
7LUZDw9AO9nnmXWa8B3OSKDyUHHJ98sTgQxs/LgSHOTR4fpy/grhsYT1bhELpXAk
JHZd2pX2V4DepVKx6YUXsjr6eN1BCYDmxHwpanUobApGpvXgKGPN4OZmyp1RauM/
t6z/cAMqz/1jJcnOu93aPxXUqIaoU7Swhzmp5J+v454vCsb+TY5I/j9Lfh0IQfCh
cHPPM7zjl77nPU2UOsweyyHoUvwL95/+iZcawQTf7dKCnf/dgUzwuM6HLnRHN7UT
DB9cO8IGi1McfCwcb3uB2m3yw7LCg808pnnVlfEjIfIxPgmiCkPC1f0+ewQuEWMl
k0thSi4XhRoh6YLWsKIHOxQDiKxQDDAHak5SZJ44gqD5TVFLty/adP4h65cwWES5
idiEkfHiniLbHf35CyTH4axfAy84RZeRxUcc+y/UQTjOsN7Wh1DKFzvU5Ja3Qmiz
SvjDWO1kJmMZZvK+M+Fs+uvkX6joI/LnVVC1xxTF+xcGhNTFv0+x3v66f9hI6Vgu
2Ul7GRdkuO/cuTCkdz7f3KNptW5cG2KR5HsrCPCc1bp8iEHlPWY4/n2qCNgq5YRV
CQA6sqxk2HH8W7oDV7rj4p1DFN7CXWSI/6c9Mwo5h43XOvff76BDf1gqs82/QPhm
mIPn2HntcCBpETZgLOdniY8/jvxoDPqk08hi+/H+RrreOkwPlV9UGWsePOK/NDef
1xezZuyfI/q4p9ANoiDkyHjwIImAO9FR8tQJQYQZx3aBK41uouKTE2FeDPQHDHFC
2cC4lejYPZVIPI0MvxI8KaTwXzO4VNkvCI/tKGx1Ikjgi+BVvLJLaWn+V7vSS1fM
X31NqLtwe6YQ8gX/v/15iUJfqqkbjBBquEDQu5XnJcIUuI/yW4kWPCustBlrvhIZ
6iWW2V3fKULELUOJG6zi/WUWo/9fm8TdXq2PZ4C4NoQiWg8LzhJXiVo9+ap+ruJo
+ZvOBguDL/JK9Oj5GcJWSQIX/DP6AjT5ifJpiTvDM4UbOX8umjonbCqGpdmreXq2
pg5O3GnldwbPCoe0Qn7Lu0vq1GZRS3paWSJMdmcFLSZlzwH9tjwUSFIEDcsqrnnS
Ei+mm2oui+RdBNopvaaxZjhG0+Oxw5WR5FEUuV+tGipwJDcvXnbw91znRhy25paH
FPbUDI7eZZV/X//dgJAweCu/NlfuxecWbBTQsxLEVEJG1WYMKLCNhwVcN73I7/65
TY08z6f4v0QnhzhupurxiKKpGmSRBlgUYNDzLV6lm6L8BaTclVcPGebXN7xBd7IP
1j/TtUCQ+SpiK1hyeQiB3JTt9THoorLw5bXRGPhGVJ/UVzVr+10myc/xF5n03qJU
UriDXZ2LprUyMqaNOIXzF3OgTUMRQhWnOcgUxzbirZ/oQzEC6G58fJZK9KF5mTFw
0a1w8uTVGw9t5CpJN2r9PVjuhHXyKAJl5+UJo1xag6gULT8ZWSoXqFh4QYkIqjwW
c3e9xrCM5AXIyaVsMuWbvaoMAVfOsD76NnVpWiEXDdcNdMofDRhwGs+vG0sWOR5X
Ta46ygDLMydKmXrym+9ofXdKUWzupjZ7nI4M523VBnjONhlLl1rfs57mTlQCpuoB
2AKfLNIPhOTbK3jXhYb8w4APOgroJpiixbJckSwt+kHi6bNkAWwejl6Wnx0u/j1A
B+gyuX8afqicXsBsx7xKJOMy2OY7kB0K+J9oj/pUrxdggUfFR5/T8EWS1/swwxCP
Z+j96yMnzLt3EEydehIflB+TU4MdziMetDPW06uZULbWA7DNf0V+CRxRws7FdhPN
vyInqvx8rXvX7cvcra/jumncpNEOzMk23uqHcNPmFYt4wFLuX1ioeDdHbhHYkvgy
CSxz2f+9vzVpTGY9nvc9of3yNEK7fu5mcmRNRngTzc3wsDsROg4NBPYFd0cZ4kL4
RIlMM/9u/2Tn2gBrusT+aMBbp+2akoedKPfTQEf1jwknu0Y1pRN7ABvhBA8NZIlE
l0i3SWNN7rY5ZNsQ1gCJ1jSToOyDFZp3fDpLvezP7fZHxRks3HLJO0wduWoW68bA
WctpKXAHp6vmN7T26e33NUzJIBOO73cRxdw2mZKJ+5G0TLZGy/Ji/TT686EMpsT5
+aLv0w+SZ7ExzqyHPLdfRmcyBAG78jTgx0oTWIRrSIc2ozZ4hhnYacv2JaiQscDs
Vmydu9BP2vHo1Xi5nCV6mAHxU6kgpuNqBSm8F2df2mC8g6If1Tj8F5r2i0SKb6kD
w955Nww6wL8IKP6LowAEQYxngw70DvHW8ebQ1wt4UPjiFxXGZe91lqVL1P9Tt7K5
b4bYZkYRyaouOdte49ezweQZuxmtlVXQo8gmh8MQ1UbJohJoPeDNztXGFB76Tz9z
1Z/wOwWShC9rdWEjJbXlk/R2SZhL+e3mO+p602cHYxVEHwB22udGxtXMSrfgGY7a
ASeUYv5qn/YgKkGIP03dpleoql3yYZu/LsuBe4CWbcnjX2yQBVTMQj93aBX5Y7TJ
aJRbn1qdRd4NkXy6+4slddPoQKYYg+8Z3brB06lzY3gDjWp2bi2nrnyvJuU9qoPt
IiZD6YjVoQUoyIVxFQnWFpgvZOE9VQOwZ+TfJV9rvX7fYhq5MOBL67143R8YrkSr
oRQr7cCPbxzCJ71OFlGghg5UDzHM6k6DOZ/nT6QfCyHKtwk4VjT7qkWLxlR7tU2d
aMWULQBNK15VItatPPF5Z3J0poa1IWly9sF0CYIqWYrZ1QAo2vR+BNZ1HbWirYON
xtUi1LH4a00Vmhg2auY1iNoUAtDtB8R7WlUCPp0z2nQtF29CgW/x0o8BP0bF7kfg
tL34gTVAvyfwVh3MfxdGsK5hUkfBiNSd3kTODbD3nSEsQPP1NeaZpADTeyO0hjA4
zUAEIr2EN1qUKDVzM8jtlYrg8p9H5EGfW+I30dh6KdsZpDGk9mTNzARvgdkiuGAO
rjZrbAPniylB8CIX/hHiaqvGgZX6fuiIWBoiYyo+HjuHaKGjYctqiNZNXld0wqrw
louxc5c4xBsfGvoNf5uB5Sw8sC+Wj6CVNOwwpSt4FquymfC+2HJJFy87hbI9SQur
4p/2Yo70T8HbKCxiHgSUHDVTKIncuyAJ4K1TJig8x74qTkCUVSas5SRymf0XTUIi
TDkzo6ZRUHH84I3gKAgC/+d27vr37jBD24+mFs13LjBGEttk9IWBBdn9dKIGsxOn
YFDQSbtvfZ0rb41RNdcJBsdpf4S9pBggV4goXkLUZOhGruQdP5CZa2Zg5l7BYMYl
Z5mPoMm1DEILXtsm1L7Ay6wcm+5uO8mcZQ4/zvLOHcVOwd1Nh114k7T4xcFShCYS
oMiXusBNQMFQ0PaSuZOrups4c/c9U2bYdSYS79LYdD7p6y+g+o6FK9ka9Iac6mI0
xKrZh1vmpvbyV8KwwHEl58aBnyL2Tj+YB5cSa8JwjOplluV+tVHRbip/V8J+Riaf
NdGd77eBdldWzZjU0PHWnAaWoEStLm3qOWGGy4JnAD/zH0eXIT5YYawGvPGOCrBT
dsvkK1B67dIkXiiARE/tiYyx6qp5NLjZLjrJUpUNryKD2fYoc+dS3btDFibOdRCT
1R3oGz5y3KAvYJnHtHu2jAoc1RhNZsVnSUHxRZGw6y37VHzk+WRfPQ4kylgNRX9W
t+IFpjlF6UzcbJT8gqp1+d5td3m532DPQm82642CkdbSUJcl3YqMjmM7H9kGjkvH
V9riLhOeuqliouWOkbxuzQjkP8CDwxbzkHbFSrlI0zskpBLcsWJvibpiltT2FboE
7Q5WQJ0vJnHc1jqIdNfJuASFoj+7rpQYODbwkyrnosPPiGXfETR3Vj7yxZpvAL4F
JMBIiVxuoBKwT0e64R8/fWh9wSq45Bc6qFvusCT4WVP++CTSUAlJNAche9tgXU2B
F76VcG06ixZX8DfayafG08vZz6ObtfOacp+xc6aTGG3PamF//zQSWwj6SHgQ6rB9
YsXhUygmy0ewA3Jn7XbscWcwzejQ1M/Uv0ldc1jR+bjo+7ZGP+dZ8QUNBvV/Anbg
YdEl+vIQtkhZXstFFj12avfe27zqOkTIaNmVVd+pOji3aePQJhCItsFZomLXzDsO
DHto3vSReAp3OifzMDwjq+6ewZjZEloTtjJoOutEIGiZ/WdmoYCIbxxS1LQyNERU
iHBEkoUXj/yw8sOO+NBvm7exdLJIPqQULgYtY0QW2x6OLV/ztJ8RjikvO//omPqo
scPvEhPajVpEmfUuDc8v3aNcN/o2dI4fonSevstkkJsF3rNERIooB6TDUaKwdi2B
XWRedMD+3C3WRZSzv5LpdUgePrwxOKnPsh5GUqRTdkTSO9R7YE7M6ztoVDi7UyLn
ZhdbaXUO7HM96M+ONLESSrVQ4DWp+chyiNlMCkhoALk39j/M5+dQQLhex9RRKtVK
eZqb9X48gugZ6+AqYLFH4hNit9T1j3E+zcSEN2qHVPu2k4Jh5WFOxZS61WqhmyJR
6EsP8DwIdnPGsImunQrqH59b4Bk15qARtDVqMvOrIc2A7yJojpWBPVmasUD//XiE
rsE26wLeoarrzVrI02RoTaBWQzzIYxk+GTgMZE4+UMorl85j0HHa3RWGHO8EkiiP
3WnbGStwk43aiPyrbvYrfUPe5Ovz/r0PBlO7alwH0VMWqLcz+4CZLAk7+KibElRf
WB/W+HC0M05nFgWlOln9XgseCq47EEWpI+Fgg8BzTltbp7y5l6XUpXTkZSOVbTca
cCj1jMnSOZkybfNSLPcbLyswhJeIQkRSobBohEsLLlX0kB6JtQfdhQbocaS4B5Tz
kSFMc1uhCbGGdT0WYQTHxchbo5BzpHg9h1vZUTIG3vSqtwgkJS5zSOApXdZRgxzr
K0VmYyzUHg9+uB0ghaBqBMPvcTdN9akih0Bzp8Dkgdfo9FzbY1kq52eO+mMph1ua
EIYiix+wasf7pwsZ9+OGL2icnKxF/xwir/OEtLo2YqAS+I+Nq2AXWIws4UnXb5bS
7HaVW9Snj0+cMV4ntxCyibReNmu/MS9wbs82Kfh0n4I2RAaeOnJ8hKXkxqgSyBn2
RIT0B3TO4uyuafFX2Lnj7D8qfDfhjNeH1i3iLZ1JGb0TKK/vX3Uk2jeTkOqbAI4z
LZ0w71kP7BBiVVNz3I4dZD9ig3Dq8M6avbCA6ONqEDjbbBfAhxYqpaoc3+cEku/N
V4x+nlXsVMtPJ/GxCmWE/ox1b9hf9Cdvchm2sXiF1zshd3odPV21DddrtY3bLRJY
1zdyO+WFIniCtzHSZg64ZiFXfIDdnjFWRbLn1SfqLyz6RivxkTbZkUjD5KfgzSHC
IHY7i5kXtrAF/ZXofNo33P3DeZyZoP1J9n3t8BQ8mPAH1XrkIJE+9/PwY3ARtLrX
i8oifKJ+DBZnDfeWSEQIhM22sPvkJZEjFvZupYWmfhyDtm0kMDLVCZxMivqZ7/Wx
x1jm2tWulxgEKjDVLUhYdJFhqKzTwcUzCfNE4n9C+ettMOJMvlHaGi9QQNFyJBr3
FseM74Lm02mYFT4BFyYRdYtF1AyJJT5WQ7e/Kv0LSTU5wt23DSjVh6laljZL05FG
pXQDfo0SlbaJHKe0UxSpx398p32slYiUX5IbPqR9ZejuqFpM15PjnQMVgHiVprQX
iSWUVjfPjGRyF+3DcL0nieREY143I1+e0LMBrvDh8WdcR+RyhnIUD+r9tNQQ/7CJ
1LfD+WGiOIPPJKSP/q05Zz7r3YVek9TQRWmU2Ar28xzLsZj9KFyuYAAIGCwYFevq
NRhR2ESye5jsmpuY7kLXvCTv8BzPOpDokLMtNkNJo/88hwMrG35ZMYu38gmzPwrQ
JhTfcrmwDb8a45LF1XnYE6TWEPH+G+CRvyvp/GDtdlbv9d5cJEE4nMtoxVr1ZcKK
Ip86bnUmVofFxZjXYZnfWzFhQWoDjEh0Rh/XTYhFhCw/DmUvrL9xUREkaxyi6fJG
4dqmMSMM0JXuwhtcGDejObKjArV8RMgj0xej0QbuY4hE1DoZxrnJM1IJ/1P3hEfk
0V8yWYUWcQ9vLvmZ73dd5/ozB2zEGsfhmxfwU7OetYqTmPQ1gkzGRRe+66MyX6G8
cF2u69tYgiL3KyF1pX1LCbXIDksmcworsrY1ih6wmHzH6598hOOtvuar01IIGbZT
Z9+tJcpmjyaBmQNFeA4knd1riPlvZ4IJZi14TGbwbupp2QqC0PtJyrbz7sK9RY/Q
333VhUEmoAO3EeSErXwqRzwjwVflLu4heRYSpbMrFmrsOu9HgcB4KrFFfMQd8GMH
yfIJee0gMNapQhzYi9wWCR/Tiu4k4wgSzo1TtPECpxsbrWvajU9KtTdiU4QkRYG/
Sb6AMGVaKB5q8IG1IaBXZxFfWDqfPyRi6OQluFnDSx3gXp5zNPsJ+C8GQTJqBxe9
Dz5TilDBlwVUjIijEKCfyMq+EuAcTZK6W1rfg0l8jevp8kJm0QbNQvaTTlce8acU
TsoxjPgue8ceQZ9P3QW6rJ23qTwsTKVPzFS+ikwTvDswrA5PLbqNLTY7COw6LiyR
xUe3baxWNwgKf9aICvV9TLVarXXjNlFwN5XdV+1INwXXATUHddyHVtnbsFsAHXQw
R2E9CpabyE9Sa2Cq7I1tCtfOB0mEx/dOepDHgCESdJwU7N5ScibO8IJZjj6G19CE
tTqH3uQYiOrOsifN7geXmips/W/nwTYMmCTMiVtP1ROfWcrvCDwhIdt25cHWoThF
UgP0wv9pwQ0r9th+r7dPb7nYTqnQ3l5KUCBiXXDAr0WjfqwNvY6jg89frloUDXH5
rPyV7AxeD4NlSzanNDDwhzSA5fHjt6VNW08h+ZiYkyaBGhRf2Wo9kFXn9KZgTNfd
M467BMvC350SAP9YklsIqYZ2TYlTUkcNDKvg4dxDwRGBvtGwH7ep+yDIum8ojcck
EsMYDsBJuKadkCC7+cZhpFukaAM0ahyXGQ8WcpuvKIqPvd7q85rWtH//juErNRx0
4kpB1LrKBRo2QwL33+McelIaUZQLr5sfrS+Vj6ba8nZOy48SijnNfzNA0P6e8rJ9
cIIOeKrkDHW4Y8HHZUCTWMwS7ZnFgziaJKL8/ZPUUFqKepRcoLGmV9PB86CrqKXP
km537LhlMWvxc/Hoeo4igjjDwj8Roq+y1/UTHCq+kcEQ6QPfOR8imY6VrSRvPQuR
5NrQcZZGIhVZTjAj3+4AzJBPD0tN6Bjm1W+plCK99yCKkCzQGTXdTxl1ynoy9hhp
qZHdFLBCLlW6HH4kUmGHxA+5PNzAGnL9ijxIKplxEZrcsxozX2U4abLqS7Ww6JMC
BjqVjSTgrU5aUyoUo2EeumxmWEqec9279+MvlSyOG8SrM1QGvWOai2zxUvGFx3pA
Q3Ir9Gg6g0KgWzWkBvHleN/aUXp/lK7DLHnjCEG+orC07v/4ScyW5Rhgmd+LsjGH
dYukHEPyDFZTZPk6lyGC22gARJswA2KOZlA12bDiIEe56qWozE4jh+PbYmCqil4m
U3kup3EwzhZmKI35nCg1tj16epZo1ip8FE7O9007hnNczU4bG5Y3mrlUOfS991LJ
Vx7GtGyFf4PKfRRqnsUOPO/MF667nhEGym/JDvqtlYQUnQKcnvMmmUhu9/hBVi0Y
94MtmxXqwaVD8zQStxYrFhkoYvhm1Z4HigjFCkOmGQxa0qDaLNgHBCB+krCHMV34
4MOMA2uPmtJzPT/aSYUQJeN1n5NT8TJdf0VKCV5RtQIbyipo+BNnwFOm1tZl5q/Q
vbtKvRHwfojJzsmWsrPiI9KU3YXz/gZNB24eJvxnomY5TEJwGUaSrF8AbvDsMRYf
aLIsnVxsphUI4qRJ9KEexgUsgzdPvmIcH0bebhliV5TB8Vn5qcFw1cDf83ARvrlT
8ThrsBwJfYjK25UWSy4bYlGIZ5GAPOU9jbMcgiizMIeStCwTm4xFyawHw7MjR1kl
soVpyzgVc7R0m2yUCs3F8Y+K+DIq2+dlHHC32869sebEHo37S1ZH9CWIjHmypZnS
NAQ+rriPdHnpDwFQHvzhjYRWtsFsx6r79BY7vgxnMEVVizI3i0MS5Bhp7FxAKUz1
3bAVvJxnZxcnco9hKmwXEGDh19bUnZPP3fN0E5P+BSDNHWDUIXkZDxbJLnSd0OHA
7RaH7gCIZPXVT1rfgdLIlF+yim2wKWCX35VAZKoCSWAhq7AjQrcQJJGLkLB1dRau
4cOIypkU4FN2rv84ERcohA+8P9ZfrZl8FiqfS7yCXg2vJHg2DfVrIg9PNnkVhHss
wLBhSBM8JQr3KjovxhQtqhRLLBiLpQrbIjsFKl27RoSjYcvI1DmR9rTLSr7GzuJU
vwPVxF9tMjMs56Fso06awIuydjWg0C9Zaqlfr3Z5yl/JwaAK6Lh19LgMqL+WUp61
hmiXIvwC3xgB1ICPNiThODX9Xx2PKOPDeB507gqdULzeSIPzFg2+lzryFp2QkRHj
YCxW5Xjj90k9rYSia8TRm+AxhS3Ff/OsA3x8uL3jPPztWTZ8IFF35JrKF5eW9Tij
6psDBjmuTQLI4WMsv+wLwpEQ8ZNTNMQm38r5GITBBNOeQItSf+mmlbda8wXX3g1U
c2zzizmiysWiYgoM2cBnm905e6xPQuZptY6O+G1CL9TAM1FkEAzbwtfD2gE60j5j
7OpDItAtPMpZO2+mf9/Ui1oQeFp4EnySc6ey321KU1KhAxQSfysekOQQLgKDlulk
wHKF3wQMtGGnYqaG4Bqg2lUOC151uqzT/p/Fp4XRmdR4e3VVrVlW+D4TRjIFFjt5
rblXGOAeRb6uw0OletsPdcrNDHaGtsMKwgEPoAp64zvDroAn5yJyWe+cto2jzGqa
LHmwxGRWu4/LHHCP9ANt6E58wXGTd00JVSW95ePnxbxYFaFtRqOPk0vsswR/YjPm
YGyuiL/3BmPgtnE+0wnXWTjzWVa8lQc45LHp4XPpApB/vL8hoMKbD3gOYIsQYS0J
mmaaZbcVEwks0VKSDk5QgY1R1BXQjjx3hRNr33Bf59IevFDjZ4mgdh2ee9KEkuvy
9Yp6UxMH+RM4RIBQ/sYkQgVvnX4KSeHmi9tkRWAotwhfxoXArprdbuv1SXCL2aMS
T+5RlrjM0VWA6LQVDId3ryvd/o5NC2fNVcqWDPiQ3dI7Kg8gTJgBHTub92BOWK7n
7WLyuuiveQxxPyv4dz2RGS8hNl91ITM4O70NtX4h2a0Rj8FHjsXFQtJug7BDorNm
sgHOFhhbarrv7uQJA5wgPfkd+Ztv1x6nxSJQHkXtevxCJ+ezCqZFLX4T00n+4dXU
vZC5/+BC/T+BQVmR6+5gNuU6GFwxMFe5zRY6Pa5totQyB1XH4VIZT7Y4nsMB7huY
WJcXWxcvJilxGNC3n/XofF0GPun1S2ocjsXWGdKlyZ9s83AEd8kHpMpPsx5JEXYd
rpQ/VOvlZc4iymwcJbDuJCeTgsPb6URAgWyCbhumMSFnDL5MbrWs1+eud1Scb3C+
sP0nAzYHAEz66WpBlKxMh+cx/GHTSroqDf3jX00er4PIClOb34v1hQEruFPN8jbb
zJcekdZDKr8aeFsD2Qtu4HAZTQs4hcpG+XtY0hNa34f+LL/QFgPzIXRuESREGd+B
q6TGxeSAoMCTzDFqnwNcX6eSddDVJBdgakWEAjiycqxVorL0eYS3ha65sjkt5xwr
WKs/54jFKp7RY1robxZyCp9pSZYu7IfF4aGyw/7KM8VwY6V0oC4YxJsvC8p890zt
0Et5JISbOVVQOXIDsPVluxh/S4GkmxSjwNfz4oBhHoupvQf1HJUTVQ/X+eBpDWBc
kESK/tHp2V9mCSx8A25J8sgWic4sHxapQ4etw3BCuQ0+XuLHUjKVgevwe2PxndE5
n12gu0bQfaz3San5Zzd/n7DRUoA/gmoTmQ0lWX1uMwN0B+3Ei8z9jhrN9wTKTuxK
0L8RsYWbVKBOY5juhCld11dEuoMERl1hirPK2CJ9z+W9gb/etfgtg4E5TkbuENMF
+F69Wq5zbTsmVzPdebIyBEFkQl7A3HDZAYiheTb5zLOvCUE0bp1qDgpD4QSfl7lB
UGFJLcqE92B3ybe8q/AR9zDMdYvtEkMSuZ2cOlCfwNzR0FQAaK130GLdNGyORlcc
fjPOEWGK8OxhVoEbXaUDz2aLZ1DnOUybWAgHgYsFVOnwuB0EgInabinCohAs9AqC
4jcTQriHmMUeiKWYLIP7oVHkuUUofBBAip89kX8VCPAdGkn2C3hYsmugS8ofc+2u
sXLqZu7SOWvDK7SdMq1KE8WIGdg+EtWXdMHqQGwho6ejvxWt3Z5mpoimxPmhGDKh
g5ZIH8qtuvO/BCmqEjMQ160wxaI03Z/jKw0eHOZ353koIPKjZ1TkGRbdl+JKKYRO
b4Scm0spykAm/EYsziK92tRbwsGguOySUxj1yiLr5Mx5F7KLml0TW9itJWO0jHWL
pH4hUb3+sBLTYSoSYneZ5s0b4agltIwYluexGzzJJAcWvN6R7ZT7UpMkU2+8ETWY
tsOr1SzWpOs6TP+NYDQ1bMXK11QAWiaF3917xN2P+s0IekpqerEiHSX7W/YCzmsm
6ewnCZGNywCPDw3tbTO+/hQ/yT70CisSUSTxSo3FGwQHJACDQKGHHIfbzudFMlTq
yBe/338OXlPLeBQBgTbYJRpOOfGU90dNZTM1viprLEAvcZ3U57RYiCI++bPA+BJ2
+JERPzwoYVLlD/ivLK7Nk3ajuIM68osVyh4uqH4HawB5/ihmv3ChncV5kMEwG07c
BZb2MG8/E9qcBbYOs/TwFaB0KmoLelmQAMJwkcz7xcYorudfVeFZyVo7e8WPcRnL
PN48tOkItBtDcKB5dmX6PkDp/zjy0gfQi6HHvNm4BlvoVT0kQiU5/3zeb/xxNyi0
dNg5nwNE3ktV8R+ym5fDRHIaplteEeE/WH8xhfTBRXpREszSoxaR3SUM/EfVTE4O
nFDGGpg6CWNQdB3B7yPF8aXaH2Fz8Z1GvG0Y0TqMFxCQ4ISuKnse+1HLOhC3Tk9m
JL2VPc34CBSVXFkUaNBp7KZnKYFngPsXwrfIp7TqSD2e9SkT7rdwL6h+ZziwZoKE
8X/7YJzrozCiZrzpG8u39iqAjZoqi1h81KsIs/CNEaQd+DJ9LXokWIW5J6KKK9ry
vb+duNLT/FICeArcdX6Fxs2ulWomMbGuQBCd8iznkp+4CiVrBiti2l9OxL1xV0+x
aXA1BOVmmTRr1aMI6VgZX4qN7YxCSV4EtHkUAeVnf66yNj+9B/50aYCvAOLM1+OV
MC0gEEA+abNdGgMECsAf29TVOwnQUxnE1lfFHabHFPNfNLaK7e30TMKfTtB6uaN+
XuuWhF1mh1rV9CzHYl/yTsNczdH4hUNW7xg+vcfqTfA8hclt9+jPOGwjK8ll16zG
yu2ZhNNiWSUFkx4rlvCx4i96eQNZcMy2NEMSVjkW8TWiiKPyYFX94d64R73Z2NRN
dZL8cBHU6ThPRektK8HWnTCm9CKdB8EwWPeohGJnDkREpUyyCCDmI/VmMiXN5Noy
c2sEfCvciFhr2Zm/PyYjfuVRR+cENtcPD11bSPkwxCx8djYslLxbvpsje0MWw0SN
hwSRid6gKGhw4k7oQJDfJiuqHckiygL07UC2UKOJNUpwU/w65qwIvbwyelSts2TS
e1Zjp031rgmlGUnmFnERei6ZT2puoQo22EPpuL1nbGEw0wSEecNoAVHa7KTkPPme
WdhjMzO6cssoQfEUz5Zru37/ciAi7CBMB/gcZuhtNCJvN8whXWsMu2y7IF8ogEK5
t93SGAyVWgIoSc89o1TArFfODZtahSMdy3a/X8Ra5wi7CpS9yfK6Cc/7W6L1zZzG
bAHhn8f5hizpaX9bgM16ZNFwjD/Lj9m8CFg7vIWBdYAF5TxAq5HhYUtfFZCdIUYm
qP5ATlb8vuxI9wNYEVvAiuq3dixkF4ycgibIk7Ws87zEVspULK0+WaL0m37PGWNQ
upe0p6G2KP51VDPLv1zS8lNy3eanPRSpI6vwVN5SnLKL6Nluc59B9oJlfltGdTik
cCRt/69xCAPFcfzJSK/7lCrZ4jn8LYDxCRrUUw4oN7n/sHyVYGcoMSn/0n1EEP7C
8CgvS1Dyu8ip8JvSFMvPC99oRP20lOiWpET6D5JuFhXEHVNl8TKH2n+z/i8empgF
arVtNQKmHOqx+4iLFN5wziqNBvcG4WwwV3E2yureaUOqAC1bADJTbBuTEUXcYrzO
8nHkBqULA5mG9vyOtAcV6bMka0yvtMVdZrlu3jIT0WkDloDLEu9K9h+QYDMkp3fM
EQH2x8Hos0OD9d+beeUvh7RHPv58MC13EEqPdM4PSQ5v5yKilws+P3FL2HEvBlns
IFvsKvIzCgH5J7pIEspPKtGXHVo7tt9EQlUJfw+Uz3FUg9uJfY5ql7w651Hwb9Ap
pcwoFrl3QR2fnVbKanbgwduXRu79dbpEaqbPhGjhDvxgs7/YQ32VWshrKScl2Y9o
h5frtPPa7Kbn4urO2uJWDY+37qL+kr5UucJurVxbytyOzknYwh7dHrivgBQSrXZO
b1kz5i0Gs9wToCi8qNED7mGiOP0n82eQCIMOcBmHmMBTN11k0mrgikNdwFeio4Qq
Rhl+TDoONvwy80DXDKXYZ0Pa9SYYyyD74PHg17NqO0EeY1rcKDwfOjTBsLbNgOMk
89rTJx362fFMN7zVxeOCCRhiaV4ulyYvzcaUpbXK0JhjPUjcCzh/uygx8MDRC9oA
BfkC1GjT9AI1mZEwVf5wQSmH5Pe+yjWq/LpREAf8UnJz+JJN24cr7PGUvBjMbSn3
P3kyVMcadCOSjCF8C2Wp2CTdsDVoOaOf6evT7Eaz4qocbTiSI1eoDB9EUThC3glV
9WM+TJWQt1m4I6oJzDSE0pnIgkB4I0wdme0ubjgPcFBsPNcUDQbDiqJkahjEKf3K
+tzZh7H2AV6NDj4yHo+xEGHj5y9D6tW3rAR+0jcXO64jJQcomqYUKIa0mi3WDaa6
yg75Ajz9+QXGSc0npIELwnnj4ZPUhGT5Rgwwcy9SiI67pZ4pv+ar/8Omed7eePMN
EjHyOS03osjAXz6XSuffgT2wTS0Vpb/7VvaOB6Iugsz2/cPkL29EUZFDzj9eue4F
pw57Y7zWGzJcYSBQ3C6e7DYE4Veeb/E4Ua5WRiNbMff+mxart1dmapo223x3H9a7
fW8LVPJFtqTaFWZSPfNGi8DP3XUf7Ds6ZshBx1QbjybFg/rJBufSuLwenJnVqUlY
fxkSXIRWGE3IHO6u5kJkuehnAZRAHOI+sbQClbPYcrKDt3S3ZFzklY60vPNQ5kUv
1J9t5M0LJ3sadWqgVeIDnQUOSYDKYY2itiFttrcNaLWcCAlX0Hv9/VQMIhrmrIbX
sc/FtBctVIty9hpfNoykH0ai+WL7J6KF6z4TZeBvOv0Ch4SRTzmg/grd7YDYcIgk
ZBGb7rjQN6OwpA3BJEhKmEmd1nuGyo+17hDqtsTG5hEiWY9ckUKA+ezlHsMldeo/
TMAJ+BITXKyBLq1uLdl/y8eZZvYLhmxrOCXKS/qf3fRbRdFE6OZ8dtRMyaDbnHoH
bKzBShudlqEpRW/D8RZExnf/Axx59aWXIKagnWqAkCWC3k+2akIFXR7km5guCu8W
r8VuPQF5dMCgSHRO2nv2kNQv+F2UhpTpvJ+GmI1PX68YPKCAGBoVncLpaJhiIet6
xXD/tPjJUMoGArZg87ovPrQQBikDEL5yk9WHj72Fs7VOQoUrynL44Bx83JBh/2/o
P4S09xODJgUYSdJCy3sr9LaJA7jFHFZ/e3UA447zcggK7oU8qGIHW1PegF5qWYas
AFtEWeNWRZ6op1N38Y90wARKNoPl9X7sBehCzU9yodFr1zz0SVRqYRD3AG9Xndni
6W+2iQT958BaDFSXaxkKXk9E953JqRXfrEEbrQ1rJ5EhRKsKzTetP0P7qEvTlmp2
o04PK6MmS33vfzOj9jW17MJ3WHhj7gqxSeOQwFe5fQnGSIVS7NmeZe7xkNr4Wmdv
saFnDIz797SlAkKgdEwWQsYw+v66XUgrOjOG3uP/xG4GmPZZ6xmP+TVYEnvCHDXk
hfM1Jo73AoPI3DGQdReoF/mAokt6ZbjkSouhED07bGLEIXEQQ0xgmJHPaac4Bf7Q
npySt/MQbHD5Op3RLgTSU55YRL+Cwt97BMY+LXKBHlRPOhYNKrN2bjlRIGyl8kBQ
/2ZJXGD9SCebVoSQ0Eq07k0q0Q29zGJGsxl93DilwwnbyRbVaFvPHwLvQl+uQ9Ml
xj9UkBmRjK4KF8Sx3QPDXCKjP9nPRTK3NPgv7tMubxT8rUn5I+FUHgW1PcacTN6G
hTSKWCWsJqv7LqH5OgHAJMWf2tUJBbWlQhWjdh6TnOoBb6Od2G724USQZWDyVmR9
nh/Q7caA/4lCK/Qu8B/VoBMLQXxDDBNFmE29QQd6rWN2ue2V3GappAWdqcYcDivi
9TVALtoxgybDomzaklxP89pfhYEgH+VI813ME2UxDbVCi/15JYfjfVDIc3nZ27XS
gwwbjqKaK5UJPWGVlse7mT7fE93emxqHnkgosjFY2A6/KiWYSJfYlxLZufrzNRqh
+yKkVynQYuM/6QrEHr0JHrUWakUNMWTEEzTkcF49vZjTk8Q731i4Dzh/axRGk8Rc
QWy1+FPO3FrKk73ALZLRNWXMvfeOo55Ia5Jopst0ZUP8muchs3arKF9gmwlemUcf
y2gIlXD95N2zFPdQNhAtnDeNjUEeaPaw5jPZ0SvKc8ukub1mpJ0o/39XT8O/49/Z
Vgj+xT73IqOaRDoE3IcEsF0WHghEKQsaX8ra9Dda9b/5AN3yrdB3ySvFOFJzJ9v0
43Y83N2RXBXjA4IeTcuzFBwxvcNZOcrIzAXIsy0IqqKNBJWwmmkM+BvRe9oCjp+J
nvSIN9RHc70oUiGVJFLuvmTlB9d3GHIpbCy5yGwpzBNmUm9+EudVkaPF9hSctql8
mH/PRNTkqJmKdXtzstwpeIh6Yj+R9GDtbtNAx1ILbMwHSmqleKbhRXln/mzAX+9N
hHZqSOyuqzSf957JNuLGfqc/nDKPwOSiLs9n2Q4ZObmVFoWGftGfNRUf6MTyh6cs
0APzE3VY31DDPGZThd8It4sFVjdZF7sNDy8A0yStzAvcJMoWcK1BxBtDK3haux0f
KeuT9aoE9/Riii+i7L3D97rWYV4PG/T7yRTgTiKbiBhRMd5c7j5WHYQ6CU9W0o5d
GyE0FxB8stzIB1ttyEMzxnG/dpWWwMssNXcpRvlXiBNSeExU8wtxW1lRjikrcSB8
N5lw5zLSaXOvAuJ7oChB5koGQJMpGApiVfrJmGRlBwVwDhlr0CVDTSQvglmoRTH4
axss3l+4G5I7Kkudbf49PPrsqdOY5VLCIN9IbaA/XkswD3CM0ByeAnDSlsffB5xq
8UPi63dO8s2nc1B47BmiUnNbyZ9olZAsAc67j9VXMOPC8z89SFP/ph33QNr/YmYr
86sZdWa8WfqFi0Kas+mwHAfOuQlhZbQ1q7kpSfto8mDcmqVH1vwHUuDQawzLcIxJ
a6fqnayhIxwVKH+XKKZ4hLiPZx8WSutoedS6axRy7ZG4oE6Cz1zgaYOMCm4A4G1M
4tLeK+ZJUXqofFOygiCaLRl/m1EQSgCIUbAQMjPQqU2dtclKNrl1/RQkxPjeAtZk
DUQ3yptfpiSfaw6j4+0F/WTnIVnYk4YQ6pnnvv8I+CD4hGWuGTbv0bi946qfNBnE
3/icEhuAQFkZs4Mej42aRD9gK2k5lOkl5i38KchCa5zDkpv+fKXM4yXHg4+9EOwD
xUneRalOwM4+YFLjkq+7sw/gtw5xCshI8mUzErog6kDWdnPdsVzH7aDzQ6/nU55L
JqyQMB1QFSU28QUmc3pBukeA/nuhhJO5/RT7NAoABKRnEqsR+IpZKwaec3obHSQe
364o8h4G4G6JKlTNm0atczomlbPB0yGrL6KqpcpOSIWf2nTCuvhIymrOmNGEdzrJ
r52zkzwOeSYenR/+NDR0MJFye4r5PylHw0MnQfcoHXyyQa/hYorGAhB8rz0a/0q6
XCplxSIZJAJkHcd7AJnRBmOaFWAL+gQCZmnlj3Rkvwel/hE6/emYbDpzJpC9AVDe
cylslVMGf3Pxw2vaaYx11wsZi6Pz36NatQhJmqKbXS5uWFjuU9NRmv2/QYScoSbG
rQ1nbWLpVTYSQ+gU48tpI/Ykk1Ay5osvcO5pOevpx5fywztE8qHZh2kFTL3wapUH
oMezsvK6ybdIp5zLLeHYY048fOREj8Tq6xJaQP+it7od243DqZbkjZkYtRZPYVCp
PyAR6/ihB4YgDxeQCMGn/Emmz7uVgzsnLv/W95XzkNX56vrCPBQOerdG6AOLbE53
1agh06rWCv2X1g+0UIZqykNKDGlluqbtRQknQ6osloOiSF1+q2s2tlxP+6ZWs1Z6
0wVJjzVmDB2qHS/UxZNBA/bVfy1YO3l7eyCexIJt7NSmXCYRN/h08stXodwAcd0N
2sHakKyGwajIINBzjTxuKCZit9l9GP+P3LxTO3tz5oDK+GIlMbd/3LWmklhKv+hi
Y8Lvp7od9vbFrorj+AfyLHnbKA+EALitAmHvIRBNHqEIREGGVzVBBe1UrZSw8qlE
vdOIq0bqm0mp6zSgyQmq6sp7EX+HX4VSlkgS7sCSkokf3IWsrjjxmib1N5V7c5Et
VLNe7UFOgLZdkVDtN5sara52RDDSNdHuHxq02boBTxS3ffTbhjKEhTqMh6lZVzPD
puVQC3au4Xhu9iymxSrtrIurwnxGc3pNJ5/M+n1fa+SD5+IZKUZTkx3xTCxZm2nn
DI+dJWijwnvJoimpFrqRYtwtvQrVrT7OL9kqOgdeyUPZ6T3yY6UhDhUnC4ffiRoc
yBpLLSVMJBrkhimLWPOalpsuQmXvFQ4w2Oxtfi28US8fbl475VpoxolvWiISOmDN
9yqabRSyPI3rzH1lF7dXU7jmVo63AI/OhoxoIXzh2SsQpsR3e9OhXPDE3fPdbdXB
5a5wDErnRT0diAQrB5qu5Zbt77/QD039ZSQiKKs0DjRbqnAP6vaS6beDGp70brMY
vKvHSs1uYEC3VNA3YvUzbbohGnU8hP2YRKmQ3djc0J92xsgNT8VXlW7z/ZaplC/r
pYvxFMXkROFweD8HFQ5zqXGBmfCuMYeMCVR7M4Xmqd5z5txXHanUgKu+2WzrNxQF
ByTk6o3KwEUcnIHtk6Vfj/Vpygy1033rk9nv8mTb9oshYG4iVPXH1iISeBhyAcMC
3y6DSzu9/CZ0jOTANTF3OJxaPbQyD89Qnwyb7+U/6iDWYU4Oy4uoKb1FPer19HAt
GH5bzNi1iTGluobfWCi4wHzv1gOWNDQnS2UyZBK7LMtVJAoX937IYoS/yMM9DaUM
osizzucYlULzxw7KaQoeI0xX0ni8JXUb0+LF7DEcvL37yBOEjgNZPtINN8+7vmcO
QbqY8k0E6FOXZzOLuJ5kxLk4zesYsuXpI7yL0S3BGS4jRYdKSxQi5PfZTnjo2Ex2
HQa/BBskbesrQhxDKSkSpytBN0YCHdNzgulahbyrW5/yGzeg6jD2ZqqRtDYKqIqQ
kjmjJ+n0lLtCIF6cGFYMzXv9iUR6ru3q8d2jrF12X1te9Mk0slF2OgkL1DVG82XI
eFJob7Pdxr9mvukZeh6NdY8v1QPOsvuXQA5Bmp3s6tWZoczMDt1Ha8ekXqiXuVhB
3G5hFXbpmYOcAh0wmW88pkEmor4NN1Uu0FRbaxPryy8i8Mnf5T9Kq8iBQQkMcvpK
xVnJOPpJPvgK2fwLQETU15oiYDGGo9TwesL0/nVnC62VaYqrpvXdOCPtZsM/vO0A
6zgLKN/OiQNCaGrxKC+BzKO7Iexdhza85WR+qlXZOKAwDTlvhpIm30H0FQAQlfNW
aEftpUD3FcOsgMUYaJ7Txtw6HOtDHdFDPREt3mn+819eDt+8Am8n9GuxyGbH0Wwl
Vv1IO0WFRupyxFqu8ad5Fnii28ht2K8pmw5z2eL99bQvebAzCj8cI3h9lG6iLRp9
kZfHwro2iZvdrWEz68nG5fwtvW2xmwPYoY31CeRTN8aNX73Bsye63eG8hyU7fRwa
6/N6rUSoDAmKBG7bsRH5sVBVc2dSSuzOFTQ/B/8HwCbDdCLIGnyYW9Tf67KMonq0
nL4T27VZE/TXTVyyteZMNkrjruQ/QEMwUQrRfnNeWF466UxW/7HBJ8wIkiqBWmCq
jgHOO557yOOY4DCLtV6rCRuJBvkfoZ4HeZWqO7VcPk3pMonD88Q3ceKjPDuUb8nI
1xboEGfQfmsD9madkBGO6LJY+ejcBU3Ti2jP4UoyFlUFxeAR0TsNrZ3bqNDvhlus
plNCYtcv4DgjjOFdnhUwLH8oQcGDX+xhHxb45O6IIRCB9LEhvw7Rr+7meBbhNGEx
5wV1aytRvUAUnht7zSqwC2m02IY41VXpbJPmeSlOBzE3/JZdRKG73tMziPA/NU0O
FHDr2WDAjYkfebDXVUy/iEO7ohKB94yWJYlk9qReE6LeYt1KlXlTyLs7dkotR9JO
vqgl7jIox8L4cec9UJP3SAz8ZLTNBmDTMJKfBDlU8bG56xkQtLlNXMdz93/1a7xP
x1rN8jAj1IbxzJwBHBN9XBgtVxA4q2ihivpFDsNxiP3VYLkYb3uBUSB2cZLAXrSD
iIbXWHIjOdxfeP9fdkzeBi9YpD/2AemgcNM8eDPmNGDxsonLKF7rggcCxksVE5MU
nZjqd5rdvSn8sHDEdqg+nWXAGxjScezKTDwZTVOtjtTZqG9q8Fya4AaF/vTr+Ex4
CpyygBBkq7iMCkVOjrGpj/yVr2Dq7ZRJ2PUzktZoiNiCl4sdFK3bJjO8//Y4rFA9
bfrqQET1TpPenrOhgOsHcQoQmGP8/na/C4ur3H4uQvRC/ptmsrvylWaB1VZTCvlD
UuwUr2hlqnnYHrm6UEzj28ZD6fFgFxv4n9hpAD5dC4ES5aTXFjO8TJ/LGWkHpcuP
UlukDzEl5aCH9MS19JWw3m6PcbABdpd7SrXR9ufTA9IpCNvyZ91jhHn7sMrPOsnn
XOw6johQeZ23hzM8/hsPkf/iEB28XHVtnY/x59kjyrYm2LCqFMuXNu4tbshibDMO
KBOm1OzCCsyEY9AoI1uJ9mLgwBW6FPaqAiSXhu/At9iA1xB2+pRV8iJIUhC7iTp0
W7ykF8l6iwmMQ6h1fcJNiiwZGQKaN/QnT/KPAiYTDauBLVBeIhbSnI6GCABBvajM
iGWbLbAj/ji+w7EP3OMUaYVfnwK7L+kFhs+6XsBPhRPUqy1p2pw2ib+w1yPrhF5E
CktnfhHkLgDrGACgv05oJAYf7Y7/zsq6uzyvgyk4r4IIrt2sd616kvOWSFlYtjgY
E45G+h534jbs/kgrPEf2STIhyZIYYWt/Pr6GfauI80R+KfsuLOCj5hfX9q93HslO
t/zz5lJ6pSrX6Ds5EUCy9YsKwYEKf/Xz85qoVI40vf390pdqKSI++Gjp1vn5/BUr
xUNjmfAnVYDknax00ti0CjRNLPiLu9fyE385zCT0c4E5SBfjQi2lXeuyYTscrJoW
7jWbiZhRcSuFcBvJqo7LOdC/KoU2vN0oRHr4svb8Mv+2wDMZ7oo5GCx4o0O4UCvG
lyFKmS5ewpHDzqhvDfA/tYoZU9wMUoxGBIMaiNjyUcwlx2LOu7CiwxeWZRcSDFuB
mWLACSya+P0fz9dCfUx6A+0B7A6y5sm9qDxZ7BN7xAk2oP31OctSvoVUAwZqF3qy
rg/cv0TJIxh53R/XInXsTwgyhAv369v/7kHvGN8G2wWAvSLP3WKadqlynbMel+Ap
h0uKwvcpHIdkhwjLdP5+gzfX4dTgY7bKUNCgu59FC76HCszLurVhsjLT2swPSf6i
uCEKV2HCFiQmiKj7bKJYlpTOEvyRHgWVgPDFYH8Hk4HIFP+2xtte8akpGCR39Vn3
Acm9zsBpwrb3o2CcgEd3VrhfCoqFbGCGjILkF/152X+Vu2QYZ+598tCi5AjOdAGC
f09gaCjPf1f4DSFMyw8IScnJjOAnfPhbpQtcN9DRyz1t8z8cgB94jyKe5EPidXhH
3cPSef1dG33ICxM2eFu0gXZrez2Z7mOhN04AHu3KrM2vbcn7MqsmwGeobGKnR5Fu
teTFRCURNkcKiD2JmeBsIwKyEwbGxkQRWmzuFDP18cNWdawYmcbZ4HLrKCmrSLNI
XeT3+y6+F0w+cm0Bj6BoXa0YReJoEypjNKncbAkl/AFs7rMEabiDc9u0FIM3EOwN
XMofgpInTm3I/JY1+DcvVbcPrh7jXtFFRFOrIRhuc5ptSqo4//8aFq5IxHGF4TpV
RV0Lvga6osOSd2PHWjFotOsC3h7B1BTlq+MZEDRZN+8dwfcLr0ju8WdqNFHs/wn/
tAti4LZni4Cjss1MC/E2fCsxLIRN78HVbqppZKH05fOAGcfDuRkzlzjIpByqc8hW
mPVPPW2zVsHEqBWf/ld0jNMTav2q6QOjHrtEr/gVl7pwtCnsb+MJkH9R5gWx37TM
L7aC9eKS3hkmh5UFhixkx7eJDiJOsQXGguMJDbscobaDfKPDqNfJIfgGZFZQtye4
1frrGxi7XFJEo6G1kvDAjqNjfBl2JHrUkmii+T0FatgXnZTnJdRR5PIJqy+jbTGw
WBxFzo7VszwW1IPUMpuOGX1UytpsOdUlzIxMFg+WK2UlgBWsTnm/NkjVcDrV4N+X
dMuNxjOS03X1EORAKkiXkQTgmDXtcDsToDutT+xp0Iq0w4cyWS8GdIfZhln8DjrK
sJN21qhMpYEnn5vLk6gH18QK87aIFU7e5e8lkcp8mc5D2cp+eOV4hQ24LLWiS5I8
rUTTrl6PaWM6QW3CKPLwMAlMRJ4b8MjNWr2s1odcrF/sO7BIcUnC8FBEmHmtIFZF
3NwXDrK2zDWjDZt7qdM71bQKuVTSkSJ80uagTz32/91NNnQAznwegNJo5QGWXc10
UpKoc9r9JzGIcP/+zKH++cmAkszhS9hVROjBocTnd7VXWr2CFX8iBkOnGVSy/cYy
EBvQJjHKdSlhmjifswlLh0ZMAiMPzwngsg6UIOgUegY4p1DkN/vEXLif6ddAx3lC
Vx9CljYQJM/AuL0BqxKrOwh2rD2DMVyl2Lp5wQvMF1Vq0oAZPgjYEobrRWJz3DJd
Yir5vz9M/Y+aC09SN0CHIbQ3cwVQwX/fnHQ0R3+uciHKbOogOilj9wsVw+Geg4qz
OzyuHShtf9irlG3SbqMcg7gz8jEJ3faYs1PE4q/SVTW0GcrLedoKGpTM+pR/7Zvu
O1qVg0J7oBw8pvzyXHOQBCulobrrlYn+McrIvF0kDqbF64ctTDrftjk6zuExJfvj
52aIO4pBEIxUZNCu87gkqEFF0UX09Lw22MxxXECn3ZfF40HYRRez6hjQ//QPh5Dp
LDGE/UPNRcHK7MyKup9i9auGzcIIpeRAuiGFI6ri7Y4GUaAUImgT+gDPKc7fBiwQ
Fq5TgB0Oop2Gq2KJ2Ee++7iiPkVJzM/bGqk4WL7reXcAbTGPMyqY6W+njaxmYtwI
NwLgHRX6nCEW9bcWN78yB93h6NSQtUlpOamV+cFJwuabwyM8It3TNghSYO7oWPdd
fYT5OEAEaw7N7DPo02g73K3FNEXJnPTnG5MktPeJOduIa9d0yQGtBmYXUee1rdon
Zhth89RrDZUuXb7L0122lVEWO0J2FVNHAKZkC8TgfcuduS+SckVF6rbLYXS0YvWb
ZHMT8AkG8+n9PXpctKX/XuYXzAKVRrovrNb732bKfCT6ISbROKWXf+UJH1Sbxm8N
FQuJpudQbKtOWSTFapxGQUBm40rwIqYNm/s9l+jXHZXaeKY5+0nZfReIFmgezMKb
w5/xIyfu0Bg506kRpN53XtX9DnezhOVd0avuD/RQRoaPbQSy+G13jcX5vN6eWmM+
0gfrRB3LF4PblwJUulLgrSvGGcvPhe7Px7r7QqnVClVkzPrDL8qAWkffGlG4NVkM
evDMnrgTJfZ2XNasOHQK0WvVwKvGtoJXyxQQ7s7C+mlsHCj9rZbFEAUDTk2SiteB
kTl91ID2a3DPYjE3v2ByHw+KnOFk+7dUDD8E7QxKzW2v9Hvi8HQxj/bLWVFQACvH
Fe+pNp+6+NMkw3Wm034ahtvWKoXRrHSAThJ3KUXrFg9FLFiYAzeJ3gdEzdHywM7l
/YpP4H6k23VmoOj5EZBtpIowx6HijU05CPFAYyXM8dujFKcmUvRGDP/bZ9L8p9Aj
7LYmQH126B8mWoB8oP5J4QUIZWopKfNMJiqOa/nKOljNtSkX9K7a2Rv2lynALSLV
OMTQ8AEpTilT2GEgeUEOMV1ct+WLnRXzxdB07zLdDFSqVU0Q0gsUFGFn6SbaqDKc
bN5hQktkjm6Qj3W7TGZNJRrhx7P+vp3K5DcdW6MnjfCUuXN0K2TdC0WXny6DCOZm
GdpEIxcqkVcFJrUfzsuq+aag9JV3KqQXmppC8HG8ilhiVSfxd8Iehed29TAi3yq2
NjaM0Yg+Q6eFfU+EQBTJ3TqseMS0h1aKAIa0e5hQItTG5opX1HWpO+UoGvomb1ol
dDpalWfjnM8CJTLFsJPhgyF4A66xkUjuCBjC7s8KQ8w7AsFUNK0dWALw1oodja+g
uf2sOVB59i+FUMfiqSHnVy0BZrY3Pf8KN/A8ZBUxHZNemsU8uEyw3u43bEaixFRL
wUwEP7A6TSfzuVfaq9Jd9RCtsGi0WjsVBAcQn9OVto4g/CMORh77PPRPB5/C7T1R
BcPzN8p/w+0FYbqr4ff/ZxCbpQ04NiAIItDQV6YNQsYZI0aXAKp0ajlKUbxk3Xvt
jA/AYqRUmTBpSJaAc+Wa+L2pQYjYSS8lKW5D1v2EGcJbHZTZ6ugaFxv2aFQGOBoV
nVRImVVEVDgD5jWbIvIT5v3S3hYk/p4xzZgG3LUM1Dkhwg+NxpptW5jqAg+AaKEU
R6vbKBTLTLIEsfr5IYuE4TgFk9ER9l/pMu6CQ1vigdepUOiu1LKPRsEqN5TBbptx
r9zeQdzJr/V9cR8qElh8fqdT6/M0pD6Yo2lJTl5iObdTWm+U5FomAsUdS1mZSUkk
vGBZ7Fxr9mr1XJXnpA90zLxD0onVCe/jCQb6sssnhmuyk7cXQnLeNsYS8Ne2k7Lb
E4g/9tieLCoGsUjcFP4v4xBrTocfif50ZNcyFJgquW3XjJvFljGmmiVtVgFAI8BH
VD+lxdz0OzhoiQ85uYc3M6oX2vkyHKMjLuqxAntcp5m5GatFIG2Nk7z4sp/sxufy
kPERz9/ED1BPuQTXrp8+X9VU4sIxTKZk2PrhB+R41LgBWzov8/zvh5BG+Q1p/ade
bSZWg/vcn/pXvbvQejsOOjzZIpUCh1ZjjVLHjMQ2QWy8TYy+1Kgv5oEchGbIQZYM
kCSQ7EedQi+IlALFjW8/rWSAWlv5gaYMT9ThJ4jkVEk3Mffj0SHTI7n/WTg+Oa/t
WlAv+3loZOD8ozHwon3lIQOnCuMgm9BqQAszNoaC0D1ey/TnzICDFJXx6wuIGSGo
IeChIQMDojEb43HLReepusFnjFLlmXqHkJSvmZ5rX7nYi5SHQH7/PVWV0YkXWJ5Q
4DChXCQ+nvkpLAeYrRZs1IW0baHJbdflEF64SdacU7vJc+W0cqVC+uxcdSL0dtEc
iXnZ5Q0WobG+eKQHumnzKiJpyOQlHSGl4D4JWnIl4llcyPg0USE15kZLil11nhgc
gsmlaMgEBQngGDV+3mhrLhIsvg3W73Y7BNHEIyS6tEixPMNNepmvkD4qE6l7jCtL
2iUc+fVw7nemlxcxygLUO4FteouiUGpGL+LyS+0HOpApgrDVRDtR6c0tWbtFxLWN
sVt3DeS2ZyAelcjh/zOZv0EfczrOQI6hy1SAV14z+7B9tCnyK83HHqxsV4KZ4jK8
WVum9XA0w6A2Api/Ei0FtQqYYD/9lPRCKhsuYDtZtQHMKAl++prNjRyu2aqzbZ/W
/DlENG0GT2Al9hrcqJgDMB35kK87UPnvOLpN9Z7xy7qz/3syLbJtIOXfbFghsxcU
/yzD+q185uDN1k3BCDzBydxu6AZrIauQoG9aix6/q7slcctsIxTkkAj7okHHFiCb
5sBvPurpBte5v8vQSIldiavkG3b1lILJsX8/7dG0zdwCO5V2pPeGmcEGE3XADI4c
A8Qtxj2ZZ4knp6mFyoA7WksLID1Ci62f4RKY2XKUT5mfmMPaO7Na9/3fl0L+Oc47
Cktfw5RCTnayR89MZqwOSjomux5ABR/p/U9QzCOXQg5W9nZAqbu9hwvSau3TZC+w
cUL4EXv29HITbSlRT0JdMGsSJrTtC3buc5bG3t8kzA7u332IbP9vxDgZt4Ql7lbq
6HOwaYucaLztc4BYnQ3+/2n97jE94vTymCdE8wDZcF0GkZFChk2J2Wk81eEytR3e
UuXz9lee+jUu5+sjJxUrLYBBthZgJQe7u1e2y6pvnzfDJAX+tUUqGjVM/MXT9o0v
52N+FLNftTE2aLL/evBSuOEQ2BuTDnh5vkGkZvawqb6iOYFf0lLEpUp2MZUH8WF9
pCLX0622Jla6V+iNMOHobWrSywTZ56qWeLUvHViFZ7NTSn+0lUbdKgIoZNGnMX+E
5+MFJGatoJpvONpdr5fAyx/37D49iSABdghBQZa2C7dyyQKVN4x47SV1u9ynBGGX
cF676njEeyOn+GwrXYK7SaacpH7IQZz/xSCiFTQecmLF7B5WmWAOBXALEvISlUpS
AoL5KRBE6z+Yr3jVnzRCWKDYXt6Hz9AeQdYJWxdqHVtL66kn0F1Y7wQ2R4eELMmA
dG1fpzv8fXV94CCg8R+uDwKUd+iOxAqw3vUl534k7adSbFqpEyFDoXIBHv1kM00H
orv6JHaw0Vtb785plQUV2TwTilbKg39/RtNraogXGkPqAfTa1xoNzQDFOyaPCjn5
UR3DSFyVX1rz4S4WYs7GBqTwVmsa/b1z/ejpYZyKo2xQBVo6Jw4GatkLMHhN7rCa
Pvub1UeV3g4pzAy6ORw7KczpeGy+rOxYLVkgYEjV7QJZhfB99n0OQrqTTudakAK8
KWP3F0TZxLTUAptqALKRcnM76EKmuSjp216dIShimh+yk2FtrENPWWmwjKek+KeC
tBUaloJkHuyp+cqtb6kLf4OW9fPcmlQuesKDbR3UoI8oG4OUl/1T40Ku40INiory
Qd2nAixZmpWYCk78tmKqwG2i6WFzRhBRbJHUznxgSD+dKo4seAWa+V1tOfQxFOYa
1QwnXD0y5f60kAyKB7xdROG7LurUs6XAVRh885DGf0Bm3B6qBhi02kZqGd9YLQgF
YYHsf1sRntkp6Kysjoj/HYhpGYLUPfYzTfNgf10CMzhbnIdZ5YZaj4trZ1qaGlpW
ZmmwdG5xkRz0oDDbiucjuiGw7d4nC5mfb676iP/owC5FMq6IrFoV8E6M+22ET4a0
VT110EvtBx3wVHPlzTm8yxSIauUJ6jPwrTMGJZMsNQhtTpe/M95vl++Bd9x8Vzrh
DENhC5d4MGAjv3rLQ/b/+DqdIO3o4zlI7nQ/SS7vIGavtkGAa8G41QRFrMrbgD7H
UdRopiFEoN6fPyV1yuDlAtMRIRz0IaLtDZx5cAVh36/hKG+DHLWVmWymLEWoa1jy
nS7OqoImdDAtm171eabV/UMdo1dguoB+0g4iYTpOTTavtMw/TI5h0Z7mwM3cLYmT
vyEs9e7IUbD8VevHGudjbNrXjoI380x6/TI4QZd1DNZo2Pig0lPxn4pnG23sPyZW
q4VonwbVDCC7A3Lpz8F9JyOIP7Rv4ymdDY73xk71BqCjr8ubr9jEojYURs8kqasJ
9KniVK0xo76qaEh4mWioA7a/262/E4pNIJSmVMxHnYgTcT7ZFoq4RsA9fj2txLMS
NJ5BaXigAZsgr3or9H5O5/mpyB1CCDy2oGubF21tAEnPgXDhYZlzQdcZDAsXz45k
UB98iMgCaOVQgdkMzhktdiQJoFdd8/VqQmtkdqLd6L199bi8C5LTU8OcMHd2USOn
WzNAZd1hNsKCV4k3EuR2Hz2RFCMqydxHwRVmja/pQS0kZfR1JQfQq1y0aid5w5Pg
aeNLlxBra+pC8TjgWZzhG1OlmtsWkyV15PCiMoI1hCszJCx7zyGBAL9RRTqrIH1G
CuMTw+nheNaPCo42NKz6Euc5TdKhxv53Jfw5SI9XBN6JbqY9emPjI7+70XhRYJkA
SYvFPUGjun1FpmQhXKylwwieIGs5ACi9eQMvmPGSdrL4W999R2RoAZR0CNTGbr0g
9aNfAAXzDAFQeS37DGkOch0UmgC5s0WCy+jag1YmDcfJeOOoh7BECxXWcoQtmbch
VT0yvpiqjtesfqpEFIQM2kS54vfkrnZ3AWsaC/JgktB/DkslgZoWp5w/UcexK20H
rcDlpYS37WIPxlixGC1ZL8JQxo/fSFCjVtImn7FUYjtZ8UhXNwwLHLMEzqraDoRP
AKrTHqTIoagIZg7umsWaVMRUeyS76wyAAP3OhwYTga+diAxWtEsm4gXoIznhvaor
Um1/kLD5v+MK3/+ubwFDx921CCi1SVba0SLi6E/tF1dbV+gTjN0FWw6QbikwBxrS
fqGdePo8XA6T88BxZnAtqwaHPX7rhhbUZXH+EcWVQXTFoSv2PLQkvyVd4AdSNfLb
ZBTiMeVxOHX/nIMWl2uxn6QsF/HyXstea1+k3/7S5wvWLoWkEeQOALsYRaivPYs9
eK5zuuW0zUfSx/aI6xIxDybElI1YHKEe+YbTlGSKH/VaHE8Q6mafnbKJFKDBllBQ
OgqDngUG9liNdUC8ekKklxDBEpet5N0j9cUWrOjqtxZ3X4SA/BQ54+QjxJTkT9ce
QRDgBkwUNFmFbHgEfaTZlm6KeXpOO3oFkk8zHhFkF69sPNNkUZHU951HYOqMraSR
qU9PXkJ5WR8a4BbIwNhIhHQDPlzDYbuj3X9WdOcZf7/oxt/fBS7t0KMJcf7b8G7V
gcZzCWcrw5xjN3AdV15+7VDQXEyMq612ahWg+9xWoDhA0pOHszPceHvrohY/z/Vo
DSGNc/GwdDpnAmQDRXIqFe6M0x8kA7SASrwrqekxjauEn0T+SXuVZK0tlOUTpms2
+fXiD0G/xfHzXhrHbT5D/yEioNbcspp2KX3z0/WQCHiGLacpUQU5+aIeetAqdL3K
nxgneHaDaVXCLs2yZiWCiFoDUX+la/xvUFwRoyf6SNyD8vZ7GqtRHr+CZFmkI7GV
ygWotGuEfs9Zj/kHqVV59QEv0Wgpu/O7x4LFimONv8kHq+a9RFFFv9HLV0TQe+hh
5Bi/zT74u7XOoqRzpZ9S3cRuDOT5qZIeG7oGoiZca/Pd5pTV2jY1wePZ6Rgc4eqd
+OJhOkRRCMRngO6i3PCfHNkRiBnBs+6H73lZLw10ln2Kcd9dVVTFLWvFAbGfSPiF
lVu4ECxxHOl9hCXc9+crC3aJUCxk1qZG5HGHqhCre/FnsO7twCP+QmSEH8UPoabG
slwayiZpBN0ilf3YSP5VKn/6AHD647cE4Y1OusJx5dZKcUIICndZ08xxBwN9XhNS
cXM9e6uPojZtVnu+ccWgQpURLvKSwOYrbbAylSADF5VJtOwzqQBTZ8q6+khF0aed
1x9qlGIAN+01Hw6OqQGsmMs6S+z3FWeRL2wSJtJ4x0sPE41ZvVfG6UXwvFROPZ3O
lDMnQGnhS8eZ9KtRSVlb97qANewIjvcmKlpQ1nyL4esZIgSqkV4QDOysBGfAWvHj
ksU+f/VaMkPHtsAqg5+ApvEESyh8Lj6v8Um0iVkAs8rTw+bdwSrD63Tm0KwNzu/m
g7OcQu95DtP+wQHvNhS/GjgSpxPWncbqk2qLMn2EVBaeOPw5GCAexyVrTzYVuHDd
P2OmaB729D+KPCyU6GXlt+ZLQwm8mX8Xs1ExojNpvOwnJjKpONduG3m8OIkj+4ZQ
VgMhMj8FpUN0qw5fAGkT3RJTd8iqb9Vp71Jof21fY5XFo5T9kv1h7nMHk/nwYQZ3
aWhX1hB10FM1EiDfckwt6SZuIbSR55xuo2fArHG7wC7h+tiQAH4i9vJ+bKEHTB2P
8BeYLmFFm8qmMKvVsgj+mOPP9mKidq8UJ4YYjYXxSqTpu62H82tKscci4YjnnQet
6p+/osCqLs91MGDe73rDQo7twwVWIbLfqUwLzWwLOehReRMcUhkwyNMSKMXYacdu
S4nVY+0OtS1dI6f793ecLVH1BlOU9nhixhlqeJZBtj5PhTUDmfa6dN7t6cq3YP+B
8J72MU/O6RBkiJKpyZcv/P27k54GsKKsOOlAFRMFzcUPELNS7JnKQ6m+0Y3wTto0
EVG5ETmEA55vZEj55t5HO3DJspg/p7DLE+u1CEiHHt1oWEU7EyxyVkP+a8MpNZVq
rsx/51jzZgAM9xcq22OCgj9r9NId9C4Drtvy9tgvbK1xY+aCVrriNkLzT9aD1GLn
/ATxzN3I9JGJra92bRQiNRVaS92GDEjNVn1Z0RZdDYrj4UgeeQHf6qdq/ipGImte
h5r2NL6B4HggK1f8CwghLodQQpzQuQ8dA6xO5UHg/MbFF/Kuooq9zr9q+WegtrD+
xu423cnK/PYuuo/CXJziN/13LbzrstiC4LznV/w+dm7T52vZRZH/3p0lzkC4Legk
qF9Q0bmeOK1lP1wuqFpM4sUwRXIsxBrvdl+y54TG6lSNgO5m4ILFBCcSwoiqlVVM
Uz+HqAyqmDs/nx+BsJ6VPJXHg4fr1vnWeTN/YfdgoGcpY4vbL5Rwn/Jt3R2XlVrZ
+Ig4VYhSKoupI3kFn0udmIo+ur9rbrgikSwGDAqc/icsfKytZ31UOddTEOxRlbaD
Jkcpd1LnH2uB6DPSZ5fVS+qFYVHqCX2f1H9NPWPUNEAXnAih5Fv77eWGfMcA7U1l
T4flo1UIutV2xSJ+Bbjqf3hSfQ9VLu8lBvTo6h+QedJOzFl9Jrtl4rEF0YJq3TzK
2Wp86grJvsRUi9B1dojb3lC8alQ3CUmTtHw5FdN0E8l/hrUiN6HxGPz2xE/sNN8N
w6uJJf0+KmQZ+LpXr8Sq7odh5h4j6RWx2mP30dWtxjba4BZg2kiXg1x/Bz151Z5k
zhrZBhQF39tsylQ4gzTbn1eV4XhXmlU+nG+CmpIW41Ah+J3GyA5KCwnNXCkCxk/4
IrPn5ZG56gqZ25Oxhi3WdvBYibRxGWBxw6isyks9cx1c5yMZ7J5gbHvKTrzi1T/c
niDegX4ZyKEWr+F2aMmcZ1Nn1q6r83rZJI2tZ/caiERni4PASImfPZJ3PHH92fK9
M+59M6IvIEYs5n3uu46YCJ3s8UDYWMnI+QxBEW5qT58iAUyVVJAy70FUaY5fEHYp
VGpmuGrHiOoXaXmKPfiQWDskfdqT27RTVTuGprS47XaDDWBQ+wluZwQVNZCU6oN7
1jLL2201UBWSFFjwizxj/eSURG4/rCyYwe9RZwDfe+mNnH9oyiPtehvv5tYAsp10
lW9ptvAbIgz1fXaQAKQKMYj9j9gGu3UFfIIXUbRabtnxXfOfMU6WeSJ6ygYrMbQj
qUx72WOOa89BaM8RSDuDhG9AYvAqEsE6K8sgCLYCAKPq6gpnDzDXGJnQEJV1TwBh
2BsFW0ps+OSvZrtNTDjzvwx+WHh/1tI6aUacEsfMTwn12BchBwRGel9YeZM8pwEn
ea0LraPYMUtYCu7Z3pD7daMVQJMcB/0g0w/9y/TiM6wAVlqTOEdrjcwlDdg5mTH0
WJqjpYMBYx8+R5UH0m3gtlWfnEY/e0OpSVlAmPjkrlZl985KyBVZgjqk/KK8dgT9
cOiaHhdRk2gJlApJAExddMPMYvC+BufTot5Mpp95rFXRpGlS3JdgfevCJ7oom+HY
teYGihWhrCGFz/6cfES7TfcBr98l7v1Vg9cPHYD5qxTIG4Jd4bQV7NbXt1fUXDAW
YMf87Q/xVIHREPj6upd/XR/a7pIJMJDZv3Z20fBXRvQd7M1wI6Ihy7JB3p4t3FFY
yJnvAf4gwyQx9T7b3Gtl5sQtkEQ3Qk0Q9JbZsRzftQgPIMwOaH9c4AuZLjrMyjLz
Y+DsPudMtzo0MiqZzzHFTyoI1pv7YMkynwQoGquVd/UwQ9mJQJKAs61UqoOCd9UT
6V6vhrbeAxa0qh+7oTpG3A2TbM3z2j5O5U8VpPjtryFncJl/tEmnwiSs9Ut5oiHz
iydWgsAWwUOUGUamXO9Fv1E9glScJSuJPGGk81naRms0/ZvfXCq9/4fj9GXouoSp
rGBF7KhxK5fcYw9N2rSGmr9bmc6A1gGUDA4c84aNhQHjQI8/PmAiCXaZhiZqoZSR
NIdCT/59n6lkFx0p/J7+hRaQD0ulpZp0BjDMrXRs0ImsfSe4xVFrEefBwQw1qDhG
YYhYInIoPSznEYInotRvxvlZjQeQv6YqR+h1rUNyO1ApMds2LtwsmiwB3VDtvtes
TFbr9TfwgI6NBJEjsCPo9Zyfh8s294s3KNnhs/FzScVI4k3NbBYfN5htbhCu8UN5
0qeeYdQpWVL8Vz+9+OxNY9gvIGCHVtAG1STEEd451NYu30pOPGDRddW3Kkvr12bZ
8aNShEotqdMWBK58iI9jk0JS9DIxov2B2GL4RZQ9GZJAGWKb+kOAESmTXdS5ALyk
MkWQVhwhp1mXLwkauSPEk8brXXxpaj9gws3E4ictaWWLdK16wfXw6CEks3gT19Ei
lQovp/5hXS5cVgQBQ9DOUfnLYD0VVzmY08ERTLv92ql4rb6xFO3da+hkc7H8yjQe
zLnDDxIDCTIOe2Oi9Vn9H3P43fARhPtwy37KULeTs5oNIQwXAR8Y69y8GjQJ6pk7
G/ykWZgDxEILijezWzeQqaO/F0IibDyLoJJxn/jGKSuS2ngJv0v8AtdzKrAPQoYY
9m4jrdnVoopLop0zrI+VvnXieP5dQPtHUvB0aH5J6A4AwlMQF9Z7EZuqvdp9WQKC
rRtO7Jbd1n4vHjKYEZweKCP1V/i4CHkmFS6TgQV2iWRz/+26PzYrogabgD6gQaD+
JneiQgqEhhjXS1zOI7InnLLYvTej8h0pxhzRX+Sc3zCG3oyqV/DdUlTeowmiKOdm
fQI0K7h+Gwdfy+sWacq75LlamE8Nn8i6lZAO+Dd+Mq2wF5/g72MUDWUu4n4Xndit
qA5LplOeVcRkJ7LMrCTe06ciNqSI/knOI8gN3afRKlQe07weHgStbfdwhx+2V9J9
wdL+/gQyS5m/TrJJwH0uCJjFU8LaqNQqGVJFKawMEXzKxETCTn87Bk4z1C2dQarG
BV3gf8/83WIz9DqNJY8sXHaocVq8+G2AUQo8P1a+UcplUKPyqXCkbuQ402n0qI2/
WfjSNG5xKTOrPiStQ47BOLKJPp8RxamBXlZ4CyR/yxjPDmrw1v2zo4xLg930h3qS
F0KsWQthY5w/8L7i8CW9+uiKWV2P0qvUZbuuImH1bymWCyA3YmskkMwHYPSTYqC3
9LIC0jBXkzUO5bzYMG+Xzyo5xjeuo2rFMXe//+R2pvnPN0DuAc/uzjE9EAdcm1Qo
ksdXjhDQOvQ8ErHYc/kvSib8bpAZE+L3sHAeNf5fa1GmbZucxPApInin9mCybZlq
aaa9S3BmxB7AWz2Nrz1KNjufe/unP1s5/xvaTzJEaWPhL2ux1oJ4xBzPeZCDDYeA
z5mTr0GRxXXgKhd5+RyXqibbSp3U8wusDjm7MFsyaS9pbUrwBqp1rWv+z5mj9428
T1Sv3yC10TqDuA1dcIowsUi4QF3UlTzPRp4bumyKTJ5UGhDT0JQy2cgjSpMRQqyr
7+WYErjXykn7q2+FnBZpx4VHR+a2fQ+T/3hxuU2PLZWIhgObFuA9GhXLIZSWN2B5
SqO8c7jdAZP5ai9jLasEJ2RwMoHbh5jLm1yx0geH0uUcneWBX22EJQWIZF6ife7B
CjonDoSuc76t1GojvE9xkcM5ExkMJsrio53JOWvflzHcM28XND54bfPeEwmeZjaZ
Rmbyaw97mOOLKI91/ZaTYF0YXCLsoUaLND8HhR3qGUSKSw280YitT1ExYUAd6L3X
iEhpLBBAq0TRtAvIr8uIBw/yDluMFJMfsO7qvFC2ksmlZKu32lsCLb3SvhSEHlQ9
nKOhuiM8A9EH1m5OCBnMuzUo+fG79HGUhzX3eAuWW/v528V3oo/TAIkTb4LNsxb7
jy+ZfGbjjEokQlTh0irPrKyiKMQ9TRk2W1gnrYk5XQQoV/ygBh2U9aD9LcY//3MS
euIZCFuQZWobuAy7cjNYD4/qKnFAP1QeMXNMOog9uNUfUJiLzOfwneeuq2mdd9kU
vQHsIg26yQ0ejBGEEnaxWhDZDBjlNy9neHexHxh8e5dpSzeG14s96FIBi3D3RP6D
kTA0C6DKziuWdsro4rGPgW5EY77B7wVCpEit8aLLMrUUHHYTkeFl8ML7OOUBUhCp
c1QPlnnbJC6ivBW8Wx8g21c6HtnWl7OM8HOo9GfIFDKq7UT+iZW+nktkEeIXTWzK
RASNet1s321OZi0KbQbhhCn/I3QaGIYp1N9cEj5ebhyyeCDUOxI+/kF84VQLlemE
BEdBVttqNbgxkkZ3QdusMRCXxuZKypCtK1bLxgOcORs3Ld0fzOu8Uus47EaKE/S+
MOAQPcq8Wsi3VnZemf+OCocd/rS6kZ0+vZgB8gKuWdtNZdPLpfgnDYc8Jd6igSbx
JciV41aXTruF4/+Nv5TzMvJDopZ4gBR3+gAqoC4PqjoG1Wt/8PScmlZ24lXvVvTv
NMhgNGvxic42iMzRPNgCXIbngHLFnw/KNYQ7Y2hJF2bE3ojiBVN5bNE787Ytq/fF
IpcztV9N/QTjnjD2bS9vurUi5NbYV+YR0DzlUz1FUomqEs+qqpY5j5Y0YpV30alk
wCrAj1maD8Xz/estW/qtAPbkLvzkE7fGGhW2xiFOeBWDTspd6jRAhkY/yeX8SQcC
n2mnlR/42XZ00YGXlFL7kxtlpdTd3rz4gfNIu/UrXjSMa/4Ow0/t4qj+gxZQUibF
2ESWMzpYF4vLFiCUg23XOwdi+mDQsMELw06bLtsZaCeX4ApdTx2Empu+C+h2Y7SZ
BKgq8N035aaKrAbFDesBlM9HnL3ceUpDVsExFD972Kr6SL2R69Hoko6SyxH3ZczJ
4RlJ+AqsQWdo1cufYrYNxoBLMh7taS3Ls7Yz1VGMw5u7kfqZ/2rQw0nUsX2x65Kn
uqMS1Cq9oJSyw4tn3SE/he/wznxx3nR09+Dokt3JGy94qMRZVnppBvqb4uzoKd9Y
DcXb/nJbXoeXS+k6hVaDpo2DGT9ElccbyzpevCAAMvJERa72l+sONqYevFzmvgts
XlqrIz3GJsnrpdxrI4q3XrVwiilhlhEp+onYVHO5NRtSazQ7yv6c2qCYKsD9P6FP
OaNr1d83z8OqPedBmFeSNPwcQnA9beGe3oNWcCAdZRaq+QcPxbMvAclRjZsGTYbY
SkVJzd9rSC0RGYXbD8MVTsYJKVX/UbOJnwGdzLx0lgIi9SM7ahcI2CqZIlIm+Jc/
92P3Bzd4l7tfN6LiREVrcclAqzleysdIxrzLwGRFdwytacJ3pzFjNDEUaXA0an++
MTmY65AjvAaxTKEoiElNgbvnmQw2t5cNKTPcoEBoEj5JnEVlY7LtSdbhcSeDetLH
bEEJ4IzIiPgaiFYgmWa6eAmx2yXRqZOaZ61GH5g0+O2DblpbvrV/t8G5xOinYZGH
33zow+hMMHJajgf+wlx87dauxWX3kqJ51ynq+GEzPttAyOvQ3nt/SWP1e13wqYW2
95Q5QRoZL4svqu764uNi+mCZrZGQ28vHaNeRGaJUubc4d0WfN3dBZgq5vBFTo4BH
WCRoVKAX8pZePljfvJ6V8lmw4vWWP9Uynw8OnuiCW3bHE3jdqh2O3oFdfgWqVMFd
MXKbwJbDnf0hnL1qgxKfFL9KIWGRwd1rNRL6P75+pE25AGD6d8T5BwzwgXTdlD56
FtjSrhff9aEYvuvoQ0MRIYbE1rnM/qm8T/etUiykIJhilX27Ss/HihgETLE3O37N
KZsNS7qv8DQeQzltnYn7kRo/H83tgKTmyyCKuPKfRR7Ulw9DHnNGqiovazoruWHf
0vC64RF9zE54q6jkNN1iF40ibL/PcpvwbRbJj0HXVvlKC1YnK4/L7K/Eqc/E9PG2
mDq48QtVYD3txrl+27UBNss5Q/Tiu6m+8QVIHbmNY++VbPuMB32D0wuMu3CZnNB8
V+7rDCBJTIinet8WvTOMOpivOeKn+bnAP09yV9NynmHLgKS4e0NzWdf7OKZVLT/2
76CsICufLaaJ3e2uHvAxg4gLjiXSx2GRTWNUAxvKWZINAcsj8oI+IQlxcZ1+Q/sR
s8dkNZvkx2B4ODKyPjt3tXswIc9FA1NVrUmQdSQPMR4Zfoza1zg3J8p6XXZ4tSix
jCKiyKiE2H4yf0qtPBfP5rIa9lLMFF13mpFMtpMvX5zTlHbAbn9kIZ56O7Ee4v0Q
3S8oHmrQGkytsyZv7EshPn0x4xyjmTnWHRhb380BK9yPQCRerNAVWWcyki+3+soN
Iub0U6GWLgTL2VEmYpATEBV2Oa6Xo4p4bz408ZJVavqJcfSTtZ0hJ7GU/jECQSob
qe2WzwxJ57jpziEBVMNVj9grq5tnf7jfBgehjJfwf4G2ALkwjTGXjbZ97eFyxS+J
zSTLP1KiZtmccUI0q/VnaEHiF5kudCr9kldEj6SQhqw9xxGdurb1YioNrU9Qxn46
f8SChubY7Mxzqt+0O+U8imWWv/ZhDStUdYyWQXQtjrjRDHiD00UrykgMvfPefO3r
g9Bb1TwM7ofpDBwWUU6RerqxxqyiNdN4j4YDc2Q0NS15YUNBxDJNN0HpQVi6xUKl
/IKcXNtpMNA9YAF6c3RI/+b0SBsikfQi2bioJJBekfQbjzC/4FVld9wn+db4CxxH
Tl4lYFgODqMgTKYr0hXjvcQtk4L7sV40gp6zutobhcKmAFCCccQJdLV8vJ3hbBvq
1vmsSuR8CF+2zMCLWHMNgy0tugq+kYQ4MgvswLMVbDRK82TjB52yvEtfCOyrWWuO
y3cy34kjmY7tJunAhivOjITnjHdukW7dunkvr4gzF/4TOFkvraTnVCy5S9g4wy17
5omDki8RLoFwKyDKLfLYlkAopVMgDgqMP5b/0PDjqGTwST1HsGniGvMSKE72UeOt
rEe3PJRFsMkCMz/pcmW5uNl/10qOH/TTLA1k6j9Z9GIzTMP0PJtpxezQynfD3KqF
mCT89WXJt34/r7wuhNDt0BQc/OIwTLVQGXK/HejH3xbPSr6eHcNwYQocEqwThtOp
GqZc/p2zcaGpQczIOdxJcR60gbyfzaA23itrsxg8TPMv9tKxXvUYe76LPPXjcJ9v
ue+BX6o/H5Fuc7qiaVnZ07rUTfvEYouMZZBwB4FCZri26LqXTi97pQ+/b4E9RHHE
kDVWsl1riUooXkuQaJ5a4ckuVPcerUirpTTfg00oaEtlloRWiGCoSX9WK+fFAWOS
CPcdRgFzMqaMb/mJEDllk/rPjhHcJmRKz9T55isyDbLdrqCbL73RLeWPLaXrKOYS
L31GHPhNdmuc42jHpX1sSwUzIpYz3B1HL6JB8uBqIpE/fCii/JeKjv9Do/qZr+g4
pcmiv1QRVzHVO9O/td9aILgvJLdmTkF/r7aFtc35FsLfw/UErUceoINn7NwLKpVs
jsjeYlV6+dkS6qS73WGCm2WnT7mKduRpwfxOW0kiQzQ/fDdxHv5uqZMHf99A/NnC
YNCjD2MLfd11Gc6WzsMf/CPjT50j1a2JVAeu4N4r+tO8aKeL6Mj4M4X23aY1S8JX
hlVSSV7GQcu/yW4u/bzASpBTue8AROd5gAuJDeu/FJVFdg7EBNDsR1AfFiFbUeEs
d16nKMWyKmcPl2FdOWgm1yfbsRgaQhmh/BBwVrzdAg7sBGtKpNucE9APHEp/uBbn
LLBb84lDN/53gaUAGmKyey2K6OBFrHRlw2n22qwm/9TaM836R+gRHN8iyMWtwRBl
+shSQkuccAaDmyyVSmd0r0PYCf6ng7w3owwqyhjfs/s6YAH1jLPsa2leA4nKRgZV
54U50nHOM1c3Ai4t92z8+VJ0hTQsc2G7sGIgeCK2y2dap1zeHD6Tk0/BwxcnOmMZ
3HIbXiTX1OEzQsBIOPKv/4BGQPUOl7bBIbDtPyzHzoXWUZ+oBPyfeKzMOVfHYgCz
kzl1xKMh88r5i+mJ4HY37tK1u5tyArqSlAzTjbR1oRhPZl8LYoNGE2y5ZPDlOqpG
sS4XVsOkW0FbPEa7mK5EuJvta7NnO2Xb+JlkZu4uI2zGuYh2w26DNfnIMuLjH9hN
95MEz9JGOWidAlkA13tGbOav14pzbQ8oPfkvNwB1qXExPrIT5djcEQLORmme0hcf
50eJ9aR292Zl969qW4pe+0DL5a8G8VoBMQlPlB34qiuKR2/lpKxyfR6IzoLZ4V9e
5Ih/BNtN0go2bRC7hvwwCgZoik24Td0OsafeWfQglpcD+gdrdsItIaQ4I8CafrOL
2pkQWY+Mc0c9YCrPc3VrL5iTA5670GwBC6HAUOExFCC+vUbxpY8xVuiep3FT3h2a
dMx7crF7vRe/yXLYrI/x9mcXuCt76Da9VUfi0+ocaFg1UNW4BMaHa6graTh1xdDh
V1uzBtizqu40WoHBm+kSB4sJ7EHZGAibIBI0O3pdDT/lsdgcH15Q53QGDtG4rw/T
5oWDo5LT6YtN0LOrys5CTMlPwfpnuq8GbxA9B2vH838y3W72iaNUYNx7KQrJbuIW
0Fr9kik1QWinOI//npBV2V4A9LopSoOWcXQKflNo+MLNDVgIWME1WsN+74nDgsrO
hvdzTy+cSFF2PeRdyco2+fbYTD8HjqvU2SGBA8a86jW58VO0K1pANHMuZt9NuksS
3+YJ6KRa1ED9Cq8fFcY8/B6egCgnFsoqtBQpIiDAinMrfzYt2Ahj9dOZLXYeDbqN
BpSXOaQkM087Ctjt61++sMPSbkhLKucyc4BVMDm6QQFz+Harc17nO8Eb9rbW6kmO
4KHg/CZVsie+yQKYAt4VSrCuBft/BK+/sSggIM365IMo4/WpPkc6pUS73Y4aMfhD
ww+Hiiwem9oqmAyHR0cFOPC7NiGJez5x8tqycJCQCfnKZNjcD5Qs2tcKLq3OxfRf
hWljzhqjI118d13vTGuqWy2G4i51PmPvvDRJ/IGApWCB3HRUl9Y4B3/IURjCRg8C
E9NH9va0HRcnsy8xE1GGu9I//yKTnj3uw6iVBHxq5cOl5cYbvk3my1NBVzOPdBaS
YmjLT5UbxuQAdkE6jLfE1QGm4HMEY4Aqpb5EWIZx0IFc4dntvzTnvGFRA5uDLBVn
0GPXghHXKegxSnfL93Vsu6MA1P2LRKQ/JaB0F9kbm+IaRABwmUEWCvx6Jkd0MtsX
jJ5pQ7pcjwZElJe3IjQL7p3xI3WFH7O4hBDVqBiu+J0TFqTPSqDhjmroU81+ote3
vIMBzoAfO4tRaq4BoonMxkG569Oa+Ghr8F6ibIYH79ZlFwKbpiOY+mBFbZ5+LKIJ
d0ESC/hRA+GSBURz4jvaXV26mdyt0SNdSEm4odUs+GBPomds41EVTl0reyE7IFAq
Typdn+WyOQV0Tu2HPhkrkcsCOXlg6q+8r5RfCPGod0ix/vBzvt25RYrwiP12keql
2Dye1qiX09SXtWy+4QzcpTMbANZasrE919YmnyDVoWtZmCeJbMDd7GJqRFaWF4Xh
ob7SKrndnO8C/uHjVos/Hmq4RIm2IK7mLqDaU0sMRJq1cpfwqxzovbLlDOqFW+J+
I8ZaCBBg7iltADU0U+5kRxAUPzFM8PKpDe62kTCKULSdrJRqAM4huvCWxq82exuR
7CS3Yszwx4BQ8mBPjBwvsqDUf3d1NIEOMmtwa5NqGn7bMi3XxWlyUN1Y2yUcijjq
2phSEz0Bw3HeukmS4VcvFlnYr9abNpKbzjhkgGW9Ej9/9TmGMCiv58g27Z01Owe3
LfBQeltWzOKhtYj+L1HmKgmn8NWeMHNyH6S/HY7oLWaN5OrvV+OgOcpkvU0P3tec
QZw3/AvPRMtZoypVX994wZ0fMWsG+pKr/JEls97xTXjoxkpQmV3Fl9Lq9wqkdrmO
de8Xv4bzR/m6+YKePeyoE9bZ1zDWY4m0fL0DqBJ7wmDq5zBARoP0f/tnN83D6dH0
tB0atyelaBA9dsmrzLhMWQtyUbIHwLO4SVWblEoXV3UAefUrKv0WsPNsLPMsuPxK
UriMIQmvn1qnMpsMnUDLRO+egaqrCzdaDE3QRC9II4yBY/t4ORNmzZVSVHBKMjWC
jDwZom9o61GBvFD8IA54iAyHWhz/VmK1lV6fsjrKvZQ1+qC4cH1ONlape1ZJRDVT
lTpLykgyGOK2JqHVEOpSZZUTjelry4zrUwu9AuUj49peiU3BR5ICYrRf71OVzSol
uBbSVQ0Yv9LCazXLLFY9ECUwCnMvrSSNj60GkUW+uPYmcGXKJbUD7hV//7B8eCsU
jZ64N9oqKV+bcr6qoXmLWLZOcE/MP7fVSwh+XZ/VlklXKsZBcxtnEcQysOoY7tvi
oYUQOIzgEDOGOGdAvOcXjoJSUR9d+rUJzmSVRWoAcB0LIqQ4WaTuHpYRQDqGInBr
1b6h/szvAj+fuaeQHH9MnURM/GhPQtH+1y7funJCf3Jb8jSwFPKo/MDOYu+uDwJQ
QjLMcmCfpeZxuBl6D/blV8OzNzx+P6Xmx54a+xHvomBRiT5CXTqoR6u8EGk9a7F3
5bNmgJpPLS9E+eZ+OaZE+ByylS/GcHgNN+IHZJ1w7QxHJ16aW5v6xUQTgjRHrrgi
9WX7etoJWX5+H7tSh3VHejz9wMpJ51PYw4LMM7KznlsseOwEk/kplhs/FThlFiJj
bQTo2CXFdMOk2TAZB2/MBBseikkZJqyO5BZoyZ+zwGZgYcbCnbaWexUopkIFP8VV
iJAP3AM5SyvliD5Fv7LLRhxXkM2DRF/VZyjER8b2cn5EdsrWVbaFR20T/pLczDe3
LUPCWdljJMBkWe9YjJ3bwDXeSimwacJ+RN1wVjkb60u0UF17jdQA07tVRE5HIxI6
HOcVil185oqg+b1JBWap22SvYRrgrKxBjqBVsJQnfCFhk6ZO6fHQkm+TUzr9Y3cu
Tq4onvOLyLpRiycjRzA1dL9I+Tk2V4uSDdVMrmE2/jyYQzD2jAUASjdXngSbufva
iCT+fUTHn0GxsRaA/5rhri5p+4LrxuqNtgAFs+IdOfDcVSf16LJsO3V+F28xNI8Y
wdHU8u0NxDWWhj3HHur7vnhOiklhjtRgHrOpqDZqxuIz6MCx0oCtDi83r9kctKsL
GoLQNkbhSLx+uUMFZrtrt23BzP6HFP0yDIbU1A8gsfeoZCIaiig8SZdEJRWn9rcV
vDwgk3hm1Ct7MyVh4jXTqNquBrQRpd/wTZJbGIDbm4+ePz2aAxtDQJgrmPalMX6+
33KJQcdD/rN76vLAzY8AaVO8t+kS0T0ZbXHfA9XS7FP/e07E5bWqqIZIbFyZsYep
fEH6OJYo5P2M4HN6yJNIPBeK/czMSLmq00KYNsswUBfTMeSZOcZ1UxdTAw52nBa2
0kjm/JOEOD0yAQHxFhTSCGkzva3RI/VFqJpSUXkFsVCCCn85l4iCTPrf5Jiobslu
IWhK6a+IolKvdW7KUCSn4d8LmH7KCVRmkddGDfU68Z1KzTOAAInvCL7fO0aqSJLN
pbnU82UH6Q/Zm66EAE3xapm77JL43qpAVfVjTMtN6+mXFBu+ZeeSwpYup5AT8e5m
7dzgKMHxXPWViLcduznfcySmjQSWmDeifdph6OFLx1CEVajQRfIt8i2+aWm5OlBX
lEaV55OOhZ5wqNKguXPqvbLk23kDoztdghfTwPm1Kep5d2zsBVRq35wiFy9tC2/W
h+gOlxQoKzQNDZXENm1m9unYJn6Q9MrNF4LHPRM/nHBTxQTm2eRRXNupaiGwymwG
2qathefLqhsibAhYC6+ft5VugCUCE+XMhK3OlHp4hHgeoUGcaZaC0ci3FBTJNsqR
6q1qYTWq8nekCj1KnUe96lMKHpjIgRWDKlMPZ5bXLvWCt4iVc3H9VwyW0aNdRocU
8Y/+5vyWE6aVtRnQi04i8jo1XxXfL+Wa2b8xCp9K5z3AHQQ3cef7/h+KC4bHOei/
MtTTRVSgY8W2FA2Oiww1z/fJDGKbFrXB4Dz22ZMw0Igwh9z7LEwaH0yroJCX3yF5
68RGCU/JQ1MYjpa4f3tXE0VtaCwqz20Oi2RFfodUg8G0f6MqfvR76suSjXBrHkOC
5NymkgExbv2K54X7IwdJB0WGRQM7D7jM7LOHGo7mRSNjTj6VtivZz6W1CDInS1rm
IKun66Wl65L4RuDWsw/S/+SXr/pf1k4lS2kEc4OE+ntehOuXK2qDutDfFIkWjpY8
KT0RzvQnena13NnSapxX4Tv+x1jZaQqDQKrNJ+dwgzP0Q50hmzxdCT8Pk2ejxX/f
HVxIVP7stBRnykwQjnOEF5X+zgzR1Ol2dnNqq1gc8JML3nDXOGGRpON5g7FA/OAm
0pTm7ntsOGNJtVYJR0oArvH7iIxKGIb9cSZMPHdUJq5IuxCREmQB5BcVg1It+x3b
vh5SdSCmoY49OFgOIzrTM0Bb83NrLeJdEUO755UIp3iLk5NAUJsVHUfD3vIeykuv
H0WuERiMyW23Plv1FykFCujU+N3nUbfE1k2tp0rbLy3HVGfSWDVZqcicwiaF4NMo
S3lL1ZrUQ310z4TGM79iGqPWwZs13X4s0qdLGvUP8cpnvTfVhYvr8wAIbM58o0FY
GefhRytr1ApxNN1engZiOUVDhxjqelenpWMXlAfFh4eVy/IRJzdyj0+lC0ZQbUxk
sEDtNoQ9WqeFmPZDE3DO7h3EBq+MiV4YNmcZtT1h9nWZIDnA5JMBdG1yswr+ejbL
UPGUYAJRTtbiAToqJpXkULsCTz8TytSvE4qrh4M5ilTqx7smM4TokUPh/ENkrhGi
F9TwCBieFjNd5rDfaqEu9IBXPrb4UBh01E6z5FW0TfPfRGCZ+uqQjrN5F8dA7bwb
zkK2FYzcb7B5DMQ5cjT8yIck1538zoCMOeoQLqQlykZLhXpm++gQu2mCD3iZGfFS
iV1rigeNHyAXkFyE+X15+bu/6dEdCQQuxNWVbpqHZWkd2UGMuaIYeQ9rMJf3kqwc
b9mjr9lNfR7BhbRVcj5yY+HoZFhL1p7cDz2tqLj3lZrMfsE1A90xYor7ooHrM9Eg
H3+Jmpos+wh9L/1/AgFAP/FaGic0uGl4jmr8DFcXoMqzwtMERNidOPCAFTubPyG9
XQy2054XcYSFDVqBazaP8IeAK7E0lfeb+z6eXTvNRre4XCB1vCPuaAJiPalLxd1Y
B6QyL2nwOpf0RJg2kVWRqNH6g/ogel/46AVpL0Y887ZEq0QS+G3XcbYK0K0W7QFP
+neWxfNjmfb4YwusZX/5pVLj5EVznIdw+HHueXnxOIMckT/ulWWjyvpm0JgdfWJx
Z8qZMdmxFjGhLXbFQ5vP/Cwym9nz+U2leNEA3sZn5X18hTKMNRJZWwnZOX9hia+f
vQ4mYHbsARzasSpcAAoT/LmetYTcSFWvq0e0UbigOoFcxOGs2+F1ocduMNGhpRVL
zDaWNK0DodYZR3dADH0e3Wa1FI79jzLTJC7+7Esewvh4DyycGXTP3ul1zvjzsHWO
8MG0n+CbC3kJ3sHeX/LKhYrkYyIVnO0/J20FHFHd+PZIZbaz2xjAfQBQ6YyVIXsd
a/BxS35iSEjJ1vwJ9kizmgPP7xAd4p8WSLGGsi5xMDWMB1fmyCYkWX+b7P33NOQ0
Xb3+YwKNEuNutzRX+eQovGXKaPUhWoJxRlTivFWTz4ZNcr/kr1V2/zmSJs8UM1N4
am3X7+RxY5f/pNdUZbA06uKpdEm/qjCxEp8s4Cv+PZjN1WXL9ehA5wwXnt/dCXy/
zHS7qwsIXir3PDPNqimlNNjaq0fE3s0izDv//L9WSCQ7t17++8j/5rN/X1DH939V
ANHY49qTJ0cs4edu12TtB59ecBtRHdtaxDFDV5bMDyRyX6PwIs0HQ4esNz6gGNuo
oMzhKmRnNH99tXqaYXhZ+BMJbfNmWh3/pwCgGPoWtU2FBviaKxu+rwUIW5zR/xaM
JhvDXY8jGJvYtlrLcVHw+nATzTZAaJBbI3ZeflICawElIe6rnfkB75HyKUju8AGo
pOXC4AWy17s3up1bs5o1htwgAwWuBT9Sb67PADgbUwc2hX1fpqIOABkchi0wpV0L
d72faAj16caX+LnyyiHb5wsQeOzhEQt8SlB1E8sY4kyGWQM5ACa+2VUKTDniJ+HA
s40vFRrM+iUALIviWbNnsYLyJ7d6ISVmmLh5TQROAXpMC8e3AScbltFvAm2FvRXd
jgvhVwo9Oj8roRGmTpiFRlh5N/RENT5dQlsctzMr1YcesO23alSkFCev8q/3w4e6
0ZdzD5VtFE+qi28NCH6yZA9xkCd7kR/1Zk6sYVNF/u2hm9aWPYN4HUWXUOr5H/Vi
Djn6eE4BGy+TotBE4OZ9Jvlqc+b124M16b1CBf8959msLMPnXKZa17/q6ib+1mKr
SJq6D4zsiLbgkutcjXXWSqK5IfendDP2HgKG12Hf0Jxlqfj7kLHnGc+jNXxMsirD
Xj3NzQXTwnnCSczqyCyyjqDjmb3zecAhRmVS4R8WKqMtgqbgcCkvZAfpAT+y8eM2
nxVFMKdXsnQNSn1j/kGPHuB7U/TxG8j7n0AFmFvAD0cxjPNR2AFAJJpHjHYX/9nD
NBY2QojzEyKIHMUkR5LPaeR+g8ZZLATwj6g8cs3G+yUExfW3udSQjlwKY6xwir2M
a/Y9XANtjLEAUax3ipKeFIuIWKrLPy9rbYsSzjp4kaXPyQYgBj80mk13OTL97GEQ
7dzGS1WkfZ6CsGR5c7AmQ+BomNCGU0EPjKxstP38iqED+1fZ5LimdWn6kZTECa/F
t5dq9FkjgTTevaXKwtG6AfsyTRoySRv2YkeaxidGIRZEUliTpdki/HpJqjsLk8Wk
PB1OXIINM+HJsM3lpTSR+nhkBGTdOaB6FlRhkOoJHijnIpy1TVfmffX7AIrNyxcW
QIOseu91buUbOIEjT1ULQqnReq3oQgpQHgoKqqDSt6T7LCOeXyrtHQB5tH61KK8i
keqW0KHacmzUUDkdlEewPSI8M6NiweY/h205dENZamYiEh3f84TNHC5DrB/+tW5H
u4Tjno/ucgheA1xtxgXxy7dDeqy62alKOR2v+Ujew/iBj5Rd/0TmG6X9SGbCn6Ow
h8PanWCSobPRN1PhuicxpOd/UTfIIMNqiC10Wy5F8gxL8WdhRiGlZdZ4oyXNclX+
lA4UzpDIBqkpcj7pbrH/q33ejpxGsTiMFQpp7GcmfBpRULFlJQhvVWUQnZ13VqHb
TrfEYkmovK0kRY0bwfbGWzXwYOtMsHTh0a8oykI9kmKAscRFqSFkkS1hkGaeA2Eg
Urs1hXawDHqmJjfWoEMJ7z2sRCwX1eRT2Lty17AAxwN3hJVudxwzH/1hmTPo67WG
5kF+VlQtWEiYj8g4pRejYodPpEeow4U7z0Fn0j5Fezk1rE8e+6oB73RGm9nLxa9/
K5N+Coig4rCqwWSCjPxl+cGb45BkyH23sspjSJIfsdldX0LgyeUpStMC865KRv6S
YsZBOfw2D/Fz5ZVWuDzR2rqzLo/KEC9X7xr2UY6RqabvhZSALqwgI45qWojaImFB
60vw+srbgYag/JqLyCiVPZb4jh7dAB/QyBJv8ZhOMOivl9kVwrAbKcBinIYtCXIK
J8H3W6qaj9jUh5qnQvbEViRyRMFuC4XP6JtIXXmXvxKw4VWO073igTMAJCqMmg8E
5K0oPJTOePm9bzX+kXvOXRfQlDAa40wbRMF0eB5FdaiJs7vAq6TWUNvgxGAS+Cpk
/qH4hm2+ucCf/G5dUjwgee9QWyDPBL/MSWOMZG1USqY4o/FLpc20kkHWnJNQm0AD
P5fxQUrMQl2UOK9Uxj1vKyehQnVbtuPsaSBEioGk0aNnTb6mPKtF4OgGBmpDSXJE
yXKLVSE6Umf+46A1+DiMv1r7TnFg4ZWxRLnBhIHrCCRhJHVFaYN56Lt+Vz/xhWMo
tBoAgFFHIKtDM0dD+apQdmc5LePG4Eu1OBWw6ZdYFl/IGePYqqw06qw5ieLPiwKZ
cptekt6ksvR5nFdmDTXyrXdLt1b+oWOhW9rF2QRBAMkwDd3LwnK+8q5OMWxVjBEw
xsih8WYVSYrokZk/2P35gEtAotEcMijUEByvXZcnKz7AZoh2TGgjtT4p4IvzbTkB
ZiUEHByXI87gKPhkdcID6zd0nAx4L8+tVa9zJrMfMRyAIQL6hIe9fGwq6rllgSoT
jYj5opEs0UOkAEUK+3uyVGAff4gjnMUVE9dAizFDOxYyVZO9lyCfVBQVeKNbxinj
a7WBkNMMLt3iPdg9W5uGZEccfZC3qk5/cmF2R4gnGONPlg7c6fr9TZf1C6jLC4ch
cI6jqeWMOTJltLDOtmgccJ4j8rvt3faZgXcKlKlED2yfUcMkJEQ3676bMh8xhtCA
2Rmzj0JUVHq3Zdm0SGbjzQEE+U99XHe2V/+cLn55NMb0q0nP1Pg5hOHAktOthwlq
gksU+Uog0eE7AjZZ40AKu6j2tX0cHXvjlqiJqN12sbRqZiDBreRu6lmexJTtAgwr
NJH0ExOcQqSgGTfYVEqJBeBbaybDMRezAJUp/C2qps83VXETHdM7/U5LRBQCuXwh
abg32oWL/M1dFKx4dwjEDdvEtwFhVGlWiI+icPOwXZASAUjV1fxf49JJ5X3/FR0P
AVOaAo/91LORL9HYgYf1xoROy8Ib+R4hzsO+ikV/dvu0Q0+MusEEjGXvQidsrZlC
U9C4FVYU/BsePVRa7576BqZwiQaWcA4Dj3CZJwC2ZOw=
`pragma protect end_protected
