`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
pqQekuZ9FcAaBCiJnZawXUsRhz+4DecJyQKTmkb9ZjUieSErjHT+76AeGM7wN1hq
/veBU6rp7j9t+eUIkTVoj+okSzMujOgmmS1pE+L9SG0kDPC245QJwqQfTQQyNbxY
QPnsr+15oyk8qgu8CZOcLhL1qViZ0c2W0rOlzXzeF/U=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2992), data_block
WedtQVPTcZPE8yl4P2obqtFpAjJSiws/31w7bIs9Co3tgBpCc+XSqFAFCdtG/lOV
TZKj3+OxBkaJzF0pHHj4xnRq3nAjUBn3GiAGFESsCfVhZhfXduj1UU6Mt71T7JDk
vhTnaoplOXUaD+DRSJkD0WraC3MYPaN9PDOiUFPSLGm9KLucx/J+Y8OwgPPkaYhY
ff4q1FShHZf1yw6VEGQ0uQTQCP0gF2SNZ0Ftrh+05/hKVwUIqNf+qjKJdZlvNNRG
DzhK85tpIeOzoDxgi6Sp5LD39pnrtSVDPUJcidr86DhY/bNSVDrm8csFcaOZgfTn
V/I3/2xaKSJwy7OsAoFCC5EFWGdlnMu7Ead/RZrOdG13iqNVUU4zVKNHR0d/eZKL
bF8XPF92xIHWrdgWHuOYbVnQtNjYVQWP69MgUmdeHHC8G6e1iIas9scV/oCrIjJ/
/enDwaZ5QC+vYqBsLIjdenUHNsoX9gjm41tx1ml+kLEaXMiHuAazt7D/UhwJNxLo
20hTucrHaqaGMAwbakVY/Pv/09j4g3ZcgtX6ZRQdH3iO4b9FiUJJDoFdF+9OxJNO
nkjmseAqdH/lKIryu4tBk4ecKigTi72py00t6s1iZHHAGMLyEMPzrESHioG/4SjV
6jCfHmKN5k3miPF23wKcDy5BxEjX/6zw5UA4h3SqUVhJP4ShESbZCIVEUsU2f2VZ
QPdq+6peRnOE37rkFUDyOtcQK0knxVLEu81J71iaOQR2vmZglwWRh/Mpcns2d9Yv
ejCaItsFcLvBfit1VOmfQpF2SkdT8XL1J0V3SW4xIbKM2KvOvLzpQpoZwLjbSvLe
a6RWbG4gvzZhYKjvHwymmxbetGo4pyyPqKIX7+1N5svQuElECkj0OZEI9yX113ca
EFaeJiRZrAOEAIppS/kl8UwqGLn+nj5k2PfMx40lTbeEGno0ilnjvOIpFblaz/y3
B8/LAg2IGTHvELryvTRHgWD+ZKPz67cx2OQnOsJXezDLH5z7h2Xgfqe4UYkzp7gp
LosP1lHANXNYpcLm1S+nGfNEmT0VDJwLsfabWybVF9pJ31FDYcC/L0yGMUE1PBId
oLdawsSLLXbv4TWWQLiXgFfX7edgTTIpOawX/lc/fkc9ZCSoyasu0EvGJEDqwgUK
HdFR1D3nz++uKwGJRK1t0RlJbHHVV3Un/veZt6zP55vqABwyDpCKFtxi7dC68oFz
GL84i3WTDO6VfAWKUbQmah5SFJNYwU86sXQ0vv1TqqQ4TmrRPN+tzn4VZkqt0WfD
hJuWyWke3opsWXndNy6OnYP6PtEkKF4ikVzrjFOiI5vv1/KhABvgJCBQY87Cm56h
mO2s71wkUzKUjneTyBmc70vYPJDA3zVf9GJYOynNkiEcWkRLmPP0Fn4q+qJBNWPg
lB3Qu1Bn+466lvIHVkVyvCRGLgzqMeqvPPVJesJs9o3ECXj4A/jMoLjrn6TLbqqx
WGbixhiwkFKsRjSw1fbnpKDau0kN+zoC1ITA4m2RbVj2PhFnA0uWK6TkQOjdje9I
ZGO8wLm1v47bQ1h/6MlnHNjSJG2QqoJI0uaxfWyLeca62gqxzlCinyPlF6ej9mpw
0HsLi2ugMlv9ebfudAbPT5tMOeVu5z4URyENuf/J6BZr9zu+TBOYsj34JR7eEq3k
D4nWgtaLTKpvOwza/VtixB5XVvVxhixeMYRCz/Rz49p6hIbLapV9JI+PI6o+S2Dm
ryDwXsdlNG9JCUawszFHl4poUpHFP14O6HDyj7VyLGAYz84D943NeqXheS1jEZNk
Tucjyr1N4284eWCkv+/yBCPhxu0wADxm4Jarsg5Ors73XUhulfdW8WU8LfG/T8iv
2Ua57Xdyb3rDOoD4PP81pcq3iC4LDogISjkpDglt3+Caj4iduOJsDFMD0iexZ6+t
5ZrnsotP5qj3tsZQLGmVfHrWuN1arNWaVW3niwESAooCIujinxqzKbQlrSuD0vuL
MCKAfSmduyKmZf7VpcAp0NSHIdmLgmASAXw/oU5FbADV7nQUiQU+WLIxSz9zRG/b
Le18qb6f5v2jiGOBaCgP4FVRxEoibDNY6tYlfAIiVxzD0MbZe4d+QvSqjRWqIRVd
p+3UrjngIZTMjjVpWml4bOJeghcZqYKDWe9zLNKqFtZpIeFUyazm4jb12XGTztZ/
Jp64YYXALsWjMiMB05v5ww/uuAmhkX1Lm9jXQ2COy7jgVN/PSigl7KSTU81mlGf1
Q/nCuqZoPCIV/7bgIgXfv0lgHX7tOozQ2ODmwMm1fbZojZqC/kKRjnX9oufJDahH
8dP/tMCf1wrKR0LnYgSTeIOWGdallco5sFjacekK+abpyK8+R3XOhkFFCDeOE/NG
lLJtoK/EPIqxlrvNMWJlJI2qtwZ7PFlXba9U6N9mrH/s2kvh1EXaQaVYteIfDVHj
4iSRCi89c62/O5nn7LxYEpmJOWthdpYdjuzkdyJhOkMsE4gP/juRddGXejwIUv1N
m5q3f9TZlPeq5664L/Y/jQriYHyiKSsRewoKvwQjKPaFeWAM1xDvTRWZ7bDUsqIt
fpeMaPwCb+cefyxku4UZdQkfjQfJCVGS9jVC2W6KMMeh62iZ7HexxYTfZ+/FYIyh
+QW3xAi21nL0F1munpJKQcNtYpch/BG4z3hJZB0HyZ13Il8JQSjuOyKBX8shMtkB
KUAr7m1C8Gk9wMfVlAA/eDZxZ89XYzuHpDv6tVQY4Aonis23gPWjdXwjp0df4hOt
M1Fl5L+wABMgW2EdEf/6ZH0rIzuo17F/2+CP8+LUNjJP20oaLzrBbB7qn0XGYP1M
LUHeP/68WEcsTM+ZSrL2V9qvb44nICHALXKS4OM2qdBenP45xttSuRMMz/N2W4lc
PJC7khXgBgFD+f/Hy8n2TQDYE64B+5mtpqS11uCfiDD4EPhjmdHAPuWrOB5H0fgD
sSatyPyvsU3OcVj4yeshqWp8KZN4XDMH1KmCPR5e0V0ekwGqnCfWCy8yNFd9oJ0P
8s55dkaRTx2mAE/gSDj4pQQGWXffvTZgaVcWITSHK2lFxb3i/m0D5ejzrXteOWC2
4d5YnbiqIuhhCCbo0J1SGRwmhAHMtcgBqx3BXWN1yFB2G5G6ZC/FV2rmCzkUCiJF
cey9Eko02gWjBQ+8bXWsz9uzjxcH/G4s8gv1VT4hpq5YttuQO7CyPASnQLuYr0/9
IONCg4jOMsnTT+F3ylsnlZOV3QY5E7ku99ZUtKSRmTvoAyxPS6gPsmJHmTRtE/ae
oi1QYrEid3MvuScuKwxVwWxnMV/5iSwAMtiHZEJEhVaQXtUoJ2+P2JXXSlHWwQ0C
wWDGeFmH5XKO/FcfOUgZ7L/anVONXtIvz/oubdhYMTwfgbCF7ZshkSbCowAhVYa4
mH7ahLvxlpMwz5C6MaE+MEjKe8O+TLV+h+iF3fSx+e8Tb6h991YowNCmcNLRDwAm
oYesgxwfap1a8MTCAnOpZSWq/6SN7PxYjjV1OUi/hZNdxlHmKEWk4H6wyaspcVko
SPm/V7U4azuvc7XKQVm6yqV2JicnWaJaremNOPJMkgJ+VySbSpAMaQQ7lUSU+LT6
1qNvUww/tBbufmKeByGOiI/9NgS6rXvX+eiBY+jlY9jRp71IV6BocaLa/0I+unWI
Rdpd+Eht8fdVmSlYCdszgQCxo07sYPsX+fZo+DgMcgPsfndgAads7gyBS4i6s8j7
1OUJJknI6kNBJchjPcKhu8aDNPMfO6lgcVO0XGhRwQNPDu4W/JopIeane/68vrw2
8tjifmJtqIorwE+vcURFd9YWi0Po3RIQZH+mkjl8HauKUYbipWWbgdSOijBrENcr
aKgy4W8nu37C1fFeUEJKu+zZDe3Bh7lq6yFs/WQzrjZyHoZQ4KBRC4QsTyn0mC9B
n/SlgWAS2/ie8xwTK5ACOPhNM+nqVqt0bxs5Nv0NLM813pkI+Da6OIZZaW+JDe+6
WMJ2kMOlG9iLtyfY5ICx0w==
`pragma protect end_protected
