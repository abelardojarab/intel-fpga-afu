// caui4_xcvr_644.v

// Generated using ACDS version 18.0.1 261

`timescale 1 ps / 1 ps
module caui4_xcvr_644 #(
		parameter rcfg_enable                                                                     = 1,
		parameter rcfg_jtag_enable                                                                = 1,
		parameter rcfg_separate_avmm_busy                                                         = 0,
		parameter dbg_embedded_debug_enable                                                       = 1,
		parameter dbg_capability_reg_enable                                                       = 1,
		parameter dbg_user_identifier                                                             = 0,
		parameter dbg_stat_soft_logic_enable                                                      = 1,
		parameter dbg_ctrl_soft_logic_enable                                                      = 1,
		parameter rcfg_emb_strm_enable                                                            = 0,
		parameter rcfg_profile_cnt                                                                = 2,
		parameter device_revision                                                                 = "14nm5cr2",
		parameter silicon_revision                                                                = "14nm5cr2",
		parameter reduced_reset_sim_time                                                          = 0,
		parameter duplex_mode                                                                     = "duplex",
		parameter channels                                                                        = 4,
		parameter enable_calibration                                                              = 1,
		parameter enable_direct_reset_control                                                     = 0,
		parameter disable_reset_sequencer                                                         = 0,
		parameter disable_digital_reset_sequencer                                                 = 0,
		parameter l_release_aib_reset_first                                                       = 1,
		parameter bonded_mode                                                                     = "not_bonded",
		parameter pcs_bonding_master                                                              = 0,
		parameter pcs_reset_sequencing_mode                                                       = "bonded",
		parameter enable_manual_bonding_settings                                                  = 0,
		parameter manual_pcs_bonding_mode                                                         = "individual",
		parameter manual_pcs_bonding_comp_cnt                                                     = 0,
		parameter manual_tx_hssi_aib_bonding_mode                                                 = "individual",
		parameter manual_tx_hssi_aib_bonding_comp_cnt                                             = 0,
		parameter manual_tx_core_aib_bonding_mode                                                 = "individual",
		parameter manual_tx_core_aib_bonding_comp_cnt                                             = 0,
		parameter manual_rx_hssi_aib_bonding_mode                                                 = "individual",
		parameter manual_rx_hssi_aib_bonding_comp_cnt                                             = 0,
		parameter manual_rx_core_aib_bonding_mode                                                 = "individual",
		parameter manual_rx_core_aib_bonding_comp_cnt                                             = 0,
		parameter plls                                                                            = 1,
		parameter number_physical_bonding_clocks                                                  = 1,
		parameter cdr_refclk_cnt                                                                  = 1,
		parameter enable_hip                                                                      = 0,
		parameter hip_cal_en                                                                      = "disable",
		parameter enable_ehip                                                                     = 0,
		parameter enable_tx_fast_pipeln_reg                                                       = 0,
		parameter enable_rx_fast_pipeln_reg                                                       = 0,
		parameter tx_coreclkin_clock_network                                                      = "dedicated",
		parameter tx_pcs_bonding_clock_network                                                    = "dedicated",
		parameter rx_coreclkin_clock_network                                                      = "dedicated",
		parameter osc_clk_divider                                                                 = 1,
		parameter enable_tx_x2_coreclkin_port                                                     = 0,
		parameter rcfg_shared                                                                     = 1,
		parameter adme_prot_mode                                                                  = "basic_enh",
		parameter adme_pma_mode                                                                   = "basic",
		parameter adme_tx_power_mode                                                              = "high_perf",
		parameter adme_data_rate                                                                  = "25781250000",
		parameter dbg_prbs_soft_logic_enable                                                      = 1,
		parameter dbg_odi_soft_logic_enable                                                       = 0,
		parameter enable_rcfg_tx_digitalreset_release_ctrl                                        = 0,
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_advanced_user_mode_rx                       = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode                       = "tx_rx_pair_enabled",
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_channel_operation_mode                      = "tx_rx_pair_enabled",
		parameter hssi_rx_pld_pcs_interface_hd_pcs8g_channel_operation_mode                       = "tx_rx_pair_enabled",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_channel_operation_mode                 = "tx_rx_pair_enabled",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_channel_operation_mode          = "tx_rx_pair_enabled",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_channel_operation_mode  = "tx_rx_pair_enabled",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_clklow_clk_hz                          = 322265625,
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_ctrl_plane_bonding_rx                  = "individual_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_fifo_mode_rx                                = "reg_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs8g_fifo_mode_rx                                 = "reg_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_fref_clk_hz                            = 322265625,
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_frequency_rules_en                     = "enable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_func_mode                              = "enable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_hclk_clk_hz                            = 0,
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_hip_en                                 = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs8g_hip_mode                                     = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_hrdrstctl_en                           = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_hrdrstctl_en                    = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx                            = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_low_latency_en_rx                           = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_low_latency_en_rx                      = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en                                      = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_lpbk_en                                     = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs8g_lpbk_en                                      = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_lpbk_en                                = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_lpbk_en                         = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_operating_voltage                      = "standard",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_ac_pwr_rules_en                    = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_pair_ac_pwr_uw_per_mhz             = 0,
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_rx_ac_pwr_uw_per_mhz               = 0,
		parameter hssi_rx_pld_pcs_interface_pcs_rx_block_sel                                      = "teng",
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel                                    = "teng_clk_out",
		parameter hssi_rx_pld_pcs_interface_pcs_rx_clk_sel                                        = "pcs_rx_clk",
		parameter hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en                                     = "hip_rx_disable",
		parameter hssi_rx_pld_pcs_interface_pcs_rx_output_sel                                     = "teng_output",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_rx_pwr_scaling_clk                 = "pma_rx_clk",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_8g_refclk_dig_nonatpg_mode_clk_hz  = 0,
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_fifo_mode_rx                       = "reg_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_pcs_refclk_dig_nonatpg_mode_clk_hz = 0,
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_rx_clk_hz                          = 0,
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_pma_dw_rx                                   = "pma_64b_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs8g_pma_dw_rx                                    = "pma_10b_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_dw_rx                              = "pma_64b_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_pma_dw_rx                       = "pma_64b_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_rx_clk_hz                          = 402832031,
		parameter hssi_rx_pld_pcs_interface_hd_g3pcs_prot_mode                                    = "disabled_prot_mode",
		parameter hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx                                 = "disabled_prot_mode_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_prot_mode_rx                                = "basic_mode_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs8g_prot_mode_rx                                 = "disabled_prot_mode_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_prot_mode_rx                           = "basic_10gpcs_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_prot_mode_rx                    = "teng_reg_mode_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_prot_mode_rx                    = "teng_basic_mode_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_prot_mode_rx            = "teng_mode_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_shared_fifo_width_rx                        = "single_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_shared_fifo_width_rx                   = "single_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_shared_fifo_width_rx    = "single_rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_sim_mode                        = "disable",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_speed_grade                            = "e2",
		parameter hssi_rx_pld_pcs_interface_hd_g3pcs_sup_mode                                     = "user_mode",
		parameter hssi_rx_pld_pcs_interface_hd_krfec_sup_mode                                     = "user_mode",
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_sup_mode                                    = "user_mode",
		parameter hssi_rx_pld_pcs_interface_hd_pcs8g_sup_mode                                     = "user_mode",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_sup_mode                               = "user_mode",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_sup_mode                        = "user_mode",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_sup_mode                        = "user_mode",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_sup_mode                = "user_mode",
		parameter hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode                                = "tx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs10g_test_bus_mode                               = "rx",
		parameter hssi_rx_pld_pcs_interface_hd_pcs_channel_transparent_pcs_rx                     = "disable",
		parameter hssi_rx_pld_pcs_interface_silicon_rev                                           = "14nm5cr2",
		parameter hssi_tx_pld_pcs_interface_hd_pcs10g_advanced_user_mode_tx                       = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode                       = "tx_rx_pair_enabled",
		parameter hssi_tx_pld_pcs_interface_hd_pcs10g_channel_operation_mode                      = "tx_rx_pair_enabled",
		parameter hssi_tx_pld_pcs_interface_hd_pcs8g_channel_operation_mode                       = "tx_rx_pair_enabled",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_channel_operation_mode                 = "tx_rx_pair_enabled",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_channel_operation_mode          = "tx_rx_pair_enabled",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_channel_operation_mode  = "tx_rx_pair_enabled",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_ctrl_plane_bonding              = "individual",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_ctrl_plane_bonding_tx                  = "individual_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs10g_fifo_mode_tx                                = "reg_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs8g_fifo_mode_tx                                 = "reg_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_frequency_rules_en                     = "enable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_func_mode                              = "enable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_hclk_clk_hz                            = 0,
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_hip_en                                 = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs8g_hip_mode                                     = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_hrdrstctl_en                           = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_hrdrstctl_en                    = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx                            = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs10g_low_latency_en_tx                           = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_low_latency_en_tx                      = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en                                      = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs10g_lpbk_en                                     = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs8g_lpbk_en                                      = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_lpbk_en                                = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_lpbk_en                         = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pcs_tx_ac_pwr_uw_per_mhz               = 0,
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel                                    = "teng_clk_out",
		parameter hssi_tx_pld_pcs_interface_pcs_tx_clk_source                                     = "teng",
		parameter hssi_tx_pld_pcs_interface_pcs_tx_data_source                                    = "hip_disable",
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en                                  = "delay1_clk_disable",
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel                                 = "pcs_tx_clk",
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl                                    = "delay1_path0",
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel                                = "one_ff_delay",
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en                                  = "delay2_clk_disable",
		parameter hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl                                    = "delay2_path0",
		parameter hssi_tx_pld_pcs_interface_pcs_tx_output_sel                                     = "teng_output",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pcs_tx_pwr_scaling_clk                 = "pma_tx_clk",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_8g_refclk_dig_nonatpg_mode_clk_hz  = 0,
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_fifo_mode_tx                       = "reg_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_pcs_refclk_dig_nonatpg_mode_clk_hz = 0,
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_tx_clk_hz                          = 0,
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_uhsif_tx_clk_hz                    = 0,
		parameter hssi_tx_pld_pcs_interface_hd_pcs10g_pma_dw_tx                                   = "pma_64b_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs8g_pma_dw_tx                                    = "pma_10b_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_dw_tx                              = "pma_64b_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_pma_dw_tx                       = "pma_64b_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_tx_clk_hz                          = 402832031,
		parameter hssi_tx_pld_pcs_interface_hd_g3pcs_prot_mode                                    = "disabled_prot_mode",
		parameter hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx                                 = "disabled_prot_mode_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs10g_prot_mode_tx                                = "basic_mode_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs8g_prot_mode_tx                                 = "disabled_prot_mode_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_prot_mode_tx                           = "basic_10gpcs_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_prot_mode_tx                    = "teng_reg_mode_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_prot_mode_tx                    = "teng_basic_mode_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_prot_mode_tx            = "teng_mode_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs10g_shared_fifo_width_tx                        = "single_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_shared_fifo_width_tx                   = "single_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_shared_fifo_width_tx    = "single_tx",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_sim_mode                        = "disable",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_speed_grade                            = "e2",
		parameter hssi_tx_pld_pcs_interface_hd_g3pcs_sup_mode                                     = "user_mode",
		parameter hssi_tx_pld_pcs_interface_hd_krfec_sup_mode                                     = "user_mode",
		parameter hssi_tx_pld_pcs_interface_hd_pcs10g_sup_mode                                    = "user_mode",
		parameter hssi_tx_pld_pcs_interface_hd_pcs8g_sup_mode                                     = "user_mode",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_sup_mode                               = "user_mode",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_sup_mode                        = "user_mode",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_sup_mode                        = "user_mode",
		parameter hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_sup_mode                = "user_mode",
		parameter hssi_tx_pld_pcs_interface_silicon_rev                                           = "14nm5cr2",
		parameter hssi_10g_tx_pcs_advanced_user_mode                                              = "disable",
		parameter hssi_10g_tx_pcs_bitslip_en                                                      = "bitslip_dis",
		parameter hssi_10g_tx_pcs_bonding_dft_en                                                  = "dft_dis",
		parameter hssi_10g_tx_pcs_bonding_dft_val                                                 = "dft_0",
		parameter hssi_10g_tx_pcs_crcgen_bypass                                                   = "crcgen_bypass_en",
		parameter hssi_10g_tx_pcs_crcgen_clken                                                    = "crcgen_clk_dis",
		parameter hssi_10g_tx_pcs_crcgen_err                                                      = "crcgen_err_dis",
		parameter hssi_10g_tx_pcs_crcgen_inv                                                      = "crcgen_inv_en",
		parameter hssi_10g_tx_pcs_ctrl_bit_reverse                                                = "ctrl_bit_reverse_dis",
		parameter hssi_10g_tx_pcs_data_bit_reverse                                                = "data_bit_reverse_dis",
		parameter hssi_10g_tx_pcs_dft_clk_out_sel                                                 = "tx_master_clk",
		parameter hssi_10g_tx_pcs_dispgen_bypass                                                  = "dispgen_bypass_en",
		parameter hssi_10g_tx_pcs_dispgen_clken                                                   = "dispgen_clk_dis",
		parameter hssi_10g_tx_pcs_dispgen_err                                                     = "dispgen_err_dis",
		parameter hssi_10g_tx_pcs_dispgen_pipeln                                                  = "dispgen_pipeln_dis",
		parameter hssi_10g_tx_pcs_distdwn_bypass_pipeln                                           = "distdwn_bypass_pipeln_dis",
		parameter hssi_10g_tx_pcs_distup_bypass_pipeln                                            = "distup_bypass_pipeln_dis",
		parameter hssi_10g_tx_pcs_dv_bond                                                         = "dv_bond_dis",
		parameter hssi_10g_tx_pcs_empty_flag_type                                                 = "empty_rd_side",
		parameter hssi_10g_tx_pcs_enc64b66b_txsm_clken                                            = "enc64b66b_txsm_clk_dis",
		parameter hssi_10g_tx_pcs_enc_64b66b_txsm_bypass                                          = "enc_64b66b_txsm_bypass_en",
		parameter hssi_10g_tx_pcs_fastpath                                                        = "fastpath_en",
		parameter hssi_10g_tx_pcs_fec_clken                                                       = "fec_clk_dis",
		parameter hssi_10g_tx_pcs_fec_enable                                                      = "fec_dis",
		parameter hssi_10g_tx_pcs_fifo_double_write                                               = "fifo_double_write_dis",
		parameter hssi_10g_tx_pcs_fifo_reg_fast                                                   = "fifo_reg_fast_dis",
		parameter hssi_10g_tx_pcs_fifo_stop_rd                                                    = "n_rd_empty",
		parameter hssi_10g_tx_pcs_fifo_stop_wr                                                    = "n_wr_full",
		parameter hssi_10g_tx_pcs_frmgen_burst                                                    = "frmgen_burst_dis",
		parameter hssi_10g_tx_pcs_frmgen_bypass                                                   = "frmgen_bypass_en",
		parameter hssi_10g_tx_pcs_frmgen_clken                                                    = "frmgen_clk_dis",
		parameter hssi_10g_tx_pcs_frmgen_mfrm_length                                              = 2048,
		parameter hssi_10g_tx_pcs_frmgen_pipeln                                                   = "frmgen_pipeln_en",
		parameter hssi_10g_tx_pcs_frmgen_pyld_ins                                                 = "frmgen_pyld_ins_dis",
		parameter hssi_10g_tx_pcs_frmgen_wordslip                                                 = "frmgen_wordslip_dis",
		parameter hssi_10g_tx_pcs_full_flag_type                                                  = "full_wr_side",
		parameter hssi_10g_tx_pcs_gb_pipeln_bypass                                                = "disable",
		parameter hssi_10g_tx_pcs_gb_tx_idwidth                                                   = "idwidth_66",
		parameter hssi_10g_tx_pcs_gb_tx_odwidth                                                   = "odwidth_64",
		parameter hssi_10g_tx_pcs_gbred_clken                                                     = "gbred_clk_en",
		parameter hssi_10g_tx_pcs_indv                                                            = "indv_en",
		parameter hssi_10g_tx_pcs_low_latency_en                                                  = "disable",
		parameter hssi_10g_tx_pcs_master_clk_sel                                                  = "master_tx_pma_clk",
		parameter hssi_10g_tx_pcs_pempty_flag_type                                                = "pempty_rd_side",
		parameter hssi_10g_tx_pcs_pfull_flag_type                                                 = "pfull_wr_side",
		parameter hssi_10g_tx_pcs_phcomp_rd_del                                                   = "phcomp_rd_del2",
		parameter hssi_10g_tx_pcs_pld_if_type                                                     = "reg",
		parameter hssi_10g_tx_pcs_prot_mode                                                       = "basic_mode",
		parameter hssi_10g_tx_pcs_pseudo_random                                                   = "all_0",
		parameter hssi_10g_tx_pcs_pseudo_seed_a                                                   = "288230376151711743",
		parameter hssi_10g_tx_pcs_pseudo_seed_b                                                   = "288230376151711743",
		parameter hssi_10g_tx_pcs_random_disp                                                     = "disable",
		parameter hssi_10g_tx_pcs_rdfifo_clken                                                    = "rdfifo_clk_en",
		parameter hssi_10g_tx_pcs_scrm_bypass                                                     = "scrm_bypass_en",
		parameter hssi_10g_tx_pcs_scrm_clken                                                      = "scrm_clk_dis",
		parameter hssi_10g_tx_pcs_scrm_mode                                                       = "async",
		parameter hssi_10g_tx_pcs_scrm_pipeln                                                     = "enable",
		parameter hssi_10g_tx_pcs_sh_err                                                          = "sh_err_dis",
		parameter hssi_10g_tx_pcs_sop_mark                                                        = "sop_mark_dis",
		parameter hssi_10g_tx_pcs_stretch_num_stages                                              = "one_stage",
		parameter hssi_10g_tx_pcs_sup_mode                                                        = "user_mode",
		parameter hssi_10g_tx_pcs_test_mode                                                       = "test_off",
		parameter hssi_10g_tx_pcs_tx_scrm_err                                                     = "scrm_err_dis",
		parameter hssi_10g_tx_pcs_tx_scrm_width                                                   = "bit64",
		parameter hssi_10g_tx_pcs_tx_sh_location                                                  = "msb",
		parameter hssi_10g_tx_pcs_tx_sm_bypass                                                    = "tx_sm_bypass_en",
		parameter hssi_10g_tx_pcs_tx_sm_pipeln                                                    = "tx_sm_pipeln_en",
		parameter hssi_10g_tx_pcs_tx_testbus_sel                                                  = "tx_fifo_testbus1",
		parameter hssi_10g_tx_pcs_txfifo_empty                                                    = "empty_default",
		parameter hssi_10g_tx_pcs_txfifo_full                                                     = "full_default",
		parameter hssi_10g_tx_pcs_txfifo_mode                                                     = "register_mode",
		parameter hssi_10g_tx_pcs_txfifo_pempty                                                   = 2,
		parameter hssi_10g_tx_pcs_txfifo_pfull                                                    = 11,
		parameter hssi_10g_tx_pcs_wr_clk_sel                                                      = "wr_tx_pma_clk",
		parameter hssi_10g_tx_pcs_wrfifo_clken                                                    = "wrfifo_clk_en",
		parameter hssi_10g_tx_pcs_silicon_rev                                                     = "14nm5cr2",
		parameter hssi_8g_rx_pcs_auto_error_replacement                                           = "dis_err_replace",
		parameter hssi_8g_rx_pcs_bit_reversal                                                     = "dis_bit_reversal",
		parameter hssi_8g_rx_pcs_bonding_dft_en                                                   = "dft_dis",
		parameter hssi_8g_rx_pcs_bonding_dft_val                                                  = "dft_0",
		parameter hssi_8g_rx_pcs_bypass_pipeline_reg                                              = "dis_bypass_pipeline",
		parameter hssi_8g_rx_pcs_byte_deserializer                                                = "dis_bds",
		parameter hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask                                            = "dis_rxvalid_mask",
		parameter hssi_8g_rx_pcs_clkcmp_pattern_n                                                 = 0,
		parameter hssi_8g_rx_pcs_clkcmp_pattern_p                                                 = 0,
		parameter hssi_8g_rx_pcs_clock_gate_bds_dec_asn                                           = "en_bds_dec_asn_clk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_cdr_eidle                                             = "en_cdr_eidle_clk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk                                           = "en_dw_pc_wrclk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_rd                                              = "en_dw_rm_rdclk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_dw_rm_wr                                              = "en_dw_rm_wrclk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_dw_wa                                                 = "en_dw_wa_clk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_pc_rdclk                                              = "en_pc_rdclk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk                                           = "en_sw_pc_wrclk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_rd                                              = "en_sw_rm_rdclk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_sw_rm_wr                                              = "en_sw_rm_wrclk_gating",
		parameter hssi_8g_rx_pcs_clock_gate_sw_wa                                                 = "en_sw_wa_clk_gating",
		parameter hssi_8g_rx_pcs_clock_observation_in_pld_core                                    = "internal_sw_wa_clk",
		parameter hssi_8g_rx_pcs_eidle_entry_eios                                                 = "dis_eidle_eios",
		parameter hssi_8g_rx_pcs_eidle_entry_iei                                                  = "dis_eidle_iei",
		parameter hssi_8g_rx_pcs_eidle_entry_sd                                                   = "dis_eidle_sd",
		parameter hssi_8g_rx_pcs_eightb_tenb_decoder                                              = "en_8b10b_ibm",
		parameter hssi_8g_rx_pcs_err_flags_sel                                                    = "err_flags_wa",
		parameter hssi_8g_rx_pcs_fixed_pat_det                                                    = "dis_fixed_patdet",
		parameter hssi_8g_rx_pcs_fixed_pat_num                                                    = 0,
		parameter hssi_8g_rx_pcs_force_signal_detect                                              = "en_force_signal_detect",
		parameter hssi_8g_rx_pcs_gen3_clk_en                                                      = "disable_clk",
		parameter hssi_8g_rx_pcs_gen3_rx_clk_sel                                                  = "rcvd_clk",
		parameter hssi_8g_rx_pcs_gen3_tx_clk_sel                                                  = "tx_pma_clk",
		parameter hssi_8g_rx_pcs_hip_mode                                                         = "dis_hip",
		parameter hssi_8g_rx_pcs_ibm_invalid_code                                                 = "dis_ibm_invalid_code",
		parameter hssi_8g_rx_pcs_invalid_code_flag_only                                           = "dis_invalid_code_only",
		parameter hssi_8g_rx_pcs_pad_or_edb_error_replace                                         = "replace_edb",
		parameter hssi_8g_rx_pcs_pcs_bypass                                                       = "dis_pcs_bypass",
		parameter hssi_8g_rx_pcs_phase_comp_rdptr                                                 = "disable_rdptr",
		parameter hssi_8g_rx_pcs_phase_compensation_fifo                                          = "register_fifo",
		parameter hssi_8g_rx_pcs_pipe_if_enable                                                   = "dis_pipe_rx",
		parameter hssi_8g_rx_pcs_pma_dw                                                           = "ten_bit",
		parameter hssi_8g_rx_pcs_polinv_8b10b_dec                                                 = "dis_polinv_8b10b_dec",
		parameter hssi_8g_rx_pcs_prot_mode                                                        = "disabled_prot_mode",
		parameter hssi_8g_rx_pcs_rate_match                                                       = "dis_rm",
		parameter hssi_8g_rx_pcs_rate_match_del_thres                                             = "dis_rm_del_thres",
		parameter hssi_8g_rx_pcs_rate_match_empty_thres                                           = "dis_rm_empty_thres",
		parameter hssi_8g_rx_pcs_rate_match_full_thres                                            = "dis_rm_full_thres",
		parameter hssi_8g_rx_pcs_rate_match_ins_thres                                             = "dis_rm_ins_thres",
		parameter hssi_8g_rx_pcs_rate_match_start_thres                                           = "dis_rm_start_thres",
		parameter hssi_8g_rx_pcs_rx_clk2                                                          = "rcvd_clk_clk2",
		parameter hssi_8g_rx_pcs_rx_clk_free_running                                              = "en_rx_clk_free_run",
		parameter hssi_8g_rx_pcs_rx_pcs_urst                                                      = "en_rx_pcs_urst",
		parameter hssi_8g_rx_pcs_rx_rcvd_clk                                                      = "rcvd_clk_rcvd_clk",
		parameter hssi_8g_rx_pcs_rx_rd_clk                                                        = "rx_clk",
		parameter hssi_8g_rx_pcs_rx_refclk                                                        = "dis_refclk_sel",
		parameter hssi_8g_rx_pcs_rx_wr_clk                                                        = "rx_clk2_div_1_2_4",
		parameter hssi_8g_rx_pcs_sup_mode                                                         = "user_mode",
		parameter hssi_8g_rx_pcs_symbol_swap                                                      = "dis_symbol_swap",
		parameter hssi_8g_rx_pcs_sync_sm_idle_eios                                                = "dis_syncsm_idle",
		parameter hssi_8g_rx_pcs_test_bus_sel                                                     = "tx_testbus",
		parameter hssi_8g_rx_pcs_tx_rx_parallel_loopback                                          = "dis_plpbk",
		parameter hssi_8g_rx_pcs_wa_boundary_lock_ctrl                                            = "sync_sm",
		parameter hssi_8g_rx_pcs_wa_clk_slip_spacing                                              = 16,
		parameter hssi_8g_rx_pcs_wa_det_latency_sync_status_beh                                   = "dont_care_assert_sync",
		parameter hssi_8g_rx_pcs_wa_disp_err_flag                                                 = "en_disp_err_flag",
		parameter hssi_8g_rx_pcs_wa_kchar                                                         = "dis_kchar",
		parameter hssi_8g_rx_pcs_wa_pd                                                            = "wa_pd_10",
		parameter hssi_8g_rx_pcs_wa_pd_data                                                       = "0",
		parameter hssi_8g_rx_pcs_wa_pd_polarity                                                   = "dont_care_both_pol",
		parameter hssi_8g_rx_pcs_wa_pld_controlled                                                = "dis_pld_ctrl",
		parameter hssi_8g_rx_pcs_wa_renumber_data                                                 = 3,
		parameter hssi_8g_rx_pcs_wa_rgnumber_data                                                 = 3,
		parameter hssi_8g_rx_pcs_wa_rknumber_data                                                 = 3,
		parameter hssi_8g_rx_pcs_wa_rosnumber_data                                                = 1,
		parameter hssi_8g_rx_pcs_wa_rvnumber_data                                                 = 0,
		parameter hssi_8g_rx_pcs_wa_sync_sm_ctrl                                                  = "gige_sync_sm",
		parameter hssi_8g_rx_pcs_wait_cnt                                                         = 0,
		parameter hssi_8g_rx_pcs_silicon_rev                                                      = "14nm5cr2",
		parameter hssi_8g_tx_pcs_bit_reversal                                                     = "dis_bit_reversal",
		parameter hssi_8g_tx_pcs_bonding_dft_en                                                   = "dft_dis",
		parameter hssi_8g_tx_pcs_bonding_dft_val                                                  = "dft_0",
		parameter hssi_8g_tx_pcs_bypass_pipeline_reg                                              = "dis_bypass_pipeline",
		parameter hssi_8g_tx_pcs_byte_serializer                                                  = "dis_bs",
		parameter hssi_8g_tx_pcs_clock_gate_bs_enc                                                = "en_bs_enc_clk_gating",
		parameter hssi_8g_tx_pcs_clock_gate_dw_fifowr                                             = "en_dw_fifowr_clk_gating",
		parameter hssi_8g_tx_pcs_clock_gate_fiford                                                = "en_fiford_clk_gating",
		parameter hssi_8g_tx_pcs_clock_gate_sw_fifowr                                             = "en_sw_fifowr_clk_gating",
		parameter hssi_8g_tx_pcs_clock_observation_in_pld_core                                    = "internal_refclk_b",
		parameter hssi_8g_tx_pcs_data_selection_8b10b_encoder_input                               = "normal_data_path",
		parameter hssi_8g_tx_pcs_dynamic_clk_switch                                               = "dis_dyn_clk_switch",
		parameter hssi_8g_tx_pcs_eightb_tenb_disp_ctrl                                            = "dis_disp_ctrl",
		parameter hssi_8g_tx_pcs_eightb_tenb_encoder                                              = "en_8b10b_ibm",
		parameter hssi_8g_tx_pcs_force_echar                                                      = "dis_force_echar",
		parameter hssi_8g_tx_pcs_force_kchar                                                      = "dis_force_kchar",
		parameter hssi_8g_tx_pcs_gen3_tx_clk_sel                                                  = "dis_tx_clk",
		parameter hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel                                             = "dis_tx_pipe_clk",
		parameter hssi_8g_tx_pcs_hip_mode                                                         = "dis_hip",
		parameter hssi_8g_tx_pcs_pcs_bypass                                                       = "dis_pcs_bypass",
		parameter hssi_8g_tx_pcs_phase_comp_rdptr                                                 = "disable_rdptr",
		parameter hssi_8g_tx_pcs_phase_compensation_fifo                                          = "register_fifo",
		parameter hssi_8g_tx_pcs_phfifo_write_clk_sel                                             = "tx_clk",
		parameter hssi_8g_tx_pcs_pma_dw                                                           = "ten_bit",
		parameter hssi_8g_tx_pcs_prot_mode                                                        = "disabled_prot_mode",
		parameter hssi_8g_tx_pcs_refclk_b_clk_sel                                                 = "tx_pma_clock",
		parameter hssi_8g_tx_pcs_revloop_back_rm                                                  = "dis_rev_loopback_rx_rm",
		parameter hssi_8g_tx_pcs_sup_mode                                                         = "user_mode",
		parameter hssi_8g_tx_pcs_symbol_swap                                                      = "dis_symbol_swap",
		parameter hssi_8g_tx_pcs_tx_bitslip                                                       = "dis_tx_bitslip",
		parameter hssi_8g_tx_pcs_tx_compliance_controlled_disparity                               = "dis_txcompliance",
		parameter hssi_8g_tx_pcs_tx_fast_pld_reg                                                  = "dis_tx_fast_pld_reg",
		parameter hssi_8g_tx_pcs_txclk_freerun                                                    = "en_freerun_tx",
		parameter hssi_8g_tx_pcs_txpcs_urst                                                       = "en_txpcs_urst",
		parameter hssi_8g_tx_pcs_silicon_rev                                                      = "14nm5cr2",
		parameter hssi_avmm1_if_pcs_arbiter_ctrl                                                  = "avmm1_arbiter_uc_sel",
		parameter hssi_avmm1_if_pcs_cal_done                                                      = "avmm1_cal_done_deassert",
		parameter hssi_avmm1_if_pcs_cal_reserved                                                  = 0,
		parameter hssi_avmm1_if_pcs_calibration_feature_en                                        = "avmm1_pcs_calibration_en",
		parameter hssi_avmm1_if_pldadapt_gate_dis                                                 = "disable",
		parameter hssi_avmm1_if_pcs_hip_cal_en                                                    = "disable",
		parameter hssi_avmm1_if_hssiadapt_nfhssi_calibratio_feature_en                            = "disable",
		parameter hssi_avmm1_if_pldadapt_nfhssi_calibratio_feature_en                             = "enable",
		parameter hssi_avmm1_if_hssiadapt_read_blocking_enable                                    = "enable",
		parameter hssi_avmm1_if_pldadapt_read_blocking_enable                                     = "enable",
		parameter hssi_avmm1_if_hssiadapt_uc_blocking_enable                                      = "enable",
		parameter hssi_avmm1_if_pldadapt_uc_blocking_enable                                       = "enable",
		parameter hssi_avmm1_if_hssiadapt_avmm_osc_clock_setting                                  = "osc_clk_div_by1",
		parameter hssi_avmm1_if_pldadapt_avmm_osc_clock_setting                                   = "osc_clk_div_by1",
		parameter hssi_avmm1_if_hssiadapt_avmm_testbus_sel                                        = "avmm1_transfer_testbus",
		parameter hssi_avmm1_if_pldadapt_avmm_testbus_sel                                         = "avmm1_transfer_testbus",
		parameter hssi_avmm1_if_hssiadapt_hip_mode                                                = "disable_hip",
		parameter hssi_avmm1_if_pldadapt_hip_mode                                                 = "disable_hip",
		parameter hssi_avmm1_if_silicon_rev                                                       = "14nm5cr2",
		parameter hssi_avmm1_if_calibration_type                                                  = "one_time",
		parameter pma_cgb_bitslip_enable                                                          = "disable_bitslip",
		parameter pma_cgb_bti_protected                                                           = "false",
		parameter pma_cgb_cgb_bti_en                                                              = "cgb_bti_disable",
		parameter pma_cgb_cgb_power_down                                                          = "normal_cgb",
		parameter pma_cgb_datarate_bps                                                            = "25781250000",
		parameter pma_cgb_initial_settings                                                        = "true",
		parameter pma_cgb_observe_cgb_clocks                                                      = "observe_nothing",
		parameter pma_cgb_pcie_gen                                                                = "non_pcie",
		parameter pma_cgb_pcie_gen3_bitwidth                                                      = "pciegen3_wide",
		parameter pma_cgb_power_rail_er                                                           = 1120,
		parameter pma_cgb_prot_mode                                                               = "basic_tx",
		parameter pma_cgb_ser_mode                                                                = "sixty_four_bit",
		parameter pma_cgb_ser_powerdown                                                           = "normal_poweron_ser",
		parameter pma_cgb_sup_mode                                                                = "user_mode",
		parameter pma_cgb_tx_ucontrol_en                                                          = "disable",
		parameter pma_cgb_tx_ucontrol_pcie                                                        = "gen1",
		parameter pma_cgb_tx_ucontrol_reset                                                       = "disable",
		parameter pma_cgb_uc_cgb_vreg_boost                                                       = "no_voltage_boost",
		parameter pma_cgb_uc_vcc_setting                                                          = "vcc_setting2",
		parameter pma_cgb_vccdreg_output                                                          = "vccdreg_nominal",
		parameter pma_cgb_vreg_sel_ref                                                            = "sel_vccer_4ref",
		parameter pma_cgb_x1_div_m_sel                                                            = "divbypass",
		parameter pma_cgb_silicon_rev                                                             = "14nm5cr2",
		parameter pma_cgb_input_select_x1                                                         = "fpll_bot",
		parameter pma_cgb_input_select_gen3                                                       = "not_used",
		parameter pma_cgb_input_select_xn                                                         = "not_used",
		parameter pma_tx_buf_pm_cr2_tx_path_analog_mode                                           = "user_custom",
		parameter pma_tx_buf_bti_protected                                                        = "false",
		parameter pma_tx_buf_calibration_en                                                       = "false",
		parameter pma_tx_buf_pm_cr2_tx_path_calibration_en                                        = "false",
		parameter pma_tx_buf_calibration_resistor_value                                           = "res_setting0",
		parameter pma_tx_buf_cdr_cp_calibration_en                                                = "cdr_cp_cal_disable",
		parameter pma_tx_buf_chgpmp_current_dn_trim                                               = "cp_current_trimming_dn_setting0",
		parameter pma_tx_buf_chgpmp_current_up_trim                                               = "cp_current_trimming_up_setting0",
		parameter pma_tx_buf_chgpmp_dn_trim_double                                                = "normal_dn_trim_current",
		parameter pma_tx_buf_chgpmp_up_trim_double                                                = "normal_up_trim_current",
		parameter pma_tx_buf_pm_cr2_tx_path_clock_divider_ratio                                   = 1,
		parameter pma_tx_buf_compensation_en                                                      = "enable",
		parameter pma_tx_buf_compensation_posttap_en                                              = "disable",
		parameter pma_tx_buf_cpen_ctrl                                                            = "cp_l1",
		parameter pma_tx_buf_datarate_bps                                                         = "25781250000",
		parameter pma_tx_buf_pm_cr2_tx_path_datarate_bps                                          = "25781250000",
		parameter pma_tx_buf_pm_cr2_tx_path_datawidth                                             = 64,
		parameter pma_tx_buf_dcc_finestep_enin                                                    = "enable",
		parameter pma_tx_buf_dcd_clk_div_ctrl                                                     = "dcd_ck_div128",
		parameter pma_tx_buf_dcd_detection_en                                                     = "disable",
		parameter pma_tx_buf_dft_sel                                                              = "dft_disabled",
		parameter pma_tx_buf_duty_cycle_correction_bandwidth                                      = "dcc_bw_2",
		parameter pma_tx_buf_duty_cycle_correction_bandwidth_dn                                   = "dcd_bw_dn_2",
		parameter pma_tx_buf_duty_cycle_correction_reference1                                     = "dcc_ref1_4",
		parameter pma_tx_buf_duty_cycle_correction_reference2                                     = "dcc_ref2_2",
		parameter pma_tx_buf_duty_cycle_correction_reset_n                                        = "reset",
		parameter pma_tx_buf_duty_cycle_cp_comp_en                                                = "cp_comp_off",
		parameter pma_tx_buf_duty_cycle_detector_cp_cal                                           = "dcd_cp_cal_disable",
		parameter pma_tx_buf_duty_cycle_detector_sa_cal                                           = "dcd_sa_cal_disable",
		parameter pma_tx_buf_duty_cycle_input_polarity                                            = "dcc_input_pos",
		parameter pma_tx_buf_duty_cycle_setting                                                   = "dcc_t32",
		parameter pma_tx_buf_duty_cycle_setting_aux                                               = "dcc2_t32",
		parameter pma_tx_buf_pm_cr2_tx_path_gt_enabled                                            = "enable",
		parameter pma_tx_buf_idle_ctrl                                                            = "id_cpen_off",
		parameter pma_tx_buf_initial_settings                                                     = "true",
		parameter pma_tx_buf_pm_cr2_tx_path_initial_settings                                      = "true",
		parameter pma_tx_buf_jtag_drv_sel                                                         = "drv1",
		parameter pma_tx_buf_jtag_lp                                                              = "lp_off",
		parameter pma_tx_buf_pm_cr2_tx_path_link                                                  = "sr",
		parameter pma_tx_buf_low_power_en                                                         = "disable",
		parameter pma_tx_buf_lst                                                                  = "atb_disabled",
		parameter pma_tx_buf_pm_cr2_tx_rx_mcgb_location_for_pcie                                  = 0,
		parameter pma_tx_buf_optimal                                                              = "true",
		parameter pma_tx_buf_pm_cr2_tx_path_optimal                                               = "true",
		parameter pma_tx_buf_pcie_gen                                                             = "non_pcie",
		parameter pma_tx_buf_pm_cr2_tx_path_pma_tx_divclk_hz                                      = "402832031",
		parameter pma_tx_buf_pm_cr2_tx_path_power_mode                                            = "high_perf",
		parameter pma_tx_buf_pm_cr2_tx_path_power_rail_eht                                        = 1800,
		parameter pma_tx_buf_power_rail_er                                                        = 0,
		parameter pma_tx_buf_pm_cr2_tx_path_power_rail_et                                         = 1120,
		parameter pma_tx_buf_powermode_ac_post_tap                                                = "tx_post_tap_ac_off",
		parameter pma_tx_buf_powermode_ac_pre_tap                                                 = "tx_pre_tap_ac_off",
		parameter pma_tx_buf_powermode_ac_tx_vod_no_jitcomp                                       = "tx_vod_no_jitcomp_ac_l0",
		parameter pma_tx_buf_powermode_ac_tx_vod_w_jitcomp                                        = "tx_vod_w_jitcomp_ac_l31",
		parameter pma_tx_buf_powermode_dc_post_tap                                                = "powerdown_tx_post_tap",
		parameter pma_tx_buf_powermode_dc_pre_tap                                                 = "powerdown_tx_pre_tap",
		parameter pma_tx_buf_powermode_dc_tx_vod_no_jitcomp                                       = "powerdown_tx_vod_no_jitcomp",
		parameter pma_tx_buf_powermode_dc_tx_vod_w_jitcomp                                        = "tx_vod_w_jitcomp_dc_l31",
		parameter pma_tx_buf_pre_emp_sign_1st_post_tap                                            = "fir_post_1t_neg",
		parameter pma_tx_buf_pre_emp_sign_pre_tap_1t                                              = "fir_pre_1t_neg",
		parameter pma_tx_buf_pre_emp_switching_ctrl_1st_post_tap                                  = 0,
		parameter pma_tx_buf_pre_emp_switching_ctrl_pre_tap_1t                                    = 0,
		parameter pma_tx_buf_prot_mode                                                            = "basic_tx",
		parameter pma_tx_buf_pm_cr2_tx_path_prot_mode                                             = "basic_tx",
		parameter pma_tx_buf_res_cal_local                                                        = "non_local",
		parameter pma_tx_buf_rx_det                                                               = "mode_0",
		parameter pma_tx_buf_rx_det_output_sel                                                    = "rx_det_pcie_out",
		parameter pma_tx_buf_rx_det_pdb                                                           = "rx_det_off",
		parameter pma_tx_buf_sense_amp_offset_cal_curr_n                                          = "sa_os_cal_in_0",
		parameter pma_tx_buf_sense_amp_offset_cal_curr_p                                          = 0,
		parameter pma_tx_buf_ser_powerdown                                                        = "normal_ser_on",
		parameter pma_tx_buf_slew_rate_ctrl                                                       = "slew_r5",
		parameter pma_tx_buf_pm_cr2_tx_path_speed_grade                                           = "e2",
		parameter pma_tx_buf_sup_mode                                                             = "user_mode",
		parameter pma_tx_buf_pm_cr2_tx_path_sup_mode                                              = "user_mode",
		parameter pma_tx_buf_swing_level                                                          = "hv",
		parameter pma_tx_buf_pm_cr2_tx_path_swing_level                                           = "hv",
		parameter pma_tx_buf_term_code                                                            = "rterm_code7",
		parameter pma_tx_buf_term_n_tune                                                          = "rterm_n7",
		parameter pma_tx_buf_term_p_tune                                                          = "rterm_p7",
		parameter pma_tx_buf_term_sel                                                             = "r_r2",
		parameter pma_tx_buf_pm_cr2_tx_path_tile_type                                             = "h",
		parameter pma_tx_buf_tri_driver                                                           = "tri_driver_disable",
		parameter pma_tx_buf_pm_cr2_tx_path_tx_pll_clk_hz                                         = "12890625000",
		parameter pma_tx_buf_tx_powerdown                                                         = "normal_tx_on",
		parameter pma_tx_buf_tx_rst_enable                                                        = "enable",
		parameter pma_tx_buf_xtx_path_xcgb_tx_ucontrol_en                                         = "disable",
		parameter pma_tx_buf_uc_gen3                                                              = "gen3_off",
		parameter pma_tx_buf_uc_gen4                                                              = "gen4_off",
		parameter pma_tx_buf_uc_tx_cal                                                            = "uc_tx_cal_on",
		parameter pma_tx_buf_uc_vcc_setting                                                       = "vcc_setting2",
		parameter pma_tx_buf_user_fir_coeff_ctrl_sel                                              = "ram_ctl",
		parameter pma_tx_buf_vod_output_swing_ctrl                                                = 31,
		parameter pma_tx_buf_vreg_output                                                          = "vccdreg_nominal",
		parameter pma_tx_buf_silicon_rev                                                          = "14nm5cr2",
		parameter pma_tx_sequencer_tx_path_rstn_overrideb                                         = "use_sequencer",
		parameter pma_tx_sequencer_xtx_path_xcgb_tx_ucontrol_en                                   = "disable",
		parameter pma_tx_sequencer_xrx_path_uc_cal_clk_bypass                                     = "cal_clk_0",
		parameter pma_tx_sequencer_silicon_rev                                                    = "14nm5cr2",
		parameter hssi_10g_rx_pcs_advanced_user_mode                                              = "disable",
		parameter hssi_10g_rx_pcs_align_del                                                       = "align_del_dis",
		parameter hssi_10g_rx_pcs_ber_bit_err_total_cnt                                           = "bit_err_total_cnt_10g",
		parameter hssi_10g_rx_pcs_ber_clken                                                       = "ber_clk_dis",
		parameter hssi_10g_rx_pcs_ber_xus_timer_window                                            = 19530,
		parameter hssi_10g_rx_pcs_bitslip_mode                                                    = "bitslip_en",
		parameter hssi_10g_rx_pcs_blksync_bitslip_type                                            = "bitslip_comb",
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_cnt                                        = 1,
		parameter hssi_10g_rx_pcs_blksync_bitslip_wait_type                                       = "bitslip_cnt",
		parameter hssi_10g_rx_pcs_blksync_bypass                                                  = "blksync_bypass_en",
		parameter hssi_10g_rx_pcs_blksync_clken                                                   = "blksync_clk_en",
		parameter hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt                                     = "enum_invalid_sh_cnt_10g",
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock                                    = "knum_sh_cnt_postlock_10g",
		parameter hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock                                     = "knum_sh_cnt_prelock_10g",
		parameter hssi_10g_rx_pcs_blksync_pipeln                                                  = "blksync_pipeln_dis",
		parameter hssi_10g_rx_pcs_clr_errblk_cnt_en                                               = "disable",
		parameter hssi_10g_rx_pcs_control_del                                                     = "control_del_none",
		parameter hssi_10g_rx_pcs_crcchk_bypass                                                   = "crcchk_bypass_en",
		parameter hssi_10g_rx_pcs_crcchk_clken                                                    = "crcchk_clk_dis",
		parameter hssi_10g_rx_pcs_crcchk_inv                                                      = "crcchk_inv_en",
		parameter hssi_10g_rx_pcs_crcchk_pipeln                                                   = "crcchk_pipeln_en",
		parameter hssi_10g_rx_pcs_crcflag_pipeln                                                  = "crcflag_pipeln_en",
		parameter hssi_10g_rx_pcs_ctrl_bit_reverse                                                = "ctrl_bit_reverse_dis",
		parameter hssi_10g_rx_pcs_data_bit_reverse                                                = "data_bit_reverse_dis",
		parameter hssi_10g_rx_pcs_dec64b66b_clken                                                 = "dec64b66b_clk_dis",
		parameter hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass                                          = "dec_64b66b_rxsm_bypass_en",
		parameter hssi_10g_rx_pcs_descrm_bypass                                                   = "descrm_bypass_en",
		parameter hssi_10g_rx_pcs_descrm_clken                                                    = "descrm_clk_dis",
		parameter hssi_10g_rx_pcs_descrm_mode                                                     = "async",
		parameter hssi_10g_rx_pcs_descrm_pipeln                                                   = "enable",
		parameter hssi_10g_rx_pcs_dft_clk_out_sel                                                 = "rx_master_clk",
		parameter hssi_10g_rx_pcs_dis_signal_ok                                                   = "dis_signal_ok_dis",
		parameter hssi_10g_rx_pcs_dispchk_bypass                                                  = "dispchk_bypass_en",
		parameter hssi_10g_rx_pcs_empty_flag_type                                                 = "empty_rd_side",
		parameter hssi_10g_rx_pcs_fast_path                                                       = "fast_path_en",
		parameter hssi_10g_rx_pcs_fec_clken                                                       = "fec_clk_dis",
		parameter hssi_10g_rx_pcs_fec_enable                                                      = "fec_dis",
		parameter hssi_10g_rx_pcs_fifo_double_read                                                = "fifo_double_read_dis",
		parameter hssi_10g_rx_pcs_fifo_stop_rd                                                    = "n_rd_empty",
		parameter hssi_10g_rx_pcs_fifo_stop_wr                                                    = "n_wr_full",
		parameter hssi_10g_rx_pcs_force_align                                                     = "force_align_dis",
		parameter hssi_10g_rx_pcs_frmsync_bypass                                                  = "frmsync_bypass_en",
		parameter hssi_10g_rx_pcs_frmsync_clken                                                   = "frmsync_clk_dis",
		parameter hssi_10g_rx_pcs_frmsync_enum_scrm                                               = "enum_scrm_default",
		parameter hssi_10g_rx_pcs_frmsync_enum_sync                                               = "enum_sync_default",
		parameter hssi_10g_rx_pcs_frmsync_flag_type                                               = "location_only",
		parameter hssi_10g_rx_pcs_frmsync_knum_sync                                               = "knum_sync_default",
		parameter hssi_10g_rx_pcs_frmsync_mfrm_length                                             = 2048,
		parameter hssi_10g_rx_pcs_frmsync_pipeln                                                  = "frmsync_pipeln_en",
		parameter hssi_10g_rx_pcs_full_flag_type                                                  = "full_wr_side",
		parameter hssi_10g_rx_pcs_gb_rx_idwidth                                                   = "idwidth_64",
		parameter hssi_10g_rx_pcs_gb_rx_odwidth                                                   = "odwidth_66",
		parameter hssi_10g_rx_pcs_gbexp_clken                                                     = "gbexp_clk_en",
		parameter hssi_10g_rx_pcs_low_latency_en                                                  = "disable",
		parameter hssi_10g_rx_pcs_lpbk_mode                                                       = "lpbk_dis",
		parameter hssi_10g_rx_pcs_master_clk_sel                                                  = "master_rx_pma_clk",
		parameter hssi_10g_rx_pcs_pempty_flag_type                                                = "pempty_rd_side",
		parameter hssi_10g_rx_pcs_pfull_flag_type                                                 = "pfull_wr_side",
		parameter hssi_10g_rx_pcs_phcomp_rd_del                                                   = "phcomp_rd_del2",
		parameter hssi_10g_rx_pcs_pld_if_type                                                     = "reg",
		parameter hssi_10g_rx_pcs_prot_mode                                                       = "basic_mode",
		parameter hssi_10g_rx_pcs_rand_clken                                                      = "rand_clk_dis",
		parameter hssi_10g_rx_pcs_rd_clk_sel                                                      = "rd_rx_pma_clk",
		parameter hssi_10g_rx_pcs_rdfifo_clken                                                    = "rdfifo_clk_en",
		parameter hssi_10g_rx_pcs_rx_fifo_write_ctrl                                              = "blklock_stops",
		parameter hssi_10g_rx_pcs_rx_scrm_width                                                   = "bit64",
		parameter hssi_10g_rx_pcs_rx_sh_location                                                  = "msb",
		parameter hssi_10g_rx_pcs_rx_signal_ok_sel                                                = "synchronized_ver",
		parameter hssi_10g_rx_pcs_rx_sm_bypass                                                    = "rx_sm_bypass_en",
		parameter hssi_10g_rx_pcs_rx_sm_hiber                                                     = "rx_sm_hiber_en",
		parameter hssi_10g_rx_pcs_rx_sm_pipeln                                                    = "rx_sm_pipeln_en",
		parameter hssi_10g_rx_pcs_rx_testbus_sel                                                  = "rx_fifo_testbus1",
		parameter hssi_10g_rx_pcs_rx_true_b2b                                                     = "b2b",
		parameter hssi_10g_rx_pcs_rxfifo_empty                                                    = "empty_default",
		parameter hssi_10g_rx_pcs_rxfifo_full                                                     = "full_default",
		parameter hssi_10g_rx_pcs_rxfifo_mode                                                     = "register_mode",
		parameter hssi_10g_rx_pcs_rxfifo_pempty                                                   = 2,
		parameter hssi_10g_rx_pcs_rxfifo_pfull                                                    = 23,
		parameter hssi_10g_rx_pcs_stretch_num_stages                                              = "one_stage",
		parameter hssi_10g_rx_pcs_sup_mode                                                        = "user_mode",
		parameter hssi_10g_rx_pcs_test_mode                                                       = "test_off",
		parameter hssi_10g_rx_pcs_wrfifo_clken                                                    = "wrfifo_clk_en",
		parameter hssi_10g_rx_pcs_silicon_rev                                                     = "14nm5cr2",
		parameter hssi_pldadapt_rx_aib_clk1_sel                                                   = "aib_clk1_pld_pcs_rx_clk_out",
		parameter hssi_pldadapt_rx_aib_clk2_sel                                                   = "aib_clk2_pld_pma_clkdiv_rx_user",
		parameter hssi_pldadapt_rx_hdpldadapt_aib_fabric_pld_pma_hclk_hz                          = 0,
		parameter hssi_pldadapt_rx_hdpldadapt_aib_fabric_rx_transfer_clk_hz                       = 805664062,
		parameter hssi_pldadapt_rx_asn_bypass_pma_pcie_sw_done                                    = "disable",
		parameter hssi_pldadapt_rx_asn_wait_for_dll_reset_cnt                                     = 64,
		parameter hssi_pldadapt_rx_asn_wait_for_fifo_flush_cnt                                    = 64,
		parameter hssi_pldadapt_rx_asn_wait_for_pma_pcie_sw_done_cnt                              = 64,
		parameter hssi_pldadapt_rx_bonding_dft_en                                                 = "dft_dis",
		parameter hssi_pldadapt_rx_bonding_dft_val                                                = "dft_0",
		parameter hssi_pldadapt_rx_chnl_bonding                                                   = "disable",
		parameter hssi_pldadapt_rx_clock_del_measure_enable                                       = "disable",
		parameter hssi_pldadapt_rx_hdpldadapt_csr_clk_hz                                          = 0,
		parameter hssi_pldadapt_rx_ctrl_plane_bonding                                             = "individual",
		parameter hssi_pldadapt_rx_ds_bypass_pipeln                                               = "ds_bypass_pipeln_dis",
		parameter hssi_pldadapt_rx_duplex_mode                                                    = "enable",
		parameter hssi_pldadapt_rx_dv_mode                                                        = "dv_mode_en",
		parameter hssi_pldadapt_rx_fifo_double_read                                               = "fifo_double_read_en",
		parameter hssi_pldadapt_rx_fifo_mode                                                      = "generic_basic",
		parameter hssi_pldadapt_rx_fifo_rd_clk_ins_sm_scg_en                                      = "enable",
		parameter hssi_pldadapt_rx_fifo_rd_clk_scg_en                                             = "disable",
		parameter hssi_pldadapt_rx_fifo_rd_clk_sel                                                = "fifo_rd_clk_pld_rx_clk1",
		parameter hssi_pldadapt_rx_fifo_stop_rd                                                   = "n_rd_empty",
		parameter hssi_pldadapt_rx_fifo_stop_wr                                                   = "n_wr_full",
		parameter hssi_pldadapt_rx_fifo_width                                                     = "fifo_double_width",
		parameter hssi_pldadapt_rx_fifo_wr_clk_del_sm_scg_en                                      = "enable",
		parameter hssi_pldadapt_rx_fifo_wr_clk_scg_en                                             = "disable",
		parameter hssi_pldadapt_rx_fifo_wr_clk_sel                                                = "fifo_wr_clk_rx_transfer_clk",
		parameter hssi_pldadapt_rx_free_run_div_clk                                               = "out_of_reset_sync",
		parameter hssi_pldadapt_rx_fsr_pld_10g_rx_crc32_err_rst_val                               = "reset_to_zero_crc32",
		parameter hssi_pldadapt_rx_fsr_pld_8g_sigdet_out_rst_val                                  = "reset_to_zero_sigdet",
		parameter hssi_pldadapt_rx_fsr_pld_ltd_b_rst_val                                          = "reset_to_one_ltdb",
		parameter hssi_pldadapt_rx_fsr_pld_ltr_rst_val                                            = "reset_to_zero_ltr",
		parameter hssi_pldadapt_rx_fsr_pld_rx_fifo_align_clr_rst_val                              = "reset_to_zero_alignclr",
		parameter hssi_pldadapt_rx_gb_rx_idwidth                                                  = "idwidth_64",
		parameter hssi_pldadapt_rx_gb_rx_odwidth                                                  = "odwidth_66",
		parameter hssi_pldadapt_rx_hip_mode                                                       = "disable_hip",
		parameter hssi_pldadapt_rx_hrdrst_align_bypass                                            = "enable",
		parameter hssi_pldadapt_rx_hrdrst_dll_lock_bypass                                         = "disable",
		parameter hssi_pldadapt_rx_hrdrst_rx_osc_clk_scg_en                                       = "disable",
		parameter hssi_pldadapt_rx_hrdrst_user_ctl_en                                             = "disable",
		parameter hssi_pldadapt_rx_indv                                                           = "indv_en",
		parameter hssi_pldadapt_rx_internal_clk1_sel1                                             = "pma_clks_or_txfiford_post_ct_mux_clk1_mux1",
		parameter hssi_pldadapt_rx_internal_clk1_sel2                                             = "pma_clks_clk1_mux2",
		parameter hssi_pldadapt_rx_internal_clk2_sel1                                             = "pma_clks_or_rxfifowr_post_ct_mux_clk2_mux1",
		parameter hssi_pldadapt_rx_internal_clk2_sel2                                             = "pma_clks_clk2_mux2",
		parameter hssi_pldadapt_rx_loopback_mode                                                  = "disable",
		parameter hssi_pldadapt_rx_low_latency_en                                                 = "disable",
		parameter hssi_pldadapt_rx_lpbk_mode                                                      = "disable",
		parameter hssi_pldadapt_rx_osc_clk_scg_en                                                 = "disable",
		parameter hssi_pldadapt_rx_phcomp_rd_del                                                  = "phcomp_rd_del2",
		parameter hssi_pldadapt_rx_pipe_enable                                                    = "disable",
		parameter hssi_pldadapt_rx_pipe_mode                                                      = "disable_pipe",
		parameter hssi_pldadapt_rx_hdpldadapt_pld_avmm1_clk_rowclk_hz                             = 0,
		parameter hssi_pldadapt_rx_hdpldadapt_pld_avmm2_clk_rowclk_hz                             = 0,
		parameter hssi_pldadapt_rx_pld_clk1_delay_en                                              = "enable",
		parameter hssi_pldadapt_rx_pld_clk1_delay_sel                                             = "delay_path13",
		parameter hssi_pldadapt_rx_pld_clk1_inv_en                                                = "disable",
		parameter hssi_pldadapt_rx_pld_clk1_sel                                                   = "pld_clk1_dcm",
		parameter hssi_pldadapt_rx_hdpldadapt_pld_rx_clk1_dcm_hz                                  = 390625000,
		parameter hssi_pldadapt_rx_hdpldadapt_pld_rx_clk1_rowclk_hz                               = 390625000,
		parameter hssi_pldadapt_rx_hdpldadapt_pld_sclk1_rowclk_hz                                 = 0,
		parameter hssi_pldadapt_rx_hdpldadapt_pld_sclk2_rowclk_hz                                 = 0,
		parameter hssi_pldadapt_rx_pma_hclk_scg_en                                                = "enable",
		parameter hssi_pldadapt_rx_powerdown_mode                                                 = "powerup",
		parameter hssi_pldadapt_rx_rx_datapath_tb_sel                                             = "cp_bond",
		parameter hssi_pldadapt_rx_rx_fastbond_rden                                               = "rden_ds_fast_us_fast",
		parameter hssi_pldadapt_rx_rx_fastbond_wren                                               = "wren_ds_del_us_del",
		parameter hssi_pldadapt_rx_rx_fifo_power_mode                                             = "full_width_full_depth",
		parameter hssi_pldadapt_rx_rx_fifo_read_latency_adjust                                    = "disable",
		parameter hssi_pldadapt_rx_rx_fifo_write_ctrl                                             = "blklock_ignore",
		parameter hssi_pldadapt_rx_rx_fifo_write_latency_adjust                                   = "disable",
		parameter hssi_pldadapt_rx_rx_osc_clock_setting                                           = "osc_clk_div_by1",
		parameter hssi_pldadapt_rx_rx_pld_8g_eidleinfersel_polling_bypass                         = "disable",
		parameter hssi_pldadapt_rx_rx_pld_pma_eye_monitor_polling_bypass                          = "disable",
		parameter hssi_pldadapt_rx_rx_pld_pma_pcie_switch_polling_bypass                          = "disable",
		parameter hssi_pldadapt_rx_rx_pld_pma_reser_out_polling_bypass                            = "disable",
		parameter hssi_pldadapt_rx_rx_prbs_flags_sr_enable                                        = "disable",
		parameter hssi_pldadapt_rx_rx_true_b2b                                                    = "b2b",
		parameter hssi_pldadapt_rx_rx_usertest_sel                                                = "enable",
		parameter hssi_pldadapt_rx_rxfifo_empty                                                   = "empty_dw",
		parameter hssi_pldadapt_rx_rxfifo_full                                                    = "full_non_pc_dw",
		parameter hssi_pldadapt_rx_rxfifo_mode                                                    = "rxgeneric_basic",
		parameter hssi_pldadapt_rx_rxfifo_pempty                                                  = 13,
		parameter hssi_pldadapt_rx_rxfifo_pfull                                                   = 51,
		parameter hssi_pldadapt_rx_rxfiford_post_ct_sel                                           = "rxfiford_sclk_post_ct",
		parameter hssi_pldadapt_rx_rxfifowr_post_ct_sel                                           = "rxfifowr_sclk_post_ct",
		parameter hssi_pldadapt_rx_sclk_sel                                                       = "sclk1_rowclk",
		parameter hssi_pldadapt_rx_hdpldadapt_speed_grade                                         = "dash_2",
		parameter hssi_pldadapt_rx_stretch_num_stages                                             = "two_stage",
		parameter hssi_pldadapt_rx_sup_mode                                                       = "user_mode",
		parameter hssi_pldadapt_rx_txfiford_post_ct_sel                                           = "txfiford_sclk_post_ct",
		parameter hssi_pldadapt_rx_txfifowr_post_ct_sel                                           = "txfifowr_sclk_post_ct",
		parameter hssi_pldadapt_rx_us_bypass_pipeln                                               = "us_bypass_pipeln_dis",
		parameter hssi_pldadapt_rx_word_align                                                     = "wa_en",
		parameter hssi_pldadapt_rx_word_align_enable                                              = "enable",
		parameter hssi_pldadapt_rx_silicon_rev                                                    = "14nm5cr2",
		parameter hssi_pldadapt_tx_aib_clk1_sel                                                   = "aib_clk1_pld_pcs_tx_clk_out",
		parameter hssi_pldadapt_tx_aib_clk2_sel                                                   = "aib_clk2_pld_pma_clkdiv_tx_user",
		parameter hssi_pldadapt_tx_hdpldadapt_aib_fabric_pld_pma_hclk_hz                          = 0,
		parameter hssi_pldadapt_tx_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                        = 805664062,
		parameter hssi_pldadapt_tx_bonding_dft_en                                                 = "dft_dis",
		parameter hssi_pldadapt_tx_bonding_dft_val                                                = "dft_0",
		parameter hssi_pldadapt_tx_chnl_bonding                                                   = "disable",
		parameter hssi_pldadapt_tx_hdpldadapt_csr_clk_hz                                          = 0,
		parameter hssi_pldadapt_tx_ctrl_plane_bonding                                             = "individual",
		parameter hssi_pldadapt_tx_ds_bypass_pipeln                                               = "ds_bypass_pipeln_dis",
		parameter hssi_pldadapt_tx_duplex_mode                                                    = "enable",
		parameter hssi_pldadapt_tx_dv_bond                                                        = "dv_bond_dis",
		parameter hssi_pldadapt_tx_dv_gen                                                         = "dv_gen_en",
		parameter hssi_pldadapt_tx_fifo_double_write                                              = "fifo_double_write_en",
		parameter hssi_pldadapt_tx_fifo_mode                                                      = "generic_basic",
		parameter hssi_pldadapt_tx_fifo_rd_clk_frm_gen_scg_en                                     = "enable",
		parameter hssi_pldadapt_tx_fifo_rd_clk_scg_en                                             = "disable",
		parameter hssi_pldadapt_tx_fifo_rd_clk_sel                                                = "fifo_rd_pma_aib_tx_clk",
		parameter hssi_pldadapt_tx_fifo_stop_rd                                                   = "n_rd_empty",
		parameter hssi_pldadapt_tx_fifo_stop_wr                                                   = "n_wr_full",
		parameter hssi_pldadapt_tx_fifo_width                                                     = "fifo_double_width",
		parameter hssi_pldadapt_tx_fifo_wr_clk_scg_en                                             = "disable",
		parameter hssi_pldadapt_tx_fpll_shared_direct_async_in_sel                                = "fpll_shared_direct_async_in_rowclk",
		parameter hssi_pldadapt_tx_frmgen_burst                                                   = "frmgen_burst_dis",
		parameter hssi_pldadapt_tx_frmgen_bypass                                                  = "frmgen_bypass_en",
		parameter hssi_pldadapt_tx_frmgen_mfrm_length                                             = 2048,
		parameter hssi_pldadapt_tx_frmgen_pipeln                                                  = "frmgen_pipeln_en",
		parameter hssi_pldadapt_tx_frmgen_pyld_ins                                                = "frmgen_pyld_ins_dis",
		parameter hssi_pldadapt_tx_frmgen_wordslip                                                = "frmgen_wordslip_dis",
		parameter hssi_pldadapt_tx_fsr_hip_fsr_in_bit0_rst_val                                    = "reset_to_one_hfsrin0",
		parameter hssi_pldadapt_tx_fsr_hip_fsr_in_bit1_rst_val                                    = "reset_to_one_hfsrin1",
		parameter hssi_pldadapt_tx_fsr_hip_fsr_in_bit2_rst_val                                    = "reset_to_one_hfsrin2",
		parameter hssi_pldadapt_tx_fsr_hip_fsr_in_bit3_rst_val                                    = "reset_to_zero_hfsrin3",
		parameter hssi_pldadapt_tx_fsr_hip_fsr_out_bit0_rst_val                                   = "reset_to_one_hfsrout0",
		parameter hssi_pldadapt_tx_fsr_hip_fsr_out_bit1_rst_val                                   = "reset_to_one_hfsrout1",
		parameter hssi_pldadapt_tx_fsr_hip_fsr_out_bit2_rst_val                                   = "reset_to_zero_hfsrout2",
		parameter hssi_pldadapt_tx_fsr_hip_fsr_out_bit3_rst_val                                   = "reset_to_zero_hfsrout3",
		parameter hssi_pldadapt_tx_fsr_mask_tx_pll_rst_val                                        = "reset_to_zero_maskpll",
		parameter hssi_pldadapt_tx_fsr_pld_txelecidle_rst_val                                     = "reset_to_zero_txelec",
		parameter hssi_pldadapt_tx_gb_tx_idwidth                                                  = "idwidth_66",
		parameter hssi_pldadapt_tx_gb_tx_odwidth                                                  = "odwidth_64",
		parameter hssi_pldadapt_tx_hip_mode                                                       = "disable_hip",
		parameter hssi_pldadapt_tx_hip_osc_clk_scg_en                                             = "enable",
		parameter hssi_pldadapt_tx_hrdrst_dcd_cal_done_bypass                                     = "disable",
		parameter hssi_pldadapt_tx_hrdrst_rx_osc_clk_scg_en                                       = "disable",
		parameter hssi_pldadapt_tx_hrdrst_user_ctl_en                                             = "disable",
		parameter hssi_pldadapt_tx_indv                                                           = "indv_en",
		parameter hssi_pldadapt_tx_loopback_mode                                                  = "disable",
		parameter hssi_pldadapt_tx_low_latency_en                                                 = "disable",
		parameter hssi_pldadapt_tx_osc_clk_scg_en                                                 = "disable",
		parameter hssi_pldadapt_tx_phcomp_rd_del                                                  = "phcomp_rd_del2",
		parameter hssi_pldadapt_tx_pipe_mode                                                      = "disable_pipe",
		parameter hssi_pldadapt_tx_hdpldadapt_pld_avmm1_clk_rowclk_hz                             = 0,
		parameter hssi_pldadapt_tx_hdpldadapt_pld_avmm2_clk_rowclk_hz                             = 0,
		parameter hssi_pldadapt_tx_pld_clk1_delay_en                                              = "enable",
		parameter hssi_pldadapt_tx_pld_clk1_delay_sel                                             = "delay_path15",
		parameter hssi_pldadapt_tx_pld_clk1_inv_en                                                = "disable",
		parameter hssi_pldadapt_tx_pld_clk1_sel                                                   = "pld_clk1_dcm",
		parameter hssi_pldadapt_tx_pld_clk2_sel                                                   = "pld_clk2_dcm",
		parameter hssi_pldadapt_tx_hdpldadapt_pld_sclk1_rowclk_hz                                 = 0,
		parameter hssi_pldadapt_tx_hdpldadapt_pld_sclk2_rowclk_hz                                 = 0,
		parameter hssi_pldadapt_tx_hdpldadapt_pld_tx_clk1_dcm_hz                                  = 390625000,
		parameter hssi_pldadapt_tx_hdpldadapt_pld_tx_clk1_rowclk_hz                               = 390625000,
		parameter hssi_pldadapt_tx_hdpldadapt_pld_tx_clk2_dcm_hz                                  = 805664062,
		parameter hssi_pldadapt_tx_hdpldadapt_pld_tx_clk2_rowclk_hz                               = 805664062,
		parameter hssi_pldadapt_tx_pma_aib_tx_clk_expected_setting                                = "x2",
		parameter hssi_pldadapt_tx_powerdown_mode                                                 = "powerup",
		parameter hssi_pldadapt_tx_sh_err                                                         = "sh_err_dis",
		parameter hssi_pldadapt_tx_hdpldadapt_speed_grade                                         = "dash_2",
		parameter hssi_pldadapt_tx_stretch_num_stages                                             = "two_stage",
		parameter hssi_pldadapt_tx_sup_mode                                                       = "user_mode",
		parameter hssi_pldadapt_tx_tx_datapath_tb_sel                                             = "cp_bond",
		parameter hssi_pldadapt_tx_tx_fastbond_rden                                               = "rden_ds_fast_us_fast",
		parameter hssi_pldadapt_tx_tx_fastbond_wren                                               = "wren_ds_fast_us_fast",
		parameter hssi_pldadapt_tx_tx_fifo_power_mode                                             = "full_width_full_depth",
		parameter hssi_pldadapt_tx_tx_fifo_read_latency_adjust                                    = "disable",
		parameter hssi_pldadapt_tx_tx_fifo_write_latency_adjust                                   = "disable",
		parameter hssi_pldadapt_tx_tx_hip_aib_ssr_in_polling_bypass                               = "disable",
		parameter hssi_pldadapt_tx_tx_osc_clock_setting                                           = "osc_clk_div_by1",
		parameter hssi_pldadapt_tx_tx_pld_10g_tx_bitslip_polling_bypass                           = "disable",
		parameter hssi_pldadapt_tx_tx_pld_8g_tx_boundary_sel_polling_bypass                       = "disable",
		parameter hssi_pldadapt_tx_tx_pld_pma_fpll_cnt_sel_polling_bypass                         = "disable",
		parameter hssi_pldadapt_tx_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                = "disable",
		parameter hssi_pldadapt_tx_tx_usertest_sel                                                = "enable",
		parameter hssi_pldadapt_tx_txfifo_empty                                                   = "empty_default",
		parameter hssi_pldadapt_tx_txfifo_full                                                    = "full_non_pc_dw",
		parameter hssi_pldadapt_tx_txfifo_mode                                                    = "txgeneric_basic",
		parameter hssi_pldadapt_tx_txfifo_pempty                                                  = 6,
		parameter hssi_pldadapt_tx_txfifo_pfull                                                   = 26,
		parameter hssi_pldadapt_tx_us_bypass_pipeln                                               = "us_bypass_pipeln_dis",
		parameter hssi_pldadapt_tx_word_align_enable                                              = "enable",
		parameter hssi_pldadapt_tx_word_mark                                                      = "wm_en",
		parameter hssi_pldadapt_tx_silicon_rev                                                    = "14nm5cr2",
		parameter cdr_pll_analog_mode                                                             = "user_custom",
		parameter cdr_pll_atb_select_control                                                      = "atb_off",
		parameter cdr_pll_auto_reset_on                                                           = "auto_reset_off",
		parameter cdr_pll_bandwidth_range_high                                                    = "1",
		parameter cdr_pll_bandwidth_range_low                                                     = "1",
		parameter cdr_pll_bbpd_data_pattern_filter_select                                         = "bbpd_data_pat_off",
		parameter cdr_pll_bti_protected                                                           = "false",
		parameter cdr_pll_bw_mode                                                                 = "mid_bw",
		parameter cdr_pll_bypass_a_edge                                                           = "bypass_a_edge_off",
		parameter cdr_pll_cal_vco_count_length                                                    = "sel_8b_count",
		parameter cdr_pll_pm_cr2_rx_path_cdr_clock_enable                                         = "cdr_clock_disable",
		parameter cdr_pll_cdr_d2a_enb                                                             = "bti_d2a_disable",
		parameter cdr_pll_cdr_odi_select                                                          = "sel_cdr",
		parameter cdr_pll_cdr_phaselock_mode                                                      = "no_ignore_lock",
		parameter cdr_pll_cdr_powerdown_mode                                                      = "power_up",
		parameter cdr_pll_chgpmp_current_dn_pd                                                    = "cp_current_pd_dn_setting4",
		parameter cdr_pll_chgpmp_current_dn_trim                                                  = "cp_current_trimming_dn_setting0",
		parameter cdr_pll_chgpmp_current_pfd                                                      = "cp_current_pfd_setting1",
		parameter cdr_pll_chgpmp_current_up_pd                                                    = "cp_current_pd_up_setting4",
		parameter cdr_pll_chgpmp_current_up_trim                                                  = "cp_current_trimming_up_setting0",
		parameter cdr_pll_chgpmp_dn_pd_trim_double                                                = "normal_dn_trim_current",
		parameter cdr_pll_chgpmp_replicate                                                        = "disable_replica_bias_ctrl",
		parameter cdr_pll_chgpmp_testmode                                                         = "cp_test_disable",
		parameter cdr_pll_chgpmp_up_pd_trim_double                                                = "normal_up_trim_current",
		parameter cdr_pll_chgpmp_vccreg                                                           = "vreg_fw0",
		parameter cdr_pll_clk0_dfe_tfall_adj                                                      = "clk0_dfe_tf0",
		parameter cdr_pll_clk0_dfe_trise_adj                                                      = "clk0_dfe_tr0",
		parameter cdr_pll_clk180_dfe_tfall_adj                                                    = "clk180_dfe_tf0",
		parameter cdr_pll_clk180_dfe_trise_adj                                                    = "clk180_dfe_tr0",
		parameter cdr_pll_clk270_dfe_tfall_adj                                                    = "clk270_dfe_tf0",
		parameter cdr_pll_clk270_dfe_trise_adj                                                    = "clk270_dfe_tr0",
		parameter cdr_pll_clk90_dfe_tfall_adj                                                     = "clk90_dfe_tf0",
		parameter cdr_pll_clk90_dfe_trise_adj                                                     = "clk90_dfe_tr0",
		parameter cdr_pll_clklow_mux_select                                                       = "clklow_mux_cdr_fbclk",
		parameter cdr_pll_datarate_bps                                                            = "25781250000",
		parameter cdr_pll_diag_loopback_enable                                                    = "no_diag_rev_loopback",
		parameter cdr_pll_disable_up_dn                                                           = "normal_mode",
		parameter cdr_pll_f_max_cmu_out_freq                                                      = "1",
		parameter cdr_pll_f_max_m_counter                                                         = "1",
		parameter cdr_pll_f_max_pfd                                                               = "350000000",
		parameter cdr_pll_f_max_ref                                                               = "800000000",
		parameter cdr_pll_f_max_vco                                                               = "14150000000",
		parameter cdr_pll_f_min_gt_channel                                                        = "8700000000",
		parameter cdr_pll_f_min_pfd                                                               = "25000000",
		parameter cdr_pll_f_min_ref                                                               = "25000000",
		parameter cdr_pll_f_min_vco                                                               = "7000000000",
		parameter cdr_pll_fref_clklow_div                                                         = 2,
		parameter cdr_pll_fref_mux_select                                                         = "fref_mux_cdr_refclk",
		parameter cdr_pll_gpon_lck2ref_control                                                    = "gpon_lck2ref_off",
		parameter cdr_pll_initial_settings                                                        = "true",
		parameter cdr_pll_lck2ref_delay_control                                                   = "lck2ref_delay_2",
		parameter cdr_pll_lf_resistor_pd                                                          = "lf_pd_setting3",
		parameter cdr_pll_lf_resistor_pfd                                                         = "lf_pfd_setting3",
		parameter cdr_pll_lf_ripple_cap                                                           = "lf_no_ripple",
		parameter cdr_pll_loop_filter_bias_select                                                 = "lpflt_bias_7",
		parameter cdr_pll_loopback_mode                                                           = "loopback_disabled",
		parameter cdr_pll_lpd_counter                                                             = 1,
		parameter cdr_pll_lpfd_counter                                                            = 2,
		parameter cdr_pll_ltd_ltr_micro_controller_select                                         = "ltd_ltr_pcs",
		parameter cdr_pll_mcnt_div                                                                = 20,
		parameter cdr_pll_n_counter                                                               = 2,
		parameter cdr_pll_ncnt_div                                                                = 2,
		parameter cdr_pll_optimal                                                                 = "true",
		parameter cdr_pll_out_freq                                                                = "12890625000",
		parameter cdr_pll_pcie_gen                                                                = "non_pcie",
		parameter cdr_pll_pd_fastlock_mode                                                        = "fast_lock_disable",
		parameter cdr_pll_pd_l_counter                                                            = 1,
		parameter cdr_pll_pfd_l_counter                                                           = 2,
		parameter cdr_pll_position                                                                = "position0",
		parameter cdr_pll_power_mode                                                              = "high_perf",
		parameter cdr_pll_powermode_ac_bbpd                                                       = "bbpd_ac_on",
		parameter cdr_pll_powermode_ac_rvcotop                                                    = "rvcotop_ac_div1",
		parameter cdr_pll_powermode_ac_txpll                                                      = "txpll_ac_off",
		parameter cdr_pll_powermode_dc_bbpd                                                       = "bbpd_dc_on",
		parameter cdr_pll_powermode_dc_rvcotop                                                    = "rvcotop_dc_div1",
		parameter cdr_pll_powermode_dc_txpll                                                      = "powerdown_txpll",
		parameter cdr_pll_primary_use                                                             = "cdr",
		parameter cdr_pll_prot_mode                                                               = "basic_rx",
		parameter cdr_pll_reference_clock_frequency                                               = "644531250",
		parameter cdr_pll_requires_gt_capable_channel                                             = "true",
		parameter cdr_pll_reverse_serial_loopback                                                 = "no_loopback",
		parameter cdr_pll_set_cdr_input_freq_range                                                = 0,
		parameter cdr_pll_set_cdr_v2i_enable                                                      = "enable_v2i_bias",
		parameter cdr_pll_set_cdr_vco_reset                                                       = "vco_normal",
		parameter cdr_pll_set_cdr_vco_speed                                                       = 0,
		parameter cdr_pll_set_cdr_vco_speed_fix                                                   = 120,
		parameter cdr_pll_set_cdr_vco_speed_pciegen3                                              = "cdr_vco_max_speedbin_pciegen3",
		parameter cdr_pll_speed_grade                                                             = "e2",
		parameter cdr_pll_sup_mode                                                                = "user_mode",
		parameter cdr_pll_tx_pll_prot_mode                                                        = "txpll_unused",
		parameter cdr_pll_txpll_hclk_driver_enable                                                = "hclk_off",
		parameter cdr_pll_rstb                                                                    = "cdr_lf_reset_off",
		parameter cdr_pll_pm_cr2_tx_rx_uc_dyn_reconfig                                            = "uc_dyn_reconfig_off",
		parameter cdr_pll_uc_ro_cal                                                               = "uc_ro_cal_off",
		parameter cdr_pll_vco_bypass                                                              = "false",
		parameter cdr_pll_vco_freq                                                                = "12890625000",
		parameter cdr_pll_vco_overrange_voltage                                                   = "vco_overrange_off",
		parameter cdr_pll_vco_underrange_voltage                                                  = "vco_underange_off",
		parameter cdr_pll_vreg_output                                                             = "vccdreg_nominal",
		parameter cdr_pll_direct_fb                                                               = "direct_fb",
		parameter cdr_pll_iqclk_sel                                                               = "power_down",
		parameter cdr_pll_silicon_rev                                                             = "14nm5cr2",
		parameter cdr_pll_pma_width                                                               = 64,
		parameter cdr_pll_cgb_div                                                                 = 1,
		parameter cdr_pll_is_cascaded_pll                                                         = "false",
		parameter pma_rx_buf_act_isource_disable                                                  = "isrc_dis",
		parameter pma_rx_buf_advanced_mode                                                        = "false",
		parameter pma_rx_buf_pm_cr2_rx_path_analog_mode                                           = "user_custom",
		parameter pma_rx_buf_bodybias_enable                                                      = "bodybias_dis",
		parameter pma_rx_buf_bodybias_select                                                      = "bodybias_sel1",
		parameter pma_rx_buf_bypass_ctle_rf_cal                                                   = "use_dprio_rfcal",
		parameter pma_rx_buf_clk_divrx_en                                                         = "normal_clk",
		parameter pma_rx_buf_const_gm_en                                                          = "cgm_en_1",
		parameter pma_rx_buf_ctle_ac_gain                                                         = 0,
		parameter pma_rx_buf_ctle_eq_gain                                                         = 0,
		parameter pma_rx_buf_ctle_hires_bypass                                                    = "ctle_hires_en",
		parameter pma_rx_buf_ctle_oc_ib_sel                                                       = "ib_oc_bw3",
		parameter pma_rx_buf_ctle_oc_sign                                                         = "add_i_2_p_eq",
		parameter pma_rx_buf_ctle_rf_cal                                                          = 1,
		parameter pma_rx_buf_ctle_tia_isel                                                        = "ib_tia_bw3",
		parameter pma_rx_buf_pm_cr2_tx_rx_cvp_mode                                                = "cvp_off",
		parameter pma_rx_buf_datarate_bps                                                         = "25781250000",
		parameter pma_rx_buf_pm_cr2_rx_path_datarate_bps                                          = "25781250000",
		parameter pma_rx_buf_pm_cr2_rx_path_datawidth                                             = 64,
		parameter pma_rx_buf_diag_lp_en                                                           = "dlp_off",
		parameter pma_rx_buf_eq_bw_sel                                                            = "eq_bw_3",
		parameter pma_rx_buf_eq_cdgen_sel                                                         = "eq_cdgen_0",
		parameter pma_rx_buf_eq_isel                                                              = "eq_isel_1",
		parameter pma_rx_buf_eq_sel                                                               = "eq_sel_3",
		parameter pma_rx_buf_pm_cr2_rx_path_gt_enabled                                            = "enable",
		parameter pma_rx_buf_initial_settings                                                     = "true",
		parameter pma_rx_buf_pm_cr2_rx_path_initial_settings                                      = "true",
		parameter pma_rx_buf_pm_cr2_rx_path_jtag_hys                                              = "hys_increase_disable",
		parameter pma_rx_buf_pm_cr2_rx_path_jtag_lp                                               = "lp_off",
		parameter pma_rx_buf_pm_cr2_rx_path_link                                                  = "sr",
		parameter pma_rx_buf_xrx_path_xcdr_deser_xcdr_loopback_mode                               = "loopback_disabled",
		parameter pma_rx_buf_loopback_modes                                                       = "lpbk_disable",
		parameter pma_rx_buf_offset_cancellation_coarse                                           = "coarse_setting_0",
		parameter pma_rx_buf_offset_rx_cal_en                                                     = "rx_oc_dis",
		parameter pma_rx_buf_optimal                                                              = "true",
		parameter pma_rx_buf_pm_cr2_rx_path_optimal                                               = "true",
		parameter pma_rx_buf_pm_cr2_tx_rx_pcie_gen                                                = "non_pcie",
		parameter pma_rx_buf_pm_cr2_tx_rx_pcie_gen_bitwidth                                       = "pcie_gen3_32b",
		parameter pma_rx_buf_pdb_rx                                                               = "normal_rx_on",
		parameter pma_rx_buf_pm_cr2_rx_path_pma_rx_divclk_hz                                      = "402832031",
		parameter pma_rx_buf_power_mode                                                           = "high_perf",
		parameter pma_rx_buf_pm_cr2_rx_path_power_mode                                            = "high_perf",
		parameter pma_rx_buf_pm_cr2_rx_path_power_rail_eht                                        = 0,
		parameter pma_rx_buf_power_rail_er                                                        = 0,
		parameter pma_rx_buf_pm_cr2_rx_path_power_rail_er                                         = 1120,
		parameter pma_rx_buf_powermode_ac_ctle                                                    = "ctle_pwr_ac4",
		parameter pma_rx_buf_powermode_ac_vcm                                                     = "vcm_pwr_ac3",
		parameter pma_rx_buf_powermode_ac_vga                                                     = "vga_pwr_ac_full",
		parameter pma_rx_buf_powermode_dc_ctle                                                    = "ctle_pwr_dc1",
		parameter pma_rx_buf_powermode_dc_vcm                                                     = "vcm_pwr_dc3",
		parameter pma_rx_buf_powermode_dc_vga                                                     = "vga_pwr_dc_full",
		parameter pma_rx_buf_prot_mode                                                            = "basic_rx",
		parameter pma_rx_buf_pm_cr2_rx_path_prot_mode                                             = "basic_rx",
		parameter pma_rx_buf_qpi_afe_en                                                           = "ctle_mode_en",
		parameter pma_rx_buf_qpi_enable                                                           = "non_qpi_mode",
		parameter pma_rx_buf_refclk_en                                                            = "disable",
		parameter pma_rx_buf_rx_atb_select                                                        = "atb_disable",
		parameter pma_rx_buf_rx_vga_oc_en                                                         = "vga_cal_off",
		parameter pma_rx_buf_sel_vcm_ctle                                                         = "vocm_eq_fixed",
		parameter pma_rx_buf_sel_vcm_tia                                                          = "vocm_tia_fixed",
		parameter pma_rx_buf_pm_cr2_rx_path_speed_grade                                           = "e2",
		parameter pma_rx_buf_sup_mode                                                             = "user_mode",
		parameter pma_rx_buf_pm_cr2_rx_path_sup_mode                                              = "user_mode",
		parameter pma_rx_buf_term_sel                                                             = "r_r4",
		parameter pma_rx_buf_term_sync_bypass                                                     = "bypass_termsync",
		parameter pma_rx_buf_term_tri_enable                                                      = "disable_tri",
		parameter pma_rx_buf_pm_cr2_tx_rx_testmux_select                                          = "setting0",
		parameter pma_rx_buf_tia_sel                                                              = "tia_sel_1",
		parameter pma_rx_buf_pm_cr2_rx_path_tile_type                                             = "h",
		parameter pma_rx_buf_pm_cr2_rx_path_uc_cal_clk_bypass                                     = "cal_clk_0",
		parameter pma_rx_buf_pm_cr2_rx_path_uc_cal_enable                                         = "rx_cal_off",
		parameter pma_rx_buf_pm_cr2_tx_rx_uc_odi_eye_left                                         = "uc_odi_eye_left_off",
		parameter pma_rx_buf_pm_cr2_tx_rx_uc_odi_eye_right                                        = "uc_odi_eye_right_off",
		parameter pma_rx_buf_pm_cr2_rx_path_uc_pcie_sw                                            = "uc_pcie_gen1",
		parameter pma_rx_buf_pm_cr2_tx_rx_uc_rx_cal                                               = "uc_rx_cal_on",
		parameter pma_rx_buf_vcm_cal_i                                                            = 4,
		parameter pma_rx_buf_vcm_current_add                                                      = "vcm_current_3",
		parameter pma_rx_buf_vcm_sel                                                              = "vcm_l0",
		parameter pma_rx_buf_vcm_sel_vccref                                                       = 6,
		parameter pma_rx_buf_vga_dc_gain                                                          = 0,
		parameter pma_rx_buf_vga_halfbw_en                                                        = "vga_half_bw_disabled",
		parameter pma_rx_buf_vga_ib_max_en                                                        = "vga_ib_max_enable",
		parameter pma_rx_buf_vga_mode                                                             = "vga_off",
		parameter pma_rx_buf_silicon_rev                                                          = "14nm5cr2",
		parameter hssi_adapt_rx_adapter_lpbk_mode                                                 = "disable",
		parameter hssi_adapt_rx_hd_hssiadapt_aib_hssi_pld_sclk_hz                                 = 0,
		parameter hssi_adapt_rx_aib_lpbk_mode                                                     = "disable",
		parameter hssi_adapt_rx_align_del                                                         = "align_del_dis",
		parameter hssi_adapt_rx_asn_bypass_clock_gate                                             = "disable",
		parameter hssi_adapt_rx_asn_bypass_pma_pcie_sw_done                                       = "disable",
		parameter hssi_adapt_rx_asn_wait_for_clock_gate_cnt                                       = 32,
		parameter hssi_adapt_rx_asn_wait_for_dll_reset_cnt                                        = 32,
		parameter hssi_adapt_rx_asn_wait_for_fifo_flush_cnt                                       = 32,
		parameter hssi_adapt_rx_asn_wait_for_pma_pcie_sw_done_cnt                                 = 32,
		parameter hssi_adapt_rx_async_direct_hip_en                                               = "disable",
		parameter hssi_adapt_rx_bonding_dft_en                                                    = "dft_dis",
		parameter hssi_adapt_rx_bonding_dft_val                                                   = "dft_0",
		parameter hssi_adapt_rx_chnl_bonding                                                      = "disable",
		parameter hssi_adapt_rx_clock_del_measure_enable                                          = "disable",
		parameter hssi_adapt_rx_control_del                                                       = "control_del_none",
		parameter hssi_adapt_rx_hd_hssiadapt_csr_clk_hz                                           = 0,
		parameter hssi_adapt_rx_ctrl_plane_bonding                                                = "individual",
		parameter hssi_adapt_rx_datapath_mapping_mode                                             = "map_10g_2x2x_2x1x_fifo",
		parameter hssi_adapt_rx_ds_bypass_pipeln                                                  = "ds_bypass_pipeln_dis",
		parameter hssi_adapt_rx_duplex_mode                                                       = "enable",
		parameter hssi_adapt_rx_dyn_clk_sw_en                                                     = "disable",
		parameter hssi_adapt_rx_fifo_double_write                                                 = "fifo_double_write_en",
		parameter hssi_adapt_rx_fifo_mode                                                         = "phase_comp",
		parameter hssi_adapt_rx_fifo_rd_clk_scg_en                                                = "disable",
		parameter hssi_adapt_rx_fifo_rd_clk_sel                                                   = "fifo_rd_pma_aib_rx_clk",
		parameter hssi_adapt_rx_fifo_stop_rd                                                      = "rd_empty",
		parameter hssi_adapt_rx_fifo_stop_wr                                                      = "n_wr_full",
		parameter hssi_adapt_rx_fifo_width                                                        = "fifo_double_width",
		parameter hssi_adapt_rx_fifo_wr_clk_scg_en                                                = "disable",
		parameter hssi_adapt_rx_fifo_wr_clk_sel                                                   = "fifo_wr_pld_pcs_rx_clk_out",
		parameter hssi_adapt_rx_force_align                                                       = "force_align_dis",
		parameter hssi_adapt_rx_free_run_div_clk                                                  = "out_of_reset_sync",
		parameter hssi_adapt_rx_fsr_pld_10g_rx_crc32_err_rst_val                                  = "reset_to_zero_crc32",
		parameter hssi_adapt_rx_fsr_pld_8g_sigdet_out_rst_val                                     = "reset_to_zero_sigdet",
		parameter hssi_adapt_rx_fsr_pld_ltd_b_rst_val                                             = "reset_to_one_ltdb",
		parameter hssi_adapt_rx_fsr_pld_ltr_rst_val                                               = "reset_to_zero_ltr",
		parameter hssi_adapt_rx_fsr_pld_rx_fifo_align_clr_rst_val                                 = "reset_to_zero_alignclr",
		parameter hssi_adapt_rx_hd_hssiadapt_hip_aib_clk_2x_hz                                    = 0,
		parameter hssi_adapt_rx_hd_hssiadapt_hip_aib_clk_hz                                       = 0,
		parameter hssi_adapt_rx_hip_mode                                                          = "disable_hip",
		parameter hssi_adapt_rx_hrdrst_dcd_cal_done_bypass                                        = "disable",
		parameter hssi_adapt_rx_hrdrst_rx_osc_clk_scg_en                                          = "disable",
		parameter hssi_adapt_rx_hrdrst_user_ctl_en                                                = "disable",
		parameter hssi_adapt_rx_indv                                                              = "indv_en",
		parameter hssi_adapt_rx_internal_clk1_sel                                                 = "pld_pma_tx_clk_out_clk1",
		parameter hssi_adapt_rx_internal_clk1_sel0                                                = "pma_clks_or_txfifowr_post_ct_or_txfiford_pre_or_post_ct_mux_clk1_mux0",
		parameter hssi_adapt_rx_internal_clk1_sel1                                                = "pma_clks_or_txfiford_pre_or_post_ct_mux_clk1_mux1",
		parameter hssi_adapt_rx_internal_clk1_sel2                                                = "pma_clks_or_txfiford_pre_ct_mux_clk1_mux2",
		parameter hssi_adapt_rx_internal_clk1_sel3                                                = "pma_clks_clk1_mux3",
		parameter hssi_adapt_rx_internal_clk2_sel                                                 = "pld_pma_tx_clk_out_clk2",
		parameter hssi_adapt_rx_internal_clk2_sel0                                                = "pma_clks_or_rxfiford_post_ct_or_rxfifowr_pre_or_post_ct_mux_clk2_mux0",
		parameter hssi_adapt_rx_internal_clk2_sel1                                                = "pma_clks_or_rxfifowr_pre_or_post_ct_mux_clk2_mux1",
		parameter hssi_adapt_rx_internal_clk2_sel2                                                = "pma_clks_or_rxfifowr_pre_ct_mux_clk2_mux2",
		parameter hssi_adapt_rx_internal_clk2_sel3                                                = "pma_clks_clk2_mux3",
		parameter hssi_adapt_rx_loopback_mode                                                     = "loopback_disable",
		parameter hssi_adapt_rx_osc_clk_scg_en                                                    = "disable",
		parameter hssi_adapt_rx_phcomp_rd_del                                                     = "phcomp_rd_del3",
		parameter hssi_adapt_rx_pipe_mode                                                         = "disable_pipe",
		parameter hssi_adapt_rx_hd_hssiadapt_pld_pcs_rx_clk_out_hz                                = 402832031,
		parameter hssi_adapt_rx_hd_hssiadapt_pld_pma_hclk_hz                                      = 0,
		parameter hssi_adapt_rx_pma_aib_rx_clk_expected_setting                                   = "x2",
		parameter hssi_adapt_rx_hd_hssiadapt_pma_aib_rx_clk_hz                                    = 0,
		parameter hssi_adapt_rx_pma_coreclkin_sel                                                 = "pma_coreclkin_pld_sel",
		parameter hssi_adapt_rx_pma_hclk_scg_en                                                   = "enable",
		parameter hssi_adapt_rx_powerdown_mode                                                    = "powerup",
		parameter hssi_adapt_rx_rx_10g_krfec_rx_diag_data_status_polling_bypass                   = "disable",
		parameter hssi_adapt_rx_rx_adp_go_b4txeq_en                                               = "enable",
		parameter hssi_adapt_rx_rx_datapath_tb_sel                                                = "cp_bond",
		parameter hssi_adapt_rx_rx_eq_iteration                                                   = "cycles_32",
		parameter hssi_adapt_rx_rx_fifo_power_mode                                                = "full_width_full_depth",
		parameter hssi_adapt_rx_rx_fifo_read_latency_adjust                                       = "disable",
		parameter hssi_adapt_rx_rx_fifo_write_latency_adjust                                      = "disable",
		parameter hssi_adapt_rx_rx_invalid_no_change                                              = "disable",
		parameter hssi_adapt_rx_rx_osc_clock_setting                                              = "osc_clk_div_by1",
		parameter hssi_adapt_rx_rx_parity_sel                                                     = "func_sel",
		parameter hssi_adapt_rx_rx_pcs_testbus_sel                                                = "direct_tr_tb_bit0_sel",
		parameter hssi_adapt_rx_rx_pcspma_testbus_sel                                             = "enable",
		parameter hssi_adapt_rx_rx_pld_8g_a1a2_k1k2_flag_polling_bypass                           = "disable",
		parameter hssi_adapt_rx_rx_pld_8g_wa_boundary_polling_bypass                              = "disable",
		parameter hssi_adapt_rx_rx_pld_pma_pcie_sw_done_polling_bypass                            = "disable",
		parameter hssi_adapt_rx_rx_pld_pma_reser_in_polling_bypass                                = "disable",
		parameter hssi_adapt_rx_rx_pld_pma_testbus_polling_bypass                                 = "disable",
		parameter hssi_adapt_rx_rx_pld_test_data_polling_bypass                                   = "disable",
		parameter hssi_adapt_rx_rx_pma_rstn_cycles                                                = "four_cycles",
		parameter hssi_adapt_rx_rx_pma_rstn_en                                                    = "disable",
		parameter hssi_adapt_rx_rx_post_cursor_en                                                 = "disable",
		parameter hssi_adapt_rx_rx_pre_cursor_en                                                  = "disable",
		parameter hssi_adapt_rx_rx_rmfflag_stretch_enable                                         = "enable",
		parameter hssi_adapt_rx_rx_rmfflag_stretch_num_stages                                     = "rmfflag_two_stage",
		parameter hssi_adapt_rx_rx_rxeq_en                                                        = "disable",
		parameter hssi_adapt_rx_rx_txeq_en                                                        = "disable",
		parameter hssi_adapt_rx_rx_txeq_time                                                      = 64,
		parameter hssi_adapt_rx_rx_use_rxvalid_for_rxeq                                           = "rxvalid",
		parameter hssi_adapt_rx_rx_usertest_sel                                                   = "direct_tr_usertest3_sel",
		parameter hssi_adapt_rx_rxfifo_empty                                                      = "empty_default",
		parameter hssi_adapt_rx_rxfifo_full                                                       = "full_dw",
		parameter hssi_adapt_rx_rxfifo_mode                                                       = "rxphase_comp",
		parameter hssi_adapt_rx_rxfifo_pempty                                                     = 2,
		parameter hssi_adapt_rx_rxfifo_pfull                                                      = 5,
		parameter hssi_adapt_rx_rxfiford_post_ct_sel                                              = "rxfiford_sclk_post_ct",
		parameter hssi_adapt_rx_rxfiford_to_aib_sel                                               = "rxfiford_sclk_to_aib",
		parameter hssi_adapt_rx_rxfifowr_post_ct_sel                                              = "rxfifowr_sclk_post_ct",
		parameter hssi_adapt_rx_rxfifowr_pre_ct_sel                                               = "rxfifowr_sclk_pre_ct",
		parameter hssi_adapt_rx_hd_hssiadapt_speed_grade                                          = "dash_2",
		parameter hssi_adapt_rx_stretch_num_stages                                                = "seven_stage",
		parameter hssi_adapt_rx_sup_mode                                                          = "user_mode",
		parameter hssi_adapt_rx_txeq_clk_scg_en                                                   = "enable",
		parameter hssi_adapt_rx_txeq_clk_sel                                                      = "txeq_pld_pcs_rx_clk_out",
		parameter hssi_adapt_rx_txeq_mode                                                         = "eq_disable",
		parameter hssi_adapt_rx_txeq_rst_sel                                                      = "txeq_pcs_rx_pld_rst_n",
		parameter hssi_adapt_rx_txfiford_post_ct_sel                                              = "txfiford_sclk_post_ct",
		parameter hssi_adapt_rx_txfiford_pre_ct_sel                                               = "txfiford_sclk_pre_ct",
		parameter hssi_adapt_rx_txfifowr_from_aib_sel                                             = "txfifowr_sclk_from_aib",
		parameter hssi_adapt_rx_txfifowr_post_ct_sel                                              = "txfifowr_sclk_post_ct",
		parameter hssi_adapt_rx_us_bypass_pipeln                                                  = "us_bypass_pipeln_dis",
		parameter hssi_adapt_rx_word_align_enable                                                 = "enable",
		parameter hssi_adapt_rx_word_mark                                                         = "wm_en",
		parameter hssi_adapt_rx_silicon_rev                                                       = "14nm5cr2",
		parameter pma_reset_sequencer_rx_path_rstn_overrideb                                      = "use_sequencer",
		parameter pma_reset_sequencer_xrx_path_uc_cal_clk_bypass                                  = "cal_clk_0",
		parameter pma_reset_sequencer_xrx_path_uc_cal_enable                                      = "rx_cal_off",
		parameter pma_reset_sequencer_silicon_rev                                                 = "14nm5cr2",
		parameter pma_tx_ser_bti_protected                                                        = "false",
		parameter pma_tx_ser_control_clks_divtx_aibtx                                             = "no_dft_control_clkdivtx_clkaibtx",
		parameter pma_tx_ser_datarate_bps                                                         = "0",
		parameter pma_tx_ser_duty_cycle_correction_mode_ctrl                                      = "dcc_disable",
		parameter pma_tx_ser_initial_settings                                                     = "true",
		parameter pma_tx_ser_pcie_gen                                                             = "non_pcie",
		parameter pma_tx_ser_power_rail_er                                                        = 1120,
		parameter pma_tx_ser_powermode_ac_ser                                                     = "ac_clk_divtx_user_33_jitcomp1p1",
		parameter pma_tx_ser_powermode_dc_ser                                                     = "dc_clk_divtx_user_33_jitcomp1p1",
		parameter pma_tx_ser_prot_mode                                                            = "basic_tx",
		parameter pma_tx_ser_ser_clk_divtx_user_sel                                               = "divtx_user_33",
		parameter pma_tx_ser_ser_aibck_enable                                                     = "enable",
		parameter pma_tx_ser_ser_aibck_x1_override                                                = "normal",
		parameter pma_tx_ser_ser_clk_mon                                                          = "disable_clk_mon",
		parameter pma_tx_ser_ser_dftppm_clkselect                                                 = "aib_dftppm",
		parameter pma_tx_ser_ser_in_jitcomp                                                       = "jitcomp_on",
		parameter pma_tx_ser_ser_powerdown                                                        = "normal_poweron_ser",
		parameter pma_tx_ser_ser_preset_bti_en                                                    = "ser_preset_bti_disable",
		parameter pma_tx_ser_sup_mode                                                             = "user_mode",
		parameter pma_tx_ser_uc_vcc_setting                                                       = "vcc_setting2",
		parameter pma_tx_ser_silicon_rev                                                          = "14nm5cr2",
		parameter pma_rx_deser_bitslip_bypass                                                     = "bs_bypass_yes",
		parameter pma_rx_deser_bti_protected                                                      = "false",
		parameter pma_rx_deser_clkdiv_source                                                      = "vco_bypass_normal",
		parameter pma_rx_deser_clkdivrx_user_mode                                                 = "clkdivrx_user_div33",
		parameter pma_rx_deser_datarate_bps                                                       = "25781250000",
		parameter pma_rx_deser_deser_aib_dftppm_en                                                = "disable",
		parameter pma_rx_deser_deser_aibck_en                                                     = "enable",
		parameter pma_rx_deser_deser_aibck_x1                                                     = "normal",
		parameter pma_rx_deser_deser_factor                                                       = "deser_64b",
		parameter pma_rx_deser_deser_powerdown                                                    = "deser_power_up",
		parameter pma_rx_deser_force_adaptation_outputs                                           = "normal_outputs",
		parameter pma_rx_deser_force_clkdiv_for_testing                                           = "normal_clkdiv",
		parameter pma_rx_deser_odi_adapt_bti_en                                                   = "deser_bti_disable",
		parameter pma_rx_deser_optimal                                                            = "true",
		parameter pma_rx_deser_pcie_g3_hclk_en                                                    = "disable_hclk_div2",
		parameter pma_rx_deser_pm_cr2_tx_rx_pcie_gen                                              = "non_pcie",
		parameter pma_rx_deser_pm_cr2_tx_rx_pcie_gen_bitwidth                                     = "pcie_gen3_32b",
		parameter pma_rx_deser_powermode_ac_deser                                                 = "deser_ac_64b_nobs",
		parameter pma_rx_deser_powermode_ac_deser_bs                                              = "deser_ac_bs_off",
		parameter pma_rx_deser_powermode_dc_deser                                                 = "deser_dc_64b_nobs",
		parameter pma_rx_deser_powermode_dc_deser_bs                                              = "powerdown_deser_bs",
		parameter pma_rx_deser_prot_mode                                                          = "basic_rx",
		parameter pma_rx_deser_rst_n_adapt_odi                                                    = "no_rst_adapt_odi",
		parameter pma_rx_deser_sd_clk                                                             = "sd_clk_disabled",
		parameter pma_rx_deser_sup_mode                                                           = "user_mode",
		parameter pma_rx_deser_tdr_mode                                                           = "select_bbpd_data",
		parameter pma_rx_deser_silicon_rev                                                        = "14nm5cr2",
		parameter pma_txpath_chnsequencer_pcie_gen                                                = "non_pcie",
		parameter pma_txpath_chnsequencer_prot_mode                                               = "basic_tx",
		parameter pma_txpath_chnsequencer_sup_mode                                                = "sup_off",
		parameter pma_txpath_chnsequencer_txpath_chnseq_enable                                    = "disable",
		parameter pma_txpath_chnsequencer_txpath_chnseq_idle_direct_on                            = "cgb_idle_direct_off",
		parameter pma_txpath_chnsequencer_txpath_chnseq_stage_select                              = 0,
		parameter pma_txpath_chnsequencer_txpath_chnseq_wakeup_bypass                             = "bypass_off",
		parameter pma_txpath_chnsequencer_silicon_rev                                             = "14nm5bcr2ea",
		parameter hssi_aibcr_rx_aib_datasel_gr0                                                   = "aib_datasel0_setting0",
		parameter hssi_aibcr_rx_aib_datasel_gr1                                                   = "aib_datasel1_setting0",
		parameter hssi_aibcr_rx_aib_datasel_gr2                                                   = "aib_datasel2_setting1",
		parameter hssi_aibcr_rx_aib_ddrctrl_gr0                                                   = "aib_ddr0_setting1",
		parameter hssi_aibcr_rx_aib_ddrctrl_gr1                                                   = "aib_ddr1_setting1",
		parameter hssi_aibcr_rx_aib_iinasyncen                                                    = "aib_inasyncen_setting2",
		parameter hssi_aibcr_rx_aib_iinclken                                                      = "aib_inclken_setting3",
		parameter hssi_aibcr_rx_aib_outctrl_gr0                                                   = "aib_outen0_setting1",
		parameter hssi_aibcr_rx_aib_outctrl_gr1                                                   = "aib_outen1_setting1",
		parameter hssi_aibcr_rx_aib_outctrl_gr2                                                   = "aib_outen2_setting1",
		parameter hssi_aibcr_rx_aib_outctrl_gr3                                                   = "aib_outen3_setting1",
		parameter hssi_aibcr_rx_aib_outndrv_r12                                                   = "aib_ndrv12_setting1",
		parameter hssi_aibcr_rx_aib_outndrv_r56                                                   = "aib_ndrv56_setting1",
		parameter hssi_aibcr_rx_aib_outndrv_r78                                                   = "aib_ndrv78_setting1",
		parameter hssi_aibcr_rx_aib_outpdrv_r12                                                   = "aib_pdrv12_setting1",
		parameter hssi_aibcr_rx_aib_outpdrv_r56                                                   = "aib_pdrv56_setting1",
		parameter hssi_aibcr_rx_aib_outpdrv_r78                                                   = "aib_pdrv78_setting1",
		parameter hssi_aibcr_rx_aib_red_rx_shiften                                                = "aib_red_rx_shift_disable",
		parameter hssi_aibcr_rx_aib_rx_clkdiv                                                     = "aib_rx_clkdiv_setting1",
		parameter hssi_aibcr_rx_aib_rx_dcc_byp                                                    = "aib_rx_dcc_byp_disable",
		parameter hssi_aibcr_rx_aib_rx_dcc_byp_iocsr_unused                                       = "aib_rx_dcc_byp_disable_iocsr_unused",
		parameter hssi_aibcr_rx_aib_rx_dcc_cont_cal                                               = "aib_rx_dcc_cal_cont",
		parameter hssi_aibcr_rx_aib_rx_dcc_cont_cal_iocsr_unused                                  = "aib_rx_dcc_cal_single_iocsr_unused",
		parameter hssi_aibcr_rx_aib_rx_dcc_dft                                                    = "aib_rx_dcc_dft_disable",
		parameter hssi_aibcr_rx_aib_rx_dcc_dft_sel                                                = "aib_rx_dcc_dft_mode0",
		parameter hssi_aibcr_rx_aib_rx_dcc_dll_entest                                             = "aib_rx_dcc_dll_test_disable",
		parameter hssi_aibcr_rx_aib_rx_dcc_dy_ctl_static                                          = "aib_rx_dcc_dy_ctl_static_setting1",
		parameter hssi_aibcr_rx_aib_rx_dcc_dy_ctlsel                                              = "aib_rx_dcc_dy_ctlsel_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_en                                                     = "aib_rx_dcc_enable",
		parameter hssi_aibcr_rx_aib_rx_dcc_en_iocsr_unused                                        = "aib_rx_dcc_disable_iocsr_unused",
		parameter hssi_aibcr_rx_aib_rx_dcc_manual_dn                                              = "aib_rx_dcc_manual_dn0",
		parameter hssi_aibcr_rx_aib_rx_dcc_manual_up                                              = "aib_rx_dcc_manual_up0",
		parameter hssi_aibcr_rx_aib_rx_dcc_rst_prgmnvrt                                           = "aib_rx_dcc_st_rst_prgmnvrt_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_core_dn_prgmnvrt                                    = "aib_rx_dcc_st_core_dn_prgmnvrt_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_core_up_prgmnvrt                                    = "aib_rx_dcc_st_core_up_prgmnvrt_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_core_updnen                                         = "aib_rx_dcc_st_core_updnen_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_dftmuxsel                                           = "aib_rx_dcc_st_dftmuxsel_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_dly_pst                                             = "aib_rx_dcc_st_dly_pst_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_en                                                  = "aib_rx_dcc_st_en_setting1",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_lockreq_muxsel                                      = "aib_rx_dcc_st_lockreq_muxsel_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_new_dll                                             = "aib_rx_dcc_new_dll_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_new_dll2                                            = "aib_rx_dcc_new_dll2_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_st_rst                                                 = "aib_rx_dcc_st_rst_setting0",
		parameter hssi_aibcr_rx_aib_rx_dcc_test_clk_pll_en_n                                      = "aib_rx_dcc_test_clk_pll_en_n_disable",
		parameter hssi_aibcr_rx_aib_rx_halfcode                                                   = "aib_rx_halfcode_enable",
		parameter hssi_aibcr_rx_aib_rx_selflock                                                   = "aib_rx_selflock_enable",
		parameter hssi_aibcr_rx_dft_hssitestip_dll_dcc_en                                         = "disable_dft",
		parameter hssi_aibcr_rx_op_mode                                                           = "rx_dcc_enable",
		parameter hssi_aibcr_rx_powermode_ac                                                      = "rxdatapath_high_speed_pwr",
		parameter hssi_aibcr_rx_powermode_dc                                                      = "powerup",
		parameter hssi_aibcr_rx_redundancy_en                                                     = "disable",
		parameter hssi_aibcr_rx_sup_mode                                                          = "user_mode",
		parameter hssi_aibcr_rx_silicon_rev                                                       = "14nm5cr2",
		parameter hssi_aibcr_tx_aib_datasel_gr0                                                   = "aib_datasel0_setting0",
		parameter hssi_aibcr_tx_aib_datasel_gr1                                                   = "aib_datasel1_setting1",
		parameter hssi_aibcr_tx_aib_datasel_gr2                                                   = "aib_datasel2_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_clkdiv                                           = "aib_dllstr_align_clkdiv_setting1",
		parameter hssi_aibcr_tx_aib_dllstr_align_dcc_dll_dft_sel                                  = "aib_dllstr_align_dcc_dll_dft_sel_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_dft_ch_muxsel                                    = "aib_dllstr_align_dft_ch_muxsel_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_dly_pst                                          = "aib_dllstr_align_dly_pst_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_dy_ctl_static                                    = "aib_dllstr_align_dy_ctl_static_setting1",
		parameter hssi_aibcr_tx_aib_dllstr_align_dy_ctlsel                                        = "aib_dllstr_align_dy_ctlsel_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_entest                                           = "aib_dllstr_align_test_disable",
		parameter hssi_aibcr_tx_aib_dllstr_align_halfcode                                         = "aib_dllstr_align_halfcode_enable",
		parameter hssi_aibcr_tx_aib_dllstr_align_selflock                                         = "aib_dllstr_align_selflock_enable",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_core_dn_prgmnvrt                              = "aib_dllstr_align_st_core_dn_prgmnvrt_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_core_up_prgmnvrt                              = "aib_dllstr_align_st_core_up_prgmnvrt_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_core_updnen                                   = "aib_dllstr_align_st_core_updnen_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_dftmuxsel                                     = "aib_dllstr_align_st_dftmuxsel_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_en                                            = "aib_dllstr_align_st_en_setting1",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_lockreq_muxsel                                = "aib_dllstr_align_st_lockreq_muxsel_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_new_dll                                       = "aib_dllstr_align_new_dll_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_new_dll2                                      = "aib_dllstr_align_new_dll2_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_rst                                           = "aib_dllstr_align_st_rst_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_st_rst_prgmnvrt                                  = "aib_dllstr_align_st_rst_prgmnvrt_setting0",
		parameter hssi_aibcr_tx_aib_dllstr_align_test_clk_pll_en_n                                = "aib_dllstr_align_test_clk_pll_en_n_disable",
		parameter hssi_aibcr_tx_aib_inctrl_gr0                                                    = "aib_inctrl0_setting1",
		parameter hssi_aibcr_tx_aib_inctrl_gr1                                                    = "aib_inctrl1_setting3",
		parameter hssi_aibcr_tx_aib_inctrl_gr2                                                    = "aib_inctrl2_setting2",
		parameter hssi_aibcr_tx_aib_inctrl_gr3                                                    = "aib_inctrl3_setting2",
		parameter hssi_aibcr_tx_aib_outctrl_gr0                                                   = "aib_outen0_setting1",
		parameter hssi_aibcr_tx_aib_outctrl_gr1                                                   = "aib_outen1_setting1",
		parameter hssi_aibcr_tx_aib_outctrl_gr2                                                   = "aib_outen2_setting1",
		parameter hssi_aibcr_tx_aib_outndrv_r12                                                   = "aib_ndrv12_setting1",
		parameter hssi_aibcr_tx_aib_outndrv_r34                                                   = "aib_ndrv34_setting1",
		parameter hssi_aibcr_tx_aib_outndrv_r56                                                   = "aib_ndrv56_setting1",
		parameter hssi_aibcr_tx_aib_outndrv_r78                                                   = "aib_ndrv78_setting1",
		parameter hssi_aibcr_tx_aib_outpdrv_r12                                                   = "aib_pdrv12_setting1",
		parameter hssi_aibcr_tx_aib_outpdrv_r34                                                   = "aib_pdrv34_setting1",
		parameter hssi_aibcr_tx_aib_outpdrv_r56                                                   = "aib_pdrv56_setting1",
		parameter hssi_aibcr_tx_aib_outpdrv_r78                                                   = "aib_pdrv78_setting1",
		parameter hssi_aibcr_tx_aib_red_dirclkn_shiften                                           = "aib_red_dirclkn_shift_disable",
		parameter hssi_aibcr_tx_aib_red_dirclkp_shiften                                           = "aib_red_dirclkp_shift_disable",
		parameter hssi_aibcr_tx_aib_red_drx_shiften                                               = "aib_red_drx_shift_disable",
		parameter hssi_aibcr_tx_aib_red_dtx_shiften                                               = "aib_red_dtx_shift_disable",
		parameter hssi_aibcr_tx_aib_red_pinp_shiften                                              = "aib_red_pinp_shift_disable",
		parameter hssi_aibcr_tx_aib_red_rx_shiften                                                = "aib_red_rx_shift_disable",
		parameter hssi_aibcr_tx_aib_red_tx_shiften                                                = "aib_red_tx_shift_disable",
		parameter hssi_aibcr_tx_aib_red_txferclkout_shiften                                       = "aib_red_txferclkout_shift_disable",
		parameter hssi_aibcr_tx_aib_red_txferclkoutn_shiften                                      = "aib_red_txferclkoutn_shift_disable",
		parameter hssi_aibcr_tx_dfd_dll_dcc_en                                                    = "disable_dfd",
		parameter hssi_aibcr_tx_dft_hssitestip_dll_dcc_en                                         = "disable_dft",
		parameter hssi_aibcr_tx_op_mode                                                           = "tx_dll_enable",
		parameter hssi_aibcr_tx_powermode_ac                                                      = "txdatapath_high_speed_pwr",
		parameter hssi_aibcr_tx_powermode_dc                                                      = "powerup",
		parameter hssi_aibcr_tx_redundancy_en                                                     = "disable",
		parameter hssi_aibcr_tx_sup_mode                                                          = "user_mode",
		parameter hssi_aibcr_tx_silicon_rev                                                       = "14nm5cr2",
		parameter hssi_aibnd_rx_aib_datasel_gr0                                                   = "aib_datasel0_setting0",
		parameter hssi_aibnd_rx_aib_datasel_gr1                                                   = "aib_datasel1_setting1",
		parameter hssi_aibnd_rx_aib_datasel_gr2                                                   = "aib_datasel2_setting1",
		parameter hssi_aibnd_rx_aib_dllstr_align_clkdiv                                           = "aib_dllstr_align_clkdiv_setting1",
		parameter hssi_aibnd_rx_aib_dllstr_align_dly_pst                                          = "aib_dllstr_align_dly_pst_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_dy_ctl_static                                    = "aib_dllstr_align_dy_ctl_static_setting1",
		parameter hssi_aibnd_rx_aib_dllstr_align_dy_ctlsel                                        = "aib_dllstr_align_dy_ctlsel_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_entest                                           = "aib_dllstr_align_test_disable",
		parameter hssi_aibnd_rx_aib_dllstr_align_halfcode                                         = "aib_dllstr_align_halfcode_enable",
		parameter hssi_aibnd_rx_aib_dllstr_align_selflock                                         = "aib_dllstr_align_selflock_enable",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_core_dn_prgmnvrt                              = "aib_dllstr_align_st_core_dn_prgmnvrt_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_core_up_prgmnvrt                              = "aib_dllstr_align_st_core_up_prgmnvrt_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_core_updnen                                   = "aib_dllstr_align_st_core_updnen_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_dftmuxsel                                     = "aib_dllstr_align_st_dftmuxsel_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_en                                            = "aib_dllstr_align_st_en_setting1",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_hps_ctrl_en                                   = "aib_dllstr_align_hps_ctrl_en_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_lockreq_muxsel                                = "aib_dllstr_align_st_lockreq_muxsel_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_new_dll                                       = "aib_dllstr_align_new_dll_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_rst                                           = "aib_dllstr_align_st_rst_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_st_rst_prgmnvrt                                  = "aib_dllstr_align_st_rst_prgmnvrt_setting0",
		parameter hssi_aibnd_rx_aib_dllstr_align_test_clk_pll_en_n                                = "aib_dllstr_align_test_clk_pll_en_n_disable",
		parameter hssi_aibnd_rx_aib_inctrl_gr0                                                    = "aib_inctrl0_setting1",
		parameter hssi_aibnd_rx_aib_inctrl_gr1                                                    = "aib_inctrl1_setting3",
		parameter hssi_aibnd_rx_aib_inctrl_gr2                                                    = "aib_inctrl2_setting2",
		parameter hssi_aibnd_rx_aib_inctrl_gr3                                                    = "aib_inctrl3_setting3",
		parameter hssi_aibnd_rx_aib_outctrl_gr0                                                   = "aib_outen0_setting1",
		parameter hssi_aibnd_rx_aib_outctrl_gr1                                                   = "aib_outen1_setting1",
		parameter hssi_aibnd_rx_aib_outctrl_gr2                                                   = "aib_outen2_setting1",
		parameter hssi_aibnd_rx_aib_outndrv_r12                                                   = "aib_ndrv12_setting1",
		parameter hssi_aibnd_rx_aib_outndrv_r34                                                   = "aib_ndrv34_setting1",
		parameter hssi_aibnd_rx_aib_outndrv_r56                                                   = "aib_ndrv56_setting1",
		parameter hssi_aibnd_rx_aib_outndrv_r78                                                   = "aib_ndrv78_setting1",
		parameter hssi_aibnd_rx_aib_outpdrv_r12                                                   = "aib_pdrv12_setting1",
		parameter hssi_aibnd_rx_aib_outpdrv_r34                                                   = "aib_pdrv34_setting1",
		parameter hssi_aibnd_rx_aib_outpdrv_r56                                                   = "aib_pdrv56_setting1",
		parameter hssi_aibnd_rx_aib_outpdrv_r78                                                   = "aib_pdrv78_setting1",
		parameter hssi_aibnd_rx_aib_red_shift_en                                                  = "aib_red_shift_disable",
		parameter hssi_aibnd_rx_dft_hssitestip_dll_dcc_en                                         = "disable_dft",
		parameter hssi_aibnd_rx_op_mode                                                           = "rx_dll_enable",
		parameter hssi_aibnd_rx_powermode_ac                                                      = "rxdatapath_high_speed_pwr",
		parameter hssi_aibnd_rx_powermode_dc                                                      = "rxdatapath_powerup",
		parameter hssi_aibnd_rx_redundancy_en                                                     = "disable",
		parameter hssi_aibnd_rx_sup_mode                                                          = "user_mode",
		parameter hssi_aibnd_rx_silicon_rev                                                       = "14nm5cr2",
		parameter hssi_aibnd_tx_aib_datasel_gr0                                                   = "aib_datasel0_setting0",
		parameter hssi_aibnd_tx_aib_datasel_gr1                                                   = "aib_datasel1_setting0",
		parameter hssi_aibnd_tx_aib_datasel_gr2                                                   = "aib_datasel2_setting1",
		parameter hssi_aibnd_tx_aib_datasel_gr3                                                   = "aib_datasel3_setting1",
		parameter hssi_aibnd_tx_aib_ddrctrl_gr0                                                   = "aib_ddr0_setting1",
		parameter hssi_aibnd_tx_aib_iinasyncen                                                    = "aib_inasyncen_setting2",
		parameter hssi_aibnd_tx_aib_iinclken                                                      = "aib_inclken_setting3",
		parameter hssi_aibnd_tx_aib_outctrl_gr0                                                   = "aib_outen0_setting1",
		parameter hssi_aibnd_tx_aib_outctrl_gr1                                                   = "aib_outen1_setting1",
		parameter hssi_aibnd_tx_aib_outctrl_gr2                                                   = "aib_outen2_setting1",
		parameter hssi_aibnd_tx_aib_outctrl_gr3                                                   = "aib_outen3_setting1",
		parameter hssi_aibnd_tx_aib_outndrv_r34                                                   = "aib_ndrv34_setting1",
		parameter hssi_aibnd_tx_aib_outndrv_r56                                                   = "aib_ndrv56_setting1",
		parameter hssi_aibnd_tx_aib_outpdrv_r34                                                   = "aib_pdrv34_setting1",
		parameter hssi_aibnd_tx_aib_outpdrv_r56                                                   = "aib_pdrv56_setting1",
		parameter hssi_aibnd_tx_aib_red_dirclkn_shiften                                           = "aib_red_dirclkn_shift_disable",
		parameter hssi_aibnd_tx_aib_red_dirclkp_shiften                                           = "aib_red_dirclkp_shift_disable",
		parameter hssi_aibnd_tx_aib_red_drx_shiften                                               = "aib_red_drx_shift_disable",
		parameter hssi_aibnd_tx_aib_red_dtx_shiften                                               = "aib_red_dtx_shift_disable",
		parameter hssi_aibnd_tx_aib_red_pout_shiften                                              = "aib_red_pout_shift_disable",
		parameter hssi_aibnd_tx_aib_red_rx_shiften                                                = "aib_red_rx_shift_disable",
		parameter hssi_aibnd_tx_aib_red_tx_shiften                                                = "aib_red_tx_shift_disable",
		parameter hssi_aibnd_tx_aib_red_txferclkout_shiften                                       = "aib_red_txferclkout_shift_disable",
		parameter hssi_aibnd_tx_aib_red_txferclkoutn_shiften                                      = "aib_red_txferclkoutn_shift_disable",
		parameter hssi_aibnd_tx_aib_tx_clkdiv                                                     = "aib_tx_clkdiv_setting1",
		parameter hssi_aibnd_tx_aib_tx_dcc_byp                                                    = "aib_tx_dcc_byp_disable",
		parameter hssi_aibnd_tx_aib_tx_dcc_byp_iocsr_unused                                       = "aib_tx_dcc_byp_disable_iocsr_unused",
		parameter hssi_aibnd_tx_aib_tx_dcc_cont_cal                                               = "aib_tx_dcc_cal_cont",
		parameter hssi_aibnd_tx_aib_tx_dcc_cont_cal_iocsr_unused                                  = "aib_tx_dcc_cal_single_iocsr_unused",
		parameter hssi_aibnd_tx_aib_tx_dcc_dft                                                    = "aib_tx_dcc_dft_disable",
		parameter hssi_aibnd_tx_aib_tx_dcc_dft_sel                                                = "aib_tx_dcc_dft_mode0",
		parameter hssi_aibnd_tx_aib_tx_dcc_dll_dft_sel                                            = "aib_tx_dcc_dll_dft_sel_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_dll_entest                                             = "aib_tx_dcc_dll_test_disable",
		parameter hssi_aibnd_tx_aib_tx_dcc_dy_ctl_static                                          = "aib_tx_dcc_dy_ctl_static_setting1",
		parameter hssi_aibnd_tx_aib_tx_dcc_dy_ctlsel                                              = "aib_tx_dcc_dy_ctlsel_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_en                                                     = "aib_tx_dcc_enable",
		parameter hssi_aibnd_tx_aib_tx_dcc_en_iocsr_unused                                        = "aib_tx_dcc_disable_iocsr_unused",
		parameter hssi_aibnd_tx_aib_tx_dcc_manual_dn                                              = "aib_tx_dcc_manual_dn0",
		parameter hssi_aibnd_tx_aib_tx_dcc_manual_up                                              = "aib_tx_dcc_manual_up0",
		parameter hssi_aibnd_tx_aib_tx_dcc_rst_prgmnvrt                                           = "aib_tx_dcc_st_rst_prgmnvrt_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_core_dn_prgmnvrt                                    = "aib_tx_dcc_st_core_dn_prgmnvrt_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_core_up_prgmnvrt                                    = "aib_tx_dcc_st_core_up_prgmnvrt_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_core_updnen                                         = "aib_tx_dcc_st_core_updnen_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_dftmuxsel                                           = "aib_tx_dcc_st_dftmuxsel_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_dly_pst                                             = "aib_tx_dcc_st_dly_pst_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_en                                                  = "aib_tx_dcc_st_en_setting1",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_hps_ctrl_en                                         = "aib_tx_dcc_hps_ctrl_en_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_lockreq_muxsel                                      = "aib_tx_dcc_st_lockreq_muxsel_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_new_dll                                             = "aib_tx_dcc_new_dll_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_st_rst                                                 = "aib_tx_dcc_st_rst_setting0",
		parameter hssi_aibnd_tx_aib_tx_dcc_test_clk_pll_en_n                                      = "aib_tx_dcc_test_clk_pll_en_n_disable",
		parameter hssi_aibnd_tx_aib_tx_halfcode                                                   = "aib_tx_halfcode_enable",
		parameter hssi_aibnd_tx_aib_tx_selflock                                                   = "aib_tx_selflock_enable",
		parameter hssi_aibnd_tx_dfd_dll_dcc_en                                                    = "disable_dfd",
		parameter hssi_aibnd_tx_dft_hssitestip_dll_dcc_en                                         = "disable_dft",
		parameter hssi_aibnd_tx_op_mode                                                           = "tx_dcc_enable",
		parameter hssi_aibnd_tx_powermode_ac                                                      = "txdatapath_high_speed_pwr",
		parameter hssi_aibnd_tx_powermode_dc                                                      = "txdatapath_powerup",
		parameter hssi_aibnd_tx_redundancy_en                                                     = "disable",
		parameter hssi_aibnd_tx_sup_mode                                                          = "user_mode",
		parameter hssi_aibnd_tx_silicon_rev                                                       = "14nm5cr2",
		parameter hssi_pipe_gen3_bypass_rx_detection_enable                                       = "false",
		parameter hssi_pipe_gen3_bypass_rx_preset                                                 = 0,
		parameter hssi_pipe_gen3_bypass_rx_preset_enable                                          = "false",
		parameter hssi_pipe_gen3_bypass_tx_coefficent                                             = 0,
		parameter hssi_pipe_gen3_bypass_tx_coefficent_enable                                      = "false",
		parameter hssi_pipe_gen3_elecidle_delay_g3                                                = 0,
		parameter hssi_pipe_gen3_ind_error_reporting                                              = "dis_ind_error_reporting",
		parameter hssi_pipe_gen3_mode                                                             = "disable_pcs",
		parameter hssi_pipe_gen3_phy_status_delay_g12                                             = 0,
		parameter hssi_pipe_gen3_phy_status_delay_g3                                              = 0,
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g12                                         = "dis_phystatus_rst_toggle",
		parameter hssi_pipe_gen3_phystatus_rst_toggle_g3                                          = "dis_phystatus_rst_toggle_g3",
		parameter hssi_pipe_gen3_rate_match_pad_insertion                                         = "dis_rm_fifo_pad_ins",
		parameter hssi_pipe_gen3_sup_mode                                                         = "user_mode",
		parameter hssi_pipe_gen3_test_out_sel                                                     = "disable_test_out",
		parameter hssi_pipe_gen3_silicon_rev                                                      = "14nm5cr2",
		parameter hssi_gen3_rx_pcs_block_sync                                                     = "bypass_block_sync",
		parameter hssi_gen3_rx_pcs_block_sync_sm                                                  = "disable_blk_sync_sm",
		parameter hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn                                          = "disable",
		parameter hssi_gen3_rx_pcs_lpbk_force                                                     = "lpbk_frce_dis",
		parameter hssi_gen3_rx_pcs_mode                                                           = "disable_pcs",
		parameter hssi_gen3_rx_pcs_rate_match_fifo                                                = "bypass_rm_fifo",
		parameter hssi_gen3_rx_pcs_rate_match_fifo_latency                                        = "low_latency",
		parameter hssi_gen3_rx_pcs_reverse_lpbk                                                   = "rev_lpbk_dis",
		parameter hssi_gen3_rx_pcs_rx_b4gb_par_lpbk                                               = "b4gb_par_lpbk_dis",
		parameter hssi_gen3_rx_pcs_rx_force_balign                                                = "dis_force_balign",
		parameter hssi_gen3_rx_pcs_rx_ins_del_one_skip                                            = "ins_del_one_skip_dis",
		parameter hssi_gen3_rx_pcs_rx_num_fixed_pat                                               = 0,
		parameter hssi_gen3_rx_pcs_rx_test_out_sel                                                = "rx_test_out0",
		parameter hssi_gen3_rx_pcs_sup_mode                                                       = "user_mode",
		parameter hssi_gen3_rx_pcs_silicon_rev                                                    = "14nm5cr2",
		parameter hssi_gen3_tx_pcs_mode                                                           = "disable_pcs",
		parameter hssi_gen3_tx_pcs_reverse_lpbk                                                   = "rev_lpbk_dis",
		parameter hssi_gen3_tx_pcs_sup_mode                                                       = "user_mode",
		parameter hssi_gen3_tx_pcs_tx_bitslip                                                     = 0,
		parameter hssi_gen3_tx_pcs_tx_gbox_byp                                                    = "bypass_gbox",
		parameter hssi_gen3_tx_pcs_silicon_rev                                                    = "14nm5cr2",
		parameter hssi_adapt_tx_aib_clk_sel                                                       = "aib_clk_pma_aib_tx_clk",
		parameter hssi_adapt_tx_hd_hssiadapt_aib_hssi_pld_sclk_hz                                 = 0,
		parameter hssi_adapt_tx_hd_hssiadapt_aib_hssi_tx_transfer_clk_hz                          = 805664062,
		parameter hssi_adapt_tx_bonding_dft_en                                                    = "dft_dis",
		parameter hssi_adapt_tx_bonding_dft_val                                                   = "dft_0",
		parameter hssi_adapt_tx_chnl_bonding                                                      = "disable",
		parameter hssi_adapt_tx_hd_hssiadapt_csr_clk_hz                                           = 0,
		parameter hssi_adapt_tx_ctrl_plane_bonding                                                = "individual",
		parameter hssi_adapt_tx_datapath_mapping_mode                                             = "map_10g_2x2x_2x1x_fifo",
		parameter hssi_adapt_tx_ds_bypass_pipeln                                                  = "ds_bypass_pipeln_dis",
		parameter hssi_adapt_tx_duplex_mode                                                       = "enable",
		parameter hssi_adapt_tx_dv_gating                                                         = "disable",
		parameter hssi_adapt_tx_dyn_clk_sw_en                                                     = "disable",
		parameter hssi_adapt_tx_fifo_double_read                                                  = "fifo_double_read_en",
		parameter hssi_adapt_tx_fifo_mode                                                         = "phase_comp",
		parameter hssi_adapt_tx_fifo_rd_clk_scg_en                                                = "disable",
		parameter hssi_adapt_tx_fifo_rd_clk_sel                                                   = "fifo_rd_pld_pcs_tx_clk_out",
		parameter hssi_adapt_tx_fifo_ready_bypass                                                 = "disable",
		parameter hssi_adapt_tx_fifo_stop_rd                                                      = "rd_empty",
		parameter hssi_adapt_tx_fifo_stop_wr                                                      = "wr_full",
		parameter hssi_adapt_tx_fifo_width                                                        = "fifo_double_width",
		parameter hssi_adapt_tx_fifo_wr_clk_scg_en                                                = "disable",
		parameter hssi_adapt_tx_free_run_div_clk                                                  = "out_of_reset_sync",
		parameter hssi_adapt_tx_fsr_hip_fsr_in_bit0_rst_val                                       = "reset_to_one_hfsrin0",
		parameter hssi_adapt_tx_fsr_hip_fsr_in_bit1_rst_val                                       = "reset_to_one_hfsrin1",
		parameter hssi_adapt_tx_fsr_hip_fsr_in_bit2_rst_val                                       = "reset_to_one_hfsrin2",
		parameter hssi_adapt_tx_fsr_hip_fsr_in_bit3_rst_val                                       = "reset_to_zero_hfsrin3",
		parameter hssi_adapt_tx_fsr_hip_fsr_out_bit0_rst_val                                      = "reset_to_one_hfsrout0",
		parameter hssi_adapt_tx_fsr_hip_fsr_out_bit1_rst_val                                      = "reset_to_one_hfsrout1",
		parameter hssi_adapt_tx_fsr_hip_fsr_out_bit2_rst_val                                      = "reset_to_zero_hfsrout2",
		parameter hssi_adapt_tx_fsr_hip_fsr_out_bit3_rst_val                                      = "reset_to_zero_hfsrout3",
		parameter hssi_adapt_tx_fsr_mask_tx_pll_rst_val                                           = "reset_to_zero_maskpll",
		parameter hssi_adapt_tx_fsr_pld_txelecidle_rst_val                                        = "reset_to_zero_txelec",
		parameter hssi_adapt_tx_hd_hssiadapt_hip_aib_clk_2x_hz                                    = 0,
		parameter hssi_adapt_tx_hd_hssiadapt_hip_aib_clk_hz                                       = 0,
		parameter hssi_adapt_tx_hd_hssiadapt_hip_aib_txeq_clk_out_hz                              = 0,
		parameter hssi_adapt_tx_hip_mode                                                          = "disable_hip",
		parameter hssi_adapt_tx_hip_osc_clk_scg_en                                                = "enable",
		parameter hssi_adapt_tx_hrdrst_align_bypass                                               = "enable",
		parameter hssi_adapt_tx_hrdrst_dcd_cal_done_bypass                                        = "disable",
		parameter hssi_adapt_tx_hrdrst_dll_lock_bypass                                            = "disable",
		parameter hssi_adapt_tx_hrdrst_rx_osc_clk_scg_en                                          = "disable",
		parameter hssi_adapt_tx_hrdrst_user_ctl_en                                                = "disable",
		parameter hssi_adapt_tx_indv                                                              = "indv_en",
		parameter hssi_adapt_tx_loopback_mode                                                     = "loopback_disable",
		parameter hssi_adapt_tx_osc_clk_scg_en                                                    = "disable",
		parameter hssi_adapt_tx_phcomp_rd_del                                                     = "phcomp_rd_del2",
		parameter hssi_adapt_tx_pipe_mode                                                         = "disable_pipe",
		parameter hssi_adapt_tx_hd_hssiadapt_pld_pcs_tx_clk_out_hz                                = 402832031,
		parameter hssi_adapt_tx_hd_hssiadapt_pld_pma_hclk_hz                                      = 0,
		parameter hssi_adapt_tx_pma_aib_tx_clk_expected_setting                                   = "x2",
		parameter hssi_adapt_tx_hd_hssiadapt_pma_aib_tx_clk_hz                                    = 0,
		parameter hssi_adapt_tx_powerdown_mode                                                    = "powerup",
		parameter hssi_adapt_tx_presethint_bypass                                                 = "enable",
		parameter hssi_adapt_tx_qpi_sr_enable                                                     = "enable",
		parameter hssi_adapt_tx_rxqpi_pullup_rst_val                                              = "reset_to_zero_rxqpi",
		parameter hssi_adapt_tx_hd_hssiadapt_speed_grade                                          = "dash_2",
		parameter hssi_adapt_tx_stretch_num_stages                                                = "seven_stage",
		parameter hssi_adapt_tx_sup_mode                                                          = "user_mode",
		parameter hssi_adapt_tx_tx_datapath_tb_sel                                                = "cp_bond",
		parameter hssi_adapt_tx_tx_fastbond_wren                                                  = "wren_ds_del2_us_del2",
		parameter hssi_adapt_tx_tx_fifo_power_mode                                                = "full_width_full_depth",
		parameter hssi_adapt_tx_tx_fifo_read_latency_adjust                                       = "disable",
		parameter hssi_adapt_tx_tx_fifo_write_latency_adjust                                      = "disable",
		parameter hssi_adapt_tx_tx_osc_clock_setting                                              = "osc_clk_div_by1",
		parameter hssi_adapt_tx_tx_qpi_mode_en                                                    = "disable",
		parameter hssi_adapt_tx_tx_rev_lpbk                                                       = "disable",
		parameter hssi_adapt_tx_tx_usertest_sel                                                   = "enable",
		parameter hssi_adapt_tx_txfifo_empty                                                      = "empty_default",
		parameter hssi_adapt_tx_txfifo_full                                                       = "full_dw",
		parameter hssi_adapt_tx_txfifo_mode                                                       = "txphase_comp",
		parameter hssi_adapt_tx_txfifo_pempty                                                     = 2,
		parameter hssi_adapt_tx_txfifo_pfull                                                      = 5,
		parameter hssi_adapt_tx_txqpi_pulldn_rst_val                                              = "reset_to_zero_txqpid",
		parameter hssi_adapt_tx_txqpi_pullup_rst_val                                              = "reset_to_zero_txqpiu",
		parameter hssi_adapt_tx_word_align                                                        = "wa_en",
		parameter hssi_adapt_tx_word_align_enable                                                 = "enable",
		parameter hssi_adapt_tx_silicon_rev                                                       = "14nm5cr2",
		parameter hssi_krfec_rx_pcs_blksync_cor_en                                                = "detect",
		parameter hssi_krfec_rx_pcs_bypass_gb                                                     = "bypass_dis",
		parameter hssi_krfec_rx_pcs_clr_ctrl                                                      = "both_enabled",
		parameter hssi_krfec_rx_pcs_ctrl_bit_reverse                                              = "ctrl_bit_reverse_en",
		parameter hssi_krfec_rx_pcs_data_bit_reverse                                              = "data_bit_reverse_dis",
		parameter hssi_krfec_rx_pcs_dv_start                                                      = "with_blklock",
		parameter hssi_krfec_rx_pcs_err_mark_type                                                 = "err_mark_10g",
		parameter hssi_krfec_rx_pcs_error_marking_en                                              = "err_mark_dis",
		parameter hssi_krfec_rx_pcs_low_latency_en                                                = "disable",
		parameter hssi_krfec_rx_pcs_lpbk_mode                                                     = "lpbk_dis",
		parameter hssi_krfec_rx_pcs_parity_invalid_enum                                           = 8,
		parameter hssi_krfec_rx_pcs_parity_valid_num                                              = 4,
		parameter hssi_krfec_rx_pcs_pipeln_blksync                                                = "enable",
		parameter hssi_krfec_rx_pcs_pipeln_descrm                                                 = "disable",
		parameter hssi_krfec_rx_pcs_pipeln_errcorrect                                             = "disable",
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_ind                                            = "enable",
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_lfsr                                           = "disable",
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_loc                                            = "disable",
		parameter hssi_krfec_rx_pcs_pipeln_errtrap_pat                                            = "disable",
		parameter hssi_krfec_rx_pcs_pipeln_gearbox                                                = "enable",
		parameter hssi_krfec_rx_pcs_pipeln_syndrm                                                 = "enable",
		parameter hssi_krfec_rx_pcs_pipeln_trans_dec                                              = "disable",
		parameter hssi_krfec_rx_pcs_prot_mode                                                     = "disable_mode",
		parameter hssi_krfec_rx_pcs_receive_order                                                 = "receive_lsb",
		parameter hssi_krfec_rx_pcs_rx_testbus_sel                                                = "overall",
		parameter hssi_krfec_rx_pcs_signal_ok_en                                                  = "sig_ok_en",
		parameter hssi_krfec_rx_pcs_sup_mode                                                      = "user_mode",
		parameter hssi_krfec_rx_pcs_silicon_rev                                                   = "14nm5cr2",
		parameter hssi_krfec_tx_pcs_burst_err                                                     = "burst_err_dis",
		parameter hssi_krfec_tx_pcs_burst_err_len                                                 = "burst_err_len1",
		parameter hssi_krfec_tx_pcs_ctrl_bit_reverse                                              = "ctrl_bit_reverse_en",
		parameter hssi_krfec_tx_pcs_data_bit_reverse                                              = "data_bit_reverse_dis",
		parameter hssi_krfec_tx_pcs_enc_frame_query                                               = "enc_query_dis",
		parameter hssi_krfec_tx_pcs_low_latency_en                                                = "disable",
		parameter hssi_krfec_tx_pcs_pipeln_encoder                                                = "enable",
		parameter hssi_krfec_tx_pcs_pipeln_scrambler                                              = "enable",
		parameter hssi_krfec_tx_pcs_prot_mode                                                     = "disable_mode",
		parameter hssi_krfec_tx_pcs_sup_mode                                                      = "user_mode",
		parameter hssi_krfec_tx_pcs_transcode_err                                                 = "trans_err_dis",
		parameter hssi_krfec_tx_pcs_transmit_order                                                = "transmit_lsb",
		parameter hssi_krfec_tx_pcs_tx_testbus_sel                                                = "overall",
		parameter hssi_krfec_tx_pcs_silicon_rev                                                   = "14nm5cr2",
		parameter hssi_pipe_gen1_2_elec_idle_delay_val                                            = 0,
		parameter hssi_pipe_gen1_2_error_replace_pad                                              = "replace_edb",
		parameter hssi_pipe_gen1_2_hip_mode                                                       = "dis_hip",
		parameter hssi_pipe_gen1_2_ind_error_reporting                                            = "dis_ind_error_reporting",
		parameter hssi_pipe_gen1_2_phystatus_delay_val                                            = 0,
		parameter hssi_pipe_gen1_2_phystatus_rst_toggle                                           = "dis_phystatus_rst_toggle",
		parameter hssi_pipe_gen1_2_pipe_byte_de_serializer_en                                     = "dont_care_bds",
		parameter hssi_pipe_gen1_2_prot_mode                                                      = "disabled_prot_mode",
		parameter hssi_pipe_gen1_2_rpre_emph_a_val                                                = 0,
		parameter hssi_pipe_gen1_2_rpre_emph_b_val                                                = 0,
		parameter hssi_pipe_gen1_2_rpre_emph_c_val                                                = 0,
		parameter hssi_pipe_gen1_2_rpre_emph_d_val                                                = 0,
		parameter hssi_pipe_gen1_2_rpre_emph_e_val                                                = 0,
		parameter hssi_pipe_gen1_2_rvod_sel_a_val                                                 = 0,
		parameter hssi_pipe_gen1_2_rvod_sel_b_val                                                 = 0,
		parameter hssi_pipe_gen1_2_rvod_sel_c_val                                                 = 0,
		parameter hssi_pipe_gen1_2_rvod_sel_d_val                                                 = 0,
		parameter hssi_pipe_gen1_2_rvod_sel_e_val                                                 = 0,
		parameter hssi_pipe_gen1_2_rx_pipe_enable                                                 = "dis_pipe_rx",
		parameter hssi_pipe_gen1_2_rxdetect_bypass                                                = "dis_rxdetect_bypass",
		parameter hssi_pipe_gen1_2_sup_mode                                                       = "user_mode",
		parameter hssi_pipe_gen1_2_tx_pipe_enable                                                 = "dis_pipe_tx",
		parameter hssi_pipe_gen1_2_txswing                                                        = "dis_txswing",
		parameter hssi_pipe_gen1_2_silicon_rev                                                    = "14nm5cr2",
		parameter hssi_common_pld_pcs_interface_dft_clk_out_en                                    = "dft_clk_out_disable",
		parameter hssi_common_pld_pcs_interface_dft_clk_out_sel                                   = "teng_rx_dft_clk",
		parameter hssi_common_pld_pcs_interface_hrdrstctrl_en                                     = "hrst_dis",
		parameter hssi_common_pld_pcs_interface_pcs_testbus_block_sel                             = "pma_if",
		parameter hssi_common_pld_pcs_interface_silicon_rev                                       = "14nm5cr2",
		parameter hssi_common_pcs_pma_interface_asn_clk_enable                                    = "false",
		parameter hssi_common_pcs_pma_interface_asn_enable                                        = "dis_asn",
		parameter hssi_common_pcs_pma_interface_block_sel                                         = "eight_g_pcs",
		parameter hssi_common_pcs_pma_interface_bypass_early_eios                                 = "true",
		parameter hssi_common_pcs_pma_interface_bypass_pcie_switch                                = "true",
		parameter hssi_common_pcs_pma_interface_bypass_pma_ltr                                    = "true",
		parameter hssi_common_pcs_pma_interface_bypass_ppm_lock                                   = "false",
		parameter hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp                            = "true",
		parameter hssi_common_pcs_pma_interface_bypass_txdetectrx                                 = "true",
		parameter hssi_common_pcs_pma_interface_cdr_control                                       = "dis_cdr_ctrl",
		parameter hssi_common_pcs_pma_interface_cid_enable                                        = "dis_cid_mode",
		parameter hssi_common_pcs_pma_interface_data_mask_count                                   = 0,
		parameter hssi_common_pcs_pma_interface_data_mask_count_multi                             = 0,
		parameter hssi_common_pcs_pma_interface_dft_observation_clock_selection                   = "dft_clk_obsrv_tx0",
		parameter hssi_common_pcs_pma_interface_early_eios_counter                                = 0,
		parameter hssi_common_pcs_pma_interface_force_freqdet                                     = "force_freqdet_dis",
		parameter hssi_common_pcs_pma_interface_free_run_clk_enable                               = "false",
		parameter hssi_common_pcs_pma_interface_ignore_sigdet_g23                                 = "false",
		parameter hssi_common_pcs_pma_interface_pc_en_counter                                     = 0,
		parameter hssi_common_pcs_pma_interface_pc_rst_counter                                    = 0,
		parameter hssi_common_pcs_pma_interface_pcie_hip_mode                                     = "hip_disable",
		parameter hssi_common_pcs_pma_interface_ph_fifo_reg_mode                                  = "phfifo_reg_mode_dis",
		parameter hssi_common_pcs_pma_interface_phfifo_flush_wait                                 = 0,
		parameter hssi_common_pcs_pma_interface_pipe_if_g3pcs                                     = "pipe_if_8gpcs",
		parameter hssi_common_pcs_pma_interface_pma_done_counter                                  = 0,
		parameter hssi_common_pcs_pma_interface_pma_if_dft_en                                     = "dft_dis",
		parameter hssi_common_pcs_pma_interface_pma_if_dft_val                                    = "dft_0",
		parameter hssi_common_pcs_pma_interface_ppm_cnt_rst                                       = "ppm_cnt_rst_dis",
		parameter hssi_common_pcs_pma_interface_ppm_deassert_early                                = "deassert_early_dis",
		parameter hssi_common_pcs_pma_interface_ppm_det_buckets                                   = "ppm_300_100_bucket",
		parameter hssi_common_pcs_pma_interface_ppm_gen1_2_cnt                                    = "cnt_32k",
		parameter hssi_common_pcs_pma_interface_ppm_post_eidle_delay                              = "cnt_200_cycles",
		parameter hssi_common_pcs_pma_interface_ppmsel                                            = "ppmsel_1000",
		parameter hssi_common_pcs_pma_interface_prot_mode                                         = "other_protocols",
		parameter hssi_common_pcs_pma_interface_rxvalid_mask                                      = "rxvalid_mask_dis",
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter                               = 0,
		parameter hssi_common_pcs_pma_interface_sigdet_wait_counter_multi                         = 0,
		parameter hssi_common_pcs_pma_interface_sim_mode                                          = "disable",
		parameter hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en                           = "false",
		parameter hssi_common_pcs_pma_interface_sup_mode                                          = "user_mode",
		parameter hssi_common_pcs_pma_interface_testout_sel                                       = "ppm_det_test",
		parameter hssi_common_pcs_pma_interface_wait_clk_on_off_timer                             = 0,
		parameter hssi_common_pcs_pma_interface_wait_pipe_synchronizing                           = 0,
		parameter hssi_common_pcs_pma_interface_wait_send_syncp_fbkp                              = 0,
		parameter hssi_common_pcs_pma_interface_silicon_rev                                       = "14nm5cr2",
		parameter hssi_rx_pcs_pma_interface_block_sel                                             = "ten_g_pcs",
		parameter hssi_rx_pcs_pma_interface_channel_operation_mode                                = "tx_rx_pair_enabled",
		parameter hssi_rx_pcs_pma_interface_clkslip_sel                                           = "pld",
		parameter hssi_rx_pcs_pma_interface_lpbk_en                                               = "disable",
		parameter hssi_rx_pcs_pma_interface_master_clk_sel                                        = "master_rx_pma_clk",
		parameter hssi_rx_pcs_pma_interface_pldif_datawidth_mode                                  = "pldif_data_10bit",
		parameter hssi_rx_pcs_pma_interface_pma_dw_rx                                             = "pma_64b_rx",
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_en                                         = "dft_dis",
		parameter hssi_rx_pcs_pma_interface_pma_if_dft_val                                        = "dft_0",
		parameter hssi_rx_pcs_pma_interface_prbs9_dwidth                                          = "prbs9_64b",
		parameter hssi_rx_pcs_pma_interface_prbs_clken                                            = "prbs_clk_dis",
		parameter hssi_rx_pcs_pma_interface_prbs_ver                                              = "prbs_off",
		parameter hssi_rx_pcs_pma_interface_prot_mode_rx                                          = "teng_basic_mode_rx",
		parameter hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion                             = "rx_dyn_polinv_dis",
		parameter hssi_rx_pcs_pma_interface_rx_lpbk_en                                            = "lpbk_dis",
		parameter hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok                               = "force_sig_ok",
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mask                                          = "prbsmask128",
		parameter hssi_rx_pcs_pma_interface_rx_prbs_mode                                          = "teng_mode",
		parameter hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel                             = "sel_sig_det",
		parameter hssi_rx_pcs_pma_interface_rx_static_polarity_inversion                          = "rx_stat_polinv_dis",
		parameter hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en                                      = "uhsif_lpbk_dis",
		parameter hssi_rx_pcs_pma_interface_sup_mode                                              = "user_mode",
		parameter hssi_rx_pcs_pma_interface_silicon_rev                                           = "14nm5cr2",
		parameter hssi_tx_pcs_pma_interface_bypass_pma_txelecidle                                 = "true",
		parameter hssi_tx_pcs_pma_interface_channel_operation_mode                                = "tx_rx_pair_enabled",
		parameter hssi_tx_pcs_pma_interface_lpbk_en                                               = "disable",
		parameter hssi_tx_pcs_pma_interface_master_clk_sel                                        = "master_tx_pma_clk",
		parameter hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx                                 = "other_prot_mode",
		parameter hssi_tx_pcs_pma_interface_pldif_datawidth_mode                                  = "pldif_data_10bit",
		parameter hssi_tx_pcs_pma_interface_pma_dw_tx                                             = "pma_64b_tx",
		parameter hssi_tx_pcs_pma_interface_pma_if_dft_en                                         = "dft_dis",
		parameter hssi_tx_pcs_pma_interface_pmagate_en                                            = "pmagate_dis",
		parameter hssi_tx_pcs_pma_interface_prbs9_dwidth                                          = "prbs9_64b",
		parameter hssi_tx_pcs_pma_interface_prbs_clken                                            = "prbs_clk_dis",
		parameter hssi_tx_pcs_pma_interface_prbs_gen_pat                                          = "prbs_gen_dis",
		parameter hssi_tx_pcs_pma_interface_prot_mode_tx                                          = "teng_basic_mode_tx",
		parameter hssi_tx_pcs_pma_interface_sq_wave_num                                           = "sq_wave_default",
		parameter hssi_tx_pcs_pma_interface_sqwgen_clken                                          = "sqwgen_clk_dis",
		parameter hssi_tx_pcs_pma_interface_sup_mode                                              = "user_mode",
		parameter hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion                             = "tx_dyn_polinv_dis",
		parameter hssi_tx_pcs_pma_interface_tx_pma_data_sel                                       = "ten_g_pcs",
		parameter hssi_tx_pcs_pma_interface_tx_static_polarity_inversion                          = "tx_stat_polinv_dis",
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock                       = "uhsif_filt_stepsz_b4lock_2",
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value                = 0,
		parameter hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock                     = "uhsif_filt_cntthr_b4lock_8",
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period                          = "uhsif_dcn_test_period_4",
		parameter hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable                             = "uhsif_dcn_test_mode_disable",
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh                          = "uhsif_dzt_cnt_thr_2",
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable                      = "uhsif_dzt_disable",
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window                          = "uhsif_dzt_obr_win_16",
		parameter hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size                             = "uhsif_dzt_skipsz_4",
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel                            = "uhsif_index_cram",
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin                               = "uhsif_dcn_margin_2",
		parameter hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value                   = 0,
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control                           = "uhsif_dft_dz_det_val_0",
		parameter hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control                             = "uhsif_dft_up_val_0",
		parameter hssi_tx_pcs_pma_interface_uhsif_enable                                          = "uhsif_disable",
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock                       = "uhsif_lkd_segsz_aflock_512",
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock                      = "uhsif_lkd_segsz_b4lock_16",
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value            = 0,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value           = 0,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value           = 0,
		parameter hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value          = 0,
		parameter hssi_tx_pcs_pma_interface_silicon_rev                                           = "14nm5cr2",
		parameter hssi_fifo_rx_pcs_double_read_mode                                               = "double_read_dis",
		parameter hssi_fifo_rx_pcs_prot_mode                                                      = "teng_mode",
		parameter hssi_fifo_rx_pcs_silicon_rev                                                    = "14nm5cr2",
		parameter hssi_fifo_tx_pcs_double_write_mode                                              = "double_write_dis",
		parameter hssi_fifo_tx_pcs_prot_mode                                                      = "teng_mode",
		parameter hssi_fifo_tx_pcs_silicon_rev                                                    = "14nm5cr2",
		parameter pma_cdr_refclk_powerdown_mode                                                   = "powerup",
		parameter pma_cdr_refclk_receiver_detect_src                                              = "iqclk_src",
		parameter pma_cdr_refclk_silicon_rev                                                      = "14nm5cr2",
		parameter pma_cdr_refclk_refclk_select                                                    = "ref_iqclk0",
		parameter pma_rx_odi_datarate_bps                                                         = "25781250000",
		parameter pma_rx_odi_enable_cdr_lpbk                                                      = "disable_lpbk",
		parameter pma_rx_odi_initial_settings                                                     = "true",
		parameter pma_rx_odi_monitor_bw_sel                                                       = "bw_1",
		parameter pma_rx_odi_optimal                                                              = "true",
		parameter pma_rx_odi_phase_steps_64_vs_128                                                = "phase_steps_64",
		parameter pma_rx_odi_phase_steps_sel                                                      = "step40",
		parameter pma_rx_odi_power_mode                                                           = "high_perf",
		parameter pma_rx_odi_prot_mode                                                            = "basic_rx",
		parameter pma_rx_odi_xrx_path_x119_rx_path_rstn_overrideb                                 = "use_sequencer",
		parameter pma_rx_odi_step_ctrl_sel                                                        = "dprio_mode",
		parameter pma_rx_odi_sup_mode                                                             = "user_mode",
		parameter pma_rx_odi_vert_threshold                                                       = "vert_0",
		parameter pma_rx_odi_vreg_voltage_sel                                                     = "vreg3",
		parameter pma_rx_odi_silicon_rev                                                          = "14nm5cr2",
		parameter pma_adapt_sequencer_rx_path_rstn_overrideb                                      = "use_sequencer",
		parameter pma_adapt_sequencer_silicon_rev                                                 = "14nm5cr2",
		parameter pma_adapt_adapt_mode                                                            = "ctle_dfe",
		parameter pma_adapt_adp_ac_ctle_cal_win                                                   = "radp_ac_ctle_cal_win_4",
		parameter pma_adapt_adp_ac_ctle_cocurrent_mode_sel                                        = "radp_ac_ctle_cocurrent_mode_sel_mode_1",
		parameter pma_adapt_adp_ac_ctle_en                                                        = "radp_ac_ctle_en_enable",
		parameter pma_adapt_adp_ac_ctle_hold_en                                                   = "radp_ac_ctle_hold_en_not_hold",
		parameter pma_adapt_adp_ac_ctle_initial_load                                              = "radp_ac_ctle_initial_load_0",
		parameter pma_adapt_adp_ac_ctle_initial_value                                             = "radp_ac_ctle_initial_value_8",
		parameter pma_adapt_adp_ac_ctle_mode_sel                                                  = "radp_ac_ctle_mode_sel_concurrent",
		parameter pma_adapt_adp_ac_ctle_ph1_win                                                   = "radp_ac_ctle_ph1_win_2p19",
		parameter pma_adapt_adp_adapt_control_sel                                                 = "radp_adapt_control_sel_from_cram",
		parameter pma_adapt_adp_adapt_start                                                       = "radp_adapt_start_0",
		parameter pma_adapt_adp_bist_datapath_en                                                  = "radp_bist_datapath_en_disable",
		parameter pma_adapt_adp_bist_errcount_rstn                                                = "radp_bist_errcount_rstn_0",
		parameter pma_adapt_adp_bist_mode_sel                                                     = "radp_bist_mode_sel_prbs31",
		parameter pma_adapt_adp_clkgate_enb                                                       = "radp_clkgate_enb_disable",
		parameter pma_adapt_adp_clkout_div_sel                                                    = "radp_clkout_div_sel_div2_4cycle",
		parameter pma_adapt_adp_ctle_bypass_ac                                                    = "radp_ctle_bypass_ac_not_bypass",
		parameter pma_adapt_adp_ctle_bypass_dc                                                    = "radp_ctle_bypass_dc_not_bypass",
		parameter pma_adapt_adp_dc_ctle_accum_depth                                               = 8,
		parameter pma_adapt_adp_dc_ctle_en                                                        = "radp_dc_ctle_en_enable",
		parameter pma_adapt_adp_dc_ctle_hold_en                                                   = "radp_dc_ctle_hold_en_not_hold",
		parameter pma_adapt_adp_dc_ctle_initial_load                                              = "radp_dc_ctle_initial_load_0",
		parameter pma_adapt_adp_dc_ctle_initial_value                                             = "radp_dc_ctle_initial_value_32",
		parameter pma_adapt_adp_dc_ctle_mode0_win_size                                            = "radp_dc_ctle_mode0_win_size_4_taps",
		parameter pma_adapt_adp_dc_ctle_mode0_win_start                                           = 0,
		parameter pma_adapt_adp_dc_ctle_mode1_h1_ratio                                            = 8,
		parameter pma_adapt_adp_dc_ctle_mode2_h2_limit                                            = 7,
		parameter pma_adapt_adp_dc_ctle_mode_sel                                                  = "radp_dc_ctle_mode_sel_mode_2",
		parameter pma_adapt_adp_dc_ctle_onetime                                                   = "radp_dc_ctle_onetime_disable",
		parameter pma_adapt_adp_dc_ctle_onetime_threshold                                         = "radp_dc_ctle_onetime_threshold_256",
		parameter pma_adapt_adp_dfe_accum_depth                                                   = 8,
		parameter pma_adapt_adp_dfe_en                                                            = "radp_dfe_en_enable",
		parameter pma_adapt_adp_dfe_fxtap_bypass                                                  = "radp_dfe_fxtap_bypass_not_bypass",
		parameter pma_adapt_adp_dfe_hold_en                                                       = "radp_dfe_hold_en_not_hold",
		parameter pma_adapt_adp_dfe_hold_sel                                                      = "radp_dfe_hold_sel_no",
		parameter pma_adapt_adp_dfe_onetime                                                       = "radp_dfe_onetime_disable",
		parameter pma_adapt_adp_dfe_onetime_threshold                                             = "radp_dfe_onetime_threshold_2048",
		parameter pma_adapt_adp_dfe_tap1_initial_load                                             = "radp_dfe_tap1_initial_load_0",
		parameter pma_adapt_adp_dfe_tap1_initial_value                                            = "radp_dfe_tap1_initial_value_0",
		parameter pma_adapt_adp_dfe_tap_sel_en                                                    = "radp_dfe_tap_sel_en_no",
		parameter pma_adapt_adp_dlev_accum_depth                                                  = 6,
		parameter pma_adapt_adp_dlev_bypass                                                       = "radp_dlev_bypass_not_bypass",
		parameter pma_adapt_adp_dlev_en                                                           = "radp_dlev_en_enable",
		parameter pma_adapt_adp_dlev_hold_en                                                      = "radp_dlev_hold_en_not_hold",
		parameter pma_adapt_adp_dlev_initial_load                                                 = "radp_dlev_initial_load_0",
		parameter pma_adapt_adp_dlev_initial_value                                                = "radp_dlev_initial_value_38",
		parameter pma_adapt_adp_dlev_onetime                                                      = "radp_dlev_onetime_disable",
		parameter pma_adapt_adp_dlev_onetime_threshold                                            = "radp_dlev_onetime_threshold_4096",
		parameter pma_adapt_adp_dlev_sel                                                          = "radp_dlev_sel_mux",
		parameter pma_adapt_adp_force_freqlock                                                    = "radp_force_freqlock_use",
		parameter pma_adapt_adp_frame_capture                                                     = "radp_frame_capture_0",
		parameter pma_adapt_adp_frame_en                                                          = "radp_frame_en_disable",
		parameter pma_adapt_adp_frame_odi_sel                                                     = "radp_frame_odi_sel_deser_err",
		parameter pma_adapt_adp_frame_out_sel                                                     = "radp_frame_out_sel_select_a",
		parameter pma_adapt_adp_load_sig_sel                                                      = "radp_load_sig_sel_from_interanl",
		parameter pma_adapt_adp_oc_accum_depth                                                    = 11,
		parameter pma_adapt_adp_oc_bypass                                                         = "radp_oc_bypass_bypass",
		parameter pma_adapt_adp_oc_en                                                             = "radp_oc_en_disable",
		parameter pma_adapt_adp_oc_hold_en                                                        = "radp_oc_hold_en_not_hold",
		parameter pma_adapt_adp_oc_initial_load                                                   = "radp_oc_initial_load_0",
		parameter pma_adapt_adp_oc_initial_sign                                                   = "radp_oc_initial_sign_0",
		parameter pma_adapt_adp_oc_onetime                                                        = "radp_oc_onetime_disable",
		parameter pma_adapt_adp_oc_onetime_threshold                                              = "radp_oc_onetime_threshold_1024",
		parameter pma_adapt_adp_odi_bit_sel                                                       = "radp_odi_bit_sel_all_bits",
		parameter pma_adapt_adp_odi_control_sel                                                   = "radp_odi_control_sel_from_cram",
		parameter pma_adapt_adp_odi_count_threshold                                               = "radp_odi_count_threshold_1e6",
		parameter pma_adapt_adp_odi_dfe_spec_en                                                   = "radp_odi_dfe_spec_en_enable",
		parameter pma_adapt_adp_odi_dlev_sel                                                      = "radp_odi_dlev_sel_0",
		parameter pma_adapt_adp_odi_en                                                            = "radp_odi_en_disable",
		parameter pma_adapt_adp_odi_mode                                                          = "radp_odi_mode_detect_errdata",
		parameter pma_adapt_adp_odi_rstn                                                          = "radp_odi_rstn_1",
		parameter pma_adapt_adp_odi_spec_sel                                                      = "radp_odi_spec_sel_0",
		parameter pma_adapt_adp_odi_start                                                         = "radp_odi_start_0",
		parameter pma_adapt_adp_pat_dlev_sign_avg_win                                             = "radp_pat_dlev_sign_avg_win_2x",
		parameter pma_adapt_adp_pat_dlev_sign_force                                               = "radp_pat_dlev_sign_force_determined_by_cram",
		parameter pma_adapt_adp_pat_dlev_sign_value                                               = "radp_pat_dlev_sign_value_1",
		parameter pma_adapt_adp_pat_spec_sign_avg_win                                             = "radp_pat_spec_sign_avg_win_256",
		parameter pma_adapt_adp_pat_spec_sign_force                                               = "radp_pat_spec_sign_force_generated_internally",
		parameter pma_adapt_adp_pat_spec_sign_value                                               = "radp_pat_spec_sign_value_0",
		parameter pma_adapt_adp_pat_trans_filter                                                  = "radp_pat_trans_filter_5",
		parameter pma_adapt_adp_pat_trans_only_en                                                 = "radp_pat_trans_only_en_enable",
		parameter pma_adapt_adp_pcie_adp_bypass                                                   = "radp_pcie_adp_bypass_no",
		parameter pma_adapt_adp_pcie_eqz                                                          = "radp_pcie_eqz_non_pcie_mode",
		parameter pma_adapt_adp_pcie_hold_sel                                                     = 0,
		parameter pma_adapt_adp_pcs_option                                                        = "radp_pcs_option_0",
		parameter pma_adapt_adp_po_actslp_ratio                                                   = "radp_po_actslp_ratio_10_percent",
		parameter pma_adapt_adp_po_en                                                             = "radp_po_en_disable",
		parameter pma_adapt_adp_po_gb_act2slp                                                     = "radp_po_gb_act2slp_288ns",
		parameter pma_adapt_adp_po_gb_slp2act                                                     = "radp_po_gb_slp2act_288ns",
		parameter pma_adapt_adp_po_initwait                                                       = "radp_po_initwait_10sec",
		parameter pma_adapt_adp_po_sleep_win                                                      = "radp_po_sleep_win_2_sec",
		parameter pma_adapt_adp_reserved                                                          = 0,
		parameter pma_adapt_adp_rstn                                                              = "radp_rstn_1",
		parameter pma_adapt_adp_status_sel                                                        = "radp_status_sel_0",
		parameter pma_adapt_adp_tx_accum_depth                                                    = 4,
		parameter pma_adapt_adp_tx_adp_accumulate                                                 = "radp_tx_adp_accumulate_0",
		parameter pma_adapt_adp_tx_adp_en                                                         = "radp_tx_adp_en_0",
		parameter pma_adapt_adp_tx_up_dn_flip                                                     = "radp_tx_up_dn_flip_0",
		parameter pma_adapt_adp_vga_accum_depth                                                   = 9,
		parameter pma_adapt_adp_vga_bypass                                                        = "radp_vga_bypass_not_bypass",
		parameter pma_adapt_adp_vga_ctle_low_limit                                                = "radp_vga_ctle_low_limit_4",
		parameter pma_adapt_adp_vga_dlev_offset                                                   = 4,
		parameter pma_adapt_adp_vga_dlev_target                                                   = 25,
		parameter pma_adapt_adp_vga_en                                                            = "radp_vga_en_enalbe",
		parameter pma_adapt_adp_vga_hold_en                                                       = "radp_vga_hold_en_not_hold",
		parameter pma_adapt_adp_vga_initial_load                                                  = "radp_vga_initial_load_0",
		parameter pma_adapt_adp_vga_initial_value                                                 = "radp_vga_initial_value_16",
		parameter pma_adapt_adp_vga_onetime                                                       = "radp_vga_onetime_disable",
		parameter pma_adapt_adp_vga_onetime_threshold                                             = "radp_vga_onetime_threshold_512",
		parameter pma_adapt_datarate_bps                                                          = "25781250000",
		parameter pma_adapt_initial_settings                                                      = "true",
		parameter pma_adapt_odi_mode                                                              = "odi_disable",
		parameter pma_adapt_optimal                                                               = "true",
		parameter pma_adapt_power_mode                                                            = "powsav_disable",
		parameter pma_adapt_prot_mode                                                             = "basic_rx",
		parameter pma_adapt_sup_mode                                                              = "user_mode",
		parameter pma_adapt_silicon_rev                                                           = "14nm5cr2",
		parameter pma_rx_dfe_adapt_bti_en                                                         = "adapt_bti_disable",
		parameter pma_rx_dfe_atb_select                                                           = "atb_disable",
		parameter pma_rx_dfe_bti_protected                                                        = "false",
		parameter pma_rx_dfe_datarate_bps                                                         = "25781250000",
		parameter pma_rx_dfe_dfe_bti_en                                                           = "dfe_bti_disable",
		parameter pma_rx_dfe_dfe_mode                                                             = "dfe_tap1_15",
		parameter pma_rx_dfe_dft_en                                                               = "dft_disable",
		parameter pma_rx_dfe_dft_hilospeed_sel                                                    = "dft_osc_lospeed_path",
		parameter pma_rx_dfe_dft_osc_sel                                                          = "dft_osc_even",
		parameter pma_rx_dfe_h1edge_bti_en                                                        = "h1edge_bti_disable",
		parameter pma_rx_dfe_initial_settings                                                     = "true",
		parameter pma_rx_dfe_latch_xcouple_disable                                                = "latch_xcouple_disable",
		parameter pma_rx_dfe_oc_sa_cdr0e                                                          = 0,
		parameter pma_rx_dfe_oc_sa_cdr0e_sgn                                                      = "oc_sa_cdr0e_sgn_0",
		parameter pma_rx_dfe_oc_sa_cdr0o                                                          = 0,
		parameter pma_rx_dfe_oc_sa_cdr0o_sgn                                                      = "oc_sa_cdr0o_sgn_0",
		parameter pma_rx_dfe_oc_sa_cdrne                                                          = 0,
		parameter pma_rx_dfe_oc_sa_cdrne_sgn                                                      = "oc_sa_cdrne_sgn_0",
		parameter pma_rx_dfe_oc_sa_cdrno                                                          = 0,
		parameter pma_rx_dfe_oc_sa_cdrno_sgn                                                      = "oc_sa_cdrno_sgn_0",
		parameter pma_rx_dfe_oc_sa_cdrpe                                                          = 0,
		parameter pma_rx_dfe_oc_sa_cdrpe_sgn                                                      = "oc_sa_cdrpe_sgn_0",
		parameter pma_rx_dfe_oc_sa_cdrpo                                                          = 0,
		parameter pma_rx_dfe_oc_sa_cdrpo_sgn                                                      = "oc_sa_cdrpo_sgn_0",
		parameter pma_rx_dfe_oc_sa_dne                                                            = 0,
		parameter pma_rx_dfe_oc_sa_dne_sgn                                                        = "oc_sa_dne_sgn_0",
		parameter pma_rx_dfe_oc_sa_dno                                                            = 0,
		parameter pma_rx_dfe_oc_sa_dno_sgn                                                        = "oc_sa_dno_sgn_0",
		parameter pma_rx_dfe_oc_sa_dpe                                                            = 0,
		parameter pma_rx_dfe_oc_sa_dpe_sgn                                                        = "oc_sa_dpe_sgn_0",
		parameter pma_rx_dfe_oc_sa_dpo                                                            = 0,
		parameter pma_rx_dfe_oc_sa_dpo_sgn                                                        = "oc_sa_dpo_sgn_0",
		parameter pma_rx_dfe_oc_sa_odie                                                           = 0,
		parameter pma_rx_dfe_oc_sa_odie_sgn                                                       = "oc_sa_odie_sgn_0",
		parameter pma_rx_dfe_oc_sa_odio                                                           = 0,
		parameter pma_rx_dfe_oc_sa_odio_sgn                                                       = "oc_sa_odio_sgn_0",
		parameter pma_rx_dfe_oc_sa_vrefe                                                          = 0,
		parameter pma_rx_dfe_oc_sa_vrefe_sgn                                                      = "oc_sa_vrefe_sgn_0",
		parameter pma_rx_dfe_oc_sa_vrefo                                                          = 0,
		parameter pma_rx_dfe_oc_sa_vrefo_sgn                                                      = "oc_sa_vrefo_sgn_0",
		parameter pma_rx_dfe_odi_bti_en                                                           = "odi_bti_disable",
		parameter pma_rx_dfe_odi_dlev_sign                                                        = "odi_dlev_pos",
		parameter pma_rx_dfe_odi_h1_sign                                                          = "odi_h1_pos",
		parameter pma_rx_dfe_optimal                                                              = "true",
		parameter pma_rx_dfe_pdb                                                                  = "dfe_enable",
		parameter pma_rx_dfe_pdb_edge_pre_h1                                                      = "cdr_pre_h1_enable",
		parameter pma_rx_dfe_pdb_edge_pst_h1                                                      = "cdr_pst_h1_enable",
		parameter pma_rx_dfe_pdb_tap_10t15                                                        = "tap10t15_dfe_enable",
		parameter pma_rx_dfe_pdb_tap_4t9                                                          = "tap4t9_dfe_enable",
		parameter pma_rx_dfe_pdb_tapsum                                                           = "tapsum_enable",
		parameter pma_rx_dfe_power_mode                                                           = "high_perf",
		parameter pma_rx_dfe_prot_mode                                                            = "basic_rx",
		parameter pma_rx_dfe_sel_oc_en                                                            = "off_canc_disable",
		parameter pma_rx_dfe_sel_probe_tstmx                                                      = "probe_tstmx_none",
		parameter pma_rx_dfe_sup_mode                                                             = "user_mode",
		parameter pma_rx_dfe_tap10_coeff                                                          = 0,
		parameter pma_rx_dfe_tap10_sgn                                                            = "tap10_sign_0",
		parameter pma_rx_dfe_tap11_coeff                                                          = 0,
		parameter pma_rx_dfe_tap11_sgn                                                            = "tap11_sign_0",
		parameter pma_rx_dfe_tap12_coeff                                                          = 0,
		parameter pma_rx_dfe_tap12_sgn                                                            = "tap12_sign_0",
		parameter pma_rx_dfe_tap13_coeff                                                          = 0,
		parameter pma_rx_dfe_tap13_sgn                                                            = "tap13_sign_0",
		parameter pma_rx_dfe_tap14_coeff                                                          = 0,
		parameter pma_rx_dfe_tap14_sgn                                                            = "tap14_sign_0",
		parameter pma_rx_dfe_tap15_coeff                                                          = 0,
		parameter pma_rx_dfe_tap15_sgn                                                            = "tap15_sign_0",
		parameter pma_rx_dfe_tap1_coeff                                                           = 0,
		parameter pma_rx_dfe_tap1_sgn                                                             = "tap1_sign_0",
		parameter pma_rx_dfe_tap2_coeff                                                           = 0,
		parameter pma_rx_dfe_tap2_sgn                                                             = "tap2_sign_0",
		parameter pma_rx_dfe_tap3_coeff                                                           = 0,
		parameter pma_rx_dfe_tap3_sgn                                                             = "tap3_sign_0",
		parameter pma_rx_dfe_tap4_coeff                                                           = 0,
		parameter pma_rx_dfe_tap4_sgn                                                             = "tap4_sign_0",
		parameter pma_rx_dfe_tap5_coeff                                                           = 0,
		parameter pma_rx_dfe_tap5_sgn                                                             = "tap5_sign_0",
		parameter pma_rx_dfe_tap6_coeff                                                           = 0,
		parameter pma_rx_dfe_tap6_sgn                                                             = "tap6_sign_0",
		parameter pma_rx_dfe_tap7_coeff                                                           = 0,
		parameter pma_rx_dfe_tap7_sgn                                                             = "tap7_sign_0",
		parameter pma_rx_dfe_tap8_coeff                                                           = 0,
		parameter pma_rx_dfe_tap8_sgn                                                             = "tap8_sign_0",
		parameter pma_rx_dfe_tap9_coeff                                                           = 0,
		parameter pma_rx_dfe_tap9_sgn                                                             = "tap9_sign_0",
		parameter pma_rx_dfe_tapsum_bw_sel                                                        = "tapsum_hibw",
		parameter pma_rx_dfe_vref_coeff                                                           = 0,
		parameter pma_rx_dfe_silicon_rev                                                          = "14nm5cr2",
		parameter pma_rx_sd_link                                                                  = "sr",
		parameter pma_rx_sd_optimal                                                               = "true",
		parameter pma_rx_sd_power_mode                                                            = "high_perf",
		parameter pma_rx_sd_prot_mode                                                             = "basic_rx",
		parameter pma_rx_sd_sd_output_off                                                         = "clk_divrx_2",
		parameter pma_rx_sd_sd_output_on                                                          = "force_sd_output_on",
		parameter pma_rx_sd_sd_pdb                                                                = "sd_off",
		parameter pma_rx_sd_sd_threshold                                                          = "sdlv_3",
		parameter pma_rx_sd_sup_mode                                                              = "user_mode",
		parameter pma_rx_sd_silicon_rev                                                           = "14nm5cr2",
		parameter pma_pcie_gen_switch_silicon_rev                                                 = "14nm5cr2"
	) (
		input  wire [3:0]   tx_analogreset,          //          tx_analogreset.tx_analogreset
		input  wire [3:0]   rx_analogreset,          //          rx_analogreset.rx_analogreset
		input  wire [3:0]   tx_digitalreset,         //         tx_digitalreset.tx_digitalreset
		input  wire [3:0]   rx_digitalreset,         //         rx_digitalreset.rx_digitalreset
		output wire [3:0]   tx_analogreset_stat,     //     tx_analogreset_stat.tx_analogreset_stat
		output wire [3:0]   rx_analogreset_stat,     //     rx_analogreset_stat.rx_analogreset_stat
		output wire [3:0]   tx_digitalreset_stat,    //    tx_digitalreset_stat.tx_digitalreset_stat
		output wire [3:0]   rx_digitalreset_stat,    //    rx_digitalreset_stat.rx_digitalreset_stat
		output wire [3:0]   tx_dll_lock,             //             tx_dll_lock.tx_dll_lock
		output wire [3:0]   tx_cal_busy,             //             tx_cal_busy.tx_cal_busy
		output wire [3:0]   rx_cal_busy,             //             rx_cal_busy.rx_cal_busy
		input  wire [3:0]   tx_serial_clk0,          //          tx_serial_clk0.clk
		input  wire         rx_cdr_refclk0,          //          rx_cdr_refclk0.clk
		output wire [3:0]   tx_serial_data,          //          tx_serial_data.tx_serial_data
		input  wire [3:0]   rx_serial_data,          //          rx_serial_data.rx_serial_data
		input  wire [3:0]   rx_seriallpbken,         //         rx_seriallpbken.rx_seriallpbken
		input  wire [3:0]   rx_set_locktodata,       //       rx_set_locktodata.rx_set_locktodata
		input  wire [3:0]   rx_set_locktoref,        //        rx_set_locktoref.rx_set_locktoref
		output wire [3:0]   rx_is_lockedtoref,       //       rx_is_lockedtoref.rx_is_lockedtoref
		output wire [3:0]   rx_is_lockedtodata,      //      rx_is_lockedtodata.rx_is_lockedtodata
		input  wire [3:0]   tx_coreclkin,            //            tx_coreclkin.clk
		input  wire [3:0]   rx_coreclkin,            //            rx_coreclkin.clk
		output wire [3:0]   tx_clkout,               //               tx_clkout.clk
		output wire [3:0]   tx_clkout2,              //              tx_clkout2.clk
		output wire [3:0]   rx_clkout,               //               rx_clkout.clk
		output wire [3:0]   rx_clkout2,              //              rx_clkout2.clk
		output wire [3:0]   rx_pma_iqtxrx_clkout,    //    rx_pma_iqtxrx_clkout.clk
		input  wire [255:0] tx_parallel_data,        //        tx_parallel_data.tx_parallel_data
		input  wire [7:0]   tx_control,              //              tx_control.tx_control
		input  wire [3:0]   tx_enh_data_valid,       //       tx_enh_data_valid.tx_enh_data_valid
		input  wire [3:0]   tx_fifo_wr_en,           //           tx_fifo_wr_en.tx_fifo_wr_en
		input  wire [47:0]  unused_tx_parallel_data, // unused_tx_parallel_data.unused_tx_parallel_data
		output wire [255:0] rx_parallel_data,        //        rx_parallel_data.rx_parallel_data
		output wire [7:0]   rx_control,              //              rx_control.rx_control
		output wire [3:0]   rx_enh_data_valid,       //       rx_enh_data_valid.rx_enh_data_valid
		output wire [3:0]   rx_data_valid,           //           rx_data_valid.rx_data_valid
		output wire [47:0]  unused_rx_parallel_data, // unused_rx_parallel_data.unused_rx_parallel_data
		input  wire [3:0]   rx_bitslip,              //              rx_bitslip.rx_bitslip
		output wire [3:0]   tx_fifo_full,            //            tx_fifo_full.tx_fifo_full
		output wire [3:0]   tx_fifo_empty,           //           tx_fifo_empty.tx_fifo_empty
		output wire [3:0]   tx_fifo_pfull,           //           tx_fifo_pfull.tx_fifo_pfull
		output wire [3:0]   tx_fifo_pempty,          //          tx_fifo_pempty.tx_fifo_pempty
		output wire [3:0]   rx_fifo_full,            //            rx_fifo_full.rx_fifo_full
		output wire [3:0]   rx_fifo_empty,           //           rx_fifo_empty.rx_fifo_empty
		output wire [3:0]   rx_fifo_pfull,           //           rx_fifo_pfull.rx_fifo_pfull
		output wire [3:0]   rx_fifo_pempty,          //          rx_fifo_pempty.rx_fifo_pempty
		input  wire [3:0]   rx_fifo_rd_en,           //           rx_fifo_rd_en.rx_fifo_rd_en
		input  wire [0:0]   reconfig_clk,            //            reconfig_clk.clk
		input  wire [0:0]   reconfig_reset,          //          reconfig_reset.reset
		input  wire [0:0]   reconfig_write,          //           reconfig_avmm.write
		input  wire [0:0]   reconfig_read,           //                        .read
		input  wire [12:0]  reconfig_address,        //                        .address
		input  wire [31:0]  reconfig_writedata,      //                        .writedata
		output wire [31:0]  reconfig_readdata,       //                        .readdata
		output wire [0:0]   reconfig_waitrequest     //                        .waitrequest
	);

	wire  [319:0] caui4_xcvr_644_rx_parallel_data; // port fragment

	generate
		// If any of the display statements (or deliberately broken
		// instantiations) within this generate block triggers then this module
		// has been instantiated this module with a set of parameters different
		// from those it was generated for.  This will usually result in a
		// non-functioning system.
		if (rcfg_enable != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_enable_check ( .error(1'b1) );
		end
		if (rcfg_jtag_enable != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_jtag_enable_check ( .error(1'b1) );
		end
		if (rcfg_separate_avmm_busy != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_separate_avmm_busy_check ( .error(1'b1) );
		end
		if (dbg_embedded_debug_enable != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_embedded_debug_enable_check ( .error(1'b1) );
		end
		if (dbg_capability_reg_enable != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_capability_reg_enable_check ( .error(1'b1) );
		end
		if (dbg_user_identifier != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_user_identifier_check ( .error(1'b1) );
		end
		if (dbg_stat_soft_logic_enable != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_stat_soft_logic_enable_check ( .error(1'b1) );
		end
		if (dbg_ctrl_soft_logic_enable != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_ctrl_soft_logic_enable_check ( .error(1'b1) );
		end
		if (rcfg_emb_strm_enable != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_emb_strm_enable_check ( .error(1'b1) );
		end
		if (rcfg_profile_cnt != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_profile_cnt_check ( .error(1'b1) );
		end
		if (device_revision != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					device_revision_check ( .error(1'b1) );
		end
		if (silicon_revision != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					silicon_revision_check ( .error(1'b1) );
		end
		if (reduced_reset_sim_time != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					reduced_reset_sim_time_check ( .error(1'b1) );
		end
		if (duplex_mode != "duplex")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					duplex_mode_check ( .error(1'b1) );
		end
		if (channels != 4)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					channels_check ( .error(1'b1) );
		end
		if (enable_calibration != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_calibration_check ( .error(1'b1) );
		end
		if (enable_direct_reset_control != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_direct_reset_control_check ( .error(1'b1) );
		end
		if (disable_reset_sequencer != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					disable_reset_sequencer_check ( .error(1'b1) );
		end
		if (disable_digital_reset_sequencer != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					disable_digital_reset_sequencer_check ( .error(1'b1) );
		end
		if (l_release_aib_reset_first != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					l_release_aib_reset_first_check ( .error(1'b1) );
		end
		if (bonded_mode != "not_bonded")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					bonded_mode_check ( .error(1'b1) );
		end
		if (pcs_bonding_master != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pcs_bonding_master_check ( .error(1'b1) );
		end
		if (pcs_reset_sequencing_mode != "bonded")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pcs_reset_sequencing_mode_check ( .error(1'b1) );
		end
		if (enable_manual_bonding_settings != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_manual_bonding_settings_check ( .error(1'b1) );
		end
		if (manual_pcs_bonding_mode != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_pcs_bonding_mode_check ( .error(1'b1) );
		end
		if (manual_pcs_bonding_comp_cnt != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_pcs_bonding_comp_cnt_check ( .error(1'b1) );
		end
		if (manual_tx_hssi_aib_bonding_mode != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_tx_hssi_aib_bonding_mode_check ( .error(1'b1) );
		end
		if (manual_tx_hssi_aib_bonding_comp_cnt != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_tx_hssi_aib_bonding_comp_cnt_check ( .error(1'b1) );
		end
		if (manual_tx_core_aib_bonding_mode != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_tx_core_aib_bonding_mode_check ( .error(1'b1) );
		end
		if (manual_tx_core_aib_bonding_comp_cnt != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_tx_core_aib_bonding_comp_cnt_check ( .error(1'b1) );
		end
		if (manual_rx_hssi_aib_bonding_mode != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_rx_hssi_aib_bonding_mode_check ( .error(1'b1) );
		end
		if (manual_rx_hssi_aib_bonding_comp_cnt != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_rx_hssi_aib_bonding_comp_cnt_check ( .error(1'b1) );
		end
		if (manual_rx_core_aib_bonding_mode != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_rx_core_aib_bonding_mode_check ( .error(1'b1) );
		end
		if (manual_rx_core_aib_bonding_comp_cnt != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					manual_rx_core_aib_bonding_comp_cnt_check ( .error(1'b1) );
		end
		if (plls != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					plls_check ( .error(1'b1) );
		end
		if (number_physical_bonding_clocks != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					number_physical_bonding_clocks_check ( .error(1'b1) );
		end
		if (cdr_refclk_cnt != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_refclk_cnt_check ( .error(1'b1) );
		end
		if (enable_hip != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_hip_check ( .error(1'b1) );
		end
		if (hip_cal_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hip_cal_en_check ( .error(1'b1) );
		end
		if (enable_ehip != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_ehip_check ( .error(1'b1) );
		end
		if (enable_tx_fast_pipeln_reg != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_tx_fast_pipeln_reg_check ( .error(1'b1) );
		end
		if (enable_rx_fast_pipeln_reg != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_rx_fast_pipeln_reg_check ( .error(1'b1) );
		end
		if (tx_coreclkin_clock_network != "dedicated")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					tx_coreclkin_clock_network_check ( .error(1'b1) );
		end
		if (tx_pcs_bonding_clock_network != "dedicated")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					tx_pcs_bonding_clock_network_check ( .error(1'b1) );
		end
		if (rx_coreclkin_clock_network != "dedicated")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rx_coreclkin_clock_network_check ( .error(1'b1) );
		end
		if (osc_clk_divider != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					osc_clk_divider_check ( .error(1'b1) );
		end
		if (enable_tx_x2_coreclkin_port != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_tx_x2_coreclkin_port_check ( .error(1'b1) );
		end
		if (rcfg_shared != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_shared_check ( .error(1'b1) );
		end
		if (adme_prot_mode != "basic_enh")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					adme_prot_mode_check ( .error(1'b1) );
		end
		if (adme_pma_mode != "basic")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					adme_pma_mode_check ( .error(1'b1) );
		end
		if (adme_tx_power_mode != "high_perf")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					adme_tx_power_mode_check ( .error(1'b1) );
		end
		if (adme_data_rate != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					adme_data_rate_check ( .error(1'b1) );
		end
		if (dbg_prbs_soft_logic_enable != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_prbs_soft_logic_enable_check ( .error(1'b1) );
		end
		if (dbg_odi_soft_logic_enable != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_odi_soft_logic_enable_check ( .error(1'b1) );
		end
		if (enable_rcfg_tx_digitalreset_release_ctrl != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_rcfg_tx_digitalreset_release_ctrl_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_advanced_user_mode_rx != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_advanced_user_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs8g_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs8g_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_clklow_clk_hz != 322265625)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_clklow_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_ctrl_plane_bonding_rx != "individual_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_ctrl_plane_bonding_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_fifo_mode_rx != "reg_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_fifo_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs8g_fifo_mode_rx != "reg_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs8g_fifo_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_fref_clk_hz != 322265625)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_fref_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_frequency_rules_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_frequency_rules_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_func_mode != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_func_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_hclk_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_hclk_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_hip_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_hip_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs8g_hip_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs8g_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_hrdrstctl_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_hrdrstctl_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_hrdrstctl_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_hrdrstctl_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_low_latency_en_rx != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_low_latency_en_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_low_latency_en_rx != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_low_latency_en_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs8g_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs8g_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_operating_voltage != "standard")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_operating_voltage_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_ac_pwr_rules_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_ac_pwr_rules_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_pair_ac_pwr_uw_per_mhz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_pair_ac_pwr_uw_per_mhz_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_rx_ac_pwr_uw_per_mhz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_rx_ac_pwr_uw_per_mhz_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_pcs_rx_block_sel != "teng")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_pcs_rx_block_sel_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel != "teng_clk_out")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_pcs_rx_clk_sel != "pcs_rx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_pcs_rx_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en != "hip_rx_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_pcs_rx_output_sel != "teng_output")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_pcs_rx_output_sel_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_rx_pwr_scaling_clk != "pma_rx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_rx_pwr_scaling_clk_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_8g_refclk_dig_nonatpg_mode_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_8g_refclk_dig_nonatpg_mode_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_fifo_mode_rx != "reg_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_fifo_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_pcs_refclk_dig_nonatpg_mode_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_pcs_refclk_dig_nonatpg_mode_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_rx_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_rx_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_pma_dw_rx != "pma_64b_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_pma_dw_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs8g_pma_dw_rx != "pma_10b_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs8g_pma_dw_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_dw_rx != "pma_64b_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_dw_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_pma_dw_rx != "pma_64b_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_pma_dw_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_rx_clk_hz != 402832031)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_rx_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_g3pcs_prot_mode != "disabled_prot_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_g3pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx != "disabled_prot_mode_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_prot_mode_rx != "basic_mode_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_prot_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs8g_prot_mode_rx != "disabled_prot_mode_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs8g_prot_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_prot_mode_rx != "basic_10gpcs_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_prot_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_prot_mode_rx != "teng_reg_mode_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_prot_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_prot_mode_rx != "teng_basic_mode_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_prot_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_prot_mode_rx != "teng_mode_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_prot_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_shared_fifo_width_rx != "single_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_shared_fifo_width_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_shared_fifo_width_rx != "single_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_shared_fifo_width_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_shared_fifo_width_rx != "single_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_shared_fifo_width_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_sim_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_sim_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_speed_grade != "e2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_speed_grade_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_g3pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_g3pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_krfec_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_krfec_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs8g_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs8g_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode != "tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs10g_test_bus_mode != "rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs10g_test_bus_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_hd_pcs_channel_transparent_pcs_rx != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_hd_pcs_channel_transparent_pcs_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pld_pcs_interface_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pld_pcs_interface_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs10g_advanced_user_mode_tx != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs10g_advanced_user_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs10g_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs10g_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs8g_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs8g_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_ctrl_plane_bonding != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_ctrl_plane_bonding_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_ctrl_plane_bonding_tx != "individual_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_ctrl_plane_bonding_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs10g_fifo_mode_tx != "reg_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs10g_fifo_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs8g_fifo_mode_tx != "reg_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs8g_fifo_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_frequency_rules_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_frequency_rules_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_func_mode != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_func_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_hclk_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_hclk_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_hip_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_hip_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs8g_hip_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs8g_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_hrdrstctl_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_hrdrstctl_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_hrdrstctl_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_hrdrstctl_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs10g_low_latency_en_tx != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs10g_low_latency_en_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_low_latency_en_tx != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_low_latency_en_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs10g_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs10g_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs8g_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs8g_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pcs_tx_ac_pwr_uw_per_mhz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pcs_tx_ac_pwr_uw_per_mhz_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel != "teng_clk_out")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_clk_source != "teng")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_clk_source_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_data_source != "hip_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_data_source_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en != "delay1_clk_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel != "pcs_tx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl != "delay1_path0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel != "one_ff_delay")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en != "delay2_clk_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl != "delay2_path0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_pcs_tx_output_sel != "teng_output")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_pcs_tx_output_sel_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pcs_tx_pwr_scaling_clk != "pma_tx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pcs_tx_pwr_scaling_clk_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_8g_refclk_dig_nonatpg_mode_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_8g_refclk_dig_nonatpg_mode_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_fifo_mode_tx != "reg_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_fifo_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_pcs_refclk_dig_nonatpg_mode_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_pcs_refclk_dig_nonatpg_mode_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_tx_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_tx_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_uhsif_tx_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_uhsif_tx_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs10g_pma_dw_tx != "pma_64b_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs10g_pma_dw_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs8g_pma_dw_tx != "pma_10b_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs8g_pma_dw_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_dw_tx != "pma_64b_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_dw_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_pma_dw_tx != "pma_64b_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_pma_dw_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_tx_clk_hz != 402832031)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_tx_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_g3pcs_prot_mode != "disabled_prot_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_g3pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx != "disabled_prot_mode_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs10g_prot_mode_tx != "basic_mode_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs10g_prot_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs8g_prot_mode_tx != "disabled_prot_mode_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs8g_prot_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_prot_mode_tx != "basic_10gpcs_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_prot_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_prot_mode_tx != "teng_reg_mode_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_prot_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_prot_mode_tx != "teng_basic_mode_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_prot_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_prot_mode_tx != "teng_mode_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_prot_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs10g_shared_fifo_width_tx != "single_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs10g_shared_fifo_width_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_shared_fifo_width_tx != "single_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_shared_fifo_width_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_shared_fifo_width_tx != "single_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_shared_fifo_width_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_sim_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_sim_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_speed_grade != "e2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_speed_grade_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_g3pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_g3pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_krfec_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_krfec_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs10g_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs10g_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs8g_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs8g_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pld_pcs_interface_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pld_pcs_interface_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_advanced_user_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_advanced_user_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_bitslip_en != "bitslip_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_bitslip_en_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_bonding_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_bonding_dft_en_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_bonding_dft_val != "dft_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_bonding_dft_val_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_crcgen_bypass != "crcgen_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_crcgen_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_crcgen_clken != "crcgen_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_crcgen_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_crcgen_err != "crcgen_err_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_crcgen_err_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_crcgen_inv != "crcgen_inv_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_crcgen_inv_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_ctrl_bit_reverse != "ctrl_bit_reverse_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_ctrl_bit_reverse_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_data_bit_reverse != "data_bit_reverse_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_data_bit_reverse_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_dft_clk_out_sel != "tx_master_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_dft_clk_out_sel_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_dispgen_bypass != "dispgen_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_dispgen_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_dispgen_clken != "dispgen_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_dispgen_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_dispgen_err != "dispgen_err_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_dispgen_err_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_dispgen_pipeln != "dispgen_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_dispgen_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_distdwn_bypass_pipeln != "distdwn_bypass_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_distdwn_bypass_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_distup_bypass_pipeln != "distup_bypass_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_distup_bypass_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_dv_bond != "dv_bond_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_dv_bond_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_empty_flag_type != "empty_rd_side")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_empty_flag_type_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_enc64b66b_txsm_clken != "enc64b66b_txsm_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_enc64b66b_txsm_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_enc_64b66b_txsm_bypass != "enc_64b66b_txsm_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_enc_64b66b_txsm_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_fastpath != "fastpath_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_fastpath_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_fec_clken != "fec_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_fec_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_fec_enable != "fec_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_fec_enable_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_fifo_double_write != "fifo_double_write_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_fifo_double_write_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_fifo_reg_fast != "fifo_reg_fast_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_fifo_reg_fast_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_fifo_stop_rd != "n_rd_empty")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_fifo_stop_rd_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_fifo_stop_wr != "n_wr_full")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_fifo_stop_wr_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_frmgen_burst != "frmgen_burst_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_frmgen_burst_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_frmgen_bypass != "frmgen_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_frmgen_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_frmgen_clken != "frmgen_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_frmgen_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_frmgen_mfrm_length != 2048)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_frmgen_mfrm_length_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_frmgen_pipeln != "frmgen_pipeln_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_frmgen_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_frmgen_pyld_ins != "frmgen_pyld_ins_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_frmgen_pyld_ins_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_frmgen_wordslip != "frmgen_wordslip_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_frmgen_wordslip_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_full_flag_type != "full_wr_side")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_full_flag_type_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_gb_pipeln_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_gb_pipeln_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_gb_tx_idwidth != "idwidth_66")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_gb_tx_idwidth_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_gb_tx_odwidth != "odwidth_64")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_gb_tx_odwidth_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_gbred_clken != "gbred_clk_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_gbred_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_indv != "indv_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_indv_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_low_latency_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_low_latency_en_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_master_clk_sel != "master_tx_pma_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_master_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_pempty_flag_type != "pempty_rd_side")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_pempty_flag_type_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_pfull_flag_type != "pfull_wr_side")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_pfull_flag_type_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_phcomp_rd_del != "phcomp_rd_del2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_phcomp_rd_del_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_pld_if_type != "reg")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_pld_if_type_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_prot_mode != "basic_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_pseudo_random != "all_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_pseudo_random_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_pseudo_seed_a != "288230376151711743")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_pseudo_seed_a_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_pseudo_seed_b != "288230376151711743")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_pseudo_seed_b_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_random_disp != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_random_disp_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_rdfifo_clken != "rdfifo_clk_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_rdfifo_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_scrm_bypass != "scrm_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_scrm_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_scrm_clken != "scrm_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_scrm_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_scrm_mode != "async")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_scrm_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_scrm_pipeln != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_scrm_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_sh_err != "sh_err_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_sh_err_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_sop_mark != "sop_mark_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_sop_mark_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_stretch_num_stages != "one_stage")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_stretch_num_stages_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_test_mode != "test_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_test_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_tx_scrm_err != "scrm_err_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_tx_scrm_err_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_tx_scrm_width != "bit64")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_tx_scrm_width_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_tx_sh_location != "msb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_tx_sh_location_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_tx_sm_bypass != "tx_sm_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_tx_sm_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_tx_sm_pipeln != "tx_sm_pipeln_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_tx_sm_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_tx_testbus_sel != "tx_fifo_testbus1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_tx_testbus_sel_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_txfifo_empty != "empty_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_txfifo_empty_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_txfifo_full != "full_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_txfifo_full_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_txfifo_mode != "register_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_txfifo_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_txfifo_pempty != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_txfifo_pempty_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_txfifo_pfull != 11)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_txfifo_pfull_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_wr_clk_sel != "wr_tx_pma_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_wr_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_wrfifo_clken != "wrfifo_clk_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_wrfifo_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_tx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_tx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_auto_error_replacement != "dis_err_replace")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_auto_error_replacement_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_bit_reversal != "dis_bit_reversal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_bit_reversal_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_bonding_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_bonding_dft_en_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_bonding_dft_val != "dft_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_bonding_dft_val_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_bypass_pipeline_reg != "dis_bypass_pipeline")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_bypass_pipeline_reg_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_byte_deserializer != "dis_bds")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_byte_deserializer_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask != "dis_rxvalid_mask")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clkcmp_pattern_n != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clkcmp_pattern_n_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clkcmp_pattern_p != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clkcmp_pattern_p_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_bds_dec_asn != "en_bds_dec_asn_clk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_bds_dec_asn_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_cdr_eidle != "en_cdr_eidle_clk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_cdr_eidle_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk != "en_dw_pc_wrclk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_dw_rm_rd != "en_dw_rm_rdclk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_dw_rm_rd_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_dw_rm_wr != "en_dw_rm_wrclk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_dw_rm_wr_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_dw_wa != "en_dw_wa_clk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_dw_wa_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_pc_rdclk != "en_pc_rdclk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_pc_rdclk_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk != "en_sw_pc_wrclk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_sw_rm_rd != "en_sw_rm_rdclk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_sw_rm_rd_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_sw_rm_wr != "en_sw_rm_wrclk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_sw_rm_wr_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_gate_sw_wa != "en_sw_wa_clk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_gate_sw_wa_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_clock_observation_in_pld_core != "internal_sw_wa_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_clock_observation_in_pld_core_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_eidle_entry_eios != "dis_eidle_eios")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_eidle_entry_eios_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_eidle_entry_iei != "dis_eidle_iei")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_eidle_entry_iei_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_eidle_entry_sd != "dis_eidle_sd")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_eidle_entry_sd_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_eightb_tenb_decoder != "en_8b10b_ibm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_eightb_tenb_decoder_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_err_flags_sel != "err_flags_wa")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_err_flags_sel_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_fixed_pat_det != "dis_fixed_patdet")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_fixed_pat_det_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_fixed_pat_num != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_fixed_pat_num_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_force_signal_detect != "en_force_signal_detect")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_force_signal_detect_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_gen3_clk_en != "disable_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_gen3_clk_en_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_gen3_rx_clk_sel != "rcvd_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_gen3_rx_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_gen3_tx_clk_sel != "tx_pma_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_gen3_tx_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_hip_mode != "dis_hip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_ibm_invalid_code != "dis_ibm_invalid_code")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_ibm_invalid_code_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_invalid_code_flag_only != "dis_invalid_code_only")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_invalid_code_flag_only_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_pad_or_edb_error_replace != "replace_edb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_pad_or_edb_error_replace_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_pcs_bypass != "dis_pcs_bypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_pcs_bypass_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_phase_comp_rdptr != "disable_rdptr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_phase_comp_rdptr_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_phase_compensation_fifo != "register_fifo")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_phase_compensation_fifo_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_pipe_if_enable != "dis_pipe_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_pipe_if_enable_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_pma_dw != "ten_bit")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_pma_dw_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_polinv_8b10b_dec != "dis_polinv_8b10b_dec")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_polinv_8b10b_dec_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_prot_mode != "disabled_prot_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rate_match != "dis_rm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rate_match_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rate_match_del_thres != "dis_rm_del_thres")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rate_match_del_thres_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rate_match_empty_thres != "dis_rm_empty_thres")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rate_match_empty_thres_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rate_match_full_thres != "dis_rm_full_thres")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rate_match_full_thres_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rate_match_ins_thres != "dis_rm_ins_thres")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rate_match_ins_thres_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rate_match_start_thres != "dis_rm_start_thres")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rate_match_start_thres_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rx_clk2 != "rcvd_clk_clk2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rx_clk2_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rx_clk_free_running != "en_rx_clk_free_run")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rx_clk_free_running_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rx_pcs_urst != "en_rx_pcs_urst")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rx_pcs_urst_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rx_rcvd_clk != "rcvd_clk_rcvd_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rx_rcvd_clk_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rx_rd_clk != "rx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rx_rd_clk_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rx_refclk != "dis_refclk_sel")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rx_refclk_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_rx_wr_clk != "rx_clk2_div_1_2_4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_rx_wr_clk_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_symbol_swap != "dis_symbol_swap")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_symbol_swap_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_sync_sm_idle_eios != "dis_syncsm_idle")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_sync_sm_idle_eios_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_test_bus_sel != "tx_testbus")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_test_bus_sel_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_tx_rx_parallel_loopback != "dis_plpbk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_tx_rx_parallel_loopback_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_boundary_lock_ctrl != "sync_sm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_boundary_lock_ctrl_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_clk_slip_spacing != 16)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_clk_slip_spacing_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_det_latency_sync_status_beh != "dont_care_assert_sync")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_det_latency_sync_status_beh_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_disp_err_flag != "en_disp_err_flag")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_disp_err_flag_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_kchar != "dis_kchar")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_kchar_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_pd != "wa_pd_10")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_pd_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_pd_data != "0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_pd_data_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_pd_polarity != "dont_care_both_pol")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_pd_polarity_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_pld_controlled != "dis_pld_ctrl")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_pld_controlled_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_renumber_data != 3)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_renumber_data_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_rgnumber_data != 3)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_rgnumber_data_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_rknumber_data != 3)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_rknumber_data_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_rosnumber_data != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_rosnumber_data_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_rvnumber_data != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_rvnumber_data_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wa_sync_sm_ctrl != "gige_sync_sm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wa_sync_sm_ctrl_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_wait_cnt != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_wait_cnt_check ( .error(1'b1) );
		end
		if (hssi_8g_rx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_rx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_bit_reversal != "dis_bit_reversal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_bit_reversal_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_bonding_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_bonding_dft_en_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_bonding_dft_val != "dft_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_bonding_dft_val_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_bypass_pipeline_reg != "dis_bypass_pipeline")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_bypass_pipeline_reg_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_byte_serializer != "dis_bs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_byte_serializer_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_clock_gate_bs_enc != "en_bs_enc_clk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_clock_gate_bs_enc_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_clock_gate_dw_fifowr != "en_dw_fifowr_clk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_clock_gate_dw_fifowr_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_clock_gate_fiford != "en_fiford_clk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_clock_gate_fiford_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_clock_gate_sw_fifowr != "en_sw_fifowr_clk_gating")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_clock_gate_sw_fifowr_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_clock_observation_in_pld_core != "internal_refclk_b")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_clock_observation_in_pld_core_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_data_selection_8b10b_encoder_input != "normal_data_path")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_data_selection_8b10b_encoder_input_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_dynamic_clk_switch != "dis_dyn_clk_switch")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_dynamic_clk_switch_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_eightb_tenb_disp_ctrl != "dis_disp_ctrl")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_eightb_tenb_disp_ctrl_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_eightb_tenb_encoder != "en_8b10b_ibm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_eightb_tenb_encoder_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_force_echar != "dis_force_echar")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_force_echar_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_force_kchar != "dis_force_kchar")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_force_kchar_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_gen3_tx_clk_sel != "dis_tx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_gen3_tx_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel != "dis_tx_pipe_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_hip_mode != "dis_hip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_pcs_bypass != "dis_pcs_bypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_pcs_bypass_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_phase_comp_rdptr != "disable_rdptr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_phase_comp_rdptr_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_phase_compensation_fifo != "register_fifo")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_phase_compensation_fifo_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_phfifo_write_clk_sel != "tx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_phfifo_write_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_pma_dw != "ten_bit")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_pma_dw_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_prot_mode != "disabled_prot_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_refclk_b_clk_sel != "tx_pma_clock")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_refclk_b_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_revloop_back_rm != "dis_rev_loopback_rx_rm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_revloop_back_rm_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_symbol_swap != "dis_symbol_swap")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_symbol_swap_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_tx_bitslip != "dis_tx_bitslip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_tx_bitslip_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_tx_compliance_controlled_disparity != "dis_txcompliance")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_tx_compliance_controlled_disparity_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_tx_fast_pld_reg != "dis_tx_fast_pld_reg")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_tx_fast_pld_reg_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_txclk_freerun != "en_freerun_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_txclk_freerun_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_txpcs_urst != "en_txpcs_urst")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_txpcs_urst_check ( .error(1'b1) );
		end
		if (hssi_8g_tx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_8g_tx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pcs_arbiter_ctrl != "avmm1_arbiter_uc_sel")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pcs_arbiter_ctrl_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pcs_cal_done != "avmm1_cal_done_deassert")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pcs_cal_done_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pcs_cal_reserved != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pcs_cal_reserved_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pcs_calibration_feature_en != "avmm1_pcs_calibration_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pcs_calibration_feature_en_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pldadapt_gate_dis != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pldadapt_gate_dis_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pcs_hip_cal_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pcs_hip_cal_en_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_hssiadapt_nfhssi_calibratio_feature_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_hssiadapt_nfhssi_calibratio_feature_en_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pldadapt_nfhssi_calibratio_feature_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pldadapt_nfhssi_calibratio_feature_en_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_hssiadapt_read_blocking_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_hssiadapt_read_blocking_enable_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pldadapt_read_blocking_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pldadapt_read_blocking_enable_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_hssiadapt_uc_blocking_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_hssiadapt_uc_blocking_enable_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pldadapt_uc_blocking_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pldadapt_uc_blocking_enable_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_hssiadapt_avmm_osc_clock_setting != "osc_clk_div_by1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_hssiadapt_avmm_osc_clock_setting_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pldadapt_avmm_osc_clock_setting != "osc_clk_div_by1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pldadapt_avmm_osc_clock_setting_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_hssiadapt_avmm_testbus_sel != "avmm1_transfer_testbus")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_hssiadapt_avmm_testbus_sel_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pldadapt_avmm_testbus_sel != "avmm1_transfer_testbus")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pldadapt_avmm_testbus_sel_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_hssiadapt_hip_mode != "disable_hip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_hssiadapt_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_pldadapt_hip_mode != "disable_hip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_pldadapt_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_avmm1_if_calibration_type != "one_time")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_avmm1_if_calibration_type_check ( .error(1'b1) );
		end
		if (pma_cgb_bitslip_enable != "disable_bitslip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_bitslip_enable_check ( .error(1'b1) );
		end
		if (pma_cgb_bti_protected != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_bti_protected_check ( .error(1'b1) );
		end
		if (pma_cgb_cgb_bti_en != "cgb_bti_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_cgb_bti_en_check ( .error(1'b1) );
		end
		if (pma_cgb_cgb_power_down != "normal_cgb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_cgb_power_down_check ( .error(1'b1) );
		end
		if (pma_cgb_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_cgb_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_initial_settings_check ( .error(1'b1) );
		end
		if (pma_cgb_observe_cgb_clocks != "observe_nothing")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_observe_cgb_clocks_check ( .error(1'b1) );
		end
		if (pma_cgb_pcie_gen != "non_pcie")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_pcie_gen_check ( .error(1'b1) );
		end
		if (pma_cgb_pcie_gen3_bitwidth != "pciegen3_wide")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_pcie_gen3_bitwidth_check ( .error(1'b1) );
		end
		if (pma_cgb_power_rail_er != 1120)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_power_rail_er_check ( .error(1'b1) );
		end
		if (pma_cgb_prot_mode != "basic_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_prot_mode_check ( .error(1'b1) );
		end
		if (pma_cgb_ser_mode != "sixty_four_bit")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_ser_mode_check ( .error(1'b1) );
		end
		if (pma_cgb_ser_powerdown != "normal_poweron_ser")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_ser_powerdown_check ( .error(1'b1) );
		end
		if (pma_cgb_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_sup_mode_check ( .error(1'b1) );
		end
		if (pma_cgb_tx_ucontrol_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_tx_ucontrol_en_check ( .error(1'b1) );
		end
		if (pma_cgb_tx_ucontrol_pcie != "gen1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_tx_ucontrol_pcie_check ( .error(1'b1) );
		end
		if (pma_cgb_tx_ucontrol_reset != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_tx_ucontrol_reset_check ( .error(1'b1) );
		end
		if (pma_cgb_uc_cgb_vreg_boost != "no_voltage_boost")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_uc_cgb_vreg_boost_check ( .error(1'b1) );
		end
		if (pma_cgb_uc_vcc_setting != "vcc_setting2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_uc_vcc_setting_check ( .error(1'b1) );
		end
		if (pma_cgb_vccdreg_output != "vccdreg_nominal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_vccdreg_output_check ( .error(1'b1) );
		end
		if (pma_cgb_vreg_sel_ref != "sel_vccer_4ref")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_vreg_sel_ref_check ( .error(1'b1) );
		end
		if (pma_cgb_x1_div_m_sel != "divbypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_x1_div_m_sel_check ( .error(1'b1) );
		end
		if (pma_cgb_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_cgb_input_select_x1 != "fpll_bot")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_input_select_x1_check ( .error(1'b1) );
		end
		if (pma_cgb_input_select_gen3 != "not_used")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_input_select_gen3_check ( .error(1'b1) );
		end
		if (pma_cgb_input_select_xn != "not_used")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cgb_input_select_xn_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_analog_mode != "user_custom")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_analog_mode_check ( .error(1'b1) );
		end
		if (pma_tx_buf_bti_protected != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_bti_protected_check ( .error(1'b1) );
		end
		if (pma_tx_buf_calibration_en != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_calibration_en_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_calibration_en != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_calibration_en_check ( .error(1'b1) );
		end
		if (pma_tx_buf_calibration_resistor_value != "res_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_calibration_resistor_value_check ( .error(1'b1) );
		end
		if (pma_tx_buf_cdr_cp_calibration_en != "cdr_cp_cal_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_cdr_cp_calibration_en_check ( .error(1'b1) );
		end
		if (pma_tx_buf_chgpmp_current_dn_trim != "cp_current_trimming_dn_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_chgpmp_current_dn_trim_check ( .error(1'b1) );
		end
		if (pma_tx_buf_chgpmp_current_up_trim != "cp_current_trimming_up_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_chgpmp_current_up_trim_check ( .error(1'b1) );
		end
		if (pma_tx_buf_chgpmp_dn_trim_double != "normal_dn_trim_current")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_chgpmp_dn_trim_double_check ( .error(1'b1) );
		end
		if (pma_tx_buf_chgpmp_up_trim_double != "normal_up_trim_current")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_chgpmp_up_trim_double_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_clock_divider_ratio != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_clock_divider_ratio_check ( .error(1'b1) );
		end
		if (pma_tx_buf_compensation_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_compensation_en_check ( .error(1'b1) );
		end
		if (pma_tx_buf_compensation_posttap_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_compensation_posttap_en_check ( .error(1'b1) );
		end
		if (pma_tx_buf_cpen_ctrl != "cp_l1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_cpen_ctrl_check ( .error(1'b1) );
		end
		if (pma_tx_buf_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_datawidth != 64)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_datawidth_check ( .error(1'b1) );
		end
		if (pma_tx_buf_dcc_finestep_enin != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_dcc_finestep_enin_check ( .error(1'b1) );
		end
		if (pma_tx_buf_dcd_clk_div_ctrl != "dcd_ck_div128")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_dcd_clk_div_ctrl_check ( .error(1'b1) );
		end
		if (pma_tx_buf_dcd_detection_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_dcd_detection_en_check ( .error(1'b1) );
		end
		if (pma_tx_buf_dft_sel != "dft_disabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_dft_sel_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_correction_bandwidth != "dcc_bw_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_correction_bandwidth_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_correction_bandwidth_dn != "dcd_bw_dn_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_correction_bandwidth_dn_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_correction_reference1 != "dcc_ref1_4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_correction_reference1_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_correction_reference2 != "dcc_ref2_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_correction_reference2_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_correction_reset_n != "reset")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_correction_reset_n_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_cp_comp_en != "cp_comp_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_cp_comp_en_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_detector_cp_cal != "dcd_cp_cal_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_detector_cp_cal_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_detector_sa_cal != "dcd_sa_cal_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_detector_sa_cal_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_input_polarity != "dcc_input_pos")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_input_polarity_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_setting != "dcc_t32")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_setting_check ( .error(1'b1) );
		end
		if (pma_tx_buf_duty_cycle_setting_aux != "dcc2_t32")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_duty_cycle_setting_aux_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_gt_enabled != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_gt_enabled_check ( .error(1'b1) );
		end
		if (pma_tx_buf_idle_ctrl != "id_cpen_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_idle_ctrl_check ( .error(1'b1) );
		end
		if (pma_tx_buf_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_initial_settings_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_initial_settings_check ( .error(1'b1) );
		end
		if (pma_tx_buf_jtag_drv_sel != "drv1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_jtag_drv_sel_check ( .error(1'b1) );
		end
		if (pma_tx_buf_jtag_lp != "lp_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_jtag_lp_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_link != "sr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_link_check ( .error(1'b1) );
		end
		if (pma_tx_buf_low_power_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_low_power_en_check ( .error(1'b1) );
		end
		if (pma_tx_buf_lst != "atb_disabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_lst_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_rx_mcgb_location_for_pcie != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_rx_mcgb_location_for_pcie_check ( .error(1'b1) );
		end
		if (pma_tx_buf_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_optimal_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_optimal_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pcie_gen != "non_pcie")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pcie_gen_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_pma_tx_divclk_hz != "402832031")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_pma_tx_divclk_hz_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_power_mode != "high_perf")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_power_mode_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_power_rail_eht != 1800)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_power_rail_eht_check ( .error(1'b1) );
		end
		if (pma_tx_buf_power_rail_er != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_power_rail_er_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_power_rail_et != 1120)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_power_rail_et_check ( .error(1'b1) );
		end
		if (pma_tx_buf_powermode_ac_post_tap != "tx_post_tap_ac_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_powermode_ac_post_tap_check ( .error(1'b1) );
		end
		if (pma_tx_buf_powermode_ac_pre_tap != "tx_pre_tap_ac_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_powermode_ac_pre_tap_check ( .error(1'b1) );
		end
		if (pma_tx_buf_powermode_ac_tx_vod_no_jitcomp != "tx_vod_no_jitcomp_ac_l0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_powermode_ac_tx_vod_no_jitcomp_check ( .error(1'b1) );
		end
		if (pma_tx_buf_powermode_ac_tx_vod_w_jitcomp != "tx_vod_w_jitcomp_ac_l31")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_powermode_ac_tx_vod_w_jitcomp_check ( .error(1'b1) );
		end
		if (pma_tx_buf_powermode_dc_post_tap != "powerdown_tx_post_tap")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_powermode_dc_post_tap_check ( .error(1'b1) );
		end
		if (pma_tx_buf_powermode_dc_pre_tap != "powerdown_tx_pre_tap")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_powermode_dc_pre_tap_check ( .error(1'b1) );
		end
		if (pma_tx_buf_powermode_dc_tx_vod_no_jitcomp != "powerdown_tx_vod_no_jitcomp")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_powermode_dc_tx_vod_no_jitcomp_check ( .error(1'b1) );
		end
		if (pma_tx_buf_powermode_dc_tx_vod_w_jitcomp != "tx_vod_w_jitcomp_dc_l31")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_powermode_dc_tx_vod_w_jitcomp_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pre_emp_sign_1st_post_tap != "fir_post_1t_neg")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pre_emp_sign_1st_post_tap_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pre_emp_sign_pre_tap_1t != "fir_pre_1t_neg")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pre_emp_sign_pre_tap_1t_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pre_emp_switching_ctrl_1st_post_tap != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pre_emp_switching_ctrl_1st_post_tap_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pre_emp_switching_ctrl_pre_tap_1t != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pre_emp_switching_ctrl_pre_tap_1t_check ( .error(1'b1) );
		end
		if (pma_tx_buf_prot_mode != "basic_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_prot_mode_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_prot_mode != "basic_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_prot_mode_check ( .error(1'b1) );
		end
		if (pma_tx_buf_res_cal_local != "non_local")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_res_cal_local_check ( .error(1'b1) );
		end
		if (pma_tx_buf_rx_det != "mode_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_rx_det_check ( .error(1'b1) );
		end
		if (pma_tx_buf_rx_det_output_sel != "rx_det_pcie_out")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_rx_det_output_sel_check ( .error(1'b1) );
		end
		if (pma_tx_buf_rx_det_pdb != "rx_det_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_rx_det_pdb_check ( .error(1'b1) );
		end
		if (pma_tx_buf_sense_amp_offset_cal_curr_n != "sa_os_cal_in_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_sense_amp_offset_cal_curr_n_check ( .error(1'b1) );
		end
		if (pma_tx_buf_sense_amp_offset_cal_curr_p != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_sense_amp_offset_cal_curr_p_check ( .error(1'b1) );
		end
		if (pma_tx_buf_ser_powerdown != "normal_ser_on")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_ser_powerdown_check ( .error(1'b1) );
		end
		if (pma_tx_buf_slew_rate_ctrl != "slew_r5")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_slew_rate_ctrl_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_speed_grade != "e2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_speed_grade_check ( .error(1'b1) );
		end
		if (pma_tx_buf_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_sup_mode_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_sup_mode_check ( .error(1'b1) );
		end
		if (pma_tx_buf_swing_level != "hv")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_swing_level_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_swing_level != "hv")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_swing_level_check ( .error(1'b1) );
		end
		if (pma_tx_buf_term_code != "rterm_code7")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_term_code_check ( .error(1'b1) );
		end
		if (pma_tx_buf_term_n_tune != "rterm_n7")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_term_n_tune_check ( .error(1'b1) );
		end
		if (pma_tx_buf_term_p_tune != "rterm_p7")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_term_p_tune_check ( .error(1'b1) );
		end
		if (pma_tx_buf_term_sel != "r_r2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_term_sel_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_tile_type != "h")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_tile_type_check ( .error(1'b1) );
		end
		if (pma_tx_buf_tri_driver != "tri_driver_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_tri_driver_check ( .error(1'b1) );
		end
		if (pma_tx_buf_pm_cr2_tx_path_tx_pll_clk_hz != "12890625000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_pm_cr2_tx_path_tx_pll_clk_hz_check ( .error(1'b1) );
		end
		if (pma_tx_buf_tx_powerdown != "normal_tx_on")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_tx_powerdown_check ( .error(1'b1) );
		end
		if (pma_tx_buf_tx_rst_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_tx_rst_enable_check ( .error(1'b1) );
		end
		if (pma_tx_buf_xtx_path_xcgb_tx_ucontrol_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_xtx_path_xcgb_tx_ucontrol_en_check ( .error(1'b1) );
		end
		if (pma_tx_buf_uc_gen3 != "gen3_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_uc_gen3_check ( .error(1'b1) );
		end
		if (pma_tx_buf_uc_gen4 != "gen4_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_uc_gen4_check ( .error(1'b1) );
		end
		if (pma_tx_buf_uc_tx_cal != "uc_tx_cal_on")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_uc_tx_cal_check ( .error(1'b1) );
		end
		if (pma_tx_buf_uc_vcc_setting != "vcc_setting2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_uc_vcc_setting_check ( .error(1'b1) );
		end
		if (pma_tx_buf_user_fir_coeff_ctrl_sel != "ram_ctl")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_user_fir_coeff_ctrl_sel_check ( .error(1'b1) );
		end
		if (pma_tx_buf_vod_output_swing_ctrl != 31)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_vod_output_swing_ctrl_check ( .error(1'b1) );
		end
		if (pma_tx_buf_vreg_output != "vccdreg_nominal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_vreg_output_check ( .error(1'b1) );
		end
		if (pma_tx_buf_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_buf_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_tx_sequencer_tx_path_rstn_overrideb != "use_sequencer")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_sequencer_tx_path_rstn_overrideb_check ( .error(1'b1) );
		end
		if (pma_tx_sequencer_xtx_path_xcgb_tx_ucontrol_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_sequencer_xtx_path_xcgb_tx_ucontrol_en_check ( .error(1'b1) );
		end
		if (pma_tx_sequencer_xrx_path_uc_cal_clk_bypass != "cal_clk_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_sequencer_xrx_path_uc_cal_clk_bypass_check ( .error(1'b1) );
		end
		if (pma_tx_sequencer_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_sequencer_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_advanced_user_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_advanced_user_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_align_del != "align_del_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_align_del_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_ber_bit_err_total_cnt != "bit_err_total_cnt_10g")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_ber_bit_err_total_cnt_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_ber_clken != "ber_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_ber_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_ber_xus_timer_window != 19530)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_ber_xus_timer_window_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_bitslip_mode != "bitslip_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_bitslip_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_blksync_bitslip_type != "bitslip_comb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_blksync_bitslip_type_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_blksync_bitslip_wait_cnt != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_blksync_bitslip_wait_cnt_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_blksync_bitslip_wait_type != "bitslip_cnt")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_blksync_bitslip_wait_type_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_blksync_bypass != "blksync_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_blksync_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_blksync_clken != "blksync_clk_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_blksync_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt != "enum_invalid_sh_cnt_10g")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock != "knum_sh_cnt_postlock_10g")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock != "knum_sh_cnt_prelock_10g")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_blksync_pipeln != "blksync_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_blksync_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_clr_errblk_cnt_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_clr_errblk_cnt_en_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_control_del != "control_del_none")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_control_del_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_crcchk_bypass != "crcchk_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_crcchk_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_crcchk_clken != "crcchk_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_crcchk_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_crcchk_inv != "crcchk_inv_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_crcchk_inv_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_crcchk_pipeln != "crcchk_pipeln_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_crcchk_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_crcflag_pipeln != "crcflag_pipeln_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_crcflag_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_ctrl_bit_reverse != "ctrl_bit_reverse_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_ctrl_bit_reverse_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_data_bit_reverse != "data_bit_reverse_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_data_bit_reverse_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_dec64b66b_clken != "dec64b66b_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_dec64b66b_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass != "dec_64b66b_rxsm_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_descrm_bypass != "descrm_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_descrm_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_descrm_clken != "descrm_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_descrm_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_descrm_mode != "async")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_descrm_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_descrm_pipeln != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_descrm_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_dft_clk_out_sel != "rx_master_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_dft_clk_out_sel_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_dis_signal_ok != "dis_signal_ok_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_dis_signal_ok_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_dispchk_bypass != "dispchk_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_dispchk_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_empty_flag_type != "empty_rd_side")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_empty_flag_type_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_fast_path != "fast_path_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_fast_path_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_fec_clken != "fec_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_fec_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_fec_enable != "fec_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_fec_enable_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_fifo_double_read != "fifo_double_read_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_fifo_double_read_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_fifo_stop_rd != "n_rd_empty")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_fifo_stop_rd_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_fifo_stop_wr != "n_wr_full")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_fifo_stop_wr_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_force_align != "force_align_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_force_align_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_frmsync_bypass != "frmsync_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_frmsync_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_frmsync_clken != "frmsync_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_frmsync_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_frmsync_enum_scrm != "enum_scrm_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_frmsync_enum_scrm_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_frmsync_enum_sync != "enum_sync_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_frmsync_enum_sync_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_frmsync_flag_type != "location_only")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_frmsync_flag_type_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_frmsync_knum_sync != "knum_sync_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_frmsync_knum_sync_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_frmsync_mfrm_length != 2048)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_frmsync_mfrm_length_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_frmsync_pipeln != "frmsync_pipeln_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_frmsync_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_full_flag_type != "full_wr_side")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_full_flag_type_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_gb_rx_idwidth != "idwidth_64")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_gb_rx_idwidth_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_gb_rx_odwidth != "odwidth_66")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_gb_rx_odwidth_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_gbexp_clken != "gbexp_clk_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_gbexp_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_low_latency_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_low_latency_en_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_lpbk_mode != "lpbk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_lpbk_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_master_clk_sel != "master_rx_pma_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_master_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_pempty_flag_type != "pempty_rd_side")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_pempty_flag_type_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_pfull_flag_type != "pfull_wr_side")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_pfull_flag_type_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_phcomp_rd_del != "phcomp_rd_del2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_phcomp_rd_del_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_pld_if_type != "reg")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_pld_if_type_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_prot_mode != "basic_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rand_clken != "rand_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rand_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rd_clk_sel != "rd_rx_pma_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rd_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rdfifo_clken != "rdfifo_clk_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rdfifo_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rx_fifo_write_ctrl != "blklock_stops")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rx_fifo_write_ctrl_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rx_scrm_width != "bit64")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rx_scrm_width_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rx_sh_location != "msb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rx_sh_location_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rx_signal_ok_sel != "synchronized_ver")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rx_signal_ok_sel_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rx_sm_bypass != "rx_sm_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rx_sm_bypass_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rx_sm_hiber != "rx_sm_hiber_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rx_sm_hiber_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rx_sm_pipeln != "rx_sm_pipeln_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rx_sm_pipeln_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rx_testbus_sel != "rx_fifo_testbus1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rx_testbus_sel_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rx_true_b2b != "b2b")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rx_true_b2b_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rxfifo_empty != "empty_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rxfifo_empty_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rxfifo_full != "full_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rxfifo_full_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rxfifo_mode != "register_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rxfifo_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rxfifo_pempty != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rxfifo_pempty_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_rxfifo_pfull != 23)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_rxfifo_pfull_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_stretch_num_stages != "one_stage")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_stretch_num_stages_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_test_mode != "test_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_test_mode_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_wrfifo_clken != "wrfifo_clk_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_wrfifo_clken_check ( .error(1'b1) );
		end
		if (hssi_10g_rx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_10g_rx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_aib_clk1_sel != "aib_clk1_pld_pcs_rx_clk_out")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_aib_clk1_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_aib_clk2_sel != "aib_clk2_pld_pma_clkdiv_rx_user")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_aib_clk2_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_aib_fabric_pld_pma_hclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_aib_fabric_pld_pma_hclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_aib_fabric_rx_transfer_clk_hz != 805664062)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_aib_fabric_rx_transfer_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_asn_bypass_pma_pcie_sw_done != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_asn_bypass_pma_pcie_sw_done_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_asn_wait_for_dll_reset_cnt != 64)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_asn_wait_for_dll_reset_cnt_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_asn_wait_for_fifo_flush_cnt != 64)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_asn_wait_for_fifo_flush_cnt_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_asn_wait_for_pma_pcie_sw_done_cnt != 64)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_asn_wait_for_pma_pcie_sw_done_cnt_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_bonding_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_bonding_dft_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_bonding_dft_val != "dft_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_bonding_dft_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_chnl_bonding != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_chnl_bonding_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_clock_del_measure_enable != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_clock_del_measure_enable_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_csr_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_csr_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_ctrl_plane_bonding != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_ctrl_plane_bonding_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_ds_bypass_pipeln != "ds_bypass_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_ds_bypass_pipeln_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_duplex_mode != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_duplex_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_dv_mode != "dv_mode_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_dv_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_double_read != "fifo_double_read_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_double_read_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_mode != "generic_basic")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_rd_clk_ins_sm_scg_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_rd_clk_ins_sm_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_rd_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_rd_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_rd_clk_sel != "fifo_rd_clk_pld_rx_clk1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_rd_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_stop_rd != "n_rd_empty")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_stop_rd_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_stop_wr != "n_wr_full")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_stop_wr_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_width != "fifo_double_width")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_width_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_wr_clk_del_sm_scg_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_wr_clk_del_sm_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_wr_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_wr_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fifo_wr_clk_sel != "fifo_wr_clk_rx_transfer_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fifo_wr_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_free_run_div_clk != "out_of_reset_sync")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_free_run_div_clk_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fsr_pld_10g_rx_crc32_err_rst_val != "reset_to_zero_crc32")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fsr_pld_10g_rx_crc32_err_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fsr_pld_8g_sigdet_out_rst_val != "reset_to_zero_sigdet")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fsr_pld_8g_sigdet_out_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fsr_pld_ltd_b_rst_val != "reset_to_one_ltdb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fsr_pld_ltd_b_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fsr_pld_ltr_rst_val != "reset_to_zero_ltr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fsr_pld_ltr_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_fsr_pld_rx_fifo_align_clr_rst_val != "reset_to_zero_alignclr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_fsr_pld_rx_fifo_align_clr_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_gb_rx_idwidth != "idwidth_64")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_gb_rx_idwidth_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_gb_rx_odwidth != "odwidth_66")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_gb_rx_odwidth_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hip_mode != "disable_hip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hrdrst_align_bypass != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hrdrst_align_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hrdrst_dll_lock_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hrdrst_dll_lock_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hrdrst_rx_osc_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hrdrst_rx_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hrdrst_user_ctl_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hrdrst_user_ctl_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_indv != "indv_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_indv_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_internal_clk1_sel1 != "pma_clks_or_txfiford_post_ct_mux_clk1_mux1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_internal_clk1_sel1_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_internal_clk1_sel2 != "pma_clks_clk1_mux2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_internal_clk1_sel2_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_internal_clk2_sel1 != "pma_clks_or_rxfifowr_post_ct_mux_clk2_mux1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_internal_clk2_sel1_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_internal_clk2_sel2 != "pma_clks_clk2_mux2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_internal_clk2_sel2_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_loopback_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_loopback_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_low_latency_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_low_latency_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_lpbk_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_lpbk_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_osc_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_phcomp_rd_del != "phcomp_rd_del2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_phcomp_rd_del_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_pipe_enable != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_pipe_enable_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_pipe_mode != "disable_pipe")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_pipe_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_pld_avmm1_clk_rowclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_pld_avmm1_clk_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_pld_avmm2_clk_rowclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_pld_avmm2_clk_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_pld_clk1_delay_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_pld_clk1_delay_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_pld_clk1_delay_sel != "delay_path13")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_pld_clk1_delay_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_pld_clk1_inv_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_pld_clk1_inv_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_pld_clk1_sel != "pld_clk1_dcm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_pld_clk1_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_pld_rx_clk1_dcm_hz != 390625000)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_pld_rx_clk1_dcm_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_pld_rx_clk1_rowclk_hz != 390625000)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_pld_rx_clk1_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_pld_sclk1_rowclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_pld_sclk1_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_pld_sclk2_rowclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_pld_sclk2_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_pma_hclk_scg_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_pma_hclk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_powerdown_mode != "powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_powerdown_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_datapath_tb_sel != "cp_bond")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_datapath_tb_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_fastbond_rden != "rden_ds_fast_us_fast")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_fastbond_rden_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_fastbond_wren != "wren_ds_del_us_del")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_fastbond_wren_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_fifo_power_mode != "full_width_full_depth")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_fifo_power_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_fifo_read_latency_adjust != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_fifo_read_latency_adjust_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_fifo_write_ctrl != "blklock_ignore")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_fifo_write_ctrl_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_fifo_write_latency_adjust != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_fifo_write_latency_adjust_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_osc_clock_setting != "osc_clk_div_by1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_osc_clock_setting_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_pld_8g_eidleinfersel_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_pld_8g_eidleinfersel_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_pld_pma_eye_monitor_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_pld_pma_eye_monitor_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_pld_pma_pcie_switch_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_pld_pma_pcie_switch_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_pld_pma_reser_out_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_pld_pma_reser_out_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_prbs_flags_sr_enable != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_prbs_flags_sr_enable_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_true_b2b != "b2b")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_true_b2b_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rx_usertest_sel != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rx_usertest_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rxfifo_empty != "empty_dw")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rxfifo_empty_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rxfifo_full != "full_non_pc_dw")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rxfifo_full_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rxfifo_mode != "rxgeneric_basic")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rxfifo_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rxfifo_pempty != 13)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rxfifo_pempty_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rxfifo_pfull != 51)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rxfifo_pfull_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rxfiford_post_ct_sel != "rxfiford_sclk_post_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rxfiford_post_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_rxfifowr_post_ct_sel != "rxfifowr_sclk_post_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_rxfifowr_post_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_sclk_sel != "sclk1_rowclk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_sclk_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_hdpldadapt_speed_grade != "dash_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_hdpldadapt_speed_grade_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_stretch_num_stages != "two_stage")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_stretch_num_stages_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_txfiford_post_ct_sel != "txfiford_sclk_post_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_txfiford_post_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_txfifowr_post_ct_sel != "txfifowr_sclk_post_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_txfifowr_post_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_us_bypass_pipeln != "us_bypass_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_us_bypass_pipeln_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_word_align != "wa_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_word_align_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_word_align_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_word_align_enable_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_rx_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_rx_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_aib_clk1_sel != "aib_clk1_pld_pcs_tx_clk_out")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_aib_clk1_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_aib_clk2_sel != "aib_clk2_pld_pma_clkdiv_tx_user")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_aib_clk2_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_aib_fabric_pld_pma_hclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_aib_fabric_pld_pma_hclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz != 805664062)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_bonding_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_bonding_dft_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_bonding_dft_val != "dft_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_bonding_dft_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_chnl_bonding != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_chnl_bonding_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_csr_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_csr_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_ctrl_plane_bonding != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_ctrl_plane_bonding_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_ds_bypass_pipeln != "ds_bypass_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_ds_bypass_pipeln_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_duplex_mode != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_duplex_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_dv_bond != "dv_bond_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_dv_bond_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_dv_gen != "dv_gen_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_dv_gen_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fifo_double_write != "fifo_double_write_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fifo_double_write_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fifo_mode != "generic_basic")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fifo_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fifo_rd_clk_frm_gen_scg_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fifo_rd_clk_frm_gen_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fifo_rd_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fifo_rd_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fifo_rd_clk_sel != "fifo_rd_pma_aib_tx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fifo_rd_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fifo_stop_rd != "n_rd_empty")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fifo_stop_rd_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fifo_stop_wr != "n_wr_full")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fifo_stop_wr_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fifo_width != "fifo_double_width")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fifo_width_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fifo_wr_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fifo_wr_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fpll_shared_direct_async_in_sel != "fpll_shared_direct_async_in_rowclk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fpll_shared_direct_async_in_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_frmgen_burst != "frmgen_burst_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_frmgen_burst_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_frmgen_bypass != "frmgen_bypass_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_frmgen_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_frmgen_mfrm_length != 2048)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_frmgen_mfrm_length_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_frmgen_pipeln != "frmgen_pipeln_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_frmgen_pipeln_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_frmgen_pyld_ins != "frmgen_pyld_ins_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_frmgen_pyld_ins_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_frmgen_wordslip != "frmgen_wordslip_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_frmgen_wordslip_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_hip_fsr_in_bit0_rst_val != "reset_to_one_hfsrin0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_hip_fsr_in_bit0_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_hip_fsr_in_bit1_rst_val != "reset_to_one_hfsrin1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_hip_fsr_in_bit1_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_hip_fsr_in_bit2_rst_val != "reset_to_one_hfsrin2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_hip_fsr_in_bit2_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_hip_fsr_in_bit3_rst_val != "reset_to_zero_hfsrin3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_hip_fsr_in_bit3_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_hip_fsr_out_bit0_rst_val != "reset_to_one_hfsrout0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_hip_fsr_out_bit0_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_hip_fsr_out_bit1_rst_val != "reset_to_one_hfsrout1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_hip_fsr_out_bit1_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_hip_fsr_out_bit2_rst_val != "reset_to_zero_hfsrout2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_hip_fsr_out_bit2_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_hip_fsr_out_bit3_rst_val != "reset_to_zero_hfsrout3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_hip_fsr_out_bit3_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_mask_tx_pll_rst_val != "reset_to_zero_maskpll")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_mask_tx_pll_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_fsr_pld_txelecidle_rst_val != "reset_to_zero_txelec")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_fsr_pld_txelecidle_rst_val_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_gb_tx_idwidth != "idwidth_66")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_gb_tx_idwidth_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_gb_tx_odwidth != "odwidth_64")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_gb_tx_odwidth_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hip_mode != "disable_hip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hip_osc_clk_scg_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hip_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hrdrst_dcd_cal_done_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hrdrst_dcd_cal_done_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hrdrst_rx_osc_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hrdrst_rx_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hrdrst_user_ctl_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hrdrst_user_ctl_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_indv != "indv_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_indv_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_loopback_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_loopback_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_low_latency_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_low_latency_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_osc_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_phcomp_rd_del != "phcomp_rd_del2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_phcomp_rd_del_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_pipe_mode != "disable_pipe")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_pipe_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_pld_avmm1_clk_rowclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_pld_avmm1_clk_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_pld_avmm2_clk_rowclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_pld_avmm2_clk_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_pld_clk1_delay_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_pld_clk1_delay_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_pld_clk1_delay_sel != "delay_path15")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_pld_clk1_delay_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_pld_clk1_inv_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_pld_clk1_inv_en_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_pld_clk1_sel != "pld_clk1_dcm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_pld_clk1_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_pld_clk2_sel != "pld_clk2_dcm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_pld_clk2_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_pld_sclk1_rowclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_pld_sclk1_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_pld_sclk2_rowclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_pld_sclk2_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_pld_tx_clk1_dcm_hz != 390625000)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_pld_tx_clk1_dcm_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_pld_tx_clk1_rowclk_hz != 390625000)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_pld_tx_clk1_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_pld_tx_clk2_dcm_hz != 805664062)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_pld_tx_clk2_dcm_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_pld_tx_clk2_rowclk_hz != 805664062)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_pld_tx_clk2_rowclk_hz_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_pma_aib_tx_clk_expected_setting != "x2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_pma_aib_tx_clk_expected_setting_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_powerdown_mode != "powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_powerdown_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_sh_err != "sh_err_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_sh_err_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_hdpldadapt_speed_grade != "dash_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_hdpldadapt_speed_grade_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_stretch_num_stages != "two_stage")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_stretch_num_stages_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_datapath_tb_sel != "cp_bond")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_datapath_tb_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_fastbond_rden != "rden_ds_fast_us_fast")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_fastbond_rden_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_fastbond_wren != "wren_ds_fast_us_fast")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_fastbond_wren_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_fifo_power_mode != "full_width_full_depth")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_fifo_power_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_fifo_read_latency_adjust != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_fifo_read_latency_adjust_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_fifo_write_latency_adjust != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_fifo_write_latency_adjust_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_hip_aib_ssr_in_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_hip_aib_ssr_in_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_osc_clock_setting != "osc_clk_div_by1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_osc_clock_setting_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_pld_10g_tx_bitslip_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_pld_10g_tx_bitslip_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_pld_8g_tx_boundary_sel_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_pld_8g_tx_boundary_sel_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_pld_pma_fpll_cnt_sel_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_pld_pma_fpll_cnt_sel_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_pld_pma_fpll_num_phase_shifts_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_pld_pma_fpll_num_phase_shifts_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_tx_usertest_sel != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_tx_usertest_sel_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_txfifo_empty != "empty_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_txfifo_empty_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_txfifo_full != "full_non_pc_dw")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_txfifo_full_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_txfifo_mode != "txgeneric_basic")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_txfifo_mode_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_txfifo_pempty != 6)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_txfifo_pempty_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_txfifo_pfull != 26)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_txfifo_pfull_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_us_bypass_pipeln != "us_bypass_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_us_bypass_pipeln_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_word_align_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_word_align_enable_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_word_mark != "wm_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_word_mark_check ( .error(1'b1) );
		end
		if (hssi_pldadapt_tx_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pldadapt_tx_silicon_rev_check ( .error(1'b1) );
		end
		if (cdr_pll_analog_mode != "user_custom")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_analog_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_atb_select_control != "atb_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_atb_select_control_check ( .error(1'b1) );
		end
		if (cdr_pll_auto_reset_on != "auto_reset_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_auto_reset_on_check ( .error(1'b1) );
		end
		if (cdr_pll_bandwidth_range_high != "1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_bandwidth_range_high_check ( .error(1'b1) );
		end
		if (cdr_pll_bandwidth_range_low != "1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_bandwidth_range_low_check ( .error(1'b1) );
		end
		if (cdr_pll_bbpd_data_pattern_filter_select != "bbpd_data_pat_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_bbpd_data_pattern_filter_select_check ( .error(1'b1) );
		end
		if (cdr_pll_bti_protected != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_bti_protected_check ( .error(1'b1) );
		end
		if (cdr_pll_bw_mode != "mid_bw")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_bw_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_bypass_a_edge != "bypass_a_edge_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_bypass_a_edge_check ( .error(1'b1) );
		end
		if (cdr_pll_cal_vco_count_length != "sel_8b_count")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_cal_vco_count_length_check ( .error(1'b1) );
		end
		if (cdr_pll_pm_cr2_rx_path_cdr_clock_enable != "cdr_clock_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_pm_cr2_rx_path_cdr_clock_enable_check ( .error(1'b1) );
		end
		if (cdr_pll_cdr_d2a_enb != "bti_d2a_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_cdr_d2a_enb_check ( .error(1'b1) );
		end
		if (cdr_pll_cdr_odi_select != "sel_cdr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_cdr_odi_select_check ( .error(1'b1) );
		end
		if (cdr_pll_cdr_phaselock_mode != "no_ignore_lock")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_cdr_phaselock_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_cdr_powerdown_mode != "power_up")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_cdr_powerdown_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_current_dn_pd != "cp_current_pd_dn_setting4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_current_dn_pd_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_current_dn_trim != "cp_current_trimming_dn_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_current_dn_trim_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_current_pfd != "cp_current_pfd_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_current_pfd_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_current_up_pd != "cp_current_pd_up_setting4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_current_up_pd_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_current_up_trim != "cp_current_trimming_up_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_current_up_trim_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_dn_pd_trim_double != "normal_dn_trim_current")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_dn_pd_trim_double_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_replicate != "disable_replica_bias_ctrl")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_replicate_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_testmode != "cp_test_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_testmode_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_up_pd_trim_double != "normal_up_trim_current")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_up_pd_trim_double_check ( .error(1'b1) );
		end
		if (cdr_pll_chgpmp_vccreg != "vreg_fw0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_chgpmp_vccreg_check ( .error(1'b1) );
		end
		if (cdr_pll_clk0_dfe_tfall_adj != "clk0_dfe_tf0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_clk0_dfe_tfall_adj_check ( .error(1'b1) );
		end
		if (cdr_pll_clk0_dfe_trise_adj != "clk0_dfe_tr0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_clk0_dfe_trise_adj_check ( .error(1'b1) );
		end
		if (cdr_pll_clk180_dfe_tfall_adj != "clk180_dfe_tf0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_clk180_dfe_tfall_adj_check ( .error(1'b1) );
		end
		if (cdr_pll_clk180_dfe_trise_adj != "clk180_dfe_tr0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_clk180_dfe_trise_adj_check ( .error(1'b1) );
		end
		if (cdr_pll_clk270_dfe_tfall_adj != "clk270_dfe_tf0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_clk270_dfe_tfall_adj_check ( .error(1'b1) );
		end
		if (cdr_pll_clk270_dfe_trise_adj != "clk270_dfe_tr0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_clk270_dfe_trise_adj_check ( .error(1'b1) );
		end
		if (cdr_pll_clk90_dfe_tfall_adj != "clk90_dfe_tf0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_clk90_dfe_tfall_adj_check ( .error(1'b1) );
		end
		if (cdr_pll_clk90_dfe_trise_adj != "clk90_dfe_tr0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_clk90_dfe_trise_adj_check ( .error(1'b1) );
		end
		if (cdr_pll_clklow_mux_select != "clklow_mux_cdr_fbclk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_clklow_mux_select_check ( .error(1'b1) );
		end
		if (cdr_pll_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_datarate_bps_check ( .error(1'b1) );
		end
		if (cdr_pll_diag_loopback_enable != "no_diag_rev_loopback")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_diag_loopback_enable_check ( .error(1'b1) );
		end
		if (cdr_pll_disable_up_dn != "normal_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_disable_up_dn_check ( .error(1'b1) );
		end
		if (cdr_pll_f_max_cmu_out_freq != "1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_f_max_cmu_out_freq_check ( .error(1'b1) );
		end
		if (cdr_pll_f_max_m_counter != "1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_f_max_m_counter_check ( .error(1'b1) );
		end
		if (cdr_pll_f_max_pfd != "350000000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_f_max_pfd_check ( .error(1'b1) );
		end
		if (cdr_pll_f_max_ref != "800000000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_f_max_ref_check ( .error(1'b1) );
		end
		if (cdr_pll_f_max_vco != "14150000000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_f_max_vco_check ( .error(1'b1) );
		end
		if (cdr_pll_f_min_gt_channel != "8700000000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_f_min_gt_channel_check ( .error(1'b1) );
		end
		if (cdr_pll_f_min_pfd != "25000000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_f_min_pfd_check ( .error(1'b1) );
		end
		if (cdr_pll_f_min_ref != "25000000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_f_min_ref_check ( .error(1'b1) );
		end
		if (cdr_pll_f_min_vco != "7000000000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_f_min_vco_check ( .error(1'b1) );
		end
		if (cdr_pll_fref_clklow_div != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_fref_clklow_div_check ( .error(1'b1) );
		end
		if (cdr_pll_fref_mux_select != "fref_mux_cdr_refclk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_fref_mux_select_check ( .error(1'b1) );
		end
		if (cdr_pll_gpon_lck2ref_control != "gpon_lck2ref_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_gpon_lck2ref_control_check ( .error(1'b1) );
		end
		if (cdr_pll_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_initial_settings_check ( .error(1'b1) );
		end
		if (cdr_pll_lck2ref_delay_control != "lck2ref_delay_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_lck2ref_delay_control_check ( .error(1'b1) );
		end
		if (cdr_pll_lf_resistor_pd != "lf_pd_setting3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_lf_resistor_pd_check ( .error(1'b1) );
		end
		if (cdr_pll_lf_resistor_pfd != "lf_pfd_setting3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_lf_resistor_pfd_check ( .error(1'b1) );
		end
		if (cdr_pll_lf_ripple_cap != "lf_no_ripple")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_lf_ripple_cap_check ( .error(1'b1) );
		end
		if (cdr_pll_loop_filter_bias_select != "lpflt_bias_7")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_loop_filter_bias_select_check ( .error(1'b1) );
		end
		if (cdr_pll_loopback_mode != "loopback_disabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_loopback_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_lpd_counter != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_lpd_counter_check ( .error(1'b1) );
		end
		if (cdr_pll_lpfd_counter != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_lpfd_counter_check ( .error(1'b1) );
		end
		if (cdr_pll_ltd_ltr_micro_controller_select != "ltd_ltr_pcs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_ltd_ltr_micro_controller_select_check ( .error(1'b1) );
		end
		if (cdr_pll_mcnt_div != 20)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_mcnt_div_check ( .error(1'b1) );
		end
		if (cdr_pll_n_counter != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_n_counter_check ( .error(1'b1) );
		end
		if (cdr_pll_ncnt_div != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_ncnt_div_check ( .error(1'b1) );
		end
		if (cdr_pll_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_optimal_check ( .error(1'b1) );
		end
		if (cdr_pll_out_freq != "12890625000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_out_freq_check ( .error(1'b1) );
		end
		if (cdr_pll_pcie_gen != "non_pcie")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_pcie_gen_check ( .error(1'b1) );
		end
		if (cdr_pll_pd_fastlock_mode != "fast_lock_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_pd_fastlock_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_pd_l_counter != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_pd_l_counter_check ( .error(1'b1) );
		end
		if (cdr_pll_pfd_l_counter != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_pfd_l_counter_check ( .error(1'b1) );
		end
		if (cdr_pll_position != "position0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_position_check ( .error(1'b1) );
		end
		if (cdr_pll_power_mode != "high_perf")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_power_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_powermode_ac_bbpd != "bbpd_ac_on")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_powermode_ac_bbpd_check ( .error(1'b1) );
		end
		if (cdr_pll_powermode_ac_rvcotop != "rvcotop_ac_div1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_powermode_ac_rvcotop_check ( .error(1'b1) );
		end
		if (cdr_pll_powermode_ac_txpll != "txpll_ac_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_powermode_ac_txpll_check ( .error(1'b1) );
		end
		if (cdr_pll_powermode_dc_bbpd != "bbpd_dc_on")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_powermode_dc_bbpd_check ( .error(1'b1) );
		end
		if (cdr_pll_powermode_dc_rvcotop != "rvcotop_dc_div1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_powermode_dc_rvcotop_check ( .error(1'b1) );
		end
		if (cdr_pll_powermode_dc_txpll != "powerdown_txpll")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_powermode_dc_txpll_check ( .error(1'b1) );
		end
		if (cdr_pll_primary_use != "cdr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_primary_use_check ( .error(1'b1) );
		end
		if (cdr_pll_prot_mode != "basic_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_prot_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_reference_clock_frequency != "644531250")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_reference_clock_frequency_check ( .error(1'b1) );
		end
		if (cdr_pll_requires_gt_capable_channel != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_requires_gt_capable_channel_check ( .error(1'b1) );
		end
		if (cdr_pll_reverse_serial_loopback != "no_loopback")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_reverse_serial_loopback_check ( .error(1'b1) );
		end
		if (cdr_pll_set_cdr_input_freq_range != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_set_cdr_input_freq_range_check ( .error(1'b1) );
		end
		if (cdr_pll_set_cdr_v2i_enable != "enable_v2i_bias")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_set_cdr_v2i_enable_check ( .error(1'b1) );
		end
		if (cdr_pll_set_cdr_vco_reset != "vco_normal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_set_cdr_vco_reset_check ( .error(1'b1) );
		end
		if (cdr_pll_set_cdr_vco_speed != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_set_cdr_vco_speed_check ( .error(1'b1) );
		end
		if (cdr_pll_set_cdr_vco_speed_fix != 120)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_set_cdr_vco_speed_fix_check ( .error(1'b1) );
		end
		if (cdr_pll_set_cdr_vco_speed_pciegen3 != "cdr_vco_max_speedbin_pciegen3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_set_cdr_vco_speed_pciegen3_check ( .error(1'b1) );
		end
		if (cdr_pll_speed_grade != "e2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_speed_grade_check ( .error(1'b1) );
		end
		if (cdr_pll_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_sup_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_tx_pll_prot_mode != "txpll_unused")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_tx_pll_prot_mode_check ( .error(1'b1) );
		end
		if (cdr_pll_txpll_hclk_driver_enable != "hclk_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_txpll_hclk_driver_enable_check ( .error(1'b1) );
		end
		if (cdr_pll_rstb != "cdr_lf_reset_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_rstb_check ( .error(1'b1) );
		end
		if (cdr_pll_pm_cr2_tx_rx_uc_dyn_reconfig != "uc_dyn_reconfig_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_pm_cr2_tx_rx_uc_dyn_reconfig_check ( .error(1'b1) );
		end
		if (cdr_pll_uc_ro_cal != "uc_ro_cal_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_uc_ro_cal_check ( .error(1'b1) );
		end
		if (cdr_pll_vco_bypass != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_vco_bypass_check ( .error(1'b1) );
		end
		if (cdr_pll_vco_freq != "12890625000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_vco_freq_check ( .error(1'b1) );
		end
		if (cdr_pll_vco_overrange_voltage != "vco_overrange_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_vco_overrange_voltage_check ( .error(1'b1) );
		end
		if (cdr_pll_vco_underrange_voltage != "vco_underange_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_vco_underrange_voltage_check ( .error(1'b1) );
		end
		if (cdr_pll_vreg_output != "vccdreg_nominal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_vreg_output_check ( .error(1'b1) );
		end
		if (cdr_pll_direct_fb != "direct_fb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_direct_fb_check ( .error(1'b1) );
		end
		if (cdr_pll_iqclk_sel != "power_down")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_iqclk_sel_check ( .error(1'b1) );
		end
		if (cdr_pll_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_silicon_rev_check ( .error(1'b1) );
		end
		if (cdr_pll_pma_width != 64)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_pma_width_check ( .error(1'b1) );
		end
		if (cdr_pll_cgb_div != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_cgb_div_check ( .error(1'b1) );
		end
		if (cdr_pll_is_cascaded_pll != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cdr_pll_is_cascaded_pll_check ( .error(1'b1) );
		end
		if (pma_rx_buf_act_isource_disable != "isrc_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_act_isource_disable_check ( .error(1'b1) );
		end
		if (pma_rx_buf_advanced_mode != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_advanced_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_analog_mode != "user_custom")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_analog_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_bodybias_enable != "bodybias_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_bodybias_enable_check ( .error(1'b1) );
		end
		if (pma_rx_buf_bodybias_select != "bodybias_sel1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_bodybias_select_check ( .error(1'b1) );
		end
		if (pma_rx_buf_bypass_ctle_rf_cal != "use_dprio_rfcal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_bypass_ctle_rf_cal_check ( .error(1'b1) );
		end
		if (pma_rx_buf_clk_divrx_en != "normal_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_clk_divrx_en_check ( .error(1'b1) );
		end
		if (pma_rx_buf_const_gm_en != "cgm_en_1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_const_gm_en_check ( .error(1'b1) );
		end
		if (pma_rx_buf_ctle_ac_gain != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_ctle_ac_gain_check ( .error(1'b1) );
		end
		if (pma_rx_buf_ctle_eq_gain != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_ctle_eq_gain_check ( .error(1'b1) );
		end
		if (pma_rx_buf_ctle_hires_bypass != "ctle_hires_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_ctle_hires_bypass_check ( .error(1'b1) );
		end
		if (pma_rx_buf_ctle_oc_ib_sel != "ib_oc_bw3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_ctle_oc_ib_sel_check ( .error(1'b1) );
		end
		if (pma_rx_buf_ctle_oc_sign != "add_i_2_p_eq")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_ctle_oc_sign_check ( .error(1'b1) );
		end
		if (pma_rx_buf_ctle_rf_cal != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_ctle_rf_cal_check ( .error(1'b1) );
		end
		if (pma_rx_buf_ctle_tia_isel != "ib_tia_bw3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_ctle_tia_isel_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_tx_rx_cvp_mode != "cvp_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_tx_rx_cvp_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_datawidth != 64)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_datawidth_check ( .error(1'b1) );
		end
		if (pma_rx_buf_diag_lp_en != "dlp_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_diag_lp_en_check ( .error(1'b1) );
		end
		if (pma_rx_buf_eq_bw_sel != "eq_bw_3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_eq_bw_sel_check ( .error(1'b1) );
		end
		if (pma_rx_buf_eq_cdgen_sel != "eq_cdgen_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_eq_cdgen_sel_check ( .error(1'b1) );
		end
		if (pma_rx_buf_eq_isel != "eq_isel_1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_eq_isel_check ( .error(1'b1) );
		end
		if (pma_rx_buf_eq_sel != "eq_sel_3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_eq_sel_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_gt_enabled != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_gt_enabled_check ( .error(1'b1) );
		end
		if (pma_rx_buf_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_initial_settings_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_initial_settings_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_jtag_hys != "hys_increase_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_jtag_hys_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_jtag_lp != "lp_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_jtag_lp_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_link != "sr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_link_check ( .error(1'b1) );
		end
		if (pma_rx_buf_xrx_path_xcdr_deser_xcdr_loopback_mode != "loopback_disabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_xrx_path_xcdr_deser_xcdr_loopback_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_loopback_modes != "lpbk_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_loopback_modes_check ( .error(1'b1) );
		end
		if (pma_rx_buf_offset_cancellation_coarse != "coarse_setting_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_offset_cancellation_coarse_check ( .error(1'b1) );
		end
		if (pma_rx_buf_offset_rx_cal_en != "rx_oc_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_offset_rx_cal_en_check ( .error(1'b1) );
		end
		if (pma_rx_buf_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_optimal_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_optimal_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_tx_rx_pcie_gen != "non_pcie")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_tx_rx_pcie_gen_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_tx_rx_pcie_gen_bitwidth != "pcie_gen3_32b")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_tx_rx_pcie_gen_bitwidth_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pdb_rx != "normal_rx_on")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pdb_rx_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_pma_rx_divclk_hz != "402832031")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_pma_rx_divclk_hz_check ( .error(1'b1) );
		end
		if (pma_rx_buf_power_mode != "high_perf")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_power_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_power_mode != "high_perf")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_power_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_power_rail_eht != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_power_rail_eht_check ( .error(1'b1) );
		end
		if (pma_rx_buf_power_rail_er != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_power_rail_er_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_power_rail_er != 1120)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_power_rail_er_check ( .error(1'b1) );
		end
		if (pma_rx_buf_powermode_ac_ctle != "ctle_pwr_ac4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_powermode_ac_ctle_check ( .error(1'b1) );
		end
		if (pma_rx_buf_powermode_ac_vcm != "vcm_pwr_ac3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_powermode_ac_vcm_check ( .error(1'b1) );
		end
		if (pma_rx_buf_powermode_ac_vga != "vga_pwr_ac_full")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_powermode_ac_vga_check ( .error(1'b1) );
		end
		if (pma_rx_buf_powermode_dc_ctle != "ctle_pwr_dc1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_powermode_dc_ctle_check ( .error(1'b1) );
		end
		if (pma_rx_buf_powermode_dc_vcm != "vcm_pwr_dc3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_powermode_dc_vcm_check ( .error(1'b1) );
		end
		if (pma_rx_buf_powermode_dc_vga != "vga_pwr_dc_full")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_powermode_dc_vga_check ( .error(1'b1) );
		end
		if (pma_rx_buf_prot_mode != "basic_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_prot_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_prot_mode != "basic_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_prot_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_qpi_afe_en != "ctle_mode_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_qpi_afe_en_check ( .error(1'b1) );
		end
		if (pma_rx_buf_qpi_enable != "non_qpi_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_qpi_enable_check ( .error(1'b1) );
		end
		if (pma_rx_buf_refclk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_refclk_en_check ( .error(1'b1) );
		end
		if (pma_rx_buf_rx_atb_select != "atb_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_rx_atb_select_check ( .error(1'b1) );
		end
		if (pma_rx_buf_rx_vga_oc_en != "vga_cal_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_rx_vga_oc_en_check ( .error(1'b1) );
		end
		if (pma_rx_buf_sel_vcm_ctle != "vocm_eq_fixed")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_sel_vcm_ctle_check ( .error(1'b1) );
		end
		if (pma_rx_buf_sel_vcm_tia != "vocm_tia_fixed")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_sel_vcm_tia_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_speed_grade != "e2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_speed_grade_check ( .error(1'b1) );
		end
		if (pma_rx_buf_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_sup_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_sup_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_term_sel != "r_r4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_term_sel_check ( .error(1'b1) );
		end
		if (pma_rx_buf_term_sync_bypass != "bypass_termsync")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_term_sync_bypass_check ( .error(1'b1) );
		end
		if (pma_rx_buf_term_tri_enable != "disable_tri")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_term_tri_enable_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_tx_rx_testmux_select != "setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_tx_rx_testmux_select_check ( .error(1'b1) );
		end
		if (pma_rx_buf_tia_sel != "tia_sel_1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_tia_sel_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_tile_type != "h")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_tile_type_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_uc_cal_clk_bypass != "cal_clk_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_uc_cal_clk_bypass_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_uc_cal_enable != "rx_cal_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_uc_cal_enable_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_tx_rx_uc_odi_eye_left != "uc_odi_eye_left_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_tx_rx_uc_odi_eye_left_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_tx_rx_uc_odi_eye_right != "uc_odi_eye_right_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_tx_rx_uc_odi_eye_right_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_rx_path_uc_pcie_sw != "uc_pcie_gen1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_rx_path_uc_pcie_sw_check ( .error(1'b1) );
		end
		if (pma_rx_buf_pm_cr2_tx_rx_uc_rx_cal != "uc_rx_cal_on")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_pm_cr2_tx_rx_uc_rx_cal_check ( .error(1'b1) );
		end
		if (pma_rx_buf_vcm_cal_i != 4)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_vcm_cal_i_check ( .error(1'b1) );
		end
		if (pma_rx_buf_vcm_current_add != "vcm_current_3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_vcm_current_add_check ( .error(1'b1) );
		end
		if (pma_rx_buf_vcm_sel != "vcm_l0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_vcm_sel_check ( .error(1'b1) );
		end
		if (pma_rx_buf_vcm_sel_vccref != 6)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_vcm_sel_vccref_check ( .error(1'b1) );
		end
		if (pma_rx_buf_vga_dc_gain != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_vga_dc_gain_check ( .error(1'b1) );
		end
		if (pma_rx_buf_vga_halfbw_en != "vga_half_bw_disabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_vga_halfbw_en_check ( .error(1'b1) );
		end
		if (pma_rx_buf_vga_ib_max_en != "vga_ib_max_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_vga_ib_max_en_check ( .error(1'b1) );
		end
		if (pma_rx_buf_vga_mode != "vga_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_vga_mode_check ( .error(1'b1) );
		end
		if (pma_rx_buf_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_buf_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_adapter_lpbk_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_adapter_lpbk_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hd_hssiadapt_aib_hssi_pld_sclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hd_hssiadapt_aib_hssi_pld_sclk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_aib_lpbk_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_aib_lpbk_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_align_del != "align_del_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_align_del_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_asn_bypass_clock_gate != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_asn_bypass_clock_gate_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_asn_bypass_pma_pcie_sw_done != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_asn_bypass_pma_pcie_sw_done_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_asn_wait_for_clock_gate_cnt != 32)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_asn_wait_for_clock_gate_cnt_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_asn_wait_for_dll_reset_cnt != 32)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_asn_wait_for_dll_reset_cnt_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_asn_wait_for_fifo_flush_cnt != 32)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_asn_wait_for_fifo_flush_cnt_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_asn_wait_for_pma_pcie_sw_done_cnt != 32)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_asn_wait_for_pma_pcie_sw_done_cnt_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_async_direct_hip_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_async_direct_hip_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_bonding_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_bonding_dft_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_bonding_dft_val != "dft_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_bonding_dft_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_chnl_bonding != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_chnl_bonding_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_clock_del_measure_enable != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_clock_del_measure_enable_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_control_del != "control_del_none")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_control_del_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hd_hssiadapt_csr_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hd_hssiadapt_csr_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_ctrl_plane_bonding != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_ctrl_plane_bonding_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_datapath_mapping_mode != "map_10g_2x2x_2x1x_fifo")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_datapath_mapping_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_ds_bypass_pipeln != "ds_bypass_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_ds_bypass_pipeln_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_duplex_mode != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_duplex_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_dyn_clk_sw_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_dyn_clk_sw_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fifo_double_write != "fifo_double_write_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fifo_double_write_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fifo_mode != "phase_comp")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fifo_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fifo_rd_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fifo_rd_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fifo_rd_clk_sel != "fifo_rd_pma_aib_rx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fifo_rd_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fifo_stop_rd != "rd_empty")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fifo_stop_rd_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fifo_stop_wr != "n_wr_full")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fifo_stop_wr_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fifo_width != "fifo_double_width")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fifo_width_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fifo_wr_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fifo_wr_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fifo_wr_clk_sel != "fifo_wr_pld_pcs_rx_clk_out")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fifo_wr_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_force_align != "force_align_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_force_align_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_free_run_div_clk != "out_of_reset_sync")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_free_run_div_clk_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fsr_pld_10g_rx_crc32_err_rst_val != "reset_to_zero_crc32")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fsr_pld_10g_rx_crc32_err_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fsr_pld_8g_sigdet_out_rst_val != "reset_to_zero_sigdet")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fsr_pld_8g_sigdet_out_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fsr_pld_ltd_b_rst_val != "reset_to_one_ltdb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fsr_pld_ltd_b_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fsr_pld_ltr_rst_val != "reset_to_zero_ltr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fsr_pld_ltr_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_fsr_pld_rx_fifo_align_clr_rst_val != "reset_to_zero_alignclr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_fsr_pld_rx_fifo_align_clr_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hd_hssiadapt_hip_aib_clk_2x_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hd_hssiadapt_hip_aib_clk_2x_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hd_hssiadapt_hip_aib_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hd_hssiadapt_hip_aib_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hip_mode != "disable_hip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hrdrst_dcd_cal_done_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hrdrst_dcd_cal_done_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hrdrst_rx_osc_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hrdrst_rx_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hrdrst_user_ctl_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hrdrst_user_ctl_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_indv != "indv_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_indv_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk1_sel != "pld_pma_tx_clk_out_clk1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk1_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk1_sel0 != "pma_clks_or_txfifowr_post_ct_or_txfiford_pre_or_post_ct_mux_clk1_mux0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk1_sel0_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk1_sel1 != "pma_clks_or_txfiford_pre_or_post_ct_mux_clk1_mux1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk1_sel1_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk1_sel2 != "pma_clks_or_txfiford_pre_ct_mux_clk1_mux2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk1_sel2_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk1_sel3 != "pma_clks_clk1_mux3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk1_sel3_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk2_sel != "pld_pma_tx_clk_out_clk2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk2_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk2_sel0 != "pma_clks_or_rxfiford_post_ct_or_rxfifowr_pre_or_post_ct_mux_clk2_mux0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk2_sel0_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk2_sel1 != "pma_clks_or_rxfifowr_pre_or_post_ct_mux_clk2_mux1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk2_sel1_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk2_sel2 != "pma_clks_or_rxfifowr_pre_ct_mux_clk2_mux2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk2_sel2_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_internal_clk2_sel3 != "pma_clks_clk2_mux3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_internal_clk2_sel3_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_loopback_mode != "loopback_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_loopback_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_osc_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_phcomp_rd_del != "phcomp_rd_del3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_phcomp_rd_del_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_pipe_mode != "disable_pipe")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_pipe_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hd_hssiadapt_pld_pcs_rx_clk_out_hz != 402832031)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hd_hssiadapt_pld_pcs_rx_clk_out_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hd_hssiadapt_pld_pma_hclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hd_hssiadapt_pld_pma_hclk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_pma_aib_rx_clk_expected_setting != "x2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_pma_aib_rx_clk_expected_setting_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hd_hssiadapt_pma_aib_rx_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hd_hssiadapt_pma_aib_rx_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_pma_coreclkin_sel != "pma_coreclkin_pld_sel")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_pma_coreclkin_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_pma_hclk_scg_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_pma_hclk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_powerdown_mode != "powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_powerdown_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_10g_krfec_rx_diag_data_status_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_10g_krfec_rx_diag_data_status_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_adp_go_b4txeq_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_adp_go_b4txeq_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_datapath_tb_sel != "cp_bond")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_datapath_tb_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_eq_iteration != "cycles_32")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_eq_iteration_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_fifo_power_mode != "full_width_full_depth")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_fifo_power_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_fifo_read_latency_adjust != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_fifo_read_latency_adjust_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_fifo_write_latency_adjust != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_fifo_write_latency_adjust_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_invalid_no_change != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_invalid_no_change_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_osc_clock_setting != "osc_clk_div_by1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_osc_clock_setting_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_parity_sel != "func_sel")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_parity_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pcs_testbus_sel != "direct_tr_tb_bit0_sel")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pcs_testbus_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pcspma_testbus_sel != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pcspma_testbus_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pld_8g_a1a2_k1k2_flag_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pld_8g_a1a2_k1k2_flag_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pld_8g_wa_boundary_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pld_8g_wa_boundary_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pld_pma_pcie_sw_done_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pld_pma_pcie_sw_done_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pld_pma_reser_in_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pld_pma_reser_in_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pld_pma_testbus_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pld_pma_testbus_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pld_test_data_polling_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pld_test_data_polling_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pma_rstn_cycles != "four_cycles")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pma_rstn_cycles_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pma_rstn_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pma_rstn_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_post_cursor_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_post_cursor_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_pre_cursor_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_pre_cursor_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_rmfflag_stretch_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_rmfflag_stretch_enable_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_rmfflag_stretch_num_stages != "rmfflag_two_stage")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_rmfflag_stretch_num_stages_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_rxeq_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_rxeq_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_txeq_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_txeq_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_txeq_time != 64)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_txeq_time_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_use_rxvalid_for_rxeq != "rxvalid")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_use_rxvalid_for_rxeq_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rx_usertest_sel != "direct_tr_usertest3_sel")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rx_usertest_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rxfifo_empty != "empty_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rxfifo_empty_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rxfifo_full != "full_dw")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rxfifo_full_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rxfifo_mode != "rxphase_comp")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rxfifo_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rxfifo_pempty != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rxfifo_pempty_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rxfifo_pfull != 5)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rxfifo_pfull_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rxfiford_post_ct_sel != "rxfiford_sclk_post_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rxfiford_post_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rxfiford_to_aib_sel != "rxfiford_sclk_to_aib")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rxfiford_to_aib_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rxfifowr_post_ct_sel != "rxfifowr_sclk_post_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rxfifowr_post_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_rxfifowr_pre_ct_sel != "rxfifowr_sclk_pre_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_rxfifowr_pre_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_hd_hssiadapt_speed_grade != "dash_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_hd_hssiadapt_speed_grade_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_stretch_num_stages != "seven_stage")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_stretch_num_stages_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_txeq_clk_scg_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_txeq_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_txeq_clk_sel != "txeq_pld_pcs_rx_clk_out")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_txeq_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_txeq_mode != "eq_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_txeq_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_txeq_rst_sel != "txeq_pcs_rx_pld_rst_n")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_txeq_rst_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_txfiford_post_ct_sel != "txfiford_sclk_post_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_txfiford_post_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_txfiford_pre_ct_sel != "txfiford_sclk_pre_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_txfiford_pre_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_txfifowr_from_aib_sel != "txfifowr_sclk_from_aib")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_txfifowr_from_aib_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_txfifowr_post_ct_sel != "txfifowr_sclk_post_ct")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_txfifowr_post_ct_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_us_bypass_pipeln != "us_bypass_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_us_bypass_pipeln_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_word_align_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_word_align_enable_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_word_mark != "wm_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_word_mark_check ( .error(1'b1) );
		end
		if (hssi_adapt_rx_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_rx_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_reset_sequencer_rx_path_rstn_overrideb != "use_sequencer")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_reset_sequencer_rx_path_rstn_overrideb_check ( .error(1'b1) );
		end
		if (pma_reset_sequencer_xrx_path_uc_cal_clk_bypass != "cal_clk_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_reset_sequencer_xrx_path_uc_cal_clk_bypass_check ( .error(1'b1) );
		end
		if (pma_reset_sequencer_xrx_path_uc_cal_enable != "rx_cal_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_reset_sequencer_xrx_path_uc_cal_enable_check ( .error(1'b1) );
		end
		if (pma_reset_sequencer_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_reset_sequencer_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_tx_ser_bti_protected != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_bti_protected_check ( .error(1'b1) );
		end
		if (pma_tx_ser_control_clks_divtx_aibtx != "no_dft_control_clkdivtx_clkaibtx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_control_clks_divtx_aibtx_check ( .error(1'b1) );
		end
		if (pma_tx_ser_datarate_bps != "0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_tx_ser_duty_cycle_correction_mode_ctrl != "dcc_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_duty_cycle_correction_mode_ctrl_check ( .error(1'b1) );
		end
		if (pma_tx_ser_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_initial_settings_check ( .error(1'b1) );
		end
		if (pma_tx_ser_pcie_gen != "non_pcie")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_pcie_gen_check ( .error(1'b1) );
		end
		if (pma_tx_ser_power_rail_er != 1120)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_power_rail_er_check ( .error(1'b1) );
		end
		if (pma_tx_ser_powermode_ac_ser != "ac_clk_divtx_user_33_jitcomp1p1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_powermode_ac_ser_check ( .error(1'b1) );
		end
		if (pma_tx_ser_powermode_dc_ser != "dc_clk_divtx_user_33_jitcomp1p1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_powermode_dc_ser_check ( .error(1'b1) );
		end
		if (pma_tx_ser_prot_mode != "basic_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_prot_mode_check ( .error(1'b1) );
		end
		if (pma_tx_ser_ser_clk_divtx_user_sel != "divtx_user_33")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_ser_clk_divtx_user_sel_check ( .error(1'b1) );
		end
		if (pma_tx_ser_ser_aibck_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_ser_aibck_enable_check ( .error(1'b1) );
		end
		if (pma_tx_ser_ser_aibck_x1_override != "normal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_ser_aibck_x1_override_check ( .error(1'b1) );
		end
		if (pma_tx_ser_ser_clk_mon != "disable_clk_mon")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_ser_clk_mon_check ( .error(1'b1) );
		end
		if (pma_tx_ser_ser_dftppm_clkselect != "aib_dftppm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_ser_dftppm_clkselect_check ( .error(1'b1) );
		end
		if (pma_tx_ser_ser_in_jitcomp != "jitcomp_on")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_ser_in_jitcomp_check ( .error(1'b1) );
		end
		if (pma_tx_ser_ser_powerdown != "normal_poweron_ser")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_ser_powerdown_check ( .error(1'b1) );
		end
		if (pma_tx_ser_ser_preset_bti_en != "ser_preset_bti_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_ser_preset_bti_en_check ( .error(1'b1) );
		end
		if (pma_tx_ser_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_sup_mode_check ( .error(1'b1) );
		end
		if (pma_tx_ser_uc_vcc_setting != "vcc_setting2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_uc_vcc_setting_check ( .error(1'b1) );
		end
		if (pma_tx_ser_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_tx_ser_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_rx_deser_bitslip_bypass != "bs_bypass_yes")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_bitslip_bypass_check ( .error(1'b1) );
		end
		if (pma_rx_deser_bti_protected != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_bti_protected_check ( .error(1'b1) );
		end
		if (pma_rx_deser_clkdiv_source != "vco_bypass_normal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_clkdiv_source_check ( .error(1'b1) );
		end
		if (pma_rx_deser_clkdivrx_user_mode != "clkdivrx_user_div33")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_clkdivrx_user_mode_check ( .error(1'b1) );
		end
		if (pma_rx_deser_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_rx_deser_deser_aib_dftppm_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_deser_aib_dftppm_en_check ( .error(1'b1) );
		end
		if (pma_rx_deser_deser_aibck_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_deser_aibck_en_check ( .error(1'b1) );
		end
		if (pma_rx_deser_deser_aibck_x1 != "normal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_deser_aibck_x1_check ( .error(1'b1) );
		end
		if (pma_rx_deser_deser_factor != "deser_64b")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_deser_factor_check ( .error(1'b1) );
		end
		if (pma_rx_deser_deser_powerdown != "deser_power_up")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_deser_powerdown_check ( .error(1'b1) );
		end
		if (pma_rx_deser_force_adaptation_outputs != "normal_outputs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_force_adaptation_outputs_check ( .error(1'b1) );
		end
		if (pma_rx_deser_force_clkdiv_for_testing != "normal_clkdiv")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_force_clkdiv_for_testing_check ( .error(1'b1) );
		end
		if (pma_rx_deser_odi_adapt_bti_en != "deser_bti_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_odi_adapt_bti_en_check ( .error(1'b1) );
		end
		if (pma_rx_deser_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_optimal_check ( .error(1'b1) );
		end
		if (pma_rx_deser_pcie_g3_hclk_en != "disable_hclk_div2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_pcie_g3_hclk_en_check ( .error(1'b1) );
		end
		if (pma_rx_deser_pm_cr2_tx_rx_pcie_gen != "non_pcie")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_pm_cr2_tx_rx_pcie_gen_check ( .error(1'b1) );
		end
		if (pma_rx_deser_pm_cr2_tx_rx_pcie_gen_bitwidth != "pcie_gen3_32b")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_pm_cr2_tx_rx_pcie_gen_bitwidth_check ( .error(1'b1) );
		end
		if (pma_rx_deser_powermode_ac_deser != "deser_ac_64b_nobs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_powermode_ac_deser_check ( .error(1'b1) );
		end
		if (pma_rx_deser_powermode_ac_deser_bs != "deser_ac_bs_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_powermode_ac_deser_bs_check ( .error(1'b1) );
		end
		if (pma_rx_deser_powermode_dc_deser != "deser_dc_64b_nobs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_powermode_dc_deser_check ( .error(1'b1) );
		end
		if (pma_rx_deser_powermode_dc_deser_bs != "powerdown_deser_bs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_powermode_dc_deser_bs_check ( .error(1'b1) );
		end
		if (pma_rx_deser_prot_mode != "basic_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_prot_mode_check ( .error(1'b1) );
		end
		if (pma_rx_deser_rst_n_adapt_odi != "no_rst_adapt_odi")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_rst_n_adapt_odi_check ( .error(1'b1) );
		end
		if (pma_rx_deser_sd_clk != "sd_clk_disabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_sd_clk_check ( .error(1'b1) );
		end
		if (pma_rx_deser_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_sup_mode_check ( .error(1'b1) );
		end
		if (pma_rx_deser_tdr_mode != "select_bbpd_data")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_tdr_mode_check ( .error(1'b1) );
		end
		if (pma_rx_deser_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_deser_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_txpath_chnsequencer_pcie_gen != "non_pcie")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_txpath_chnsequencer_pcie_gen_check ( .error(1'b1) );
		end
		if (pma_txpath_chnsequencer_prot_mode != "basic_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_txpath_chnsequencer_prot_mode_check ( .error(1'b1) );
		end
		if (pma_txpath_chnsequencer_sup_mode != "sup_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_txpath_chnsequencer_sup_mode_check ( .error(1'b1) );
		end
		if (pma_txpath_chnsequencer_txpath_chnseq_enable != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_txpath_chnsequencer_txpath_chnseq_enable_check ( .error(1'b1) );
		end
		if (pma_txpath_chnsequencer_txpath_chnseq_idle_direct_on != "cgb_idle_direct_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_txpath_chnsequencer_txpath_chnseq_idle_direct_on_check ( .error(1'b1) );
		end
		if (pma_txpath_chnsequencer_txpath_chnseq_stage_select != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_txpath_chnsequencer_txpath_chnseq_stage_select_check ( .error(1'b1) );
		end
		if (pma_txpath_chnsequencer_txpath_chnseq_wakeup_bypass != "bypass_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_txpath_chnsequencer_txpath_chnseq_wakeup_bypass_check ( .error(1'b1) );
		end
		if (pma_txpath_chnsequencer_silicon_rev != "14nm5bcr2ea")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_txpath_chnsequencer_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_datasel_gr0 != "aib_datasel0_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_datasel_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_datasel_gr1 != "aib_datasel1_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_datasel_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_datasel_gr2 != "aib_datasel2_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_datasel_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_ddrctrl_gr0 != "aib_ddr0_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_ddrctrl_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_ddrctrl_gr1 != "aib_ddr1_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_ddrctrl_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_iinasyncen != "aib_inasyncen_setting2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_iinasyncen_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_iinclken != "aib_inclken_setting3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_iinclken_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outctrl_gr0 != "aib_outen0_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outctrl_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outctrl_gr1 != "aib_outen1_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outctrl_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outctrl_gr2 != "aib_outen2_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outctrl_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outctrl_gr3 != "aib_outen3_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outctrl_gr3_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outndrv_r12 != "aib_ndrv12_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outndrv_r12_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outndrv_r56 != "aib_ndrv56_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outndrv_r56_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outndrv_r78 != "aib_ndrv78_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outndrv_r78_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outpdrv_r12 != "aib_pdrv12_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outpdrv_r12_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outpdrv_r56 != "aib_pdrv56_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outpdrv_r56_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_outpdrv_r78 != "aib_pdrv78_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_outpdrv_r78_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_red_rx_shiften != "aib_red_rx_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_red_rx_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_clkdiv != "aib_rx_clkdiv_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_clkdiv_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_byp != "aib_rx_dcc_byp_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_byp_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_byp_iocsr_unused != "aib_rx_dcc_byp_disable_iocsr_unused")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_byp_iocsr_unused_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_cont_cal != "aib_rx_dcc_cal_cont")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_cont_cal_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_cont_cal_iocsr_unused != "aib_rx_dcc_cal_single_iocsr_unused")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_cont_cal_iocsr_unused_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_dft != "aib_rx_dcc_dft_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_dft_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_dft_sel != "aib_rx_dcc_dft_mode0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_dft_sel_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_dll_entest != "aib_rx_dcc_dll_test_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_dll_entest_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_dy_ctl_static != "aib_rx_dcc_dy_ctl_static_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_dy_ctl_static_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_dy_ctlsel != "aib_rx_dcc_dy_ctlsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_dy_ctlsel_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_en != "aib_rx_dcc_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_en_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_en_iocsr_unused != "aib_rx_dcc_disable_iocsr_unused")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_en_iocsr_unused_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_manual_dn != "aib_rx_dcc_manual_dn0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_manual_dn_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_manual_up != "aib_rx_dcc_manual_up0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_manual_up_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_rst_prgmnvrt != "aib_rx_dcc_st_rst_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_rst_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_core_dn_prgmnvrt != "aib_rx_dcc_st_core_dn_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_core_dn_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_core_up_prgmnvrt != "aib_rx_dcc_st_core_up_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_core_up_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_core_updnen != "aib_rx_dcc_st_core_updnen_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_core_updnen_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_dftmuxsel != "aib_rx_dcc_st_dftmuxsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_dftmuxsel_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_dly_pst != "aib_rx_dcc_st_dly_pst_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_dly_pst_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_en != "aib_rx_dcc_st_en_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_en_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_lockreq_muxsel != "aib_rx_dcc_st_lockreq_muxsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_lockreq_muxsel_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_new_dll != "aib_rx_dcc_new_dll_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_new_dll_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_new_dll2 != "aib_rx_dcc_new_dll2_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_new_dll2_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_st_rst != "aib_rx_dcc_st_rst_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_st_rst_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_dcc_test_clk_pll_en_n != "aib_rx_dcc_test_clk_pll_en_n_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_dcc_test_clk_pll_en_n_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_halfcode != "aib_rx_halfcode_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_halfcode_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_aib_rx_selflock != "aib_rx_selflock_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_aib_rx_selflock_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_dft_hssitestip_dll_dcc_en != "disable_dft")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_dft_hssitestip_dll_dcc_en_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_op_mode != "rx_dcc_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_op_mode_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_powermode_ac != "rxdatapath_high_speed_pwr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_powermode_ac_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_powermode_dc != "powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_powermode_dc_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_redundancy_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_redundancy_en_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_aibcr_rx_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_rx_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_datasel_gr0 != "aib_datasel0_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_datasel_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_datasel_gr1 != "aib_datasel1_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_datasel_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_datasel_gr2 != "aib_datasel2_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_datasel_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_clkdiv != "aib_dllstr_align_clkdiv_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_clkdiv_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_dcc_dll_dft_sel != "aib_dllstr_align_dcc_dll_dft_sel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_dcc_dll_dft_sel_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_dft_ch_muxsel != "aib_dllstr_align_dft_ch_muxsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_dft_ch_muxsel_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_dly_pst != "aib_dllstr_align_dly_pst_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_dly_pst_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_dy_ctl_static != "aib_dllstr_align_dy_ctl_static_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_dy_ctl_static_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_dy_ctlsel != "aib_dllstr_align_dy_ctlsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_dy_ctlsel_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_entest != "aib_dllstr_align_test_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_entest_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_halfcode != "aib_dllstr_align_halfcode_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_halfcode_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_selflock != "aib_dllstr_align_selflock_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_selflock_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_core_dn_prgmnvrt != "aib_dllstr_align_st_core_dn_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_core_dn_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_core_up_prgmnvrt != "aib_dllstr_align_st_core_up_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_core_up_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_core_updnen != "aib_dllstr_align_st_core_updnen_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_core_updnen_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_dftmuxsel != "aib_dllstr_align_st_dftmuxsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_dftmuxsel_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_en != "aib_dllstr_align_st_en_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_en_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_lockreq_muxsel != "aib_dllstr_align_st_lockreq_muxsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_lockreq_muxsel_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_new_dll != "aib_dllstr_align_new_dll_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_new_dll_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_new_dll2 != "aib_dllstr_align_new_dll2_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_new_dll2_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_rst != "aib_dllstr_align_st_rst_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_rst_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_st_rst_prgmnvrt != "aib_dllstr_align_st_rst_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_st_rst_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_dllstr_align_test_clk_pll_en_n != "aib_dllstr_align_test_clk_pll_en_n_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_dllstr_align_test_clk_pll_en_n_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_inctrl_gr0 != "aib_inctrl0_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_inctrl_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_inctrl_gr1 != "aib_inctrl1_setting3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_inctrl_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_inctrl_gr2 != "aib_inctrl2_setting2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_inctrl_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_inctrl_gr3 != "aib_inctrl3_setting2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_inctrl_gr3_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outctrl_gr0 != "aib_outen0_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outctrl_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outctrl_gr1 != "aib_outen1_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outctrl_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outctrl_gr2 != "aib_outen2_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outctrl_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outndrv_r12 != "aib_ndrv12_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outndrv_r12_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outndrv_r34 != "aib_ndrv34_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outndrv_r34_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outndrv_r56 != "aib_ndrv56_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outndrv_r56_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outndrv_r78 != "aib_ndrv78_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outndrv_r78_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outpdrv_r12 != "aib_pdrv12_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outpdrv_r12_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outpdrv_r34 != "aib_pdrv34_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outpdrv_r34_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outpdrv_r56 != "aib_pdrv56_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outpdrv_r56_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_outpdrv_r78 != "aib_pdrv78_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_outpdrv_r78_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_red_dirclkn_shiften != "aib_red_dirclkn_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_red_dirclkn_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_red_dirclkp_shiften != "aib_red_dirclkp_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_red_dirclkp_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_red_drx_shiften != "aib_red_drx_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_red_drx_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_red_dtx_shiften != "aib_red_dtx_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_red_dtx_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_red_pinp_shiften != "aib_red_pinp_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_red_pinp_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_red_rx_shiften != "aib_red_rx_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_red_rx_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_red_tx_shiften != "aib_red_tx_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_red_tx_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_red_txferclkout_shiften != "aib_red_txferclkout_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_red_txferclkout_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_aib_red_txferclkoutn_shiften != "aib_red_txferclkoutn_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_aib_red_txferclkoutn_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_dfd_dll_dcc_en != "disable_dfd")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_dfd_dll_dcc_en_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_dft_hssitestip_dll_dcc_en != "disable_dft")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_dft_hssitestip_dll_dcc_en_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_op_mode != "tx_dll_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_op_mode_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_powermode_ac != "txdatapath_high_speed_pwr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_powermode_ac_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_powermode_dc != "powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_powermode_dc_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_redundancy_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_redundancy_en_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_aibcr_tx_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibcr_tx_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_datasel_gr0 != "aib_datasel0_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_datasel_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_datasel_gr1 != "aib_datasel1_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_datasel_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_datasel_gr2 != "aib_datasel2_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_datasel_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_clkdiv != "aib_dllstr_align_clkdiv_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_clkdiv_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_dly_pst != "aib_dllstr_align_dly_pst_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_dly_pst_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_dy_ctl_static != "aib_dllstr_align_dy_ctl_static_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_dy_ctl_static_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_dy_ctlsel != "aib_dllstr_align_dy_ctlsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_dy_ctlsel_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_entest != "aib_dllstr_align_test_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_entest_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_halfcode != "aib_dllstr_align_halfcode_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_halfcode_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_selflock != "aib_dllstr_align_selflock_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_selflock_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_core_dn_prgmnvrt != "aib_dllstr_align_st_core_dn_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_core_dn_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_core_up_prgmnvrt != "aib_dllstr_align_st_core_up_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_core_up_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_core_updnen != "aib_dllstr_align_st_core_updnen_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_core_updnen_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_dftmuxsel != "aib_dllstr_align_st_dftmuxsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_dftmuxsel_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_en != "aib_dllstr_align_st_en_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_hps_ctrl_en != "aib_dllstr_align_hps_ctrl_en_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_hps_ctrl_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_lockreq_muxsel != "aib_dllstr_align_st_lockreq_muxsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_lockreq_muxsel_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_new_dll != "aib_dllstr_align_new_dll_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_new_dll_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_rst != "aib_dllstr_align_st_rst_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_rst_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_st_rst_prgmnvrt != "aib_dllstr_align_st_rst_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_st_rst_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_dllstr_align_test_clk_pll_en_n != "aib_dllstr_align_test_clk_pll_en_n_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_dllstr_align_test_clk_pll_en_n_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_inctrl_gr0 != "aib_inctrl0_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_inctrl_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_inctrl_gr1 != "aib_inctrl1_setting3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_inctrl_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_inctrl_gr2 != "aib_inctrl2_setting2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_inctrl_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_inctrl_gr3 != "aib_inctrl3_setting3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_inctrl_gr3_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outctrl_gr0 != "aib_outen0_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outctrl_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outctrl_gr1 != "aib_outen1_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outctrl_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outctrl_gr2 != "aib_outen2_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outctrl_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outndrv_r12 != "aib_ndrv12_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outndrv_r12_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outndrv_r34 != "aib_ndrv34_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outndrv_r34_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outndrv_r56 != "aib_ndrv56_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outndrv_r56_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outndrv_r78 != "aib_ndrv78_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outndrv_r78_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outpdrv_r12 != "aib_pdrv12_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outpdrv_r12_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outpdrv_r34 != "aib_pdrv34_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outpdrv_r34_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outpdrv_r56 != "aib_pdrv56_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outpdrv_r56_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_outpdrv_r78 != "aib_pdrv78_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_outpdrv_r78_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_aib_red_shift_en != "aib_red_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_aib_red_shift_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_dft_hssitestip_dll_dcc_en != "disable_dft")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_dft_hssitestip_dll_dcc_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_op_mode != "rx_dll_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_op_mode_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_powermode_ac != "rxdatapath_high_speed_pwr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_powermode_ac_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_powermode_dc != "rxdatapath_powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_powermode_dc_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_redundancy_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_redundancy_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_aibnd_rx_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_rx_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_datasel_gr0 != "aib_datasel0_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_datasel_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_datasel_gr1 != "aib_datasel1_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_datasel_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_datasel_gr2 != "aib_datasel2_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_datasel_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_datasel_gr3 != "aib_datasel3_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_datasel_gr3_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_ddrctrl_gr0 != "aib_ddr0_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_ddrctrl_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_iinasyncen != "aib_inasyncen_setting2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_iinasyncen_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_iinclken != "aib_inclken_setting3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_iinclken_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_outctrl_gr0 != "aib_outen0_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_outctrl_gr0_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_outctrl_gr1 != "aib_outen1_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_outctrl_gr1_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_outctrl_gr2 != "aib_outen2_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_outctrl_gr2_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_outctrl_gr3 != "aib_outen3_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_outctrl_gr3_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_outndrv_r34 != "aib_ndrv34_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_outndrv_r34_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_outndrv_r56 != "aib_ndrv56_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_outndrv_r56_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_outpdrv_r34 != "aib_pdrv34_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_outpdrv_r34_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_outpdrv_r56 != "aib_pdrv56_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_outpdrv_r56_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_red_dirclkn_shiften != "aib_red_dirclkn_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_red_dirclkn_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_red_dirclkp_shiften != "aib_red_dirclkp_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_red_dirclkp_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_red_drx_shiften != "aib_red_drx_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_red_drx_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_red_dtx_shiften != "aib_red_dtx_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_red_dtx_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_red_pout_shiften != "aib_red_pout_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_red_pout_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_red_rx_shiften != "aib_red_rx_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_red_rx_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_red_tx_shiften != "aib_red_tx_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_red_tx_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_red_txferclkout_shiften != "aib_red_txferclkout_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_red_txferclkout_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_red_txferclkoutn_shiften != "aib_red_txferclkoutn_shift_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_red_txferclkoutn_shiften_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_clkdiv != "aib_tx_clkdiv_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_clkdiv_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_byp != "aib_tx_dcc_byp_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_byp_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_byp_iocsr_unused != "aib_tx_dcc_byp_disable_iocsr_unused")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_byp_iocsr_unused_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_cont_cal != "aib_tx_dcc_cal_cont")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_cont_cal_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_cont_cal_iocsr_unused != "aib_tx_dcc_cal_single_iocsr_unused")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_cont_cal_iocsr_unused_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_dft != "aib_tx_dcc_dft_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_dft_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_dft_sel != "aib_tx_dcc_dft_mode0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_dft_sel_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_dll_dft_sel != "aib_tx_dcc_dll_dft_sel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_dll_dft_sel_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_dll_entest != "aib_tx_dcc_dll_test_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_dll_entest_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_dy_ctl_static != "aib_tx_dcc_dy_ctl_static_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_dy_ctl_static_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_dy_ctlsel != "aib_tx_dcc_dy_ctlsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_dy_ctlsel_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_en != "aib_tx_dcc_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_en_iocsr_unused != "aib_tx_dcc_disable_iocsr_unused")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_en_iocsr_unused_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_manual_dn != "aib_tx_dcc_manual_dn0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_manual_dn_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_manual_up != "aib_tx_dcc_manual_up0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_manual_up_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_rst_prgmnvrt != "aib_tx_dcc_st_rst_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_rst_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_core_dn_prgmnvrt != "aib_tx_dcc_st_core_dn_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_core_dn_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_core_up_prgmnvrt != "aib_tx_dcc_st_core_up_prgmnvrt_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_core_up_prgmnvrt_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_core_updnen != "aib_tx_dcc_st_core_updnen_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_core_updnen_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_dftmuxsel != "aib_tx_dcc_st_dftmuxsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_dftmuxsel_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_dly_pst != "aib_tx_dcc_st_dly_pst_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_dly_pst_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_en != "aib_tx_dcc_st_en_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_hps_ctrl_en != "aib_tx_dcc_hps_ctrl_en_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_hps_ctrl_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_lockreq_muxsel != "aib_tx_dcc_st_lockreq_muxsel_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_lockreq_muxsel_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_new_dll != "aib_tx_dcc_new_dll_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_new_dll_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_st_rst != "aib_tx_dcc_st_rst_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_st_rst_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_dcc_test_clk_pll_en_n != "aib_tx_dcc_test_clk_pll_en_n_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_dcc_test_clk_pll_en_n_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_halfcode != "aib_tx_halfcode_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_halfcode_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_aib_tx_selflock != "aib_tx_selflock_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_aib_tx_selflock_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_dfd_dll_dcc_en != "disable_dfd")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_dfd_dll_dcc_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_dft_hssitestip_dll_dcc_en != "disable_dft")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_dft_hssitestip_dll_dcc_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_op_mode != "tx_dcc_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_op_mode_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_powermode_ac != "txdatapath_high_speed_pwr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_powermode_ac_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_powermode_dc != "txdatapath_powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_powermode_dc_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_redundancy_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_redundancy_en_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_aibnd_tx_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_aibnd_tx_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_bypass_rx_detection_enable != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_bypass_rx_detection_enable_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_bypass_rx_preset != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_bypass_rx_preset_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_bypass_rx_preset_enable != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_bypass_rx_preset_enable_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_bypass_tx_coefficent != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_bypass_tx_coefficent_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_bypass_tx_coefficent_enable != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_bypass_tx_coefficent_enable_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_elecidle_delay_g3 != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_elecidle_delay_g3_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_ind_error_reporting != "dis_ind_error_reporting")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_ind_error_reporting_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_mode != "disable_pcs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_mode_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_phy_status_delay_g12 != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_phy_status_delay_g12_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_phy_status_delay_g3 != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_phy_status_delay_g3_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_phystatus_rst_toggle_g12 != "dis_phystatus_rst_toggle")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_phystatus_rst_toggle_g12_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_phystatus_rst_toggle_g3 != "dis_phystatus_rst_toggle_g3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_phystatus_rst_toggle_g3_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_rate_match_pad_insertion != "dis_rm_fifo_pad_ins")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_rate_match_pad_insertion_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_test_out_sel != "disable_test_out")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_test_out_sel_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen3_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen3_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_block_sync != "bypass_block_sync")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_block_sync_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_block_sync_sm != "disable_blk_sync_sm")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_block_sync_sm_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_lpbk_force != "lpbk_frce_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_lpbk_force_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_mode != "disable_pcs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_mode_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_rate_match_fifo != "bypass_rm_fifo")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_rate_match_fifo_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_rate_match_fifo_latency != "low_latency")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_rate_match_fifo_latency_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_reverse_lpbk != "rev_lpbk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_reverse_lpbk_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_rx_b4gb_par_lpbk != "b4gb_par_lpbk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_rx_b4gb_par_lpbk_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_rx_force_balign != "dis_force_balign")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_rx_force_balign_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_rx_ins_del_one_skip != "ins_del_one_skip_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_rx_ins_del_one_skip_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_rx_num_fixed_pat != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_rx_num_fixed_pat_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_rx_test_out_sel != "rx_test_out0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_rx_test_out_sel_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_gen3_rx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_rx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_gen3_tx_pcs_mode != "disable_pcs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_tx_pcs_mode_check ( .error(1'b1) );
		end
		if (hssi_gen3_tx_pcs_reverse_lpbk != "rev_lpbk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_tx_pcs_reverse_lpbk_check ( .error(1'b1) );
		end
		if (hssi_gen3_tx_pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_tx_pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_gen3_tx_pcs_tx_bitslip != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_tx_pcs_tx_bitslip_check ( .error(1'b1) );
		end
		if (hssi_gen3_tx_pcs_tx_gbox_byp != "bypass_gbox")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_tx_pcs_tx_gbox_byp_check ( .error(1'b1) );
		end
		if (hssi_gen3_tx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_gen3_tx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_aib_clk_sel != "aib_clk_pma_aib_tx_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_aib_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_aib_hssi_pld_sclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_aib_hssi_pld_sclk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_aib_hssi_tx_transfer_clk_hz != 805664062)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_aib_hssi_tx_transfer_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_bonding_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_bonding_dft_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_bonding_dft_val != "dft_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_bonding_dft_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_chnl_bonding != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_chnl_bonding_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_csr_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_csr_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_ctrl_plane_bonding != "individual")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_ctrl_plane_bonding_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_datapath_mapping_mode != "map_10g_2x2x_2x1x_fifo")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_datapath_mapping_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_ds_bypass_pipeln != "ds_bypass_pipeln_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_ds_bypass_pipeln_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_duplex_mode != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_duplex_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_dv_gating != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_dv_gating_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_dyn_clk_sw_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_dyn_clk_sw_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fifo_double_read != "fifo_double_read_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fifo_double_read_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fifo_mode != "phase_comp")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fifo_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fifo_rd_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fifo_rd_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fifo_rd_clk_sel != "fifo_rd_pld_pcs_tx_clk_out")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fifo_rd_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fifo_ready_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fifo_ready_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fifo_stop_rd != "rd_empty")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fifo_stop_rd_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fifo_stop_wr != "wr_full")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fifo_stop_wr_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fifo_width != "fifo_double_width")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fifo_width_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fifo_wr_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fifo_wr_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_free_run_div_clk != "out_of_reset_sync")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_free_run_div_clk_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_hip_fsr_in_bit0_rst_val != "reset_to_one_hfsrin0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_hip_fsr_in_bit0_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_hip_fsr_in_bit1_rst_val != "reset_to_one_hfsrin1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_hip_fsr_in_bit1_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_hip_fsr_in_bit2_rst_val != "reset_to_one_hfsrin2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_hip_fsr_in_bit2_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_hip_fsr_in_bit3_rst_val != "reset_to_zero_hfsrin3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_hip_fsr_in_bit3_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_hip_fsr_out_bit0_rst_val != "reset_to_one_hfsrout0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_hip_fsr_out_bit0_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_hip_fsr_out_bit1_rst_val != "reset_to_one_hfsrout1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_hip_fsr_out_bit1_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_hip_fsr_out_bit2_rst_val != "reset_to_zero_hfsrout2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_hip_fsr_out_bit2_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_hip_fsr_out_bit3_rst_val != "reset_to_zero_hfsrout3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_hip_fsr_out_bit3_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_mask_tx_pll_rst_val != "reset_to_zero_maskpll")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_mask_tx_pll_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_fsr_pld_txelecidle_rst_val != "reset_to_zero_txelec")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_fsr_pld_txelecidle_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_hip_aib_clk_2x_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_hip_aib_clk_2x_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_hip_aib_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_hip_aib_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_hip_aib_txeq_clk_out_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_hip_aib_txeq_clk_out_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hip_mode != "disable_hip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hip_osc_clk_scg_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hip_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hrdrst_align_bypass != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hrdrst_align_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hrdrst_dcd_cal_done_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hrdrst_dcd_cal_done_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hrdrst_dll_lock_bypass != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hrdrst_dll_lock_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hrdrst_rx_osc_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hrdrst_rx_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hrdrst_user_ctl_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hrdrst_user_ctl_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_indv != "indv_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_indv_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_loopback_mode != "loopback_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_loopback_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_osc_clk_scg_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_osc_clk_scg_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_phcomp_rd_del != "phcomp_rd_del2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_phcomp_rd_del_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_pipe_mode != "disable_pipe")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_pipe_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_pld_pcs_tx_clk_out_hz != 402832031)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_pld_pcs_tx_clk_out_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_pld_pma_hclk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_pld_pma_hclk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_pma_aib_tx_clk_expected_setting != "x2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_pma_aib_tx_clk_expected_setting_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_pma_aib_tx_clk_hz != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_pma_aib_tx_clk_hz_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_powerdown_mode != "powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_powerdown_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_presethint_bypass != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_presethint_bypass_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_qpi_sr_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_qpi_sr_enable_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_rxqpi_pullup_rst_val != "reset_to_zero_rxqpi")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_rxqpi_pullup_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_hd_hssiadapt_speed_grade != "dash_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_hd_hssiadapt_speed_grade_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_stretch_num_stages != "seven_stage")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_stretch_num_stages_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_tx_datapath_tb_sel != "cp_bond")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_tx_datapath_tb_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_tx_fastbond_wren != "wren_ds_del2_us_del2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_tx_fastbond_wren_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_tx_fifo_power_mode != "full_width_full_depth")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_tx_fifo_power_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_tx_fifo_read_latency_adjust != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_tx_fifo_read_latency_adjust_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_tx_fifo_write_latency_adjust != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_tx_fifo_write_latency_adjust_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_tx_osc_clock_setting != "osc_clk_div_by1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_tx_osc_clock_setting_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_tx_qpi_mode_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_tx_qpi_mode_en_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_tx_rev_lpbk != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_tx_rev_lpbk_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_tx_usertest_sel != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_tx_usertest_sel_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_txfifo_empty != "empty_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_txfifo_empty_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_txfifo_full != "full_dw")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_txfifo_full_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_txfifo_mode != "txphase_comp")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_txfifo_mode_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_txfifo_pempty != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_txfifo_pempty_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_txfifo_pfull != 5)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_txfifo_pfull_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_txqpi_pulldn_rst_val != "reset_to_zero_txqpid")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_txqpi_pulldn_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_txqpi_pullup_rst_val != "reset_to_zero_txqpiu")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_txqpi_pullup_rst_val_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_word_align != "wa_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_word_align_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_word_align_enable != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_word_align_enable_check ( .error(1'b1) );
		end
		if (hssi_adapt_tx_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_adapt_tx_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_blksync_cor_en != "detect")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_blksync_cor_en_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_bypass_gb != "bypass_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_bypass_gb_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_clr_ctrl != "both_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_clr_ctrl_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_ctrl_bit_reverse != "ctrl_bit_reverse_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_ctrl_bit_reverse_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_data_bit_reverse != "data_bit_reverse_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_data_bit_reverse_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_dv_start != "with_blklock")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_dv_start_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_err_mark_type != "err_mark_10g")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_err_mark_type_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_error_marking_en != "err_mark_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_error_marking_en_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_low_latency_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_low_latency_en_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_lpbk_mode != "lpbk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_lpbk_mode_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_parity_invalid_enum != 8)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_parity_invalid_enum_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_parity_valid_num != 4)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_parity_valid_num_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_blksync != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_blksync_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_descrm != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_descrm_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_errcorrect != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_errcorrect_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_errtrap_ind != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_errtrap_ind_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_errtrap_lfsr != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_errtrap_lfsr_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_errtrap_loc != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_errtrap_loc_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_errtrap_pat != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_errtrap_pat_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_gearbox != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_gearbox_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_syndrm != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_syndrm_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_pipeln_trans_dec != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_pipeln_trans_dec_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_prot_mode != "disable_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_receive_order != "receive_lsb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_receive_order_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_rx_testbus_sel != "overall")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_rx_testbus_sel_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_signal_ok_en != "sig_ok_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_signal_ok_en_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_krfec_rx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_rx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_burst_err != "burst_err_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_burst_err_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_burst_err_len != "burst_err_len1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_burst_err_len_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_ctrl_bit_reverse != "ctrl_bit_reverse_en")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_ctrl_bit_reverse_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_data_bit_reverse != "data_bit_reverse_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_data_bit_reverse_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_enc_frame_query != "enc_query_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_enc_frame_query_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_low_latency_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_low_latency_en_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_pipeln_encoder != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_pipeln_encoder_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_pipeln_scrambler != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_pipeln_scrambler_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_prot_mode != "disable_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_transcode_err != "trans_err_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_transcode_err_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_transmit_order != "transmit_lsb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_transmit_order_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_tx_testbus_sel != "overall")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_tx_testbus_sel_check ( .error(1'b1) );
		end
		if (hssi_krfec_tx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_krfec_tx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_elec_idle_delay_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_elec_idle_delay_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_error_replace_pad != "replace_edb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_error_replace_pad_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_hip_mode != "dis_hip")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_ind_error_reporting != "dis_ind_error_reporting")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_ind_error_reporting_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_phystatus_delay_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_phystatus_delay_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_phystatus_rst_toggle != "dis_phystatus_rst_toggle")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_phystatus_rst_toggle_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_pipe_byte_de_serializer_en != "dont_care_bds")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_pipe_byte_de_serializer_en_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_prot_mode != "disabled_prot_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rpre_emph_a_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rpre_emph_a_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rpre_emph_b_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rpre_emph_b_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rpre_emph_c_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rpre_emph_c_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rpre_emph_d_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rpre_emph_d_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rpre_emph_e_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rpre_emph_e_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rvod_sel_a_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rvod_sel_a_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rvod_sel_b_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rvod_sel_b_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rvod_sel_c_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rvod_sel_c_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rvod_sel_d_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rvod_sel_d_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rvod_sel_e_val != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rvod_sel_e_val_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rx_pipe_enable != "dis_pipe_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rx_pipe_enable_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_rxdetect_bypass != "dis_rxdetect_bypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_rxdetect_bypass_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_tx_pipe_enable != "dis_pipe_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_tx_pipe_enable_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_txswing != "dis_txswing")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_txswing_check ( .error(1'b1) );
		end
		if (hssi_pipe_gen1_2_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pipe_gen1_2_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_common_pld_pcs_interface_dft_clk_out_en != "dft_clk_out_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pld_pcs_interface_dft_clk_out_en_check ( .error(1'b1) );
		end
		if (hssi_common_pld_pcs_interface_dft_clk_out_sel != "teng_rx_dft_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pld_pcs_interface_dft_clk_out_sel_check ( .error(1'b1) );
		end
		if (hssi_common_pld_pcs_interface_hrdrstctrl_en != "hrst_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pld_pcs_interface_hrdrstctrl_en_check ( .error(1'b1) );
		end
		if (hssi_common_pld_pcs_interface_pcs_testbus_block_sel != "pma_if")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pld_pcs_interface_pcs_testbus_block_sel_check ( .error(1'b1) );
		end
		if (hssi_common_pld_pcs_interface_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pld_pcs_interface_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_asn_clk_enable != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_asn_clk_enable_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_asn_enable != "dis_asn")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_asn_enable_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_block_sel != "eight_g_pcs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_block_sel_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_bypass_early_eios != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_bypass_early_eios_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_bypass_pcie_switch != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_bypass_pcie_switch_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_bypass_pma_ltr != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_bypass_pma_ltr_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_bypass_ppm_lock != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_bypass_ppm_lock_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_bypass_txdetectrx != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_bypass_txdetectrx_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_cdr_control != "dis_cdr_ctrl")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_cdr_control_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_cid_enable != "dis_cid_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_cid_enable_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_data_mask_count != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_data_mask_count_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_data_mask_count_multi != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_data_mask_count_multi_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_dft_observation_clock_selection != "dft_clk_obsrv_tx0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_dft_observation_clock_selection_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_early_eios_counter != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_early_eios_counter_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_force_freqdet != "force_freqdet_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_force_freqdet_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_free_run_clk_enable != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_free_run_clk_enable_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_ignore_sigdet_g23 != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_ignore_sigdet_g23_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_pc_en_counter != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_pc_en_counter_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_pc_rst_counter != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_pc_rst_counter_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_pcie_hip_mode != "hip_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_pcie_hip_mode_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_ph_fifo_reg_mode != "phfifo_reg_mode_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_ph_fifo_reg_mode_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_phfifo_flush_wait != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_phfifo_flush_wait_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_pipe_if_g3pcs != "pipe_if_8gpcs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_pipe_if_g3pcs_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_pma_done_counter != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_pma_done_counter_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_pma_if_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_pma_if_dft_en_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_pma_if_dft_val != "dft_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_pma_if_dft_val_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_ppm_cnt_rst != "ppm_cnt_rst_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_ppm_cnt_rst_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_ppm_deassert_early != "deassert_early_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_ppm_deassert_early_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_ppm_det_buckets != "ppm_300_100_bucket")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_ppm_det_buckets_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_ppm_gen1_2_cnt != "cnt_32k")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_ppm_gen1_2_cnt_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_ppm_post_eidle_delay != "cnt_200_cycles")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_ppm_post_eidle_delay_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_ppmsel != "ppmsel_1000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_ppmsel_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_prot_mode != "other_protocols")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_rxvalid_mask != "rxvalid_mask_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_rxvalid_mask_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_sigdet_wait_counter != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_sigdet_wait_counter_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_sigdet_wait_counter_multi != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_sigdet_wait_counter_multi_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_sim_mode != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_sim_mode_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_testout_sel != "ppm_det_test")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_testout_sel_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_wait_clk_on_off_timer != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_wait_clk_on_off_timer_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_wait_pipe_synchronizing != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_wait_pipe_synchronizing_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_wait_send_syncp_fbkp != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_wait_send_syncp_fbkp_check ( .error(1'b1) );
		end
		if (hssi_common_pcs_pma_interface_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_common_pcs_pma_interface_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_block_sel != "ten_g_pcs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_block_sel_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_clkslip_sel != "pld")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_clkslip_sel_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_master_clk_sel != "master_rx_pma_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_master_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_pldif_datawidth_mode != "pldif_data_10bit")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_pldif_datawidth_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_pma_dw_rx != "pma_64b_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_pma_dw_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_pma_if_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_pma_if_dft_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_pma_if_dft_val != "dft_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_pma_if_dft_val_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_prbs9_dwidth != "prbs9_64b")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_prbs9_dwidth_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_prbs_clken != "prbs_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_prbs_clken_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_prbs_ver != "prbs_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_prbs_ver_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_prot_mode_rx != "teng_basic_mode_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_prot_mode_rx_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion != "rx_dyn_polinv_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_rx_lpbk_en != "lpbk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_rx_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok != "force_sig_ok")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_rx_prbs_mask != "prbsmask128")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_rx_prbs_mask_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_rx_prbs_mode != "teng_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_rx_prbs_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel != "sel_sig_det")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_rx_static_polarity_inversion != "rx_stat_polinv_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_rx_static_polarity_inversion_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en != "uhsif_lpbk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_rx_pcs_pma_interface_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_rx_pcs_pma_interface_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_bypass_pma_txelecidle != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_bypass_pma_txelecidle_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_channel_operation_mode != "tx_rx_pair_enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_channel_operation_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_lpbk_en != "disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_lpbk_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_master_clk_sel != "master_tx_pma_clk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_master_clk_sel_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx != "other_prot_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_pldif_datawidth_mode != "pldif_data_10bit")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_pldif_datawidth_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_pma_dw_tx != "pma_64b_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_pma_dw_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_pma_if_dft_en != "dft_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_pma_if_dft_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_pmagate_en != "pmagate_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_pmagate_en_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_prbs9_dwidth != "prbs9_64b")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_prbs9_dwidth_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_prbs_clken != "prbs_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_prbs_clken_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_prbs_gen_pat != "prbs_gen_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_prbs_gen_pat_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_prot_mode_tx != "teng_basic_mode_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_prot_mode_tx_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_sq_wave_num != "sq_wave_default")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_sq_wave_num_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_sqwgen_clken != "sqwgen_clk_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_sqwgen_clken_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_sup_mode_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion != "tx_dyn_polinv_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_tx_pma_data_sel != "ten_g_pcs")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_tx_pma_data_sel_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_tx_static_polarity_inversion != "tx_stat_polinv_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_tx_static_polarity_inversion_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock != "uhsif_filt_stepsz_b4lock_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock != "uhsif_filt_cntthr_b4lock_8")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period != "uhsif_dcn_test_period_4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable != "uhsif_dcn_test_mode_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh != "uhsif_dzt_cnt_thr_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable != "uhsif_dzt_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window != "uhsif_dzt_obr_win_16")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size != "uhsif_dzt_skipsz_4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel != "uhsif_index_cram")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin != "uhsif_dcn_margin_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control != "uhsif_dft_dz_det_val_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control != "uhsif_dft_up_val_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_enable != "uhsif_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_enable_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock != "uhsif_lkd_segsz_aflock_512")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock != "uhsif_lkd_segsz_b4lock_16")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value_check ( .error(1'b1) );
		end
		if (hssi_tx_pcs_pma_interface_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_tx_pcs_pma_interface_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_fifo_rx_pcs_double_read_mode != "double_read_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_fifo_rx_pcs_double_read_mode_check ( .error(1'b1) );
		end
		if (hssi_fifo_rx_pcs_prot_mode != "teng_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_fifo_rx_pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_fifo_rx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_fifo_rx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_fifo_tx_pcs_double_write_mode != "double_write_dis")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_fifo_tx_pcs_double_write_mode_check ( .error(1'b1) );
		end
		if (hssi_fifo_tx_pcs_prot_mode != "teng_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_fifo_tx_pcs_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_fifo_tx_pcs_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_fifo_tx_pcs_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_cdr_refclk_powerdown_mode != "powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cdr_refclk_powerdown_mode_check ( .error(1'b1) );
		end
		if (pma_cdr_refclk_receiver_detect_src != "iqclk_src")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cdr_refclk_receiver_detect_src_check ( .error(1'b1) );
		end
		if (pma_cdr_refclk_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cdr_refclk_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_cdr_refclk_refclk_select != "ref_iqclk0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_cdr_refclk_refclk_select_check ( .error(1'b1) );
		end
		if (pma_rx_odi_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_rx_odi_enable_cdr_lpbk != "disable_lpbk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_enable_cdr_lpbk_check ( .error(1'b1) );
		end
		if (pma_rx_odi_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_initial_settings_check ( .error(1'b1) );
		end
		if (pma_rx_odi_monitor_bw_sel != "bw_1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_monitor_bw_sel_check ( .error(1'b1) );
		end
		if (pma_rx_odi_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_optimal_check ( .error(1'b1) );
		end
		if (pma_rx_odi_phase_steps_64_vs_128 != "phase_steps_64")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_phase_steps_64_vs_128_check ( .error(1'b1) );
		end
		if (pma_rx_odi_phase_steps_sel != "step40")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_phase_steps_sel_check ( .error(1'b1) );
		end
		if (pma_rx_odi_power_mode != "high_perf")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_power_mode_check ( .error(1'b1) );
		end
		if (pma_rx_odi_prot_mode != "basic_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_prot_mode_check ( .error(1'b1) );
		end
		if (pma_rx_odi_xrx_path_x119_rx_path_rstn_overrideb != "use_sequencer")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_xrx_path_x119_rx_path_rstn_overrideb_check ( .error(1'b1) );
		end
		if (pma_rx_odi_step_ctrl_sel != "dprio_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_step_ctrl_sel_check ( .error(1'b1) );
		end
		if (pma_rx_odi_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_sup_mode_check ( .error(1'b1) );
		end
		if (pma_rx_odi_vert_threshold != "vert_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_vert_threshold_check ( .error(1'b1) );
		end
		if (pma_rx_odi_vreg_voltage_sel != "vreg3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_vreg_voltage_sel_check ( .error(1'b1) );
		end
		if (pma_rx_odi_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_odi_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_adapt_sequencer_rx_path_rstn_overrideb != "use_sequencer")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_sequencer_rx_path_rstn_overrideb_check ( .error(1'b1) );
		end
		if (pma_adapt_sequencer_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_sequencer_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_adapt_adapt_mode != "ctle_dfe")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adapt_mode_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ac_ctle_cal_win != "radp_ac_ctle_cal_win_4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ac_ctle_cal_win_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ac_ctle_cocurrent_mode_sel != "radp_ac_ctle_cocurrent_mode_sel_mode_1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ac_ctle_cocurrent_mode_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ac_ctle_en != "radp_ac_ctle_en_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ac_ctle_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ac_ctle_hold_en != "radp_ac_ctle_hold_en_not_hold")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ac_ctle_hold_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ac_ctle_initial_load != "radp_ac_ctle_initial_load_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ac_ctle_initial_load_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ac_ctle_initial_value != "radp_ac_ctle_initial_value_8")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ac_ctle_initial_value_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ac_ctle_mode_sel != "radp_ac_ctle_mode_sel_concurrent")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ac_ctle_mode_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ac_ctle_ph1_win != "radp_ac_ctle_ph1_win_2p19")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ac_ctle_ph1_win_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_adapt_control_sel != "radp_adapt_control_sel_from_cram")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_adapt_control_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_adapt_start != "radp_adapt_start_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_adapt_start_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_bist_datapath_en != "radp_bist_datapath_en_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_bist_datapath_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_bist_errcount_rstn != "radp_bist_errcount_rstn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_bist_errcount_rstn_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_bist_mode_sel != "radp_bist_mode_sel_prbs31")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_bist_mode_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_clkgate_enb != "radp_clkgate_enb_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_clkgate_enb_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_clkout_div_sel != "radp_clkout_div_sel_div2_4cycle")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_clkout_div_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ctle_bypass_ac != "radp_ctle_bypass_ac_not_bypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ctle_bypass_ac_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_ctle_bypass_dc != "radp_ctle_bypass_dc_not_bypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_ctle_bypass_dc_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_accum_depth != 8)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_accum_depth_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_en != "radp_dc_ctle_en_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_hold_en != "radp_dc_ctle_hold_en_not_hold")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_hold_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_initial_load != "radp_dc_ctle_initial_load_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_initial_load_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_initial_value != "radp_dc_ctle_initial_value_32")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_initial_value_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_mode0_win_size != "radp_dc_ctle_mode0_win_size_4_taps")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_mode0_win_size_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_mode0_win_start != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_mode0_win_start_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_mode1_h1_ratio != 8)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_mode1_h1_ratio_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_mode2_h2_limit != 7)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_mode2_h2_limit_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_mode_sel != "radp_dc_ctle_mode_sel_mode_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_mode_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_onetime != "radp_dc_ctle_onetime_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_onetime_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dc_ctle_onetime_threshold != "radp_dc_ctle_onetime_threshold_256")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dc_ctle_onetime_threshold_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_accum_depth != 8)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_accum_depth_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_en != "radp_dfe_en_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_fxtap_bypass != "radp_dfe_fxtap_bypass_not_bypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_fxtap_bypass_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_hold_en != "radp_dfe_hold_en_not_hold")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_hold_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_hold_sel != "radp_dfe_hold_sel_no")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_hold_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_onetime != "radp_dfe_onetime_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_onetime_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_onetime_threshold != "radp_dfe_onetime_threshold_2048")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_onetime_threshold_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_tap1_initial_load != "radp_dfe_tap1_initial_load_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_tap1_initial_load_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_tap1_initial_value != "radp_dfe_tap1_initial_value_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_tap1_initial_value_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dfe_tap_sel_en != "radp_dfe_tap_sel_en_no")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dfe_tap_sel_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dlev_accum_depth != 6)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dlev_accum_depth_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dlev_bypass != "radp_dlev_bypass_not_bypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dlev_bypass_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dlev_en != "radp_dlev_en_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dlev_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dlev_hold_en != "radp_dlev_hold_en_not_hold")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dlev_hold_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dlev_initial_load != "radp_dlev_initial_load_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dlev_initial_load_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dlev_initial_value != "radp_dlev_initial_value_38")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dlev_initial_value_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dlev_onetime != "radp_dlev_onetime_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dlev_onetime_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dlev_onetime_threshold != "radp_dlev_onetime_threshold_4096")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dlev_onetime_threshold_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_dlev_sel != "radp_dlev_sel_mux")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_dlev_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_force_freqlock != "radp_force_freqlock_use")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_force_freqlock_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_frame_capture != "radp_frame_capture_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_frame_capture_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_frame_en != "radp_frame_en_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_frame_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_frame_odi_sel != "radp_frame_odi_sel_deser_err")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_frame_odi_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_frame_out_sel != "radp_frame_out_sel_select_a")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_frame_out_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_load_sig_sel != "radp_load_sig_sel_from_interanl")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_load_sig_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_oc_accum_depth != 11)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_oc_accum_depth_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_oc_bypass != "radp_oc_bypass_bypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_oc_bypass_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_oc_en != "radp_oc_en_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_oc_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_oc_hold_en != "radp_oc_hold_en_not_hold")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_oc_hold_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_oc_initial_load != "radp_oc_initial_load_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_oc_initial_load_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_oc_initial_sign != "radp_oc_initial_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_oc_initial_sign_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_oc_onetime != "radp_oc_onetime_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_oc_onetime_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_oc_onetime_threshold != "radp_oc_onetime_threshold_1024")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_oc_onetime_threshold_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_bit_sel != "radp_odi_bit_sel_all_bits")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_bit_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_control_sel != "radp_odi_control_sel_from_cram")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_control_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_count_threshold != "radp_odi_count_threshold_1e6")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_count_threshold_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_dfe_spec_en != "radp_odi_dfe_spec_en_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_dfe_spec_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_dlev_sel != "radp_odi_dlev_sel_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_dlev_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_en != "radp_odi_en_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_mode != "radp_odi_mode_detect_errdata")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_mode_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_rstn != "radp_odi_rstn_1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_rstn_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_spec_sel != "radp_odi_spec_sel_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_spec_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_odi_start != "radp_odi_start_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_odi_start_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pat_dlev_sign_avg_win != "radp_pat_dlev_sign_avg_win_2x")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pat_dlev_sign_avg_win_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pat_dlev_sign_force != "radp_pat_dlev_sign_force_determined_by_cram")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pat_dlev_sign_force_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pat_dlev_sign_value != "radp_pat_dlev_sign_value_1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pat_dlev_sign_value_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pat_spec_sign_avg_win != "radp_pat_spec_sign_avg_win_256")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pat_spec_sign_avg_win_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pat_spec_sign_force != "radp_pat_spec_sign_force_generated_internally")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pat_spec_sign_force_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pat_spec_sign_value != "radp_pat_spec_sign_value_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pat_spec_sign_value_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pat_trans_filter != "radp_pat_trans_filter_5")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pat_trans_filter_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pat_trans_only_en != "radp_pat_trans_only_en_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pat_trans_only_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pcie_adp_bypass != "radp_pcie_adp_bypass_no")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pcie_adp_bypass_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pcie_eqz != "radp_pcie_eqz_non_pcie_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pcie_eqz_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pcie_hold_sel != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pcie_hold_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_pcs_option != "radp_pcs_option_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_pcs_option_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_po_actslp_ratio != "radp_po_actslp_ratio_10_percent")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_po_actslp_ratio_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_po_en != "radp_po_en_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_po_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_po_gb_act2slp != "radp_po_gb_act2slp_288ns")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_po_gb_act2slp_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_po_gb_slp2act != "radp_po_gb_slp2act_288ns")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_po_gb_slp2act_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_po_initwait != "radp_po_initwait_10sec")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_po_initwait_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_po_sleep_win != "radp_po_sleep_win_2_sec")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_po_sleep_win_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_reserved != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_reserved_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_rstn != "radp_rstn_1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_rstn_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_status_sel != "radp_status_sel_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_status_sel_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_tx_accum_depth != 4)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_tx_accum_depth_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_tx_adp_accumulate != "radp_tx_adp_accumulate_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_tx_adp_accumulate_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_tx_adp_en != "radp_tx_adp_en_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_tx_adp_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_tx_up_dn_flip != "radp_tx_up_dn_flip_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_tx_up_dn_flip_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_accum_depth != 9)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_accum_depth_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_bypass != "radp_vga_bypass_not_bypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_bypass_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_ctle_low_limit != "radp_vga_ctle_low_limit_4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_ctle_low_limit_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_dlev_offset != 4)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_dlev_offset_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_dlev_target != 25)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_dlev_target_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_en != "radp_vga_en_enalbe")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_hold_en != "radp_vga_hold_en_not_hold")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_hold_en_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_initial_load != "radp_vga_initial_load_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_initial_load_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_initial_value != "radp_vga_initial_value_16")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_initial_value_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_onetime != "radp_vga_onetime_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_onetime_check ( .error(1'b1) );
		end
		if (pma_adapt_adp_vga_onetime_threshold != "radp_vga_onetime_threshold_512")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_adp_vga_onetime_threshold_check ( .error(1'b1) );
		end
		if (pma_adapt_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_adapt_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_initial_settings_check ( .error(1'b1) );
		end
		if (pma_adapt_odi_mode != "odi_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_odi_mode_check ( .error(1'b1) );
		end
		if (pma_adapt_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_optimal_check ( .error(1'b1) );
		end
		if (pma_adapt_power_mode != "powsav_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_power_mode_check ( .error(1'b1) );
		end
		if (pma_adapt_prot_mode != "basic_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_prot_mode_check ( .error(1'b1) );
		end
		if (pma_adapt_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_sup_mode_check ( .error(1'b1) );
		end
		if (pma_adapt_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_adapt_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_adapt_bti_en != "adapt_bti_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_adapt_bti_en_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_atb_select != "atb_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_atb_select_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_bti_protected != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_bti_protected_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_datarate_bps != "25781250000")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_datarate_bps_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_dfe_bti_en != "dfe_bti_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_dfe_bti_en_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_dfe_mode != "dfe_tap1_15")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_dfe_mode_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_dft_en != "dft_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_dft_en_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_dft_hilospeed_sel != "dft_osc_lospeed_path")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_dft_hilospeed_sel_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_dft_osc_sel != "dft_osc_even")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_dft_osc_sel_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_h1edge_bti_en != "h1edge_bti_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_h1edge_bti_en_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_initial_settings_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_latch_xcouple_disable != "latch_xcouple_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_latch_xcouple_disable_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdr0e != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdr0e_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdr0e_sgn != "oc_sa_cdr0e_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdr0e_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdr0o != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdr0o_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdr0o_sgn != "oc_sa_cdr0o_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdr0o_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdrne != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdrne_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdrne_sgn != "oc_sa_cdrne_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdrne_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdrno != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdrno_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdrno_sgn != "oc_sa_cdrno_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdrno_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdrpe != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdrpe_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdrpe_sgn != "oc_sa_cdrpe_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdrpe_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdrpo != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdrpo_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_cdrpo_sgn != "oc_sa_cdrpo_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_cdrpo_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_dne != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_dne_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_dne_sgn != "oc_sa_dne_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_dne_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_dno != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_dno_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_dno_sgn != "oc_sa_dno_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_dno_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_dpe != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_dpe_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_dpe_sgn != "oc_sa_dpe_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_dpe_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_dpo != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_dpo_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_dpo_sgn != "oc_sa_dpo_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_dpo_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_odie != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_odie_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_odie_sgn != "oc_sa_odie_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_odie_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_odio != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_odio_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_odio_sgn != "oc_sa_odio_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_odio_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_vrefe != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_vrefe_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_vrefe_sgn != "oc_sa_vrefe_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_vrefe_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_vrefo != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_vrefo_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_oc_sa_vrefo_sgn != "oc_sa_vrefo_sgn_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_oc_sa_vrefo_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_odi_bti_en != "odi_bti_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_odi_bti_en_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_odi_dlev_sign != "odi_dlev_pos")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_odi_dlev_sign_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_odi_h1_sign != "odi_h1_pos")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_odi_h1_sign_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_optimal_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_pdb != "dfe_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_pdb_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_pdb_edge_pre_h1 != "cdr_pre_h1_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_pdb_edge_pre_h1_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_pdb_edge_pst_h1 != "cdr_pst_h1_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_pdb_edge_pst_h1_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_pdb_tap_10t15 != "tap10t15_dfe_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_pdb_tap_10t15_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_pdb_tap_4t9 != "tap4t9_dfe_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_pdb_tap_4t9_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_pdb_tapsum != "tapsum_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_pdb_tapsum_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_power_mode != "high_perf")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_power_mode_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_prot_mode != "basic_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_prot_mode_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_sel_oc_en != "off_canc_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_sel_oc_en_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_sel_probe_tstmx != "probe_tstmx_none")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_sel_probe_tstmx_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_sup_mode_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap10_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap10_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap10_sgn != "tap10_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap10_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap11_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap11_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap11_sgn != "tap11_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap11_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap12_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap12_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap12_sgn != "tap12_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap12_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap13_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap13_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap13_sgn != "tap13_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap13_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap14_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap14_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap14_sgn != "tap14_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap14_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap15_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap15_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap15_sgn != "tap15_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap15_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap1_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap1_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap1_sgn != "tap1_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap1_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap2_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap2_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap2_sgn != "tap2_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap2_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap3_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap3_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap3_sgn != "tap3_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap3_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap4_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap4_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap4_sgn != "tap4_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap4_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap5_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap5_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap5_sgn != "tap5_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap5_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap6_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap6_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap6_sgn != "tap6_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap6_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap7_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap7_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap7_sgn != "tap7_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap7_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap8_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap8_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap8_sgn != "tap8_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap8_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap9_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap9_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tap9_sgn != "tap9_sign_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tap9_sgn_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_tapsum_bw_sel != "tapsum_hibw")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_tapsum_bw_sel_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_vref_coeff != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_vref_coeff_check ( .error(1'b1) );
		end
		if (pma_rx_dfe_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_dfe_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_rx_sd_link != "sr")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_link_check ( .error(1'b1) );
		end
		if (pma_rx_sd_optimal != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_optimal_check ( .error(1'b1) );
		end
		if (pma_rx_sd_power_mode != "high_perf")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_power_mode_check ( .error(1'b1) );
		end
		if (pma_rx_sd_prot_mode != "basic_rx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_prot_mode_check ( .error(1'b1) );
		end
		if (pma_rx_sd_sd_output_off != "clk_divrx_2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_sd_output_off_check ( .error(1'b1) );
		end
		if (pma_rx_sd_sd_output_on != "force_sd_output_on")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_sd_output_on_check ( .error(1'b1) );
		end
		if (pma_rx_sd_sd_pdb != "sd_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_sd_pdb_check ( .error(1'b1) );
		end
		if (pma_rx_sd_sd_threshold != "sdlv_3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_sd_threshold_check ( .error(1'b1) );
		end
		if (pma_rx_sd_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_sup_mode_check ( .error(1'b1) );
		end
		if (pma_rx_sd_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_rx_sd_silicon_rev_check ( .error(1'b1) );
		end
		if (pma_pcie_gen_switch_silicon_rev != "14nm5cr2")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					pma_pcie_gen_switch_silicon_rev_check ( .error(1'b1) );
		end
	endgenerate

	ex_100g_altera_xcvr_native_s10_htile_180_m3pnzmq #(
		.rcfg_enable                                                                     (1),
		.rcfg_jtag_enable                                                                (1),
		.rcfg_separate_avmm_busy                                                         (0),
		.dbg_embedded_debug_enable                                                       (1),
		.dbg_capability_reg_enable                                                       (1),
		.dbg_user_identifier                                                             (0),
		.dbg_stat_soft_logic_enable                                                      (1),
		.dbg_ctrl_soft_logic_enable                                                      (1),
		.rcfg_emb_strm_enable                                                            (0),
		.rcfg_profile_cnt                                                                (2),
		.device_revision                                                                 ("14nm5cr2"),
		.silicon_revision                                                                ("14nm5cr2"),
		.reduced_reset_sim_time                                                          (0),
		.duplex_mode                                                                     ("duplex"),
		.channels                                                                        (4),
		.enable_calibration                                                              (1),
		.enable_direct_reset_control                                                     (0),
		.disable_reset_sequencer                                                         (0),
		.disable_digital_reset_sequencer                                                 (0),
		.l_release_aib_reset_first                                                       (1),
		.bonded_mode                                                                     ("not_bonded"),
		.pcs_bonding_master                                                              (0),
		.pcs_reset_sequencing_mode                                                       ("bonded"),
		.enable_manual_bonding_settings                                                  (0),
		.manual_pcs_bonding_mode                                                         ("individual"),
		.manual_pcs_bonding_comp_cnt                                                     (0),
		.manual_tx_hssi_aib_bonding_mode                                                 ("individual"),
		.manual_tx_hssi_aib_bonding_comp_cnt                                             (0),
		.manual_tx_core_aib_bonding_mode                                                 ("individual"),
		.manual_tx_core_aib_bonding_comp_cnt                                             (0),
		.manual_rx_hssi_aib_bonding_mode                                                 ("individual"),
		.manual_rx_hssi_aib_bonding_comp_cnt                                             (0),
		.manual_rx_core_aib_bonding_mode                                                 ("individual"),
		.manual_rx_core_aib_bonding_comp_cnt                                             (0),
		.plls                                                                            (1),
		.number_physical_bonding_clocks                                                  (1),
		.cdr_refclk_cnt                                                                  (1),
		.enable_hip                                                                      (0),
		.hip_cal_en                                                                      ("disable"),
		.enable_ehip                                                                     (0),
		.enable_tx_fast_pipeln_reg                                                       (0),
		.enable_rx_fast_pipeln_reg                                                       (0),
		.tx_coreclkin_clock_network                                                      ("dedicated"),
		.tx_pcs_bonding_clock_network                                                    ("dedicated"),
		.rx_coreclkin_clock_network                                                      ("dedicated"),
		.osc_clk_divider                                                                 (1),
		.enable_tx_x2_coreclkin_port                                                     (0),
		.rcfg_shared                                                                     (1),
		.adme_prot_mode                                                                  ("basic_enh"),
		.adme_pma_mode                                                                   ("basic"),
		.adme_tx_power_mode                                                              ("high_perf"),
		.adme_data_rate                                                                  ("25781250000"),
		.dbg_prbs_soft_logic_enable                                                      (1),
		.dbg_odi_soft_logic_enable                                                       (0),
		.enable_rcfg_tx_digitalreset_release_ctrl                                        (0),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_advanced_user_mode_rx                       ("disable"),
		.hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode                       ("tx_rx_pair_enabled"),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_channel_operation_mode                      ("tx_rx_pair_enabled"),
		.hssi_rx_pld_pcs_interface_hd_pcs8g_channel_operation_mode                       ("tx_rx_pair_enabled"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_channel_operation_mode                 ("tx_rx_pair_enabled"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_channel_operation_mode          ("tx_rx_pair_enabled"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_channel_operation_mode  ("tx_rx_pair_enabled"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_clklow_clk_hz                          (322265625),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_ctrl_plane_bonding_rx                  ("individual_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_fifo_mode_rx                                ("reg_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs8g_fifo_mode_rx                                 ("reg_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_fref_clk_hz                            (322265625),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_frequency_rules_en                     ("enable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_func_mode                              ("enable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_hclk_clk_hz                            (0),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_hip_en                                 ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs8g_hip_mode                                     ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_hrdrstctl_en                           ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_hrdrstctl_en                    ("disable"),
		.hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx                            ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_low_latency_en_rx                           ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_low_latency_en_rx                      ("disable"),
		.hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en                                      ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_lpbk_en                                     ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs8g_lpbk_en                                      ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_lpbk_en                                ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_lpbk_en                         ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_operating_voltage                      ("standard"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_ac_pwr_rules_en                    ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_pair_ac_pwr_uw_per_mhz             (0),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_rx_ac_pwr_uw_per_mhz               (0),
		.hssi_rx_pld_pcs_interface_pcs_rx_block_sel                                      ("teng"),
		.hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel                                    ("teng_clk_out"),
		.hssi_rx_pld_pcs_interface_pcs_rx_clk_sel                                        ("pcs_rx_clk"),
		.hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en                                     ("hip_rx_disable"),
		.hssi_rx_pld_pcs_interface_pcs_rx_output_sel                                     ("teng_output"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pcs_rx_pwr_scaling_clk                 ("pma_rx_clk"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_8g_refclk_dig_nonatpg_mode_clk_hz  (0),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_fifo_mode_rx                       ("reg_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_pcs_refclk_dig_nonatpg_mode_clk_hz (0),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_rx_clk_hz                          (0),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_pma_dw_rx                                   ("pma_64b_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs8g_pma_dw_rx                                    ("pma_10b_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_dw_rx                              ("pma_64b_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_pma_dw_rx                       ("pma_64b_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_rx_clk_hz                          (402832031),
		.hssi_rx_pld_pcs_interface_hd_g3pcs_prot_mode                                    ("disabled_prot_mode"),
		.hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx                                 ("disabled_prot_mode_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_prot_mode_rx                                ("basic_mode_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs8g_prot_mode_rx                                 ("disabled_prot_mode_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_prot_mode_rx                           ("basic_10gpcs_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_prot_mode_rx                    ("teng_reg_mode_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_prot_mode_rx                    ("teng_basic_mode_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_prot_mode_rx            ("teng_mode_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_shared_fifo_width_rx                        ("single_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_shared_fifo_width_rx                   ("single_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_shared_fifo_width_rx    ("single_rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_sim_mode                        ("disable"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_speed_grade                            ("e2"),
		.hssi_rx_pld_pcs_interface_hd_g3pcs_sup_mode                                     ("user_mode"),
		.hssi_rx_pld_pcs_interface_hd_krfec_sup_mode                                     ("user_mode"),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_sup_mode                                    ("user_mode"),
		.hssi_rx_pld_pcs_interface_hd_pcs8g_sup_mode                                     ("user_mode"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_sup_mode                               ("user_mode"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pld_if_sup_mode                        ("user_mode"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_pma_if_sup_mode                        ("user_mode"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_sup_mode                ("user_mode"),
		.hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode                                ("tx"),
		.hssi_rx_pld_pcs_interface_hd_pcs10g_test_bus_mode                               ("rx"),
		.hssi_rx_pld_pcs_interface_hd_pcs_channel_transparent_pcs_rx                     ("disable"),
		.hssi_rx_pld_pcs_interface_silicon_rev                                           ("14nm5cr2"),
		.hssi_tx_pld_pcs_interface_hd_pcs10g_advanced_user_mode_tx                       ("disable"),
		.hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode                       ("tx_rx_pair_enabled"),
		.hssi_tx_pld_pcs_interface_hd_pcs10g_channel_operation_mode                      ("tx_rx_pair_enabled"),
		.hssi_tx_pld_pcs_interface_hd_pcs8g_channel_operation_mode                       ("tx_rx_pair_enabled"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_channel_operation_mode                 ("tx_rx_pair_enabled"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_channel_operation_mode          ("tx_rx_pair_enabled"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_channel_operation_mode  ("tx_rx_pair_enabled"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_ctrl_plane_bonding              ("individual"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_ctrl_plane_bonding_tx                  ("individual_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs10g_fifo_mode_tx                                ("reg_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs8g_fifo_mode_tx                                 ("reg_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_frequency_rules_en                     ("enable"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_func_mode                              ("enable"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_hclk_clk_hz                            (0),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_hip_en                                 ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs8g_hip_mode                                     ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_hrdrstctl_en                           ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_hrdrstctl_en                    ("disable"),
		.hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx                            ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs10g_low_latency_en_tx                           ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_low_latency_en_tx                      ("disable"),
		.hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en                                      ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs10g_lpbk_en                                     ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs8g_lpbk_en                                      ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_lpbk_en                                ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_lpbk_en                         ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pcs_tx_ac_pwr_uw_per_mhz               (0),
		.hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel                                    ("teng_clk_out"),
		.hssi_tx_pld_pcs_interface_pcs_tx_clk_source                                     ("teng"),
		.hssi_tx_pld_pcs_interface_pcs_tx_data_source                                    ("hip_disable"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en                                  ("delay1_clk_disable"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel                                 ("pcs_tx_clk"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl                                    ("delay1_path0"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel                                ("one_ff_delay"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en                                  ("delay2_clk_disable"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl                                    ("delay2_path0"),
		.hssi_tx_pld_pcs_interface_pcs_tx_output_sel                                     ("teng_output"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pcs_tx_pwr_scaling_clk                 ("pma_tx_clk"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_8g_refclk_dig_nonatpg_mode_clk_hz  (0),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_fifo_mode_tx                       ("reg_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_pcs_refclk_dig_nonatpg_mode_clk_hz (0),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_tx_clk_hz                          (0),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_uhsif_tx_clk_hz                    (0),
		.hssi_tx_pld_pcs_interface_hd_pcs10g_pma_dw_tx                                   ("pma_64b_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs8g_pma_dw_tx                                    ("pma_10b_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_dw_tx                              ("pma_64b_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_pma_dw_tx                       ("pma_64b_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_tx_clk_hz                          (402832031),
		.hssi_tx_pld_pcs_interface_hd_g3pcs_prot_mode                                    ("disabled_prot_mode"),
		.hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx                                 ("disabled_prot_mode_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs10g_prot_mode_tx                                ("basic_mode_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs8g_prot_mode_tx                                 ("disabled_prot_mode_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_prot_mode_tx                           ("basic_10gpcs_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_prot_mode_tx                    ("teng_reg_mode_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_prot_mode_tx                    ("teng_basic_mode_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_prot_mode_tx            ("teng_mode_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs10g_shared_fifo_width_tx                        ("single_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_shared_fifo_width_tx                   ("single_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_shared_fifo_width_tx    ("single_tx"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_sim_mode                        ("disable"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_speed_grade                            ("e2"),
		.hssi_tx_pld_pcs_interface_hd_g3pcs_sup_mode                                     ("user_mode"),
		.hssi_tx_pld_pcs_interface_hd_krfec_sup_mode                                     ("user_mode"),
		.hssi_tx_pld_pcs_interface_hd_pcs10g_sup_mode                                    ("user_mode"),
		.hssi_tx_pld_pcs_interface_hd_pcs8g_sup_mode                                     ("user_mode"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_sup_mode                               ("user_mode"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pld_if_sup_mode                        ("user_mode"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_pma_if_sup_mode                        ("user_mode"),
		.hssi_tx_pld_pcs_interface_hd_pcs_channel_share_fifo_mem_sup_mode                ("user_mode"),
		.hssi_tx_pld_pcs_interface_silicon_rev                                           ("14nm5cr2"),
		.hssi_10g_tx_pcs_advanced_user_mode                                              ("disable"),
		.hssi_10g_tx_pcs_bitslip_en                                                      ("bitslip_dis"),
		.hssi_10g_tx_pcs_bonding_dft_en                                                  ("dft_dis"),
		.hssi_10g_tx_pcs_bonding_dft_val                                                 ("dft_0"),
		.hssi_10g_tx_pcs_crcgen_bypass                                                   ("crcgen_bypass_en"),
		.hssi_10g_tx_pcs_crcgen_clken                                                    ("crcgen_clk_dis"),
		.hssi_10g_tx_pcs_crcgen_err                                                      ("crcgen_err_dis"),
		.hssi_10g_tx_pcs_crcgen_inv                                                      ("crcgen_inv_en"),
		.hssi_10g_tx_pcs_ctrl_bit_reverse                                                ("ctrl_bit_reverse_dis"),
		.hssi_10g_tx_pcs_data_bit_reverse                                                ("data_bit_reverse_dis"),
		.hssi_10g_tx_pcs_dft_clk_out_sel                                                 ("tx_master_clk"),
		.hssi_10g_tx_pcs_dispgen_bypass                                                  ("dispgen_bypass_en"),
		.hssi_10g_tx_pcs_dispgen_clken                                                   ("dispgen_clk_dis"),
		.hssi_10g_tx_pcs_dispgen_err                                                     ("dispgen_err_dis"),
		.hssi_10g_tx_pcs_dispgen_pipeln                                                  ("dispgen_pipeln_dis"),
		.hssi_10g_tx_pcs_distdwn_bypass_pipeln                                           ("distdwn_bypass_pipeln_dis"),
		.hssi_10g_tx_pcs_distup_bypass_pipeln                                            ("distup_bypass_pipeln_dis"),
		.hssi_10g_tx_pcs_dv_bond                                                         ("dv_bond_dis"),
		.hssi_10g_tx_pcs_empty_flag_type                                                 ("empty_rd_side"),
		.hssi_10g_tx_pcs_enc64b66b_txsm_clken                                            ("enc64b66b_txsm_clk_dis"),
		.hssi_10g_tx_pcs_enc_64b66b_txsm_bypass                                          ("enc_64b66b_txsm_bypass_en"),
		.hssi_10g_tx_pcs_fastpath                                                        ("fastpath_en"),
		.hssi_10g_tx_pcs_fec_clken                                                       ("fec_clk_dis"),
		.hssi_10g_tx_pcs_fec_enable                                                      ("fec_dis"),
		.hssi_10g_tx_pcs_fifo_double_write                                               ("fifo_double_write_dis"),
		.hssi_10g_tx_pcs_fifo_reg_fast                                                   ("fifo_reg_fast_dis"),
		.hssi_10g_tx_pcs_fifo_stop_rd                                                    ("n_rd_empty"),
		.hssi_10g_tx_pcs_fifo_stop_wr                                                    ("n_wr_full"),
		.hssi_10g_tx_pcs_frmgen_burst                                                    ("frmgen_burst_dis"),
		.hssi_10g_tx_pcs_frmgen_bypass                                                   ("frmgen_bypass_en"),
		.hssi_10g_tx_pcs_frmgen_clken                                                    ("frmgen_clk_dis"),
		.hssi_10g_tx_pcs_frmgen_mfrm_length                                              (2048),
		.hssi_10g_tx_pcs_frmgen_pipeln                                                   ("frmgen_pipeln_en"),
		.hssi_10g_tx_pcs_frmgen_pyld_ins                                                 ("frmgen_pyld_ins_dis"),
		.hssi_10g_tx_pcs_frmgen_wordslip                                                 ("frmgen_wordslip_dis"),
		.hssi_10g_tx_pcs_full_flag_type                                                  ("full_wr_side"),
		.hssi_10g_tx_pcs_gb_pipeln_bypass                                                ("disable"),
		.hssi_10g_tx_pcs_gb_tx_idwidth                                                   ("idwidth_66"),
		.hssi_10g_tx_pcs_gb_tx_odwidth                                                   ("odwidth_64"),
		.hssi_10g_tx_pcs_gbred_clken                                                     ("gbred_clk_en"),
		.hssi_10g_tx_pcs_indv                                                            ("indv_en"),
		.hssi_10g_tx_pcs_low_latency_en                                                  ("disable"),
		.hssi_10g_tx_pcs_master_clk_sel                                                  ("master_tx_pma_clk"),
		.hssi_10g_tx_pcs_pempty_flag_type                                                ("pempty_rd_side"),
		.hssi_10g_tx_pcs_pfull_flag_type                                                 ("pfull_wr_side"),
		.hssi_10g_tx_pcs_phcomp_rd_del                                                   ("phcomp_rd_del2"),
		.hssi_10g_tx_pcs_pld_if_type                                                     ("reg"),
		.hssi_10g_tx_pcs_prot_mode                                                       ("basic_mode"),
		.hssi_10g_tx_pcs_pseudo_random                                                   ("all_0"),
		.hssi_10g_tx_pcs_pseudo_seed_a                                                   ("288230376151711743"),
		.hssi_10g_tx_pcs_pseudo_seed_b                                                   ("288230376151711743"),
		.hssi_10g_tx_pcs_random_disp                                                     ("disable"),
		.hssi_10g_tx_pcs_rdfifo_clken                                                    ("rdfifo_clk_en"),
		.hssi_10g_tx_pcs_scrm_bypass                                                     ("scrm_bypass_en"),
		.hssi_10g_tx_pcs_scrm_clken                                                      ("scrm_clk_dis"),
		.hssi_10g_tx_pcs_scrm_mode                                                       ("async"),
		.hssi_10g_tx_pcs_scrm_pipeln                                                     ("enable"),
		.hssi_10g_tx_pcs_sh_err                                                          ("sh_err_dis"),
		.hssi_10g_tx_pcs_sop_mark                                                        ("sop_mark_dis"),
		.hssi_10g_tx_pcs_stretch_num_stages                                              ("one_stage"),
		.hssi_10g_tx_pcs_sup_mode                                                        ("user_mode"),
		.hssi_10g_tx_pcs_test_mode                                                       ("test_off"),
		.hssi_10g_tx_pcs_tx_scrm_err                                                     ("scrm_err_dis"),
		.hssi_10g_tx_pcs_tx_scrm_width                                                   ("bit64"),
		.hssi_10g_tx_pcs_tx_sh_location                                                  ("msb"),
		.hssi_10g_tx_pcs_tx_sm_bypass                                                    ("tx_sm_bypass_en"),
		.hssi_10g_tx_pcs_tx_sm_pipeln                                                    ("tx_sm_pipeln_en"),
		.hssi_10g_tx_pcs_tx_testbus_sel                                                  ("tx_fifo_testbus1"),
		.hssi_10g_tx_pcs_txfifo_empty                                                    ("empty_default"),
		.hssi_10g_tx_pcs_txfifo_full                                                     ("full_default"),
		.hssi_10g_tx_pcs_txfifo_mode                                                     ("register_mode"),
		.hssi_10g_tx_pcs_txfifo_pempty                                                   (2),
		.hssi_10g_tx_pcs_txfifo_pfull                                                    (11),
		.hssi_10g_tx_pcs_wr_clk_sel                                                      ("wr_tx_pma_clk"),
		.hssi_10g_tx_pcs_wrfifo_clken                                                    ("wrfifo_clk_en"),
		.hssi_10g_tx_pcs_silicon_rev                                                     ("14nm5cr2"),
		.hssi_8g_rx_pcs_auto_error_replacement                                           ("dis_err_replace"),
		.hssi_8g_rx_pcs_bit_reversal                                                     ("dis_bit_reversal"),
		.hssi_8g_rx_pcs_bonding_dft_en                                                   ("dft_dis"),
		.hssi_8g_rx_pcs_bonding_dft_val                                                  ("dft_0"),
		.hssi_8g_rx_pcs_bypass_pipeline_reg                                              ("dis_bypass_pipeline"),
		.hssi_8g_rx_pcs_byte_deserializer                                                ("dis_bds"),
		.hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask                                            ("dis_rxvalid_mask"),
		.hssi_8g_rx_pcs_clkcmp_pattern_n                                                 (0),
		.hssi_8g_rx_pcs_clkcmp_pattern_p                                                 (0),
		.hssi_8g_rx_pcs_clock_gate_bds_dec_asn                                           ("en_bds_dec_asn_clk_gating"),
		.hssi_8g_rx_pcs_clock_gate_cdr_eidle                                             ("en_cdr_eidle_clk_gating"),
		.hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk                                           ("en_dw_pc_wrclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_dw_rm_rd                                              ("en_dw_rm_rdclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_dw_rm_wr                                              ("en_dw_rm_wrclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_dw_wa                                                 ("en_dw_wa_clk_gating"),
		.hssi_8g_rx_pcs_clock_gate_pc_rdclk                                              ("en_pc_rdclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk                                           ("en_sw_pc_wrclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_sw_rm_rd                                              ("en_sw_rm_rdclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_sw_rm_wr                                              ("en_sw_rm_wrclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_sw_wa                                                 ("en_sw_wa_clk_gating"),
		.hssi_8g_rx_pcs_clock_observation_in_pld_core                                    ("internal_sw_wa_clk"),
		.hssi_8g_rx_pcs_eidle_entry_eios                                                 ("dis_eidle_eios"),
		.hssi_8g_rx_pcs_eidle_entry_iei                                                  ("dis_eidle_iei"),
		.hssi_8g_rx_pcs_eidle_entry_sd                                                   ("dis_eidle_sd"),
		.hssi_8g_rx_pcs_eightb_tenb_decoder                                              ("en_8b10b_ibm"),
		.hssi_8g_rx_pcs_err_flags_sel                                                    ("err_flags_wa"),
		.hssi_8g_rx_pcs_fixed_pat_det                                                    ("dis_fixed_patdet"),
		.hssi_8g_rx_pcs_fixed_pat_num                                                    (0),
		.hssi_8g_rx_pcs_force_signal_detect                                              ("en_force_signal_detect"),
		.hssi_8g_rx_pcs_gen3_clk_en                                                      ("disable_clk"),
		.hssi_8g_rx_pcs_gen3_rx_clk_sel                                                  ("rcvd_clk"),
		.hssi_8g_rx_pcs_gen3_tx_clk_sel                                                  ("tx_pma_clk"),
		.hssi_8g_rx_pcs_hip_mode                                                         ("dis_hip"),
		.hssi_8g_rx_pcs_ibm_invalid_code                                                 ("dis_ibm_invalid_code"),
		.hssi_8g_rx_pcs_invalid_code_flag_only                                           ("dis_invalid_code_only"),
		.hssi_8g_rx_pcs_pad_or_edb_error_replace                                         ("replace_edb"),
		.hssi_8g_rx_pcs_pcs_bypass                                                       ("dis_pcs_bypass"),
		.hssi_8g_rx_pcs_phase_comp_rdptr                                                 ("disable_rdptr"),
		.hssi_8g_rx_pcs_phase_compensation_fifo                                          ("register_fifo"),
		.hssi_8g_rx_pcs_pipe_if_enable                                                   ("dis_pipe_rx"),
		.hssi_8g_rx_pcs_pma_dw                                                           ("ten_bit"),
		.hssi_8g_rx_pcs_polinv_8b10b_dec                                                 ("dis_polinv_8b10b_dec"),
		.hssi_8g_rx_pcs_prot_mode                                                        ("disabled_prot_mode"),
		.hssi_8g_rx_pcs_rate_match                                                       ("dis_rm"),
		.hssi_8g_rx_pcs_rate_match_del_thres                                             ("dis_rm_del_thres"),
		.hssi_8g_rx_pcs_rate_match_empty_thres                                           ("dis_rm_empty_thres"),
		.hssi_8g_rx_pcs_rate_match_full_thres                                            ("dis_rm_full_thres"),
		.hssi_8g_rx_pcs_rate_match_ins_thres                                             ("dis_rm_ins_thres"),
		.hssi_8g_rx_pcs_rate_match_start_thres                                           ("dis_rm_start_thres"),
		.hssi_8g_rx_pcs_rx_clk2                                                          ("rcvd_clk_clk2"),
		.hssi_8g_rx_pcs_rx_clk_free_running                                              ("en_rx_clk_free_run"),
		.hssi_8g_rx_pcs_rx_pcs_urst                                                      ("en_rx_pcs_urst"),
		.hssi_8g_rx_pcs_rx_rcvd_clk                                                      ("rcvd_clk_rcvd_clk"),
		.hssi_8g_rx_pcs_rx_rd_clk                                                        ("rx_clk"),
		.hssi_8g_rx_pcs_rx_refclk                                                        ("dis_refclk_sel"),
		.hssi_8g_rx_pcs_rx_wr_clk                                                        ("rx_clk2_div_1_2_4"),
		.hssi_8g_rx_pcs_sup_mode                                                         ("user_mode"),
		.hssi_8g_rx_pcs_symbol_swap                                                      ("dis_symbol_swap"),
		.hssi_8g_rx_pcs_sync_sm_idle_eios                                                ("dis_syncsm_idle"),
		.hssi_8g_rx_pcs_test_bus_sel                                                     ("tx_testbus"),
		.hssi_8g_rx_pcs_tx_rx_parallel_loopback                                          ("dis_plpbk"),
		.hssi_8g_rx_pcs_wa_boundary_lock_ctrl                                            ("sync_sm"),
		.hssi_8g_rx_pcs_wa_clk_slip_spacing                                              (16),
		.hssi_8g_rx_pcs_wa_det_latency_sync_status_beh                                   ("dont_care_assert_sync"),
		.hssi_8g_rx_pcs_wa_disp_err_flag                                                 ("en_disp_err_flag"),
		.hssi_8g_rx_pcs_wa_kchar                                                         ("dis_kchar"),
		.hssi_8g_rx_pcs_wa_pd                                                            ("wa_pd_10"),
		.hssi_8g_rx_pcs_wa_pd_data                                                       ("0"),
		.hssi_8g_rx_pcs_wa_pd_polarity                                                   ("dont_care_both_pol"),
		.hssi_8g_rx_pcs_wa_pld_controlled                                                ("dis_pld_ctrl"),
		.hssi_8g_rx_pcs_wa_renumber_data                                                 (3),
		.hssi_8g_rx_pcs_wa_rgnumber_data                                                 (3),
		.hssi_8g_rx_pcs_wa_rknumber_data                                                 (3),
		.hssi_8g_rx_pcs_wa_rosnumber_data                                                (1),
		.hssi_8g_rx_pcs_wa_rvnumber_data                                                 (0),
		.hssi_8g_rx_pcs_wa_sync_sm_ctrl                                                  ("gige_sync_sm"),
		.hssi_8g_rx_pcs_wait_cnt                                                         (0),
		.hssi_8g_rx_pcs_silicon_rev                                                      ("14nm5cr2"),
		.hssi_8g_tx_pcs_bit_reversal                                                     ("dis_bit_reversal"),
		.hssi_8g_tx_pcs_bonding_dft_en                                                   ("dft_dis"),
		.hssi_8g_tx_pcs_bonding_dft_val                                                  ("dft_0"),
		.hssi_8g_tx_pcs_bypass_pipeline_reg                                              ("dis_bypass_pipeline"),
		.hssi_8g_tx_pcs_byte_serializer                                                  ("dis_bs"),
		.hssi_8g_tx_pcs_clock_gate_bs_enc                                                ("en_bs_enc_clk_gating"),
		.hssi_8g_tx_pcs_clock_gate_dw_fifowr                                             ("en_dw_fifowr_clk_gating"),
		.hssi_8g_tx_pcs_clock_gate_fiford                                                ("en_fiford_clk_gating"),
		.hssi_8g_tx_pcs_clock_gate_sw_fifowr                                             ("en_sw_fifowr_clk_gating"),
		.hssi_8g_tx_pcs_clock_observation_in_pld_core                                    ("internal_refclk_b"),
		.hssi_8g_tx_pcs_data_selection_8b10b_encoder_input                               ("normal_data_path"),
		.hssi_8g_tx_pcs_dynamic_clk_switch                                               ("dis_dyn_clk_switch"),
		.hssi_8g_tx_pcs_eightb_tenb_disp_ctrl                                            ("dis_disp_ctrl"),
		.hssi_8g_tx_pcs_eightb_tenb_encoder                                              ("en_8b10b_ibm"),
		.hssi_8g_tx_pcs_force_echar                                                      ("dis_force_echar"),
		.hssi_8g_tx_pcs_force_kchar                                                      ("dis_force_kchar"),
		.hssi_8g_tx_pcs_gen3_tx_clk_sel                                                  ("dis_tx_clk"),
		.hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel                                             ("dis_tx_pipe_clk"),
		.hssi_8g_tx_pcs_hip_mode                                                         ("dis_hip"),
		.hssi_8g_tx_pcs_pcs_bypass                                                       ("dis_pcs_bypass"),
		.hssi_8g_tx_pcs_phase_comp_rdptr                                                 ("disable_rdptr"),
		.hssi_8g_tx_pcs_phase_compensation_fifo                                          ("register_fifo"),
		.hssi_8g_tx_pcs_phfifo_write_clk_sel                                             ("tx_clk"),
		.hssi_8g_tx_pcs_pma_dw                                                           ("ten_bit"),
		.hssi_8g_tx_pcs_prot_mode                                                        ("disabled_prot_mode"),
		.hssi_8g_tx_pcs_refclk_b_clk_sel                                                 ("tx_pma_clock"),
		.hssi_8g_tx_pcs_revloop_back_rm                                                  ("dis_rev_loopback_rx_rm"),
		.hssi_8g_tx_pcs_sup_mode                                                         ("user_mode"),
		.hssi_8g_tx_pcs_symbol_swap                                                      ("dis_symbol_swap"),
		.hssi_8g_tx_pcs_tx_bitslip                                                       ("dis_tx_bitslip"),
		.hssi_8g_tx_pcs_tx_compliance_controlled_disparity                               ("dis_txcompliance"),
		.hssi_8g_tx_pcs_tx_fast_pld_reg                                                  ("dis_tx_fast_pld_reg"),
		.hssi_8g_tx_pcs_txclk_freerun                                                    ("en_freerun_tx"),
		.hssi_8g_tx_pcs_txpcs_urst                                                       ("en_txpcs_urst"),
		.hssi_8g_tx_pcs_silicon_rev                                                      ("14nm5cr2"),
		.hssi_avmm1_if_pcs_arbiter_ctrl                                                  ("avmm1_arbiter_uc_sel"),
		.hssi_avmm1_if_pcs_cal_done                                                      ("avmm1_cal_done_deassert"),
		.hssi_avmm1_if_pcs_cal_reserved                                                  (0),
		.hssi_avmm1_if_pcs_calibration_feature_en                                        ("avmm1_pcs_calibration_en"),
		.hssi_avmm1_if_pldadapt_gate_dis                                                 ("disable"),
		.hssi_avmm1_if_pcs_hip_cal_en                                                    ("disable"),
		.hssi_avmm1_if_hssiadapt_nfhssi_calibratio_feature_en                            ("disable"),
		.hssi_avmm1_if_pldadapt_nfhssi_calibratio_feature_en                             ("enable"),
		.hssi_avmm1_if_hssiadapt_read_blocking_enable                                    ("enable"),
		.hssi_avmm1_if_pldadapt_read_blocking_enable                                     ("enable"),
		.hssi_avmm1_if_hssiadapt_uc_blocking_enable                                      ("enable"),
		.hssi_avmm1_if_pldadapt_uc_blocking_enable                                       ("enable"),
		.hssi_avmm1_if_hssiadapt_avmm_osc_clock_setting                                  ("osc_clk_div_by1"),
		.hssi_avmm1_if_pldadapt_avmm_osc_clock_setting                                   ("osc_clk_div_by1"),
		.hssi_avmm1_if_hssiadapt_avmm_testbus_sel                                        ("avmm1_transfer_testbus"),
		.hssi_avmm1_if_pldadapt_avmm_testbus_sel                                         ("avmm1_transfer_testbus"),
		.hssi_avmm1_if_hssiadapt_hip_mode                                                ("disable_hip"),
		.hssi_avmm1_if_pldadapt_hip_mode                                                 ("disable_hip"),
		.hssi_avmm1_if_silicon_rev                                                       ("14nm5cr2"),
		.hssi_avmm1_if_calibration_type                                                  ("one_time"),
		.pma_cgb_bitslip_enable                                                          ("disable_bitslip"),
		.pma_cgb_bti_protected                                                           ("false"),
		.pma_cgb_cgb_bti_en                                                              ("cgb_bti_disable"),
		.pma_cgb_cgb_power_down                                                          ("normal_cgb"),
		.pma_cgb_datarate_bps                                                            ("25781250000"),
		.pma_cgb_initial_settings                                                        ("true"),
		.pma_cgb_observe_cgb_clocks                                                      ("observe_nothing"),
		.pma_cgb_pcie_gen                                                                ("non_pcie"),
		.pma_cgb_pcie_gen3_bitwidth                                                      ("pciegen3_wide"),
		.pma_cgb_power_rail_er                                                           (1120),
		.pma_cgb_prot_mode                                                               ("basic_tx"),
		.pma_cgb_ser_mode                                                                ("sixty_four_bit"),
		.pma_cgb_ser_powerdown                                                           ("normal_poweron_ser"),
		.pma_cgb_sup_mode                                                                ("user_mode"),
		.pma_cgb_tx_ucontrol_en                                                          ("disable"),
		.pma_cgb_tx_ucontrol_pcie                                                        ("gen1"),
		.pma_cgb_tx_ucontrol_reset                                                       ("disable"),
		.pma_cgb_uc_cgb_vreg_boost                                                       ("no_voltage_boost"),
		.pma_cgb_uc_vcc_setting                                                          ("vcc_setting2"),
		.pma_cgb_vccdreg_output                                                          ("vccdreg_nominal"),
		.pma_cgb_vreg_sel_ref                                                            ("sel_vccer_4ref"),
		.pma_cgb_x1_div_m_sel                                                            ("divbypass"),
		.pma_cgb_silicon_rev                                                             ("14nm5cr2"),
		.pma_cgb_input_select_x1                                                         ("fpll_bot"),
		.pma_cgb_input_select_gen3                                                       ("not_used"),
		.pma_cgb_input_select_xn                                                         ("not_used"),
		.pma_tx_buf_pm_cr2_tx_path_analog_mode                                           ("user_custom"),
		.pma_tx_buf_bti_protected                                                        ("false"),
		.pma_tx_buf_calibration_en                                                       ("false"),
		.pma_tx_buf_pm_cr2_tx_path_calibration_en                                        ("false"),
		.pma_tx_buf_calibration_resistor_value                                           ("res_setting0"),
		.pma_tx_buf_cdr_cp_calibration_en                                                ("cdr_cp_cal_disable"),
		.pma_tx_buf_chgpmp_current_dn_trim                                               ("cp_current_trimming_dn_setting0"),
		.pma_tx_buf_chgpmp_current_up_trim                                               ("cp_current_trimming_up_setting0"),
		.pma_tx_buf_chgpmp_dn_trim_double                                                ("normal_dn_trim_current"),
		.pma_tx_buf_chgpmp_up_trim_double                                                ("normal_up_trim_current"),
		.pma_tx_buf_pm_cr2_tx_path_clock_divider_ratio                                   (1),
		.pma_tx_buf_compensation_en                                                      ("enable"),
		.pma_tx_buf_compensation_posttap_en                                              ("disable"),
		.pma_tx_buf_cpen_ctrl                                                            ("cp_l1"),
		.pma_tx_buf_datarate_bps                                                         ("25781250000"),
		.pma_tx_buf_pm_cr2_tx_path_datarate_bps                                          ("25781250000"),
		.pma_tx_buf_pm_cr2_tx_path_datawidth                                             (64),
		.pma_tx_buf_dcc_finestep_enin                                                    ("enable"),
		.pma_tx_buf_dcd_clk_div_ctrl                                                     ("dcd_ck_div128"),
		.pma_tx_buf_dcd_detection_en                                                     ("disable"),
		.pma_tx_buf_dft_sel                                                              ("dft_disabled"),
		.pma_tx_buf_duty_cycle_correction_bandwidth                                      ("dcc_bw_2"),
		.pma_tx_buf_duty_cycle_correction_bandwidth_dn                                   ("dcd_bw_dn_2"),
		.pma_tx_buf_duty_cycle_correction_reference1                                     ("dcc_ref1_4"),
		.pma_tx_buf_duty_cycle_correction_reference2                                     ("dcc_ref2_2"),
		.pma_tx_buf_duty_cycle_correction_reset_n                                        ("reset"),
		.pma_tx_buf_duty_cycle_cp_comp_en                                                ("cp_comp_off"),
		.pma_tx_buf_duty_cycle_detector_cp_cal                                           ("dcd_cp_cal_disable"),
		.pma_tx_buf_duty_cycle_detector_sa_cal                                           ("dcd_sa_cal_disable"),
		.pma_tx_buf_duty_cycle_input_polarity                                            ("dcc_input_pos"),
		.pma_tx_buf_duty_cycle_setting                                                   ("dcc_t32"),
		.pma_tx_buf_duty_cycle_setting_aux                                               ("dcc2_t32"),
		.pma_tx_buf_pm_cr2_tx_path_gt_enabled                                            ("enable"),
		.pma_tx_buf_idle_ctrl                                                            ("id_cpen_off"),
		.pma_tx_buf_initial_settings                                                     ("true"),
		.pma_tx_buf_pm_cr2_tx_path_initial_settings                                      ("true"),
		.pma_tx_buf_jtag_drv_sel                                                         ("drv1"),
		.pma_tx_buf_jtag_lp                                                              ("lp_off"),
		.pma_tx_buf_pm_cr2_tx_path_link                                                  ("sr"),
		.pma_tx_buf_low_power_en                                                         ("disable"),
		.pma_tx_buf_lst                                                                  ("atb_disabled"),
		.pma_tx_buf_pm_cr2_tx_rx_mcgb_location_for_pcie                                  (0),
		.pma_tx_buf_optimal                                                              ("true"),
		.pma_tx_buf_pm_cr2_tx_path_optimal                                               ("true"),
		.pma_tx_buf_pcie_gen                                                             ("non_pcie"),
		.pma_tx_buf_pm_cr2_tx_path_pma_tx_divclk_hz                                      ("402832031"),
		.pma_tx_buf_pm_cr2_tx_path_power_mode                                            ("high_perf"),
		.pma_tx_buf_pm_cr2_tx_path_power_rail_eht                                        (1800),
		.pma_tx_buf_power_rail_er                                                        (0),
		.pma_tx_buf_pm_cr2_tx_path_power_rail_et                                         (1120),
		.pma_tx_buf_powermode_ac_post_tap                                                ("tx_post_tap_ac_off"),
		.pma_tx_buf_powermode_ac_pre_tap                                                 ("tx_pre_tap_ac_off"),
		.pma_tx_buf_powermode_ac_tx_vod_no_jitcomp                                       ("tx_vod_no_jitcomp_ac_l0"),
		.pma_tx_buf_powermode_ac_tx_vod_w_jitcomp                                        ("tx_vod_w_jitcomp_ac_l31"),
		.pma_tx_buf_powermode_dc_post_tap                                                ("powerdown_tx_post_tap"),
		.pma_tx_buf_powermode_dc_pre_tap                                                 ("powerdown_tx_pre_tap"),
		.pma_tx_buf_powermode_dc_tx_vod_no_jitcomp                                       ("powerdown_tx_vod_no_jitcomp"),
		.pma_tx_buf_powermode_dc_tx_vod_w_jitcomp                                        ("tx_vod_w_jitcomp_dc_l31"),
		.pma_tx_buf_pre_emp_sign_1st_post_tap                                            ("fir_post_1t_neg"),
		.pma_tx_buf_pre_emp_sign_pre_tap_1t                                              ("fir_pre_1t_neg"),
		.pma_tx_buf_pre_emp_switching_ctrl_1st_post_tap                                  (0),
		.pma_tx_buf_pre_emp_switching_ctrl_pre_tap_1t                                    (0),
		.pma_tx_buf_prot_mode                                                            ("basic_tx"),
		.pma_tx_buf_pm_cr2_tx_path_prot_mode                                             ("basic_tx"),
		.pma_tx_buf_res_cal_local                                                        ("non_local"),
		.pma_tx_buf_rx_det                                                               ("mode_0"),
		.pma_tx_buf_rx_det_output_sel                                                    ("rx_det_pcie_out"),
		.pma_tx_buf_rx_det_pdb                                                           ("rx_det_off"),
		.pma_tx_buf_sense_amp_offset_cal_curr_n                                          ("sa_os_cal_in_0"),
		.pma_tx_buf_sense_amp_offset_cal_curr_p                                          (0),
		.pma_tx_buf_ser_powerdown                                                        ("normal_ser_on"),
		.pma_tx_buf_slew_rate_ctrl                                                       ("slew_r5"),
		.pma_tx_buf_pm_cr2_tx_path_speed_grade                                           ("e2"),
		.pma_tx_buf_sup_mode                                                             ("user_mode"),
		.pma_tx_buf_pm_cr2_tx_path_sup_mode                                              ("user_mode"),
		.pma_tx_buf_swing_level                                                          ("hv"),
		.pma_tx_buf_pm_cr2_tx_path_swing_level                                           ("hv"),
		.pma_tx_buf_term_code                                                            ("rterm_code7"),
		.pma_tx_buf_term_n_tune                                                          ("rterm_n7"),
		.pma_tx_buf_term_p_tune                                                          ("rterm_p7"),
		.pma_tx_buf_term_sel                                                             ("r_r2"),
		.pma_tx_buf_pm_cr2_tx_path_tile_type                                             ("h"),
		.pma_tx_buf_tri_driver                                                           ("tri_driver_disable"),
		.pma_tx_buf_pm_cr2_tx_path_tx_pll_clk_hz                                         ("12890625000"),
		.pma_tx_buf_tx_powerdown                                                         ("normal_tx_on"),
		.pma_tx_buf_tx_rst_enable                                                        ("enable"),
		.pma_tx_buf_xtx_path_xcgb_tx_ucontrol_en                                         ("disable"),
		.pma_tx_buf_uc_gen3                                                              ("gen3_off"),
		.pma_tx_buf_uc_gen4                                                              ("gen4_off"),
		.pma_tx_buf_uc_tx_cal                                                            ("uc_tx_cal_on"),
		.pma_tx_buf_uc_vcc_setting                                                       ("vcc_setting2"),
		.pma_tx_buf_user_fir_coeff_ctrl_sel                                              ("ram_ctl"),
		.pma_tx_buf_vod_output_swing_ctrl                                                (31),
		.pma_tx_buf_vreg_output                                                          ("vccdreg_nominal"),
		.pma_tx_buf_silicon_rev                                                          ("14nm5cr2"),
		.pma_tx_sequencer_tx_path_rstn_overrideb                                         ("use_sequencer"),
		.pma_tx_sequencer_xtx_path_xcgb_tx_ucontrol_en                                   ("disable"),
		.pma_tx_sequencer_xrx_path_uc_cal_clk_bypass                                     ("cal_clk_0"),
		.pma_tx_sequencer_silicon_rev                                                    ("14nm5cr2"),
		.hssi_10g_rx_pcs_advanced_user_mode                                              ("disable"),
		.hssi_10g_rx_pcs_align_del                                                       ("align_del_dis"),
		.hssi_10g_rx_pcs_ber_bit_err_total_cnt                                           ("bit_err_total_cnt_10g"),
		.hssi_10g_rx_pcs_ber_clken                                                       ("ber_clk_dis"),
		.hssi_10g_rx_pcs_ber_xus_timer_window                                            (19530),
		.hssi_10g_rx_pcs_bitslip_mode                                                    ("bitslip_en"),
		.hssi_10g_rx_pcs_blksync_bitslip_type                                            ("bitslip_comb"),
		.hssi_10g_rx_pcs_blksync_bitslip_wait_cnt                                        (1),
		.hssi_10g_rx_pcs_blksync_bitslip_wait_type                                       ("bitslip_cnt"),
		.hssi_10g_rx_pcs_blksync_bypass                                                  ("blksync_bypass_en"),
		.hssi_10g_rx_pcs_blksync_clken                                                   ("blksync_clk_en"),
		.hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt                                     ("enum_invalid_sh_cnt_10g"),
		.hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock                                    ("knum_sh_cnt_postlock_10g"),
		.hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock                                     ("knum_sh_cnt_prelock_10g"),
		.hssi_10g_rx_pcs_blksync_pipeln                                                  ("blksync_pipeln_dis"),
		.hssi_10g_rx_pcs_clr_errblk_cnt_en                                               ("disable"),
		.hssi_10g_rx_pcs_control_del                                                     ("control_del_none"),
		.hssi_10g_rx_pcs_crcchk_bypass                                                   ("crcchk_bypass_en"),
		.hssi_10g_rx_pcs_crcchk_clken                                                    ("crcchk_clk_dis"),
		.hssi_10g_rx_pcs_crcchk_inv                                                      ("crcchk_inv_en"),
		.hssi_10g_rx_pcs_crcchk_pipeln                                                   ("crcchk_pipeln_en"),
		.hssi_10g_rx_pcs_crcflag_pipeln                                                  ("crcflag_pipeln_en"),
		.hssi_10g_rx_pcs_ctrl_bit_reverse                                                ("ctrl_bit_reverse_dis"),
		.hssi_10g_rx_pcs_data_bit_reverse                                                ("data_bit_reverse_dis"),
		.hssi_10g_rx_pcs_dec64b66b_clken                                                 ("dec64b66b_clk_dis"),
		.hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass                                          ("dec_64b66b_rxsm_bypass_en"),
		.hssi_10g_rx_pcs_descrm_bypass                                                   ("descrm_bypass_en"),
		.hssi_10g_rx_pcs_descrm_clken                                                    ("descrm_clk_dis"),
		.hssi_10g_rx_pcs_descrm_mode                                                     ("async"),
		.hssi_10g_rx_pcs_descrm_pipeln                                                   ("enable"),
		.hssi_10g_rx_pcs_dft_clk_out_sel                                                 ("rx_master_clk"),
		.hssi_10g_rx_pcs_dis_signal_ok                                                   ("dis_signal_ok_dis"),
		.hssi_10g_rx_pcs_dispchk_bypass                                                  ("dispchk_bypass_en"),
		.hssi_10g_rx_pcs_empty_flag_type                                                 ("empty_rd_side"),
		.hssi_10g_rx_pcs_fast_path                                                       ("fast_path_en"),
		.hssi_10g_rx_pcs_fec_clken                                                       ("fec_clk_dis"),
		.hssi_10g_rx_pcs_fec_enable                                                      ("fec_dis"),
		.hssi_10g_rx_pcs_fifo_double_read                                                ("fifo_double_read_dis"),
		.hssi_10g_rx_pcs_fifo_stop_rd                                                    ("n_rd_empty"),
		.hssi_10g_rx_pcs_fifo_stop_wr                                                    ("n_wr_full"),
		.hssi_10g_rx_pcs_force_align                                                     ("force_align_dis"),
		.hssi_10g_rx_pcs_frmsync_bypass                                                  ("frmsync_bypass_en"),
		.hssi_10g_rx_pcs_frmsync_clken                                                   ("frmsync_clk_dis"),
		.hssi_10g_rx_pcs_frmsync_enum_scrm                                               ("enum_scrm_default"),
		.hssi_10g_rx_pcs_frmsync_enum_sync                                               ("enum_sync_default"),
		.hssi_10g_rx_pcs_frmsync_flag_type                                               ("location_only"),
		.hssi_10g_rx_pcs_frmsync_knum_sync                                               ("knum_sync_default"),
		.hssi_10g_rx_pcs_frmsync_mfrm_length                                             (2048),
		.hssi_10g_rx_pcs_frmsync_pipeln                                                  ("frmsync_pipeln_en"),
		.hssi_10g_rx_pcs_full_flag_type                                                  ("full_wr_side"),
		.hssi_10g_rx_pcs_gb_rx_idwidth                                                   ("idwidth_64"),
		.hssi_10g_rx_pcs_gb_rx_odwidth                                                   ("odwidth_66"),
		.hssi_10g_rx_pcs_gbexp_clken                                                     ("gbexp_clk_en"),
		.hssi_10g_rx_pcs_low_latency_en                                                  ("disable"),
		.hssi_10g_rx_pcs_lpbk_mode                                                       ("lpbk_dis"),
		.hssi_10g_rx_pcs_master_clk_sel                                                  ("master_rx_pma_clk"),
		.hssi_10g_rx_pcs_pempty_flag_type                                                ("pempty_rd_side"),
		.hssi_10g_rx_pcs_pfull_flag_type                                                 ("pfull_wr_side"),
		.hssi_10g_rx_pcs_phcomp_rd_del                                                   ("phcomp_rd_del2"),
		.hssi_10g_rx_pcs_pld_if_type                                                     ("reg"),
		.hssi_10g_rx_pcs_prot_mode                                                       ("basic_mode"),
		.hssi_10g_rx_pcs_rand_clken                                                      ("rand_clk_dis"),
		.hssi_10g_rx_pcs_rd_clk_sel                                                      ("rd_rx_pma_clk"),
		.hssi_10g_rx_pcs_rdfifo_clken                                                    ("rdfifo_clk_en"),
		.hssi_10g_rx_pcs_rx_fifo_write_ctrl                                              ("blklock_stops"),
		.hssi_10g_rx_pcs_rx_scrm_width                                                   ("bit64"),
		.hssi_10g_rx_pcs_rx_sh_location                                                  ("msb"),
		.hssi_10g_rx_pcs_rx_signal_ok_sel                                                ("synchronized_ver"),
		.hssi_10g_rx_pcs_rx_sm_bypass                                                    ("rx_sm_bypass_en"),
		.hssi_10g_rx_pcs_rx_sm_hiber                                                     ("rx_sm_hiber_en"),
		.hssi_10g_rx_pcs_rx_sm_pipeln                                                    ("rx_sm_pipeln_en"),
		.hssi_10g_rx_pcs_rx_testbus_sel                                                  ("rx_fifo_testbus1"),
		.hssi_10g_rx_pcs_rx_true_b2b                                                     ("b2b"),
		.hssi_10g_rx_pcs_rxfifo_empty                                                    ("empty_default"),
		.hssi_10g_rx_pcs_rxfifo_full                                                     ("full_default"),
		.hssi_10g_rx_pcs_rxfifo_mode                                                     ("register_mode"),
		.hssi_10g_rx_pcs_rxfifo_pempty                                                   (2),
		.hssi_10g_rx_pcs_rxfifo_pfull                                                    (23),
		.hssi_10g_rx_pcs_stretch_num_stages                                              ("one_stage"),
		.hssi_10g_rx_pcs_sup_mode                                                        ("user_mode"),
		.hssi_10g_rx_pcs_test_mode                                                       ("test_off"),
		.hssi_10g_rx_pcs_wrfifo_clken                                                    ("wrfifo_clk_en"),
		.hssi_10g_rx_pcs_silicon_rev                                                     ("14nm5cr2"),
		.hssi_pldadapt_rx_aib_clk1_sel                                                   ("aib_clk1_pld_pcs_rx_clk_out"),
		.hssi_pldadapt_rx_aib_clk2_sel                                                   ("aib_clk2_pld_pma_clkdiv_rx_user"),
		.hssi_pldadapt_rx_hdpldadapt_aib_fabric_pld_pma_hclk_hz                          (0),
		.hssi_pldadapt_rx_hdpldadapt_aib_fabric_rx_transfer_clk_hz                       (805664062),
		.hssi_pldadapt_rx_asn_bypass_pma_pcie_sw_done                                    ("disable"),
		.hssi_pldadapt_rx_asn_wait_for_dll_reset_cnt                                     (64),
		.hssi_pldadapt_rx_asn_wait_for_fifo_flush_cnt                                    (64),
		.hssi_pldadapt_rx_asn_wait_for_pma_pcie_sw_done_cnt                              (64),
		.hssi_pldadapt_rx_bonding_dft_en                                                 ("dft_dis"),
		.hssi_pldadapt_rx_bonding_dft_val                                                ("dft_0"),
		.hssi_pldadapt_rx_chnl_bonding                                                   ("disable"),
		.hssi_pldadapt_rx_clock_del_measure_enable                                       ("disable"),
		.hssi_pldadapt_rx_hdpldadapt_csr_clk_hz                                          (0),
		.hssi_pldadapt_rx_ctrl_plane_bonding                                             ("individual"),
		.hssi_pldadapt_rx_ds_bypass_pipeln                                               ("ds_bypass_pipeln_dis"),
		.hssi_pldadapt_rx_duplex_mode                                                    ("enable"),
		.hssi_pldadapt_rx_dv_mode                                                        ("dv_mode_en"),
		.hssi_pldadapt_rx_fifo_double_read                                               ("fifo_double_read_en"),
		.hssi_pldadapt_rx_fifo_mode                                                      ("generic_basic"),
		.hssi_pldadapt_rx_fifo_rd_clk_ins_sm_scg_en                                      ("enable"),
		.hssi_pldadapt_rx_fifo_rd_clk_scg_en                                             ("disable"),
		.hssi_pldadapt_rx_fifo_rd_clk_sel                                                ("fifo_rd_clk_pld_rx_clk1"),
		.hssi_pldadapt_rx_fifo_stop_rd                                                   ("n_rd_empty"),
		.hssi_pldadapt_rx_fifo_stop_wr                                                   ("n_wr_full"),
		.hssi_pldadapt_rx_fifo_width                                                     ("fifo_double_width"),
		.hssi_pldadapt_rx_fifo_wr_clk_del_sm_scg_en                                      ("enable"),
		.hssi_pldadapt_rx_fifo_wr_clk_scg_en                                             ("disable"),
		.hssi_pldadapt_rx_fifo_wr_clk_sel                                                ("fifo_wr_clk_rx_transfer_clk"),
		.hssi_pldadapt_rx_free_run_div_clk                                               ("out_of_reset_sync"),
		.hssi_pldadapt_rx_fsr_pld_10g_rx_crc32_err_rst_val                               ("reset_to_zero_crc32"),
		.hssi_pldadapt_rx_fsr_pld_8g_sigdet_out_rst_val                                  ("reset_to_zero_sigdet"),
		.hssi_pldadapt_rx_fsr_pld_ltd_b_rst_val                                          ("reset_to_one_ltdb"),
		.hssi_pldadapt_rx_fsr_pld_ltr_rst_val                                            ("reset_to_zero_ltr"),
		.hssi_pldadapt_rx_fsr_pld_rx_fifo_align_clr_rst_val                              ("reset_to_zero_alignclr"),
		.hssi_pldadapt_rx_gb_rx_idwidth                                                  ("idwidth_64"),
		.hssi_pldadapt_rx_gb_rx_odwidth                                                  ("odwidth_66"),
		.hssi_pldadapt_rx_hip_mode                                                       ("disable_hip"),
		.hssi_pldadapt_rx_hrdrst_align_bypass                                            ("enable"),
		.hssi_pldadapt_rx_hrdrst_dll_lock_bypass                                         ("disable"),
		.hssi_pldadapt_rx_hrdrst_rx_osc_clk_scg_en                                       ("disable"),
		.hssi_pldadapt_rx_hrdrst_user_ctl_en                                             ("disable"),
		.hssi_pldadapt_rx_indv                                                           ("indv_en"),
		.hssi_pldadapt_rx_internal_clk1_sel1                                             ("pma_clks_or_txfiford_post_ct_mux_clk1_mux1"),
		.hssi_pldadapt_rx_internal_clk1_sel2                                             ("pma_clks_clk1_mux2"),
		.hssi_pldadapt_rx_internal_clk2_sel1                                             ("pma_clks_or_rxfifowr_post_ct_mux_clk2_mux1"),
		.hssi_pldadapt_rx_internal_clk2_sel2                                             ("pma_clks_clk2_mux2"),
		.hssi_pldadapt_rx_loopback_mode                                                  ("disable"),
		.hssi_pldadapt_rx_low_latency_en                                                 ("disable"),
		.hssi_pldadapt_rx_lpbk_mode                                                      ("disable"),
		.hssi_pldadapt_rx_osc_clk_scg_en                                                 ("disable"),
		.hssi_pldadapt_rx_phcomp_rd_del                                                  ("phcomp_rd_del2"),
		.hssi_pldadapt_rx_pipe_enable                                                    ("disable"),
		.hssi_pldadapt_rx_pipe_mode                                                      ("disable_pipe"),
		.hssi_pldadapt_rx_hdpldadapt_pld_avmm1_clk_rowclk_hz                             (0),
		.hssi_pldadapt_rx_hdpldadapt_pld_avmm2_clk_rowclk_hz                             (0),
		.hssi_pldadapt_rx_pld_clk1_delay_en                                              ("enable"),
		.hssi_pldadapt_rx_pld_clk1_delay_sel                                             ("delay_path13"),
		.hssi_pldadapt_rx_pld_clk1_inv_en                                                ("disable"),
		.hssi_pldadapt_rx_pld_clk1_sel                                                   ("pld_clk1_dcm"),
		.hssi_pldadapt_rx_hdpldadapt_pld_rx_clk1_dcm_hz                                  (390625000),
		.hssi_pldadapt_rx_hdpldadapt_pld_rx_clk1_rowclk_hz                               (390625000),
		.hssi_pldadapt_rx_hdpldadapt_pld_sclk1_rowclk_hz                                 (0),
		.hssi_pldadapt_rx_hdpldadapt_pld_sclk2_rowclk_hz                                 (0),
		.hssi_pldadapt_rx_pma_hclk_scg_en                                                ("enable"),
		.hssi_pldadapt_rx_powerdown_mode                                                 ("powerup"),
		.hssi_pldadapt_rx_rx_datapath_tb_sel                                             ("cp_bond"),
		.hssi_pldadapt_rx_rx_fastbond_rden                                               ("rden_ds_fast_us_fast"),
		.hssi_pldadapt_rx_rx_fastbond_wren                                               ("wren_ds_del_us_del"),
		.hssi_pldadapt_rx_rx_fifo_power_mode                                             ("full_width_full_depth"),
		.hssi_pldadapt_rx_rx_fifo_read_latency_adjust                                    ("disable"),
		.hssi_pldadapt_rx_rx_fifo_write_ctrl                                             ("blklock_ignore"),
		.hssi_pldadapt_rx_rx_fifo_write_latency_adjust                                   ("disable"),
		.hssi_pldadapt_rx_rx_osc_clock_setting                                           ("osc_clk_div_by1"),
		.hssi_pldadapt_rx_rx_pld_8g_eidleinfersel_polling_bypass                         ("disable"),
		.hssi_pldadapt_rx_rx_pld_pma_eye_monitor_polling_bypass                          ("disable"),
		.hssi_pldadapt_rx_rx_pld_pma_pcie_switch_polling_bypass                          ("disable"),
		.hssi_pldadapt_rx_rx_pld_pma_reser_out_polling_bypass                            ("disable"),
		.hssi_pldadapt_rx_rx_prbs_flags_sr_enable                                        ("disable"),
		.hssi_pldadapt_rx_rx_true_b2b                                                    ("b2b"),
		.hssi_pldadapt_rx_rx_usertest_sel                                                ("enable"),
		.hssi_pldadapt_rx_rxfifo_empty                                                   ("empty_dw"),
		.hssi_pldadapt_rx_rxfifo_full                                                    ("full_non_pc_dw"),
		.hssi_pldadapt_rx_rxfifo_mode                                                    ("rxgeneric_basic"),
		.hssi_pldadapt_rx_rxfifo_pempty                                                  (13),
		.hssi_pldadapt_rx_rxfifo_pfull                                                   (51),
		.hssi_pldadapt_rx_rxfiford_post_ct_sel                                           ("rxfiford_sclk_post_ct"),
		.hssi_pldadapt_rx_rxfifowr_post_ct_sel                                           ("rxfifowr_sclk_post_ct"),
		.hssi_pldadapt_rx_sclk_sel                                                       ("sclk1_rowclk"),
		.hssi_pldadapt_rx_hdpldadapt_speed_grade                                         ("dash_2"),
		.hssi_pldadapt_rx_stretch_num_stages                                             ("two_stage"),
		.hssi_pldadapt_rx_sup_mode                                                       ("user_mode"),
		.hssi_pldadapt_rx_txfiford_post_ct_sel                                           ("txfiford_sclk_post_ct"),
		.hssi_pldadapt_rx_txfifowr_post_ct_sel                                           ("txfifowr_sclk_post_ct"),
		.hssi_pldadapt_rx_us_bypass_pipeln                                               ("us_bypass_pipeln_dis"),
		.hssi_pldadapt_rx_word_align                                                     ("wa_en"),
		.hssi_pldadapt_rx_word_align_enable                                              ("enable"),
		.hssi_pldadapt_rx_silicon_rev                                                    ("14nm5cr2"),
		.hssi_pldadapt_tx_aib_clk1_sel                                                   ("aib_clk1_pld_pcs_tx_clk_out"),
		.hssi_pldadapt_tx_aib_clk2_sel                                                   ("aib_clk2_pld_pma_clkdiv_tx_user"),
		.hssi_pldadapt_tx_hdpldadapt_aib_fabric_pld_pma_hclk_hz                          (0),
		.hssi_pldadapt_tx_hdpldadapt_aib_fabric_pma_aib_tx_clk_hz                        (805664062),
		.hssi_pldadapt_tx_bonding_dft_en                                                 ("dft_dis"),
		.hssi_pldadapt_tx_bonding_dft_val                                                ("dft_0"),
		.hssi_pldadapt_tx_chnl_bonding                                                   ("disable"),
		.hssi_pldadapt_tx_hdpldadapt_csr_clk_hz                                          (0),
		.hssi_pldadapt_tx_ctrl_plane_bonding                                             ("individual"),
		.hssi_pldadapt_tx_ds_bypass_pipeln                                               ("ds_bypass_pipeln_dis"),
		.hssi_pldadapt_tx_duplex_mode                                                    ("enable"),
		.hssi_pldadapt_tx_dv_bond                                                        ("dv_bond_dis"),
		.hssi_pldadapt_tx_dv_gen                                                         ("dv_gen_en"),
		.hssi_pldadapt_tx_fifo_double_write                                              ("fifo_double_write_en"),
		.hssi_pldadapt_tx_fifo_mode                                                      ("generic_basic"),
		.hssi_pldadapt_tx_fifo_rd_clk_frm_gen_scg_en                                     ("enable"),
		.hssi_pldadapt_tx_fifo_rd_clk_scg_en                                             ("disable"),
		.hssi_pldadapt_tx_fifo_rd_clk_sel                                                ("fifo_rd_pma_aib_tx_clk"),
		.hssi_pldadapt_tx_fifo_stop_rd                                                   ("n_rd_empty"),
		.hssi_pldadapt_tx_fifo_stop_wr                                                   ("n_wr_full"),
		.hssi_pldadapt_tx_fifo_width                                                     ("fifo_double_width"),
		.hssi_pldadapt_tx_fifo_wr_clk_scg_en                                             ("disable"),
		.hssi_pldadapt_tx_fpll_shared_direct_async_in_sel                                ("fpll_shared_direct_async_in_rowclk"),
		.hssi_pldadapt_tx_frmgen_burst                                                   ("frmgen_burst_dis"),
		.hssi_pldadapt_tx_frmgen_bypass                                                  ("frmgen_bypass_en"),
		.hssi_pldadapt_tx_frmgen_mfrm_length                                             (2048),
		.hssi_pldadapt_tx_frmgen_pipeln                                                  ("frmgen_pipeln_en"),
		.hssi_pldadapt_tx_frmgen_pyld_ins                                                ("frmgen_pyld_ins_dis"),
		.hssi_pldadapt_tx_frmgen_wordslip                                                ("frmgen_wordslip_dis"),
		.hssi_pldadapt_tx_fsr_hip_fsr_in_bit0_rst_val                                    ("reset_to_one_hfsrin0"),
		.hssi_pldadapt_tx_fsr_hip_fsr_in_bit1_rst_val                                    ("reset_to_one_hfsrin1"),
		.hssi_pldadapt_tx_fsr_hip_fsr_in_bit2_rst_val                                    ("reset_to_one_hfsrin2"),
		.hssi_pldadapt_tx_fsr_hip_fsr_in_bit3_rst_val                                    ("reset_to_zero_hfsrin3"),
		.hssi_pldadapt_tx_fsr_hip_fsr_out_bit0_rst_val                                   ("reset_to_one_hfsrout0"),
		.hssi_pldadapt_tx_fsr_hip_fsr_out_bit1_rst_val                                   ("reset_to_one_hfsrout1"),
		.hssi_pldadapt_tx_fsr_hip_fsr_out_bit2_rst_val                                   ("reset_to_zero_hfsrout2"),
		.hssi_pldadapt_tx_fsr_hip_fsr_out_bit3_rst_val                                   ("reset_to_zero_hfsrout3"),
		.hssi_pldadapt_tx_fsr_mask_tx_pll_rst_val                                        ("reset_to_zero_maskpll"),
		.hssi_pldadapt_tx_fsr_pld_txelecidle_rst_val                                     ("reset_to_zero_txelec"),
		.hssi_pldadapt_tx_gb_tx_idwidth                                                  ("idwidth_66"),
		.hssi_pldadapt_tx_gb_tx_odwidth                                                  ("odwidth_64"),
		.hssi_pldadapt_tx_hip_mode                                                       ("disable_hip"),
		.hssi_pldadapt_tx_hip_osc_clk_scg_en                                             ("enable"),
		.hssi_pldadapt_tx_hrdrst_dcd_cal_done_bypass                                     ("disable"),
		.hssi_pldadapt_tx_hrdrst_rx_osc_clk_scg_en                                       ("disable"),
		.hssi_pldadapt_tx_hrdrst_user_ctl_en                                             ("disable"),
		.hssi_pldadapt_tx_indv                                                           ("indv_en"),
		.hssi_pldadapt_tx_loopback_mode                                                  ("disable"),
		.hssi_pldadapt_tx_low_latency_en                                                 ("disable"),
		.hssi_pldadapt_tx_osc_clk_scg_en                                                 ("disable"),
		.hssi_pldadapt_tx_phcomp_rd_del                                                  ("phcomp_rd_del2"),
		.hssi_pldadapt_tx_pipe_mode                                                      ("disable_pipe"),
		.hssi_pldadapt_tx_hdpldadapt_pld_avmm1_clk_rowclk_hz                             (0),
		.hssi_pldadapt_tx_hdpldadapt_pld_avmm2_clk_rowclk_hz                             (0),
		.hssi_pldadapt_tx_pld_clk1_delay_en                                              ("enable"),
		.hssi_pldadapt_tx_pld_clk1_delay_sel                                             ("delay_path15"),
		.hssi_pldadapt_tx_pld_clk1_inv_en                                                ("disable"),
		.hssi_pldadapt_tx_pld_clk1_sel                                                   ("pld_clk1_dcm"),
		.hssi_pldadapt_tx_pld_clk2_sel                                                   ("pld_clk2_dcm"),
		.hssi_pldadapt_tx_hdpldadapt_pld_sclk1_rowclk_hz                                 (0),
		.hssi_pldadapt_tx_hdpldadapt_pld_sclk2_rowclk_hz                                 (0),
		.hssi_pldadapt_tx_hdpldadapt_pld_tx_clk1_dcm_hz                                  (390625000),
		.hssi_pldadapt_tx_hdpldadapt_pld_tx_clk1_rowclk_hz                               (390625000),
		.hssi_pldadapt_tx_hdpldadapt_pld_tx_clk2_dcm_hz                                  (805664062),
		.hssi_pldadapt_tx_hdpldadapt_pld_tx_clk2_rowclk_hz                               (805664062),
		.hssi_pldadapt_tx_pma_aib_tx_clk_expected_setting                                ("x2"),
		.hssi_pldadapt_tx_powerdown_mode                                                 ("powerup"),
		.hssi_pldadapt_tx_sh_err                                                         ("sh_err_dis"),
		.hssi_pldadapt_tx_hdpldadapt_speed_grade                                         ("dash_2"),
		.hssi_pldadapt_tx_stretch_num_stages                                             ("two_stage"),
		.hssi_pldadapt_tx_sup_mode                                                       ("user_mode"),
		.hssi_pldadapt_tx_tx_datapath_tb_sel                                             ("cp_bond"),
		.hssi_pldadapt_tx_tx_fastbond_rden                                               ("rden_ds_fast_us_fast"),
		.hssi_pldadapt_tx_tx_fastbond_wren                                               ("wren_ds_fast_us_fast"),
		.hssi_pldadapt_tx_tx_fifo_power_mode                                             ("full_width_full_depth"),
		.hssi_pldadapt_tx_tx_fifo_read_latency_adjust                                    ("disable"),
		.hssi_pldadapt_tx_tx_fifo_write_latency_adjust                                   ("disable"),
		.hssi_pldadapt_tx_tx_hip_aib_ssr_in_polling_bypass                               ("disable"),
		.hssi_pldadapt_tx_tx_osc_clock_setting                                           ("osc_clk_div_by1"),
		.hssi_pldadapt_tx_tx_pld_10g_tx_bitslip_polling_bypass                           ("disable"),
		.hssi_pldadapt_tx_tx_pld_8g_tx_boundary_sel_polling_bypass                       ("disable"),
		.hssi_pldadapt_tx_tx_pld_pma_fpll_cnt_sel_polling_bypass                         ("disable"),
		.hssi_pldadapt_tx_tx_pld_pma_fpll_num_phase_shifts_polling_bypass                ("disable"),
		.hssi_pldadapt_tx_tx_usertest_sel                                                ("enable"),
		.hssi_pldadapt_tx_txfifo_empty                                                   ("empty_default"),
		.hssi_pldadapt_tx_txfifo_full                                                    ("full_non_pc_dw"),
		.hssi_pldadapt_tx_txfifo_mode                                                    ("txgeneric_basic"),
		.hssi_pldadapt_tx_txfifo_pempty                                                  (6),
		.hssi_pldadapt_tx_txfifo_pfull                                                   (26),
		.hssi_pldadapt_tx_us_bypass_pipeln                                               ("us_bypass_pipeln_dis"),
		.hssi_pldadapt_tx_word_align_enable                                              ("enable"),
		.hssi_pldadapt_tx_word_mark                                                      ("wm_en"),
		.hssi_pldadapt_tx_silicon_rev                                                    ("14nm5cr2"),
		.cdr_pll_analog_mode                                                             ("user_custom"),
		.cdr_pll_atb_select_control                                                      ("atb_off"),
		.cdr_pll_auto_reset_on                                                           ("auto_reset_off"),
		.cdr_pll_bandwidth_range_high                                                    ("1"),
		.cdr_pll_bandwidth_range_low                                                     ("1"),
		.cdr_pll_bbpd_data_pattern_filter_select                                         ("bbpd_data_pat_off"),
		.cdr_pll_bti_protected                                                           ("false"),
		.cdr_pll_bw_mode                                                                 ("mid_bw"),
		.cdr_pll_bypass_a_edge                                                           ("bypass_a_edge_off"),
		.cdr_pll_cal_vco_count_length                                                    ("sel_8b_count"),
		.cdr_pll_pm_cr2_rx_path_cdr_clock_enable                                         ("cdr_clock_disable"),
		.cdr_pll_cdr_d2a_enb                                                             ("bti_d2a_disable"),
		.cdr_pll_cdr_odi_select                                                          ("sel_cdr"),
		.cdr_pll_cdr_phaselock_mode                                                      ("no_ignore_lock"),
		.cdr_pll_cdr_powerdown_mode                                                      ("power_up"),
		.cdr_pll_chgpmp_current_dn_pd                                                    ("cp_current_pd_dn_setting4"),
		.cdr_pll_chgpmp_current_dn_trim                                                  ("cp_current_trimming_dn_setting0"),
		.cdr_pll_chgpmp_current_pfd                                                      ("cp_current_pfd_setting1"),
		.cdr_pll_chgpmp_current_up_pd                                                    ("cp_current_pd_up_setting4"),
		.cdr_pll_chgpmp_current_up_trim                                                  ("cp_current_trimming_up_setting0"),
		.cdr_pll_chgpmp_dn_pd_trim_double                                                ("normal_dn_trim_current"),
		.cdr_pll_chgpmp_replicate                                                        ("disable_replica_bias_ctrl"),
		.cdr_pll_chgpmp_testmode                                                         ("cp_test_disable"),
		.cdr_pll_chgpmp_up_pd_trim_double                                                ("normal_up_trim_current"),
		.cdr_pll_chgpmp_vccreg                                                           ("vreg_fw0"),
		.cdr_pll_clk0_dfe_tfall_adj                                                      ("clk0_dfe_tf0"),
		.cdr_pll_clk0_dfe_trise_adj                                                      ("clk0_dfe_tr0"),
		.cdr_pll_clk180_dfe_tfall_adj                                                    ("clk180_dfe_tf0"),
		.cdr_pll_clk180_dfe_trise_adj                                                    ("clk180_dfe_tr0"),
		.cdr_pll_clk270_dfe_tfall_adj                                                    ("clk270_dfe_tf0"),
		.cdr_pll_clk270_dfe_trise_adj                                                    ("clk270_dfe_tr0"),
		.cdr_pll_clk90_dfe_tfall_adj                                                     ("clk90_dfe_tf0"),
		.cdr_pll_clk90_dfe_trise_adj                                                     ("clk90_dfe_tr0"),
		.cdr_pll_clklow_mux_select                                                       ("clklow_mux_cdr_fbclk"),
		.cdr_pll_datarate_bps                                                            ("25781250000"),
		.cdr_pll_diag_loopback_enable                                                    ("no_diag_rev_loopback"),
		.cdr_pll_disable_up_dn                                                           ("normal_mode"),
		.cdr_pll_f_max_cmu_out_freq                                                      ("1"),
		.cdr_pll_f_max_m_counter                                                         ("1"),
		.cdr_pll_f_max_pfd                                                               ("350000000"),
		.cdr_pll_f_max_ref                                                               ("800000000"),
		.cdr_pll_f_max_vco                                                               ("14150000000"),
		.cdr_pll_f_min_gt_channel                                                        ("8700000000"),
		.cdr_pll_f_min_pfd                                                               ("25000000"),
		.cdr_pll_f_min_ref                                                               ("25000000"),
		.cdr_pll_f_min_vco                                                               ("7000000000"),
		.cdr_pll_fref_clklow_div                                                         (2),
		.cdr_pll_fref_mux_select                                                         ("fref_mux_cdr_refclk"),
		.cdr_pll_gpon_lck2ref_control                                                    ("gpon_lck2ref_off"),
		.cdr_pll_initial_settings                                                        ("true"),
		.cdr_pll_lck2ref_delay_control                                                   ("lck2ref_delay_2"),
		.cdr_pll_lf_resistor_pd                                                          ("lf_pd_setting3"),
		.cdr_pll_lf_resistor_pfd                                                         ("lf_pfd_setting3"),
		.cdr_pll_lf_ripple_cap                                                           ("lf_no_ripple"),
		.cdr_pll_loop_filter_bias_select                                                 ("lpflt_bias_7"),
		.cdr_pll_loopback_mode                                                           ("loopback_disabled"),
		.cdr_pll_lpd_counter                                                             (1),
		.cdr_pll_lpfd_counter                                                            (2),
		.cdr_pll_ltd_ltr_micro_controller_select                                         ("ltd_ltr_pcs"),
		.cdr_pll_mcnt_div                                                                (20),
		.cdr_pll_n_counter                                                               (2),
		.cdr_pll_ncnt_div                                                                (2),
		.cdr_pll_optimal                                                                 ("true"),
		.cdr_pll_out_freq                                                                ("12890625000"),
		.cdr_pll_pcie_gen                                                                ("non_pcie"),
		.cdr_pll_pd_fastlock_mode                                                        ("fast_lock_disable"),
		.cdr_pll_pd_l_counter                                                            (1),
		.cdr_pll_pfd_l_counter                                                           (2),
		.cdr_pll_position                                                                ("position0"),
		.cdr_pll_power_mode                                                              ("high_perf"),
		.cdr_pll_powermode_ac_bbpd                                                       ("bbpd_ac_on"),
		.cdr_pll_powermode_ac_rvcotop                                                    ("rvcotop_ac_div1"),
		.cdr_pll_powermode_ac_txpll                                                      ("txpll_ac_off"),
		.cdr_pll_powermode_dc_bbpd                                                       ("bbpd_dc_on"),
		.cdr_pll_powermode_dc_rvcotop                                                    ("rvcotop_dc_div1"),
		.cdr_pll_powermode_dc_txpll                                                      ("powerdown_txpll"),
		.cdr_pll_primary_use                                                             ("cdr"),
		.cdr_pll_prot_mode                                                               ("basic_rx"),
		.cdr_pll_reference_clock_frequency                                               ("644531250"),
		.cdr_pll_requires_gt_capable_channel                                             ("true"),
		.cdr_pll_reverse_serial_loopback                                                 ("no_loopback"),
		.cdr_pll_set_cdr_input_freq_range                                                (0),
		.cdr_pll_set_cdr_v2i_enable                                                      ("enable_v2i_bias"),
		.cdr_pll_set_cdr_vco_reset                                                       ("vco_normal"),
		.cdr_pll_set_cdr_vco_speed                                                       (0),
		.cdr_pll_set_cdr_vco_speed_fix                                                   (120),
		.cdr_pll_set_cdr_vco_speed_pciegen3                                              ("cdr_vco_max_speedbin_pciegen3"),
		.cdr_pll_speed_grade                                                             ("e2"),
		.cdr_pll_sup_mode                                                                ("user_mode"),
		.cdr_pll_tx_pll_prot_mode                                                        ("txpll_unused"),
		.cdr_pll_txpll_hclk_driver_enable                                                ("hclk_off"),
		.cdr_pll_rstb                                                                    ("cdr_lf_reset_off"),
		.cdr_pll_pm_cr2_tx_rx_uc_dyn_reconfig                                            ("uc_dyn_reconfig_off"),
		.cdr_pll_uc_ro_cal                                                               ("uc_ro_cal_off"),
		.cdr_pll_vco_bypass                                                              ("false"),
		.cdr_pll_vco_freq                                                                ("12890625000"),
		.cdr_pll_vco_overrange_voltage                                                   ("vco_overrange_off"),
		.cdr_pll_vco_underrange_voltage                                                  ("vco_underange_off"),
		.cdr_pll_vreg_output                                                             ("vccdreg_nominal"),
		.cdr_pll_direct_fb                                                               ("direct_fb"),
		.cdr_pll_iqclk_sel                                                               ("power_down"),
		.cdr_pll_silicon_rev                                                             ("14nm5cr2"),
		.cdr_pll_pma_width                                                               (64),
		.cdr_pll_cgb_div                                                                 (1),
		.cdr_pll_is_cascaded_pll                                                         ("false"),
		.pma_rx_buf_act_isource_disable                                                  ("isrc_dis"),
		.pma_rx_buf_advanced_mode                                                        ("false"),
		.pma_rx_buf_pm_cr2_rx_path_analog_mode                                           ("user_custom"),
		.pma_rx_buf_bodybias_enable                                                      ("bodybias_dis"),
		.pma_rx_buf_bodybias_select                                                      ("bodybias_sel1"),
		.pma_rx_buf_bypass_ctle_rf_cal                                                   ("use_dprio_rfcal"),
		.pma_rx_buf_clk_divrx_en                                                         ("normal_clk"),
		.pma_rx_buf_const_gm_en                                                          ("cgm_en_1"),
		.pma_rx_buf_ctle_ac_gain                                                         (0),
		.pma_rx_buf_ctle_eq_gain                                                         (0),
		.pma_rx_buf_ctle_hires_bypass                                                    ("ctle_hires_en"),
		.pma_rx_buf_ctle_oc_ib_sel                                                       ("ib_oc_bw3"),
		.pma_rx_buf_ctle_oc_sign                                                         ("add_i_2_p_eq"),
		.pma_rx_buf_ctle_rf_cal                                                          (1),
		.pma_rx_buf_ctle_tia_isel                                                        ("ib_tia_bw3"),
		.pma_rx_buf_pm_cr2_tx_rx_cvp_mode                                                ("cvp_off"),
		.pma_rx_buf_datarate_bps                                                         ("25781250000"),
		.pma_rx_buf_pm_cr2_rx_path_datarate_bps                                          ("25781250000"),
		.pma_rx_buf_pm_cr2_rx_path_datawidth                                             (64),
		.pma_rx_buf_diag_lp_en                                                           ("dlp_off"),
		.pma_rx_buf_eq_bw_sel                                                            ("eq_bw_3"),
		.pma_rx_buf_eq_cdgen_sel                                                         ("eq_cdgen_0"),
		.pma_rx_buf_eq_isel                                                              ("eq_isel_1"),
		.pma_rx_buf_eq_sel                                                               ("eq_sel_3"),
		.pma_rx_buf_pm_cr2_rx_path_gt_enabled                                            ("enable"),
		.pma_rx_buf_initial_settings                                                     ("true"),
		.pma_rx_buf_pm_cr2_rx_path_initial_settings                                      ("true"),
		.pma_rx_buf_pm_cr2_rx_path_jtag_hys                                              ("hys_increase_disable"),
		.pma_rx_buf_pm_cr2_rx_path_jtag_lp                                               ("lp_off"),
		.pma_rx_buf_pm_cr2_rx_path_link                                                  ("sr"),
		.pma_rx_buf_xrx_path_xcdr_deser_xcdr_loopback_mode                               ("loopback_disabled"),
		.pma_rx_buf_loopback_modes                                                       ("lpbk_disable"),
		.pma_rx_buf_offset_cancellation_coarse                                           ("coarse_setting_0"),
		.pma_rx_buf_offset_rx_cal_en                                                     ("rx_oc_dis"),
		.pma_rx_buf_optimal                                                              ("true"),
		.pma_rx_buf_pm_cr2_rx_path_optimal                                               ("true"),
		.pma_rx_buf_pm_cr2_tx_rx_pcie_gen                                                ("non_pcie"),
		.pma_rx_buf_pm_cr2_tx_rx_pcie_gen_bitwidth                                       ("pcie_gen3_32b"),
		.pma_rx_buf_pdb_rx                                                               ("normal_rx_on"),
		.pma_rx_buf_pm_cr2_rx_path_pma_rx_divclk_hz                                      ("402832031"),
		.pma_rx_buf_power_mode                                                           ("high_perf"),
		.pma_rx_buf_pm_cr2_rx_path_power_mode                                            ("high_perf"),
		.pma_rx_buf_pm_cr2_rx_path_power_rail_eht                                        (0),
		.pma_rx_buf_power_rail_er                                                        (0),
		.pma_rx_buf_pm_cr2_rx_path_power_rail_er                                         (1120),
		.pma_rx_buf_powermode_ac_ctle                                                    ("ctle_pwr_ac4"),
		.pma_rx_buf_powermode_ac_vcm                                                     ("vcm_pwr_ac3"),
		.pma_rx_buf_powermode_ac_vga                                                     ("vga_pwr_ac_full"),
		.pma_rx_buf_powermode_dc_ctle                                                    ("ctle_pwr_dc1"),
		.pma_rx_buf_powermode_dc_vcm                                                     ("vcm_pwr_dc3"),
		.pma_rx_buf_powermode_dc_vga                                                     ("vga_pwr_dc_full"),
		.pma_rx_buf_prot_mode                                                            ("basic_rx"),
		.pma_rx_buf_pm_cr2_rx_path_prot_mode                                             ("basic_rx"),
		.pma_rx_buf_qpi_afe_en                                                           ("ctle_mode_en"),
		.pma_rx_buf_qpi_enable                                                           ("non_qpi_mode"),
		.pma_rx_buf_refclk_en                                                            ("disable"),
		.pma_rx_buf_rx_atb_select                                                        ("atb_disable"),
		.pma_rx_buf_rx_vga_oc_en                                                         ("vga_cal_off"),
		.pma_rx_buf_sel_vcm_ctle                                                         ("vocm_eq_fixed"),
		.pma_rx_buf_sel_vcm_tia                                                          ("vocm_tia_fixed"),
		.pma_rx_buf_pm_cr2_rx_path_speed_grade                                           ("e2"),
		.pma_rx_buf_sup_mode                                                             ("user_mode"),
		.pma_rx_buf_pm_cr2_rx_path_sup_mode                                              ("user_mode"),
		.pma_rx_buf_term_sel                                                             ("r_r4"),
		.pma_rx_buf_term_sync_bypass                                                     ("bypass_termsync"),
		.pma_rx_buf_term_tri_enable                                                      ("disable_tri"),
		.pma_rx_buf_pm_cr2_tx_rx_testmux_select                                          ("setting0"),
		.pma_rx_buf_tia_sel                                                              ("tia_sel_1"),
		.pma_rx_buf_pm_cr2_rx_path_tile_type                                             ("h"),
		.pma_rx_buf_pm_cr2_rx_path_uc_cal_clk_bypass                                     ("cal_clk_0"),
		.pma_rx_buf_pm_cr2_rx_path_uc_cal_enable                                         ("rx_cal_off"),
		.pma_rx_buf_pm_cr2_tx_rx_uc_odi_eye_left                                         ("uc_odi_eye_left_off"),
		.pma_rx_buf_pm_cr2_tx_rx_uc_odi_eye_right                                        ("uc_odi_eye_right_off"),
		.pma_rx_buf_pm_cr2_rx_path_uc_pcie_sw                                            ("uc_pcie_gen1"),
		.pma_rx_buf_pm_cr2_tx_rx_uc_rx_cal                                               ("uc_rx_cal_on"),
		.pma_rx_buf_vcm_cal_i                                                            (4),
		.pma_rx_buf_vcm_current_add                                                      ("vcm_current_3"),
		.pma_rx_buf_vcm_sel                                                              ("vcm_l0"),
		.pma_rx_buf_vcm_sel_vccref                                                       (6),
		.pma_rx_buf_vga_dc_gain                                                          (0),
		.pma_rx_buf_vga_halfbw_en                                                        ("vga_half_bw_disabled"),
		.pma_rx_buf_vga_ib_max_en                                                        ("vga_ib_max_enable"),
		.pma_rx_buf_vga_mode                                                             ("vga_off"),
		.pma_rx_buf_silicon_rev                                                          ("14nm5cr2"),
		.hssi_adapt_rx_adapter_lpbk_mode                                                 ("disable"),
		.hssi_adapt_rx_hd_hssiadapt_aib_hssi_pld_sclk_hz                                 (0),
		.hssi_adapt_rx_aib_lpbk_mode                                                     ("disable"),
		.hssi_adapt_rx_align_del                                                         ("align_del_dis"),
		.hssi_adapt_rx_asn_bypass_clock_gate                                             ("disable"),
		.hssi_adapt_rx_asn_bypass_pma_pcie_sw_done                                       ("disable"),
		.hssi_adapt_rx_asn_wait_for_clock_gate_cnt                                       (32),
		.hssi_adapt_rx_asn_wait_for_dll_reset_cnt                                        (32),
		.hssi_adapt_rx_asn_wait_for_fifo_flush_cnt                                       (32),
		.hssi_adapt_rx_asn_wait_for_pma_pcie_sw_done_cnt                                 (32),
		.hssi_adapt_rx_async_direct_hip_en                                               ("disable"),
		.hssi_adapt_rx_bonding_dft_en                                                    ("dft_dis"),
		.hssi_adapt_rx_bonding_dft_val                                                   ("dft_0"),
		.hssi_adapt_rx_chnl_bonding                                                      ("disable"),
		.hssi_adapt_rx_clock_del_measure_enable                                          ("disable"),
		.hssi_adapt_rx_control_del                                                       ("control_del_none"),
		.hssi_adapt_rx_hd_hssiadapt_csr_clk_hz                                           (0),
		.hssi_adapt_rx_ctrl_plane_bonding                                                ("individual"),
		.hssi_adapt_rx_datapath_mapping_mode                                             ("map_10g_2x2x_2x1x_fifo"),
		.hssi_adapt_rx_ds_bypass_pipeln                                                  ("ds_bypass_pipeln_dis"),
		.hssi_adapt_rx_duplex_mode                                                       ("enable"),
		.hssi_adapt_rx_dyn_clk_sw_en                                                     ("disable"),
		.hssi_adapt_rx_fifo_double_write                                                 ("fifo_double_write_en"),
		.hssi_adapt_rx_fifo_mode                                                         ("phase_comp"),
		.hssi_adapt_rx_fifo_rd_clk_scg_en                                                ("disable"),
		.hssi_adapt_rx_fifo_rd_clk_sel                                                   ("fifo_rd_pma_aib_rx_clk"),
		.hssi_adapt_rx_fifo_stop_rd                                                      ("rd_empty"),
		.hssi_adapt_rx_fifo_stop_wr                                                      ("n_wr_full"),
		.hssi_adapt_rx_fifo_width                                                        ("fifo_double_width"),
		.hssi_adapt_rx_fifo_wr_clk_scg_en                                                ("disable"),
		.hssi_adapt_rx_fifo_wr_clk_sel                                                   ("fifo_wr_pld_pcs_rx_clk_out"),
		.hssi_adapt_rx_force_align                                                       ("force_align_dis"),
		.hssi_adapt_rx_free_run_div_clk                                                  ("out_of_reset_sync"),
		.hssi_adapt_rx_fsr_pld_10g_rx_crc32_err_rst_val                                  ("reset_to_zero_crc32"),
		.hssi_adapt_rx_fsr_pld_8g_sigdet_out_rst_val                                     ("reset_to_zero_sigdet"),
		.hssi_adapt_rx_fsr_pld_ltd_b_rst_val                                             ("reset_to_one_ltdb"),
		.hssi_adapt_rx_fsr_pld_ltr_rst_val                                               ("reset_to_zero_ltr"),
		.hssi_adapt_rx_fsr_pld_rx_fifo_align_clr_rst_val                                 ("reset_to_zero_alignclr"),
		.hssi_adapt_rx_hd_hssiadapt_hip_aib_clk_2x_hz                                    (0),
		.hssi_adapt_rx_hd_hssiadapt_hip_aib_clk_hz                                       (0),
		.hssi_adapt_rx_hip_mode                                                          ("disable_hip"),
		.hssi_adapt_rx_hrdrst_dcd_cal_done_bypass                                        ("disable"),
		.hssi_adapt_rx_hrdrst_rx_osc_clk_scg_en                                          ("disable"),
		.hssi_adapt_rx_hrdrst_user_ctl_en                                                ("disable"),
		.hssi_adapt_rx_indv                                                              ("indv_en"),
		.hssi_adapt_rx_internal_clk1_sel                                                 ("pld_pma_tx_clk_out_clk1"),
		.hssi_adapt_rx_internal_clk1_sel0                                                ("pma_clks_or_txfifowr_post_ct_or_txfiford_pre_or_post_ct_mux_clk1_mux0"),
		.hssi_adapt_rx_internal_clk1_sel1                                                ("pma_clks_or_txfiford_pre_or_post_ct_mux_clk1_mux1"),
		.hssi_adapt_rx_internal_clk1_sel2                                                ("pma_clks_or_txfiford_pre_ct_mux_clk1_mux2"),
		.hssi_adapt_rx_internal_clk1_sel3                                                ("pma_clks_clk1_mux3"),
		.hssi_adapt_rx_internal_clk2_sel                                                 ("pld_pma_tx_clk_out_clk2"),
		.hssi_adapt_rx_internal_clk2_sel0                                                ("pma_clks_or_rxfiford_post_ct_or_rxfifowr_pre_or_post_ct_mux_clk2_mux0"),
		.hssi_adapt_rx_internal_clk2_sel1                                                ("pma_clks_or_rxfifowr_pre_or_post_ct_mux_clk2_mux1"),
		.hssi_adapt_rx_internal_clk2_sel2                                                ("pma_clks_or_rxfifowr_pre_ct_mux_clk2_mux2"),
		.hssi_adapt_rx_internal_clk2_sel3                                                ("pma_clks_clk2_mux3"),
		.hssi_adapt_rx_loopback_mode                                                     ("loopback_disable"),
		.hssi_adapt_rx_osc_clk_scg_en                                                    ("disable"),
		.hssi_adapt_rx_phcomp_rd_del                                                     ("phcomp_rd_del3"),
		.hssi_adapt_rx_pipe_mode                                                         ("disable_pipe"),
		.hssi_adapt_rx_hd_hssiadapt_pld_pcs_rx_clk_out_hz                                (402832031),
		.hssi_adapt_rx_hd_hssiadapt_pld_pma_hclk_hz                                      (0),
		.hssi_adapt_rx_pma_aib_rx_clk_expected_setting                                   ("x2"),
		.hssi_adapt_rx_hd_hssiadapt_pma_aib_rx_clk_hz                                    (0),
		.hssi_adapt_rx_pma_coreclkin_sel                                                 ("pma_coreclkin_pld_sel"),
		.hssi_adapt_rx_pma_hclk_scg_en                                                   ("enable"),
		.hssi_adapt_rx_powerdown_mode                                                    ("powerup"),
		.hssi_adapt_rx_rx_10g_krfec_rx_diag_data_status_polling_bypass                   ("disable"),
		.hssi_adapt_rx_rx_adp_go_b4txeq_en                                               ("enable"),
		.hssi_adapt_rx_rx_datapath_tb_sel                                                ("cp_bond"),
		.hssi_adapt_rx_rx_eq_iteration                                                   ("cycles_32"),
		.hssi_adapt_rx_rx_fifo_power_mode                                                ("full_width_full_depth"),
		.hssi_adapt_rx_rx_fifo_read_latency_adjust                                       ("disable"),
		.hssi_adapt_rx_rx_fifo_write_latency_adjust                                      ("disable"),
		.hssi_adapt_rx_rx_invalid_no_change                                              ("disable"),
		.hssi_adapt_rx_rx_osc_clock_setting                                              ("osc_clk_div_by1"),
		.hssi_adapt_rx_rx_parity_sel                                                     ("func_sel"),
		.hssi_adapt_rx_rx_pcs_testbus_sel                                                ("direct_tr_tb_bit0_sel"),
		.hssi_adapt_rx_rx_pcspma_testbus_sel                                             ("enable"),
		.hssi_adapt_rx_rx_pld_8g_a1a2_k1k2_flag_polling_bypass                           ("disable"),
		.hssi_adapt_rx_rx_pld_8g_wa_boundary_polling_bypass                              ("disable"),
		.hssi_adapt_rx_rx_pld_pma_pcie_sw_done_polling_bypass                            ("disable"),
		.hssi_adapt_rx_rx_pld_pma_reser_in_polling_bypass                                ("disable"),
		.hssi_adapt_rx_rx_pld_pma_testbus_polling_bypass                                 ("disable"),
		.hssi_adapt_rx_rx_pld_test_data_polling_bypass                                   ("disable"),
		.hssi_adapt_rx_rx_pma_rstn_cycles                                                ("four_cycles"),
		.hssi_adapt_rx_rx_pma_rstn_en                                                    ("disable"),
		.hssi_adapt_rx_rx_post_cursor_en                                                 ("disable"),
		.hssi_adapt_rx_rx_pre_cursor_en                                                  ("disable"),
		.hssi_adapt_rx_rx_rmfflag_stretch_enable                                         ("enable"),
		.hssi_adapt_rx_rx_rmfflag_stretch_num_stages                                     ("rmfflag_two_stage"),
		.hssi_adapt_rx_rx_rxeq_en                                                        ("disable"),
		.hssi_adapt_rx_rx_txeq_en                                                        ("disable"),
		.hssi_adapt_rx_rx_txeq_time                                                      (64),
		.hssi_adapt_rx_rx_use_rxvalid_for_rxeq                                           ("rxvalid"),
		.hssi_adapt_rx_rx_usertest_sel                                                   ("direct_tr_usertest3_sel"),
		.hssi_adapt_rx_rxfifo_empty                                                      ("empty_default"),
		.hssi_adapt_rx_rxfifo_full                                                       ("full_dw"),
		.hssi_adapt_rx_rxfifo_mode                                                       ("rxphase_comp"),
		.hssi_adapt_rx_rxfifo_pempty                                                     (2),
		.hssi_adapt_rx_rxfifo_pfull                                                      (5),
		.hssi_adapt_rx_rxfiford_post_ct_sel                                              ("rxfiford_sclk_post_ct"),
		.hssi_adapt_rx_rxfiford_to_aib_sel                                               ("rxfiford_sclk_to_aib"),
		.hssi_adapt_rx_rxfifowr_post_ct_sel                                              ("rxfifowr_sclk_post_ct"),
		.hssi_adapt_rx_rxfifowr_pre_ct_sel                                               ("rxfifowr_sclk_pre_ct"),
		.hssi_adapt_rx_hd_hssiadapt_speed_grade                                          ("dash_2"),
		.hssi_adapt_rx_stretch_num_stages                                                ("seven_stage"),
		.hssi_adapt_rx_sup_mode                                                          ("user_mode"),
		.hssi_adapt_rx_txeq_clk_scg_en                                                   ("enable"),
		.hssi_adapt_rx_txeq_clk_sel                                                      ("txeq_pld_pcs_rx_clk_out"),
		.hssi_adapt_rx_txeq_mode                                                         ("eq_disable"),
		.hssi_adapt_rx_txeq_rst_sel                                                      ("txeq_pcs_rx_pld_rst_n"),
		.hssi_adapt_rx_txfiford_post_ct_sel                                              ("txfiford_sclk_post_ct"),
		.hssi_adapt_rx_txfiford_pre_ct_sel                                               ("txfiford_sclk_pre_ct"),
		.hssi_adapt_rx_txfifowr_from_aib_sel                                             ("txfifowr_sclk_from_aib"),
		.hssi_adapt_rx_txfifowr_post_ct_sel                                              ("txfifowr_sclk_post_ct"),
		.hssi_adapt_rx_us_bypass_pipeln                                                  ("us_bypass_pipeln_dis"),
		.hssi_adapt_rx_word_align_enable                                                 ("enable"),
		.hssi_adapt_rx_word_mark                                                         ("wm_en"),
		.hssi_adapt_rx_silicon_rev                                                       ("14nm5cr2"),
		.pma_reset_sequencer_rx_path_rstn_overrideb                                      ("use_sequencer"),
		.pma_reset_sequencer_xrx_path_uc_cal_clk_bypass                                  ("cal_clk_0"),
		.pma_reset_sequencer_xrx_path_uc_cal_enable                                      ("rx_cal_off"),
		.pma_reset_sequencer_silicon_rev                                                 ("14nm5cr2"),
		.pma_tx_ser_bti_protected                                                        ("false"),
		.pma_tx_ser_control_clks_divtx_aibtx                                             ("no_dft_control_clkdivtx_clkaibtx"),
		.pma_tx_ser_datarate_bps                                                         ("0"),
		.pma_tx_ser_duty_cycle_correction_mode_ctrl                                      ("dcc_disable"),
		.pma_tx_ser_initial_settings                                                     ("true"),
		.pma_tx_ser_pcie_gen                                                             ("non_pcie"),
		.pma_tx_ser_power_rail_er                                                        (1120),
		.pma_tx_ser_powermode_ac_ser                                                     ("ac_clk_divtx_user_33_jitcomp1p1"),
		.pma_tx_ser_powermode_dc_ser                                                     ("dc_clk_divtx_user_33_jitcomp1p1"),
		.pma_tx_ser_prot_mode                                                            ("basic_tx"),
		.pma_tx_ser_ser_clk_divtx_user_sel                                               ("divtx_user_33"),
		.pma_tx_ser_ser_aibck_enable                                                     ("enable"),
		.pma_tx_ser_ser_aibck_x1_override                                                ("normal"),
		.pma_tx_ser_ser_clk_mon                                                          ("disable_clk_mon"),
		.pma_tx_ser_ser_dftppm_clkselect                                                 ("aib_dftppm"),
		.pma_tx_ser_ser_in_jitcomp                                                       ("jitcomp_on"),
		.pma_tx_ser_ser_powerdown                                                        ("normal_poweron_ser"),
		.pma_tx_ser_ser_preset_bti_en                                                    ("ser_preset_bti_disable"),
		.pma_tx_ser_sup_mode                                                             ("user_mode"),
		.pma_tx_ser_uc_vcc_setting                                                       ("vcc_setting2"),
		.pma_tx_ser_silicon_rev                                                          ("14nm5cr2"),
		.pma_rx_deser_bitslip_bypass                                                     ("bs_bypass_yes"),
		.pma_rx_deser_bti_protected                                                      ("false"),
		.pma_rx_deser_clkdiv_source                                                      ("vco_bypass_normal"),
		.pma_rx_deser_clkdivrx_user_mode                                                 ("clkdivrx_user_div33"),
		.pma_rx_deser_datarate_bps                                                       ("25781250000"),
		.pma_rx_deser_deser_aib_dftppm_en                                                ("disable"),
		.pma_rx_deser_deser_aibck_en                                                     ("enable"),
		.pma_rx_deser_deser_aibck_x1                                                     ("normal"),
		.pma_rx_deser_deser_factor                                                       ("deser_64b"),
		.pma_rx_deser_deser_powerdown                                                    ("deser_power_up"),
		.pma_rx_deser_force_adaptation_outputs                                           ("normal_outputs"),
		.pma_rx_deser_force_clkdiv_for_testing                                           ("normal_clkdiv"),
		.pma_rx_deser_odi_adapt_bti_en                                                   ("deser_bti_disable"),
		.pma_rx_deser_optimal                                                            ("true"),
		.pma_rx_deser_pcie_g3_hclk_en                                                    ("disable_hclk_div2"),
		.pma_rx_deser_pm_cr2_tx_rx_pcie_gen                                              ("non_pcie"),
		.pma_rx_deser_pm_cr2_tx_rx_pcie_gen_bitwidth                                     ("pcie_gen3_32b"),
		.pma_rx_deser_powermode_ac_deser                                                 ("deser_ac_64b_nobs"),
		.pma_rx_deser_powermode_ac_deser_bs                                              ("deser_ac_bs_off"),
		.pma_rx_deser_powermode_dc_deser                                                 ("deser_dc_64b_nobs"),
		.pma_rx_deser_powermode_dc_deser_bs                                              ("powerdown_deser_bs"),
		.pma_rx_deser_prot_mode                                                          ("basic_rx"),
		.pma_rx_deser_rst_n_adapt_odi                                                    ("no_rst_adapt_odi"),
		.pma_rx_deser_sd_clk                                                             ("sd_clk_disabled"),
		.pma_rx_deser_sup_mode                                                           ("user_mode"),
		.pma_rx_deser_tdr_mode                                                           ("select_bbpd_data"),
		.pma_rx_deser_silicon_rev                                                        ("14nm5cr2"),
		.pma_txpath_chnsequencer_pcie_gen                                                ("non_pcie"),
		.pma_txpath_chnsequencer_prot_mode                                               ("basic_tx"),
		.pma_txpath_chnsequencer_sup_mode                                                ("sup_off"),
		.pma_txpath_chnsequencer_txpath_chnseq_enable                                    ("disable"),
		.pma_txpath_chnsequencer_txpath_chnseq_idle_direct_on                            ("cgb_idle_direct_off"),
		.pma_txpath_chnsequencer_txpath_chnseq_stage_select                              (0),
		.pma_txpath_chnsequencer_txpath_chnseq_wakeup_bypass                             ("bypass_off"),
		.pma_txpath_chnsequencer_silicon_rev                                             ("14nm5bcr2ea"),
		.hssi_aibcr_rx_aib_datasel_gr0                                                   ("aib_datasel0_setting0"),
		.hssi_aibcr_rx_aib_datasel_gr1                                                   ("aib_datasel1_setting0"),
		.hssi_aibcr_rx_aib_datasel_gr2                                                   ("aib_datasel2_setting1"),
		.hssi_aibcr_rx_aib_ddrctrl_gr0                                                   ("aib_ddr0_setting1"),
		.hssi_aibcr_rx_aib_ddrctrl_gr1                                                   ("aib_ddr1_setting1"),
		.hssi_aibcr_rx_aib_iinasyncen                                                    ("aib_inasyncen_setting2"),
		.hssi_aibcr_rx_aib_iinclken                                                      ("aib_inclken_setting3"),
		.hssi_aibcr_rx_aib_outctrl_gr0                                                   ("aib_outen0_setting1"),
		.hssi_aibcr_rx_aib_outctrl_gr1                                                   ("aib_outen1_setting1"),
		.hssi_aibcr_rx_aib_outctrl_gr2                                                   ("aib_outen2_setting1"),
		.hssi_aibcr_rx_aib_outctrl_gr3                                                   ("aib_outen3_setting1"),
		.hssi_aibcr_rx_aib_outndrv_r12                                                   ("aib_ndrv12_setting1"),
		.hssi_aibcr_rx_aib_outndrv_r56                                                   ("aib_ndrv56_setting1"),
		.hssi_aibcr_rx_aib_outndrv_r78                                                   ("aib_ndrv78_setting1"),
		.hssi_aibcr_rx_aib_outpdrv_r12                                                   ("aib_pdrv12_setting1"),
		.hssi_aibcr_rx_aib_outpdrv_r56                                                   ("aib_pdrv56_setting1"),
		.hssi_aibcr_rx_aib_outpdrv_r78                                                   ("aib_pdrv78_setting1"),
		.hssi_aibcr_rx_aib_red_rx_shiften                                                ("aib_red_rx_shift_disable"),
		.hssi_aibcr_rx_aib_rx_clkdiv                                                     ("aib_rx_clkdiv_setting1"),
		.hssi_aibcr_rx_aib_rx_dcc_byp                                                    ("aib_rx_dcc_byp_disable"),
		.hssi_aibcr_rx_aib_rx_dcc_byp_iocsr_unused                                       ("aib_rx_dcc_byp_disable_iocsr_unused"),
		.hssi_aibcr_rx_aib_rx_dcc_cont_cal                                               ("aib_rx_dcc_cal_cont"),
		.hssi_aibcr_rx_aib_rx_dcc_cont_cal_iocsr_unused                                  ("aib_rx_dcc_cal_single_iocsr_unused"),
		.hssi_aibcr_rx_aib_rx_dcc_dft                                                    ("aib_rx_dcc_dft_disable"),
		.hssi_aibcr_rx_aib_rx_dcc_dft_sel                                                ("aib_rx_dcc_dft_mode0"),
		.hssi_aibcr_rx_aib_rx_dcc_dll_entest                                             ("aib_rx_dcc_dll_test_disable"),
		.hssi_aibcr_rx_aib_rx_dcc_dy_ctl_static                                          ("aib_rx_dcc_dy_ctl_static_setting1"),
		.hssi_aibcr_rx_aib_rx_dcc_dy_ctlsel                                              ("aib_rx_dcc_dy_ctlsel_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_en                                                     ("aib_rx_dcc_enable"),
		.hssi_aibcr_rx_aib_rx_dcc_en_iocsr_unused                                        ("aib_rx_dcc_disable_iocsr_unused"),
		.hssi_aibcr_rx_aib_rx_dcc_manual_dn                                              ("aib_rx_dcc_manual_dn0"),
		.hssi_aibcr_rx_aib_rx_dcc_manual_up                                              ("aib_rx_dcc_manual_up0"),
		.hssi_aibcr_rx_aib_rx_dcc_rst_prgmnvrt                                           ("aib_rx_dcc_st_rst_prgmnvrt_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_st_core_dn_prgmnvrt                                    ("aib_rx_dcc_st_core_dn_prgmnvrt_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_st_core_up_prgmnvrt                                    ("aib_rx_dcc_st_core_up_prgmnvrt_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_st_core_updnen                                         ("aib_rx_dcc_st_core_updnen_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_st_dftmuxsel                                           ("aib_rx_dcc_st_dftmuxsel_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_st_dly_pst                                             ("aib_rx_dcc_st_dly_pst_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_st_en                                                  ("aib_rx_dcc_st_en_setting1"),
		.hssi_aibcr_rx_aib_rx_dcc_st_lockreq_muxsel                                      ("aib_rx_dcc_st_lockreq_muxsel_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_st_new_dll                                             ("aib_rx_dcc_new_dll_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_st_new_dll2                                            ("aib_rx_dcc_new_dll2_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_st_rst                                                 ("aib_rx_dcc_st_rst_setting0"),
		.hssi_aibcr_rx_aib_rx_dcc_test_clk_pll_en_n                                      ("aib_rx_dcc_test_clk_pll_en_n_disable"),
		.hssi_aibcr_rx_aib_rx_halfcode                                                   ("aib_rx_halfcode_enable"),
		.hssi_aibcr_rx_aib_rx_selflock                                                   ("aib_rx_selflock_enable"),
		.hssi_aibcr_rx_dft_hssitestip_dll_dcc_en                                         ("disable_dft"),
		.hssi_aibcr_rx_op_mode                                                           ("rx_dcc_enable"),
		.hssi_aibcr_rx_powermode_ac                                                      ("rxdatapath_high_speed_pwr"),
		.hssi_aibcr_rx_powermode_dc                                                      ("powerup"),
		.hssi_aibcr_rx_redundancy_en                                                     ("disable"),
		.hssi_aibcr_rx_sup_mode                                                          ("user_mode"),
		.hssi_aibcr_rx_silicon_rev                                                       ("14nm5cr2"),
		.hssi_aibcr_tx_aib_datasel_gr0                                                   ("aib_datasel0_setting0"),
		.hssi_aibcr_tx_aib_datasel_gr1                                                   ("aib_datasel1_setting1"),
		.hssi_aibcr_tx_aib_datasel_gr2                                                   ("aib_datasel2_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_clkdiv                                           ("aib_dllstr_align_clkdiv_setting1"),
		.hssi_aibcr_tx_aib_dllstr_align_dcc_dll_dft_sel                                  ("aib_dllstr_align_dcc_dll_dft_sel_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_dft_ch_muxsel                                    ("aib_dllstr_align_dft_ch_muxsel_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_dly_pst                                          ("aib_dllstr_align_dly_pst_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_dy_ctl_static                                    ("aib_dllstr_align_dy_ctl_static_setting1"),
		.hssi_aibcr_tx_aib_dllstr_align_dy_ctlsel                                        ("aib_dllstr_align_dy_ctlsel_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_entest                                           ("aib_dllstr_align_test_disable"),
		.hssi_aibcr_tx_aib_dllstr_align_halfcode                                         ("aib_dllstr_align_halfcode_enable"),
		.hssi_aibcr_tx_aib_dllstr_align_selflock                                         ("aib_dllstr_align_selflock_enable"),
		.hssi_aibcr_tx_aib_dllstr_align_st_core_dn_prgmnvrt                              ("aib_dllstr_align_st_core_dn_prgmnvrt_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_st_core_up_prgmnvrt                              ("aib_dllstr_align_st_core_up_prgmnvrt_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_st_core_updnen                                   ("aib_dllstr_align_st_core_updnen_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_st_dftmuxsel                                     ("aib_dllstr_align_st_dftmuxsel_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_st_en                                            ("aib_dllstr_align_st_en_setting1"),
		.hssi_aibcr_tx_aib_dllstr_align_st_lockreq_muxsel                                ("aib_dllstr_align_st_lockreq_muxsel_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_st_new_dll                                       ("aib_dllstr_align_new_dll_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_st_new_dll2                                      ("aib_dllstr_align_new_dll2_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_st_rst                                           ("aib_dllstr_align_st_rst_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_st_rst_prgmnvrt                                  ("aib_dllstr_align_st_rst_prgmnvrt_setting0"),
		.hssi_aibcr_tx_aib_dllstr_align_test_clk_pll_en_n                                ("aib_dllstr_align_test_clk_pll_en_n_disable"),
		.hssi_aibcr_tx_aib_inctrl_gr0                                                    ("aib_inctrl0_setting1"),
		.hssi_aibcr_tx_aib_inctrl_gr1                                                    ("aib_inctrl1_setting3"),
		.hssi_aibcr_tx_aib_inctrl_gr2                                                    ("aib_inctrl2_setting2"),
		.hssi_aibcr_tx_aib_inctrl_gr3                                                    ("aib_inctrl3_setting2"),
		.hssi_aibcr_tx_aib_outctrl_gr0                                                   ("aib_outen0_setting1"),
		.hssi_aibcr_tx_aib_outctrl_gr1                                                   ("aib_outen1_setting1"),
		.hssi_aibcr_tx_aib_outctrl_gr2                                                   ("aib_outen2_setting1"),
		.hssi_aibcr_tx_aib_outndrv_r12                                                   ("aib_ndrv12_setting1"),
		.hssi_aibcr_tx_aib_outndrv_r34                                                   ("aib_ndrv34_setting1"),
		.hssi_aibcr_tx_aib_outndrv_r56                                                   ("aib_ndrv56_setting1"),
		.hssi_aibcr_tx_aib_outndrv_r78                                                   ("aib_ndrv78_setting1"),
		.hssi_aibcr_tx_aib_outpdrv_r12                                                   ("aib_pdrv12_setting1"),
		.hssi_aibcr_tx_aib_outpdrv_r34                                                   ("aib_pdrv34_setting1"),
		.hssi_aibcr_tx_aib_outpdrv_r56                                                   ("aib_pdrv56_setting1"),
		.hssi_aibcr_tx_aib_outpdrv_r78                                                   ("aib_pdrv78_setting1"),
		.hssi_aibcr_tx_aib_red_dirclkn_shiften                                           ("aib_red_dirclkn_shift_disable"),
		.hssi_aibcr_tx_aib_red_dirclkp_shiften                                           ("aib_red_dirclkp_shift_disable"),
		.hssi_aibcr_tx_aib_red_drx_shiften                                               ("aib_red_drx_shift_disable"),
		.hssi_aibcr_tx_aib_red_dtx_shiften                                               ("aib_red_dtx_shift_disable"),
		.hssi_aibcr_tx_aib_red_pinp_shiften                                              ("aib_red_pinp_shift_disable"),
		.hssi_aibcr_tx_aib_red_rx_shiften                                                ("aib_red_rx_shift_disable"),
		.hssi_aibcr_tx_aib_red_tx_shiften                                                ("aib_red_tx_shift_disable"),
		.hssi_aibcr_tx_aib_red_txferclkout_shiften                                       ("aib_red_txferclkout_shift_disable"),
		.hssi_aibcr_tx_aib_red_txferclkoutn_shiften                                      ("aib_red_txferclkoutn_shift_disable"),
		.hssi_aibcr_tx_dfd_dll_dcc_en                                                    ("disable_dfd"),
		.hssi_aibcr_tx_dft_hssitestip_dll_dcc_en                                         ("disable_dft"),
		.hssi_aibcr_tx_op_mode                                                           ("tx_dll_enable"),
		.hssi_aibcr_tx_powermode_ac                                                      ("txdatapath_high_speed_pwr"),
		.hssi_aibcr_tx_powermode_dc                                                      ("powerup"),
		.hssi_aibcr_tx_redundancy_en                                                     ("disable"),
		.hssi_aibcr_tx_sup_mode                                                          ("user_mode"),
		.hssi_aibcr_tx_silicon_rev                                                       ("14nm5cr2"),
		.hssi_aibnd_rx_aib_datasel_gr0                                                   ("aib_datasel0_setting0"),
		.hssi_aibnd_rx_aib_datasel_gr1                                                   ("aib_datasel1_setting1"),
		.hssi_aibnd_rx_aib_datasel_gr2                                                   ("aib_datasel2_setting1"),
		.hssi_aibnd_rx_aib_dllstr_align_clkdiv                                           ("aib_dllstr_align_clkdiv_setting1"),
		.hssi_aibnd_rx_aib_dllstr_align_dly_pst                                          ("aib_dllstr_align_dly_pst_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_dy_ctl_static                                    ("aib_dllstr_align_dy_ctl_static_setting1"),
		.hssi_aibnd_rx_aib_dllstr_align_dy_ctlsel                                        ("aib_dllstr_align_dy_ctlsel_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_entest                                           ("aib_dllstr_align_test_disable"),
		.hssi_aibnd_rx_aib_dllstr_align_halfcode                                         ("aib_dllstr_align_halfcode_enable"),
		.hssi_aibnd_rx_aib_dllstr_align_selflock                                         ("aib_dllstr_align_selflock_enable"),
		.hssi_aibnd_rx_aib_dllstr_align_st_core_dn_prgmnvrt                              ("aib_dllstr_align_st_core_dn_prgmnvrt_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_st_core_up_prgmnvrt                              ("aib_dllstr_align_st_core_up_prgmnvrt_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_st_core_updnen                                   ("aib_dllstr_align_st_core_updnen_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_st_dftmuxsel                                     ("aib_dllstr_align_st_dftmuxsel_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_st_en                                            ("aib_dllstr_align_st_en_setting1"),
		.hssi_aibnd_rx_aib_dllstr_align_st_hps_ctrl_en                                   ("aib_dllstr_align_hps_ctrl_en_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_st_lockreq_muxsel                                ("aib_dllstr_align_st_lockreq_muxsel_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_st_new_dll                                       ("aib_dllstr_align_new_dll_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_st_rst                                           ("aib_dllstr_align_st_rst_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_st_rst_prgmnvrt                                  ("aib_dllstr_align_st_rst_prgmnvrt_setting0"),
		.hssi_aibnd_rx_aib_dllstr_align_test_clk_pll_en_n                                ("aib_dllstr_align_test_clk_pll_en_n_disable"),
		.hssi_aibnd_rx_aib_inctrl_gr0                                                    ("aib_inctrl0_setting1"),
		.hssi_aibnd_rx_aib_inctrl_gr1                                                    ("aib_inctrl1_setting3"),
		.hssi_aibnd_rx_aib_inctrl_gr2                                                    ("aib_inctrl2_setting2"),
		.hssi_aibnd_rx_aib_inctrl_gr3                                                    ("aib_inctrl3_setting3"),
		.hssi_aibnd_rx_aib_outctrl_gr0                                                   ("aib_outen0_setting1"),
		.hssi_aibnd_rx_aib_outctrl_gr1                                                   ("aib_outen1_setting1"),
		.hssi_aibnd_rx_aib_outctrl_gr2                                                   ("aib_outen2_setting1"),
		.hssi_aibnd_rx_aib_outndrv_r12                                                   ("aib_ndrv12_setting1"),
		.hssi_aibnd_rx_aib_outndrv_r34                                                   ("aib_ndrv34_setting1"),
		.hssi_aibnd_rx_aib_outndrv_r56                                                   ("aib_ndrv56_setting1"),
		.hssi_aibnd_rx_aib_outndrv_r78                                                   ("aib_ndrv78_setting1"),
		.hssi_aibnd_rx_aib_outpdrv_r12                                                   ("aib_pdrv12_setting1"),
		.hssi_aibnd_rx_aib_outpdrv_r34                                                   ("aib_pdrv34_setting1"),
		.hssi_aibnd_rx_aib_outpdrv_r56                                                   ("aib_pdrv56_setting1"),
		.hssi_aibnd_rx_aib_outpdrv_r78                                                   ("aib_pdrv78_setting1"),
		.hssi_aibnd_rx_aib_red_shift_en                                                  ("aib_red_shift_disable"),
		.hssi_aibnd_rx_dft_hssitestip_dll_dcc_en                                         ("disable_dft"),
		.hssi_aibnd_rx_op_mode                                                           ("rx_dll_enable"),
		.hssi_aibnd_rx_powermode_ac                                                      ("rxdatapath_high_speed_pwr"),
		.hssi_aibnd_rx_powermode_dc                                                      ("rxdatapath_powerup"),
		.hssi_aibnd_rx_redundancy_en                                                     ("disable"),
		.hssi_aibnd_rx_sup_mode                                                          ("user_mode"),
		.hssi_aibnd_rx_silicon_rev                                                       ("14nm5cr2"),
		.hssi_aibnd_tx_aib_datasel_gr0                                                   ("aib_datasel0_setting0"),
		.hssi_aibnd_tx_aib_datasel_gr1                                                   ("aib_datasel1_setting0"),
		.hssi_aibnd_tx_aib_datasel_gr2                                                   ("aib_datasel2_setting1"),
		.hssi_aibnd_tx_aib_datasel_gr3                                                   ("aib_datasel3_setting1"),
		.hssi_aibnd_tx_aib_ddrctrl_gr0                                                   ("aib_ddr0_setting1"),
		.hssi_aibnd_tx_aib_iinasyncen                                                    ("aib_inasyncen_setting2"),
		.hssi_aibnd_tx_aib_iinclken                                                      ("aib_inclken_setting3"),
		.hssi_aibnd_tx_aib_outctrl_gr0                                                   ("aib_outen0_setting1"),
		.hssi_aibnd_tx_aib_outctrl_gr1                                                   ("aib_outen1_setting1"),
		.hssi_aibnd_tx_aib_outctrl_gr2                                                   ("aib_outen2_setting1"),
		.hssi_aibnd_tx_aib_outctrl_gr3                                                   ("aib_outen3_setting1"),
		.hssi_aibnd_tx_aib_outndrv_r34                                                   ("aib_ndrv34_setting1"),
		.hssi_aibnd_tx_aib_outndrv_r56                                                   ("aib_ndrv56_setting1"),
		.hssi_aibnd_tx_aib_outpdrv_r34                                                   ("aib_pdrv34_setting1"),
		.hssi_aibnd_tx_aib_outpdrv_r56                                                   ("aib_pdrv56_setting1"),
		.hssi_aibnd_tx_aib_red_dirclkn_shiften                                           ("aib_red_dirclkn_shift_disable"),
		.hssi_aibnd_tx_aib_red_dirclkp_shiften                                           ("aib_red_dirclkp_shift_disable"),
		.hssi_aibnd_tx_aib_red_drx_shiften                                               ("aib_red_drx_shift_disable"),
		.hssi_aibnd_tx_aib_red_dtx_shiften                                               ("aib_red_dtx_shift_disable"),
		.hssi_aibnd_tx_aib_red_pout_shiften                                              ("aib_red_pout_shift_disable"),
		.hssi_aibnd_tx_aib_red_rx_shiften                                                ("aib_red_rx_shift_disable"),
		.hssi_aibnd_tx_aib_red_tx_shiften                                                ("aib_red_tx_shift_disable"),
		.hssi_aibnd_tx_aib_red_txferclkout_shiften                                       ("aib_red_txferclkout_shift_disable"),
		.hssi_aibnd_tx_aib_red_txferclkoutn_shiften                                      ("aib_red_txferclkoutn_shift_disable"),
		.hssi_aibnd_tx_aib_tx_clkdiv                                                     ("aib_tx_clkdiv_setting1"),
		.hssi_aibnd_tx_aib_tx_dcc_byp                                                    ("aib_tx_dcc_byp_disable"),
		.hssi_aibnd_tx_aib_tx_dcc_byp_iocsr_unused                                       ("aib_tx_dcc_byp_disable_iocsr_unused"),
		.hssi_aibnd_tx_aib_tx_dcc_cont_cal                                               ("aib_tx_dcc_cal_cont"),
		.hssi_aibnd_tx_aib_tx_dcc_cont_cal_iocsr_unused                                  ("aib_tx_dcc_cal_single_iocsr_unused"),
		.hssi_aibnd_tx_aib_tx_dcc_dft                                                    ("aib_tx_dcc_dft_disable"),
		.hssi_aibnd_tx_aib_tx_dcc_dft_sel                                                ("aib_tx_dcc_dft_mode0"),
		.hssi_aibnd_tx_aib_tx_dcc_dll_dft_sel                                            ("aib_tx_dcc_dll_dft_sel_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_dll_entest                                             ("aib_tx_dcc_dll_test_disable"),
		.hssi_aibnd_tx_aib_tx_dcc_dy_ctl_static                                          ("aib_tx_dcc_dy_ctl_static_setting1"),
		.hssi_aibnd_tx_aib_tx_dcc_dy_ctlsel                                              ("aib_tx_dcc_dy_ctlsel_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_en                                                     ("aib_tx_dcc_enable"),
		.hssi_aibnd_tx_aib_tx_dcc_en_iocsr_unused                                        ("aib_tx_dcc_disable_iocsr_unused"),
		.hssi_aibnd_tx_aib_tx_dcc_manual_dn                                              ("aib_tx_dcc_manual_dn0"),
		.hssi_aibnd_tx_aib_tx_dcc_manual_up                                              ("aib_tx_dcc_manual_up0"),
		.hssi_aibnd_tx_aib_tx_dcc_rst_prgmnvrt                                           ("aib_tx_dcc_st_rst_prgmnvrt_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_st_core_dn_prgmnvrt                                    ("aib_tx_dcc_st_core_dn_prgmnvrt_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_st_core_up_prgmnvrt                                    ("aib_tx_dcc_st_core_up_prgmnvrt_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_st_core_updnen                                         ("aib_tx_dcc_st_core_updnen_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_st_dftmuxsel                                           ("aib_tx_dcc_st_dftmuxsel_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_st_dly_pst                                             ("aib_tx_dcc_st_dly_pst_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_st_en                                                  ("aib_tx_dcc_st_en_setting1"),
		.hssi_aibnd_tx_aib_tx_dcc_st_hps_ctrl_en                                         ("aib_tx_dcc_hps_ctrl_en_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_st_lockreq_muxsel                                      ("aib_tx_dcc_st_lockreq_muxsel_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_st_new_dll                                             ("aib_tx_dcc_new_dll_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_st_rst                                                 ("aib_tx_dcc_st_rst_setting0"),
		.hssi_aibnd_tx_aib_tx_dcc_test_clk_pll_en_n                                      ("aib_tx_dcc_test_clk_pll_en_n_disable"),
		.hssi_aibnd_tx_aib_tx_halfcode                                                   ("aib_tx_halfcode_enable"),
		.hssi_aibnd_tx_aib_tx_selflock                                                   ("aib_tx_selflock_enable"),
		.hssi_aibnd_tx_dfd_dll_dcc_en                                                    ("disable_dfd"),
		.hssi_aibnd_tx_dft_hssitestip_dll_dcc_en                                         ("disable_dft"),
		.hssi_aibnd_tx_op_mode                                                           ("tx_dcc_enable"),
		.hssi_aibnd_tx_powermode_ac                                                      ("txdatapath_high_speed_pwr"),
		.hssi_aibnd_tx_powermode_dc                                                      ("txdatapath_powerup"),
		.hssi_aibnd_tx_redundancy_en                                                     ("disable"),
		.hssi_aibnd_tx_sup_mode                                                          ("user_mode"),
		.hssi_aibnd_tx_silicon_rev                                                       ("14nm5cr2"),
		.hssi_pipe_gen3_bypass_rx_detection_enable                                       ("false"),
		.hssi_pipe_gen3_bypass_rx_preset                                                 (0),
		.hssi_pipe_gen3_bypass_rx_preset_enable                                          ("false"),
		.hssi_pipe_gen3_bypass_tx_coefficent                                             (0),
		.hssi_pipe_gen3_bypass_tx_coefficent_enable                                      ("false"),
		.hssi_pipe_gen3_elecidle_delay_g3                                                (0),
		.hssi_pipe_gen3_ind_error_reporting                                              ("dis_ind_error_reporting"),
		.hssi_pipe_gen3_mode                                                             ("disable_pcs"),
		.hssi_pipe_gen3_phy_status_delay_g12                                             (0),
		.hssi_pipe_gen3_phy_status_delay_g3                                              (0),
		.hssi_pipe_gen3_phystatus_rst_toggle_g12                                         ("dis_phystatus_rst_toggle"),
		.hssi_pipe_gen3_phystatus_rst_toggle_g3                                          ("dis_phystatus_rst_toggle_g3"),
		.hssi_pipe_gen3_rate_match_pad_insertion                                         ("dis_rm_fifo_pad_ins"),
		.hssi_pipe_gen3_sup_mode                                                         ("user_mode"),
		.hssi_pipe_gen3_test_out_sel                                                     ("disable_test_out"),
		.hssi_pipe_gen3_silicon_rev                                                      ("14nm5cr2"),
		.hssi_gen3_rx_pcs_block_sync                                                     ("bypass_block_sync"),
		.hssi_gen3_rx_pcs_block_sync_sm                                                  ("disable_blk_sync_sm"),
		.hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn                                          ("disable"),
		.hssi_gen3_rx_pcs_lpbk_force                                                     ("lpbk_frce_dis"),
		.hssi_gen3_rx_pcs_mode                                                           ("disable_pcs"),
		.hssi_gen3_rx_pcs_rate_match_fifo                                                ("bypass_rm_fifo"),
		.hssi_gen3_rx_pcs_rate_match_fifo_latency                                        ("low_latency"),
		.hssi_gen3_rx_pcs_reverse_lpbk                                                   ("rev_lpbk_dis"),
		.hssi_gen3_rx_pcs_rx_b4gb_par_lpbk                                               ("b4gb_par_lpbk_dis"),
		.hssi_gen3_rx_pcs_rx_force_balign                                                ("dis_force_balign"),
		.hssi_gen3_rx_pcs_rx_ins_del_one_skip                                            ("ins_del_one_skip_dis"),
		.hssi_gen3_rx_pcs_rx_num_fixed_pat                                               (0),
		.hssi_gen3_rx_pcs_rx_test_out_sel                                                ("rx_test_out0"),
		.hssi_gen3_rx_pcs_sup_mode                                                       ("user_mode"),
		.hssi_gen3_rx_pcs_silicon_rev                                                    ("14nm5cr2"),
		.hssi_gen3_tx_pcs_mode                                                           ("disable_pcs"),
		.hssi_gen3_tx_pcs_reverse_lpbk                                                   ("rev_lpbk_dis"),
		.hssi_gen3_tx_pcs_sup_mode                                                       ("user_mode"),
		.hssi_gen3_tx_pcs_tx_bitslip                                                     (0),
		.hssi_gen3_tx_pcs_tx_gbox_byp                                                    ("bypass_gbox"),
		.hssi_gen3_tx_pcs_silicon_rev                                                    ("14nm5cr2"),
		.hssi_adapt_tx_aib_clk_sel                                                       ("aib_clk_pma_aib_tx_clk"),
		.hssi_adapt_tx_hd_hssiadapt_aib_hssi_pld_sclk_hz                                 (0),
		.hssi_adapt_tx_hd_hssiadapt_aib_hssi_tx_transfer_clk_hz                          (805664062),
		.hssi_adapt_tx_bonding_dft_en                                                    ("dft_dis"),
		.hssi_adapt_tx_bonding_dft_val                                                   ("dft_0"),
		.hssi_adapt_tx_chnl_bonding                                                      ("disable"),
		.hssi_adapt_tx_hd_hssiadapt_csr_clk_hz                                           (0),
		.hssi_adapt_tx_ctrl_plane_bonding                                                ("individual"),
		.hssi_adapt_tx_datapath_mapping_mode                                             ("map_10g_2x2x_2x1x_fifo"),
		.hssi_adapt_tx_ds_bypass_pipeln                                                  ("ds_bypass_pipeln_dis"),
		.hssi_adapt_tx_duplex_mode                                                       ("enable"),
		.hssi_adapt_tx_dv_gating                                                         ("disable"),
		.hssi_adapt_tx_dyn_clk_sw_en                                                     ("disable"),
		.hssi_adapt_tx_fifo_double_read                                                  ("fifo_double_read_en"),
		.hssi_adapt_tx_fifo_mode                                                         ("phase_comp"),
		.hssi_adapt_tx_fifo_rd_clk_scg_en                                                ("disable"),
		.hssi_adapt_tx_fifo_rd_clk_sel                                                   ("fifo_rd_pld_pcs_tx_clk_out"),
		.hssi_adapt_tx_fifo_ready_bypass                                                 ("disable"),
		.hssi_adapt_tx_fifo_stop_rd                                                      ("rd_empty"),
		.hssi_adapt_tx_fifo_stop_wr                                                      ("wr_full"),
		.hssi_adapt_tx_fifo_width                                                        ("fifo_double_width"),
		.hssi_adapt_tx_fifo_wr_clk_scg_en                                                ("disable"),
		.hssi_adapt_tx_free_run_div_clk                                                  ("out_of_reset_sync"),
		.hssi_adapt_tx_fsr_hip_fsr_in_bit0_rst_val                                       ("reset_to_one_hfsrin0"),
		.hssi_adapt_tx_fsr_hip_fsr_in_bit1_rst_val                                       ("reset_to_one_hfsrin1"),
		.hssi_adapt_tx_fsr_hip_fsr_in_bit2_rst_val                                       ("reset_to_one_hfsrin2"),
		.hssi_adapt_tx_fsr_hip_fsr_in_bit3_rst_val                                       ("reset_to_zero_hfsrin3"),
		.hssi_adapt_tx_fsr_hip_fsr_out_bit0_rst_val                                      ("reset_to_one_hfsrout0"),
		.hssi_adapt_tx_fsr_hip_fsr_out_bit1_rst_val                                      ("reset_to_one_hfsrout1"),
		.hssi_adapt_tx_fsr_hip_fsr_out_bit2_rst_val                                      ("reset_to_zero_hfsrout2"),
		.hssi_adapt_tx_fsr_hip_fsr_out_bit3_rst_val                                      ("reset_to_zero_hfsrout3"),
		.hssi_adapt_tx_fsr_mask_tx_pll_rst_val                                           ("reset_to_zero_maskpll"),
		.hssi_adapt_tx_fsr_pld_txelecidle_rst_val                                        ("reset_to_zero_txelec"),
		.hssi_adapt_tx_hd_hssiadapt_hip_aib_clk_2x_hz                                    (0),
		.hssi_adapt_tx_hd_hssiadapt_hip_aib_clk_hz                                       (0),
		.hssi_adapt_tx_hd_hssiadapt_hip_aib_txeq_clk_out_hz                              (0),
		.hssi_adapt_tx_hip_mode                                                          ("disable_hip"),
		.hssi_adapt_tx_hip_osc_clk_scg_en                                                ("enable"),
		.hssi_adapt_tx_hrdrst_align_bypass                                               ("enable"),
		.hssi_adapt_tx_hrdrst_dcd_cal_done_bypass                                        ("disable"),
		.hssi_adapt_tx_hrdrst_dll_lock_bypass                                            ("disable"),
		.hssi_adapt_tx_hrdrst_rx_osc_clk_scg_en                                          ("disable"),
		.hssi_adapt_tx_hrdrst_user_ctl_en                                                ("disable"),
		.hssi_adapt_tx_indv                                                              ("indv_en"),
		.hssi_adapt_tx_loopback_mode                                                     ("loopback_disable"),
		.hssi_adapt_tx_osc_clk_scg_en                                                    ("disable"),
		.hssi_adapt_tx_phcomp_rd_del                                                     ("phcomp_rd_del2"),
		.hssi_adapt_tx_pipe_mode                                                         ("disable_pipe"),
		.hssi_adapt_tx_hd_hssiadapt_pld_pcs_tx_clk_out_hz                                (402832031),
		.hssi_adapt_tx_hd_hssiadapt_pld_pma_hclk_hz                                      (0),
		.hssi_adapt_tx_pma_aib_tx_clk_expected_setting                                   ("x2"),
		.hssi_adapt_tx_hd_hssiadapt_pma_aib_tx_clk_hz                                    (0),
		.hssi_adapt_tx_powerdown_mode                                                    ("powerup"),
		.hssi_adapt_tx_presethint_bypass                                                 ("enable"),
		.hssi_adapt_tx_qpi_sr_enable                                                     ("enable"),
		.hssi_adapt_tx_rxqpi_pullup_rst_val                                              ("reset_to_zero_rxqpi"),
		.hssi_adapt_tx_hd_hssiadapt_speed_grade                                          ("dash_2"),
		.hssi_adapt_tx_stretch_num_stages                                                ("seven_stage"),
		.hssi_adapt_tx_sup_mode                                                          ("user_mode"),
		.hssi_adapt_tx_tx_datapath_tb_sel                                                ("cp_bond"),
		.hssi_adapt_tx_tx_fastbond_wren                                                  ("wren_ds_del2_us_del2"),
		.hssi_adapt_tx_tx_fifo_power_mode                                                ("full_width_full_depth"),
		.hssi_adapt_tx_tx_fifo_read_latency_adjust                                       ("disable"),
		.hssi_adapt_tx_tx_fifo_write_latency_adjust                                      ("disable"),
		.hssi_adapt_tx_tx_osc_clock_setting                                              ("osc_clk_div_by1"),
		.hssi_adapt_tx_tx_qpi_mode_en                                                    ("disable"),
		.hssi_adapt_tx_tx_rev_lpbk                                                       ("disable"),
		.hssi_adapt_tx_tx_usertest_sel                                                   ("enable"),
		.hssi_adapt_tx_txfifo_empty                                                      ("empty_default"),
		.hssi_adapt_tx_txfifo_full                                                       ("full_dw"),
		.hssi_adapt_tx_txfifo_mode                                                       ("txphase_comp"),
		.hssi_adapt_tx_txfifo_pempty                                                     (2),
		.hssi_adapt_tx_txfifo_pfull                                                      (5),
		.hssi_adapt_tx_txqpi_pulldn_rst_val                                              ("reset_to_zero_txqpid"),
		.hssi_adapt_tx_txqpi_pullup_rst_val                                              ("reset_to_zero_txqpiu"),
		.hssi_adapt_tx_word_align                                                        ("wa_en"),
		.hssi_adapt_tx_word_align_enable                                                 ("enable"),
		.hssi_adapt_tx_silicon_rev                                                       ("14nm5cr2"),
		.hssi_krfec_rx_pcs_blksync_cor_en                                                ("detect"),
		.hssi_krfec_rx_pcs_bypass_gb                                                     ("bypass_dis"),
		.hssi_krfec_rx_pcs_clr_ctrl                                                      ("both_enabled"),
		.hssi_krfec_rx_pcs_ctrl_bit_reverse                                              ("ctrl_bit_reverse_en"),
		.hssi_krfec_rx_pcs_data_bit_reverse                                              ("data_bit_reverse_dis"),
		.hssi_krfec_rx_pcs_dv_start                                                      ("with_blklock"),
		.hssi_krfec_rx_pcs_err_mark_type                                                 ("err_mark_10g"),
		.hssi_krfec_rx_pcs_error_marking_en                                              ("err_mark_dis"),
		.hssi_krfec_rx_pcs_low_latency_en                                                ("disable"),
		.hssi_krfec_rx_pcs_lpbk_mode                                                     ("lpbk_dis"),
		.hssi_krfec_rx_pcs_parity_invalid_enum                                           (8),
		.hssi_krfec_rx_pcs_parity_valid_num                                              (4),
		.hssi_krfec_rx_pcs_pipeln_blksync                                                ("enable"),
		.hssi_krfec_rx_pcs_pipeln_descrm                                                 ("disable"),
		.hssi_krfec_rx_pcs_pipeln_errcorrect                                             ("disable"),
		.hssi_krfec_rx_pcs_pipeln_errtrap_ind                                            ("enable"),
		.hssi_krfec_rx_pcs_pipeln_errtrap_lfsr                                           ("disable"),
		.hssi_krfec_rx_pcs_pipeln_errtrap_loc                                            ("disable"),
		.hssi_krfec_rx_pcs_pipeln_errtrap_pat                                            ("disable"),
		.hssi_krfec_rx_pcs_pipeln_gearbox                                                ("enable"),
		.hssi_krfec_rx_pcs_pipeln_syndrm                                                 ("enable"),
		.hssi_krfec_rx_pcs_pipeln_trans_dec                                              ("disable"),
		.hssi_krfec_rx_pcs_prot_mode                                                     ("disable_mode"),
		.hssi_krfec_rx_pcs_receive_order                                                 ("receive_lsb"),
		.hssi_krfec_rx_pcs_rx_testbus_sel                                                ("overall"),
		.hssi_krfec_rx_pcs_signal_ok_en                                                  ("sig_ok_en"),
		.hssi_krfec_rx_pcs_sup_mode                                                      ("user_mode"),
		.hssi_krfec_rx_pcs_silicon_rev                                                   ("14nm5cr2"),
		.hssi_krfec_tx_pcs_burst_err                                                     ("burst_err_dis"),
		.hssi_krfec_tx_pcs_burst_err_len                                                 ("burst_err_len1"),
		.hssi_krfec_tx_pcs_ctrl_bit_reverse                                              ("ctrl_bit_reverse_en"),
		.hssi_krfec_tx_pcs_data_bit_reverse                                              ("data_bit_reverse_dis"),
		.hssi_krfec_tx_pcs_enc_frame_query                                               ("enc_query_dis"),
		.hssi_krfec_tx_pcs_low_latency_en                                                ("disable"),
		.hssi_krfec_tx_pcs_pipeln_encoder                                                ("enable"),
		.hssi_krfec_tx_pcs_pipeln_scrambler                                              ("enable"),
		.hssi_krfec_tx_pcs_prot_mode                                                     ("disable_mode"),
		.hssi_krfec_tx_pcs_sup_mode                                                      ("user_mode"),
		.hssi_krfec_tx_pcs_transcode_err                                                 ("trans_err_dis"),
		.hssi_krfec_tx_pcs_transmit_order                                                ("transmit_lsb"),
		.hssi_krfec_tx_pcs_tx_testbus_sel                                                ("overall"),
		.hssi_krfec_tx_pcs_silicon_rev                                                   ("14nm5cr2"),
		.hssi_pipe_gen1_2_elec_idle_delay_val                                            (0),
		.hssi_pipe_gen1_2_error_replace_pad                                              ("replace_edb"),
		.hssi_pipe_gen1_2_hip_mode                                                       ("dis_hip"),
		.hssi_pipe_gen1_2_ind_error_reporting                                            ("dis_ind_error_reporting"),
		.hssi_pipe_gen1_2_phystatus_delay_val                                            (0),
		.hssi_pipe_gen1_2_phystatus_rst_toggle                                           ("dis_phystatus_rst_toggle"),
		.hssi_pipe_gen1_2_pipe_byte_de_serializer_en                                     ("dont_care_bds"),
		.hssi_pipe_gen1_2_prot_mode                                                      ("disabled_prot_mode"),
		.hssi_pipe_gen1_2_rpre_emph_a_val                                                (0),
		.hssi_pipe_gen1_2_rpre_emph_b_val                                                (0),
		.hssi_pipe_gen1_2_rpre_emph_c_val                                                (0),
		.hssi_pipe_gen1_2_rpre_emph_d_val                                                (0),
		.hssi_pipe_gen1_2_rpre_emph_e_val                                                (0),
		.hssi_pipe_gen1_2_rvod_sel_a_val                                                 (0),
		.hssi_pipe_gen1_2_rvod_sel_b_val                                                 (0),
		.hssi_pipe_gen1_2_rvod_sel_c_val                                                 (0),
		.hssi_pipe_gen1_2_rvod_sel_d_val                                                 (0),
		.hssi_pipe_gen1_2_rvod_sel_e_val                                                 (0),
		.hssi_pipe_gen1_2_rx_pipe_enable                                                 ("dis_pipe_rx"),
		.hssi_pipe_gen1_2_rxdetect_bypass                                                ("dis_rxdetect_bypass"),
		.hssi_pipe_gen1_2_sup_mode                                                       ("user_mode"),
		.hssi_pipe_gen1_2_tx_pipe_enable                                                 ("dis_pipe_tx"),
		.hssi_pipe_gen1_2_txswing                                                        ("dis_txswing"),
		.hssi_pipe_gen1_2_silicon_rev                                                    ("14nm5cr2"),
		.hssi_common_pld_pcs_interface_dft_clk_out_en                                    ("dft_clk_out_disable"),
		.hssi_common_pld_pcs_interface_dft_clk_out_sel                                   ("teng_rx_dft_clk"),
		.hssi_common_pld_pcs_interface_hrdrstctrl_en                                     ("hrst_dis"),
		.hssi_common_pld_pcs_interface_pcs_testbus_block_sel                             ("pma_if"),
		.hssi_common_pld_pcs_interface_silicon_rev                                       ("14nm5cr2"),
		.hssi_common_pcs_pma_interface_asn_clk_enable                                    ("false"),
		.hssi_common_pcs_pma_interface_asn_enable                                        ("dis_asn"),
		.hssi_common_pcs_pma_interface_block_sel                                         ("eight_g_pcs"),
		.hssi_common_pcs_pma_interface_bypass_early_eios                                 ("true"),
		.hssi_common_pcs_pma_interface_bypass_pcie_switch                                ("true"),
		.hssi_common_pcs_pma_interface_bypass_pma_ltr                                    ("true"),
		.hssi_common_pcs_pma_interface_bypass_ppm_lock                                   ("false"),
		.hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp                            ("true"),
		.hssi_common_pcs_pma_interface_bypass_txdetectrx                                 ("true"),
		.hssi_common_pcs_pma_interface_cdr_control                                       ("dis_cdr_ctrl"),
		.hssi_common_pcs_pma_interface_cid_enable                                        ("dis_cid_mode"),
		.hssi_common_pcs_pma_interface_data_mask_count                                   (0),
		.hssi_common_pcs_pma_interface_data_mask_count_multi                             (0),
		.hssi_common_pcs_pma_interface_dft_observation_clock_selection                   ("dft_clk_obsrv_tx0"),
		.hssi_common_pcs_pma_interface_early_eios_counter                                (0),
		.hssi_common_pcs_pma_interface_force_freqdet                                     ("force_freqdet_dis"),
		.hssi_common_pcs_pma_interface_free_run_clk_enable                               ("false"),
		.hssi_common_pcs_pma_interface_ignore_sigdet_g23                                 ("false"),
		.hssi_common_pcs_pma_interface_pc_en_counter                                     (0),
		.hssi_common_pcs_pma_interface_pc_rst_counter                                    (0),
		.hssi_common_pcs_pma_interface_pcie_hip_mode                                     ("hip_disable"),
		.hssi_common_pcs_pma_interface_ph_fifo_reg_mode                                  ("phfifo_reg_mode_dis"),
		.hssi_common_pcs_pma_interface_phfifo_flush_wait                                 (0),
		.hssi_common_pcs_pma_interface_pipe_if_g3pcs                                     ("pipe_if_8gpcs"),
		.hssi_common_pcs_pma_interface_pma_done_counter                                  (0),
		.hssi_common_pcs_pma_interface_pma_if_dft_en                                     ("dft_dis"),
		.hssi_common_pcs_pma_interface_pma_if_dft_val                                    ("dft_0"),
		.hssi_common_pcs_pma_interface_ppm_cnt_rst                                       ("ppm_cnt_rst_dis"),
		.hssi_common_pcs_pma_interface_ppm_deassert_early                                ("deassert_early_dis"),
		.hssi_common_pcs_pma_interface_ppm_det_buckets                                   ("ppm_300_100_bucket"),
		.hssi_common_pcs_pma_interface_ppm_gen1_2_cnt                                    ("cnt_32k"),
		.hssi_common_pcs_pma_interface_ppm_post_eidle_delay                              ("cnt_200_cycles"),
		.hssi_common_pcs_pma_interface_ppmsel                                            ("ppmsel_1000"),
		.hssi_common_pcs_pma_interface_prot_mode                                         ("other_protocols"),
		.hssi_common_pcs_pma_interface_rxvalid_mask                                      ("rxvalid_mask_dis"),
		.hssi_common_pcs_pma_interface_sigdet_wait_counter                               (0),
		.hssi_common_pcs_pma_interface_sigdet_wait_counter_multi                         (0),
		.hssi_common_pcs_pma_interface_sim_mode                                          ("disable"),
		.hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en                           ("false"),
		.hssi_common_pcs_pma_interface_sup_mode                                          ("user_mode"),
		.hssi_common_pcs_pma_interface_testout_sel                                       ("ppm_det_test"),
		.hssi_common_pcs_pma_interface_wait_clk_on_off_timer                             (0),
		.hssi_common_pcs_pma_interface_wait_pipe_synchronizing                           (0),
		.hssi_common_pcs_pma_interface_wait_send_syncp_fbkp                              (0),
		.hssi_common_pcs_pma_interface_silicon_rev                                       ("14nm5cr2"),
		.hssi_rx_pcs_pma_interface_block_sel                                             ("ten_g_pcs"),
		.hssi_rx_pcs_pma_interface_channel_operation_mode                                ("tx_rx_pair_enabled"),
		.hssi_rx_pcs_pma_interface_clkslip_sel                                           ("pld"),
		.hssi_rx_pcs_pma_interface_lpbk_en                                               ("disable"),
		.hssi_rx_pcs_pma_interface_master_clk_sel                                        ("master_rx_pma_clk"),
		.hssi_rx_pcs_pma_interface_pldif_datawidth_mode                                  ("pldif_data_10bit"),
		.hssi_rx_pcs_pma_interface_pma_dw_rx                                             ("pma_64b_rx"),
		.hssi_rx_pcs_pma_interface_pma_if_dft_en                                         ("dft_dis"),
		.hssi_rx_pcs_pma_interface_pma_if_dft_val                                        ("dft_0"),
		.hssi_rx_pcs_pma_interface_prbs9_dwidth                                          ("prbs9_64b"),
		.hssi_rx_pcs_pma_interface_prbs_clken                                            ("prbs_clk_dis"),
		.hssi_rx_pcs_pma_interface_prbs_ver                                              ("prbs_off"),
		.hssi_rx_pcs_pma_interface_prot_mode_rx                                          ("teng_basic_mode_rx"),
		.hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion                             ("rx_dyn_polinv_dis"),
		.hssi_rx_pcs_pma_interface_rx_lpbk_en                                            ("lpbk_dis"),
		.hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok                               ("force_sig_ok"),
		.hssi_rx_pcs_pma_interface_rx_prbs_mask                                          ("prbsmask128"),
		.hssi_rx_pcs_pma_interface_rx_prbs_mode                                          ("teng_mode"),
		.hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel                             ("sel_sig_det"),
		.hssi_rx_pcs_pma_interface_rx_static_polarity_inversion                          ("rx_stat_polinv_dis"),
		.hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en                                      ("uhsif_lpbk_dis"),
		.hssi_rx_pcs_pma_interface_sup_mode                                              ("user_mode"),
		.hssi_rx_pcs_pma_interface_silicon_rev                                           ("14nm5cr2"),
		.hssi_tx_pcs_pma_interface_bypass_pma_txelecidle                                 ("true"),
		.hssi_tx_pcs_pma_interface_channel_operation_mode                                ("tx_rx_pair_enabled"),
		.hssi_tx_pcs_pma_interface_lpbk_en                                               ("disable"),
		.hssi_tx_pcs_pma_interface_master_clk_sel                                        ("master_tx_pma_clk"),
		.hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx                                 ("other_prot_mode"),
		.hssi_tx_pcs_pma_interface_pldif_datawidth_mode                                  ("pldif_data_10bit"),
		.hssi_tx_pcs_pma_interface_pma_dw_tx                                             ("pma_64b_tx"),
		.hssi_tx_pcs_pma_interface_pma_if_dft_en                                         ("dft_dis"),
		.hssi_tx_pcs_pma_interface_pmagate_en                                            ("pmagate_dis"),
		.hssi_tx_pcs_pma_interface_prbs9_dwidth                                          ("prbs9_64b"),
		.hssi_tx_pcs_pma_interface_prbs_clken                                            ("prbs_clk_dis"),
		.hssi_tx_pcs_pma_interface_prbs_gen_pat                                          ("prbs_gen_dis"),
		.hssi_tx_pcs_pma_interface_prot_mode_tx                                          ("teng_basic_mode_tx"),
		.hssi_tx_pcs_pma_interface_sq_wave_num                                           ("sq_wave_default"),
		.hssi_tx_pcs_pma_interface_sqwgen_clken                                          ("sqwgen_clk_dis"),
		.hssi_tx_pcs_pma_interface_sup_mode                                              ("user_mode"),
		.hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion                             ("tx_dyn_polinv_dis"),
		.hssi_tx_pcs_pma_interface_tx_pma_data_sel                                       ("ten_g_pcs"),
		.hssi_tx_pcs_pma_interface_tx_static_polarity_inversion                          ("tx_stat_polinv_dis"),
		.hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock                       ("uhsif_filt_stepsz_b4lock_2"),
		.hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value                (0),
		.hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock                     ("uhsif_filt_cntthr_b4lock_8"),
		.hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period                          ("uhsif_dcn_test_period_4"),
		.hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable                             ("uhsif_dcn_test_mode_disable"),
		.hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh                          ("uhsif_dzt_cnt_thr_2"),
		.hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable                      ("uhsif_dzt_disable"),
		.hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window                          ("uhsif_dzt_obr_win_16"),
		.hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size                             ("uhsif_dzt_skipsz_4"),
		.hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel                            ("uhsif_index_cram"),
		.hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin                               ("uhsif_dcn_margin_2"),
		.hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value                   (0),
		.hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control                           ("uhsif_dft_dz_det_val_0"),
		.hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control                             ("uhsif_dft_up_val_0"),
		.hssi_tx_pcs_pma_interface_uhsif_enable                                          ("uhsif_disable"),
		.hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock                       ("uhsif_lkd_segsz_aflock_512"),
		.hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock                      ("uhsif_lkd_segsz_b4lock_16"),
		.hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value            (0),
		.hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value           (0),
		.hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value           (0),
		.hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value          (0),
		.hssi_tx_pcs_pma_interface_silicon_rev                                           ("14nm5cr2"),
		.hssi_fifo_rx_pcs_double_read_mode                                               ("double_read_dis"),
		.hssi_fifo_rx_pcs_prot_mode                                                      ("teng_mode"),
		.hssi_fifo_rx_pcs_silicon_rev                                                    ("14nm5cr2"),
		.hssi_fifo_tx_pcs_double_write_mode                                              ("double_write_dis"),
		.hssi_fifo_tx_pcs_prot_mode                                                      ("teng_mode"),
		.hssi_fifo_tx_pcs_silicon_rev                                                    ("14nm5cr2"),
		.pma_cdr_refclk_powerdown_mode                                                   ("powerup"),
		.pma_cdr_refclk_receiver_detect_src                                              ("iqclk_src"),
		.pma_cdr_refclk_silicon_rev                                                      ("14nm5cr2"),
		.pma_cdr_refclk_refclk_select                                                    ("ref_iqclk0"),
		.pma_rx_odi_datarate_bps                                                         ("25781250000"),
		.pma_rx_odi_enable_cdr_lpbk                                                      ("disable_lpbk"),
		.pma_rx_odi_initial_settings                                                     ("true"),
		.pma_rx_odi_monitor_bw_sel                                                       ("bw_1"),
		.pma_rx_odi_optimal                                                              ("true"),
		.pma_rx_odi_phase_steps_64_vs_128                                                ("phase_steps_64"),
		.pma_rx_odi_phase_steps_sel                                                      ("step40"),
		.pma_rx_odi_power_mode                                                           ("high_perf"),
		.pma_rx_odi_prot_mode                                                            ("basic_rx"),
		.pma_rx_odi_xrx_path_x119_rx_path_rstn_overrideb                                 ("use_sequencer"),
		.pma_rx_odi_step_ctrl_sel                                                        ("dprio_mode"),
		.pma_rx_odi_sup_mode                                                             ("user_mode"),
		.pma_rx_odi_vert_threshold                                                       ("vert_0"),
		.pma_rx_odi_vreg_voltage_sel                                                     ("vreg3"),
		.pma_rx_odi_silicon_rev                                                          ("14nm5cr2"),
		.pma_adapt_sequencer_rx_path_rstn_overrideb                                      ("use_sequencer"),
		.pma_adapt_sequencer_silicon_rev                                                 ("14nm5cr2"),
		.pma_adapt_adapt_mode                                                            ("ctle_dfe"),
		.pma_adapt_adp_ac_ctle_cal_win                                                   ("radp_ac_ctle_cal_win_4"),
		.pma_adapt_adp_ac_ctle_cocurrent_mode_sel                                        ("radp_ac_ctle_cocurrent_mode_sel_mode_1"),
		.pma_adapt_adp_ac_ctle_en                                                        ("radp_ac_ctle_en_enable"),
		.pma_adapt_adp_ac_ctle_hold_en                                                   ("radp_ac_ctle_hold_en_not_hold"),
		.pma_adapt_adp_ac_ctle_initial_load                                              ("radp_ac_ctle_initial_load_0"),
		.pma_adapt_adp_ac_ctle_initial_value                                             ("radp_ac_ctle_initial_value_8"),
		.pma_adapt_adp_ac_ctle_mode_sel                                                  ("radp_ac_ctle_mode_sel_concurrent"),
		.pma_adapt_adp_ac_ctle_ph1_win                                                   ("radp_ac_ctle_ph1_win_2p19"),
		.pma_adapt_adp_adapt_control_sel                                                 ("radp_adapt_control_sel_from_cram"),
		.pma_adapt_adp_adapt_start                                                       ("radp_adapt_start_0"),
		.pma_adapt_adp_bist_datapath_en                                                  ("radp_bist_datapath_en_disable"),
		.pma_adapt_adp_bist_errcount_rstn                                                ("radp_bist_errcount_rstn_0"),
		.pma_adapt_adp_bist_mode_sel                                                     ("radp_bist_mode_sel_prbs31"),
		.pma_adapt_adp_clkgate_enb                                                       ("radp_clkgate_enb_disable"),
		.pma_adapt_adp_clkout_div_sel                                                    ("radp_clkout_div_sel_div2_4cycle"),
		.pma_adapt_adp_ctle_bypass_ac                                                    ("radp_ctle_bypass_ac_not_bypass"),
		.pma_adapt_adp_ctle_bypass_dc                                                    ("radp_ctle_bypass_dc_not_bypass"),
		.pma_adapt_adp_dc_ctle_accum_depth                                               (8),
		.pma_adapt_adp_dc_ctle_en                                                        ("radp_dc_ctle_en_enable"),
		.pma_adapt_adp_dc_ctle_hold_en                                                   ("radp_dc_ctle_hold_en_not_hold"),
		.pma_adapt_adp_dc_ctle_initial_load                                              ("radp_dc_ctle_initial_load_0"),
		.pma_adapt_adp_dc_ctle_initial_value                                             ("radp_dc_ctle_initial_value_32"),
		.pma_adapt_adp_dc_ctle_mode0_win_size                                            ("radp_dc_ctle_mode0_win_size_4_taps"),
		.pma_adapt_adp_dc_ctle_mode0_win_start                                           (0),
		.pma_adapt_adp_dc_ctle_mode1_h1_ratio                                            (8),
		.pma_adapt_adp_dc_ctle_mode2_h2_limit                                            (7),
		.pma_adapt_adp_dc_ctle_mode_sel                                                  ("radp_dc_ctle_mode_sel_mode_2"),
		.pma_adapt_adp_dc_ctle_onetime                                                   ("radp_dc_ctle_onetime_disable"),
		.pma_adapt_adp_dc_ctle_onetime_threshold                                         ("radp_dc_ctle_onetime_threshold_256"),
		.pma_adapt_adp_dfe_accum_depth                                                   (8),
		.pma_adapt_adp_dfe_en                                                            ("radp_dfe_en_enable"),
		.pma_adapt_adp_dfe_fxtap_bypass                                                  ("radp_dfe_fxtap_bypass_not_bypass"),
		.pma_adapt_adp_dfe_hold_en                                                       ("radp_dfe_hold_en_not_hold"),
		.pma_adapt_adp_dfe_hold_sel                                                      ("radp_dfe_hold_sel_no"),
		.pma_adapt_adp_dfe_onetime                                                       ("radp_dfe_onetime_disable"),
		.pma_adapt_adp_dfe_onetime_threshold                                             ("radp_dfe_onetime_threshold_2048"),
		.pma_adapt_adp_dfe_tap1_initial_load                                             ("radp_dfe_tap1_initial_load_0"),
		.pma_adapt_adp_dfe_tap1_initial_value                                            ("radp_dfe_tap1_initial_value_0"),
		.pma_adapt_adp_dfe_tap_sel_en                                                    ("radp_dfe_tap_sel_en_no"),
		.pma_adapt_adp_dlev_accum_depth                                                  (6),
		.pma_adapt_adp_dlev_bypass                                                       ("radp_dlev_bypass_not_bypass"),
		.pma_adapt_adp_dlev_en                                                           ("radp_dlev_en_enable"),
		.pma_adapt_adp_dlev_hold_en                                                      ("radp_dlev_hold_en_not_hold"),
		.pma_adapt_adp_dlev_initial_load                                                 ("radp_dlev_initial_load_0"),
		.pma_adapt_adp_dlev_initial_value                                                ("radp_dlev_initial_value_38"),
		.pma_adapt_adp_dlev_onetime                                                      ("radp_dlev_onetime_disable"),
		.pma_adapt_adp_dlev_onetime_threshold                                            ("radp_dlev_onetime_threshold_4096"),
		.pma_adapt_adp_dlev_sel                                                          ("radp_dlev_sel_mux"),
		.pma_adapt_adp_force_freqlock                                                    ("radp_force_freqlock_use"),
		.pma_adapt_adp_frame_capture                                                     ("radp_frame_capture_0"),
		.pma_adapt_adp_frame_en                                                          ("radp_frame_en_disable"),
		.pma_adapt_adp_frame_odi_sel                                                     ("radp_frame_odi_sel_deser_err"),
		.pma_adapt_adp_frame_out_sel                                                     ("radp_frame_out_sel_select_a"),
		.pma_adapt_adp_load_sig_sel                                                      ("radp_load_sig_sel_from_interanl"),
		.pma_adapt_adp_oc_accum_depth                                                    (11),
		.pma_adapt_adp_oc_bypass                                                         ("radp_oc_bypass_bypass"),
		.pma_adapt_adp_oc_en                                                             ("radp_oc_en_disable"),
		.pma_adapt_adp_oc_hold_en                                                        ("radp_oc_hold_en_not_hold"),
		.pma_adapt_adp_oc_initial_load                                                   ("radp_oc_initial_load_0"),
		.pma_adapt_adp_oc_initial_sign                                                   ("radp_oc_initial_sign_0"),
		.pma_adapt_adp_oc_onetime                                                        ("radp_oc_onetime_disable"),
		.pma_adapt_adp_oc_onetime_threshold                                              ("radp_oc_onetime_threshold_1024"),
		.pma_adapt_adp_odi_bit_sel                                                       ("radp_odi_bit_sel_all_bits"),
		.pma_adapt_adp_odi_control_sel                                                   ("radp_odi_control_sel_from_cram"),
		.pma_adapt_adp_odi_count_threshold                                               ("radp_odi_count_threshold_1e6"),
		.pma_adapt_adp_odi_dfe_spec_en                                                   ("radp_odi_dfe_spec_en_enable"),
		.pma_adapt_adp_odi_dlev_sel                                                      ("radp_odi_dlev_sel_0"),
		.pma_adapt_adp_odi_en                                                            ("radp_odi_en_disable"),
		.pma_adapt_adp_odi_mode                                                          ("radp_odi_mode_detect_errdata"),
		.pma_adapt_adp_odi_rstn                                                          ("radp_odi_rstn_1"),
		.pma_adapt_adp_odi_spec_sel                                                      ("radp_odi_spec_sel_0"),
		.pma_adapt_adp_odi_start                                                         ("radp_odi_start_0"),
		.pma_adapt_adp_pat_dlev_sign_avg_win                                             ("radp_pat_dlev_sign_avg_win_2x"),
		.pma_adapt_adp_pat_dlev_sign_force                                               ("radp_pat_dlev_sign_force_determined_by_cram"),
		.pma_adapt_adp_pat_dlev_sign_value                                               ("radp_pat_dlev_sign_value_1"),
		.pma_adapt_adp_pat_spec_sign_avg_win                                             ("radp_pat_spec_sign_avg_win_256"),
		.pma_adapt_adp_pat_spec_sign_force                                               ("radp_pat_spec_sign_force_generated_internally"),
		.pma_adapt_adp_pat_spec_sign_value                                               ("radp_pat_spec_sign_value_0"),
		.pma_adapt_adp_pat_trans_filter                                                  ("radp_pat_trans_filter_5"),
		.pma_adapt_adp_pat_trans_only_en                                                 ("radp_pat_trans_only_en_enable"),
		.pma_adapt_adp_pcie_adp_bypass                                                   ("radp_pcie_adp_bypass_no"),
		.pma_adapt_adp_pcie_eqz                                                          ("radp_pcie_eqz_non_pcie_mode"),
		.pma_adapt_adp_pcie_hold_sel                                                     (0),
		.pma_adapt_adp_pcs_option                                                        ("radp_pcs_option_0"),
		.pma_adapt_adp_po_actslp_ratio                                                   ("radp_po_actslp_ratio_10_percent"),
		.pma_adapt_adp_po_en                                                             ("radp_po_en_disable"),
		.pma_adapt_adp_po_gb_act2slp                                                     ("radp_po_gb_act2slp_288ns"),
		.pma_adapt_adp_po_gb_slp2act                                                     ("radp_po_gb_slp2act_288ns"),
		.pma_adapt_adp_po_initwait                                                       ("radp_po_initwait_10sec"),
		.pma_adapt_adp_po_sleep_win                                                      ("radp_po_sleep_win_2_sec"),
		.pma_adapt_adp_reserved                                                          (0),
		.pma_adapt_adp_rstn                                                              ("radp_rstn_1"),
		.pma_adapt_adp_status_sel                                                        ("radp_status_sel_0"),
		.pma_adapt_adp_tx_accum_depth                                                    (4),
		.pma_adapt_adp_tx_adp_accumulate                                                 ("radp_tx_adp_accumulate_0"),
		.pma_adapt_adp_tx_adp_en                                                         ("radp_tx_adp_en_0"),
		.pma_adapt_adp_tx_up_dn_flip                                                     ("radp_tx_up_dn_flip_0"),
		.pma_adapt_adp_vga_accum_depth                                                   (9),
		.pma_adapt_adp_vga_bypass                                                        ("radp_vga_bypass_not_bypass"),
		.pma_adapt_adp_vga_ctle_low_limit                                                ("radp_vga_ctle_low_limit_4"),
		.pma_adapt_adp_vga_dlev_offset                                                   (4),
		.pma_adapt_adp_vga_dlev_target                                                   (25),
		.pma_adapt_adp_vga_en                                                            ("radp_vga_en_enalbe"),
		.pma_adapt_adp_vga_hold_en                                                       ("radp_vga_hold_en_not_hold"),
		.pma_adapt_adp_vga_initial_load                                                  ("radp_vga_initial_load_0"),
		.pma_adapt_adp_vga_initial_value                                                 ("radp_vga_initial_value_16"),
		.pma_adapt_adp_vga_onetime                                                       ("radp_vga_onetime_disable"),
		.pma_adapt_adp_vga_onetime_threshold                                             ("radp_vga_onetime_threshold_512"),
		.pma_adapt_datarate_bps                                                          ("25781250000"),
		.pma_adapt_initial_settings                                                      ("true"),
		.pma_adapt_odi_mode                                                              ("odi_disable"),
		.pma_adapt_optimal                                                               ("true"),
		.pma_adapt_power_mode                                                            ("powsav_disable"),
		.pma_adapt_prot_mode                                                             ("basic_rx"),
		.pma_adapt_sup_mode                                                              ("user_mode"),
		.pma_adapt_silicon_rev                                                           ("14nm5cr2"),
		.pma_rx_dfe_adapt_bti_en                                                         ("adapt_bti_disable"),
		.pma_rx_dfe_atb_select                                                           ("atb_disable"),
		.pma_rx_dfe_bti_protected                                                        ("false"),
		.pma_rx_dfe_datarate_bps                                                         ("25781250000"),
		.pma_rx_dfe_dfe_bti_en                                                           ("dfe_bti_disable"),
		.pma_rx_dfe_dfe_mode                                                             ("dfe_tap1_15"),
		.pma_rx_dfe_dft_en                                                               ("dft_disable"),
		.pma_rx_dfe_dft_hilospeed_sel                                                    ("dft_osc_lospeed_path"),
		.pma_rx_dfe_dft_osc_sel                                                          ("dft_osc_even"),
		.pma_rx_dfe_h1edge_bti_en                                                        ("h1edge_bti_disable"),
		.pma_rx_dfe_initial_settings                                                     ("true"),
		.pma_rx_dfe_latch_xcouple_disable                                                ("latch_xcouple_disable"),
		.pma_rx_dfe_oc_sa_cdr0e                                                          (0),
		.pma_rx_dfe_oc_sa_cdr0e_sgn                                                      ("oc_sa_cdr0e_sgn_0"),
		.pma_rx_dfe_oc_sa_cdr0o                                                          (0),
		.pma_rx_dfe_oc_sa_cdr0o_sgn                                                      ("oc_sa_cdr0o_sgn_0"),
		.pma_rx_dfe_oc_sa_cdrne                                                          (0),
		.pma_rx_dfe_oc_sa_cdrne_sgn                                                      ("oc_sa_cdrne_sgn_0"),
		.pma_rx_dfe_oc_sa_cdrno                                                          (0),
		.pma_rx_dfe_oc_sa_cdrno_sgn                                                      ("oc_sa_cdrno_sgn_0"),
		.pma_rx_dfe_oc_sa_cdrpe                                                          (0),
		.pma_rx_dfe_oc_sa_cdrpe_sgn                                                      ("oc_sa_cdrpe_sgn_0"),
		.pma_rx_dfe_oc_sa_cdrpo                                                          (0),
		.pma_rx_dfe_oc_sa_cdrpo_sgn                                                      ("oc_sa_cdrpo_sgn_0"),
		.pma_rx_dfe_oc_sa_dne                                                            (0),
		.pma_rx_dfe_oc_sa_dne_sgn                                                        ("oc_sa_dne_sgn_0"),
		.pma_rx_dfe_oc_sa_dno                                                            (0),
		.pma_rx_dfe_oc_sa_dno_sgn                                                        ("oc_sa_dno_sgn_0"),
		.pma_rx_dfe_oc_sa_dpe                                                            (0),
		.pma_rx_dfe_oc_sa_dpe_sgn                                                        ("oc_sa_dpe_sgn_0"),
		.pma_rx_dfe_oc_sa_dpo                                                            (0),
		.pma_rx_dfe_oc_sa_dpo_sgn                                                        ("oc_sa_dpo_sgn_0"),
		.pma_rx_dfe_oc_sa_odie                                                           (0),
		.pma_rx_dfe_oc_sa_odie_sgn                                                       ("oc_sa_odie_sgn_0"),
		.pma_rx_dfe_oc_sa_odio                                                           (0),
		.pma_rx_dfe_oc_sa_odio_sgn                                                       ("oc_sa_odio_sgn_0"),
		.pma_rx_dfe_oc_sa_vrefe                                                          (0),
		.pma_rx_dfe_oc_sa_vrefe_sgn                                                      ("oc_sa_vrefe_sgn_0"),
		.pma_rx_dfe_oc_sa_vrefo                                                          (0),
		.pma_rx_dfe_oc_sa_vrefo_sgn                                                      ("oc_sa_vrefo_sgn_0"),
		.pma_rx_dfe_odi_bti_en                                                           ("odi_bti_disable"),
		.pma_rx_dfe_odi_dlev_sign                                                        ("odi_dlev_pos"),
		.pma_rx_dfe_odi_h1_sign                                                          ("odi_h1_pos"),
		.pma_rx_dfe_optimal                                                              ("true"),
		.pma_rx_dfe_pdb                                                                  ("dfe_enable"),
		.pma_rx_dfe_pdb_edge_pre_h1                                                      ("cdr_pre_h1_enable"),
		.pma_rx_dfe_pdb_edge_pst_h1                                                      ("cdr_pst_h1_enable"),
		.pma_rx_dfe_pdb_tap_10t15                                                        ("tap10t15_dfe_enable"),
		.pma_rx_dfe_pdb_tap_4t9                                                          ("tap4t9_dfe_enable"),
		.pma_rx_dfe_pdb_tapsum                                                           ("tapsum_enable"),
		.pma_rx_dfe_power_mode                                                           ("high_perf"),
		.pma_rx_dfe_prot_mode                                                            ("basic_rx"),
		.pma_rx_dfe_sel_oc_en                                                            ("off_canc_disable"),
		.pma_rx_dfe_sel_probe_tstmx                                                      ("probe_tstmx_none"),
		.pma_rx_dfe_sup_mode                                                             ("user_mode"),
		.pma_rx_dfe_tap10_coeff                                                          (0),
		.pma_rx_dfe_tap10_sgn                                                            ("tap10_sign_0"),
		.pma_rx_dfe_tap11_coeff                                                          (0),
		.pma_rx_dfe_tap11_sgn                                                            ("tap11_sign_0"),
		.pma_rx_dfe_tap12_coeff                                                          (0),
		.pma_rx_dfe_tap12_sgn                                                            ("tap12_sign_0"),
		.pma_rx_dfe_tap13_coeff                                                          (0),
		.pma_rx_dfe_tap13_sgn                                                            ("tap13_sign_0"),
		.pma_rx_dfe_tap14_coeff                                                          (0),
		.pma_rx_dfe_tap14_sgn                                                            ("tap14_sign_0"),
		.pma_rx_dfe_tap15_coeff                                                          (0),
		.pma_rx_dfe_tap15_sgn                                                            ("tap15_sign_0"),
		.pma_rx_dfe_tap1_coeff                                                           (0),
		.pma_rx_dfe_tap1_sgn                                                             ("tap1_sign_0"),
		.pma_rx_dfe_tap2_coeff                                                           (0),
		.pma_rx_dfe_tap2_sgn                                                             ("tap2_sign_0"),
		.pma_rx_dfe_tap3_coeff                                                           (0),
		.pma_rx_dfe_tap3_sgn                                                             ("tap3_sign_0"),
		.pma_rx_dfe_tap4_coeff                                                           (0),
		.pma_rx_dfe_tap4_sgn                                                             ("tap4_sign_0"),
		.pma_rx_dfe_tap5_coeff                                                           (0),
		.pma_rx_dfe_tap5_sgn                                                             ("tap5_sign_0"),
		.pma_rx_dfe_tap6_coeff                                                           (0),
		.pma_rx_dfe_tap6_sgn                                                             ("tap6_sign_0"),
		.pma_rx_dfe_tap7_coeff                                                           (0),
		.pma_rx_dfe_tap7_sgn                                                             ("tap7_sign_0"),
		.pma_rx_dfe_tap8_coeff                                                           (0),
		.pma_rx_dfe_tap8_sgn                                                             ("tap8_sign_0"),
		.pma_rx_dfe_tap9_coeff                                                           (0),
		.pma_rx_dfe_tap9_sgn                                                             ("tap9_sign_0"),
		.pma_rx_dfe_tapsum_bw_sel                                                        ("tapsum_hibw"),
		.pma_rx_dfe_vref_coeff                                                           (0),
		.pma_rx_dfe_silicon_rev                                                          ("14nm5cr2"),
		.pma_rx_sd_link                                                                  ("sr"),
		.pma_rx_sd_optimal                                                               ("true"),
		.pma_rx_sd_power_mode                                                            ("high_perf"),
		.pma_rx_sd_prot_mode                                                             ("basic_rx"),
		.pma_rx_sd_sd_output_off                                                         ("clk_divrx_2"),
		.pma_rx_sd_sd_output_on                                                          ("force_sd_output_on"),
		.pma_rx_sd_sd_pdb                                                                ("sd_off"),
		.pma_rx_sd_sd_threshold                                                          ("sdlv_3"),
		.pma_rx_sd_sup_mode                                                              ("user_mode"),
		.pma_rx_sd_silicon_rev                                                           ("14nm5cr2"),
		.pma_pcie_gen_switch_silicon_rev                                                 ("14nm5cr2")
	) caui4_xcvr_644 (
		.tx_analogreset                    (tx_analogreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   input,    width = 4,       tx_analogreset.tx_analogreset
		.rx_analogreset                    (rx_analogreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   input,    width = 4,       rx_analogreset.rx_analogreset
		.tx_digitalreset                   (tx_digitalreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //   input,    width = 4,      tx_digitalreset.tx_digitalreset
		.rx_digitalreset                   (rx_digitalreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //   input,    width = 4,      rx_digitalreset.rx_digitalreset
		.tx_analogreset_stat               (tx_analogreset_stat),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //  output,    width = 4,  tx_analogreset_stat.tx_analogreset_stat
		.rx_analogreset_stat               (rx_analogreset_stat),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //  output,    width = 4,  rx_analogreset_stat.rx_analogreset_stat
		.tx_digitalreset_stat              (tx_digitalreset_stat),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //  output,    width = 4, tx_digitalreset_stat.tx_digitalreset_stat
		.rx_digitalreset_stat              (rx_digitalreset_stat),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //  output,    width = 4, rx_digitalreset_stat.rx_digitalreset_stat
		.tx_dll_lock                       (tx_dll_lock),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //  output,    width = 4,          tx_dll_lock.tx_dll_lock
		.tx_cal_busy                       (tx_cal_busy),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //  output,    width = 4,          tx_cal_busy.tx_cal_busy
		.rx_cal_busy                       (rx_cal_busy),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //  output,    width = 4,          rx_cal_busy.rx_cal_busy
		.tx_serial_clk0                    (tx_serial_clk0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   input,    width = 4,       tx_serial_clk0.clk
		.rx_cdr_refclk0                    (rx_cdr_refclk0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   input,    width = 1,       rx_cdr_refclk0.clk
		.tx_serial_data                    (tx_serial_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //  output,    width = 4,       tx_serial_data.tx_serial_data
		.rx_serial_data                    (rx_serial_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   input,    width = 4,       rx_serial_data.rx_serial_data
		.rx_seriallpbken                   (rx_seriallpbken),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //   input,    width = 4,      rx_seriallpbken.rx_seriallpbken
		.rx_set_locktodata                 (rx_set_locktodata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //   input,    width = 4,    rx_set_locktodata.rx_set_locktodata
		.rx_set_locktoref                  (rx_set_locktoref),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //   input,    width = 4,     rx_set_locktoref.rx_set_locktoref
		.rx_is_lockedtoref                 (rx_is_lockedtoref),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //  output,    width = 4,    rx_is_lockedtoref.rx_is_lockedtoref
		.rx_is_lockedtodata                (rx_is_lockedtodata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //  output,    width = 4,   rx_is_lockedtodata.rx_is_lockedtodata
		.tx_coreclkin                      (tx_coreclkin),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //   input,    width = 4,         tx_coreclkin.clk
		.rx_coreclkin                      (rx_coreclkin),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //   input,    width = 4,         rx_coreclkin.clk
		.tx_clkout                         (tx_clkout),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //  output,    width = 4,            tx_clkout.clk
		.tx_clkout2                        (tx_clkout2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //  output,    width = 4,           tx_clkout2.clk
		.rx_clkout                         (rx_clkout),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //  output,    width = 4,            rx_clkout.clk
		.rx_clkout2                        (rx_clkout2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //  output,    width = 4,           rx_clkout2.clk
		.rx_pma_iqtxrx_clkout              (rx_pma_iqtxrx_clkout),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //  output,    width = 4, rx_pma_iqtxrx_clkout.clk
		.tx_parallel_data                  ({tx_fifo_wr_en[3],unused_tx_parallel_data[47:41],tx_parallel_data[255:224],unused_tx_parallel_data[40:38],tx_enh_data_valid[3],unused_tx_parallel_data[37:36],tx_control[7:6],tx_parallel_data[223:192],tx_fifo_wr_en[2],unused_tx_parallel_data[35:29],tx_parallel_data[191:160],unused_tx_parallel_data[28:26],tx_enh_data_valid[2],unused_tx_parallel_data[25:24],tx_control[5:4],tx_parallel_data[159:128],tx_fifo_wr_en[1],unused_tx_parallel_data[23:17],tx_parallel_data[127:96],unused_tx_parallel_data[16:14],tx_enh_data_valid[1],unused_tx_parallel_data[13:12],tx_control[3:2],tx_parallel_data[95:64],tx_fifo_wr_en[0],unused_tx_parallel_data[11:5],tx_parallel_data[63:32],unused_tx_parallel_data[4:2],tx_enh_data_valid[0],unused_tx_parallel_data[1:0],tx_control[1:0],tx_parallel_data[31:0]}),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //   input,  width = 320,     tx_parallel_data.tx_parallel_data
		.rx_parallel_data                  ({caui4_xcvr_644_rx_parallel_data[319],caui4_xcvr_644_rx_parallel_data[318:312],caui4_xcvr_644_rx_parallel_data[311:280],caui4_xcvr_644_rx_parallel_data[279:277],caui4_xcvr_644_rx_parallel_data[276],caui4_xcvr_644_rx_parallel_data[275:274],caui4_xcvr_644_rx_parallel_data[273:272],caui4_xcvr_644_rx_parallel_data[271:240],caui4_xcvr_644_rx_parallel_data[239],caui4_xcvr_644_rx_parallel_data[238:232],caui4_xcvr_644_rx_parallel_data[231:200],caui4_xcvr_644_rx_parallel_data[199:197],caui4_xcvr_644_rx_parallel_data[196],caui4_xcvr_644_rx_parallel_data[195:194],caui4_xcvr_644_rx_parallel_data[193:192],caui4_xcvr_644_rx_parallel_data[191:160],caui4_xcvr_644_rx_parallel_data[159],caui4_xcvr_644_rx_parallel_data[158:152],caui4_xcvr_644_rx_parallel_data[151:120],caui4_xcvr_644_rx_parallel_data[119:117],caui4_xcvr_644_rx_parallel_data[116],caui4_xcvr_644_rx_parallel_data[115:114],caui4_xcvr_644_rx_parallel_data[113:112],caui4_xcvr_644_rx_parallel_data[111:80],caui4_xcvr_644_rx_parallel_data[79],caui4_xcvr_644_rx_parallel_data[78:72],caui4_xcvr_644_rx_parallel_data[71:40],caui4_xcvr_644_rx_parallel_data[39:37],caui4_xcvr_644_rx_parallel_data[36],caui4_xcvr_644_rx_parallel_data[35:34],caui4_xcvr_644_rx_parallel_data[33:32],caui4_xcvr_644_rx_parallel_data[31:0]}), //  output,  width = 320,     rx_parallel_data.rx_parallel_data
		.rx_bitslip                        (rx_bitslip),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //   input,    width = 4,           rx_bitslip.rx_bitslip
		.tx_fifo_full                      (tx_fifo_full),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //  output,    width = 4,         tx_fifo_full.tx_fifo_full
		.tx_fifo_empty                     (tx_fifo_empty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //  output,    width = 4,        tx_fifo_empty.tx_fifo_empty
		.tx_fifo_pfull                     (tx_fifo_pfull),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //  output,    width = 4,        tx_fifo_pfull.tx_fifo_pfull
		.tx_fifo_pempty                    (tx_fifo_pempty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //  output,    width = 4,       tx_fifo_pempty.tx_fifo_pempty
		.rx_fifo_full                      (rx_fifo_full),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //  output,    width = 4,         rx_fifo_full.rx_fifo_full
		.rx_fifo_empty                     (rx_fifo_empty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //  output,    width = 4,        rx_fifo_empty.rx_fifo_empty
		.rx_fifo_pfull                     (rx_fifo_pfull),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //  output,    width = 4,        rx_fifo_pfull.rx_fifo_pfull
		.rx_fifo_pempty                    (rx_fifo_pempty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //  output,    width = 4,       rx_fifo_pempty.rx_fifo_pempty
		.rx_fifo_rd_en                     (rx_fifo_rd_en),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //   input,    width = 4,        rx_fifo_rd_en.rx_fifo_rd_en
		.reconfig_clk                      (reconfig_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //   input,    width = 1,         reconfig_clk.clk
		.reconfig_reset                    (reconfig_reset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   input,    width = 1,       reconfig_reset.reset
		.reconfig_write                    (reconfig_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   input,    width = 1,        reconfig_avmm.write
		.reconfig_read                     (reconfig_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //   input,    width = 1,                     .read
		.reconfig_address                  (reconfig_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //   input,   width = 13,                     .address
		.reconfig_writedata                (reconfig_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //   input,   width = 32,                     .writedata
		.reconfig_readdata                 (reconfig_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //  output,   width = 32,                     .readdata
		.reconfig_waitrequest              (reconfig_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //  output,    width = 1,                     .waitrequest
		.tx_aibreset                       (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_aibreset                       (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rcfg_tx_digitalreset_release_ctrl (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // (terminated),                                    
		.tx_transfer_ready                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_transfer_ready                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.osc_transfer_en                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_fifo_ready                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_fifo_ready                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_digitalreset_timeout           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_digitalreset_timeout           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.avmm_busy                         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_serial_clk1                    (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_serial_clk2                    (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_serial_clk3                    (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_bonding_clocks                 (24'b000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      // (terminated),                                    
		.tx_bonding_clocks1                (24'b000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      // (terminated),                                    
		.tx_bonding_clocks2                (24'b000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      // (terminated),                                    
		.tx_bonding_clocks3                (24'b000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      // (terminated),                                    
		.rx_cdr_refclk1                    (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // (terminated),                                    
		.rx_cdr_refclk2                    (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // (terminated),                                    
		.rx_cdr_refclk3                    (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // (terminated),                                    
		.rx_cdr_refclk4                    (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // (terminated),                                    
		.rx_pma_clkslip                    (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_adapt_reset                    (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_adapt_start                    (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_pma_qpipulldn                  (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_pma_qpipulldn                  (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_pma_qpipullup                  (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_pma_rxfound                    (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_pma_txdetectrx                 (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_pma_elecidle                   (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_x2_coreclkin                   (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_clkout_hioint                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_clkout2_hioint                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_clkout_hioint                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_clkout2_hioint                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.delay_measurement_clkout          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.delay_measurement_clkout2         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_pma_iqtxrx_clkout              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.latency_sclk                      (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.clk_delay_sclk                    (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_fifo_latency_pulse             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_fifo_latency_pulse             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_pcs_fifo_latency_pulse         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_pcs_fifo_latency_pulse         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_fifo_latency_adj_ena           (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_fifo_latency_adj_ena           (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_prbs_err_clr                   (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_prbs_done                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_prbs_err                       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_fifo_insert                    (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_fifo_del                       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_fifo_align_clr                 (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_pcs_fifo_full                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_pcs_fifo_empty                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_pcs_fifo_full                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_pcs_fifo_empty                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_std_bitrev_ena                 (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_std_byterev_ena                (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_polinv                         (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_polinv                         (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_std_bitslipboundarysel         (20'b00000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated),                                    
		.rx_std_bitslipboundarysel         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_std_wa_patternalign            (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_std_wa_a1a2size                (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_std_rmfifo_full                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_std_rmfifo_empty               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_std_signaldetect               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_enh_frame                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_enh_frame_burst_en             (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.tx_enh_frame_diag_status          (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       // (terminated),                                    
		.rx_enh_frame                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_enh_frame_lock                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_enh_frame_diag_status          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_enh_crc32_err                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_enh_highber                    (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_enh_highber_clr_cnt            (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_enh_clr_errblk_count           (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated),                                    
		.rx_enh_blk_lock                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_enh_bitslip                    (28'b0000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pipe_sw_done                      (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             // (terminated),                                    
		.pipe_sw                           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pipe_hclk_in                      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // (terminated),                                    
		.pipe_hclk_out                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pipe_rx_eidleinfersel             (12'b000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pipe_rx_elecidle                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pcs_bonding_bot_data_in           (120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     // (terminated),                                    
		.pcs_bonding_bot_data_out          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pcs_bonding_top_data_in           (120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     // (terminated),                                    
		.pcs_bonding_top_data_out          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pld_aib_bond_tx_ds_in             (20'b00000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated),                                    
		.pld_aib_bond_tx_us_in             (20'b00000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated),                                    
		.pld_aib_bond_tx_ds_out            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pld_aib_bond_tx_us_out            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pld_aib_bond_rx_ds_in             (20'b00000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated),                                    
		.pld_aib_bond_rx_us_in             (20'b00000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated),                                    
		.pld_aib_bond_rx_ds_out            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pld_aib_bond_rx_us_out            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hssi_aib_bond_tx_ds_in            (28'b0000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hssi_aib_bond_tx_us_in            (28'b0000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hssi_aib_bond_tx_ds_out           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hssi_aib_bond_tx_us_out           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hssi_aib_bond_rx_ds_in            (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // (terminated),                                    
		.hssi_aib_bond_rx_us_in            (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // (terminated),                                    
		.hssi_aib_bond_rx_ds_out           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hssi_aib_bond_rx_us_out           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hip_aib_data_in                   (404'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         // (terminated),                                    
		.hip_aib_data_out                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hip_pcs_data_in                   (368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             // (terminated),                                    
		.hip_pcs_data_out                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hip_aib_fsr_in                    (16'b0000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // (terminated),                                    
		.hip_aib_ssr_in                    (160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             // (terminated),                                    
		.hip_aib_fsr_out                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hip_aib_ssr_out                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hip_cal_done                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.hip_in_reserved_out               (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       // (terminated),                                    
		.pld_pmaif_mask_tx_pll             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.pldadapt_out_test_data_b10        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.ehip_aib_data_in                  (420'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         // (terminated),                                    
		.ehip_aib_data_out                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.ehip_aib_pld_tx_data_out          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.ehip_pcs_pld_tx_data_in           (588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 // (terminated),                                    
		.ehip_pcs_pld_rx_data_out          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.tx_pldpcs_clkout                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.rx_pldpcs_clkout                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // (terminated),                                    
		.out_pma_aib_tx_clk                ()                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   // (terminated),                                    
	);

	assign rx_parallel_data = { caui4_xcvr_644_rx_parallel_data[311:280], caui4_xcvr_644_rx_parallel_data[271:240], caui4_xcvr_644_rx_parallel_data[231:200], caui4_xcvr_644_rx_parallel_data[191:160], caui4_xcvr_644_rx_parallel_data[151:120], caui4_xcvr_644_rx_parallel_data[111:80], caui4_xcvr_644_rx_parallel_data[71:40], caui4_xcvr_644_rx_parallel_data[31:0] };

	assign unused_rx_parallel_data = { caui4_xcvr_644_rx_parallel_data[318:312], caui4_xcvr_644_rx_parallel_data[279:277], caui4_xcvr_644_rx_parallel_data[275:274], caui4_xcvr_644_rx_parallel_data[238:232], caui4_xcvr_644_rx_parallel_data[199:197], caui4_xcvr_644_rx_parallel_data[195:194], caui4_xcvr_644_rx_parallel_data[158:152], caui4_xcvr_644_rx_parallel_data[119:117], caui4_xcvr_644_rx_parallel_data[115:114], caui4_xcvr_644_rx_parallel_data[78:72], caui4_xcvr_644_rx_parallel_data[39:37], caui4_xcvr_644_rx_parallel_data[35:34] };

	assign rx_data_valid = { caui4_xcvr_644_rx_parallel_data[319], caui4_xcvr_644_rx_parallel_data[239], caui4_xcvr_644_rx_parallel_data[159], caui4_xcvr_644_rx_parallel_data[79] };

	assign rx_control = { caui4_xcvr_644_rx_parallel_data[273:272], caui4_xcvr_644_rx_parallel_data[193:192], caui4_xcvr_644_rx_parallel_data[113:112], caui4_xcvr_644_rx_parallel_data[33:32] };

	assign rx_enh_data_valid = { caui4_xcvr_644_rx_parallel_data[276], caui4_xcvr_644_rx_parallel_data[196], caui4_xcvr_644_rx_parallel_data[116], caui4_xcvr_644_rx_parallel_data[36] };

endmodule
