// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// MLAB based synchronizer of width 16.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_sync16m #(
    parameter SIM_EMULATE = 1'b0
) (
    input din_clk,
    input [15:0] din,
    input dout_clk,
    output [15:0] dout
);

wire [15:0] dout_w;
alt_e100s10_mlab16a1r1w1 m0 (
    .rclk(dout_clk),
    .wclk(din_clk),
    .waddr(1'b0),
    .din(din),
    .raddr(1'b0),
    .dout(dout_w)
);
defparam m0 .SIM_EMULATE = SIM_EMULATE;

generate
genvar i;
for (i=0; i<16; i=i+1)
begin : sync
       alt_e100s10_altera_std_synchronizer_nocut #(
                    .depth(3),
                    .rst_value(16'b0)
            )  synchronizer_nocut_inst  (
                    .clk(dout_clk),
                    .reset_n(1'b1),
                    .din(dout_w[i]),
                    .dout(dout[i])
       );
end
endgenerate

endmodule

