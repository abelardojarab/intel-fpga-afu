// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// 4 bit counter.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_cnt4i #(
    parameter SIM_EMULATE = 1'b0
) (
    input clk,
    input inc,
    output [3:0] dout
);

wire [3:0] dout_w;

alt_e100s10_lut6 t0 (
    .din({6'h0 | dout | ({6{inc}} & 6'h20)}),
    .dout(dout_w[0])
);
defparam t0 .MASK = 64'h55555555aaaaaaaa;
defparam t0 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 t1 (
    .din({6'h0 | dout | ({6{inc}} & 6'h20)}),
    .dout(dout_w[1])
);
defparam t1 .MASK = 64'h66666666cccccccc;
defparam t1 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 t2 (
    .din({6'h0 | dout | ({6{inc}} & 6'h20)}),
    .dout(dout_w[2])
);
defparam t2 .MASK = 64'h78787878f0f0f0f0;
defparam t2 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 t3 (
    .din({6'h0 | dout | ({6{inc}} & 6'h20)}),
    .dout(dout_w[3])
);
defparam t3 .MASK = 64'h7f807f80ff00ff00;
defparam t3 .SIM_EMULATE = SIM_EMULATE;

reg [3:0] dout_r = 4'b0 /* synthesis preserve_syn_only dont_replicate */;
always @(posedge clk) dout_r <= dout_w;
assign dout = dout_r;

endmodule

