// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// Pulse stretch to 16 cycles.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_pulse16 #(
    parameter SIM_EMULATE = 1'b0
) (
    input clk,
    input din,
    output dout
);

reg [4:0] cntr = 5'b0;
wire [5:0] cntr_w;

alt_e100s10_lut6 t0 (
    .din(6'h0 | {cntr,din}),
    .dout(cntr_w[0])
);
defparam t0 .MASK = 64'hbbbbbbbabbbbbbba;
defparam t0 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 t1 (
    .din(6'h0 | {cntr,din}),
    .dout(cntr_w[1])
);
defparam t1 .MASK = 64'h1414141414141414;
defparam t1 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 t2 (
    .din(6'h0 | {cntr,din}),
    .dout(cntr_w[2])
);
defparam t2 .MASK = 64'h1540154015401540;
defparam t2 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 t3 (
    .din(6'h0 | {cntr,din}),
    .dout(cntr_w[3])
);
defparam t3 .MASK = 64'h1555400015554000;
defparam t3 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 t4 (
    .din(6'h0 | {cntr,din}),
    .dout(cntr_w[4])
);
defparam t4 .MASK = 64'h1555555440000000;
defparam t4 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 t5 (
    .din(6'h0 | {cntr,din}),
    .dout(cntr_w[5])
);
defparam t5 .MASK = 64'hfffffffefffffffe;
defparam t5 .SIM_EMULATE = SIM_EMULATE;

reg dout_r = 1'b0;
always @(posedge clk) {dout_r,cntr} <= cntr_w;
assign dout = dout_r;

endmodule

