`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oP/yiOPnyBBP7LuOUq6SHs0gtIFKQ3mpKh7OlSuXqQZGYy0gVTRzLBFPMJffDTtJ
K7/oeYvetaedx1vPQqKVcID4RFPkv+m/67E3/V/qXb0QmtxZAOqHJFnC6FQxSF4N
0D7e6CGiPKdy964BHLIHceIZ8av2uMuqw7Tc5NnKvv4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6224)
rMv3LRhnI25CIQIHpYT/IYo8wpxuuUwZ3Sel9ospi3GsxeeBmC10UoLjv1CwP9fZ
dH8yB12Cboi2rrinxevjvh8V5klIXiV49ueQddsJabB43mxGK6sd7BmleFLKxhSo
uMH02gijZCYXWihvrmqgki9XauKrMpLbwgOOJxtHl9ogpcOsjJtD8/EBmjKE3rAu
nP+BUHZZ6LWMSKvh6bwTjta9wSwP+LZNOuEg3cYPiTqR31U15SUsw/le0wEhntLX
+RSFn0+iST5Hi97+euOzd5lMigT7fj09hLwSLeCQkbNNLU2iY/0MfyGDPA2uY3PB
Ls8P7z2ok6+Zo/OQ1irqIZobUgNZ+2anKePQvBpgA7sXFlgc3I/l61vOzQwAmmbP
pOfrB1JbEqZ1T9LDKGdEbm5sJnEBGri0OiSFkKitVKC9iM8M49JbDkuMR96IDu5I
lAC0qOeQcOaOgRf0PQcfaR3j2DlT7Oto+IkPw/i5GoF9k039+VRiXkpydl+Xsqog
rCtPJphwvQHnImItwlXxVEiA6/V4FL44v+XPBFI4q0PN+fBcpo/z6+dUmMFX0Ifv
Vj3F0Vf38GRSs2Q9OD+Bpag1cBDzUbgVfALCpYGgs34wwFPXwyHQQIwgbrSnc4jn
/86kFTW0/cQdgSWqjBUZGEZ1Jdlk71NVVeoWFSeUzhTvvxs1LvYi9jd8lakFZ9bh
bI8OmkzJTO0dw+ukCMv8w6vXut7CZgoHE1/BzHXC+8gbIfOeWPP3ShL2qcHX6vs7
3NtKdrWmGI4ienge/ckbTk+joouJok73r/LCVDyW1hd7gxU2qtpvt9NyySe6pYiT
fldRV7J37M2x9JfLoK1As0moCJ5OnZDITOEug+6lgk1xho+r3nKyWsF/7e0Wmilb
CdQwmk7AUREzwHlvJy/vVxC1Sh0pWk3ANGy5AVMEb2cYuclFanxK00olZokuPhe1
ZhwOs5VAWdkBnILPRxPkDCODL1RpyoSYc5D8JEeAcSID5EihcA5QlkSu69ec67JI
bJgYqUbvpxqfG/8whJVhSLZvwIC+YX1DVPzH+E/uS0PNIoGQ8PVdy6F9OTX0Z5ZS
QUvqhsJJAeuyOVs7cnALuKG62V4nolvos6oUEwWcuO0VwEhUsQQUN5i0f5gahTOr
cNGs0oP8lDCk0FK7+nAYfnTfzfle8lwSqSvS4oPehuCcbhkAg8rDxCK3+FHzetWw
aWqgIOP9W2uITrahTxupU/3byCECe/NyKjjrM/1IEiIW9hrd6Se/ILj2hcxEcmTS
SF+V0+NOmS4TfEXppl15NzsKinFp98+gpzadHiJJZQjAdSXS+gStD2xs44FpB02d
/i6kYR+Owmz8UA9P+gn7RpxkPglcFYhle6nw9JUsbe+UA9fhb7WfT1T8RtvuF1b3
LskQomkYUPCsYpbAHibjmikWAMYcOZwmpSx+eq12mR9v5aaRU/D1X6ZjIgkcVi4C
9Dcbj1POydxU3l/dXpFObzTCS8N4cRpxu0hpfr9DchAvJ036Y95HGp28WYG5/kqP
LOZht8pu0cie7xHoENW9ai8AZQDToBE9BOBFboUmrWMH9q61BAPBFRKvU/DjjO0M
CBVfIFU4kNvs2MLAobMt/ZjFOjFXIraCd7C8Um7zoExr4Q1VdTfRnGiucAj22/B3
KrPMwOT9v5aIE20TR1obeTsd1FcA8/WaE6d8PitECrIDj+MQnWAhR4k93gDdi62Z
EfKiNfYL45c0OlkkgjRHaVLsr+5QXyfzh1JyvxsJW5RCQZuk6tTCD0lzgMLOwiU+
A2ZKvHC2xTm52c0LT+jj9ULIk6tokQS3c2ILwSxtxPXylajE2icNt/HajBHolBw5
9RQN6f5cNTY6pJ/SexW3vnCDBVbcPsHrJd0YyYxy/IiZit7G7hdboAFRAKROeFdd
1YtIDIotP+gpOpB5gDGHWWhvRK0u+tmPwP4LiKORCRI2GUAshKsxPSD+m5KjXraC
bGAhY703pnjF7rWQeEfq6KPOHq+FenHvlErochNNZhAA0/qI6DZq67DD1GNFl4mH
KdHNnJlG9tecSOsCIgQfm045390WxP/MxyMFZO06KJPx8NjZH27AKFZ5sZ1wYt3j
H9O8kht9LVF5+zoF1nsEMfTc+TJfdIh7sDnAkvn+MqXa3LhbuNtk7SkgrjXwRvW6
XRV8LnQvUhvN13cgd2NQAgujYjkXeaSvllrqI3tMvzYmusb8aHMwXITkgnHQeo1Y
sb27H/H57SS9NSmWNh9xyUgLK9uOYKNaTPi+itbn+Wjodu5OLxu3f0amcugaKx4F
PpbhlXkRKMZsyAUJlBrvoWpmwFAp9sSFZBZLF7C+dy/dwuZjd2dovwieC+9Z3kEj
7uCfVbUd9uJtM+VwcrRaZ7JD6NrtMxdBZ+8LE8QkIVeIlBOZWpQyzXSN+biFbwOj
SAE6FJAFCgE0dehnItAPhhSdlxG03qebETKdCLv27e4pDlBXZfbTRmv1baMIudU6
/FnxokET9cfjoTpuw7hbB56l/bnw+1TndfyXJDldcT7GizbCruQr2e0MFzGvlZu9
OEI3GUMB1YoI996LW3pQnHJ5Ive5l/aEtdkzz8V4+tXf677qug2exxHhF7p2l5m0
5QLtMhZDlAbh6ZkEEovcYd4UQyp94+cMUDPzP8j0Aa1zjJJhh7NNRJs1F5Uvgpw3
UKNGojojt7/lMcd0KZsKgJ0v5V5zAX1l3HsUqpNrH+xKiqd0C8pZt0wga/GPzk6/
klzCr273fz9PFcZ6Mo2NDM8a0bIFygOqlcmyTJEG7lAWaVjeVPlC3EhpgFYbjWsy
D8vBPJXxnAoyAmsWwO8yD4P7mqMs1CcF9L0b1f5HYcwn1jUqX6GrUe2mdPBje63u
RoxHgMcykjgpUHrL8zP0+HXh4v3/hv4peJx4gJaVyA15ejGLXDXXb2Z4WPyrLug5
tCjzxnc8zAMaA+vTx/RYIWYq+Xy7lhqeer3LiZtwOrnojBQNfNj9zRy3FGSg327N
7YiCfX93ejKD5qDeXiZDggo+KVLM+tfdySNSrt3lde6v3f4JAPHKgCmktPZELrui
QX8pDe8HofsZNQarxb4hVD6PyzzhlPZYgc7+Qp4NXjG0aWpIy74T6GrbgN8ksyHj
qxfFHDU6DTdUoybVHWJV/mkAk78qQRwtcBGl6f4umfXOUJdiTYeqECV0ctpuUo2D
0XfA/FB1N6MFpcrheXeH3rLzuB41unwo07ADLWftJpt5lQbS8xuloS0iK+qU1eSU
zNUZNvu3qmt1u66tEuVbdYpces+SaKSPEYrYReziHtTMAczAYD7UurtJ18IUtmoA
Hbz6YYWhxM+RdSK1oCogexRtxC9UlrCayxVnPY8kE8+MqbHik87ZN+qKN4ELaVTG
am9Kg7YHRNMuIU+/409KdI3i5duKG78eNuAqCPxwF8toLYpaLa5FjJ8K7H5ZceIV
8Dm92BAkBSwG89THZyMWivpeEg3FBgLMhYlNylPfw/jX8Lo4I15iLyG6XVu5YNef
68q4icG549ZDCeNsuqww3N6djNzReCmn+G+j7vo/q9mf9oCFjwYaXtNwpLb1fVZQ
P2Q2aSSEWFu/wA2r04bPo3AxevC7gZf1hl5lIf0TE3khUawLi30UjF8eVW+qvEbD
Oaz4HKhlHqI7WD3xP4r/VNonxJbkR9EBxBoP5wb8KiyrzuT21CKH1Tymak7OiXTw
L8IvvA+csoECUn2T5a5uhWLr3bBAME8LKjq4FjxoBfUakrA/zxCIsGcRtzN+yqL2
Se9iNQ7dciKOkQ2YwDe2c/N8AgSS82gRdSrXHFfrhOzEW3WJBZS/x9TgkufV39Be
aFflLgZfL7D8vFUdMzJxAwWPjRuL1XYp/qQtU3eRhRbyVGr4p1Z/Aw3cJ1aPsrYJ
ocPo4HaQofbmAhG9xeD1fDT8raxHF4PbtM9OerIb/3puDtL4w21W6HCO/vfVtgJK
6aKWfjjC/aZNft3w/HwvEBXvZSwyulXRFA7XinKAx+Ch3Em2o1hga5E8xqCdp+Fz
oqHf9lzScKmj27wy5Bz92e1OZxabKudc8NfuSOSOGqsK+o9jebP6z9R5W0dFcRG2
abbrT5RtGQw0nE3PJ8bXXNZ75NLRtorHVpC7MLlslkxo77+eFmLRhG/2N4bHN+SK
sd3CqobDge0dJtMvqPBEBXIeKbX90ySCXtj2mEly40SK2LPq/R85RNV4qyIBe1Ux
+tZ3Yb6KnKSFE1vYT8p8H3MZernsB5CiT67UQNRDMa4eQEaLm22f3bHY4B1JJaMN
HcISuw8xkxR/lB/swaC7vMmqCV68h0jxjp2t3nFysPDItkKr5ZIxeYavOCiy0Fua
K9K30nSeYt5vW+uhRpxQZ5FrtSjN4AsqFBWJ5R0qA5bTHrLEmBdYfiGalNyhZsSp
5vUM6FTGjlHT/bslzKh5vS4f9M+NCrb/rt7WPdoV+joQDHvaiZ6Z5pubMGcmlLIL
5NxCh/w6gHkFcVXmI1jFX0mbavjRKNMA8qys2kdWY7Bn5icw5QIZ/JC0Y268VVnS
SMURSPLuhCRpZf2sNQXrrDRsnukTttBFUk5A0GzTgZ6hCNtqyRuq23v6PjJdPS8J
gyyM+wpqiApGlYNMpt3F1qzvvZEBdzkTNpQlUN5pP5Wa+lF4/hkZvby/XvE3+TRG
6gSZaNh+AN8bVo6nsCDobxwsZM60/b5aGhaH5iMqx65AISlC1URj2I4/r3yPq2NK
zCD4djeSgcKMJ/s1BpvcVMSsBLg7K7aJbYqsTWY78DV4wEiAfAT+vFhgd4nAplQF
gVJe70QQIw0QXHROoNxIm5EFm7OGo84/0alBGXWD81CkUEZssVuSVC5l6mnNQp5y
uRW93uQtnCl98AulkAYAegj63P/hzJsl8Ha9Im1vKq1Q9/R73YABnhhj8eRzxAjx
+JjRAK0ddBkXaCKRMa+tgtb9CEIqQEfyLJnBuRhrOER/D0gu8VqUsTZjShzqGMkR
3tBM9qJ8Vg8oMJOqFDATMElE4s2i97Arzv2VDrrrvHipITAqZuoB6B4reREUfzC4
3iO29GBvjaqjTOIqs8Sfd55fF2iTrgA4uNvFz1axKRNR8xUvBzhTSClOatG5diCl
rv1+mP6J1o5Fp7aDvQW6FpWpBNHe/XE0Nd9fKJlrhYTBuFtF6RPKCdxMRi9exBfL
dAUU52vGxqFlVWQGRrAHNJVe0yItIpW27M6DVi5wHLxMU1mKYeGKkK/Ea9CzB+PB
/v/iUnfFNm++RgxeQGL51Q01WvPo8Sv+yutBWIl24j6WBT2hC2OrMAw83Ov7Ej7v
yhA6qmFv6c0AsaB1iL/mmf4t3T6ZwtReECEc9K7M7F1JdnhPXi/yanA2sW/G33GP
Kb6ROUt4JhAuEEsNjDg/IxHIsEy/0SeZ1JHdCSnMxfB00AelNPiP5B1b10Azjy/x
71b3gm025hiRZwRjhepjx8tQV7PX1c4QrK5bwc9IrDhDHJHsJAhNvxshQy4etVl1
jAPLlslxSJ2Sn9Iyfpt/DoP8WYBojKzTbunONqziFsMPuKlNuAbhM0/YYCEUEaHI
u4drjPpyQCvrN7ssWr8cO62IJBiPBnk9g0yofzWyGNJHkOrCK8ZcXykk/eNTV5sQ
/ky5CRTR3/nTrdEVNSnT9sB2tzaDbR+/RaIm83KqYdV8F3pdPGgR3O8bwPMALB1z
GDGa9RWaQo5qcn2QLH5Pu01D0f0QysXKjDL3khzf22tzEtAJ5bj6DwofscAM2Eh7
6IcloobEiLoRkWqeicRFiBckTbHntfZ6fR7EjVUaR1085k13sqrW8jdBa0goQCjL
PC6lSUKrDHBKLI9Qd+Shnkx8xXA9aWBRt++kGuDLYJW08InGzmTbs25I2PxYzc5y
Iz159QHTT5HOVP8sKDfTVo+yLHbFMO/TEjBEFh38MJXGq2lJjhM0k6KaHGhuZm5F
AJLCbsNPS7rSNeIa/VJBab+7yABueuYfPxMBb9KFwuEUKEChVu8foV7qSz4L8s6g
3aA1V8bm769oMnZ0Ep9dYGydBdNhcOQD5fADPdfEx1q+M8QAYeQRMzQAuFTtdX2w
iYnvnVf0DLCOQuj4rkUtjCqoIXAHCT0XLnlJl7jwaEHY8Yv6MgsvGv222Lx38LtF
GKZgC2YprggG00j5XuJOlIBXFkIEXwrICEaM1rCAyhALmuHaQZmodsTi5pP0dPo7
aTe/PmJaN04OOSXpOjDcXYE+uSCB6GOLQkW0uyQFrfykltczP17iILmqAh1DNvl7
iQJ0CSIvCQRgIMjyucGEHJv71eie+hj3I4dUGPofr0G02i+EFqE/+SQHs+ss6Kfr
yQRpLCOHZhbh49YIqlnThMvZVqeN7u5r/FKahDEIsErIwIgH3bUGaHkiQdM+8JCL
uuS4+6P98Z8RdcRfoiGT7lbw4beHuNOU9NIVg+20QahbtfnLB2wh7kmdbdTP55tx
vVCk6NN5Hvpxc7c7PdegsKKkN3IVOKZdPQnnPVx6UNg8a8H2Lg/zhZf+EHGiLUPd
ABrNrVgQoYOaV1Qj6HR++cnmm5x/QBmX5Kn7SpaMJSOunnW8afmuglS+4dPzIUbH
AXS6cG0Siu4/fcaypFI8el+dGDjPV67mnkFR0i/Q4ZRY5RGTl10QCIYD8rd5Srlz
yjnHtf3GtMbCLwS0ZpwwkoL6SYmGTKKNYkwJ1CPv6EHbZ6pND153B7mH2ryok2Yu
i0TlnhKZqBi6fnf1DtkeVRs5Imw08EIrixG5mLbmIzndDIjmSfib/O8C9Mw9aqWn
QKNti9x+Gdc1v488W7O80jhsGTUqTY9KOvIQdHFsG/LJOxIiI2BRZIaWlwOBom3k
P8xW289cWofo4vSu+MMCTqLf7UPD11WxVahLQBuoAtBCWZK29XO8glrHDc7ph39d
rgUi1vCjNb4sXP1u9so2WZBOx+qprxipj4MzcQqIYgqb3PIMDn70ozmW5ZuuumGo
Bf4uoVSvO/hIBaol5fpQS1YpfV5NkcZ4NCyRSxawYks5gOKtmc6bANfDpRL6+KSh
lWKWFZ2gyaba+aI5frKP2WYDLb7EBMtK0biNUX4C+ws+23TCJ12U2cXNJZiEa0O8
UJp0SfI41gYI1zjMB/3vQ4HuhLEvJGkYIwmWx3GEvotwyj1KgynLxzsTjbri9GzZ
fh4Vbp1K3yRN0UexkCzcQRCJ34JmnYG/GbNxWt2tJgAskOxa4j0skN69qEw5bCXU
OeBYrg6oxs5M7icSJvW3jsWfdgsMcikLV4DnR69VlEY/A2+Hl7ttERWd0P/gEs7Q
6x0GMKTR6+TQKu3+F8Ja0G4F/H6AUcdJhUAk/K9gBNFGyMi2M/B8vXQCgzufgI4F
zg6yZHegE2p+HpbrFuZreuN7anYVBi6hyLyDi2jKEVXuDcV5QFaIAaaCm0H3Ydm3
eq54OwTCrFbx291z91+uw/+99urBTEAFLHjBzbDa6mWQ/z0pzOw7EkcWKhysi6Yd
Ns++3/E7TZz7OaVZBUpsWgF47Te8/H+GQGoyWx2gioI2KlXY1fieW+c0fA2Y1Dqs
rodZYxKVKLvGN1La7G2LoIgOi7UfiFCAtk498S+ZpfAkYT6QyVMGd1dKTrH4Rjus
0fe/m9G8g+LiX8I0/d/IZ3lZVzEDUpRCc8Zxz1xSUySNwhuZfYPtfjxVpT7ndIro
qxcP98naVWz3Hr+LjKVSHgeYAzjJfXTST9kdQIiWfoJQSryjSwuJc1yeArm7mv38
9BDufgmnNtjT8JyW69SS55luwKbzDMHs35anjdfDKErLOp7Qy998hiTJExfoYNW+
5nbAT+1KBloUlgCJUZZVapvQVMPf4sy48DlSP55wTVTXLa5VKjra30XMKeXd36A+
34+agGa0NCFnpS8xzubwJ9oTzaMk1o6JRlIJPx8pz7GsHlu+NuD6Blwc+Neq9VoK
SMcWMLGKazEaxb8JhwOdn4WB659Uk2BBMrn9j3Eu0LeHK5Wjbc3XrIbSF7fdxuTk
6p3NYKexolH5TzcZoQ/WSCd85Tg7XjRCyM5A0n1oPGaSgSEtEdk3TxtFxgimbWYM
C42BT8Oj9ppcJpiPtHz+AbpODpSWzvgPoABB6+/kuAY2vrcbq/7ocTBt72HK7rTg
TtNHODYnadMODWMFuS5QNvltuE/OjLuNdqcg/NH8Mts1LcDAvLCmfp3r5ZpANtW5
lXIe2kB3wgArpjioOzag2aDy1tC63EVH8dbLgYhoX+gB95qP9EAzftuj8xp6jVED
7ZdR2153bW9PrBBGiU2S1KKIQi9p8byhUuvrO6dQaww=
`pragma protect end_protected
