`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
ilovciy3WhisHf5j/GAJxk9LmJn5Zg5MmvF9X2hnTWNS0SynsgGUb+X+We4/tHrV
Svx8EsB383L6fD5hROBORnLjB6dhcqV7q5D9O/O77NmzFG0obj2Y5wPiQfm2VPpC
fDDYLaxHfK3CDQ+M1URI4K30KZINWOSR0QJ3+SQlhL0=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4080), data_block
cN5g83qFj+Q6RmEpeML5nD0YHJQLjDZvh5SjJXy/ImX4yONKK1M0k+WTR2xZr5cQ
cZZzyv8sGpT4U3PK6NirEAK/x+2Vrd6s8YvLyKMaGu6KfTXA1RCyOSmqwa14aUu+
Q6Xd+bafsVCm1Dm5ENrQdXnTl6RdsXnGBWI0LBEwDn/D8OIGAwKiLiiWPa2uQ7Al
6lHn4iFcYo96+nOU/LtbXE1Lqxa4XrXdCp8IOqy/Y4yPcAcBdBWxZ1OPzJ5HBwyq
0H6LmM4Ue+4o76Qbw07NSYdFMONcUWIw2dSvo75SThq7uUhWfWetc2NTw0c59YKv
j4V1VMZjCNI8JS3zFrMgPUi8Y1q35aLnYSlpUbid/pN4telkplRb31L0MlmZXRiG
1drHHmoYANgcDRSxI/JiYD45/glxm5yj8yYidrzoGEN04mG/YSDBp9aIwpUWHsJg
Dm7OqIoh9bwMyqdKZk7BjO1tdBLycI4dxDdl2cfiYdWo/O0zKfSYCEVQo64M1XSh
gjC7A7vhcMzTDs7Bu9h/3GEufOtmliU3RI0Hopw4bFiLZbM40rkxWNjCfz8MKtnc
MIdrh4R3pc5346V6o5pS3E1aXZdWZA94YT0NUYjrcC7yf4nJj8rr/xj89WgbtykS
0a2Quy/G4q3J4JnvdcWsUorCYP2BOFmvzsJ9wRMh9Yb3LuCi6RSIEjMnBQ56BJze
qrJv6lMHBdeV5L6tcrTjLzPQYjVnXKeZvXy6MR97HRXi4darpALTQ5TDZmeCXcEM
QWNUNM9SCUSbA+nVnfmcm9T8bc6DvL7Zf8J6mL+p9Mv08BEAWGaS+wyYBKPBh/0p
TDcw331JgWQ1aKcCb9U04vY23NoRDiOZa+9KwU/vkrgC+LMACvzAun9Ad7ip2bsd
rDmfehwrThT1RkNiDKdaKtET0EJ9Tkev22bU57b3Zh8fzdKS9Oo6pczIGvJfKC/W
JRlcySlghFrJWP1UJfh7C0UyPbHYeiOxHd5Zn63ErXWYpMy2WBFpYYElcs2bbGYj
S/tg5WP+HebVQZZXhNerccpWqYPvS3hezJ7agPCnfib+XXHXcoeDTI3T1Ia34zlN
9pHBXrD/4ZBtHM3JRLiIGLKwcusJ/OK60FDULuXDPBs29hfVK/dHWMCqnyFRrrJS
kUsNwZLj+ip8//7JdvALBEUJR97BjTvFZSPKUEH6wEhtE0Y7wF71gOq33MMQv0Q8
um4ClsKAO4h+6n5/HrDWdrPcNBAJDxjrL1TF66fXkUd+s4VKbV0cZclVM0oOwpgV
83LOIWcPeBIt63obVFdle8Y4URhAX4jFoPdHzDnXwmJIvCuPQvblRLMzoBMExqUi
+2FqtmbsSAZcLxBHmoXjNUPJVdIGpXPtTKnY4rCZxY7LUCOnaHdcUgbE5mNDaIG1
mLb+JY2R2nagaWMXLDtmD/nsS1+M9ZWhiZJgvoPDQgJcONahYpa1W7UJYFuBP97U
heWaDbAo1OHkHWC5WH/KcEhJ7TOqibdmAI5riN3lMkM9zj/PR4SkQyyX/MhCGRAp
tYMWlB5lb9h+jooWj2UkWQwry5v8r8X1y2QYoOUsJn4G2Rz8Mhr0MuVADoWPndu7
wsQ4AXRLq617nXTTWkcc+6V61eUv9VFHQc2GofIBYH3isvha3e+QQ6d/g5aJR5v1
j50U1ylmMWCQAWungFusXmShTWIOXu9YBv78nUTzOkKsscg4kYu0w4Tp5+KrSd05
0M99pPI0qd5OrvPGfn/iqbfXZN7+potdC9Obg68oNDsHhkVJJKK6PQaxZZ9/w6FI
aSnnDukzYf/hUbj4LrqqgYh2dZmtM7T28l5QDKSNXD2gxhc8nLymqI3uji+FRpyi
UiXr7a7nwEgZ9LT9DfBhZNAyBYhaltgojPXb5Tmd6EyyikUFelR1wz6A3/hdXY8J
Q4TwXnBiKrs91E4GoCugRpIN4laU+qf0EvutdxaSJkK+t1mQeuPD3+HcWK3IonBt
H6hFPXNtkr+hjRVVUYK28rxvC3iFsgbDtKG+p7Xy81bjv1FHkTpBRk8ShbO6QvWQ
tCaD22oMfR2cZrIBDxuTFkQVxpTKMi4VkPd+6D/LEddHN5FMtp1qRZvBKzCqGn5y
bV/6sFaTS/L4ygNet9yaH2aUJdP2d6bUTsjG+TyAmdGf937Yw49wtsxiPPObiZge
s+MCs3znoC1jWLSrLoFlCNUeJANJMrwkGwr8QShHuInq/x05KswaPpXnaQ9LFyII
X37tfem4PRgJdwCbQnld+SGWPbeC92t0hynPIoMgFDyi7XQa+IbM2kVVgfXUb/us
YMR5ItNbo/V/PQw0q6LPOL8wBAr1VKisYUP1ZWI9C9KMILnkm4ckGcXcDIINVEny
9z8CYTScxnjltO/PhHEDszGM35rHMvk3OwIsGusKGqFw6g2sU4PoDazR/cpwGbaj
jcS5bFqCyQw2eAfaLZhlQd5zUD9oACbmNYjRsYLSLcghOA8XWU3uxobFvelKrym3
Q4RzAyAUBXpZQ6z41qqn+xcfcmtGx/ZOOLcpM1qt8qDe3g64yL0LNuRj8TIytZAi
6Wh733Q1GQYWg3pUeTJFcE2T4BLyk4LEFzaaBQM6x3HemtvTk7Fb+JttM3q6NwOO
X+9Wgmx14HcXm1zI7kA3SA2bpNk57TzpAGjtmR7jv8lT6L2I8qs9/7gV+pzKO7Sf
cfQ0gJZbCCq4JGFa6b+RWDb5kLez0/kGzq+E5n8XInW6qylmp2+Xl3Y8+psWWpuk
LZ9FmPvNAGI/YxxrI21JdWwmc1SiXFGf40jU6+CQwJWHoBhYncoK+5rYqdb/G/M8
ePe5KUoSrfGV/K0AyG2E1TQwAnA1U3nDpPUJU8Nizv/+S9oton5kfpuibGjh1O29
4Ob0rRjq8tOnpxyQZQyXNw/HWhmJPe1bqaf2jMaxUq4hv7TNrsjKGhYIkUrykQ33
Pbd/g8x5UBmWZwCRIgEhKdjce8w8Ko2DArv3DoBvYMpDFmZbHWrhQNod9lB/FBY4
ofQ6aqlfD+ji8wZeSgU0zywPL8Whh5+Lwm0nru2itwBU9cX+Bry0BYI4SLlGhILS
c8QVPEn7weIiT6bNDR+Z4ueVY1oAqrai6tMNJQN+RBeiSYa6QqyLw96TWlYtcoqK
FWahbXATc5dIN1jrAfn/Ht94iOlQr26RO2WT6M3VkpBN0zkgRAVIrcBgyJJQwe4a
B08IVasNcr2vwxKGjo5zv2usH5v9stRJYyfbS/qatrJhwIFnwcYhldNCjPoc15ia
hglihJhWl5RTCA1KqdzpcmBot/XGDf/ZrwkjemkU/wpJWoWgTCtZPKT4QxXEsCfK
HUrkPzApBuLOLk34QjUHnbs1tcGhLw/A33UNUC6+INu6yb1Jl/FNprQWiz/RSJbF
oZwtDcV0dxPeTw4NfSK0fXBmUJOWlb+xIN5I/UijKeMxMQNPf9pv7ouWQoBCOx57
+aSqcfuoD6fyJ4sQKQ7TQl/caDwYNhw67laO7MXZqUVGDBh7Ilp09V0FQ2oCs/HN
XMK0c1tMnIEyGNwpkDwpQQZEcH0q50eb4y7fg+4EAhc2pC66ZSxrWsn9t8nclxwt
yK8NNCz9hDe3GE8q1z68giRcQgyWAgcGu7e3F+ChdfXVlEBdlRBX0jVenlO6ZN9l
VGnTUsHLQ4mC3Y9NzOi1xbcKHm1Er1FeOzgLeyyU9o9NVOv7j8S6A04v9fnZL7YG
7yv3m7FKBCKXgTLUeyzEbqV+EsiGz1CO31t+Du3W2EHFEwz+UG4bl4jMeF8h6u6F
DodSe7mmlr3ot+qQZvu6oH2i4OFdjjVoPsU487pdv9uDywbeURKWSFxZSyX5xv0t
d5iMz1KWH6OCiKM8BABpAPodqC8tMqufbVKCnihbr6HYGxbEO7NQW7UBoAV7IEFk
orrd7ITkoVZJfkGErsFxOm72EGJinygYHdvDBwh1rmDjCEyKwHkUAELHurEhtc/l
bDpMwl2d8LzlL3bJ9j7RKijIZow5IDBsAWbDR4KVTbOg8qBC/kUsX1Pa2D+JDFOA
hFfolKxZ1+vVQloqjeCHVzBC54EDHIAucVrNb1HFmsdlEPII5niYM0UMQXxooyN6
+Y54aaCciZNaEXaCoBfPI72UiMhNCeyJLF7l7bvW+SnN3Jf7P+195SHOtzU+Q2rY
sYxH20DfNBvB5z9d7bv/LAS+ruX0Nvcu0GqYgH+zmdfN0tPd6PmYAFkoeP+gV2pS
tKXZbfpubtUj33ZQDNWxQBFc1ZO5JlphXACoU/Xjr5Ym2s0IzSfmjaRoySRIOU9n
ohLwBNg+0IoRGane1ZbWKJTJi5IxLrxEK0r4fXe0uszlw76Ow6Zz8mKBqdTWROuc
wp5o+iOiglMeBglENKt/bPiaDcA4ygpiGpITjqjRG2sws6fyb1UQXvozeDgzktgk
IUernOvyGXuPH1GGMCucz0+A7P4MV2L+TCwxLB++9pxDYC2K0Q7cvWjQNpiTmgqk
SU4wVFyJSKUnZAfobWviRLOLGZZvT8dW4382pcI5aXK50T8Dvd6ZUx5vLVstfEGk
2KUSgvE7Kin0fOe3kb1SyvhCRGFFQ+IUX4S6sna+taPV+JgbaEEwyaCHd8qfFUew
o4mwmh2q1blzb20z7DWB6u8xAMlU74I+MCLmoytFVGMreBflCVqCJZ7/3yZKDT4y
JWAZWjBM41U/tPWFqrLzpZXuBzfRivecNTaxJdFAwrovSHsr4z0pCYPE9gRLcbdl
kGqavFFEdgEusFVPpo6EQ1craJHeNi7uSX5fDWbQvWklCUT0MgE8A1Ag+/FgeDmu
tB1PHXrrTYf67o1MHdhLAjlnSqQyQbKOoggUOJ/vg9A/dF8EG8s6w1Qxuf3KuBGo
3YnCSyM3+uN1hhYQBCvcV8rWYBWWIzoyDTs4Z63sCjohNp8cZxVdLbtpo35ovaO2
KWCNSpde8ltFpV0s+oaeVIeKxGxEnca6lBp0epTO626VG6/GHAYi1Ckx8Fb0wHOX
9yJuWINKwRunqBG7mHNa/s4l93rcCN2HDF1LR7A5EU9H4HbQQ46fT4Jht6EsX7X9
+jqiYI7IKzDefB834Te1ULSFekKEs0NKiGhXiDqnbm+8riMolvprApwkT0MjY0Fb
FH9kUE3QhyMwiyvsYICqfCDQyqwbVVrimPTZ+QK1HGzkG3hY821tREQ7ko/bCuwJ
1Sm07seedayVwTI+LxUJMS/Nu/DUbl/L4/THZjqtGacxpzovyx6DIrnar+UlCZ3Z
TB47pDIuP5Daju9N2LKj6luWJjPiXXRJEuEYggic0q4YK3UU2Wwxanp3SSnyj+bi
EYhIDF1iAeXyH6NTrhE7wAz2Ek53HHXTIZuOkx1NS4g/FtFtj03lOSmYun/c09ON
55rqhKWuZU09bYkz2qV5fdHbwNLo8T1V+ZVrrTYS13rdbpGs7njvPjv8xPZ15ezm
`pragma protect end_protected
