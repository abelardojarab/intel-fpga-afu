`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YZi05o3tPGSQ3b5ObijRHiKsX+MPoBXAbom9oa/HhGuCdMlYdVqawenGdwJJPmo4
fRBSN+cZKGl6wh63l6kuA6Fp95kwng09lGsoTY8sPM/CWrCzzmMAahZH9idy3r8U
qZeCAqsjyvaTMAmqBepmJTYLjJlPZ/UQp/ciIBq383I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34480)
APrFetBcZ/zZcvPvV29lJ6f+uYFP6xIhPkim2UbJawgsk25uvjH8tWdIZON/Gxna
bVTk9SHm1ZtvQ7/k3RL41d/2DjFbHslrlOe/7zru1PHSyt07aJ2plRNdTv116zgp
ULeVatEOrsnjeP5ozNPMxYnZAuzb/sHtjX9UECl0b+wTkDR9xiih/zjGkf0YJjCk
QqSiSP/+JEKQsnvu8Ir6YLOwtnk4of5oKQgPDoWjy2cwwIeTyr4U5hgMuuoIUn5a
noacyCSkZNZspjEBowW4jBGlBNlh1Hym/Rrxbg15sHYiaeQI5NYZilKThTJ0/jbL
vk9xgO3CyHF49Hx/PPizzpidw4RxbW7yDhyA9usB/Lbun6ov6p0Z25f+VN7izZ0s
77F+tuZeF7h4UnBmA1IjCyOGgeKIttwh3ECTUue3F/E+IWr0IYNWZkHHdQcrITnY
TN5uDDtKEhAUhL8uX/DXiS7kohhWXJM36r7CEl3VVdMJ0ktD0kYitKwnbeEQydWA
qrwUXskcvOcPva7uBD7i7+Y6oun1VqtRRWUCj7mE+oG5zNzCsVHUebukgKkvVw25
OInRujXGXRY/qaSccFewvPKzrIncAgfzyog8tCHMWfObINDss9y/PbUMN+AkYD00
iHRkgNpgdeT4a4y6+zt6g2QoyM4/9+18slJQcbIRaOX1H1bQAREYt/hQHAqdMA1D
tU06lnCviMDYt+Kl6a7ZywuzQloJrUvQSUJMkrsxWllHgzF6R0QKs0bKXiXF6yTK
vO2g9DXz9BYbIIAu68KO/MJWfQnLKuSVLSCxGnipwpfmhZPXWKzZgpKpkERD4fNW
8zEwh9+FyDeRkYRpzx+fssGy2u42RakO0of0yhxfcPqNB4Ajevvvye38ERMH8Qqw
cknx29bd9Ndawox74AF161Yh6tw058W5sSCT0MLChx3sy/mxyn733b7mcZfoj5Ia
HM39RiW/0JGNcvDbxzt2twvqbqcQ8StwUwqFQdpCJt+TaFcsa1gicmydetYyWWdl
wUDSWd1WM4ERJDLsVuQQHtigh+8KPQ0mfqYLfcjS/jAbXtqkAAhqC6CtXHLXeITz
ecg4c3n30RZ3nBTBJGiUoaqI0+Gxk1oqP50Rf3RnZHlR8/U6WEIWjJwSFDCpEWdY
liv3Pm1ihHDMrTZMLrz1ic4ftsVBAfMW+5aAMFDr62rMF//nD0AVCULV2unzUBwB
thDAwuJu45HnVC9cu0ZpNY1ZnAlHGYUfORIVF5xSjUB5yQQ6ypi1o5W5XqWNdL2T
2Rp2WEGbDEdHmObXwXcC2IK0O2s2ltrjzOyQahbG4is8yvZllclzoiQkrO4rS1JH
NXvoIYHuFi/Hvxo04aWWfewIRVaU6KzddndXuC4cNTmoVA1dQanwIyvplOk9Uu5+
fbHG24LCgzyDxqVQ2WSOYg7BiL+k11vGTQ7GSK2Yww57//aa2QcBPBzjRR0mVcHA
CNWBFZkWA4Rdx072VfGoZK03zzIO0fcX2SDUTfeK6j1J7RKBtFsUR5EWGkhJ10M+
VwX5Xhw6P5kmSgjuVU+SRxgeRzfnhonC5NrIVhTjf8HG+la1fA+bpCDu5f1AfjbF
VfKzaicQ/Oknom8A0dP3KV32s7qcXGVcekJ0tn91AoWVhz8OuUMENTGViCFcKHiF
Q7ebSjUHhLvmfx1UghxP+yW/9ShZuzvtJAdolmqVRR9ZF9MArernBCnaHHbFwQZT
3zu1jLD5musv0G2eouQ98Q23rHxuDcIeKmB7ncWkJjJRq5HpOBf0q8wX4XLJ0wGl
ZGa5ovZpPBSM5nxoJY9VVdFzKrZsQg5F+UHbKHYQdyGppnVaJM29R//YlpKWiBpx
M4nm3r0zCr2+n4ITBTX0MkxslWXDOX+mKUYhsIAAd8sfrGtZsNZ3GOmRNsl1GhAA
yWNAO3qOmIU8MfVdk4LbJl81e54njVBdAaWnZbH6pO7oNxpH7NuX+2gIMdmuMx9G
vS8/cJeRqvdelSKLRe6Pe+u8B1POp0jVaQIHKtTW8H6rJSSbFO3YP7t8e+wkHr4L
GXMTG+jvrNJ3alvh1oO5OZQqJ8x6D9Nj5kOAYMeUfu4WBU2xaD84P/MEeMII7BKB
tqtRghar1HmiJprLO3ooHpkadJWpD/tUu1ATJt5Lzln4nfkFtqpkeFN7y+z9IaPt
rdi6T5089c3XXVgyAOzGZRteTNIeOoodib6g7JtY1TEwLSSLkCQoikij9wY8Viez
T9cpu4iD8iLIROX94LAWvQpDNQCmoGj/iPV/WLQcsO9nI1mXZtKfPYB9sFOiM04D
gcFWHFy+uL58EfEJvUq7q8znqCpB4PeRxa1rdXqiPYNJ0XnMQrbMP8Fp9TGpLsdG
iSotfdhc42caz1liU5i61gqLlxoZ8EGMEbAEOaEU1UUJu4u+3mscZoSj7/y88WpY
ejKgj5Ey24EK5r4kkxCiTodFw4eF+UNEuH+8+CcbTXpUSzfqNk/gEL472Zhms6gV
tO/cXQ3jeNsdnoKHN82TFz6gr46qb6ErTy9ulXXfqQkYvKwLR9ORkGPjo2wKvo8y
SeqnwOeIi235UzGoilHmmnoX/yexXD+QMjoish+e8WAH/V00Vvj9JmiYKeeTr6t7
x2GZGBMGc97NW5O4EVnFLJYcJMhdcumUALn0gMCnM5zutRo/ovwIvP3UWKcVHEZ/
btnklJeSiQFm320gB6NvCBfTpNf6ahrAP9RA9xQfm5osZYrC44TCF2jqOXZD8+Zn
/Ed74xyMPhJHNjmuig5z51fC/iIz+HgfJrNMLTeBNlErCzq+BeIgOkkfHvbMEKsg
SHiJll/C7tkaoe9q9pt55VF/ammgxMjsQaS/7UFNqubUuFUu5SrTN7Lulo3TlexA
Ah3ZB+2QELhx1LilkCefQ4dbj0h710iWANgJLmC3aJ3z4SJzT69fkNsat9kNUu0l
vCFRvlcZGHu36fSZOobb59VtFyKpoGed6LzyHhn7RkvlLSXP4K+CjvrVfyaBoCgd
VzbKLVseLQsZX+Lqqer2dBtfgFX70CPNhhmMDHlJnQ1Bj5P0MztEtwVvdylRERXJ
Mi9PfVbaNHwwS17I8MK9Uxi9w4Xbhaj2u5R176HhWaJl4J7pAssqyabGUMvROWws
EWMmP84H7i92CLqeiKNRzVOoO71RY3EssEs+IC7u0jVpYaU8DlSnPlKKQLQt+7Ly
6SZbJj+uHi8LgG8kQOroW/LazJ7MOsbonMyV5mdU34/NBkmzcisValDGJsLiwFBt
qIvHdtg34kTOR+6GuLHhagdv7LtugkZvR9FhBrz0Rp3AbB164AAUKQhOeFNc7lgL
rdXc7LfRoOR6NJauU7NehKoWRVn/lM5oPrZ5NxHO+m7jaT4NTLPbK3QKX8bn+VnP
P5pXVI2HcQssuob7/dG8jkhn+qi9xG75VA5a5/0rEqtjnRoHlfVN+R6y0g2j9pLz
KFMlBvUHOhOidGtLrqY5HykJ0o6sjIJ8h04dXe/EaDPZVDuI1vcOvl9uRpm43vx+
I/QmhkDHutaW6l622kTVImP5L2FIQ/pLLfZsQ/6q/qEPqp3OsD3PCBX/vf+1f7d0
SVvxB1TGFn84Rx/F1wnZqaK/nNfVVZw69W7UkJ1WYjJTYKmr0dDaBWkmJOURZ+FB
gRxqvfdPWP99scH8zfFny4xGXGYyvQrQqwqwc5pRLVB3K8zxDP0TLAmWb1Q40aXq
WJ3Aui4D4YS2ZTpiFRCJryixJxriNpyO12khFyvRmqJLNCsITSHfLpvnEVt2kRh2
b6CvZGnHDwH/wWTPnQhHv+u8IZQ/pliFDelqVRL75/63LeLR+XBROJTkVjkoqSSD
7dloh+hEL1hUgEErTJxIDloBvAobvBUubj2GzNc4vf+UVT9t6hm0Lfhzt2OsFQb4
ag3o49C1crUpbvFMh5bjKkn0ikfvJ2a2xIsbR9BGTwuHYeSZTozdGtusQjoe/HoQ
n4ru14tL2UF5OwSnW18343ENgjppT2kzb7OKCBSggNs6s7G7b5/L68dWOgLJIIEe
lvhUhhzyZ8FTNcHoyBHtpG9UlQe+GMwPQPnDs4MEG+enBaakcC8OPX2Z9VveFD0o
zxBrk4G6ZRUfV9XXZPn1s3zw0+2hMSKyRba6CkScpSOG6YD+mfZq/LdQ/POTS0i4
fjovdqq48Y2GSauEodGRtnJc3I2qMXb9Z9+8nU6HQJ9zw7U2X6bBn7I3GgY8MjSx
XkMrCkI8MceVx6Ioc1r2iLsdau9SzHlZL0cp5aAN3b6yaJg/XylWiqw8TsHZDAGf
84SxQmzEwE0IrqsGURrzR62ELCNy797fhnNj2i4EYeyO43i0CT99wVt5hUZJktQf
ziOFYKWxZkxjfsVnLOT1uzxHMk85f+ll5fS/10Kl4AxDhKdBtDfpTHbbLcbPvFCW
LpiOVwDFmNEXksrOk6gUXedhgSrn+5lEn+R94F3d1uEr2wdqSadyTwgI6n8b9aMd
3uqheu3ZDTgG1D39lPHjiEFcdhRBEpoN1hyJxnn2HycvqVNUkCtNqJjeU81l82QF
SaGsf/AzKv3StwSl54O74g1jeaPUpDb8k+hyRhsSPIFMvc6G62kFmrM9DZKb3+7H
uQAwdTZXLRrB6NNiKGbkrl0gpPLgSZHCEqzeAgzFaOQ2MqzO2updXSuvwwLCJNyf
/ZaUWhzgf1Gnc3Vk8IBZrsAtqhGEV2BkFOpoHZRLGh0JGz05U1wl6QPIqPrTeXtK
SETdQ9ez1kKNozmCuEfhc1HMZ94Mex+7rgmyJl84OwAeCATXRql338XYkJ4xHN7e
NGiiyzs0hT4Vb4BhScJBj3+iNf9b4JprHAyhTM+b/03rvgIptEcFymuw0Poh83Lp
xyCTanivrN7c41yZi5SfXkWhrcy7lbXhT6S69HGbhefywMrsxS9/VFc6jhnWaLCI
w5M9yHwqAVtV9BdZ0xUcVgiWnqbmB4tCUvmeu+ZTcbmtyJfS7t3xrs7daS3zTe2j
Wzj6yS+xvljcDZ5IlA4aQs001werO7IX0zHZomuykMeKEpKpCtasViSPc8ENrk9q
e0W9CqHW4A0rFe7iJTQHZdb3JX81nX/9QeuD1WbA1ozz/KLLLLCbOi+KKDxljJr6
VU3rD3oQpJi4wSmpkmZ8Z7o4rwXBiRTsOZC/ja/d6tuycfYOo3caVtBle+0HCYq6
PWKFhWeUssAH9cvZZzyxwljL4WciSLw1GxkUmbq5uPCkCP5xBydAX2uxr5Hb5h9H
BRTf7/dKvewY/4sC7wGWqWvRc9mOzEhX+wx/gdQUEDDYJeXuggMYWFUT+/zpCQt+
uxSwjsZrLpIAH9kbZuIHqIXYBIyGTK4R/xxRQo6xX8t8wrqGts7Nszch4xm1tXZB
HAG2U4MrcW0/ZQnktSX5fR5koAtuV1T/4EFYBYd3gdJgtemXilgixT3oDZVWKLnj
OUzuOoMB5WTyjo0JoYCzSXQ+qKss1NcHntz+S8Zhezvr1AxTq0e2dWzjTcBKQw0y
aNfsg/BEv+PNan0IfmlwmMO2pUX0Tgecw9gIJjLzwO9x3CjQk2vWKUSJFNSKkRLb
S9NbJY86blwDgduv+xEAxTargxE+eIraJ0UUs3EdNp6BnjOm9WXkzzoYqtm5A4Im
37X77Sw0M8fa4y2617lrgXp9/iQDCyId9caE/z+EMNuDWa0bh11zQMs9yvNpOn4z
oidWeKu/eAOudNHNSctkRtoPPuyzM615t5t2O2YIRwVuequvCgwceggsr6M3LxFo
L2keMXhhkgbLdc8Pnq7BBGhp7WdCi1My5SXAfwyURcVkWcKDV1qSI1JmOnvpQymE
TXLPeh1LG2mTIpVgDbt/Nud/le11A3agbKpdtiXL2P7Vg2lkHUaExnvIlMsOVHbF
Q6jXvn2BZxbnVXVcRY8LaqdC8XTUt/UZtHhio5OfL/d9UMCokG4X/1sfpmbX+qth
r1AZLJCLtCadeP305XktrGtTK8gPT0R9C0ZQZu78UgZzloouLnwVp/1S2Ba2lmfT
oYcM+uBpQeObhnbV6d2MwGlloXY3lUCiC7ZayQTwtAI7dXaM39v7dKOcwb3/Hm6R
BKj3E7WkD7maUHFQHUqmGszZsd5eFMtYZyHqYHY5gwbhTvq8XEnjjeqW0bmUJnAP
iwnbu6x7LVpESme5DYDPGjNgfkuMgRxe6rCwfDEEIxscfAgPjkxWgsXPI3km6JTq
19Xhf2LNtEQhzUFDSn5Tk5jIn8PiO/37JQWeKA8Ejt/3zeVX0OU7ydX40Q8eouXM
jykmzHVoVuesp5fZr/cNbcQEkDQQm9b63Qh7JQpxLvQVx99iWnDNq/uuwg3QdhXF
MtAXkfwpvfhXyvuYVoMef8Y0XfdDVjB+8Z6bvXN4QNeXfXz/H7pqF1WDczdHCqLC
F6h60bMUHoITY6DQ9JAY34AnCrYNOqq24lWfuOXrnsRTDufI766LoGGEKXaG/5yv
h0Y+M5mqQ1ffB974IZuHFr2pQWHlerDx4EXWOh5vjQhk0hw3dbX3i2UTDmU0gV0+
Z8x9V4eBDr5UdRYOzf2ZCJn0dXtXOA8ifnzefVqteefY630nVGYmm+/0e2j6wwWT
mBe8M2lLUOr9C9weTQuCYiIAtCAwXuWXM2Cb0D2zgAcRIN3zc/Q77O6rppFGtInM
WdzXSai1U/HrNWra75g8wlyo8n6zLhpNpoetxvKTkPgGwFqJpJssdaBZA/fkmwtP
YgblGbVQ3QCNEOfyS25xZdlKBm1HCcG8qEckESA9XfSSfefIIgswwgE7kZlq4ynb
YmxzbBvWvU/A7lJsvU924WY+Irw6nUFR19l9g49Kj3JtXs3oKkMeZSvJgDRlMIRu
960R9m0yQiA2lh+1hr6q5Q6BMsGnnmFSEzpU2tZuYKfQdxNnVx1lnkSpagpDT2k5
14yWEbj2FERRQwDZx9Tq2f712aGDm7aNpE8UdazV10PF6nl5u0EbgUWnqLR8c8wV
XO3FLBK3X1UOO7TXECRHAI77a77OPXU6FH0WKPE94QhkM1Wrw+69jGRdsvOcbIFQ
fWzricvKeRAbwtUkFqH8UCSzAaTxY3ZKf2b0Fh9vdeLmhCs3hbZVHYSwJepkZCSX
YEhJU5w8osnIUiloPzHIZu9WcA3ToLarKFngulVBdPolAymJcW700KkYyqIV0iUS
Q0dHsNPJonWvNeaOUqux3UVPxWqcMe8iAWdND+Kgrxj8gWSr5dkWrtMEJu6pJAZu
6U2S0Y49vdpoARqgZeY1MdNz5Xmfbn6lgcGpw5WUJYGb79HXm01Zryi66DuK8No9
okPP9jsL9t/jZ8d/SshZFxkB7PIiF3r/ZQR3J0q51JEbERZcZhVUCDMDQCpVyG6I
UCCDwIdZiz9ynF4TayD+th9McbCvLCSFkohjwI1G8Da/WBnHmlKauylua4k8X7pL
BQafpPW3tjOmNCsVQ2NdM1v7tuEXxAv46WvhvX0v4sfBFunQ/4a9UCcxUYo+8A43
e1OSUZiA+OwrgZ1wiJQgRjv+mhhSZbKLfNrHNv5JlJT17KrxtAI3ajRmjd7kBm88
RGufpUoW6p1QoU8bK7F58FqUPdR4lObiu9g0BUoHJ3dVGnPVOzDHqPYSjLQEj0ql
J2wI34BghGj6hus9SPwk+JMFkhjmpH4vP/G+FP3co5UScsQHl1n8OUfffSnOt9UI
PqEk+Xphn5iW115E+YH+v/ldBWGJR6LRSqpUNURCp1sipVmlRM1L7Vf026/pwK20
36H8GJdhojEukw5cy2ZLy4McB0NviQt+zCrrEIj8ZLxphX8j3fc2NeMjgca5U8rF
psUvjh0BArwx3vSw/yhALdl1K2fOhJYhStZl7HwrqWdU/D14n2ESZXd8dJacIxPv
mjA7j59plxYGX+RK9j2g1SpmCGx6WPsODxmNSI/38PJmebimIXR+6ktq/TM13L67
A3aGWa+FVEy2ooKUwpcksmLZKTqJXYNWK5kV+O0ctlRup6Rhl0pOSm3rXfpzW4I6
QoiAOvg0ulOZOzrjQGhZVgy/CWdZi0C6Fc0yUyobSNDq4Bq8/261HxCACneZbBCq
l9xSg0TEjsXL7egySmZJ1KI9lqiiFxlXPAKtkMSGPWGPi/Cm4jfHs8tB2XV3AQ8A
U106yz3fXAdSj/erFzoPA+trrqw7Rm4BJMsF19xMm1LC/LUq2EQJqiSQNWyzq7Ad
gK69EZttzS2/QX+/oyVEkM6S8CgwP3zq/tjv71+RXBJtiazkT7faczMI6VmlLqaG
YVKFq0l4rBoBWgaGlJhCglbCNIJw0FJIXMRp3bdfHeHHZoQBzXgDo/YocZE3audt
7np0uAR7vpy5XZBGcBmgNdrtVwOWW+PwS2sNDG7g2TjGgVfHqmMny3fafdoVq6d1
3mb4RfVatBlvkRWrTVik+1Yu+V5V19sbR64QdJlg0iZ1Su4ogg3Di2mit9fG/0wH
R7lr2auYKMfvDpWDku/uVvNZ8uzwkT8qQf3FLNjXy9wojtQAtrtxMmqN90WdMfvq
+T0iDDA5GKAPrzIz+FmQLULCCXAKIIBYlpxetVNrYCASD7gmtbkieUmLNkFnmbN/
LIBI5gXkJHjuRh7TM5UTm1FNc/PapBpY0wngQwiMcqdA4XWMtLlKqXVMkz3aoNnn
ODCRxw28vTOLWDOtFiMpLwg48Augh5YahxOszTfNKu4Gmr50yt5db+NhzKticmng
wkcx6l3thqlW8y0HGfW5f/8/RtQwPV0RpSZY675fIIcc9xC7pFkV8cp9jwtLmIWn
qrOFN3Wo7oykg7hSTfGHqVWunijqLO0BZk7JDRuaxLW23uebRMLjrA0iP+AVJv2Z
VHcm3Y2XYssRUrObni+fsWAsZat9AYPkvb3V8gwfwtiHxGzdr5VFhoZRB83xbvlo
cv4UBape37IHHU168ePTbrJbHaP+6bT+kndF2W+mzGqEZir2Vv6EsKqT1THNZN9W
VI6NN4Y5QQ0DHDfEb7n5RKJJyU6fkbZMwwDFDki0kUtiVpaYdYcFNYX8/e+HsFS2
lHskDkf5fEcIoQs/A2eSK1TwNgp0PeLYheHolXAfGWDeAkHDmrrlbbQSMZsWmzH9
58ifs6cYS320647atWNm01NRHXJTiubK7ordQyPf5aWZATkyOTG3u7XOy02BNhr8
yVvnevwJNVgxsBubi/XVVcNRR3uVL7Qxdc8+WJf0CavN6PPVG38n3WYaZWadKghK
rmfYSGNUcUlcg4p+k/8YJepjeUfHDFprUTqoyZ8NE8aZFOZqA0EPr+iWnejQ509N
/Zr+qvJTkeozxRd5te64xjpP417hWGtLkgU3zs5CdWpDEiDJr6oxrltopmNfiegR
VxCeD/Ib+X6fynmHCTJnZOBNJxbIljL5QjC8R2jvqd07Tk2yz1c7rWG2IbhIFedl
z7Yd28Q0hho+86iZV/IpkGtrJXfC9N1CythPB4MmqQnnSThOfhvfjRZjnJPnfGOS
BoBN/Ynupz6Vy63VTUxtrhVGvCMmOOVMw5KFR+wSfgR2jWnF2XzqK/+M1iLIpIFf
nVW2yp6nI4e5Dh8LGtC2MLLGY7Qp9qPXcydnSYdaMW0Nme8JIYELlbfbwyur6szI
E9OxiwoOWqED26EcMPgacOX372hYJW6dx/Ug/xfk4tFTIZXgHARFY3ksX1Vba9IA
TRlvHH4iqIxxAQ61gauBivYwS31yvoyejgB6OigWS031CB870YSzNLNxMjKkdFe3
b2Ip0R46EW5qaHkyZB+wXMYxUi5IKW2q1Sx4RHBp/u6/wZPma5tprL5qnAdGco9r
y1LekiYJXjs0rWkWzanEPo8BnGma2XDmYSpHxRzO4v0vnlzwiokOFM9HLAj/u6TW
Y8ZO5p4OsIV1ubHvF/OOPSP8F4kb3wNU4nlUuB8L9u7wbTYa+9g4LMC6wgc7I0T9
REj2yjP13sFx/utudvVZ6GFjtDSJXJck4dgPbBzXj8M/FqErIy1wRhTnqQBqG3L4
80zBpHc0cYKiKtoEyrbvqeJKpLEzfrcy+bODVX6tNNMhLEAi+gWwMvvRXMOEo8Y9
MPUpkNrSp63d4aWG7LLDQMUV+5pPy0pJ1GVhV0hltxtQhMXZuI3duGIlgQfv6E9A
cLBN5OoEpdiskDtbcUbQq+4dGi6VW3fW55+/k1cfcR/v/DriC4Tbtj7C6Be3/H89
Lo9RZ9ScupvFrPt2KQfYcvLh58nSlO5l3e8XBDXAwwF71LpMb5N+znDaxpg0RlNt
e7qI4QU/7lvXepvkR5DqpjIXKl17xfVIZ/qsDNUaNgGNla58w/8oy7BIR7ReAX5+
NZ7Ag/tUumsttlGLm3tPrTg4CIqJZ1PcfXInBaTYaP6n238yl0nCd26Fytwtpts3
Yed+0Bo34gTfpVmKK8byeTSlLB0+tUQMslXKjJM9/Cw+TnBoTMScK8kSVDxgJCYW
bLHPg4s21YmMzh34m3RePw2Y9K8HxJBgIs3FMZ7SbG/sYZODYzEjWzkqY2ZmhKZC
ZyfQdZ47EBWA3yOKhmyifX27AgEDbj08ax4BzPT3OWu9DteIpdb5mMBl0G5ouwX5
ys68t7m0nn5zsGSRWMgob5DArFRANOfSTeYBSATV5zqpfGP0EhLAwOVTnBBKGw1r
X9dBxzYygWejZDwaqtqvA3WzDBWvGemGRyMppJAqLfsnU/vKbAmZN6K18ay/O2pQ
gC8CW3mdXcp8gJbO4qcERef0bZiYg0Ew/bexHF3jg/eRmVw0p7opqmd0e5qdoPrD
pTKqnUF+dvwC+8E1aNQYAG15AVImtBbAgWwwS4j/xAG06/pbtC90smtjvetu2fJ9
jzdXEEhNsbAVD1Z/PxEwQusP7Lwzx4zvGJCP1pW0opV7swXNMzkyuZpHRaRSTQBh
5t5vcKo0g8Mi0+DEZZ/h0bfiTwJBgbDDtY8b/i/X/8Mnl3yGcYqEZbEE5ATWdnOy
0/fHd8253bGzVpvhZDriZ2vjoJKnsNTuKUzHyEyHti7KTl2ywZegQ4N4etLQma+X
IqVQz1HU8XN6/NZaZf1csCz7FawJMaOLx3cfmI+AncyUxaWRVtptxWwTo7VfqEFV
juW1xe8Zlv/wtGuGjWKNWkZhIDvJ1fBAo3/+KiPnVajwDbc/1l6SJtjE6GNPYR8D
umJpbg58vrNAg7EFBQUZ5Nl68yJWkTICB5XxrS0BTg2qfYwuWsYrNobctFxiRYBU
OR2UQMJlu5ULeWnOiG5V0+LZKf7Ut6DTpI3OMUygB6LEBGF3fv7nSvc4ORgSvGrA
eWSFAkAJX8dzk0PlBjRyZas403JRps346S4uySUBPhiDXVXAcXJLIDITwTbeVe6t
346jPzvMNu5ZS98Gr7GT0WupF5nJk2GdYtgAyYr8Sm71cYpW/UDbOOv66kGlGTvX
edbzSga+6n6C8y45vHeRM2K274JBLMngL1vp3trWBLGYhK1KQ1iCZKl4v3uYwn5l
2hCqFTho2KGtoXQzzdMpEHEMsdmoLtkdB7Wg1tszSWybNA1dmF3aSLiGgXZ8la06
rh9l4Xuvdqz/EwwhxdnTc858Rtec3D9+fJ45fY8RxarLhr3jBhzg45nRkicpwoys
ykM7A42v6vYEYSsszppv4MFEgE4L2dvN4KUKAg2wxHATOy/3H7sXP7WZgsdeVGPO
0TU5nyqlVttLwe88Gt3PH14AlyiLIA/40iQO+lFrJL3P3orGK3fDKBLY3opBGp6+
SBJ4NoDCSNy7jCEIx0gWqb+1QNV/nilAtdk7Dgm9kSFlckvoM58n/KX5SkqDKamt
VGUBKEjFa92KuoEv7a76B1B9hz5Xt5Uf1BaNZdi4hkhJ8BWLet87ngRl0c1Tk+hI
NS0Uph3kg4e3jin/WnnPYSqxpWzHkjIf5UDeWYqM+0w7t4wCnEWgfw/PDeMpH5DE
Z9Y6pskm7iS51+Cyz9d2RnzP1SiQw8AVppSRE2LIpFLIVDpOe8FSulJMUlC/lIb4
knOa4pDXNP0qlcAuF1hm26d6/Oy0ntHjWEqN1HwSauvGpQCE0diTbG4rbtLZ9enM
EJPDkaWBX3ZAyvRD4k7b9r/cVPHafnfjkugxoZ9GgKpQYJe44KCliuhsn5LK4lKk
RKImolzqMqhiL6tNpiJ+U5qhx01WzyuXRNuNk2H3uRbRvgOlUE6Eq10sUoU+qPYZ
aUjMNWldkcYR1bfLkkBiZKdUr4Ps/83QB51haJmMCLhL6S6ZjJ1raGlZMPKVdRA4
6ylsc0OiGuXn4Ip5NNGlxgv00HvnWOt9ye5vzyhjcN2z4Ogy6WlWeMOeLQ+Og9im
oW9+8hEE/tSUqFy1WLAxBXy+YFSRzeW5Hnh2+H990/ZkxTyPSYveaBQPrFmHA/pV
xtb4bjTFr9TVCFUkSuetwK504J1ay8rfIHdwMlkSwcVCUj7LL9f1ZdCx02qyEDIY
72skYgrO/mIl5kQ8ukwzaWNNuY3FZTkomj19Sguj2bvJb6L+lidDNBuDsm7uVjzw
QCiaAa1T5mL/tCE8on4CYlfp8VdGbT5BtxViI2ZcKTAbrgo1ZCzQfJpOcRVs0GGp
qSUt808ka3VLXtT93PyyZarrbJjanMlelwlCgGk9bNaEvkxymOnyok1LBbc6G3ZO
WEK380jsGBZxJajuQ1XiCEgrHm/hq1DP06v7Hv24lNRbjS7QS6tnXrbrDMy0j2CD
PunrOVraD5qFoULW+wuxaMLhT3B09mcHV2j8FOSoGRPTGHYJO2Q3/edb+6bVQ+M3
D8MAss+9lm0diniwjjYFeAULnCUmCdW01Sldme91BEr6CYCw6ObUxkkfzXpKY2Ci
yTjD339q61Hsb6NIrZ7fy7WpPuxRbi+bW61Ua1tXdRXtxKdTcMLFlCvKU+cJd3ZY
0BCGQuPYcURh6bO1uV1oQHzT7lf90YS9ABH59T4+uN6xoXH62tb/4HBUhqKveVAh
o0kJwTJCvcq+tOr0+eNdBD2l2a3ZL/vD8IiyuXgtTJSfIKZmxlaa2BgStwZpE3Mn
78I9vZ2CFLyiCdftOQW7wKjpdXW/uwINnXvcJI4st0c7MgC2IsnoMraHgCElDpjs
BrF95WOiKzoRfAuk4+DhzxGHNELB9+DjJpY0AZMh0To8eWceSv42psO1r3woP0MK
KJ4Ek8r6t3AoUoWWp+/G/zpAZm0PbSDHcrCM0bgqW+DEkOlV1YGrWB+i0efuyzcY
Pf4aa6g+qYZBxr9P2wje+igh/3zcQhtekrRnmKbbrNZTwxR6Ho5DRwIUMDHWRLrh
h75P5O4IAxglN9iJoo+xdJL44dZspswA3f9t5OedLsbFX5hqcoSyNGHjkSelsEQE
Zu7m7a1gBNpt2hctkhftGY3YWOOz3gIPmR26AdA7YyP74egwGdY6cjqOq7HQCKBP
+eC1Z8XoNN2lYpRgCUiuuNt25U7jj+Tt87/rN9DBnQ33SA78R2Le0HkCcKFOLPGn
fym4CgQj5XEL17M6I60knHtuiMY0ijwUkdD4rgc0DZ0ZbSCk1ACwxUoSogBO5b1p
BZkl8vALOrbaC5qJhkFkGF3BuE2lQyIvKcWHXv2RHGkF4er5RZhGmu0canx+S3Bm
6G/o0keR366zCexX+mR7H+cQeu8Qgm7gY0sX2jt9rRu+dtKJ6JEI/VSkjgLBdUGU
UXF/WYOx701834srmPW1YRAmLXXDLnKHyhHxzVZaDYiRjctBdFoQ90lUU7XxCU2v
RJPesqld3iawj4miyjY7CJsA3gJoCiuA1v0k1HiR5Epx+jiqjiW3MrqQKVJ/Fimc
K2b4gTl7wOTeZgB8DzZcB2AupYvr1NtCMavU473yNodkkaeWHy7keM/D4KfBGgZx
2MA+2xfHXHE5xC1VPgGIUDSPj2JMYg9TgyCM/gn2E3AJPuJJ9ZSaTH6TBFaU7RHZ
QMGBsmJvx3X7HCYR0Rb+zQaigEpncSi7SBhwxzTH1zT881aoZs4wdrgqd6qC99gc
jpm7p4c1bKZgaW2EKFm5k2K8nWbesb3DZwRDYPd+dMZ3lvTakM3NBQIxZzhZQA2o
138OEnRlLLTKyRHfiFWxXtBGut4tM+DhPBtk82MsKMRPz9e6ELCqHgTRJRuII1vY
UYg3/tPVMwsaG0T9EG59IvYNoH9Gohnr0L804h1UzHPoaC+uN/GZ4N4ZHEB2z0Rd
NS3dEQt4KCfVI5wqMB6h0XItWRiCkN9rHJi9cdx4rx88c8LDuyiIeDJsVjYhOV/4
O99WWnw8GJXnShn14QCh/Y53ysxIKThTXnFKaE8JGfrJZnvoOGqVNpFCbLmYUHPV
f/Ww05XhAIeuTJ6l6IYeUDaqx9NmLnNZb8SMlg7B+sX0KT0QYfGBvMxoPL35d+Vh
dY0RuelL68AUUMsUX/nmonp3bdkZtgZROAEDJ2J6dQcTkR1Oq/akuk/Hso8VDQcy
Z6m6O0+9R2+aoEX7BdCRxcEJ13MVJsAxrG+aGcewPTgPCDinsbGxs2t9bKk+5FoR
SHwB1wy9+CjLf9CFcaKP3Z8NMCkyX9HXch7ULoNzZvkfQALNx8zrAq96fMKg4945
UgB1lsbBP0KAbINCEI+smrDhoyL4K8cG56cewc3Zd3AT7SN6R9hMCtHsEdZl8SUq
wx2src3pQ2K5oB6j0UUiAn6v77jgLnPjBKKE7u2lAlinE/urL+TkwJW0VS2pbQ3F
X4CQWLnImmpkcoTs/QPim0KZ9N4O6UlUoBOwFsf7SJWEa8trLZqOqpiHZ1HruX3Q
xjdniNKB5gFwprKAp3BfxHXSc7ntWz3LmQuQg/Db9EPW/TVTMwi4lF46WcaJjCZZ
OZkf3bM/QdkMdbuTGV2eFDVo2ENQtuPENYx7mvZnDWvQkdNc36iswW3zDp36ndxL
Hv5X6MU9eaDkvNjkMZuOT2ubWwTn/Fz746jqWq9ZPz9nio2brI4CSqoPM8kyAf6Y
wTRmebhXoWBnF1Y8JVDlKnlNdJeH2mKMo9cO2Cx+zWnrqYCECtYun4b7Z82bHTMQ
SEqWw3XrzkcsiH/VJMtYTWUXqo9BToTM06j4ZN4YENNdQZhIO0p/nREab7rxHikv
ZjU5IHySt+2MmI0OnB21b4ImArr5HqmXntE7dYZb6nrmiBZPhoE3X83rDv8O1L9k
v+I7N6H7Iu83Cq+ddaXhKn+uCKGt2ZKv9+27u79ZK0Q4vDPCLOm5+5FezjQhNY3U
rFzW9AlZF/wJlFb8bzNMHft925oQYZSaJ9CUdRUQGlLXBzlzq0sPLFEj8+LT8NIX
4D5OMcNIG5XmKNtbc1+BlxOVsEZ/wEpZO65GSgXmu2glruaxgBmXrOoLPgFJtKcC
ijPvk9hsXFgDIipuvnuHxViVSof4AJ2jEUozPy7Sq6cjNfOltsoUGmj3hycrE3y/
qUHs9u9dPKKhM3d+rkXXmR8AXpfVhxEcZ7qJdoY6HCxUU9YazyKqDXf6Uez2NLz/
F5KkpkCQUy+C7fyNFYdolBmFzWhbETbDjJI6Rfuiv1lHWs1VPP/u6J8S+hiDFNZ3
ZicrosYjQKn8sSKxIzVspl0X5vthkPYvoz6CXDWk+OpJCM0RxCeNXBevWyUCT/zp
DFkv1/I8oMPfuMbDJsC/MR4azaw37B53SvcHOkm3tgPxOeWLiTwF2r7X1s7Uau1l
GyXfp+3HrsF9PQIcHiUIQwro3Ot20M9Rn4wZlPvyIzvmh1b+XR79CSxkrD4Qy/Li
lbTl0DuTNvEtO+/gl1A0zCXLNsANTY1l3cgUiOXo5OdrgLu1g3WqZ51s/ARFNAlt
/qxCD7Omt+8frIj9rALB2rV2EHhhAZbM4eQ8Pdnm+vvekwSiwnHhE3AHbmpzZ2GR
5GPWRVFbOtoPNHBdfNm3ozwmjwg5aFkVZkTmRvNXLLEUjoy1wiDV1JfD2FhICvWX
tNIlVBxmJ6Ay66Zu01jNZcaZUX3mjwgxzNRx7STtIfu/3XTXJCMekb6PaBCc29gF
zARUaFf63akWtKmwgnyN8UdzrwBALcMbCadun7McgQQC02mFC40YiEPtBwzeVUqx
3+I2IBOF20ltaqixVMsXyyWssgr2axCBvzSs0hIfJq74ZTZkOoU4U6rdiBjJ4NQh
u1QFw+0gjVyAjpK32zuC6/ZqoH9k6ezboXaQOqjmPx3uK7AiZ6ay8VBJYyuRNR6k
wcVLMU9ZOW4YBO19ntOTH0gN0uJ2q9kIGCv8D0MHAt09tuJFGFC/DBb8Rln6CkUa
siw6Bw1dLQDBrbRh/1Jjgv4Sd9ZUO3Xe/SkGoqir+g9bJyBrerCG1KJr+o/o6Gey
XBA6JvgNIkPc8XYPu3TvLZk11NJU0ddVjbchPnXFMdq4IM8RTqI1JmOfdP5cxQZN
+fFvlN64BkxdBbXvd8KzVVgllZx2tbFQCNlSv7AbB2GiQ6LltHYzYBawHqh+QOQr
kyhdQeV0EmSJTi/xjitv4A0i4g2NF09NtOxMpa18GkDO3UFv2LmpmbpYpY9WgU53
4O7/lgUahev4qfbTT0LLi7M3HX46ZLsYTgeQgwGYBCGb/ujXpkka4Hw9c4WXdfwQ
HjR8W3cNtLdNOMbUqeUSNiuwdAW8M7v7q07uLaij9X9si7uGWPIr6WvuoO+FzENe
wpMtTl7La50qBcoccbmiOCEI67qmw9AcgEZzku80PK8wyCkkHICpkFpPavz1H4dC
NaiJHhBQSIQTROtPYsv2ZLL8iBLGY4tglni6LJdlv6GVjXy5fsOgxl6XDLJ1l0td
vF4yHYbBLZzX9xwWGX6BIZfEPw4lLNIYNBVEZgj225a9ewo0JlKdyA6tDNZY+dP1
4tMyxnBfo/HbzcyoFGDVwRiMH3siPU6ooKGXrEJVWwi29C+F3YGSvmdGBS3dnGqm
XR0i91bsMZl/WDvOsmCi2BYsNmxkSnDTjq7/QnwsaDxhHQrN2hcGUcMUgl+5XpR0
UR2eQ8qfmqtYvYKRZ6T/UR0nZausw6J+B6c1sPukixj/ubDmxorroINekbV3UYQf
w+z4buuFbxuic8OXwtF9ndR4Td3+gRyDErOriT+cIMpTtUAHM0tO5CnQrtWNkark
eVYqeSULy+lnsavXei1cf6RA4QHWpiF09rkfhd1tKWwLB646ykGG8/3N0Uru8FLO
iwV/H5tIDmbv1LN2+XMTEqjlzCPKuCTRiaZIRDFpDvJ0KpJsCTVxoCmSgYZeSIKa
atKEBoFsynn5I5eK5uxueWml/Wl7bTakDWtWkRvh5FfMJo8qU+tJxeEFpr8BwPPS
a1DxE3Q5n6ONXDtq0XW/rn4d4S7y5CdeoWKNRUfI/Rzib3PQYdJwVGgevb6712k9
8WcNi85psMq5JoJPA5fkUcnwHuhXhHV9ARxiR9/rkcSccNOQ1V2p/8mpG7STYAVw
B4Ht3f/Uz4cR0Mmooc0s4Q2ofohMs3tUp1sdhhM2AhBlOcCs4mqhx2pKg/g+lwAU
L1UlE2ZwAC/YQgymyAEit6UwPZm2rqyCrwnMaJPQR57SPWG8gFf0xJAjyhB7M6z0
hJKXFRs3nT3Sb0CNt1mgJ4oNc2Dpm6zeiOoF+9moldbYLEmOt4lVibJFIovgtIhq
qcXHKSnci1cMhcotijjzKUhK0hKcTbgpdhwanJmtM2QTKzF8vAZ6Q/6b7Oq1am3s
sgzb/7JCr6aDTypoLTQWN49YPOPfaqTTbXgb+F41uGz5ZoSMti+FBRCfYdktjus7
YAnZE5C5iwC4alpULkmUR8sy1ClB1hSMqT0gwoduYooCi3p8NIP2ezq8JcTko+VL
SQGEm1nZsYiSoPUnzPfasd7o8fliKMvEZE3UuTCE0xp/ZRJhKi7EHVsV03qi2JlA
DW0Ar4rUeGgzed7QefutUdM43FcCUCc06NzGU7EKFx3FHdKtBjyjDmAPrFExs2Gs
9kvvSuEQ/fxCarXV/Tl0qlsOKb20uVIY7CBRmoN+1DZVdCTm9/SXPvcLqtJRroYd
p9FgE7h24F9v69QHfgNIjWSyktxkjd4XYKZx7TmkmHlGvCbrcFp1VIUfe8pJfcUc
d8ujLWd2zmZZBSweMsc4JZBFPCGb870ttUHZq9UjsmzAFq5/3SJhnYxc+5tBb9Y7
4TdqybZvvARTDJJzwXzEzXZKKJTB4Sv84iQ8bowHS4BAi4pKsTh5wqOuHjQiNCyY
bdy8FkkimWd4f9KRh0E7zQquYADkTV65FcfZOGGuMpp+I+vaoQNMbbt82OPCXBlU
dkivNvM2YYUr83oUnFBIlVn4GiVo9wHj6JLdWU93OGevQOHYxz5eIoNjB6++spxP
MmBH/r9EIXrWKDcilDj0wJuGMRAZHp83pKzsNPcIBZIDfZlf1eykBnCsNcC6J2Nf
A6xSikybwjNJxqX0FUYKzFFsitxOvI+UFbQ3jwUJvEkG5NaZ/UHtMUWEWg5q2tUv
U/rdI2YDknL8wlQAFTwNjz8RGHCW9MbetY36PEcEOlmC67zgFm6BdCE58TSX3IVo
Pz6SWgU4w4FSPzVSbZ1O9Wzk9fsG46Z1WUHQAdLHgrVq5N+jW78hTGxaF2gwfazJ
HDmefOtkdwqW8Ao+cQW3PHujXt7YrrKCFgDTEWGdWkHfT80AFH3jpaJi+A0KyzR+
02NE5Qmvenz70K/ykmF6GNw/Q14jxwCCO6dg0KMcjDY/aV8Bevy5PY/U5yrIfZfo
ADUfLIGStuf8D3/6tthoUl8np+tQWGco55yFkrQaW/WiyQUzPrFw19HnBxGLC2xG
4FEcpU2vl9FbVKj2tylZI55xKujyBLfKuod/doHlw7gQlGTZen+F8OHkyrfoZ4bK
/+2JjZ20XWhx2abqglokdyxtyAPIMAAWC5qNKQtZn+LVVVSBe4SMbp+fRjelv+Wa
PAJ/1Dv5Fn+R4ffbJODoPkzb2VKkFOj5Hw86aaNZ9YMP9EhtnXMkStGSocfvun1n
mfJeOndOj1jUQwaDYwNItSBmuVzmpwwwHDljdO9sJIHxbMqyGIDBlJnhm+ak3uqw
wh35Y0YoJaKe7TVUemtScH71LGgE0McUdK9YUV/Rf9qsWzRGoYKNb6Nl+s3BVpd4
QWbbFTrGSksPSGDa/4KqtdlTRb5jqcEf+IPGSKUFYpG7FO/vbQN4SdmTG+pm9Gj/
2OyEJ9nE2GKhfMIIk9Ca9b06RtkzXcAP9A7QCBCXad/syyyJvEet60jwl8pvKIE2
HdYbfV0lHXwTLijokU0XJE/qydxW+hcta8ZSfS0Pr/gPqNdh3h6NXx19LYNXe4AJ
QVYHMrZfp4TNMUXlbfJJ1wie+xqi3jkLVLVD8LYjYN0BeFew2Vnb56DX0MZMrV2q
XwY7yt1/hHmGidXxfWyqFiHqINeZTYGSxtOwCeqOGniIO7jPUlInNgS6f/iXsR6F
fgo5h5kCr6AO7+oQ01QLCEzlZ5YsQ/On8XbeyZXpsvVkkoK8GdBX0epeVb7BUOXK
ddBK8srOnvRfgz8G2+Z2pcuv3MBkU9kVc9yYCmGHEvOVAjyhPem9j2WCgY6xjCJj
CVtbFa1hZys8IkjhxxwhE69lzMPZu0/WIRzP09OwR7ZMd2qkUEdDfU1dLGG6PKeo
9kVNg0bwCAbdMW9ezfzFewhkLOEZUXajDqIu8SxtCLNHXojQ0vSkN8Wry38Nu3to
g1Ia/22jOIFRuYCh5npTIdlRS/YzxXRdDY3AnjRWQc9P/sWaIJ5HvlRshnASgxUX
OPfEzQd6fTbT0tzKgopnMXpGZj1Yt4r57nIBmZrAEmNxFqQ5ogfJbrurj9ACxYQq
XPrn3xNVOOcNjlbwow2UnHyYvN/rQHrtPkvnnB4OT/c4cCli1ekgLey0WcLO3rbP
9FFD/KvSyGlRwhYvqP0QDQJQazwfaABWWjOaXgOehwN9OKCF2p/naaW5GHKR6kzp
SFyXGIfXDfnTtmWqC2oZFREc12/Os/UNBEq8adI4akxLUB4oyhlOMHggkbA62aNK
wIUzrtiQkKiXsJnHZPx5lYzCoIu4iK/PBpl86y+QT+QbrmJyw1CjN1/CvfSTvYJZ
QZctmiM5mHiG9gBIdN2af8jMvz3YdNV4IymJbTNCS2pLhekchzs+yOIrO5ovjtdf
TeZsGL/dgyYKZEiXP55Wy9xLrnSFXZ6M2BSTUnqE4uAYQJAl8YMqwy5pfXf1qT8B
RsI+OUOnzQ3w2N4UmMg6sKQ/RxEtVBzZedMR0qYBb17kSK92scNY3PXwcOsyKzsg
ZXp0RHELuI2mdr1+qxoPlaMUR3pieeyIeIsL47pBCE2M57aeMNw3kxuFbFFWcvH+
7K3KiksDCpLQNnGrDKP+8CLSwrj6f3s6yDwN3YWpdm9iEnEMehThdH0qMzZOoyxj
Smt+mfb9X6gRuuDv0fAavjBd36OkK89rqynCk01z7ZJHrR3c3TfZtA6k+MsvHSNL
RsP9ftN4gKz9DDQiddE3kdHY11Wuv9v30BdsuWuwHOKxV+Bxw4pYHlQCE4BLmqzA
hmmaFtSE5HDrlEOyvNYyhgVKb6s1Pa4TKMdSax/+b8uoNd7MZ3apmLc2a3GjZYJz
tNfFmHYMMwqbqECyaMY/33Aa48kA+YEek/X3sGR0ZLYDWXA9HCi9S0ytvXrXn18W
p+eSTZa5nfGWaEmlbRyINcUnZx/lntvPooHLL1tJ8eWzfuO70jdvJBCe2dITxA8X
aBzuHebp0tI3LCe+iovvp+VuG+TLxxT+TNIQrjuThBPCoB/eq4AKscPqIN+eEr6s
SQuqmKOKMDtSYMmq1rGpVTdQrdW2uE0s98IGv8gOT9wePbCYxgtTPKnyi8vpDnBI
9DoI1c9//FxO0MXnH0u214m3i2UKCQFo3g6ibJbd/GNOoYwXJcDVZ7MGFWPI1StS
Qnk69PpD5eC16JBBQDrR3I0dppnyit91udvn9+37H+L+A/+9skdHvif94C9jz/Zi
2tnreIaVKL5nxbRcXonIZcGdbDv/SrtohiuDG1ilkF6XuF8kDsPBhoieJEzjpx0M
MTDA4duR0MqjoysSxfwGKn9oHj76jh08s5jSwjcbk2zFN3ASdK+nJ8vgqN2/HEM9
a5uDs2CXIjRe7ai63WMH3uRhsyu1OlA28HilygRSsIgPlhpj9OUJfltaa1LoArrh
kqbV+cFKYSbSZ0BKY6ruCT9vxKPK/OGZqscfV7+vB6AnNhL9LWyFoXvoZQZAL8jH
aVZXdArTV3iXHnzs4qA4PzZ4/mdmVOKzvUiwX3h5/gTZ1iNNVcGdCgj5MDA+mZHO
/RZEZSQ8rzJom3+OerGgDaqCHa15UG0bAUCzcKo4IhMrEuLGo+dSkPWHEh6yDxDc
Vfw6VR3yalj6kG+dyf+9b/XbyNimJlYX+Q2GkyTvetnheLU3s6M+X/8UpfTUpIIV
Fj1FS3Lzoi+QcUVIbjd8ewJhqBpy5mb1x3BXGLHc6q+CwFzaR/WoI4NslmVOIS4E
g2jcbOYVYeRYQ1r7mdl4aEXgNGV258BjX4x7PL/scCwjIs4jn75oWtbU070o2emo
vFwmE+5Y1HK2RZ5vekI5IHtN0uygHmlKNxWMavOJIkH3FMfQI6pCBKLU9M4Ek+px
Ycd4cvfWD9JWVc1hlmq/ppQ1vGV905hS+mRoJdbTYgdN1JI7AmQ+sHw8xvshzwLb
xgAOVqQ5RAzVA8Mpv75e+vwT36GG0P44/O3KuhTpnlPkQJUFE6GqI+IPR5zhHJYB
bxYOSwiNAQlkdvG6x34ZIohZUos/CeX94l0+Z6knQG58siHPta9hUFRwVy08uTJd
RP9g1d5xqQxqf62HbmgLPc49l23WOLcg63Ah2x4PI1NbkwXn/uRwSfcnpsbmAg/o
bIaFcl8GDzn4NnfomjZ/dG7hwWKnx5fn+zqpPHCuuwmA8CQVYDyMcVMCvk/YcnN6
v38XxIu4o8B7dijqRrj8bMbfWXM6r8jjtyW6c/jtoReNbvA1pbQlLjag0QXNB9ao
xyaC3CGRvrsj6Ec/5EvVIyCboCoHn0aG0jeqWqzoGo50hTeNHkgFxJI02pcpJ4vy
TPPtmrxhLi+IeX7HxEZcznypyyr7HKhrHNPAbDUQgMVYm9nNTJ0VwkOSVnC5akqZ
f8/NfhhGxGAtBu5gKC7l29Xui7Qam8L58eI9bchAiVD0d8YABi8PdGk56gCCDC+j
PjsJoZmBRjEXfYn81EX9b/69YFmn2ESAQt2/5vOW5T+oXSlWJJ59wxmxCBUVi8hz
XdTYAXqrf+UytNyR5fdzYLlw+jf30QSSQIZ/RkfEv9E8tfusNp6Z8+VAI0WTTxwX
fdR4g+n3KpDiSXjPaU9mCLePaP+PSdg0Ut/ybk0QuNHSDRd42Rv140BDlzfsxcPz
A4R3N2LOc0pBVU43BYmyCe/5z9ybYFjLh/iYhxLmLU60ly2bI4yzCAK1oVAt91jX
J+Vc4u4WJQF2JgOss3scev7g89v/N+18zce9ZUeIIxGD8glqf3vMFK4KadmrkklA
PRI2TdIp1UBReBtnM4jnfZ/jUsLhIajehm/JNMGa3fJXNsLzVeyt5a5rnM5hyh7D
4e+8bI7/hAQ+FX+oOk5y+7IJtZhX+vpP5i61lNBf/KyyKKBCPsKKB1UW4Y+C3VzZ
ptoAaIznGK5pPmdtTu8eroQd+uAGu1aWqBiuxuNrVqF/u4YOItNem2MJLGz+6t4E
HnSzN87p7V+Fnu3UKJjBN4Rp1ss85hkemKLUnppS7b9uAll4xjsOAqCT4FS/9jAj
Lo5tHSTtk506fpWvX6H9tmX5SPLNsVx+yAKGuTfHSGNmItnNnyRScw7lxy3v8dVc
EjQrVzG/3XFyecc2nI/FOFA25+Y6gebBRKrYJ6BLPY6/sznIxmx6HeAgfhEtkp7t
hdhSQm0aOGBomgnR5xapqbPM6kCaibwUh9aXkhut+lVVA80aFk+UCofw4ZYRm7Wn
MguGy/PsfahiqVPEYgat1iL1+1h1MXiO+wERfHXkYxodQArZZozCQQs8+f04CFza
oAa6T2NF7YK5p1YUJHE0A16EEGCfCGAgB9qeKOeWS9xdvY8VgpE3x9grCxDWLAk2
5Q1ScPLGdFrtjQnCHmtB6og/DHFUhJHTVpaNhgDzO0a3qfgCg+w+bhrsnOjRtKQo
/upsnKcBNHgujPdjNoVK2t8SYMVnmWHGTJtb4V9a0Ag0u9kauc+uRKv873xvPPMN
wQ5UxzECh0awMh0OqNYyk/njGJcz1PofPbqglR9tEQO7OqtDuCbrTx5fWrQJQ2qX
aK/j6kNdIjvcwprQE4tOqYF2ijuBvWp6+KTU++rau95rjD5+nwlHve+nV5+lY+G1
MV1yVcbex7Drt+eU9vlsbWkjcxLueWr5wTBZXHAdNAvAaY35mFFJu4OUNqEZ+Y+r
xEAHjwlEGd0FkQQB21LyZsYu/PtWmQdSl7aPS1do1d6E51A7MeZBqiEP8Ogluxta
LNCvnvzgUoWiDR0V8pniq77eBV2rEVEoTAkHRjcEwnInBNDJVEUr0xT+642dF7s5
iVLf2fQCS1g6ptYX7qvZ/nDXrJan4DW8pWyD3le19a0ioUFWzdPD421kjIJ0SPza
Jc2c5SG+yIFyaGo14k51g6KSlxDwRQekgWhOfztaoqC0U/bGUoB/4V3ViJDqAY2M
f/vXrY37hcVU7vV4TThx+t+Ir6ty4bALjA7xah601IhEM1e4LP156Mds8fKjeTE4
naeGaU9cleJ3u6j3xEakolXyS8nJygdbYCVH3el/jLMVQ+/tOGhHP5DO1lPPhoe7
ZcqzE/h+LJqr8L8zpUj70IhiREko9wbwOfTf/tE5W8eHghZUMA8k4/uTyu1m/mVv
LUpePwH9b4ZnxNrXYie9i5YZRnYCJDGqGP3NBtJLoZyrAlFCHcxEt9L7AU+iq0bW
XhcEe0+KlLBsWfcIP9HiwVtxp2BSF7iS+Fc28NPI9CfXFru/KYccXYFrRbY5XL9k
ihCK17cZp20B0/dG3OsOgqC4JJ847jUK13w4HovB3lenVCF0NvIxL3LqYOm8mEOF
g4ID141dwKK06D8qAFtPhBFR1GWK+kn/KBk4j0ro1hWFTupNucMUFu4j1jKv1Hb4
c5RDSkFcwo3pxISp22DhRPZolcyZr892T6XoQmF2AqgU/wRKE7T2Z202t/RuWfBT
SKqyHlaDUg8qeqP01m9azAJTI+eStzXzwpYiBmKbrDq8xfWMsVOpqnlI8EZ4ISPa
GsG/58ZaVal7cKZIutvCutCSc5GNo7JwPQYOojHT6iN3IBt7OIvQPqxtFTQW5v82
7lnE99U6YFzeEEo2fmlrzeHkmsi3AiRn5cxdgxNqHQZHO+6Zc3ViU2/3fRH5Kj4G
Bppcbjqm09IenUzMdBJ+JxaLguR/aDCbDQoIElEt6NXF0TvhAaowOoQIjDnltnEH
4gH0Qj3BuVH5hxvr8nWFmAcn0iIM/icjGehf4UfXOtm6emwbfmR4a6Q4d0Y+lATs
jR0MuyFYTyWN6tK+wHU0ZZTP4tv+v52T85p1REyr9xWzHXWKcreyWJoS20TCPPAz
Zl+80Rf5Mt8dvSysVUvjgyXftDChkAnfYNCUb1AjPpH4h+m8u60sEWjqzTiwkcY6
FxSFS9GRfNU37oYfgtEEIOtb20nord+ZGxfAnSvKq1cv6rrwr6d9NH5HYMvAJMS5
H6ZJrCROieizm21f2Bq8LwcTIXfuggjoqpbUVbwCwUBuO4pFZFUuKYv7PXAl6zf/
s49uJLFQQLdbLKwOK3d3Gv7jDkNYho4Ena62Znj1PCcrZ70JrmJRMaQBKibpMO0f
NkiGgRWlAlw/XM1k2ULHRDloPofcBs1IYWS+U8fEDohRYiDhA/J0qSNXdnh/5KfO
wY4sVT3TckFAZaRfoKozz7stOS+I5U/w/m8BTMywEA6R1Gav1nqIzZgGSR+vv9Dq
H4PYdXtYqjdnZJiLQeeQe+tLVnuzZHfhozvD2tJzA30DSllz+/1q07hhNBKabtF7
npfin2/lZJENJ9wfhSjDz/UNC3zsK8NZBXvIyrb1oYxv7S908Um3nQfCsS4pu3WX
on60cD6U8Ax0gIDywxfCdheSDZyP3d8s/4lVILrHepwun7lD+jmUHKyQSLsCrWDJ
E+kufgNM8ig/vVHYaWcr/iccLwB1Kw6yzFuvwOYIcaW2p41Ov+WXRmMS/UuBAKTE
Aj6g9y1RPhDI8QnHly497/M6FZNQ+P+7W/t5zqB6JKWQRR7Ua66ZbTFgmr/BjxYz
1LF8LaEpFsbYZ2ibmVosIK3HBcaZRIlPRL15XM2PoAyexocFrZZB7Z9MSinpiZOn
hwJcbo23eD48GXxyuCMajMFiPKePB/NhqQ5pIxigzUU2QogaX3W65KXkAB/vUi1B
2trLasetKOhFBNlD2gLb4xlkh4DOD32ytK1FuKbSfnrd9DMogJjl3LAkCFrVvwFH
uAotM0rcSJ9fvQuQ1nnUx7E9Rat41aClWB788KO8CiwImdtHayRZpgJgo+mKteFL
M858Jm0razV+H9CRQZp/KNpBPWT03zkvnTV7a3LseLMlMr0T/Zytlit9Dtl1vK8z
36V9FkeiaGT7R6+bU5LjwIV8815itzmIs/sHKN9VxGCkYmNrAa+XLqLTWBDCzGDO
xA2hpId3wdRBT9eBTmFitzrpkBkiRZ6ZSzB4T+YKPdx0wiCcMycLmMeTP7io8cbF
kFq+/KcYd0SxnIiJYAMpX79LHGj2/KXrwdIll+Wiaoe09gwJk4NvbtD/sxvJeUjX
MLKQdSXQzDaEIb/oJBjcmpUBlfHQv/g8nbYpRasC9zVnYq/dxL5SM39iIzo1TZme
B/hm26aekAsyq78yvfqTZu60aenexJFa6C58ceN/Ex46qnElEyo90JItZ8CZZzbh
jv2uGYoSUH0bssJ/Gn3yE/h2I0xBicjJV5bkIyg8KtTVzSSTtkx0ki+FysPH0CWe
xavAsbtZtE1KKV5WD3g4xXczEUA5EyeBWGS83sAdXfpo+4ZELfoL2a2vkMVgppBm
ppQ4u0hd/aTt1cpfYY1JuNubKCIncFoj4DapsG3L279Nc0ebcOPSeUPrs1Q7xHMK
+1TN//j7KHfgDa4hQbgA3BGkg5RuDWFgPORlEpZU68L0P9lsMC+A/VaPGfAo9wSc
VuujaNEb5QeZePJ1yyZX4gXXyiTj+Rrd4KpYWpQiK7XL4x4WPWZofsip3zlchtGM
59JEAUiPNJ+gauPrpx3N1w3jCOUOo+NVnW6rGsMU6igl8FVT6+GkSzOWFdBJUHl7
HyjEmKn3GrPEQ6QBogfAelbiJqrRHNOBXA6KkBXCNG3D/L61bnV8TxrloUwFQ9mE
AXrIwH6L9IdOMizrcmtXCryDy6NmxHmc+9XVrcSQmcnlBPTCUSJj5AMEUXHoR5zn
gpaiSGZX7pXiAOKFW9TbONNmBkyqM/4JhQSgCjopcorJraMtxZfY2yjZ1jwxuvTS
gOnvDe2C7oDl27VTAl2hVLknzd8OklvJ1qRyhN4vJTq3+lMVdYp7P68Umvh0hQyl
q/Nyx3mp9zxujx1HjH3xt2rVsKwPo1uy0lsQNkOasmPtWW3FDAXbBEt70wL6sic0
7rWiYnSfL4jS4vZTBMLS3qiHwFrX/8CMHOI4Cu3Zu0QP/ImUY0hNMafJ/t6z1XCt
aS5FGXYpOKrVXgjIjevjcPiV/2mAk2v6gzvjDu33i/GA5NxtaB5g8foGDwqO203Y
t0O7CVYU4oclE/YuNkNC4E2OafFRfPpj7WEGH1bJj7eQxc110NADf+2yzW6PihHj
7CCnKQlMHdzI5EgcP77FPdKs/Uvshhh7yJlo1KaDWhkFh5hNLHHECuqvlItlxwVT
UN0TmM1gHK9dHsgZ53lUC3ZmVxEcpf/h+r1dQbBBcCybihSaLq/B70Jljth6dtbh
IEt4RelUvs7TyW3m2O4HMGXsf3GcWglg7RI4lUAbTfQ5gNrb3gcc7VouEW+Ot/9S
XgrvL6dqBkbeB3IbxgtUpPn8mZVdN6uJ7fO+qJQjIr7x9jELW8+/o/3ojUPwbBPq
V9fJFOrcW7jUqYaeI+W/bUkyYAZWm03lL+pK86OesTY8Fq3it/FdTMbA+e3BA+tw
ZwP+TtGChNKddfRJ+xryB6Hhqh3tQVWdpgCRXDmkyoke8ofR04hOJ6beSG1Nr7Qv
FWsJjNP2/lQc6DeZXU/6hav1kWCyWxN6TTipZboOjJl0Mw0setsY3B+BKNPbeQ0G
vjxkxgc1fPVtPX5KFj4eax31aLpkLDleExdepyLZ84iqwUvutfOZJoDaNsr9JgnP
WDQ+HBLBOq43c8sb9hqCxro+ovKiR1gGAb0jIpTEH/Y8nFWu39avrys0mfwGthyz
jxbftbauM2xI8ldCXM80SBzzdZIFaZF8c92FsU6qL/Pqw+ohUrgVwHZ0ijglPmqz
7pbLaTv3j0ywnApzVELJXN+tvT1V/+b4lMAoWQeG4OUD+bhlTSSk0xyuPC0+5Qg4
lFE601jimlFYgdoijSf1+WMZREMnqmj1CWmXQHg/SlL5syH0fR2xfjoD2c1z+EQD
kruPHQpJxVxHuajq3j6aN47MNDx072FQWtM4Cs5IzsUhoVsakYLVogx7NNuXNWhq
o82z5YrJ/oJuGjBtxSBE01nOzX53CQQQofRWYHBNyKyRs3D8qZMgplLx9FvmtdrB
HO/n9pU9Z/bhANL/fYPh5PsCBatMCD0gFzzcskvlahUL8d6KdJT9F9QnOmx2/LN4
aw7y/XVg4kLx1ibm8vzNO3BdBELpdgSrcDc0LLSYiXHPlQn/9LsSrO0faF1IFSiQ
U6nyovSfP3a8C/RGAgdv54MhK8zk6fi3PkBfSg9+zlg8rJ2L6zx2/FlSmkUEr6po
SqHj/uuT0JnSeaweEWiKrLnTAT6Hd08n8pYJldYMgv3EPH8xbD+w8u+ljZJe3w9d
8K4SeSS3x+G8flbyi2eSI1ZOsDrOnwgqaON9WJojZkXDOLHzv1F8ti3OSAADsff4
q8lVRfkam4uVWbo2DHKuq4pDfgKnk2bxyM2rpt6NLQNarx9veFlVQNI1wkhpWWz6
38qyAj01P5GeEem+WEgQJr/1q2zrOoTeY6zLH7ry8LzChTWtzhm6kijAsUAoUM7e
RTTyGB1N31srw1mFpKQJDTzlKWoZr3yBS80ie+34+lPvhXvECDkjM1MASLeJLVD+
yMyEtgmoW4iIDNywECMUKwgx3BwZ9uRIM29Kd1/Q9eKYUsMb3MkFuFhYXElGgQSs
9mBq56YIPSRMDk+xvGbeD9SvTlL87XOjM/fjqdJfZcXR7bG1Rx/0wA3i6hNmtxAV
B/tOqL8aznRCHEb2Gu/quexaSeM4WIdExAz/54e9zqAk6Sa2iFZOe5xpeYh64+ke
9S/WiEdDXP0ZIvKBgjski+yTwkH9/ZYFBMV25dGwi8y34xc+8e60etVUbYTQo38E
U+7FieVMeuWXUY33W8U5efihh6CpQt79ANXmPrJUe6myf6l+9QTcK1YtIfgn/rBX
elgwRRdzZ+yvOihnNwiT4NyXTDFQj+p/9mRsu51+VMg14U01rV6hAkIHAxgppbk/
e4RXq4Yyop+11Zd1mYTigxVQNoSEbm2RSmwSYF8LJ1RPaEJTYaQTN2Wvj0jM51SG
SHi5uE94RX7yKzG5G7ATCV0AXM5H21As9ic7EmY0QIGqJ0/3SaUyQs0titfzT7tV
4lsH2Yk7MmkUgtpPxymatGf6+Krkq76FptrpPkK79jd5Paicq1Psl6uZROBGQaKW
5sSyVZO8ns0CCJVd/HD2L1DzyfNTfF52MJIrVNCEDeuBoIdmGSCX3cRbo1pIw+PY
JedwapJPQ3HydRTlE2jXmTXFzzi4Kj9IhyKZk/1vsc6SaAPiVZEp8vO2pOlfxccI
3xpq1tNd5KU0+DsqNlThKCXroHRx0uW8FeFslvRM44T/nuukyUoXpQhqKhC3POGN
sftZoB8UZOlQz+NjmV9pKopdEMt0xZqQaQf9rzHtq8KBo5i0iv4mCP8htfDN4XqE
SKqzKcte4Jkz8R+SRR9wdzNXnFC6WE719X3I2aRrywuC6CsVMYaPGEGTHL/F1P/p
7yFTnnkKyhXxHRrO6FmY8+Dx/L3aQ+2qEdOSUOFWhaYxEh3jbCiASBeAEi2ep+qD
sCPanU8WLQCAHdRRyofo1KhbgCzfyLI7Vhb8bQ7gAL7jMEZQka+3yv93Gl4dlXG9
fWoOIaDrX8Pm2nUYIxx0Kmi0DoEH9nDi1f3EVZTI+asti7DU/Qn3kggSEZ9KR5sX
DP9mTiNshwfs9Rly0ZwNUkNbmTTb/61tckjZUsjhOKc/MisChc8e+rY8f9zsIpeM
CwGujWJTPaXEe9poYT2CuM8xPAMdaq0aAWwio3ZRIoGoFHia4aU5UoAmYA3yUMdD
46NNCRIm8Br+CKTJTic5ZNo0L2NVohhFcqHDvWXIM6nKCOSthpYUbeiqlknU8ZQw
9/vd+y4jYYfRcTBERFhVi6jfpApj5rfgtTUI7iCu+XgCUaD6MlPAZHjDBthDXo7x
osfUNebg6aYuCqRSoXFJVAqi1fGRXNGn90y/mAz6vqkJ2u5NajoclKlduCPoar8u
eAdzTWAGM4Auo01F0TOmJVAJV2IjycUvlEfoKyQ3I2bMXd0KMNPiQ3IJ1/bN5Nq0
V/s2D//4RSCDkKFfd3YshT98PuhJX1jblmhBIwuIc01kefrDOQ3Y0kg5s3VjjQnY
Wo2u5nXGUjm2ushWazZJVyaeZlTw1p0sufqPd3/yZBBOF49/Zg56juPl8qhft324
oOKy3WH23bJ1cXqB35XbHOo0wTgrQ522eDVpS7m3XjtB/nCAq49ZkAJKNwGgrkvb
Unx8zEedM9bCsuQux8zoqb7oQ+IMZQoAuZgH0q26JJSJVBwDFyI3do8PIsBCkH7j
DzDf9QQdh00tIpL1duGquDlI47siG7y8bOtTfLcJ0bb9X4wF/ByrLtNmcBtEgx2t
5dxPMIoRSVXIEs2f+FQIA1PVkwb8LJmIpxGfRDM6Rl4QMhhQulBXLPml/HoAlI4l
dPfcBBKKU2tvK4OgUbzETZFEoGx7NtFJmPxHisZiA2VmGb6wVU6PSRhXf2Elw79G
3C8dEB4GviYLkqmkofn/XnwJVyBBMkj844kgOgnwjM1I0cbSMw6I6maMVBn5gm3N
lV0MQNAkifD4HnyjpDXFCmc/je/rcj6sj7/F/vX/3wzDHc9JzWdMEC5p0i1VKDAL
JHcKP5Tstn4YCk110V9h51dVTApiQwX9QDmTfMYFqncTF99z9OqtUQ7Qs3amweC/
df7P+pu4IRkwVFfA7UbH2fPPr6sqhjNuQYqKvMFf8LUcpwDyT4PRsmA1gPWchlbY
XiN2l7d247GLf4vWB1taCVFmRj1+K9pP8hAboa9yoypLM5rhr+eOq5V4lgx25UwO
4V6MJrIMwKmalFRD3whKZz4FEKoPOF8bTVJt/U7fojZhRNTgiTxy9gdVhYVR2VVR
F4HwLbUh+NfPUIR/sFfn2NeoCOlwEofEjcAz3dwrFUvOfkFlz8sVZwtCrviX6RCR
WiRXxKpoq3v0olgDCsy5Etv2BXUqewz2aQDuDQRJ+z14mNfdvLE9lpRutArPZZ3E
vJVxdGuedhXlsYjWLYsZJudLhuPyvZFA4XY+LywsGDTpoTdyrTNtBXRzEaXv/l+K
GAY7Eje5x/52XSq+xQTFyQQsL/xFEGL/kMi++C8NgcP3HmH6BALbuR3TQT6nkSDT
gpyiDJook7TQdLpRKiB5YrMPFcWvYfO1+T5Car7+Btlb05kt2GPSIzkPNhY2ZfnG
9gG+gsGfmo7xtllF3BqZEK4utfRU+UI+xNantcrfS3QS21Y9ueyV7dAQwZvEaGoJ
WH8ZZ8eaVeDkjrg+17/TW2EJDI+fVA928jQBNBiZAUBVrcEYaJ4cpwAIsoqZX6FA
PUqwSn+MjotgDic13did9bTvKkn4kzmplHgs4x63p0GX3C5K9R8Gjf9nS3+qUSBm
KHUKDnN9Aknbe09gG+HLTPLAjGvB0L2r3ZDjlmSJ81f0zPx4WodWZaP2KLP90Ms7
Kd1bSFQGUedVWj5iIHW30l76wuqKInCvG9gN0Zg0PQgZhLP9/H3XDgIgoL5VCNku
225+a5ai6d1iT/lCUEVCBm+FkvoxRBKW07Os2r78ub7HRfJHU+Wkvhei87G1B3tS
qmYZzQwIJh76XF2zvzLHTLD0MHkQ4jX4cGVgVJ7GsXRhSkhuEM7XkNkeXIlf0Pzs
I1G/hpqKz83KROf8eztUOeEkVBKV2hAnjyTbbmjbOYuDX+OSKtiIeroOx6fabxqa
AwJsUeWPSjDFeA4ULiFw9LcqGqk8nE/+O+uQ58H+4/UmKH9ZvvLOK11XsieiwFXx
c7GnKSPrOXnQG4A4zFazhSSIgSnqP+9c6f41Gw4Us9NV+NQJmhdx5reUcXK7p1Xw
lZWsihnZBefhz3on7wlO82qbMchDldD3/KO/7y2aCzyoQMpcOYfnXPZDPTPm/ird
QHlCB7+PpVH0tKG7ewjFwC86fG1sJ2bTWmgZPcubrWxWQSkQ5N/NYTJrWcNHFB2R
B0NdrUQIXRfns72WQt054bBAeyaf5y298tN63r3obUPFZ4a/9YavRGLcOYkl+sVO
XgUu1AxlcFiiRhUvx7EWD+Hb7aCnDYDKg7guFJpJkxs+T6DiiDRA6lG7RHMxyKxn
u4MB+hDztdB0lwCPxhuKbcQcUSJ1cx+Qz88WjrLGAqnP3JeGRXiNiGoBHs8xb48K
oeOGUhcowyfRcZLPPakbfAKwYoAtsfzl7/vNgQrqZ84pir/0w1jtyvyoerje1Ml+
s7uWowwDlHvnlzFk28HYzG0wGqeI7YRKp1bAs1tYGlvKRehkmx+MwoDWiFz7eJR0
c5yiETKinYpoKG3SX/qWQzIZADiMxfboG3bG+nwrZl44j0XoZ4y1zpzMP+ZpNVrr
KtOOaCONGU0aqTVHS99c10bI9Hr/eYw2K/KOfP8vcnX3DZSwBuas/fJj01hNBcpf
9emjG0IBUXYo2BBItrxw1+y20jvhUqLehnj8fMvEf+n1Wi8XW+0hjRG2AgFJJwlA
2SOWnVoKzolj4iqYOMbGMTrNjmej3excNLR8CZN2GUmqq2uYukZfznlO6c6VRTsV
15tOD3JNoXvN3xkuDm23G1j//Cr6uNmruO3JMs3HBmtjjWn3YxcDDmycyhXuTPD+
+91qJLRvQ9Qj4nQGNwqT+1ik4oIwAaz2rpSJihQUs4Z2bRsebg9kWk+mGAsFGN8v
TjFF75kgJgMOirohQHL6BTLIuDNTphTE+mj7w+RCFSNBE2X4T/uMH442GchGJvq3
4XmkiHPjiGUHb4DujVSvsIYhp1dt1C69+OqAKIBlc7clXHxYmxsWQVHiUYiM6bCd
zAHMaV+/5BhG+AdQi7upZisk+qhEVUVarmqqF4HmYuevvSGGDVQ1GZ6BF+Vp65Vb
WuFXTYK8tI3XJ/eSrCx6hqaWCWPRiKay+dZlsAhTwS91BPOI6hGeJs8c5NV/PTwh
22TJFwIY2XMZ2SuwHDdvV/oePjLqameTlVRzJ/56Lk7FpuriX7Q7gk2n7Tp6wQ4t
o3Cu9S3Rn4bjLzeNtpsTLszswUVMCB8lVPODtWKbpsz1dOgdTox1McsVov9mBm3X
AdjCy6XNTdi3fQcYU15NRsAPMc4D+OhJnF4OIMj5pX2SNAwaPXAKcSN+TWbcahUg
77df/dg/XmlqVqkBvKBGCqakOmzzDz1sNHlCpx6WylNeF5RHe7o9XmbYAjXEz/L3
kIoHwntNA+OtxjgJoubWgSYA8LyW88RsLnm8bNbEAUgFuYB+ZExTfmeqz1MstvR4
0lQmyNGcG52dfOJiP4K3cVxxFtu9C+/Up8H9EHpFaFpBTWWJG06l12Xgf/imaco2
poSm4uWT8/8a6HOgMI2Q+9AVQUfJ8PSMt6qzcJWUHvsLpyMrUH1n9AfhLyjRm9Qc
VMM++tTS//pNUgyDc3agmilVlDshzlYgOlcUsZ5pxCEJtM2AETsGyI/J6OxPAgaU
NhtGYnteIsAk5xmXTHrzdVZOfmsNvqWH642q3nmxQS4uS/KEgaMw9osVZcFQo8qD
4+F8UME7c7QOmuN3BMHV+sxAfk91FiLeW7Th1mEzgGZ8Cmhs/c/GqP1whaw+nkYC
y8D1JwZXswMLCeYZBA9Ii21bvSLmavrI+5eT2ElG9fr0FNtuXbozT8LVBVVeRyUF
CM4Hp+v3bG5M3oUOopMJe5VqD/XXf7o0JUr1nuv1W6p529KQ49U9knqgDOo5hUKe
ABdKYOnGdtqdb0/YO3KbLskeBouIQFtICfm2ep7M7kBwU+7lIMIFsBNqCtf6yUg1
qolyny+U6N91J64OAcriZRcfaEITIMS9r2rPCMkyqhl8hC+EHCmNLN3DAqIHbpQq
uAO2YbMMwgbnwS4ASd3PZwhy4wLPtyeyyR8lgGjA6Uk5MyPyxN1qAnR0Vj6qT7sm
Rc9ik7ETNY9ZXa98N2DH4THdpI4eyAgEyU96fuqHphwXYLHeFa3gDRFkWMrhZcM2
ZIgOqsEk+odaEKtwkApBdkzJ2YIKRJWB69a9EFh4NBb+Hy/xaJReg0uDc74QHdWM
Fb/ZkNdeXIgouHKPM+J5SsKmEMeQTo08tvmshkG1FjDfYJWyqth2dVNQKRdBcPHu
L2BOdopoyHY9Lqpjd6elqAkh4sv3Rgh9sQRSpRjiqUKP7Y0Xd8Kn+d8ZLhYbkqVi
gk/9BO5+JMFQKqlXaceqCPZ/8oORlufs2EYVFGtYbFZuwxX3+P7wi44rR4lNp1kN
uFos6Z42dSw89wuASBivnUKbv9Br7IlbOXKrFMR1ITAzzcopD9UjU+BcsSoLmc2j
9Gdjgb3Wvbw87zVLNOnJJVIrEquZQ0moUYanClbbGgvPIQFvDRb2+2s3q6jOpegQ
myFln6oS/sE6MjhDWzf/NOlM12JJjqglvpPDCYOhxyCiO9DKpMjLb+v25VJRz5J3
1J958eQzMAasmn9DGWasn34q8yJ9zswMUlmPheAYGWjyGtODXjJ18z9saiKlv0Sb
4tKgqPtdc+2ORRBNBOFFZYLcLFbBypRxuC1mXVz5hO6msfGlvs2k9kdREHhqqOIK
uqJVYlj4flaHS19ZVzYqU4HJMuAAyHzKLGiumj9FwlLLfMFl/oe7CWorf154xCe1
jLxGdTo/VYmD/SlVVK274MElh0ugfRTmREyyxmczmHYl8RnBjm+c+v0D3Kb5RqGd
rFeIAZC3qxeJnCQC99YQj43OxORzQeDSiQkXMtvLhNeHJr8Pz/Ypime40LfH/JAD
fNpyu0HfeUIuaRkfuCyH0urX9/27xOhh1n90FRaI+DwykzsJGtWSz/ymPXJMn6jd
ywXjBxH0XPzLInUoQCWzZfnA2SokK7M+FBrKVqFVGExZ4ZBGYZwCqVCjfNffLMul
aWQMFnLATpZjjKvA3JfkAqUcBgJlBPcjyT3w0DvoP+jQr74x52V9/v3rhCYA0xh4
3u38lH5AePprwE63IeIFgUntVcpetPTFx3z+epjdHLkDay5RQI00yonlQ11fZ8qU
rDbaEy5PdBysU+KQUgR9J88NuL4Mu+hDQo+xDhrFjwdGgnpo2eZ67pUMzonmwmwj
XzEeYHRb26QX58FI+ebNgba0rUdGIeUHOrutGjxKMMRCitqyVOEOe1bZaaDxvpt6
NL8PcBLue4172AipIy/UagMG2HVOECcm2JaboP+RG1ABhg0HGiCziRJN6Elmc50D
hNcjb1a7c3MLC5XgwzBVbFvB2qayCgQVYBruaR/i+gTOGOvy5E1jS3w/v4JRBzmi
wBIx0PKm4M+njvlmF8/W3l840tRkENpCQoZBi1/K7BoKh9KeE96VXiLBRTy+GJEz
SjSJ2dCC+mOy3zR18Ci8QUJIjTVnICqBIZKv8eEgs7ae/CtWPMLneo9gcbKsDhjX
TIqGNmYM0iYE8Q8ofoXamjoqwFfRCNyjcdDhlOZITjag96A6LEUHS021973fV82K
GYxYwtPviI8N0JSnmtsB3nL5Yvw6vxhuKwQBSLOnJmnuz1WgwQIrZjaKnMU3sbeL
jQNUueJsTgGj4TqNLGnvdIJjisvyXehHaaPpvy8fGR9bBipaW7MYn34cFezP/Noh
oL/953ZmJ2b3Gx/YpDeqFICKhv2CPPaLDjfwY1UAeXcoMIZbZCu5vGhZt6q9XoU5
skq5MW//T6RKVq9spTIPqsKBvkfIeoB3OD4JZ0ALBerqctOwqyVkxGT+8gmxHqeY
HuJ6uAfknKRQaWPOUzn6F9cO7QfXyq50BZZFyqV350LTX8nOhMH5tjuZwbo34sps
R8zjImiPlkGd3UOqRcw+Nd9+1bdmltXqMDPOF6MXbovLdgag7DUhOG2302CPOc48
nu3+VR2KcLDy56/7cHj2JwPiHU3PkPPp8QBfix5evwpAEibjG+SXHIpvr1R6tnnu
4qOzMSStmw108T2ZaYxgiCvBWSX8Lk2+33v1sAy0/2T557C0uwfuus+fGjbBYkxg
v6q1iwSbiLnF1myHwKEb4eXMdResxIC/IGbPeqogmzg5EffanHqtI/5IeS4StMQE
CirDa/OrMuuRKmFBrrE8uoRL6VJkIwKRedQTNirI/UKkSQ7nbAZ7h9jxc1Y20er2
85XVfWgWkpE+ttqfGcT5BhoAfr8UjYwb2zdSySDmwbgYYpCeYGkGXOQMNqnrPLnM
lg0y13z+Kidl2EbTeff5nWSfVmm2tXTHf9s5KX6cdtpJqEL6WjLaUGe2c0v7RiwO
sbN65gORUwMcXSPpDT1wWOZMRAdNyRf975U7H4JFYXk/6KgNzvsz3rvRdOWEYxUj
CbUYrle+w62k92z6LCmhRGQKShVkXwx8JRAV9cDKvSh9ibuTkMU4YhAm10SFBbxn
60LYmvb2BwUowOtSTbhAG/hMkd1BLg4qPxskVoE1/Cv8P35QcaHgsT2MdAAjoU6Y
12ma+BcKmY+p2LKTOa+aQjN5mBA64C/VcR1OZ6TElu9COo9Ryr2sAQZG1EEAOosM
4CgOQrlCPnQYBRvpEymPAAZQyzh+vt3Od1vmNS1JHhfnSA07Ik3seGQBRqaifbeB
34d/XcHruZh6d3XV2DtIkrZbCopGmA4mbVVO4wSJN5G58u5IVvf0PX5tR94bdSys
Q2cUBmoZv1XWPsH8yNyb6l8jJDeb9kvCtKBgL5c21/9GefKElTGwhJcDqElStz2S
x8sOApLJL1/Hc3xZoU8rp3+zlWgr2pvFoIwCsgTxzEeboyNncMEPTiEOjX+PayOn
hbgb7Y9f/CP4JpXUTKs4VE2u71iVranPUG1yFRv37b09/DpZM91yAzSVEDzNzKb/
zkrQ2WTaVToGggaynA6ng/zBqU0MQ3b8zr/upZrPmsvwNUIbp3QbhSimf2fdY204
IV9UGKpMi5NUlrUBH3gemhdRxAUE3XjNicfjdb+r20tbf52ipC3eZu30wOvZZ2dO
k6TXOz1KxhiLVWaAkWkU080YonoPhpH/LBcupVMFuMaj7RW4BjeUbFoRwDKGJJr4
I9yRJeCKGNBcAixdkG6Q8xfvs9C2/SQ7qH/7c8PiTuOLEIflouEF4EiaRsLqRvlK
BQOVV5j+BW1QHu9CpC9iL1gMV9NC2YI+BkNm9ZJBy3SnaaLCWjuA6FT0FjuJz2zi
1VUTOHtvHszPIOwhynKpLBewlmjBBjusaerpyox+gjRnE4dwbRcV5X57svcVUMbs
5qKvlUKSPMMTkRAGD/7U6HiuwzRVDEOHMuL+VXuTI2cMQwhogNpmWaI2gczkWm+z
2yQ3a+cDD4/1N6ZVz54/+LqhiPhPKf6PFzlkS/1pVF4w/VT+QE8KvIHO557HI1yS
bgwbcsIusCkLDYJAqIjUDd8c+jZQwwWK73F9v9Uugs8ZjKWfboEppJUQgkNkI5i+
GvbsiZcQA2dRTTbS8ABlLeGE4m0ypO91zP5xyFQ3So4F54N542n29oo+w+NnmD5M
znkvRVPa9RVsDcN59XCgasZzjXDR0KPYmrM1/cdrhracRav6rEHpCNEt1+Vl0VhL
p2OkzOBCWGMRioGeABa1lTXQr1y1SD4A8b8736Ela0agOwvZpRkLEBwZjFGxWcwQ
dO/ahjTC6LYz2Mu+1k7/5SGLD4thKN/ogFrJCLZtIGbhFBXZVZ9tPz4zbqOgeEPe
5lsDdt9KuuP6mwIqJ4DMsgON8+cPTppJzmCpZCv8dGafs+hsKZhF/yh5mMYhUobV
NUBjeK0TazmihHSC1JWz/wp4UhIYJr5k1DnyAhMPV+0ATPyt1RNFun0X5vMQtMIx
6Xhljfy7pvFw17Ua3JhG5lpMIIoE/pWX1jLIJrnBVn1epD89eiE2ReF2dk/Uz1QL
ccKumEM0enoqhBhdRTS1nXMlTsfk9Xn0I7ZJzUGhnaY4fbGLfhBHw+rQ2e1KRjXX
TPwnWDg+kmlF+U5hJxq8DJelP+0pTNGS2BfU3gdB+pOhk30oECEgN2CVlVp2xdZI
QrNomvGlT0Lwql5/aGEIWfWe02HmJ23uMNDYdGaHEDiecj80a1xbh3GEbkd+5nII
aKiPpThIlkrlaksdDsy7PHvUEokRcAScnW6/oTj3urqTaOsPoOWb6ObN2b9N0h8t
e24NazHCO4y8+lgmHzVCM7xhhgpcE1F6sA6IdhWv0+TS3SsGcEw3QHvbSEhL5/kr
eEA6nSvQRZxV+dQ4uHJ4xHJVE/c4oj3CDTMVulyM3AQ2O6dSV29Lmx0LkBoR0/7H
92b9paVOBF513U+CqickaXBNjSXmjX4MLPgm2Tb/C4K0WraGDjEi2rr2fe5SKdr4
YfIQanEsceAaezq8DP/BbtJO9zB2jFJahcR+E5UdkoTnXkq5PUZndw4Oqyr/7H7n
MzthC2LZD9H99jGjJQSe8daR7bT8ZGT7yl4ypqD5d9pXnm5rywc3hfHQyBcChd99
ys3wTlNnpO8UWW3c4+Ah3vthbJYcspm4MQk65G0ub/6VEaFE0EB0lx4ONChWgt9d
84g8JR3SOZ5fxD8oP3CaOUnv/iBBJLZ8Rto2JnhJwlUiXzEMTv4X0YWHKnXIu+fi
9vt18Vat5rd/YmxBUkHIhWyBnD9GyFHeN4PeEHp3ojY5nZjMYCHERAdzx26HdRqs
eC69QY2RBJUf3L/0ohwbwH7UL9S/MHf+dsbvoH/G35QAXghQb06U9oG0CJQatlA6
zWH+VJ3YXvtB0UaZQfWy/KbVc9hE8xkG04igkvlFaHbRjByA+2Y4kH6jIjc9byRz
n53w/QaeF+NmSjnNjwrP/O8NTgivxM+rTwWeVI5RC822WNohLxxdPGMLuh9TgdeW
FBAl435OKd+IU5FPjv1VbuSVzShldDJZQ8XxcKg85N47O9RxcoCUVO4umCuQ0ztf
Ae1nqBfroq/vNEhm+qkQkbCnJVf9i0z7o+qbL1+ia/puoG/fsghXopl6w/dXuWPV
xfvk45+U/p6PbxQgrkbVt5dd2eB7J7K/ysfeHhdp0qcNPyJjROPt/dDYfW864HXN
no+xuMvWM1Kh3h4TySrvrh7lzps7vQb4yAwLgxqXynbbepuTZuUIBnzLWnuJgfjU
SXLkP9BUX4nlYckNleRQqfJRUnAGVfwxJokQhTVNBQ3zFvqzzFLiQSl3NIem/Xhc
TJqFlsh/QzBecpEhTvEjH/6U84+4bQXBEp8q8SoZ5mDJerpssbl6hY/E1xRdySW5
1gkyjJf/+mmomC19UC+P9WuOg7tg7TH2Y/n8Pei8tS4RMifsszvYCBhMMTzwSET+
zB6B8cRWPPzqG012oPC1eD1LnbQcmyVgWfs4Jr0b19foG/m8H4L+J7ACS+CIaSQ+
ax0yZYOxvn0oZVB9B8wg2grp8odVHSn4y1aF6QB/ola8c1mcWHqC4wxfgD/lJfd8
d6uSwJD2/Eo9TRtGopa1i9BwbpFiaxEfzb+MPZisUO5G0ujFASxVHPlcNqaLf9mc
Uvjx+smkWtpN/f5XwDj+fftupe2M2lVJ4CNODd3ZbY6o1KT3JzBa0G463cFMYJB4
b7tv4dujVpMTG4DT+7mlQbfmZDBGlAO14bUdrwppYA9XqOv0aF271JPwOwp6QVTd
FKAei68egXaAW6eorVfVX4smvhlz5Rdv4uGZWuwwqHKPFMK7DBRWYRaHjM3S3L8q
GuIdiB00zZzodyrDWfzIvvwYCZHjTj3Kw9iwrHTusQ4ElSjxQL6faOakN66x3bKk
cER7VY+driXElyn/f0l9XG1wuZJdqSeoGONC8dCvt1IkrL2dekMF+CadOoeyXUpx
Tnm4je17xTEcLKhaew6QG48pZHiZTqYXBU1h1yHBOkzdFrUZZqlcbsFbWa91kOF4
hMFz2Ta3y6PXdIU6OEu/lYKciO3QNcbKWJ7rBtOxd8/zA0/CbhzJHPlY8BpnPZd2
pDohd97SJfizM3NwHmHvgs5pGc7HstnWsKgpaQTdsdA0K0LsRxsKXlra0stMja6S
S3TAu3Orjtlayg2UECyCEj1P50TgzcGrb2boOyKNLukkXf3DkNpYc+gdA/A7oEN5
l7cxhfHbfCOBAMz3MLOKZDv3jswxnkIE2SAHmQqyGwlIG8zw5qVaqYNpILfsIdq1
HmyCD5GxfCs449xXnFIHj365HOGxmwfe7fcCf5io980xdUzJiUgzsf7WOf3tp8w6
b5hzc/oLPFCorJOR+bUxYLFRPDf/G0EBqjXA0r5Rc2644CPo9eU0iDRJ1+NwVKyg
1XCN+tU5DFqzRYIBT0Ia8aMMqONiFVaizEhrJUgsHDiP1ZE0VMkdmsgYBH/tkNXr
eLgxHzaW+gayxCHN8LTuHFe3DT05ilUeWeWvoJpUxX4TqS8w8NTWWa4sloUrnDg9
Zoxs2bVMsCq3Af3P4ASgTxTaV9D/J47qKxtnH4kxec8YRLJ/zGUleZ16SPf7KvrG
BmlkpmptBvQiqNCA4fbM65YYM5P+k8GG8sAxHj3Kma8n9ecXx3/AqcWs32dySx4I
QS0O2Tg20m+yLs+82Chhn1nw8lAE0aIPnTMDCKVI9ZKeiwuB2/cLD/5wsFq0RnBU
vLtGRtTYBY01EPHBQgUXAothyTxANTwISnAbpA3WZ2X7MVPTde2Tus5IMEBs2cHk
Mwdk/VhYuDoJo0+gm508l3lSzkblbx2HdPsSFZTMwEh5SSaicLWngpKEY09xjqZK
he929ohREmc7Iq7U/SSFYNg2tSkDWGaLng0HeFSI3YtMjxA+WtoKmyfO9o+RNTkl
fNByhHepdjk814YLrIiUI3xwhuLuiwEH5f0I49OI20+EAiPtWmtURWmlAnXs0kNw
lR5UxkoEwCoOwGgcR4ZbK0L1FIyhJFVXzFg7LuKw0KaVeSKmgRF6XCAg+CyX+C0T
KodT9RkjABEh0JgGsAW9sRDfd+QF5zS//HsH/Jt2GUDXd184rBf8XYKuG5MAAzGo
dhFaCFGgGtTcZOQAeSHYtdVHjRw5K2DWfItOf9WJajzBQeunHH8e9F93AlqhirCR
EtvNEUSKau1ZPdAkYsnonTXy7OxUqpRo8rFPBSO18hjU56bDZj9zGWBbkZcOfyEb
iO2Rcy2lkMYYcEpedw/us4G3UnOtx3l75mkrS29vF0Bq+KDmKuwKkkLi17RgXLDa
LZf2+tMQ3clLoihUoCBFYIC/bKV0ZdqFE028VhWIv/3tGC3f3voYGHehyHM0+nMD
R+L7apAX6AlcfNwIN8g6FHJl2UxNACHeR7LQiOT5V4kY81sQIrx/cUSvxGTv3hqG
DDx4L/5iMkp/eFHo8RxemrrysZNdHYSuTXO1J8ULW3zFf8QJQUpJ8MwUq4XyXJkn
zoD0n+Mqqnvl685rXHZKqpFEK1c3bA7VitBgkzIU3mNJHNyMlLYqLejs3TP/eAkr
V92js6iLXhZrePlQsnw6JdN/ugPv7WZ80Lb6k7FVSrb4Ifr+hgB2CB4708cK4A7j
8Q8ATCsXADbvqKfk2IfLP/BTorl/93Zs8M4TuRWcPx+ozOCwSRKvvKbHEPwL5zmO
aLAxfezvKxCgpjfUeTAEvadR2VZexnahPLg6rxnIYvGMTWlrRT+obIIGacLUqJyU
4+xgtlwk2XmuuObsU25q4NG3q0QoXi/1bMNgEnU5M84fyYWZK4JS7xCdpOhqyAP3
eE1RKZj+nAqHVIhUFAsxRbm79hu1qPjxatdADXwE107qjn+alCg8ykQd/H6KShla
Nxc6XWW1+YngACLWPQzfZTKqV62CrRgy24nqLykqXjlLioq5FuDTh3TiM2wgAi2q
WSfJb8YyDEge09Hvx/CMuQ9nwB6LutKl/inip2RrEu/2UictyQ0r9hN5R+qKSOGb
2LCkRuouX+WQ4aEcO0hm8ltze7LSddbLZgzX9SoQCVUs/Wi/KCskOOIpJYGoOg1J
+npMUG7U+q+tyh/0iLo7q2roA0ahiZPxZWSz89EBLyL50drrhRWcCJJ5zoP4iObs
z1G0l1yViUMLCRdhqh8KBRfLy+HS1nk4ylUbpG9S788CGY3TLETLrlWXTDYoYojL
DYrgWvOfT3ZQV/Dgl5wGBZYrogrmcjkhgNw2Vb8NJ3fqj9l7TkRDPg8kg8eLfDdz
Qv/N7iz7Gj1VYwc6vj7kfV8jgsuEugJIPkJNt9sgTUGe3WZGv0s0fMg9suRVIGMG
voYkFvs43b70PlGuBTgoxeBWXKG6/feriy6FuedXKoX6GuVZPXX5gS6vIqSX27qV
uYShsET87khFQDflrJt2Ecw5PEl/UVGIC7RFxgyXWA1nHftWHkIu5abdr8x9hhC/
NEZG2j5/SXb6E+gbn3GVjl0k9M7bzZZUMFMXA6Bmbh1vnINbt8N5TPBkSzaiJuRx
2Y4STiHoSIDZrCy8Arn1RYf5VmfeMHNAhF/LZA/VqVBraLrg1KPxjH560K8SGaJX
jbTbqIguUn0kyybtMoMD3cY85GEKT1M70+up1z583F+xrl9E20GBKTQM2jycMwFe
KuMDyU8AaWOLhUERpnl/RRsmcimJMFCQp8XrZVhm60DSoUXimvAZjcVy8jnE8EDe
cv/JNrTQjcuY0EIrkFNvquwlhJyhSoxN8Yl9qdUUqn1Ej901Yk7ka7XlAKyU1bFT
QqwRqs5m+Y69MiWSkR/uCntCiuL2NCRTlPKHMCwjcNzIIZP39os7r0SgL2nbeSKJ
jU1whp0ph08FYUIjJYcRHGp+RMwd4DU0U9XX2bgxj+CrAhlbZdSaUEhj/ZIttZrx
80j0H0rq+mu5gpvImH261IkVzGc8EAHhiKhveGV5D6Ii9uqCeSV4/G/FEWN/WakO
SS4L4scJnOml0ihioNuNVnPXGSd4knRWttgLL9BPPzHNSyzVvR343p9SWkBO1ZRN
UmJ4klaAxkxv0CcT2NljcEw1w+R0+ekP+lthXZ0HBo0pOr7Fx5cNzu2i7Rql1Kdb
jJSxhU6nSHjNET/VzMsF9+ZK5cIpxAU+FQv2Sq7E0spUkTQlnqIpZbQf1+D38cPe
+8sYqkAQ7SHe8EivV0Z1I4WE2ryWa/Vk97ZpQ0CFF00/cRlHSn6rBgVtyI8BX59+
wbie+v+4lZbmWtH95wqnaAqBaw/hYxsOATyWGwy/zgjvsFi+hicLKx0lYIsng0gI
hSBjg0D88JsDY4AaMcSzOo66sjXnyXh55M1kZ7cbSc/U8QbLsVbs+xRAII7roXKW
kEVARXYXrZC8N6VwkU1PLMH1wl5uW/3zGtfgVZe+B2BRBimeUm+W/Hc7pqMKJkAG
fL8GRFDpgTQypUZYrJEVh68VNP4StNmh4oSjG3rt0ivgNnvgbE0lh44HrlS9PAQb
DNp480P6MGGMhuXmcMQgeeIkS+PjHk2qKzP7yD2ZpvS06dT2T+TTI9AjtWZ5TZMt
I1YKeiAm/g4dtsbsIrBSfGC1QAREo4yEdF3oU/OF9UhEKJVBdcejJw8d4NO0hDzI
klDo5YcUrXTLsfRNeXxLl36STQr4ihHL3yfpT9yZn0q6SgKRkbrtUv8R3k6779nz
ipSPIxNYiigqzHYdwxp/Tx/a/OSSfOSVzrg6ynaDuyFaoBCHZwipSGVZ7pAm1dZo
3b/KutAKQbOAqABEhQnHe4YszXqzZKzcTFz0vT2Nw03Ek5iBz2pogV0jy9Lex0FO
GqWDy5zGqGSbgvayXd2FkD7kXZ1iTqVb9CJUNGq+y+I2TnSwX7gGBnoerVsqlz++
P+seu0U6qfItNug/I9PgcS/wdeYjgbbx905Z2ccGypC03B/9T6e3X4equm3NrLfS
lv6YnUa4n5+Li6GVSWXm1+8FRDhGNXs22azx0Ch3s+PG86Bf3RQvQsVr62jDIE5V
4QWDz2AwKUJVYHHoq5FNhifN7Wd8F4ET9DaC+2kPbmqu6UgvwQMWZKAHDtF7QhhU
o/7Vz3UkA8gYVmp60E4I+m4MQSdy9sNK2/4INocPcdzkLPw1SlIkpnD25+55fz7n
gfZP4OBrBOY4aa2KC2jrAY8LUXCLoR6bqF2KXEhUDYvjTNJdugwq0wkAXU54uCFO
hkGyfh8htPgVQhymDwKBLKMs9hwWNlECEzvdRC9s4nHnZtH6U8aQuwpgYEmPAo34
HlJrARi42QN+KwbQtyXPVjziGahQpWoPpfyt/zv3gJ7fSVnr1nvSgxqSX6AWf1dT
W+XdIiXMjmVcvQvXJ5iwFhyNRSwXGG2cAwtoyHNCWHINnK0xIXnJhmkZube4Qnxg
PTpT3RqmX3OobpTjk/bgpKZEsnDZg9j5YykJjt0LsdTgOdGuTed9rN6Vw3WbOyb6
VE/GvyvL4SFp96NZX/47eTBLA+H5PpTFvpkli7DKNrXP9MCHOKxl9GqpNcMYp9a3
XxCGpqBcKKORPhwO+JzcTweyT1UhtuHzAWhQDvJ/LCuOVHhw+VUzLIks4GTNUwSq
hym88k9gyovJ+26ZtcTHPf/9jNUifgq3GWX4XKwlKOtMQB0k7S1algH4WfNgD3CS
As0UwCudAwNU1Od5R3mvTWLg772GdddcNsLGSd7QU1v3JlR+3oIxkMvXk7ie3DbF
UFPWkx8A8R0KA8ZpAiE1nnY9pO0AInyl6nBIZdH1bjiip+AWQz5LkiXfW93dzT/5
h8ZTP8Xc3DHKSQvVolxPygKumOiZ3WEN/UA/z/vo+H8IkEkT7t0wXs6I3gCI9Khq
+3Cf/RWn7Wtt49PThBjMX61CxtZk5mnj1UiOIZGYPgwUzAavvw+61i3ljtrA79AQ
rJEZZWMgx6FGf8wTq5PsLAUaKpAkU3a08pkChWhbY8BQMK4UUZ9Ic466Et/+3IUF
KBntPbrIa9j4FpO/OKH7LqHRMaKu3t8Gf5pP7ZSNe7mZxQuWsM6WhaCi+MREHV1C
2YL98cixvVziQUPBq7/y5ww6GRWe2kmdx1SPcHW2aczqyR6uBVPtP9/6H5Zo/8yF
wzB5sGNIbRVkKFG7eqeZp++GsxLEjbEdRbCoaUXBzfCWssSy0KzyVcWH1VUXcEL4
IJtd5QQdJ/k6sMttfxrnyZ4TiK85q8c7+0rcX/IYA9Kmjs0DZiV4Lx0VYSZ5aK0r
+75yOVr/K2FdJ5bEZLMXjPBp0bMUw7Y5EH0a6m19mPrfXoAH35gS8i/gvRXx08V/
PEOizAlTWilonKrIA0AbXkxH9vcwccBqfLE3iZk0ZPSrrV+r5m6Fmfg0/J2RW35U
YuhCaUWUcWHC4YWs2uVslUgYvyZQxNChGujdHR6mAS3cNAHvCjTUq1LGN2os4Vie
Id85Uvs6FJA2hXAqprnKe/aw6SRHFnaIrO84fVVsdm9GQ7UuJcEURpB3uvO8krJa
nQ4ucHnzjsDw6pPh9rd82xMnMKJDA3QNugcIH67uCAi/PXCdazBMGVuAwh5kukK4
3e7xqr4a7ctKiuAGbJ3yOluKq5jSqNLIe41L96UARdHXpQhj44w8ybhuRIdDb5Fx
21MaC47Y4Y0j3W0QbLXk5Tj6YjpELYcr7y6Io7wAW64mUXLNmbt0qkFbPHyP/DPW
V96tFI5lkLfzD4/5nDByD9HNMJ01wXjGRj5rNwbVhKtYTHWBVJfYGr01RsE+cMlu
fh6nCO0sSCFyUW/0kcTnlUSzCQKxmp2K2SAsN9MwcLX82BSpQ5N3AWOy5YVAMJ5G
LElvuN5Fl+rnkNUDy4L76dXSIcbhadiLz7CzMjBSuGiG/YAG2LiYbsniNx3nMtSh
CabZ49DrZ1IDLsJVSUa8lentUwrI/1lXjs1vST4sd161cYw348NGLdWsaO5uZ47d
emBIvIAGh6pvpWtNNqGyBXxLgLUZise658OsPbm2DvniKhfm2gWWuEK7L82uJ3uw
cbLWkQzSQ0+8KUJ0/R+uZaWHwKt52cN2YA8rfn5xnA4HRXDBBGFyjwlGNNBG2EuY
ikUr920j8DHYmAw7cAQzZjBLPvylValX+NUITX+DqFgCzHDeIaJzTNz8BrG/7ECY
ucpdJGMqPLIuU2VXetBl6xK4qF6Fg7PQhapoqEZ2tauiVCbJzslkNDf94uicq4qD
hLKDzpJ87Lfci6nfVqJPEaC+ILvFttNL3aTam4kgkRIHLUEPmb5qC817w7rGS5PP
yQLwq8BTeBwKWmzVVxUkisx9uXTtX2dbNoS2uqdRzFv/4C/hQfgFAMsF8cXT0IEE
NN7R3HFsxBYGaCKEt1MURcisqLebVKdyOs5YytXz4jdMx2P7b/KFhyYQSLZJLQsP
iNqGWfA+0KRYUuLlsVkR/8T5iKCB7ADHyXuJvEIewGJ5S/207oL4SY7o3Zco9RqT
fvOB3BHEmeV13LVgKz2Q0hdh3xMhzz+NYf7TU2bFj7SAXALtGy3PI4rKmPkkcK1u
m2j1z0LdVVLZkQXurEUBxf7cFKOu6Cce2eY448lBnTqweaFkSLxTDSEVn2gAbGMY
X6fkqzMaRegXLyuY3Z9QRYc3S5GiNih89eOuWKF/RdWz7GFYprvlbRUDrOGRjmxM
f5KX7tPA6oDcDwN+oTzrg0HQw1GL9WryCmgvAHiVQPpTjKXccFNW70wzO1NW5a3F
jbTQHQfAeRzF35rtd7X39Q==
`pragma protect end_protected
