// ed_synth_tg_0.v

// Generated using ACDS version 17.0 290

`timescale 1 ps / 1 ps
module ed_synth_tg_0 (
		input  wire         amm_ready_0,           //       ctrl_amm_0.waitrequest_n
		output wire         amm_read_0,            //                 .read
		output wire         amm_write_0,           //                 .write
		output wire [31:0]  amm_address_0,         //                 .address
		input  wire [575:0] amm_readdata_0,        //                 .readdata
		output wire [575:0] amm_writedata_0,       //                 .writedata
		output wire [6:0]   amm_burstcount_0,      //                 .burstcount
		output wire [63:0]  amm_byteenable_0,      //                 .byteenable
		input  wire         amm_readdatavalid_0,   //                 .readdatavalid
		input  wire         emif_usr_clk,          //     emif_usr_clk.clk
		input  wire         emif_usr_reset_n,      // emif_usr_reset_n.reset_n
                output logic [3:0]  fsm_state,
		output wire         traffic_gen_pass_0,    //      tg_status_0.traffic_gen_pass
		output wire         traffic_gen_fail_0,    //                 .traffic_gen_fail
		output wire         traffic_gen_timeout_0  //                 .traffic_gen_timeout
	);

	altera_emif_avl_tg_top #(
		.PROTOCOL_ENUM                      ("PROTOCOL_DDR4"),
		.PHY_PING_PONG_EN                   (0),
		.MEGAFUNC_DEVICE_FAMILY             ("ARRIA 10"),
		.NUM_OF_CTRL_PORTS                  (1),
		.SEPARATE_READ_WRITE_IFS            (0),
		.GENERATE_LOCAL_RESET_SYNC          (1),
		.CTRL_AVL_PROTOCOL_ENUM             ("CTRL_AVL_PROTOCOL_MM"),
		.USE_AVL_BYTEEN                     (0),
		.AMM_WORD_ADDRESS_WIDTH             (26),
		.AMM_WORD_ADDRESS_DIVISIBLE_BY      (1),
		.AMM_BURST_COUNT_DIVISIBLE_BY       (1),
		.USE_SIMPLE_TG                      (0),
		.TEST_DURATION                      ("SHORT"),
		.PORT_CTRL_AMM_ADDRESS_WIDTH        (32),
		.PORT_CTRL_AMM_RDATA_WIDTH          (576),
		.PORT_CTRL_AMM_WDATA_WIDTH          (576),
		.PORT_CTRL_AMM_BCOUNT_WIDTH         (7),
		.PORT_CTRL_AMM_BYTEEN_WIDTH         (64),
		.PORT_CTRL_MMR_MASTER_ADDRESS_WIDTH (10),
		.PORT_CTRL_MMR_MASTER_RDATA_WIDTH   (32),
		.PORT_CTRL_MMR_MASTER_WDATA_WIDTH   (32),
		.PORT_CTRL_MMR_MASTER_BCOUNT_WIDTH  (2)
	) tg_0 (
		.emif_usr_reset_n                (emif_usr_reset_n),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      // emif_usr_reset_n.reset_n
		.emif_usr_clk                    (emif_usr_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //     emif_usr_clk.clk
		.amm_ready_0                     (amm_ready_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       ctrl_amm_0.waitrequest_n
		.amm_read_0                      (amm_read_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                 .read
		.amm_write_0                     (amm_write_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                 .write
		.amm_address_0                   (amm_address_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                 .address
		.amm_readdata_0                  (amm_readdata_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                 .readdata
		.amm_writedata_0                 (amm_writedata_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                 .writedata
		.amm_burstcount_0                (amm_burstcount_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                 .burstcount
		.amm_byteenable_0                (amm_byteenable_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                 .byteenable
		.amm_readdatavalid_0             (amm_readdatavalid_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                 .readdatavalid
		.traffic_gen_pass_0              (traffic_gen_pass_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //      tg_status_0.traffic_gen_pass
                .fsm_state                       (fsm_state),
		.traffic_gen_fail_0              (traffic_gen_fail_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                 .traffic_gen_fail
		.traffic_gen_timeout_0           (traffic_gen_timeout_0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                 .traffic_gen_timeout
		.amm_beginbursttransfer_0        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_beginbursttransfer_1        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_beginbursttransfer_2        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_beginbursttransfer_3        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_beginbursttransfer_4        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_beginbursttransfer_5        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_beginbursttransfer_6        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_beginbursttransfer_7        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.emif_usr_reset_n_sec            (1'b1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.emif_usr_clk_sec                (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_ready_1                     (1'b1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_read_1                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_write_1                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_address_1                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdata_1                  (576'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //      (terminated)
		.amm_writedata_1                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_burstcount_1                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_byteenable_1                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdatavalid_1             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_ready_2                     (1'b1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_read_2                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_write_2                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_address_2                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdata_2                  (576'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //      (terminated)
		.amm_writedata_2                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_burstcount_2                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_byteenable_2                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdatavalid_2             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_ready_3                     (1'b1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_read_3                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_write_3                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_address_3                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdata_3                  (576'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //      (terminated)
		.amm_writedata_3                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_burstcount_3                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_byteenable_3                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdatavalid_3             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_ready_4                     (1'b1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_read_4                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_write_4                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_address_4                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdata_4                  (576'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //      (terminated)
		.amm_writedata_4                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_burstcount_4                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_byteenable_4                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdatavalid_4             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_ready_5                     (1'b1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_read_5                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_write_5                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_address_5                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdata_5                  (576'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //      (terminated)
		.amm_writedata_5                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_burstcount_5                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_byteenable_5                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdatavalid_5             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_ready_6                     (1'b1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_read_6                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_write_6                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_address_6                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdata_6                  (576'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //      (terminated)
		.amm_writedata_6                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_burstcount_6                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_byteenable_6                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdatavalid_6             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_ready_7                     (1'b1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.amm_read_7                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_write_7                     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_address_7                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdata_7                  (576'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //      (terminated)
		.amm_writedata_7                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_burstcount_7                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_byteenable_7                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.amm_readdatavalid_7             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.traffic_gen_pass_1              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_fail_1              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_timeout_1           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_pass_2              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_fail_2              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_timeout_2           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_pass_3              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_fail_3              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_timeout_3           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_pass_4              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_fail_4              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_timeout_4           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_pass_5              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_fail_5              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_timeout_5           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_pass_6              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_fail_6              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_timeout_6           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_pass_7              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_fail_7              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.traffic_gen_timeout_7           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.ctrl_user_priority_hi_0         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.ctrl_user_priority_hi_1         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.ctrl_auto_precharge_req_0       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.ctrl_auto_precharge_req_1       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.ctrl_ecc_user_interrupt_0       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.ctrl_ecc_user_interrupt_1       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.mmr_master_waitrequest_0        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.mmr_master_read_0               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_write_0              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_address_0            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_readdata_0           (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.mmr_master_writedata_0          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_burstcount_0         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_beginbursttransfer_0 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_readdatavalid_0      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.mmr_master_waitrequest_1        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.mmr_master_read_1               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_write_1              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_address_1            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_readdata_1           (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //      (terminated)
		.mmr_master_writedata_1          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_burstcount_1         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_beginbursttransfer_1 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //      (terminated)
		.mmr_master_readdatavalid_1      (1'b0)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //      (terminated)
	);

endmodule
