`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
roq4UVfIJ2gLynm9XgN/spygvmAi/tjCYdc0U4PGkhs+h+5uFnJkTqm94nbxw8f5
YJeEijJ8iY9N2RD2zHusbhQtB6uhWS0rfARDoqSSvVyH6oaIeS/qHmujbwain6Kj
oWO+HX9/haxTwFuCZMoSKAb+7FRvMLhdArMFG276tfQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2992), data_block
jIHaNCvGrHfL2EFncbly4WvpZsljYhn/AoGPmSCWjzxjJbDTeuFYUb9HT7WRq0oK
FMWhEAI9lMewQEfgtQu8AzcRJp/JoEBvUb6oQjwFj2EBEHQRXNOLTr0TvL79Yxgw
mvg19ec3E+QOI0NukfETPlSafd8Dwgv9GPwGN2xICGspEite+f9ZBAJpedkwM2FB
Xw1LYamThtpOhoyhC/zJdsyWSc6mqGgxx9S1IMuBN8eJRwdVWPERZjsX0XdX9ywg
6TP0XhC/FO4AgBPay+7EL6bOnkaPqvRtymAgfMP+XCqJwy4bLWAJNhnZeb3jTCdo
KM+KMRxx9r2N1cdIzeU6ucO+wlrTIu3cWy8WDMfDS+rRqzuo9Mzpvo//7OeKlpYT
rmBjC8l/J+gcATvIX/JMlmWDNqRlYmHE93gZAUCb1BYlI8zoay77A+zJDC39oYi5
VdpgMgop98dOgRl/5t2sb4F0xu8YJFDCTsOFHvxu7UsW5oFTVLrmZBWcNlVvIVSh
n70WyKtmZ7LN/Vf/ugMufZiVkb+ULn8Bv6qDOzqGBv4qarkmqRZVRHeyNnPhs76p
3MnNNrq7Kdd/izHi59xpDGSyxiA2Rtgr6ryy7pAx8tEiurhoMTXlFuqt9vSXq2QL
VqT5K7NQ+1UqqhPNTvFtlzzZmj+QBpZqn4WmoMS8dYBXY0jhWsIwehiVkTsWf/1+
NR3V9dTEl8veapwHk7gTGdcmV1i2HXHTgP3e5MPhCHeGD/qSsBwxXMGNyeR2bXem
ZG/hBQ9p5iIQC561jR828SZPtiJwn2HhIZRzIvZxmeCgs/E7Oi5iS/+qtw7ZTIOX
YVwvvlvzFTiMaZyV8jH9py+vAZoonrH7bsz7pSwwztaihWh0fONb5DjZ0hRj/qml
8p+BJBnE+E8ata6nvo2vl9iNQW3V2cKS0D4rwpm3LIMM9GVG+pu4WxX4DLljziGS
v5phu95MKvgx/9TNpYRqVdY2j5AIed/VJkmdzmGPXT0BRsNMXhaK6a1A8EMNvSY6
MKWyJd9zLRxrxz7SWGRNobLaL9bl3W0Hfb/lC6yOC1hX0FK06813gb/JhXNn5cQN
I2T8rByYIXW28XeI9HeLicS1hVzF8Gz5BfMMXIDFIlFkyNAXHgM86XN+SDL/aTwe
fPda24sQFJQPKHQk3XXSUJScRnKyfwLf3EZTQi7Gg0+baKmVrod0FIqFlmfq0QPu
gbbQ39jBEA5/RV8BiKngPcfrpdWCiv8M8IndPXn0736wbbFGHNidSV/MDEN44fSU
N9d1mTTA0OXgSiyJuZ79szADYNcqAKhcz+gW79fp7xtDatXGpW4yshlaNTqRRvBN
zESa5rtwpfPai3zVg1C7KoIgD3+NWS6So6TAWn+SJ5ldLt3xITKMySWogZSzsCDq
b1Ur3U9VGfxu/5rxEcOJX8wugrw4RpU5TML/DLGkDa4WVORf84IYC3a0BFOaY4Gf
HiDVEAAaduhNpm4WuWUo3KwByNAcETpJu+JcPzF320othRVdjQiwG2VEtFwnlKHf
YDjEIW/TapW4XvbZiLrB9blg8MUdCl6Am+nloY6Ni0VuEg7zDRoBnnwca75Vrz7w
i2U+Nm4R2Yf1XPIZffBflrIx4R8reLi+lm3a78TSeeC3/eXJYbpsO2sa2Alk5la0
ILzIbNKfN/6hq68RSBZfNl7t5Vgkm2sLAKwhUmub2LvpxWep2pXsHlFi4dKQSKZQ
2fihKj3shQa7aLijsvWbvVmbJCxz2WzPlRhS7HAK2C1gUwAYOvfj9Php47svmfL6
fCAnZTjofQJKc7G6X7qd7DOv2Tni+nqzOY2gZmUB7dJkGfXkwTPXJ+LOVM/qNXIH
HXXmCJfi9X4n+eRGUmR14mjcGm953e4G1k1NVVO5nhv09DCsoGv9yP9282RDMCJv
QzNjwUwsgwc76ogkGcXIDfkhvY05SgJar2JmyTa/2kdSo0nt9cpM/F7YxPuKUmaM
z607zsn1ruUbFkhiKviQdy9f5CsPK0y9ErW8jX6CoOjjMZjpk+Sb9+Dx8SIbOcKu
VuvZi1UcBBmV0ZzNaq4vw2J0xUzrsuHk/OBKQpDQeA+j1D7rpDGNNWa3a8LHc84d
r9Ac5R7HfvVtSUimzt2UeWP9CjVEYX7FBfNGaBhPBD4RRVXJg3e65NH1UGU5M6v9
Heh9dMKaBiNFnrT+/XqIkJtI3F9h14Fb7N9zVbV4E2RfiIUX6SRPQwtB68YG6dSg
fmSoULF+iqIDx10P0oxOd0X6yO9c65iaN7gbpktXk8ECsR32UmQn17KORPKP4EAf
16SaiuTsDH2ZANRg3xGzHDxHN9VN99PrkjTTdVP0y1oE8Xpl2R0eEjbJvWKK7mPv
6jy0gRpRKcbhDExDKcfRDBdpOnE241m4keN/NvE6dcUDbCPCTGvW5P4BMOfCAvYr
471JQhAEjS2Q14K3qVIBnd24wrOJRAIxyP5Ybvx2YP9OrKLTZV2llXDHjh1Z7IYJ
Nw2GBmiapUfnRTZBZ+cq4lR9CeidAMEhfJlpcRdJENOQFnRdf8ESNIoc1Oa8mTzD
H4WyoZyqJYU7pcbnTY1Jbyt8knx3/UXm/TO/MfwLCmfA0GUIxA5CDdie8gRqoa3c
Ov4UuIRKhTKAEj7In84WOYhjExIBCgp9rXrviqxMKKqVdoMLiCBhPVa4KQbwMHfZ
2scrEayMrzRs2MOiKz0/tVUCTmo+8RcVm4Iww6ODymkCbC+IUN7H15dJLC6Y91AC
k2UCD/cspeOaSvvOCPY4kUNWEiuDZMyi2UsqRh0kEBfqrTVZ+trcnuQ7WdOkf1rQ
JZHoQgFhLntD4cDiXQxBpi18aCw8+UKM92F+5Em2h5P2ON9CRIzhvmdptm/Ru12o
BZBMJeXosrDIHUu6YT0jv/snFkikh3y6EpmK6DYJyKRsqQwGvhBTfpcDCnnJAO2v
LuEpre3N/8G3V9PW4BrLSJHYRIyidMhXuooTuIvqfZwr+StB+cZY2yYecbRp+vGu
YmuHhAg+E64YKqe+tVRbt8dExtmTeqahKMklL7yDvN3OdMXKZjowV0rlAosfMNWB
+Q6sOWcGgs17Jr3BxY+Ji9zMUyS+vaz0BMBd1ltR+A0W8nwYZjM0yUFnPx8mmHsM
NOkQNbPrLaJnhpWY/hcFGEyUIYJuBf4dvnJoEoXBfGZU6HZW47LUOIH8GnU7/lSl
nzCe7QR8hv0GArcbo8SRYaoTw7bvVzaoOKPG3Gha3EWYooldWeNx/CVDBJkgEaiO
8FuCLDuLQou5h1+jDiQAujseVhW25qC8ziF1msfxBzzOm9MA63V4pXArEnLftiLJ
IYGEwmBXEbwW14OtRJpat4xI5/hEm3L1XKwk+4aafGkd9ZPN7hGAnHO3Kl6fvxZA
6i1FqiTWUy/i1vO+ymsNHiDP2f0pCqBH0ZDSPsJ9zmgTXFu11tx6trlQXvHItP9u
7j5Wud4WcrIQT3VPu/0hfBPE8xzve2hO98UrsEhCthoUzLmfpYPBK8Hqu/r/i3/h
C19BLzLcpvGSQdRFBYkqDrVLQlVQZ2qZk3ox7tXlNAWSvopeZjCwQNtvMyXPks6h
iPzgG/MDkYFr+voLYW3uxaIXFWsKfbbuVsCaxUeO5FHAuephVHnD8ILHon+JHfa1
d2mbSQiXAWMvbh8K/qyYwjbi4MYlEsPNE/0UH5yoqQ3jLy8bRp2MGs6MRHWBf+0Y
X/fchMejr3pY9HECxGjraWXtK2vy6mjbCQnPT4pgbEoDJnMnEwEDIBHao2h9DHzj
PUVZIEKN/BFN2IAk88qw4JcHWe8B9MlcWd6Vf1WE7od38IIsdGsWoF1ezd1lP/Ei
cWk5em9PZVOpZ8C1NQwE3Msg5A/90iuZ3fjldWvXDDNyungiRArMCB8aGuRuHVz9
Ux5gGFe9Va2PYB3mURYWPLDS//K/7tJmprX33Aw1psJISsVJVa99EwEa7Y923qJ1
zz5rU8CxAdr8vIGKWHdSvA==
`pragma protect end_protected
