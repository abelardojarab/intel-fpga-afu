`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oVDRIdOp4aN0BLi7X0JoC2LYb8yabLnLlN7Zl4RfNfLgBw7trw1sJ3ES/Yws3z3v
FWXoSYGv/NHdfzHsB0TQDGWfSbVP/uSzOMRxPC7j5Pi01NSP+s1BxL53tJ0ba1RR
WsWnwbzeOqGKFYpbXre7n9PlOHoTAcl63GEx7OPTPzc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21472)
qlrEPd+GuIIOLF8rTiCxFD6Qch+NB97hVtu1up88EaxdWie+Gq+z49D0/PNL8+mQ
liJR7S2ImvHhF6CYldoU9ZdlKNDxmong2Rs8lMKolmgxzKRbtqrlRDUHRSjSal2e
cZicoe9pb7V34Ex9rxdbcwysyWzW0B03WT/jbddeiKf/YaLXQcs6rwUW32NEPTjz
ahf9DNykhBmid/9G0yEzZKrC9CS2lQ+xKMutAxJ8DZkuiTi3SComVJoZ+aTUfl7D
qhevCFQNCg11iBbqO56bL0XoEgfl7m7zA8VIoVSlVB2SDs9XNLsJfKfBUeA6Tosr
6IbGuPgHlDrQWb1gJOvueh57W/K06aH68a15XmlSu60MkhQR+aC7JOb2Eecc3jln
wrnkMpuGcbYbn5BL3gMs+DlMHq02g3oQs+g/WVxgALTqLGcyBB3thzkPkyZsvxyW
RpneRotbklKZfbuESiyIQY0Pr3mYt8b05rFckYCbp6XfiEDyvCdDdK3Eku2uE0bi
xC7wVQof+g1CKYVy1XvR9N+AxlL6NCdrNCr8GKGIlRHKraKqbk5XEak8Ef9f1Rhl
UZ7i5pu/jtqW/1bJFPPLK5bgXOlAArHKPwuv84AJGDI2hcObJIZOwjjH6JkCyUEN
cP7rx6DnccVzF67qqdagN6H1WpxyGWuQSlQWScCxj5bJvWypnjnzAbG7/QIH5LIl
GgAoK8nBECn6EgZFIJp1xYyY2e5nJMwK+vCDPNeRjSyFhsb64Wf7zisxh2lIWbDW
NDRDUO037C8cGQdmaAlalPOxqaEOKG684UhgVtFf/y8W500O3XR+r2G++JhNku2B
zmqFddMG0CIN567QJ8mQdR1RFfJwjCVbuian+KGNTRT68z8HiHEDv/nNVH8kpS9x
v5LtVyh0zUP2OAg10nuZ1yXl+B4IUzyyZcNY5ALpuZfBO++JO2XZ8n6k22EY3KWD
gn58eGSlDMw9k5XNhn6Yxxk8YqSKv4HkAz+z4XurDAZNu/k6r5Zn6GDNMNK8eVvS
d2RFkpGQz8gfDYl2v7ghBqECs0L6nwPJskV7aJIlSlN/Gt3/b6PcEkY6eXzKJ3q3
COWqEweCc2kQ//pFH5KAlD+7Z6FHuKxsVhBs3Mxwe4N9CRSceYBE+KS88e9gfm6K
N0dGIGHXkJUNsgcMJeaz6yxIVyrcmJwqH8HdQK4+KMtxXDA7jLHj2tqeuLH3YrYm
zoYTuU56P2QYpWAwED1TMuNTNBuFdfKa2TmMkwAHvPXS83jg/6ioCZeFeKabrpih
QZdxPLDJ/a7kwhCVQ0QFxiSt09lhqRWpaNYAUOMoKLdFwTnLwEfN8XMyKxTZ8kOS
CVnZci2yJfzNo12t43V1tmyqf7N2u3o3PZybYxG9uonjQut/TXZnCvWBUMFSkx+3
1g7XuG8CtBmgg1rh+2hjHvbP1CNTWQOeCoSV//q+2S8cPn1T9lPGcFBe3PaOalcu
0aK9ESqN6W7AnKooJN30Lc5baYN9STDfeHRa7wKa2gkmktaI/ihhmKIhoBwdWWfH
up91HvpOO8+cIKV9Xr+3zUizh7XBFiRh6IzArQQPNVJJDKQpWyTRXMbcFSjTYy8g
UB6/Wfoxn8FpaSoBjl5qXS9uZhuU1mUJraVY0EqLp1GXQalRYfrO7nYuV5WiL2Za
kRstq528wqzwEznim/ip4X69whwlvEj7fAy9+93XLolwCWvmydVTsvXOY7spon5K
9QKWYgKyyFNeuWKkE4OaS4qBv6sRPjg9OPB1n+rWbX/92sTguwDLoT/pFFwLGJAJ
i0MTKKjIlPPreJV7PoHAiZNvp/h44U1sCN/cewudx09kLDNCD5iEchSELgg9nFsP
eUyVCs+ITtglk1vodGn/1QshH851yydlSHAl3In0w9uz/aqgn3mGYU7QrouwBnqw
dA2+pnGAyZtowm0u8Cu4Kab+tcSsprh6K9YCWCW6/0WfBToxrik0SrhnrDUfiqKX
kJBcBOl4fO/JhHt7E5NIHCxNeTE/9C/9sxldePqFgskXRKEgzJL8Gc28DdZwUmjp
e17DUug5311P6oSVWfycqsaNguYURy7e88g9ss94/FFewBRCaFUa6blPzotyIMnu
2ioIVubWaD4ODYFlh5Yswgz6n4U0LxRojEh9ukeJZIRM/wCpGBR0xGa1jUCYsOki
k54PILMsNEb0yg+p3boXtfsjl/eFpWK5RVMqK27fqtWlmb6kh5WMdCE6T+FLq5Of
C4wIyTtWO0Yu/ef+3dGhs0S1f6f5xh0sGMeHyiofJJ10/IkXehDNAEOerVZkL8GF
DgQ06UkoLi2fZSmvKKCBp861HUoMkEsNYoPnBEL6KvEN9G4dYZ6OIdz9PCocFXzs
fZJrwoRp76sSvyQ04rkUwN8/m82yKQblLd6LzW9TFHV0+3VMIkQwxNjybtn453BY
lpH8M4UtHRnEtfiZxC8YgzZ9boNzjRUEgSnPM70d469YIQSi9IBWa1cqzKXUn4L4
VQK8tMWozuu7tIBfvcCxJVd/VDLGYAMjy7lnyJaqv9yETw6ndApjSo9JESvXP348
vxa+RoFNEPEPn9YQewUY1Jfv/ERuL5835/CS1PtYOI25IpchkjF0Aa0FoD/iqYkt
1D+YCshLFBJLbbxcRfScdceRMIAdTFZdlMHboLJ3nmHE8fybDY6MlwiIDMR8waKN
u2yTxPRKf8FBw5AsiN7hVD89UCfwAsuo5eChr7l7thX7Q8WXlwQx076vNFGRrFCt
s5d2l2PaDX5IY/XL8fLDzR1AiMpm4ha9Rb5rNPTGxd0Hg75zUAMKIB3PF0/EzlqO
rEm7uFfU7Wbjourn8mM2dfDvm3W0gN2Lo4SNR4wyTpweT46esvsEZimingygpSzR
Esl36uCJFRJrcr81G2OHq0A/Drd3Dv6++mvHJhIyiU5eyyZr4ypWY131zge+psff
FQfEQgP0Caj571JAozZmtfSEdE/c307s3Wb3EBeQ+f7J66CIk6NpGvpJG3gInwvL
PAq1c2eZ2zdobUjTdFyvpgiVxdUhrmXcdQCeJyItPI7cOgZR+nsQzPqGE1Lg/8oo
KzuLXfr8MtFz+LhKiGbLrZLU8REakrvoA203U9ZgGuXkWKSsCSNdkSN4SyE2ND2L
OOUI8aNWVZXbLujnIQZCXndjvwPCka4IaV6EM778M2VIivqesrUcjjlitv25Omsm
jIbjGPeq5RYN2HrV0M/LyqiZkDo8Gh9ZLB62d6e4Df+/jigtlxfgP8Oe0jnXpaIB
UTsXzGUuo6DgY9OHF+OE58TStY/a71yP/z8mghmYg69+xUrsTq8H0DeAkzskBgYi
NL5yqh17cVDdixXw7hL2wUgGZWy/vC/rsZrCTIQ5CaoK8N5YD31YI1AcGxFLmHkN
tubX+cp1L7MJf2pRhN4nNjxTpS8v3tm7HMPwKIxYrn/bzsTOAhaVh6CxlPLUJBGI
G2r5qrhaa48o+d8+2Tp5Agbse59Ot3X/7L2iLl442plslh3el4+M2LegxkHLTTMV
TNdBxDQWhQ6Vrq7W+ZLY/3LwHZnnqKsAav7BwJlkO3Q6S/FvVpjqexfKcVgGy0Ut
8CmIYxWrVHdAedZ3cRUXw0TTBZRbdnvsbpOuazk7tL4qc7l6xcd+0bF3HJgmI7K3
gdzqWFBFfDooJQu+VlQOJbfqU7qw9Bj2gcjWrMRjpPjVnuOKGANOKdXRs9gXwwwk
SW+GbsM63iKjQcSAatZDMoeGpuYwfThR2BjIHLKjRAwqz8IQApztMasAX+kSsAJ6
30uCnXkUivhEFG/IXRXLlW3zlfnp6TdgnwcX3H+V2PpLLB6k9hp8yOIyu+fIanbc
XCdZ4D+qgiwn7SjwpQQcexak3+b5DAb+z85gRxgXTBUkznKW/nMZcWcKZTKXt5Jg
f+MszsRW5p1cOtQhPEgaK3AoZnHsW3vSbeUHDJTQegMRvAsHQX9uMDuxxYprRT/q
2eHzFtkRBXFAS6pWBOrwtMr4jvfH41bkppa2bLrjolUQQ+iHkmZAoVaxgKpuVr15
ukOTtefn3YA2POv4wFyHhPHHCQUuFTlpd1nHxnDOn2Fh1XkY0UxnUb2cYDfwJ2/i
Gl7Zf9Ezw7vs7jQV1TaYJ3H8TfXzBiytgoJl7lIO4X5LgJkETw370mTT0eS0zrdh
55asXOkGPS70o6PjDP7DTw5go+Tqhx15JR3e1FvL6KxpMlUmTjRtquINYe7zP3CV
QdHzl1QBarUOVqYxMccgt8tokVxqIUQ0q8qASMqkko07V1Sem4q4eJYJPrwAZj7/
5/Shf85bY3B6uQD2ehzGbdfqH/8WOkWXfdXUuoX5vmsfEvYr1w9+Frgzea3yOff9
M838ETCo3BhuPg1AF7Funcf+MaEBr295axV0xgTu/xHJovPptkf0chOihmzNpBtG
c+kIVGYWGKikTnMV0yvdF7FtUQvSnt2vgMpYIoa3ucpqnyHHGGujkGdeXZwSzBN0
2cUU82qkTCIq0u8cyz3WVqoyhY1m9aWArLn6LiCHzUwbG91gp/a8GfYSbLp8x83k
W4k/1neNgnKz0RM8hB/UHXnC0vzoG8JO5xBqyL1ZK5fTMG3DXdcgc/WsfwCMsEIZ
C0RqLbyAqmpkKArSE/7LLerMI6Ens8B6MvMy/OWuAfseW/cE+mzG1W17TNIYEWnG
Ns5TRoH2mBjuaApYUew7WYXLKWhTq0KeXn/tZPX36D9qXhN+M3tR+X0AJYMuD4ZG
d3r6prm6njW/LHpWzbyS1pgcuYS3xox+cxEJtHcD0TLNGbjMNVqFtvIXvqtu7iqt
IEv1woh+Oy2Xw1GV7iMLfCU2EHl4MxB3RM+u9bLH6jIHvvWMqyj1t3xzw1/XCIjx
SzzVKqIStKtReXfahz8zPW484cI2kd8ybtvHSE8JnGhLFDDqOfxrEpj/0ZE3ODuk
RyS4D8mlUzyM+ruNHd0NiIkQVnv8dk698DspVDAhRRJ3Cb4ZJjd6idSkwIiwC/kd
fAM3M0BiLdzfphrh3nfNp9fr8X0wy+M6LRY1IW9E/nfbbG87nRtHn9sL4SmqnfVa
d1GjoIOOkmwM9yVCrzZrgR2oeeJLOc+ry6R+pggj1MshCZ7NL3senijhHLS5Q5dI
xlhvi92g6VhRw1aJG6cqCWD3yWayL1yIZbUWavly8uTv4eCdZEX+hW8uKi9O/bBT
VQXiwOuffzRyuyubdo+FwHySmT1WFTJ1AqY9tAhWNRM45hhdUwoUPbtUKPCQhcW3
AICENNqrVFerTl7PAnLzsybRFdY0jG7bY55v5k+Rq6kxVPi0S58MolaVt4h4QHga
Ssoa+EyWJTwEG8QYCzTYfETsfRAjm1FeAdUWevVEalbcuvcaJDGvoYarbtH/uePe
u+QHIQKF8umDe9+FEUQkH6wZle3v6S++THMXPpD05o0KGtNzPjANsVA9unhhnnju
UUbmWiyRUMJWPC9O44kC9rs0qfSWKmljIILkEU3f5PP24BUNjZk4D5psFNhdN0i9
wxEDol0Gm6/+dgLcR8EFCCG6G5kHFDxRRL/8/LNE7EjpBYqG0CWkUh+5UPxkMjLb
ablDVJgWYOnRtAvvVd2B2ymjwjj1glhUoP5W6difLi1pFJ7tLICbRDrNvnjGvsFw
IZe+pDTmFl22/16SFZgOXmF03q4FOsKT2kk/CfmnU0/w4x1C82pEUysnq51DI+BM
+bOIKlZFOLDK+1JW6GD++l+Zz9Szyn3oQb0p1d6UHh/S+Va+cMOye+m/8EGnEcpR
jT1AFRrBFCpfPQ2grx6zrgDGJ/RIcuDJyQcibiEA14OLSXzZW20h16ilSFxcEHhc
0fLX0gvkMHXG68D5DnWB7Thy06ax9v5rAZx500ggnXPq25WdmKa9rdAAb3itcJQ9
vIbAZTIPENRgJ+fFurCPIyII6nP6yR92tLPylBaAfGaMD+ybmP6JgmhkkkarBxN6
TCLmdTsYkpPSeQwmEorS5nK9BTvjqfZMp8EuCtrrQuzaDA9nL5U9hUBlPbAP3eR1
5IPPAhuJ4+1q6A23KaLxDLQLVCFQhF+7595PNS/Fj6r5StSZ0s1zeP7eus0elu6E
8X/UHlLHO5JdSwFlOUPl42W2k+h1qPdey7Y5q+xmDftdZDL4vRTu+K40ITD/5fJZ
xNZg5hs3dB64THF6jr9JLqw94GrDK8esOxk2MHTtxTJwS2zr+4EaGjqv1YMN2Uo1
U4NynJtUN2RxdZNfvzM+4jhtLdiCerbpwDWssfVDNLK6szIeEG3URcDuwtfcuPMy
cJJ49QYI4wUnaSRAsFrC7/+OD+DCifJsFtQlGoCWfvInhXTWNdAlMsRNxEwkPBjp
npDROHtQaZL754YNKmBLginoz4enxFR7TZumLdDe/NtoOa4EplxPV8AnUiGm1FYX
LdEtT2rFHz1pNLeqGYVC09znALYDPEvHds2f/u5W41EUGLGbNYJeW+I/oqgovDWQ
t+xBDChAFdloMQ8zC2Rnp6koFNzdYsiNWvr+dpmn1+UVvkF52axzzvuExTe6vLO1
/HQNhy9sf0CcA/f2QTHWiilGWPh6vwN5M/ul+WqX07ir4Y6bG5yyhAFuG3Qt5w9y
sahWJjqIUBifXWyk1D2nl3OziSG/67jzMmMesUlFPC+EK7u4a0zn4VWkPiqSTSWd
nXWF5dphn9yh9POhBr1t+dnhrDmIMo32ojdkjuiTeB/f2CHYf5hSwuNaA5+QdBYj
vNbdyIHdTKIR83nZXv1jokdO4rYxtzZf7rEjBie/iHk9dqg8pypHC7HKDGNCFQip
yRQd3qvjAhuom5XelVW+mLjZjTLcmWWh6SzWWsy6efuaJsIDaQv9yAvlmoAYkTTu
8D/sEScXT2vrhRkmzFOWlWINwMp/aWSJJyckE3dJ428XxtYnWwi5vljN7tfea8dj
L9Vg3nv29cv/dvG3Cf/mbxud/dpA4QCpOits8IDIol4EPDJKCrPEUbzWsX1DzQn4
G++/6eeLwsSIz8Ij/TxhQfKcmkyP6Aa6x0nzG2WIUKBkwz7SMMg+HHKvLv3PE8nF
AM8yTSe7QEPqJRPnsD4vrbDgzerQR5QtNr98c01E4KfD1Wo5NJBYxZhZBip5WfjF
084xMdXTxCR6CmXLMZoq9XuO27n8MzhYt40SjQH7FuQvSu/TV2AXMiBX+byuQXMW
R5xDCMmvrnMR1KEEhks+DLvazvOJFKNB9Msld26WIHZ6u1aGVcbtUAdScHPzy0ca
mmALkbadfnrAupKqrOCo9eM5pcAM3CGOzKxohdNNDbxHcRMxwMSjOudb0HUaqkPS
T98qc+b+m3awjMV1W6RFOxsqtrIE/1BbXBn4H//2BE4JXvEWdrAHhEWJ/iP9gBc2
agPX1+F8zPoL/gb5drcJQQzX8niqJakrkP/tM0ammWMf6lFMPh3GmBck8HOIQTxi
iBh5Efuv1jYttmiTzLG9YsDa3ioKkwW+u84LyLo4lIL7H1VlniuIdpGMhsSusyrm
HLqANKfQoOBmoZTXPMBaEcveH9t7uCme9SguZRBVU/lliIquufEa82WldT3agfsh
Z5gqoe+Qeb45DpwF4B3hqeEOQ5mFTUfK6c//LN4UY2uTzQG4U372W6QthkZqJYKm
sDO/g0jS89Yxw/10tkMj4SAlOqcNRLOtqow3KCzuOrSEh9N08yWiOUML41WKdU0+
/Yf+UiI9mk9IR4D7sKLZXMRnlSpEOfMb7pswL1X8CD1HyUdz6uQdmFVqLUQi1bQ7
vdL9q8A3R4kz2m2kb34wGOwfhYlWdJW/BRJqSk5P79UXA1hw4IzP8rIckjcQTvdQ
f3eTvccCQF0+jzJhYMEuH3JwXTpyVLdRZ6UqkDimfcztvNx+q+w1qi+WVi6NdT++
PJOFHT2c352teShBkgOj3ZZ71Pd6AH96kfdoMAZY0fLrDOcpGuN+8iTfeV3S88l+
RzInaGxQXOhKS5xNaogklIBWlJUbcjWqqkvw3mlf0Zv0Gx22rk4T+ZmXsTux7e3w
/aH85fd30Lk7UIX+zM+N3xrOS49HjzTG40d9dK2BSxdj2lMEJ3hBmI7zY7oPF9pK
91VhlBDy/cCsrs2RHDpbFmdyEwlnGi5BIei8oKBn028khEuYTJ2VuU4Wk091PUbZ
ZFAkhCmEAOq7zOEPKcEXef05ZmKUqr63hcomLkDRcmkYjm1H2HwYgIV/+9XRYf2M
3Ue/OK40AaF/fkUqPosuJma8xvX4tAJ1KlNWrmnVLDeXJUgVnp2o5eXx47435M6q
IU7Yl/9jrNVFHiGwkcTKcIfWie42IBUk+PFHrE+MVOAu09nkH4g8IV5nokDY3130
SxffblrxLBNF9MEul1qqbEGGg5fdNR33Pt2JlfWPQRzAZmxd7HDdPLT/RdPPS3RK
SDFsgjFP+mrCtizttFDIax4WevM3xEWJscB2zJc2RtLefaQ6jWn0ibAIkagUuk0Y
ZjtBDxmYFqsewwd0XaLBM5laGzaGyBch6VteNM633n0xIptyUPQzSgg0PMtFNaqN
h4FwMhFU6DYeNWhyVVbE8ZpmgtRCIYMRJ+5N1/7qnsyKLBgfopwSduXlEpM6k+kB
G8RtGU/65d39aSO6wEgfu7zlOOnnCiTopbOpVMtR5aZwj+HyrM32zWaT199NQp4d
nt1VVck5qcLUd7leYDxioHJaKNic9pYZ7wjlFoIXkdhgOFl1M4N+DXK3BDRRF2BP
s6rqKoYY8Oxshv2KhP48XoLnacpfFFANODCVrMq/JwNVfKXdhaEiWx139zhBZr4O
yqs/QlTicm8wmbjBF2iji3w3ndIiwXShhKFpiEmKTEdVo0DjMFINVsr66dcVIlkJ
BoIrViOk+jpMFo0DvGpDQruKCdR8qxQPsco4Dq0yCgvxyrf8hdTtuj1XRw851viE
cskJ0ZkgNA5E63Q0MhtMHF0KQatN6tRdbFE/dwU5IxODzcp+JLiOYUk8k/GYsPhT
shsi3iwiJxBtjgP2WagZV9X5/pkNUYdGzFOJ20DUNwkOOohZ12oZ5AhwTCs1H1bd
tpSpkunDQ9aFClkLtc4Ou2rX8fyjYJHh4bSp0i5ES7XV8dQapzf+jbq7HKURlsOk
j2XJm5zypGs06a6xQVYwlMkiLTuYiEsDIRQ871MQUfYNLZFViACjDqlEE9hsk9/c
oQ2IldFb2vkFaowzdJjgY9qTZf4qA7delPa7e3KpEXqQhFPpeAut098eoefFYWBv
jI5jL8JLh/cvNaQ3uzk7RlU8+Cz0v9GBI9sB2PAdIAMvgWDhHEYMie0ZDKE88xUK
GtbEARSzZv9Yz8UdN/qi6vhAk77rmDtSHROTQKPNr7Uy3SnjPa8ggb+oVNKFXvPi
iypLbJkKUURHWvzFe6Msz+QmN4okS4am3mHDVOsL1nOX3k/7OwfhX8body2QdUpC
e+Qyi4j9Yqz/nswKZuyvgEOqbfUusP0BfLg2d/LF9ag/nEVrdk4oe4bKHoZdyQFC
JBOn3Cuz2bwXoCUGt0csIrsSm391KrEpd3oXbLhuYrGAh+t4Sek4P4eAkfIIwayV
W47cJGBkM+KshTPknFqFxpzKTjtvM0JbDPJVj55RVdc/Dtbv0lTCfhmCOG/U6vmu
LQVU/c86UjbML17ETGVFhnAsPFlYyjLhEjgI21hyit4CLNNja0syG5W6gG44rrLz
XcVzUm1ViOJeqJ8AHuuVYIykZ6cyo9ny+mZisXO60EIuv2AzmwT5ifGav0nhVSBc
EnpvoDlor6eG723BMQzPOf2tZ4tDcc5sVhdhu11VoJa/xc7mtkkeccpln4+XLVUK
8shLjMaV3R9kh7cub9r9HP6ELZwgkeP/9fvESjybJVBzGdB7sXwD1NOlPWMq+as0
GQfszam7s5pMsHN9QZhgKmvGylR8ez+OL7YVWfjfWOfqFG++9QjAMlpJ3OlF78RK
fso8JKq2DQ7yiMEkTmJarGRwhADdwNj9wUGG8oxd7tLQqSVX3JnfQe8Fhg2jB6VI
mLpaFeReVNwXUPkFa4uQ7lqnapegyQErpcl7IrHDFrlnmAHjtb5X4YRXT0MAgCpN
scwCFQN+NS5IYlkS+g/YsQFyYMYDZ7UPfvBiKi8DyAu5Gq01GI2Ec2CYy2KYYZil
GRY8+3pAqZlYozQby4goZVJN0QnMhWiQOeXZD0vVpeH6Y3wrWG3fIBKoay3AwkID
hld+kFQlwfQxMyZvNrj5lftmo83YsqaVZrNzbQBL8tGB+FLtG6G++dh+/2hFfIqA
w5qYItlLHdcfV/RDSTFevvp5H4BG1Esd7EoGBj3ll7eeKGdtpnFvcbktyySVKY79
1myPd/QjZ8+tizqFBwNKm+JrJzYO8yZvvqtOmxHeLCxsReny1g7Y1TskFBsiY3VM
VcYamu60J62kygTy7IRsYRYS38x1e6gFE1tz3XpB2SXyE+xLebUpJ3y6UUhsurOM
cofIYePmwPbavk7fYmywwxhc50ryO9qvzzUunOB5tzRJI0OCAXL3sq/f+gVTHaSp
rif/gmKdY2fjYGv+52Tujvr2xFhyF2ABXa+dCvw7OLyL05HpGKAEIDpWbd/370vj
ygF/UlwE9ddr+LKbMdllB/ZhZBXHadDGmf3JTctN81A1PrEY5XdiEVN1ST3vTWJ/
L5NKAms1qGzPZBd+TpK6wjsbFT4Vn2K5SSnUKmhaqmge+TO1vZNjCJZpW1EFQeKp
gRGIIwuXY0uQQm7I+j0G6QWyCVobk1LF/0VynsXzbOkH82dQg17xJSpmPe9N/yo/
doBrEXxjyoSz4XU8B9W8Hjx2oZ13ayq2IObcjp9rz+Zp24b3NGAI1kv3Nzq/+ljs
hVDeVZ9jUII72Jaoa2/Ir3h4sNOI84/l+ETIKA+0rZH2N69qcz4eK242TO5B2bIr
jPoFXji9zW3x1p0RFiR1xtu35amqAxHQ/8BbQe7VVOUHH7ZYHZXz6bBJRUmoJA+R
bXLU56pO4vZprbpgs53lugKgR+1+9q3tWqWIM51jzBcKskO6Exe9suzoik/7h2MR
HNkotQvvaOAS+D+hDbvjZnEzmKqWkkGwYW+ZQsDG4dKTIA/m7GmqncoOXXip92+p
1ooMXUSzs3A0SICLljcKSsfYCwZ6OPIuSElb8ouTWiMXwrjJj5Hxo4GqfNqoQgUc
1h6QTd/UeUWn1NHjdWvvuOxv3qEKmscKzAQooDFKt56u0T+lIWK6OUKSxr2sZU0/
F4P2WAQIQ+NtPpQ66vTT+ASbBbWUWb34JESC//eXfEgViQwppHYWoCTWpgORg1sk
qM1kamQhBQ0nAXzHIUfe0G92ED4nf+RLHx3BzGYoCX+sS+2XzCIQDCxcHMM4DQhM
5+9t2doSj9NJ1tE3sOuWaqXIHVxCIhqBFFHSYq6y2p0cQg1UCKqo6ZmpPoYN7h2m
elKNSoJ+qZc2J2/3ERp4Y4A62qtbYBXf1WpqFCNzidtT6QMEFxmbKDrvQEmDp/uM
AKOjFh0rhIeN6eszp1kPtCHbpc447UlHpPlXotNEC7OObiZpf5g5ky9FcfmiIetC
yQDRbJFLyxRkKmuPQrgGn9ZtxnHJMigTf4I70ZKbj9OxLmtsH0IRj8q1Rg2cwSMT
ulAPdsyK/IlG4mS/E7Clx9t2RKpWsXp1Bw4Q5M9GCD5wkUg5nw1jS1/ySOwNP6Tg
as6loF/Ls+0RZGpD7AY5BAjl61CRLmxv5iz7FebLmF2kcwbgy8thJi6lveH04Jvj
027yVyeTR3FW3fY/7D7RlTPB7onqa4eQS3aK8p0HTk7TN8OZAWidAtseHxoTzUfd
nBF4ludbKovaWvL+xWC6KIEC5fUS0Eot8CivQgldKg2kz+0Fizy2NzU4pmSWTwGH
JNc4TkzSinMnyADLcdTiHVo8LlNntpQHRcdO4TlNGDEWQvgwKGlBOKsPmoNulQTB
bHxar/zQ8mdlshFIln5PZ1NGWiMxRUhprU0loJPrXDfCRUcLAGBCRXN+awNv7/Nr
YpK9AM/EK3lTOnn0aSXMRp5LegCkdvDgCdEJSLAM8TUGyF+cZ7xyxu7oIli4KvCR
WbP2XoLoT6e+yBQCBh2SLoCCx9E+ajIxCYlMmSgXArUBIXkWFtQ8Ql4+wCsy1xdK
e4u0UE/iFIbCmbGEji9fk41/lb08BlZr9ZuFj8YYN94PrR5DyunA1dWn4O6y72Sj
X3YHeI069x4rsJ+jap8N45oaw+yylgp431iwmhPKsYJVXEijMELrxN//FDRjVMY+
yXGFOZterctaamEB7edDAiDl+eKSDMnnBzMFBKbHzqvrBFHpiwC/vCAoU5Nh5+rf
kf106VlSE2V6O8LFmhHVffICr2OalabFy0FZMSmf0iQbLe4w/Vk+kKvrkTbR6qrr
WgZyY/vJw+1xu0aoTiaxkb0ZOa0S446lAUSocAAuJVuQR/xReGYfpTeBJI6Dbt14
XFMo0rVwABzBOST3P+fzzzkd9VHbWMPtyKWYXaDKtjFnawrSBBN78TKkPl4AcBaF
Sw2TGaSmrxS2IDeGbNd97ydKeK0Sr1DiturzCkQFd/+uBqugupo4/s+UE8rMOiUm
eput9dgrrgLwDInqszHApi/LjXGrIg3MjSrv4xknhydszYzh6SCogHqT6PAAc2DG
qn68f8ueoyrI/HfHVM5afqvfGt/E8+UhpsGiLOmUcu1VJz8SahKOP+hE6/eafGgb
9aaTVoykcddmtGC+nB6CWtwmUE90cOFsXpy+B6nGF0VwhW/5/WV4Qs++c9EeyO1h
zxtafnijHdVfGv+VmB6LFHfGv3NX5uQxlZ3KSi1jzxfvrrYEEYjbW4v1VfxcTYCA
4jfDiJB5HU6afOQBsoTAwQKQMt6Omyjytg7bqdiQiKnTCnqmiwFcy2Fw1i6oHr5C
Oo9ECtjT74duoam3WKNKln8TuyqQhSDFuSvR7g68RzJ1lndsL6P4B0MHHHjFKTlm
6ixXywet6ygk5iQYD4OyMv+Rjg8J2h1K5F9Wa+GnlbzdgKW8FJywx2pd7kDQwtx+
f6rk6JFmBQjL4U6jGv5LtDVBMgiglST/O1rS5OxMiFQP9qXuJi73Nq2nty2U8IG+
SfRhOyk6mJHFwINj1MdFtKLn4IFbwMkXquezeVGFl+jV0MDVMTNQJ1TWz3gjKNR1
PLhzxVYrEKjeQsR17yALX51I6Ur8UVpBb3vNBSai9zzLrocR+iLxvuwKlv+HMBIW
2Dcmh8bsDP7a3JUBgPaccKfksAlGnRL4su/2uph8fApBwNwhmZHs36QMWD4NjGTh
ZTXK0VbrrU85PPcgyFbG0euV+j0LZ+DvlO3vLEX92tAe82iJNTia/GAfTihZcDkU
noK1bj9gvcxHedzxsVI/sfwTczybX30BprvQTLDQS7VT0oyo1MTwb28sfenT9n/z
cYcHTnxFD1i9v0YfjlZZXbbETsz24RI18hELLLmdQmSQ+37TjRAu+pEPhiWe5K50
v8U+l+qGmqmF9t0BjgI9iDRsIZGgnE37Kj1Z8mLt9A91C4A1PBS1O/E/aUVp8MbU
ICfFwty3SQ83rQ5jwuMNiNDPlXy9QqFRBp/5uC7zr2RYrV5PVAakoYiDcVBDSBNO
cE0cwGdjXY/aFj0xVcN+4c/WUb+2jOIDVl8dSGRbd0u2u2heeYmsWPbCGWiWAuhH
++va213V16jvZSK+UECngyOizAuD18ARG+ODOBGikmUZLN5ycHZmUhckQcwQM9vY
b/cciHa08puWtpzPJsqn0ZU/F/IN/t8t//mmtM2lNtIHytuTYkoJaoVg8Gxx/Y5N
UOiWho1TB51EcwDgzIx/GanQjjCmTet3+7Zf4PCKZq0KKeoK8Y7RQziY8QRaHCka
WGBlLtvhikJV24WRekZReGAeYNQTWyWPZsM2OylMabcJHZnSBZNXw7z9ZpE/DOme
PmU2kpgYS7nURyftXdML1IazrPnGubSMoQthiPyYoaxFYtf4CEbm8SaSiAdMv5Vi
E+KXj+93fNx6l8pWd087WfB8u+S1zGShTwRDWgc0BoH0T9D/9CuB0eHM0aJXtR/8
i0V+y3hiKFnvZpSyLFR3ryobcEI7XhsYdxGDqWv5uFahC23ucughCF0XO13cJ7X5
XSUYqiaa1ZHDZbuMz3XyMjfzVbwUMEBTzf+niJZhlrySTg5CVxV+Bb1EyXja/NOi
Y55XYa4YIAk+eUfnd5r9EFBaMOp1E+RRP0oO6Npg38YMUaRtdSgoJ3srv6dW3O8E
6u4vY1HVGIak7Tb9N8TQY9VFkdTE5O7vOC5Ds1hxQxvlEWbastVL2MSVxRWslP6V
yxWr+Rup7FcVnfCpi421C5/S8Wba95v4tFYrhEnSvgttRvk5quAIa2j1N23UiZHn
ZU8Tcyyew3960eEtWy+hH54EssIDdYT9mqNLmaz70nGbG8hJh9gliG0km8JWbDIF
zfDes5D7i+Whb/kgBCirfHPzpmvbnffKW9Rb+jfvL51aaSzdpD1mbf6zWI3hJmXT
XDVvgmLExMQ/TJEbuFzvixddLzJOMs04a58l95Yk+iP82mTGQ2eLFBxRzw5pHTjI
cUM12mEmSdvgbLXVPuYv4MwcIG3PGN2VGRwNgEmWTS292u2rrujqKm/T0Ub13PzL
TrFfUljdivPw/c+A/ZHovKvHb337mUMKIOqdtWwk88tRjaTioAG36FphCkeSy8UN
cXT3pYl/hx0KXN12wzk5Vau+zFaLDVBOKL3IQFnNzTPsw+84jXDt3ZSDj+pfc8Yp
kV2NIN3UY6BxsjgfblRiYTxVLyhpcsz3gr/64YN9FlwMf8BwilgD8fBThjhhCfl5
JpDOAI82ykUKGxFksr6LhdZAifq+w9vC9hF4ZABtO5vcGVYGHfAB8HEMiwXI9AIZ
yMGpAQOxQrylnl2XzYicm7N798v5gX+7BkYAni+loNmq8siK6AGBitas9plW7dbI
6LZ4MXMyniFP+hX78Wyr2sVYEGEkRdliObmMxZIT4T5zAxmleXyLUVaZAfyXwc0O
T9scx0lqfhdmzvSybjZB01Pj3NMjrGMGynzfvpaV2glNWReQKq1eyzx9QnUD2QEG
ftHwkPL20EhkyVI74Htsq/gHcqSoIk6ZavBqYrzInWo6aW7eFeqJH26mMgkpFX5y
3sOFWeeEPpqBDFAUDwq8iY6/yRbmMeDUmx/G2x2kw7h27wQs1XyxtzKQ/jdwdE3V
+zn3WWo8pyHxxwqwvp8HbJttCfYap4VhYwGWOBu0AFF4g8l3dEh3d06bzVj+epU9
K+7J8uhL0aKxMgObfygxn4d65jtCWzaot6A627VLBPe6rfX9dt1695+80Gf7Zj1m
daC4XiugNgsgbhX7vs5gxnW6YRao0tzpylFLtNRlx1ihacoRaAYcWSuyJXS7ztCn
6Javw10mmHBT/1BQWB/p2p3jH89bC4cPcm6t/uTfVpLLgEXDR3XRMET+t++Jtg13
H3cVV4FMhOcNWUepXdjOj/M3vQi4JooPTzAQ12AiZ4yYudPc0OvHkF3hnreDZthS
VkJX23GwFDyiSZiBpkYpVHJFCz7S1V4v1LzkeB1esoiDeaVMoaRc8hY7QO/NsV/V
jTv3GGePmfDzbtJe70bOIXH24EKTNy/XozHkbLr8PiaIygyhOFxesvrXVrgfOsT+
Hn+1ZNTxVqeVlsRYnm/WIKNAcEefGojKeODFAP4xtnksYDkvuz7cMSIQrFAHK4Zg
9rVBsbUzRswKQinjqHE4aOwDLBVxAJ1lrDRrGW3+DWAwJIjd5ZcGoW7+H+IFhk+e
0T9gc4wJwPrTIY790ZNKIccjc9Ww2bNWrSl+zQgED+P/JxwhvissR55Ee0frjl5O
RVeLv0xggYoRUABEWTKkj6W3OCUS08PxPeRM3bushEXe40yKw+0aR96qOZvfRG3M
v8yDIjx0p7rBkDS+6elmBGdKawy+ejzxC3rKZlgJK77O9iP0ozRmypOIjB6LH5ff
3qiwNTX0ybzRNcU+6EpkfYRbZWQSjAADaFGh2SDwEzM2gg6DY5V+f5exlEOlNwQ+
HYoF3gm4rfrdKu1nAHAiM4NX1kQMjnoY6viZWJclXdZFoTOaHLkhbXpQsYu0GgNa
eHnaSSf3XaoNP/K/45THg46ATZ6fI2J1UIO5vgU52EGMCOIb+7TEWqrpeh5rQYOj
13zfyTqcs82WHfJU6ROp0lJvcUViz1sWMVRzn7oPn8iO5ws+0v5KKqRxM3ZAarkB
TPjVn6XRJtcOOZ1xVSI9c+66eRaXB64oYs0DKlFvbM1MgqZTS+JkfCnl8DzR+wOi
tmaXGAyPVC0tjWKI5YebM9zSQtB4CC4P0Mdi7cfAAmxfBUgItxpJfwHRvUIXXlGg
FXW//e6mQ2bIlBNuOJdXG9hZcXC4D1xL8EwH+aCvjfOlI2KhiPsPkHHHo/cJ74y0
HuLZ6W1l9QYn66raIQHoMxHALriJkTZCxcaUQ49JHXmEu4psb2DuMv0vaX8obe+g
/3t6HB9k275TfgXYqCc914tCdcAeBngoSm2z6cwrBt1M8zfPBlGftpG4DaSb5ETq
aC7LTew2u3rw27uyUdD5EKuXeaIzSSeOLJMSihgpxkueDXjt4XsotYAhSPQQaE4a
L9SJE/fMOApixrCo0h0eBfHx0m9Wc48UMzetcDWiGHby25v/nPoHGuj6lKVnFaX3
uUKlKvHqFBBjgtbzBZhlaH/BiNbQhV16CjCAEZnQ+/K0vn43SA9EhcehN6HK3yix
Zb71k5OspAKuUyfXnN62WoitBGP+wqpxR7OrD9RFZKDTLGFGGaTEZfQYmuDoYWF2
zJgk5nx1eW+JyIpt/8fatP2tKlvcprvwlbnheFZkYXz6gcj35I+zi6iBfz/2NFw8
U0OwezsgHQCtK5qSM0EaeDJ977yWAMqYoz72yIRBLginhRUDExp5Q9EPX/l/b/Rm
u3j06AZso4KqMlhT+Up9yeXb74Vx6vnADmO+sCbntoHuR+YrmfV0lyldjxVcLG5C
OhvFq6ZbPQ6+OvPfGtEKEG8B33VNcSw3YE1ILlejubUKRyz8l5IOOTvwsENR8vVS
16qicAH00mYsusE7gHYF7vCYICz9DwelV3GSfafEjqnqeOpzbD0+ZkL37yHkbczQ
FbUyuQE4vemrTF27iQO4Q4r4uEVPvOIy8xVEbNQcnm7WJtEKW4HtpaOnEdOIms3W
1O4ldZeMqFC46A7CHcKhqPNXnU2V2q/DF3Q8yA0qjppGe/olZx8+5EP7zsQn6T53
BV1JwnGoZK0nI255OscgTkiW8YSMfekXkj97LE28ETjKTMJdfTCP0331c1qPD39f
B94YKksMlP3tg2d5B6q7kEh0oYPEb/CBQlreutwngoZpGSBSD0qq7ouAoFkuhVv3
rZ8orEVF0W8uEWGiQ2gAsSOkWiP6+dwBbMXRXdJDKLkiPqpFJtmq/zQjK5BtXPWv
5CFbnz0PGKsA0kN2mpMY/dLkiG4bYLk8Vrw/nPuiTCtdFNaL6QD41LxmbigsE9+y
AYld0wmaJgCsLKT82DpjN9jWrjy8AQ4iU+Xjn5dXWy3tIGmFCdpDqHf4EAjyWEUU
VH42n8giTzPA909ubzUVpzim6uhdCmZfLROWR6Nsyezdr7vNYZ+Br8aua4XvasEy
S9gaBd2DIWWrB0jZzjVgOSGM3zGwoXdCZvP+vyZdAHwL4vwm70BNdBzAMW5G0HMY
nC5RWV2mZajFB9a2gaBGkdoyiigslY2v/G2yDVt4zBIYY6m/L4UBX/NT0oFKsv9j
3I1C1Maqpl5yqgZ/70Gagkj5XQvNPHkvD+cdf8ZgamLTyZq/Yy+erMsn6Gc/gl8e
OPKYuTqBZClQqng23GfdIe0EYfXGLh0mXlRpPhtZyDlojNjCAAUFDE0mQkHIUnyl
G0kL1Y4WT1gaNU+ZPH3ezcmf1Qk49aZg6R8w98dbhbWx/YnFdXI1m2DERyCF0mqI
C/xJ6tvE6NQ/whOcoijTj6MlhP8omiT0poD5Tx6mdO32ePxx34MfddTHN/j0qQVE
NdW7ARzp3AhD+rZJ+qiWrXmF2pI8xgCmlzy2hQy1tIk9w4ZMFI4voGNqtBYT9zp2
+MLO761M57wIdEUAEvkzFDfzBSfxyB8iHjNRhsxa7YBKowo+P0iQm2NdTQbV65tN
0H8o53sYi9PMDB6nMnSRcevEr4ECz2pwp1VPnjUz4V7Asz9shxR9lJpTLvMkQf84
Yz1P/Yyjxr9jLbTE3jkzu4/umG1Nt5W7RICNRoauAWiyx6XRsOdHJgoi664G8zbZ
HCo8wAGDoQTekE0dtKc2KY/qrx5FsOiWAQede8aK/iF0Xn0YYM76Ung7tHgiOXLK
MWHnQd+KVqDfWgrHmWeOj0rs1C59T845c4CfJpOs2dn0zm/WIgv3ZAOYKhTlU8iO
BLHuQzENlMEUcrqKIgdKooDFUbh+Zo9X60PxrXC0susj3umYHulOm/mQSPjy+NkS
Dou1vBnbMeAl+A6wCh2cp/E9nHjK6oaEW9nvZXpCp3O5bcOeHUDaPXL8LEpVcUVk
PMZXfN89DSkBnWthNdfKQBsICnEnrHyyVzYyQntdVBx3sIlloEtp8Lr06O5fBvEV
pokAeqrqTtLR8cIFP6+SHnnMLatQWTwWfMOxFFsI9LefRGtXpbpzTHn6OzQgsep+
pFoITT/mk2zVrxMGmSAYWI7RFdosu+SG2cJqonXIIdvr7XnGyi+VGfnAR9ubQG4O
KkOHyLPEQ5eXNhTDf8jaG5YDx+oXFrIwrD0uQ8MxuE/RFknkRIIfM42iPHmSW8F1
9O92sW+tr7FciXGPkJArMGp2WgIPZJzqqE56b8tvhkw8likyt+/+6tWhbgRaTqXL
MM0F/P+LWQbOMc4I/k+3/4UaNzLLGFMPESLab68bORa61uvnIXY4o1eEH9JoYY9O
2wkNPk7RNw1gSHwB7cP/yXMZzto7+NdAbvfVRiOCDdGT3JwQh8ZQ8wg9nTSGBC/4
f46J16rU9EaoY/ElCR1B5oVm3lK8MTS5Gm/ZB11FPHIbCcI6fTJP3HZm6XLkBbvW
Ld5BhwmAI2teEu5yj2g9IWKWqVuE/e31rj7onZpOPjfsz1KyN5oS8TiixHakceIA
Jgnz0Mr8D2sHIjLVngcZvrKbERNJlPU0PUqpM8D5cG/XopVsVbvdgaBXyDJaBK3D
42fSksMIQZD5B089axC1l4ImQIdZRz8+x12Vem2Yk9oKbXAMfLJlLbev8ZFhWn/P
LxP9Cy59qgGyKcq8sSxfqLrOtERaiS4lvWJDMiA86WXlXI5ExrJ5TF6cdQUu/WOX
QMJDtkmVGwq3NDfrs6mRUrgRdsb5bBZIqlMDfxAa63HPzu/zWURFccUxSJjGWPYK
q8XgFhvWMpfDu7y0Rc9W3niaD+GftJfbNvJtAltdXwy/WcDbDznzV+ToUhsMdJxx
NTT6LiAtx0F4wji7vYvqc4XDfY6+R4qMaqBLdMI3SFaMpQylhgZjMKY9gh5gbeH/
Jl64ANgb1q1oq4Br4AjidodG0YjJpo76zIe191KcNtzoXZufB+alISO8Jq4KMiXr
G+2gE4FVts/gGYMbqgEYuRZo8p8bYNln+n9wT4c5BuRLXBXarNyg0w4cKpzbVhpt
SrbxzahxRbV7ZgO0mPXDAz+iVC9t+B9XBG/rJU4BCCsnOQynmMzxeSybC5FTpP/R
Cc44237yE77lP95uKekWiiq584q3VzJ3Yx1OIp8+7xgMp2d+bnpDzTAG/Wj9nBhJ
SYR8Lup0i+OuWsHQBgS6ZX/+rDnXBxjUYnX4+o1Vm0EB8QGsJippY/8hO7K6P0ER
AvvcUuete2X1mnXeXc7EObM63S36RgxZ46ovAovuxQ+nqRmjccpJ0+09T7whjDU8
R9a5tTxHR/KyQimcE5/Li30wKRZMJN6DdSTlWj8XkTe96FCWagg0prLbzyaUPkGV
jKV9MmTbzdYWgLA3FJJrG1hLG0HZTT+vYIxovbTtCsmaoHmXh5nofCUUzWAyFMX7
R0FcA67xQN3TQJpAUOsqAh+j4smUQcoxzpHJq+k4y+WJ0lv0KyvyjRK7CkRMP8Z9
/ldxmrUgFmNKwpv7gAbyneHp584Qn3BzC7UnEdC2Jzrucff7mid3mhVkcbF/gIeY
vohHfgYBz++gip+sccRjhfvOhe9wV/pkKiij+hohjhQG0goTxU1J4LDurgLchdeB
aTeznq62XNsNQJ0kM8W/eFoc+9F1L5fh7V5A6H1yJ0fEYZfW0sQnmyCHUYp237o7
jdXT3qfCeno1QyqvHu04r9LuWC9Gg+cFkmUNt5cJGxHu96iQVbT4P2RrExD9MA2w
yvZVFivwH1P7hZiSNx2rWERcMbDkYDZvL5rDHDMhrpmz6eCcu3VkI5xlR3r/9qvJ
ina0KfJXs6+pbBiJ+9sfMVasPgZvLNwBpxeOEHq9NjhLzD0LtSyCKubPpb1Ih3XG
Nk/m+49N1EqfPXQzQ5RQGsiz7eUZb3RsoaAlZfYRbLqPgd0/eSsje77KSIOk/55N
X/enXSlEMaumqEn5jpbqRqSpJBLZ8Qh0NrDu6/yqHg/JdZmP2TA+GG+Zma21Vkju
N0HPMTpk2BIwCTYxqhaNKdTMYlnJ6PijdqPVjLTtXQCJ9SRF3m57bkOxbdgBAjbm
4oMKQC0M5HfYYhCkcqSY0kJBWGwtAuWsgWRTq3fW0J0BsgWcFTm9lFTkbZbenMQ2
l2ewiiCCcHfZU86zgAH1pBsvpINNeO/kY2RuhNs3cvKlumFYpzkjF8dmT6LQbBgD
tRzX2emMX1twQjk+KfNcnrehIArTHwcLqTgQf7UxOD9uGFyuIPqcFBeU9RyXvAhj
zXQZTQpWBbYNLVT3fqB6KRegk8E8j4Cu7ZankDWcQf2yC+G9UCMpCIbLnW+Lc/qj
CebJm+shNtvaG1gqBTa6/65w64u1eI6RjunhSvqu8evgx7lol4Hujx9MnvvCYPDQ
0wIMcFtIWMoNVVEZeSGPvUv5+EYGjd7jviV95RwdnFkKsiOd8IXQ54ykV3lj2xk+
KADmr9iEd/76bmJ8cjLSmbQpeVlSZpHDisSx2MrUbhHIB8+sUM46zQjRxwyp9L/+
P4GzUTsrWfFmjRCDFxZajvwIKQbEZRi1LCbN5KQfGKCsC5mqHbjXgHjLE6znjdkZ
trWlezVGosGUo8Mi1XsEHZfcQgMhoglHTFYy0NMfTW56Yi9xDiwHzBtgxQHYFOX7
E9xkHlPbVPtnJgDVRzpSuCP8tH2qykTls/uffTtDXL4jvkOOkGwoJH54n1Z38DLx
p3ltdxT24TyJ0pCZz7DDBzWpRM0sdCGSO19DVjiJ4DaQUROmfS7B4Kj++yHOR4CR
BZ2LG9nB+Lrl/w+Fd4fEiHPQ8BqFV3kG8YWOmf6ky+P05XvGjbj7aN9ynDS7ezec
+o1+cCPoakH9R5NXhRDbcfcp3+/L22AtMXJhNN0riPAAeZfJ/4iT+KBUtyYaBUHM
VK8JQfQzL7nBYUM64pDN/BcJ0Gp/kDDzqHWgysWZ0IeRa9Zj4J37GpkDrbJ8Upyw
DUDJEbUJ7tAbLRSUa7qWJMgxSzstqKvpIMUg5xsh49CHXXl+G+cjGwxM5DqeLuNa
SJ3baLkZ7C4EL0wiZdSXRdfj/WbkqeZUqsbC2nrxY9i0ey4Tb7sOOou+9vUik+Vl
GBWhWpafKnZR+lLPPUVi/rC5y1b/SahBm2Hek2IF0UrPiYlO18Ff2kcJwe5ViiCb
uyozsFA8t4R1jegLGPQ/VpS6T1DeYs3mncRZqmcDmnJdkcOf8Nbo5O9uxhwLlh0X
Kcb/88lHO0C7k9JvRfoCPOOj3OzB5RhUKLFz1trVgwXnbgCcJ/1dsbHuhhkwuW55
xs20WQAxab50SMj9ISwtT5+V2p52C81KLnIzwr2WUjoy1ny62RJ+KVOSx/Fti2dh
S8iv61e7poMLNd/U6v8WPlwRhDsOrfqwS0kvQ3qEpi/KRDNgXiL0PtxP4YUVPM5E
++7yd7lZWyy3f1WUYdqLd8N/IIL8MZA/m9AgSd2K0+b999FUSh9Uo9uxTvZQmSLg
1i/hvFkgOHTqolsTfiG3inP6NEp9S0niny433yCit3lVEQ7CMRrhzl1t3SIiU3xt
/kD1J2KU9BQpzNLrDDvmgKCbs7s0rdTATOtJ1Wg4IHh1fyfibnaVhZizuZpOf+G0
cQuVmld6Ahi9ShiRLW03i7cfhEXU4zZNIComuswR1JBE+3C4Cq6+Qp+HrOmx5V85
gKnoBUiagFj2MPmiTBhbefdWcYg6OwPllUcoHafoXxgjqHJgB8bR0u0n7XH60Noj
3g1AqHISM+6NkvOSqxKymV4whbYKY9Z+f7YFbdYHTBkjWQdaJ+tlLkLfl/PV8tuC
CIt1Xox4VUE3KMeEIdZuxTuhpIUE/f5X4aLnkiAsP2N8MBzzWwhioNuCdXSeQIdQ
cxzHHLRivEgQNicQ4Sw56EsEDhpx6bbJ0WILK0ASjIvOCYFK4Wt1yLCw6W8+3VTJ
ULr1hYVMqTjehG4G059MwZ2oKbpEtNJwD3L/pRnO7wgkYgNVA8Cq6xbXcOJpcwK4
+P658dR+w5w+CqT/aCR2oWeuxRkX7H9+bXGhbunP48Eutt8fVU+vPPI2aQy23e/0
3bauImGSczxsgjGBAH0jNcGosBDvloYUXMPDuBC1R/ndGUfgYD77ZfjISMuGGIHc
U6u4Y4iEP40pE3RcmLDkFE5+v9hg//d1p55pzXhCdWibJgKdzEbZTGCrvw0qLdaP
dnbHpKP37RXWQ3ETAObsk1jdYwu2sfXBBarSc4f54WohbWPyP7N4HIkG1HpR+Vak
xjwhQUDfwM/IEqzW5Ssyr77DxO2RUp1/pd6YcXw0Y5P6HZdS6Cyu36fAxdsV1sU7
u/3h3u25uR59Qw06Dy8mpXd7jO7JCWle25AoDy8XvWSvXXfjfxnQzpGIJqNC1je6
rHmudmUwapd9+BF3nGyBKungeTH8yTZNqO626Hr+c7ZzpIsnbE+OP8CmSI+E6uWc
sdd8dkLWGFiDp87PWE4KvZslz3Af47hz3mBfDn3x/qhnyP3lEeGMHF1RPHHsirA/
8YZK4jR0lgOyoiENCMiLeSISXwIrd2IrDRdJCSMu7nDsdQjWssd8k6Jnt57h6I09
9ISWTi0dBsdKzw9QJu73LjiLdN0dUS9T0MvUyFCHBacHeJnOWwV7g5TR8PSgqnKf
r/MQGrOyuIXQr4Hep25r195ga7gi0dkjy8J9OsR9f9KT9rfLXBHcY2mO/VApYJe7
+1h93L6hAayBIG2V2pghssJVGUINnOuZrLZeHYpgrUipGeqh/Sp+4c8JQQjWGhph
teWK7Fo3aHpUlqp5xJhfGDeWvyKibX7lAjko2IeKKEyXYoLDQ4+pWlZzTq9uWu5M
0cwS6AHinvvE6cUeDZ5Vs4F8EbSiVaHiBLdSiHfHZHOOXJqRzJhN1oLQ1BjOBNBn
svUUgOfm2CtMhOSNTXJC1pWu8TPbItszJyIv8u8eoY1ee4mdvl7nRR2Z4HTRYllq
RHmp8PUPyhZtfe7H5ZkrxjBiucdx9iMODMw41noWoQkMdCJoiepC0bUMeZaroIEe
MQR6hu3SYbXMosQD6TtporSr2dX5q1dCHRPurchqIrl8vMrOBbjmJo4uVHMiPLhG
AlUXvb2Qp2oElPnB6LfPUF0lmI9QoDeyikPhnatlhezVf00/1Vn3iuMc2f0hxBQs
cYWAw2NKqIGxWN7UWdf0I/x+Ck+Gd9nCrhT+pr/GZPOOmiZoK8Hf/RYv1V2da3vb
7JgBx5Af3UO+qYGDYi7QZqecj9eRfrlKPN3Jeb8M2HIF1gepYl84hp7c6qAHl20/
e+1NnlgkaoRPzrdoTCSqO3CkIKjn3KW5ErpMJMGybB8N23sq9GoX+3tyGvaQ986R
BpOfQ4y8A8xjx3PKezFmz5l06B5ihTSvgfbfLflWLHlIgmnbS4OBST8y8SWVSZiL
wydWHPFvbdPofSjgBmO/3QKgerC2uNR3zdKXkY3Opc7vkpMvXQGz+D3hfkQ+9NCS
pzWrK5J4NWah3G68JxFnfx5K61vmINqzGYC86hjv1UR875wS6bXjxPG9CWmBrLT4
WJ7gHC+vu7fYaYlSEvhlNxj0UhxhjFt/68MEmwjhErWkxeefyXbNpB09rbRDispq
srgDwMTDTipXOrJvynnyEorvnUkTqLakzz7zC/VyQRxyEICS+FAdbNLKc+FniM2m
t/tGyJukXJWIZ8P2FW6ZqKIvlUmHspbIDaO7hMezQ6zJC2KPs8CI5/T8M/21ANvT
cVDpQdKyvStnSVsB/VeyUPsTa64U4/DVRFK6ZRGwo2nT6orHlaWK2RpiLWdaFRfk
aa5/UQ62V7rfuSUI1n/wMYvqbSh+w/g2joWmjADF+MeM5zeOpVCwqFBdiwWK+46W
eoQgCVcZs21Jm4q6OiNtes+/uv4NpMNHsM4mRBsB2jzgvCmumybqrWNDmZiv6Wr5
cauo4NSGpbBwNBOuPY9htYvT2O++6HzpBZ9CiwlJJ6tbBybCqHhI/XFkQw6tohG+
rrnuMGyMfmr/Fmj544sw8TigDCzGxvKAwBAGjh0KYF1/MyR26epWObTBNRyWdFUc
YPS/kvSqtkRNBK56CgcwRF2x1hPe4n0uNhMBzzBU9HjSMwBkLyU/hEuzk0YT9560
Nh0II55HmnJDat0Z5BUYF08e6m4jEPMHanPkvObJ3DvxYLlkkTtfN2+zU4fvFtkA
sPQIDj2Hs5HuO/S1WuOviHCfV2ZxlBh5ZtlviAU0kjExPKk5vBCzxjxGhEPXtUE3
QeRvkYxWtoakGRSp7mvIiFmSH1yzvu6WgoGTiDYvcZLcDVtPwTz8OM1PCK+gqb+a
ytMVAhR8HaBpggOOEJGW3T/I5t4j+p5UIra32IplqaTkR9WgGcRM/4eHIdZSsuV8
JpO/UQqha5afZd/3XYRT1phvBHZvtGrPXcSnatN/SWZ04q/IF9KHACzGXhedhAXj
oVBkKrHpGmDasETXVdcQZHgVurlIVPkoHF1ZTtNvS5Wfpu2mjQmZnF5KyTbOHS6i
8M5bfW2NqTKb12zd/0lFfWSNcAa9O5+0fnbhNBYOT81MjxeCWyFMVa8a0U7mdCRD
LcdqUWDxA0NpnZDE7h/aN2mMw6dGbtXPFnl7Zf0WTzzapsHsPRRhYAdolMDXIcbL
8/uIAc1vglf/GX/og+rQrzIFkyHtwvwUDpPUpi++RZrapKM1sWSBFZUvYOJE2+pX
QkwjSAzz9CPNkARuqOU4N1luZRggB7ouq5Pnkr3GB4qWlbWcjp8Sy4y+Vs/OHuSo
RFsmIRasdamL5K8OBMMOWwizoXxOjgrCrJNt74oiYrfGX4XIJjgTAac7z1cZCFb5
KZu78yYTrwQX5e2b8ySknKckzrS2ALAPovyxAvn8+sznX3L+qZZEmDqLiiyRiOhc
bCxClOJk18eF69b5sxjLMyYWNMbNEmAKbAOMGyyzSWZ+f4CigmXF0iRmWDSc1WPT
wItGDoNYtypYRB8ybKaaJSCrC4B8a/h2erkBTIG8K2g3h0zRwWH5SFtnkXgEWx1I
nS3cH1HnJi+G2++Nys+NlmJe8Rb84j90mU3SjcvpyQ6nAsIBowrIQkKvsMeVeUuD
hjbekC5HX1e37BgJIDKenTmVAM756wsI2evcBsEZHmQnNqg8H1JrPMmFglOqufyn
I/Meqn9zjU8lNZutXc2z3xODpO7vcoa1RfOKTvZk5NHN43sYhpsImJOMLZj9YRk7
WtqFSLjfdfu1+KtvjgABtFE/3Qs9HFp7E/a0upBRYQndrCjly/BirPvqlm2XufMq
xO5DYUzspBlM6B5/z/Qx6lK7DFPvVAli6QNL/fccf6ZxD3K1r2vQXzOFoI61UD2T
+Wxcak0jxdRU7pZMyApu8puYnTv0knK+B9OeyiLtPv6r5IFwm07ww4X0tpH1wmQT
Z42ZGiYrNHODOE7yQQzCW3Oe7rT/l1W9MAIIBzmOYTiUL/4Z0vnPF1cxtN6KNa7Z
cQTIpIJn5PW+5RghvOx1E4dIJ49llwXY4LNHEd8hpa31gakw6A/OY2FjVaY8vlv4
fjb9fsTnEEkrbTk3dqB8Q1j2x4+yVIx8VI9mFz3xsvNia+ZPBXo8YBscCapOWPAf
I60GaqYyAweFMT43VLPIxGw2TIc9YdS6atEwSSVK00fqcm2BQN+7P4hdK+y89Onj
xweez19qaYRnfBLI+apInLZiFuOBHixUbiurokimXPr8ybHc5W8FH0W21c/vgg7x
/3+rcQfruTN7gnZw7IUWu2TK5Mc3baLom4SLPXi4raKz9TV5prysrvUS+V40Lf03
Lk7NEFJiouMIzf2roikzpaEcF+TkdvSZcYTqHgwY6gMd+EMBZx5FCF2W7MXfLTeH
gbt7mf5X9Vqk/efICH+IWyKkt41AO1nfEH4TATOzNZiPIStCpFxTVhy92IYZzsRR
i24wHkH7631mmfZfUPC7CXXFdQMM+wlCUvBgQUNuFf+pYL9UxlvDdX5f4VimthCw
5roEuJLggp/zg7RfEnlSOBr5+CRsgooFp7rS76egLJluB69ZEoTUdNxGvOEsiuiG
ywySvd/ToKC/HaXlShCqS5CCotyPvVD+bBCpiUpMtDvUPpEwzNm7wQhJ+MOe7NT0
xFiudm/X7Hriop4ZFB+gLCNMG1cWX8/Hu9jHHCTfT54ju++aWoTd1UNkTibUN4L3
ZZd4Kf3tM5my209cWUFS0uy/SGasNP+4kTJbmXjAF+elEnK/O4GwyZzeOw6s2y4u
Pc7m6df2cKI9ncOLR7sg5IFYYUa0o7Hb8XwCaC/NMiXH98KFyhQ6rNsG8ztk/c2X
G0zalEQyuXh77hOBS/jtq9P5jZapiXu8FE9FK9mGeHLnTphnwDAyylOaTXLoMyEe
CWZWlwVuuL7CU5e9x20tlXixBALpWQemGcqV/O5SKh8dnh1ewVhSrqWkmz8Q1tJQ
toScbrS+wUhS19DVNSo43z0fwXHs04mw3Vhf5OyboFJVvdJb2edib+EQUKffyQG3
mbDLu468R27qGm1iUzXVb2Oo/aYYX+ZBwLprnpjtiaPZ41ff1niVXO2iLhMUpR64
K3aR20oXhG/HbvSrluQ9fMFqu88hvvfehU6Fa+sSP68+Wv1v3RKaQXqrtxpCc4ab
d5OKFHJD4DYp0i3dEqiXNwMekARLRd4INbVnNbdH/X+ZUi50aB8dsx0DDIcGcz1/
ffw1qzKK3NW7CtORTkZ9UNab1IeTusrZyMvP9iBjR0Q0skUKrycfwtXAUrzLinMu
gRPNXQ/ZiSXN1XY21xs1d+UJsjr6M/YKtRDNdxi5Z/L2llxUax4EQtsaaNM3mJw/
ZqEsRQ/NHyp0iZyGFzj/Z5+ouE8BQ4ayj89+42o3cNmunhyU7tz10jaucdth0b6K
6VuQoXmKC6bsT57jn3yF4oTl7DVf3GMlqB4Yzrm+3XoF3jg6s7y236L0XlGmO7uB
btiZpSEDfTKdanP54xODdlsbmpPcmDdTu0kZH4mHJ79VuWPv/xRlzSz7QvZ8lFmt
DijIhAO6EuHfcPf0M1y8BwnKJGp9h1UgotHiJqSKnOd/rBifhq+OWvepzwm/ia9D
AA5k/4esNl+yFDoFgylOAhBblruYDkbwrSZnrVp7r9qWnujTM77CrYw0LCCpoRB4
EvmMlJq4rY8fj4D98MiEqwr1A99BzyRKdVbNqUjsJ/D/N6Z8CKxssqhjq4BrVVrT
d7AtEPIEDWWMIlOWyc+jG5DjxVuXeGYyzMMGcxLaPtU38v8RAlyE2Q21YlLWvw+a
OwlBQe6L+058F35emSOxksOMvnGWFD+N7aPVhpmcILVezHc5+m99yu0kFqHnk+vY
DJ6eaOlQagDTk+3rXGAxmcIQ/qrAt/C/ptj9gcOwX0kNkEO6boM7NyqYa2dOOVPY
Bts2tWR9vh3c7SUnzh7mzwfJVzJK17jvOngHSE0pkL9eyDvt4m09zS20no0ehI/t
RDyEHBd5H05F1nKXwtZkLf9DehkhiT9L94oEIujKsxSuicXOCIMCl8HAcq458nzI
VFh9MFMX68gcBoOsNzZTXiksMEL1pGX7MiNTSgcHtBG2DCatezuncyHY5/d9zwHq
m7ZJwkiwkX0e3pVxPtblh1VzhG2kqRfHFtzMDGXni/OOT5dzmc1SzIxe0LNmWrOg
pvsmQNIpeSnMGxshBTrYCuHzGencO0L6CebfuqIsFqyt6Y68q3jTot2qt2PKgdJ4
YnNIP7suiN3NpgRJJCMSWoFpCI/l58K0TZNzokqLGdAFJTK4ECJIWPYBFqkDKPMw
WcvfMM4GWRRrYxxtmN3Q+krKwVneLsJFXQPsvsVzuNbThJbWPBI6fcHbsfP5tVm6
fNympzNMh8UJkCXF/V/tMXEPFr/KbCCbjxY5xNnSPNfH7w1SgAnqeHUPS5gzzvak
gA/eWlDEVdP8k1ydOySssXZbwacG9I5DHPgon9oD5yio8Ncl1JK5fUdJph4dTRYf
LFIZGgladKNs+k6u3TRxgR571DacoYmM+KrcbObS3yi0LS1swgZBO7TcoUfWg+HZ
+wPjO/Z9/AZ35+A8G1HfBE2APmXh3Uj+J2721phB9wF7GmGLOZ9vxuUStai3u5fq
MkNF6aqoodnWpBD+iZrRiQ==
`pragma protect end_protected
