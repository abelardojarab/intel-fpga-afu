`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BfXvw4ZUnUGyB7MD5UiBvFcWV50wrV0WLf+zhd3Z4cbifykTEQOwDSKBHsWnTE1K
GLLOCsTr0HmlXPze3Ud1+JxKYEnmIJz9rZk3BbbbNQ8x/ZEHu2uCZXEI1RJtwVKG
oKVzkGaqmowd1/bASexmd5lIx1IW+WvH1hQIGt196W0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2809888)
isRogiIEoS5lRqWE1h7BJW62q1Xah51tC80nUhd6iq/1ioGHGGcbNhMZf9h8nlKL
1QABeUB3CfyYh4FHWQ2RPFZrIeaLHqWcacBTZAU5X6WY7Smu2LjJaHyqSoHsZ/TM
QHycadYY2koF35JBwR3HzOU7zUiQ83kU/0fugTnRNQEZJzVh91BMOr+hArlugLOm
oO0w5/BFkyB164NqC4wyxxjqHlf7zS5qABwHu1rgHUZZKw1VdZr5JVWIMWqAXh+I
6+YWHfkb9Q4NSYCfxg31h4+CYL3JncRYgQlJk1l0N9xKohhbMygm//cohO/I+c2i
wTIWsWQ8hKzXApiY/IwxL8bBG+3dhDQKOkkHnVByivsoiLuPKhcrHkH25HxGgK5t
PJ/5Nwzi6hYMXzWuEjDEinsagEor20F9ox+McXZPJElQe0IOZ7KPIxDxaewtWvof
GyyQyXy/RVYzgEWW5FZh/oNXXKpao+HrxF8X+FPjpXpQok45zYdLWAZ3oimAVnqN
QfITCOxHSLUnjFbkHajoDQlxDFA+20khsPBJfa78uU5sjkCDRztvAJsFuQD4zqFg
FiLqyw81190lx8Jf2jEdIb0IDj+lK+lOumAZVIo94lhPogqu0Fs/BCD6rbD9Y34x
sf9hXhGlbaV9tKhp7VhgAenKg4CNOMly2pkpN2/HDMeh/mFPyavbbDKy8SKqns48
HzVtOnuI19Ajn2VgVjX98FW0AptvXwgI2hKGEzMOiUWeFKEW5blbO7z0KKmK5EgG
1FmwqE6QwZQilunsR9TpljPCuqdtx/9EZO6Dob+5bKIVYDkgw0Aeu7cuoFzrR85t
wc5ZKFl8DbdTA4baJ7Hki8cDgxo+mhN/Zz/pdAgxOfgAURxWU/RsTuictCajrepP
M1Iqirk6X3W/F6XcSw1O8X20GtKFQGorLAidDB0GIp9LkDPy6gS8bz6BZADafNBm
69ckIm5YcERZP8gDwBSOuRkzDFRUWJXo1I9EukcujGkwd/9GvZazk8ctq1zBmLdP
9QnsI0pQBuHqjjfnXknSqr3OmepxYvrtRqW1TxSRZIN/FQbrd8lsY1l+NoF6MCMh
V7cAy351ZCJ6ufOEwI5QdoBJfwYayoPoJQsVeqnZsSPrJRWA4uTPLrgkWbRa4O9F
CAkTgOWZcVCkYOYukY+q59yhz/aYHgkefjvcnyFg5MaeU6L5TCO3QAjbvCEbE9G1
IVxxDFvmGiwSI8z0/v+WgMeRR7FDypGffKjXnn2IUFBhM7lSPPRvUMnt8fUsDBxc
77aaTKdfVPNmJd0MZz5bxmAOSxhCPqPdBsxoll47P2hzCR5AMkvnyOD5j85DPnh+
Gajkq9Z+7DR0KKzCPx8+jNxO32Uv8jGz+84JHAszubtNqF+UKA3RytLMpL8E0ODk
j7okvtHQTZrn9RAlbnTfHUFkOJn88oID7Xfj5SJ/PKX09EkI0s+W4pgOdD2a0sgG
WNQ5xskj0HXUAv2HNWUfYC1v/Tz2q+VaWlX9AaDkAy7oECDJpAnXvE3hxPZdIjpZ
DaK7i/F6a95sKTKh1xzlM5xKuEvDC7YTPs2N4XQV3cPQtbSuWZi1IRhJv5ANFAJD
VNRFpX+qZGfef0tDRksZB7oDNAGXOHAJRjKjUIjnE7qHUaqHNUQlYvc23rMKksct
fyoeNxb2TXom+3PFaJAtzRuHPEcvF6llrMIDoEGA7rSTCL6z6jXst14Bxu7ebZX2
eoR2llkhf1FsGGtJ+ahq/+W1RFpO+TR4+gCiG612rrJOugFBuxvdRWlTtx6VY42X
gvbqSUfQvlVR8vScbM4ILTGowBuU6H6cCljS7fpJ9kIHtg7u6TYBskkuLT2DbV9z
l/vXwDmSNQeucdMqK/TW4TZosqJ07SEIjhlHxgWLAwIaHFZuIR2BH+LzViDJUiaH
muVth0WBLSoSkA0GdvIj47E0DXVHgQu8xB8+O9dzS1oTsvxQlfD3zqBeJWmkqL4p
cxFLuqwfuZhhIFNGROngsF73T/8nD80QK85ek6xw5K8410u7MPbbMUmQxP5ozDGs
1PCcAjQCaPPZ3+H7TCCQ+HuCU/gvVMqm5p+lfzIaYGT8a40ceCo/Ht6AULIEIMbf
jvJvpMogqlaXFMPgvJyQWPkXoN/UyM6e96ijLpQNoKM3yVuANJ9XEUPjJqAHm8QL
rxxiZE2dsdLHW6NdQSA1b1mdh2gAZ6wSIX4PABLQEcvvERtKoMdu5/4CUCiyjOj7
ztvfeO8jtzIQn3OQStIjJNcmFmeT1Hf2iHHSw3lRmQIvZW+oIwR8CdatdrWGxRMo
GSjQDFEHAQvjs/cTzuOevrEL+Kl7/ZSZjifmNbmxy+A5MRBvjgGpbeq+nKvAKWbB
eGxV82hMQFvBP9NWY+fK0S9b3CDfg4rkvKVgVOEl1fv39ncCz5LfwUKXxvov3/KD
aMA3vvs1wJFFR1KKsXjyWv/GDpYFT8XM+eVpwjXl/8l+Npt3g0Lbalna1xCGdq9a
eRjG9h5XRAq5sB0utvyx+E+8t101EtbgHGHcJIXPDKpyXaH6t3WuIZrk45PtU8QI
zwJFGg1cUMeKf8UYsT17/0iU5EM8FgNXlHq1nzrSr07w2Lg9sjrdv5FlpGR3T3ti
XIcCPm9F8toZhq3iwBRz9dH+GR+er5FGS4jkHEgZbfgCRQSlPLXskZ5ulzMm7Jnb
v6dA51xPC9r6lkTUXvNXUtCcaY1yR6Md3iPy+9gUyfgzlnfCMpQrPU17mdfu/rn4
BgB2xfd/moJYsRQfvEQq+MgtKxC2LyQFTL5/ZyHrmoQ5wvdcGj5Jn+SdZMe4RpBY
FwdE2PA+amCbt2wrJQHIdnZHPpr5M1YM8L5gQ5G/L9TO7+IxKxlqRgJ6YHaHCWKu
VuEsCf29rruQPdgTQm6qgwV5XSFzKA34cJ77hY3Lj6jOjVaJaazgaJWDViRrPkhn
mhWi+t68+TRNh0AGXORgL5JrcmG/r/hKiTMBUUku9bIUk33GccYjFiaS+F65sRRd
leB8lDWJPjNqmTGS6Jl2cHROUidpF9K0CWxsnv/nI1mRFF1L0fvoYQyKCdxsCkP7
okweDjcWmke8ECraLaj63KnnhFchS5Jypx0i07iBSbXekMtoU3aXwxQ6Iy1XkwS1
WDRKxFAuI7HTkMg22tfVMP5r3xiHzG3eo8M5tFIVzflDu+g8KVcumJDriL8xmGK3
zvHoHvR7zNDrBrsk8xuKUmbHC1FtUaWwXOPu37nxEtelmirmPCoNE9/iakDjuoZ9
8j5tF9QEMwSPUWaAEMIaxBDxhf0uVkhhaBGGL8rsnn6Ysw/+8khXA74+mf/KeATp
ZEo/GaC05DUycotojUvjXQCUDwEj1Lvp5Wak1RZ86yFf3KffYyY35pfkveiWFXr1
bw495PjX4JEmZQEf1t+cBumeBZMgtT3T7AKsJdVa4Jv91pntSuZZYdM2NaQjdETy
TV+S1z6eLVrkwuNHL5Pe1PyCJHGwMqGSNS8bkqZjR1GDzZeVmsZmiqckGpbw2bIO
wICfsRrhM5M3wXCzLTtx2OCaqaZfTywWpurRUbW03qntTIUO6j518Yh6J7lplbL/
CljU2/XlAo810dub/Xr0q8W4g2fOoNkd4ZAPFbncw6tDj8N5ws5zKOmWOKfzj0Ct
DARAKDmpN5b72n+lIE1tIAJ8knZwC8NWbxcCH0aBDnQojHqgaDrx6yLrh7w3XdPH
B1nTrQUlFFeHyqBpf0mpq8pZlqlPg0CtAeUDAd+kFEioeM51sK9agVw9paEZvSAS
I3+U9RmT+61aH8rgvQdGt7Aff+DjtJyQ7iajZIPQgsywLcuRJdV8vFz0IWFC0dnC
polRoc2mWjRPoXmuqOAq9ndN1RRp+75tQdmYGkozllV4DYxuzKvzkaiLQAhpJOMz
55Cgs+8tN2U3wvY8Smy7Ceji45Rg8WXz/5l9F6uSGmZYDRPDF/VZxTs/t5pn0zk+
fS/AZAK7fKHD6SevQ3pUQQcrCog/2T4hmEYopMzzpBzBg2/LdIE84C6DI9B2DAOr
08Qty64qoevA1Ydk5rHquog0KELyLhWxkOt98s7uU2gwVAl2OTTy/gMwIfDV6FYO
cr/sDoHrhQSvrSB9sH2idBbY2zAcNGztTME/HOTJUnr+gqfyoYdJeQ63wIywLE21
prtnIYk0Qdy1uwlpPz9Zu+CCYmUowoTw5apYsWLzfiLGzg5183yxifOkyiXzA+UW
rcZf95jZXVbzHXj+HF2A2PJXTsgeaRA1LxO4yj7KmCngUkBt2n1zXizY0WnIpjo9
NpW6Zh/qQLW9NC7cUghS8wJXGX1sagr0iTpROlQW0qrkoF8bpbyILgcY6yuIlNUP
W4+Fy1kJOxjNDU8EQge2lDl0p8w6iVvAtdbqo2dTK1LVcShG5kKcGf8p8CVFG/MV
HlqesEvis6xgDPw+JKZaaKcA1a3ghGj3LJFmulvcCOtOehD263lv5UUKDaHz9F0b
/7lu+barRYCcrDjKsnwGubvUIWcgK2Put6QG5vzXBIw7+I3TcdK+3mWHkU5mfrEO
dXD8LcFFjUdC0NFMBEb1mFQfUHnXKxa/t+TKg0tunwzgcFCQC5sRwdGGA34syblf
eo1Xe4O19XJa1C18kLPktNqjdI/hbDkJ4KU/o0hZ45ci0c5ttE93EWrsl43CZPsF
O8bj+/EuJjusbW9LrnR33fsYIBTbbur01/4JxrDhKlcy9QOVQxz9xKnJ1pU+Ma5D
LlNVkFYRY8nkwD5IA3MJT2KOF/jU+SxT/Z/eHwsqjvYyw5Hlp6DCJ3FiSuunN7Fs
YkJAqgmaeZof1mLDhj62f/TKNMI4kW43jVh1GEVYyMHIIfOiH3fLGf1WXjFcnkyH
mqAzYNMcRoBdiXObs4/m5AFokVJuSIUCGIzoDi2L0k9h3tpubzpMeHGAoOjnpLq8
5aLlAlc0hojpBwobi3Z3JGMqZPIbvtKJEK6lbNx4A04QqUJltQZMSllBGWbBHsg/
0ec+I7RmJOloRBK2hRRSYeGK0rGUxJjVTT3WQ8BhEKem9bYFsw1ujS9Q3v9lTfca
EXpaNmUDpuxAzzmS1UZD+9PJ88IkRR/Sav9dU0o3QJsgArMOtuHRNzVlgLDzY/Fo
S58DYwaABLhqlZ0UYPA/10c9lrPG7UANmaeuCKYsDMOtPSxditvWEB0HIVwN5AW4
uSEwtZ0BCGfMrHW4IWK6QUqUe933kqXHPY+A1/CkCSp1i2R3nHpq0xQdsTQZOb3N
WQdykgXlTvc4P80LZu5Ex1e+JMiPHLN/wB1lb858owKUncPv84Y0NKMo9bWslLzO
6r+o9b4rEJiZbvtI63NBvy5AGFTS/vDx7AmFwb1xKTE8DNLXTBszdJAvuEnNCVhC
HMm79hkhKhxMojQ0I3wkJpFHCd9IorR+9zg97+N0Tuf4hpUdNUG6dozC1b0Fsomf
MFlz1cql9Mfs0BiEzDsGKw9KU2JQ6SnS1xgWcNTFeaQxW1eya4E6lmxU+1fjzg//
F91WLTU6VWnh+GHdDGgNwZm/l8TrfIwyZgpEGy+YQT4BRC+IY2Ev1BgZo9DVeR8D
HHfgTDChz1DSsyMPFTThHWBF1oosWWZYSSIyDYN+a6rsFqWMFN63Gttjn4lwLBne
HsHOE937n2VVtJO46JOKNy5aVDJyHSNboEO/TrzzWTG2qNMR1+OKTdn3gX+MP1t+
h3UWwQ2HaADFU4Loq4RuosMyz/F2Iacahm/rnKc4voCzslqUN+EhYMkSBp9OvaOy
Fn9ZPRnUvWZQ+f7Qoq403pcGm8sxkiMHadc193NGvnX8WMqL3xHA+00hBTHfCYSB
iBI2eEfmH6EpCJiA5Ri81HTFJCDiKSMxSlppeRUClKlDr2VTJfPmt5BtOCMOSX1C
U7rbjCqa/g8MCkUH8vZHAjW0mWeVx0StxSYUwg8FRG0SNuz+qXA3l1o3e7QZs2cU
MpDPzzcG3gcU4Ih9/PD4hDXXDFBMckduzV/60YYMbCdnUt/OiMQz6BKEJOozQdef
ihngulwSEvOUmeV6VmavYsMv9NO3X5cHhkPuvHzUS3cO1LjMD3SpLjTkJ7Fo7md6
zfc6tAjLRkRHVP6fYGywhGUd4qSdsWNzXwrcHdVZVjs+JqlKuBpyE5C9MgKuspO+
mrdvkHGXYpI04ProiXpzKdjUsvQsbgPO1oOODlCNpZQD7McRLnDudtLATDEEYZsM
oKBjjnulvLXG/0XYUk91rBzl+MK86DtQcdxjYIVphEgB+eF8oNNoSHlomoLLE7XN
QI/UCU+3SSjufSAH3RUE+IulLxFydFXUriKjABlUtdGiKIANwim8r+61uuOpRU+T
t2chG7wUiB4e1b6MkVAmDQiy1Uz+VyAnsUEqRAHrBHmAMvKxru/tuKIa8PpMdk/n
IIIL4Ew1ySSy7HQsLcH+BOVbjWtCmW+Lqfu64ljJDPJypBiYfu8k6D5l+sKfp7KE
WW1a4L6BInR9RWGGONNeFcNfcpKOaqQ4LYdEUoNLViXI9OrkDmIKDCPRBwkse9oU
FcczKxzFwLRi5x+SRLlFWgyuDkIIGLZLqIkhahf0IgLI60uLdoMbcgTjjLXpTzF8
zbxPLUP/KSzg6MnawM7RtWQKIX7VTGX2iifqLQVXcmoYNobiKINaanyU6Qdu1W9f
483/SjsWvdq9HS4Z7WGOGTzjfBLnBo5MolfYqOm5qE1RikmLJT/mRfDe7mJOV0QQ
ittsmw7wmOivs4xap8DOTg2vAW27w3OnqTIiLbzWYfBCOW3Gjgr80dX0/OttxRHO
8oL5oH/OofYf2M1qqf3tmpjkNDRXadbnj2BDHs4BXRGhkqsdv8s5ae+GqN+eGaoP
gqIcWIsKC80c4kxf/2KQjQ3JiQ4y4q5MN8r+ux359wX+WGfQrwCN8rH8Fe9EkDgb
nNWHg7jw2tNuBZCHpdznfUPshYRsBk8pU0WGUnqiTlp5Siwx+aSuF5BgIr1ZaFkl
x0EuVYbwRX8PQnjajFu38B8N4BM3T8g49DkJb00R8vKQBoQ2OboqEywpqGQ7LOOF
pU/fGEpzBsExBFdp+4kimBUpku9Hkt9q+FvBxEVSN7GX0ckCCcCk+Y3rIPdMq8xR
xwz6CTh4L/C8IUEXpfpZKVMxPm2KGkq2xrSWTVkMt2TuVhcdj9WymXpw+eXIpNjo
qkbE0EA/OvYCL9UbbUHllqnpXoUD9KFMQUiKGTlRzPnKi5iJCOAP1+AEVZ+TGCiJ
wtSfGeFa3sIFi3xLMf+KYlQdBCN03H0fxcSEO4d8UWXd5Hc3T65qaF/t6/VpoP02
jMRt2GFGTY+ujUs9jK4Grj93DgrNQZzIXeQ/ZvupbppIGA5HQ+hd3w5AAEvw/LLB
De4PQSF7vufLbygBARy9YUvTDBVWoz1Cg7rEdtsynFDh35ioZ/2zYBfy1h+WvJSZ
N9bfQ+jHbWLucKfbqsxyIEqwYE3VVoRyYIgpTfCTvVorbYO2584GJhKV5mnrf/Fy
iWkgmkeImhuUxa7wCYL40mSH1QqzyRNAuFNKDai00OHzEYB81D+A8ZpgC0iG+gIB
GQkvXmy1mXiaXb4P5ZkDIvK5LW2W/GYoeIAQB3EbCqTpRP7Fc5+GQE3tOeES/mp0
8fWCQ3tcoU7e0VT/VA1xfbhnR7H3ERzaTFyDvijDjzDTp43CWvEjne/xfbEZF/h/
hqpIEG1TRAzWa/YghogcMGu3hUnoSaJtv/9f8O2WRVgb3hyRx6FX4u3INaWu5oa+
KSdt9zwwLZ0doWMkpIhKFdv4rMwm1kvLbmQCX92lbj4N70EQaHVlt57LVSOF1Cq2
QAoru2NrxWInntpoSDs3wkiIlZrnXo/eWoDSvatnEUOlQGqKqIt545R+IS3WrhGt
7E+XP02lSwlIkx2Wjk9wVwDaYnwTM8kSxjAvauSIYKdaEMoWsi5ci4jFDc5CMdPc
G602lJdnNzkWCNk4VzE6H66XWfqnF6rX+UOBCsWa2dCZJg6p3zIGBj2FjFPn5xPk
0IkOzsT3phfjjmqNV3ZAOMHUJVEAUwA2TXnO/5O9i0vg6EnemPxkFOPVP/tchWaU
rtr4h6KvxiZrU7UBOlUEULlz8P3mxobM77RJkd9yfykCk+ogC/peORDy0r83oelA
XsszzTM2W63HJGJu1gBtTvjy6DjWAnrHH3mjiveZzDoR6aVRK06avJukGYBjKb6H
UITFpgB3GhDJ6CP9r2+X1AH/orf63+6txRTACAkpDfMtLA+VQE5oGSgYDcI//cjV
QbPDVV5XutJS6k+XpShsU/WBlqM9+zlN5pQs+6AHSoxwRCjs7D2LqwoKXT4Dr6l0
WQf1XwqKSXh2mmO7DFT6SJ5ANO1Seam2VTGIGmFPNqgiHiSl/tefiX3gEUZx2LZe
FRwyLSLHSW80Ey5IrQBzWG7KcIfxSrLwZYnkqk8nu+p57Ts11oljGHKY/5rxhvDS
DKjUs+a224c3tUBp4DsZXoMAJDLL76VJ4qajCfymGTw7Q3/ZuhicH4H9CP6j49rf
TxOwcCUH6FLntx6RB57YeKArA3DPdZVA9bR3nQsZUDpQGB/IS4PJmqH8T5vhSa68
E4wuemTGH1QwX5RsG8B//EVPFtKTLx/Icbecg5aWmGEfjRpEWol+9OETvlfXwxlv
fRsZpUiWGqFP4yfeQh7YSATKYRyHZUUL979ozyca/Oy9EH0RGftIsS3FFDAIziJs
tVytXCcOf6HMNa2DPbzTNUvxX8YqOnh8ISvKAe6yzsXWcOhoFhBlgl233xQLkwUu
506KsBZ/w5eX3AY2NbyUdyGM6phM1Gb8aZNqzoJ2WY4EwYAhw+SZBIEBo9wky5ow
GJcEUVTmEwGETIhMk8PJoKYRL6aoJwJ5XcvCu+PgmS+651DpLDmz7paZJVpDy7Or
ybN+Ubxs6EjXQig7N4pndAiXHfsjWjhGvk+1fGkCxf0+Ai501W7FroPLRWAa0bzh
8Cj4PD3VJkhLflJ0gHJc2XaLocekZqsAGIe215jJncL9eAQxH/WcsCQfrVCCw/ru
Jro4+TJ/DYoN/DQOzVQE2V06Ppjrrg+ynbzcffIAW3V0f4bEZEIVx5NFmDJUyGcz
iW6/EIZW68Wnq1m41/Vc3TYapWlXTzsE8SBUtOpaLtiYXkn3VSZeLFQb5ue34i80
lGYQBbr2extGr2rgEgV2vJepqIQ3NGkEINHT7PwIbAgQ5+O9HLtiqy5rHWItLus4
H1OjzSKbux4xnBBbsoyeHMPKxzb5MXNatPhmo47E356HzTwCMEgVKGw2tUBAjzKw
irBLFk5y59WhCJEibyheEWG/wnCgyuSrC+5YG/pCgk2nTWw74IX68yLhu42HQu9y
mAOAAINqHN1BW7mHJaKgB8hPDDzuVMJHNvnmYlBqZ+eW6AK67n02WtjmQBUjn/1J
Ld4utdH/HhMX2eC0pjOaNLUy1IE/g0l0jBLKrnuSFsz53HqS+SRDrWHQVGFvssf7
xINss+PdRM88bCszwI4VujhoFKsJr3fZB2K73ZlgMbPK697QQCICRL/uyxpWP4co
TnkhjkBbD5kqibX0oBXM+FguOU+aAM+KMRehQwz0uKB1IUqbwET5WIneQF2aLEbR
GkbkJjkgLO6UVB220O+8VTHmOAhLkMA7GAMxAassxZTLMnRuGKqPWwwAttgqmDa5
nLt8NKlvpJk45Sqcb9JEqMHabgi/hFo4v4o7lVX3cxcmCx8vy7ncdCUkNiNwDlau
IexG7nlmkSCjX5VnmzZY3h1IWSFPeP6rEzSwN+eBpTDk4iT42wz390sYOlEML6RF
c1chpqnyvtvANDYEU4IEy/V5YJaxZAmvhahzQpHrY0egnJDV2WwKSsjCrddgAlxY
d6lSFIwC8dkmogHKVZo9UGjTL/KGbQHclVZPeQsPedPpPYQH44Jy0xX4uwPHzpa/
q8zCmR1SdNy02pNaduyYme6+X47chLkLovxV2YqXj3c+HrN88OkqqXipjsy9SCyC
VdXHEiIiE/LFe+cH4c18YYtrZni05XZm50Lrf5aczAL/mYbm+n5DxlrbWOy8HPWp
6r1ufADvtn/JbIgaGvDhvpfQwb7TwCBKPBR08R+QlrLYdlWlJtbiL20z0XW21OOw
OBLQLnAoQeECohJZ/9g/Y9R4b2qGp44IrG84zeR0BWFXiSZ3muKOXZnTHz/muSIC
yS+N4QhjoVAfx0u4XJxOc5mK9rHYSMNE1Cb/uwj1LcqgSg+cAhK85J9JPWBdS6iV
/Ovdye7wXhEwIMTpcOHVlMFuZFlCaT9J3IMOSyIf65t+Ql5otGfTY6lVPEugXgIn
fHVGufwiEupDLA0zmxUiqBfKLFhnRe8rtZ1Fluqr8MLhXbcGQOKZ5sO5GWfoHBvF
U7o9oPqZRJfx/1+7AvYLpvMW9aJRMS0bmhvqOIrX4Zqza92X3m2rOhq3oEnyEjnk
xSCJWruNsCRLqpvEZ2mp0N0Ep6B/YAVCl4OW5XPWwbgxxDGGa5lXr5p3AuWZkMfy
+k4r1cDDctkte1QU2hotbW4HU3asxtW5ugGN6Zit8flIp4hPsI0gkwfm9XhKB4sS
n54XE2TT24Oo8n26FZzv/uNQNXzyRlNDuNVx9f2m/Lhijx8JQI04Ecu/PZUhajfL
onGswqhJcb8wvIAkCS19xUFNS3GjVEDS0CW5jJpO+nRr0xHuAgPnGGI35bS1n4Cq
/pVHaMvyBytU7m/h23XskTz1/VxsNzMM17kOJdKiy+p9xn8v8VYUV4rtk4ah6tfH
iLeOidLAe9xkCLXn2o5a/oFD/5naaV2I741tWxh4ObfTzv60JT4SxchEXvpU/zV6
iN4Zrj6+lbMsQMHGrYSh43o5vqpJB8PyHukLVHCXy4u3OjoYIyun1JqiHAC/Vt5P
NvO6q7dClxBmObawbkvh1oOZKYiNWZGwXFz5uR20/1F3Il7kyQrcVot24/z32FZy
P0eDHJjSfVHgJ4qd99JIiOAFNgwqPVPfm/Z0GIkmlRzvmY3fy6xUI2PBh+t6kcCe
RLKnAEfE8FIL2XF4n4pZB5AlXnuBSMSRJIJ4VAvSvq3O9iHA/h38Dono8hFmLqiC
YvptxCDqnU4wvhHjjaAvwRg1a8EZfQsl6NFuOTXQlJJTPuMsxRLjakoAbLXzW2JP
jyhjYWs0UExnXnUnQrd3482Wl3lfCmwA8RM6koShEgrZkSoJn6oX8WyLC50nhMZc
DtLuOhDjJ9HWNEhiBASfX6LJaaj/+F66MzcdLzrSA4ikYjvBGhKKGlnZhomCUcU7
QYfjrlD2StF3uS1QgMnuRG42fwbHs1q/kbC3wGcy8tJOJJojfQC+Vb/1hzCh/Zhu
yolvu4eYRcI8Ne0IEyquxy6xEQuoYpwLyHrH6PXu1XMRS2aTZywHL+c1HNCleM2R
3YELfFlhlUHOI+CHxG2vWF0ab+Y8WqZ7QJb9eKdfWmUbre69IeNRRhGSz3Jda9TB
GgmfjAf72AvEZnXuhqwH4hDc7WcsJsVFgKK7VVCRRKCBDTwOGm4ebvqdgf3XJYlt
uOQOLfyXKSiqL8P3qPJI2HJxEjXCgZfMTwqNCpVu0OGrQmO3/cnoiacg29DC+Po5
jx5jIruZ5Y+OmCtx0izUTF4yZzX9dpK/5db6CCtRd/cBiOrwaHrsTXcEp8KuXNcA
sVGUtUpowLzmL+CLZR8fFFCgjyCqzyCuE7AwSscV6D34kfmGyrLTxgluaNFdVoE2
J9xI7RqQ8FCw+pIpwOnlXeeCas8dmSirXBUJloZ2p6uFrupm5MHUK/YRIYRJJRZz
BwA6yDoTSDJ39ejqHpZcoYHpHCCk4vBBcMLm9WPJrywBmf4L7KpPnw1jMiJLJspl
hNfiawPOyEE99SLN2LtS5/XqOtkbKYEsvfYJvte6H6mQNa9cw4H0/VeGptOwkNoE
jPxMIM+YiajrK8vML18NdvstHc5ssxYI1Vaw5E5TUWVFXRx7hajvhFNv8QdqUvUg
ZSdt65ekiKy6z0bTzpnSC5w848hRCHHdtdCIJUfHAtDWyJ7BaqKBzrNdiRLRkvrk
8TB/i98aqlL/rqzTbsDnX8pKYC6sFJEYEIC/rHl/cQKT0jMS/VKSXw2USNFpOqny
3J4WzpiSkwLYdpSokCMVPtjaq18N3boVjkHvZvv7RnsSGs6C/dzVPGp3OFUP/zH6
ulM62lnOef5nBZUjwiEX2jSrLJhhzrCU4Nuc/VshYeNEJXxAqh3D+3KtxD/+W2aI
0arSPS05xDWc8QtaRHWkt7AfCAaKlTpn+xKIepBtK8EcV0VlIudPw1wnJWPHO0lT
cQiUDHU9H+GxLV/q2RP6g7SfP3Gs/F6YHUFY+w29RuEIDIaT7DRizfSFXdXoZyl7
ZOxHktlOWU0+OuhXmIDRIoxjv6SiAZd0uvpSDxp16Iw99MNEEGvvl/hgIQzryfQ/
ZMgs7RShMMhWAq+Foh0IPk5SdGgQrNSd7qDu3OliFudoAVYB+unFwhgSbVfFHvjq
zLAC/ZuYY7NKHJYFg93jZGZ8+i4I3yL+EGgMTPg+AHPbSzqtagWnKJWFl2ZpjQ4+
t63CVTCvf8Yb6yDk4oNwAouCmuELQhhie2Z2JH47GM62ySJTw1SGVOYMnrBUY/ih
Trw0RIrYTSTtu3HxL1wI1KWX+zdr1J5AgdbMPNGp8W+DBh3OmJYUK7rvRJbn4V5h
Zksniq8LVKWSpJJbC8nQhqdKD4HOvCXdDOIMG6zLJrxj9olXSKceMNAVu+dxMutf
vOKHcgFn1YydrvMhOTmHr2WJLj4YmCsNneHef80AirRQDBC+FJkI2Ibw/6kE+k+0
AO/U6xoAx4zLWdj19GfGpRTfX2nYSnfyncfnR2BegGB/Mc82ToHb0RkWi3VZfouO
2n9cV8Fv76vjNqPmqXAauPrIcxG46XXQCelao+S4tAIHUoYMAkyxX5vmEk86g5ID
AiyV+wzIbJibiSjetYz9iDhHbMLaJ9ztP6rmi2y2PooBri3gvd9ohgiwZ7K6JggI
e2f+ilIDaw9HFnlS1HB09wQsMV7z2gGaoGPT0p2fGNfsaKDhpa6T/hIma7BZqZ1U
yZMO/de1fobveKXlgiH89m9aftDv1b35F9+6Sreq2CPyxhKozKdgv7AoV73elK48
el39y4+TQ3LO2U5DCLkUI2RUNWkTL8N+RB+UOdoECTd+sTKLHCVnR+KjusQLPYdv
aH67HcOQn7pRXmaWhQh7YKow3yBWmv0mF0SszXQmOUIhlASJSyC/OxoELvN+0PA6
hpsMnoPpGGj26cn0njnh1l9qEgTxZB+u4v+uv16MOKoZhVMCBx7+lPOSpJz6RZvu
tY5UNpjWm2p6mtmXl/66Bl04TOuM8+g4hkRR4J47+XQ+eHA9dgWTThv9GfO3NY1w
aMNvjkqSnTBo+pusi9GraV62gam95E0L/d8HPxEmbAa6d/0pyNGumJTaHZz+OJ0n
vUxFma5o9VDicRLRevNqSrKQq/d6MEkenCt9S2BkAosYYIXytoGhyusSLYotOEWy
HfP9NtUVy3m0AydOH5cWRxGayj/SEjNzrLpotIhT07Q2OrKZfy0WwFSBPtuBnjhP
uercW/yS71Rt3nbVBQx4LseclekS98pyHX6uFgWDF3+f4jKZFdIqh+llhqDYa/AQ
CS5Yf3CPLFvLmc4BquUpr/+EUpzogPS+PSK2Vi39DURqlnbaTspuCwVAj0yTYynH
UMTSvFjHc4k2BR5bBOPrBM1T0reknT8sMJQyvnmFSqa7OQNCim6zgRfAsZQcAK7D
M5h4+InnnVLlLoMq0njA+DLzPporXtFibvdImaj9M86RG8FpslKupYnlXdYAS1iM
aa/yOqMJg9b1gcA2Ytan0h6gcVTucEEWdRyFFjmymWvq622qks9iWxHVM96yK/8+
/tuwFDaeG9xpngtzZOg+S5efJN1lRfcWU0V16wkLcYHFld0ewGKspiklGxnh1Qy5
C6isEFwFqNq+H0P1izlY5qFly0JWK/dPJZPeOW4c8sPZyqpQV4YJEDAlUq/SimRC
m3ioajxNybCyl265XMygxejZYxzOG4K2MzDhASWIIbmUIARye5MahDCOxrGL3teD
10Duu7hT5kLiTXBfdWf+kn6eP5PnLRciO1VeCoICBG48B/eU2pQKWw4ZwIoWqnq3
0u0Octux3GHZ1yDDb5EmC6FF92ePIFaPktoQ2e7dWnUi3jm2CEw+28KuUG3pNMPc
7g/YOFlGqn1sy7H3yWYXQ7W0v6UXgFDPX6vzGkCiZVg/8IH/QcDptnFQ8VMS1jay
EFjvvAk3bx229f5+uiaCWuAc8hwaTGVDZ/UM8oN5YWN5sQ1CoZwJK6BA4u4UImkG
QV0+jzLJO91JYIzLs7dXTAQrxvmLEGBx9UKMJORkwDUTVxqY75ioLAn3PPHyixB/
22y9z/pdfRsFds4Us1cecNsqSIQsPemqDHMnxXmZOQj7/gZzoyLE5y9+VXE40wyK
dah9NXbtBf2RrQB8gY5/FxQdWpmlytChI9CO1cm0Mi1xgpbvV+52xCA2XIAFIF6g
4hRiyULNKoaCeWu19RIYa8bwL9cU3Zj5prBgOrWJyUoz3nxGTgIqZa39UgomoKqd
mzAyg/30zZVCUtr6y5wHLMmaNYYXDxIiVqHOXdI8dxxA/Nsfp9OZY5Pnbih7wLHv
rAS/cm5lfvCuLS5hjF1xKQ8GFB6ktlu+UW5D91zdySQhP2lcNWRhrDhFsBVJmatb
yv1AEdZANypGLbzEtavRhXEIoeArtQwKxETLO3njVn1kBIh7m9Ay5a5zkTdGdOzl
BS9NvtChJUkmtTQghWo/HUtDknXQ96QUIP5JLi3RlCdUkjWEo8vyaJIHJWOFARg6
xn9cKUSqAvrw8C6qKjNKClRVe3ZD0tbNIB2Z8jreVCXMZxCVQKZEzCS+F8ZVDymu
nFU88y9e+8s8AgT0a9gi5PxPC+aOOCgF9fACf/hgn86xOUSdp4NBp+QhRWA4lupC
Rlyr+HjDFLoxCrF5zkB6K0RA9KEgwoRHIe9FNFBaSVXGqQM1gwJ0xvyfowmQYneb
7v9MMkC4IN+UY49goVguEgWU7CBywf1iE16MWJS8P/XzWMe0T6BZHC9bgxUoCv4n
QMNT7zhdDVmQP0HMrnyeh9BnBMuXx7VsXDEy4MK3541lwNnwPoSCWQF3MhklFWzu
qKrgAGh9LtVxbdpwr/AxAqmbcOFnfkiNNbp17BLt3KnIKshWYFyUOx7dl+mCGFQX
2+ZrVHO+HmgrmlILyBe4r+LeLzKhIpIEJvuYDPLBAY+9DgrCpft961dbuAqL0IKP
y4y4I13Bx/oe7tv8mrizHhVzXY4UTdXnwRlUg09qHYSs0Eu14QiBbbOv1N6WIJSB
XE1Pqzxhc/oLyS/2GWnI/76jPL5j/B5xLJjimTFh5HGmyUrkgPlXp1XIr4juXD/L
8XMz6ct8Hfvd2L0SA+rUvdjzXerUMxjPWo5uT2g+jxQ7P5fdTwBqZpcEyqnOLJnp
TaL+WwlcFSM3MGEnF6iTwUd3DVWlkTH+/m0rDFTSJuvTXjeFIp7tRmeFIAwlWWJQ
Hef5PsUFv1lA33IQEzr9m9kAUp26J4NHqlDhCbZ8lERsI1buIftrPX1Kme7kwCK1
nwnOqpxCe7m4hbOgi+X82MzjIXO0JXPiTqK7bctyD8T/k1B1TEbckCV4z3OHvlTy
5zG6lUAHCjB28qrwwSHrI23+8Cepa16JPnuvwyq89GgHhXK3sWo0PEShlD4YTOL2
JGzjNq+6RatPdoudhoXk1rdrNNmNX7lHtZwVzbUxq7V75ugBE0lVP8jmdfAfZAGi
rpx4Vk7UscJpDvOQQxmYC2qUXIhrwurFmH5VdajwdUhHwZtMvCuNn/AXTgTknEVz
1tjz4VpGSOBWi9T7/gS2H7CraeJ2HdweHAPHGRVZOMhs7MI4H5SNqxpZ0rc0bRLK
aHutaG21BeWl42dJTd0+0nVncWhAMuvqnoMxWNWD+toEt96AmIPJ9S7lp1vxMKDe
PLQlxq+qKPxnN8RHV7m/22uBp+dY677HNN7KKRSABi/2P4R31tOZB+1UCm/8vHXC
saWbWYpEkQZmp2ql7F15WI1EaPcpo8mW0cX7ggbcK+z3j4Q58IIpGhDM250Zzps3
21CNx6htN4fXoe23mOjrbG9/PM4D5hoWC9XktxDmlUzxsgbnAY/DAeonSIMY9ZCO
hOmVbpSG/zArY2+NUlxS+eUf810+ECXv/EZ88N4W3aYl3HCBf9MDnufb+WIbbFBM
jpPvFqVFeMkhqnRNnsoAmK6+i3wsIsHciYt/A4u5I65SikZA4UaPezSSkOKlCXuL
MII69bxJJhQJSnT2va/oB6LSBPXsgtASSn9XNmqGPIqrtdGV9ccOo1+wzl3NFbz5
Q1E7mnfQb9Zz/ys6E49H93vq+B/+qvcJU0cKQBPVx7WdBxcFKZqcFPh47s6BXjB2
xNHviy5VDb5NjzBZ1ayQj+MEzgSx+kvK0MoryuuUI/spbJBZWeBOssi/zsWoXWSY
q/+I+Z5Hc6ugcYl+Ajn5mPd8crBVaBWIU1gU4jX8NfwgX+/MBGOU06QYcAmr549d
A9wDSOF4H2XZTThDbyka1/YTshex6R0qs7sMu/ofMIdkWKv9YsdrfRdNfy3GStbQ
i5vB0tzXwSUTlXuNvOs7udynM8maNaG3bZPQQjlF3cbWWy86MBv2tbhP0bnfYpkS
W3+Tlg/ix6oGUjtgSacPq8xgCNcZmwVbl/hfwNK13jU1OHibuY75hOljzGwLudj5
8Z/pd+xgokOH3GxfjbT6gJ2Ljk6w3TGNhEW1Dq3eDdI44EWOY80bfABgsqOsg1XU
9ZfgzcG/ul4cTJhmoR9Ap/+6e7bI7WnybSzz9BCMRMZZuAXZwrQ3eYsiH7P/ktSG
Kc0lUBirdxTeAsJ/HYJsYjmN0d+Kl45XQUrmEHpMlAwNWsoW8SWrg/HQEXgt/mwZ
nUCJFGp/sTSIFw0b1/fqyfaV87+F/GoeiaFsuumjhWK+04XZZPzcb/U9D0H0Ow9Y
y6Uca0ouVVsAhTq2S/QCyTPI6hyLo6ipvc3mMwz+jyR0slZBAzoBwb1N3nseo2n9
RqloLDtOeJVXtyb+kwLWmYXYSPcIGLQRdpBKyx3wGYZShobGp3hcVZ3FZ7JxxmNx
VlUJQB71zpDqPs/uUoNoGNSB7P514SOzCP+R5EWXDjR1csD0DYR5nc/e8mrWPdqH
or2IvVxntSEwEnMgO95nnVr+hdq1ov+bIj8P2eHUJjAzY9C7djJq20S77UcpK/Gp
a9Bs4inFgpAQa1gfgXZmZn79Pc8m7MNSZpzGqQqX38HId7CPHB0lKkUEn+i7y3ec
fSrmoLTvr6YPQpCc2x09sY9WuO/6lzGCO+TfQSXF3qbK/lu2RdG9qmj0lT6hu8g/
AgN8wj2omveyBhNvgos0kHh24BXsjHR260pUlF8zKSt+DuHKLeeER+s7h6/3eFex
+LcgKNHkodsXWUQV6WG1xvsCVN8q7x8cOMK1c5y9Ja3/0O6yy2w/D9h4zUy1pegH
0i+5wk7rVtgYFiql80aFc+YhQvAMOJsoX1kpDf72pcY6DhPmYoDakJbx70njGxGF
JHLkLRMSaUrsbzSxJDCncN1ObC3FrkPXXyMsX936nuE3nSHJJrxaKfLNigqp3QPa
L9antaKUmzlzFu2Y4WBBshizBdy5WRuiSaEgOeXPVF+2rwXgHZ0tI3ASgX/r26UA
E+byAb2nU9bXCmYmN4eXcaHJPvmD8cNlyf/LBnRDlrwOcDW5T4U/uaGCmLyAefEH
AI79o1kQZLYuuXAWPWwKHY/BbBgu0xnnzLa61GlZeyhTKHYVuPL3NIhVdK8UpJav
gZkWpj0Y75wwDsPfzbLIhk4ST+9EzrPL7pgn9ZFJ69uoyEIIWEUCMyG8rygc8COd
tRZO8HFAXBCXf3uRWPvFhBOq4qYoKsGZ3bzjpsKBqpvxBqriqGfAeD4P3ZJNSmpY
TWA1FwgqNgQw3uR2hk6y2G4on7pRjTX5vxCSWJKr7cKfbKrpaL7chvJs57JswCKt
0oZEFKzqIhrxMCaOl4JYOUJsYdhmiW5VE3wLk9kpmFcCe7L/2dYFAoh7p/FsO8Qd
yIIwzJ/52S4p4r/n9CKkFlUI5nOvFcz11+1PW8sSsElkT1xvcNr2gOOOGT/xvyyQ
v2FnyZjcX8oXsNzW/k/8a385ByRVzEjRt5gG55FwnYejUsHVJwHPV4EO2QcqbODK
NeYiD9dYIkEpyPU/1UvLrswzcl+k/U+wxryN7+Ttk4f8nKCtLHxDT0vivOfSRUxs
9q9NSKAMTGGJiEiymmqC6eYflVsOGSQHU3Jaav17tUJrK0LQ/RasLQQqCqrk7HkM
gyvgpFGWrxEXMMlpqF8inhplKo3HX+M7zBOWSZZBEnRg1yuC6Gp3Cn1X5i2qAjeL
8CQqWaVfp4cm9rfjUKu5U/UUWQAUXVr8joJ71XabKFUl945FEBk7iYOKdYZAIY6i
gjV988Tit8t1z1gcszAZFA/0SP7jv4Os/bJDCcng8PUWm88EuJrtPDeDG4bIlQx/
1etegvIKeHKdPpzLkmvR1dDge3QEk4Kj6CN7KyrG478cFY6ggOyJaLj+GO8qyj7l
5zTVI0qegx0AJKzr4Ho7ggLmKIVzfQHY7f1NyQZpG+8JVp9uiwA1p9Yk6ejazBgc
y/J+r5HJHzJvsR6F6nQFgiVQ4NB1l+5LS/JAKjOKTwTp3oEn4MhRsuG+HDhF20mn
Gu1TKbsZCnPXCwEiOnwc32lfAQOc+Brqy/nOEvimyH/DvfSgPZTb2seXV9mzemJn
ZbMu4t2cdZTEw/FuqCSECB0XkN3S1pyfZDjbk/Ic+ujd2RhSplAg/LaTgo75Ig11
/RhiP4Tv25fk+E3CPKPb3NOro9OcWKbKgh6/eu+0HE5QtZSr6YW8MdMVtT+M9ziD
kBOvBlQLHmiw1Z85ks+XKOps+/abcTtelli36HKR+VvPXhdxHVgwygNu/jHhylMO
Oblj0FSY+Ph1A45QrLIr6iP8AHUiNg+cZF/Y6CbOM161Fv88O3bmrR05STemUsKV
seqwJAnVzkFHn0lUJv7sIg4pCts+Tfls4Xzk3oja6RuGR3ShT6Ldq0vw6wYFNkRT
WwY9Gn+lyrfsXE0gOB2WbFs0EzW/Z8NHdf2INDAniANbLCEhFRc4PT/5KImzBBka
m1SshyzSfiFK6unn2shXnbZYFRzzhiaaHeD7rzyeAliTZjTKe+NDNcEuEDv89Yci
w6FpNLUM5kvxqN+fZ4y/eI+4UMo/TgErgvzHFNni+vpd2mDh1IhMqD/mX9i39Kkx
3zyv1aj/E0oLuvKYACPxJ/hz7Qd1rOtCja1hFWFLFe2aK9fUWzroGhEZoK66O3xz
9xDh0XySfrMe/4jFSc5d0Tji3a0gq3/Qz7Ia2Ew1Z+opk8HH6NsKwLRy/21miVWQ
oGFoZ0JsOEWi1qGCwdJ/BN0YkQzDeFcXbpkMc5WNmvjW/Wv9SCQgr4i8s5tcQCWU
U/MkEIP7h/mf6HgffDRtHOhW8wWQCfhDrSwIOkM6yIXutfXUXY18Nby2SVwYE3UX
g+gFKe7DUJ5xx1UKvNYFCng1Wha4o6HnyxtNa1ihGBIXtEwgQJc56fp8gL5zNS20
JzuvgyuK4j+kU2ZbtYMUiu8ee2IKUM04XWgHKxe36GdINdC48ej/gQw6xKkNNVKU
e8aVrJFprSy5ClaZGk9VnNYlSL6JP15KXp84r6pe/5maIsuqai73MbVg/IinJDZw
pjoI4msBVxonazsx/cczCENHJ/DTqIs8FxKZK5UFt+nhr+R1U3XQUw2d9ltk2ADw
Wa4+FKBnZUT8dKmyGnV4wx7N7mVtgQieJw/gPnZf78MqtbpPgBGDojsa214DThqM
gwadWppIqKoyxHEwC1w+GvcKRdLjlVFTJm5pW/UabQykDCPpVaxjfqp5Ev7of72g
BSVMScmILoTsV5UZJ66ebAlZF8r7jbxJ77lN+ZNcKSAzzE1QlJKPkuzguUaBeH8O
W6xP/m7yBDmIrd/p4skRXgq4K36BHsor6qNQJINvlCCA+rOYcSJUkL8A0Tvz0wl3
RvbRWWKq/CSlyPVVUDxZDbUDVsEucQfvzKReaFFmi+NMM85ehcIIyA3hQxEgDzGP
MQjDcVu69251BiGVfHWqYjHYIVn8lNsDOaJ/0Ith1GB7Zk1LVJ8QvwPTSRejeA2e
7BL4q6IMmvXNgBfgpWLgv0VUttJFR2YHB8vMmHcwghGkDGZ7/DHT5MUxROCCri0W
L0XROZjVUmIXfV7/fBcFgHaqrY3d/+onSfaH8lF4u0uAU9jeh2sVsPe2mBLJRCp/
7GRHk5pMqinefjk5QN9M9JqiKZ49w0tbUqXqDzcnI+m9X3tkSQwjwQQo351Ek2Cu
QE09RpYK+HPYsqoFUW659IGijhctV7ATgSzYNacMKUV2A8WWMwX/bHotfD9gdz2t
tnB5wU2MjAfKjKFI9x/o1oJ4QHLGmGbapvx9n6BFkvfFqcNFoVKy2D5w9BIchRAY
lYrRDzs5/An0foo/mvYgwqSuez3SdW8F7Zmaj/mjUwkSnBv8iPC1uCSbmhKjRHyR
g+cSh4VX8gK7DhYTaUE2Eo+mxllu1WWAzzFFTiFnp5WOQdqbWJ5EKeFX3qjrqTel
+jJHBCshIgvpH5jWR7w8Hs2/AR45FP/rpEgak8i5ohtXEfcLWUlV7DL57CQHwtd7
bCc5vJcBtUVF+xL47kYIDWJuELCp4vVkbzzyUa4nYU7QN3C6xtE5aLRe/AICS3cU
bVTDWVKNDJBc0ru4GqlTHQY9kMZGVxMwIKafhkigrABolYtdrog/BCr6HLcBX/ZM
UzckjWN+X7myN3jP1WwlO46U5yMTFkaV+l1B6mVm8YXbU27v+VFwPjl1QFWsptRS
Mrub2VN6sh0ohRFJzkP8gu4qPuUbSvSgy9hUFGBC+Qb/l7M/QM6NuRGw1sCbDzdi
okGHXyuIsP2iSJ/kfNSdk3iloae4guog1Vc1hgccBiCPa9QfqfsXRu2zRmLFIzxl
RqdhXsSDIkmp+C+Bfw+cAFDsfPPxj3DWVhsZdZWyzKrMb0my/hYmOFpLKqVyIblm
1DXJZ/BOLnLaMVX6ltV3jYWsZPndLDaBaIjUZhpDf28LR390ibjxA41lix84fIIW
fb9eHMRNCu4R6JnDddue98L+WDHw6LAC/BwRvobqR4EUW4KTUAevt0kqDhISvLz8
WQnHoPrVEq/6RQjA0THnVT/Um8qFu9RUA8Xs4kDEH6sM6cYcZp+SC/ywINW5dXCW
xFhgISKTTILaWABdiljBdSTHNp+2WNt0u7wUTmrsF28P2w8JxjX2AbZAlP9SPrFI
w2HOpVvN7j6JFzrOQ+l57xyOrSm4r2oE4CRT3v7HhSgrGhcKomYB9YzR5I39ZtSE
phFlfBu6gtG46eVrOesCkvoFf0KL0vPhuYjhTYwQNU7eu60drvXKLlXHdsnRTLMe
EQSmOnFVvV05kvmzwqssjFaSOxqor6Gxy1OMsjQzd+G3EHbihM6usqfyKkC1hm/n
tb8T1zkS4cQ9jWlxZcnWHqBH41e0l14gJ2nGZWd2CmQaLyvaimM3PSE1muQld4xb
uxwe0mFMwtMrQ9iX4N7tS+B6U3AUF+JYeUVUieELEKpu5jzweltDlnJorhMNkiW5
+NJYDx8tLPYzneHUe7b7xF3aw8WnqfuWkZ0TFmONAANB0KcAKJvhR8Ye+2hVPZlh
cl058Q1LpobFaVVZeRpDcAB9Tr1hDmp6wIJ9DOMUJddEWufLVsknxQJx4aOtAW7a
mSDr6Ak8sSAzJO72rwBviTx1oKKGeYMDbHEIBmL0UnCh98rCI8WeMUwcrUfCkPY7
LmydHHYexVstY3aISGGNAxACDZRJCe7G0lapPTI8Bb0WBeagSNreVd2ZZWDTwKMy
MtdgKV1tirA7xshflBRUsD3aLj1LwaKrWL2tuubyIDuebBvKryIXHJ7S4dxUl2gt
i4gArOuO+Uaj1dOxAGt3gPus/KR8f+pfmQSHpkexfDdAGnQh26jhkmtN6ppWnTBH
Im6OHp4U4eSnDRkiC8e87M9o14cDn9HyR0Zg+8xzisa4TL8Ate02sIGmC4lkr8mG
LIjeJ/JL9HWynE7B5QueQahMkuVkjvlIPV+/+VQ30NLLUiOAs8yqsTvnmqc/Q6BK
e3Wrhv4WXXLhgqDAhADNWJ5lEe2nzm8ZoKkmkgunUKVYHS49IIgjmMgsgVbga81G
BJaAUUhSfI0l2iIie50wFxRP86PbPJqy5LnzHFs1B/rgbF5Dn1uNAQmK2ipRrdX7
+5t76DvA2w3775ly8DjbIiZtDUkSqyQ1mBpAHm+4vylyDkFEuq+b4J7xgzx/68Ih
rWSM0ObReOhRU5TUlzF0+6i1SOtlLOsAhEpdTKg4CREruuDNAKgWPVoa7ObtW7wc
7IHwbbFlfg8VVb2ONRe3GD08ASlnozzFcqDjwps4KixZ1EPJRVo5iPF2gMa2wDgA
vjCvn0PteT8I1Ty+2S6FXXpV4QkRa65yyM49Om0yVmgqzlpnhwkDgKkqoCuNF00H
/CN56bn2GM6SJRoeJZDjy80eYsmNnuXt2CujDozWWjXBGHzKzs7/DaHjPEuEWQ3m
UvlxfsPXk4eb0t9or36o8XAoXeD/RmIRqC21liQkI11rFrLOKAX2S0hyfT7vCrYn
vgZizmCydUIPImEbt+2x+41cRn2KloygTZjQvykhOo8b9MUo2GiInKClpr0xMP5Y
8zP70wt97tpTb6GNce0wM1iEhm3Gt/RNiLeNT7dawySAjzJRVigXauvQ8zf+TBfu
WPdlWtcjgrDThnw5hP/h6xFglGgeAD0RNGdDRRXW+GsAZ5dmFasse2kXD70BvC42
VBAYHO1AROcYpTNW5YLcJMPueSL2nZm26hbj5xah9WBNQhF/EzKIcYWp1MIhItUi
fssvBFI2/sVTeTpXlDsEI9y3vA6clLDlIbMUn53KTnn7IsROWaKXdM9okXQ332cC
T7J7YpcfLD3v85Kk1xBe2sVDyUyjt3XzEKqu6isJrKNgRKsYdep3A6fTtd+H4Z3x
0//AXNu+19U2YaqRF5GU8BSknkx5/rddmvZDTV8z+5dC64haBjrrt9Svq2C5tBk5
//s3L69bErGRTjtrfpNdqoslt+gPOMWcVDCZJ9QDFMSM+N2kAXzuvp3efv2BiWmq
l9twzzoJ57ciZPPMt3bXlnOxRvAsPlMIoPYWFtOmKqm0Or2prv50hhFFZVJP8XKf
3kpXBCbcjUsQUZ7U4sRcSn1VyqsigrCubv/QrYjEIumaZYRmwYwD04EiOKkF62b4
zkvfKskA8ucnTpScViwqiBiJhEkzCNKl9orGo1XN9TLQkpgLxLROQ1JByrcZjmVi
9UIQbytV57zuKNgq1nnd9QXjqDO4FMr64T/fykfrwBY/k+JGRCqCdGruMhWgyL8G
ToLp84aG1AD+MwSHlbiGnIn3x7G3AqEc6USGkfjmh9MVIUDVLstBt/khOXxfWg7g
Z0FCGZTT0Q0RvqO1TIA0XmfsjNvyZtnS3dxCI86nhdaqpDZhJFf+CtY8HysXhbdv
EuClvVaK/F0I9ot09GYqyzEadwIjend4gy90QCU2KLKmE8r/4HFdfeGFOOidibeZ
Yzf+ZCLomDSwxh7P5+KHLzw3beKq4A0Gg9kc0ZSg/fKFaH0TF7HzdvOaoO7+fhwW
ETU/bIGOVucUN6GVmb39XfB1UGBY8CJCCTUA8n5ChOWkCnpIJ7MmThgR2O66hNZz
qfr2HmP9RfV18F4gr0s/Mh+CECw6FGiRLhQJ+BPeJP9jazfnjLDn0GXXfXRTysAh
uPPTj7EHVSHz7JpUsdpQo7clo+J8N5zS2LwNJO9TNrSesMsQmT36CyBQE/YgCZKn
HMNxj3yyu18xB/2x8/ekfn7MzSpaEXNP7zao3Nb5/PT5ua8BgSU4KFfnE64qFS1c
/jYnJjDPwxOEvXMChULJify872TcWpQqWL+JiPZfPJ3aPpr3eq43Thsh++qPvXVi
IofdAuoIOMtRAQpIpavRiAqDfQveI3VyV3DzYRkOCl8HS3WlHOyxwNV3c5OUGCGz
emIJxLZ+B1tQ+MfXPR5+p/C8PphQZX9LNQcZTFBZ/u3i4BKnze+nzAHnFQDqi8hq
MrdxUm7p/2xk2lRVkOIQda/3lIRwKA0hbDbqUdPtWGxdgzEWdk6Bx0Vhc618bBQt
WhHBUBrK/GamZaKLqSQOWLCuG9UXuS0J58JrkHfoEoMm/85QZizp+WsF0NylJ7D5
KHJjv7Mi/Q7veJjO9zJrymmdFfcazFjMODSMc2h0sDjVtMDJiNRysOoeGuYX5Umy
TE3n92u6Wc4M8PYvFiqZC1foHu6b3Yy9HUpV+MlbyET+wahMjbYA03Q10MwWgDPs
O1ii89ceeBJIlJXQ3muZ48XDK/1Fue0XN0cgow3Vi8oXFOr9/heAUqGuwEnxW2nq
bKFW7DApIUCMlpWWG9ySlQg2YJdJRgLvuzijOivWNS5qFahWnJenFOlp4aVLQ8CU
AoVcU4DnwJsmp+zXvGTG+G82crCGMimodvQ3NQWMxsdh3hyGuESToupYkwi0JS48
nYG6R8D3IJvpWeXbV7BhJ73Cfa3a8kOq/kcthHQxjIe2r7DJB93rOOb60aK99tWR
Dxdty06FWABU/EvKqenxhkvrF6Q/bNyWPcr0yGa/mi8qvmTGgqSEtdS5cn2Qsp1z
/y1GG9tulF04d3glmCd9ZhfrStXJWm/FMLCtzzX/ux8Wmf0XWSfFumsZ7rP627u8
/rUmkq3q2AEBC6hNCVzcA8qpmN9yirMVgILe8AmtL+lC0BVQBfjBCQ1zarylb6zK
TjyEAK4VJ+ekaa07y4HihaRh3ioDwwDcqS7gHzIjj1KXopI9NKYB40k0Fhktkhr1
5uX1BDQ2m4Jcwj2BVn2iZkOq5d+c0Ed4x0sxwOy5Km/POVUthT3Xb+Fb9Kqgpsuw
tudQOk7F+csQImLuN4t/yL/98Q4JIUVyTOpI/qSKaAKp5h5NiM/TxfxVNajKMDjU
3SjLg/7MEP7PU0s6951+SB9qprHI5HoOv37Ksk9NORHoDpuos2MHc0VmintXA8l+
S++ne2K12GdLWZm898OHFqBh/39o7zm+ce6L5akgVsfNQqAyQgyolvC3UVh8XT31
SIxPAqLEPjkFkOaxf9POPLIEcCy8vOe2tV3z6oHGgqzf9+b1NjSlbZN2RCP1lNMV
obnmbrqiF9MMAuSEFOGQ89vPJgm2qvN0DuHwK80dVFHRlhdJBeq7xBW0ag3hesCI
hrNEsoz8Q9vBPS2NxytghgfKGX+StYvIDrNgozSjP5UKMMfLvC9Urecv/vNH25Tl
8HX1q2UNzK2yZDKJXNhkhA1NPBWUltT90Vu2QY66WKaVazIdEO46gkk4XV6y5+qO
+8vuiHp0xKnktZnN7Ut3Ft+Qyi+sib4TxbKFEJUq4B5yiXvA683v5p2WjEkmdrsZ
yqN1SgOR2qTkWxf4rc347cYPMpJkrP3EhCFMKF7cFAuhyuyUwX7fOC+Tdj/4mnHK
I7AbaXWxTprmQJ5yjOFifcePHJKmZaMnETCXksecYHbI3+Yjjc319DtO4DHwPZwE
4oEPYiz1efOvyoAmMyOOkGB5WRyB+KZiPzegwVTFc/eDjLJNQymImIpbf8qUNQ7g
gh6sITQEuVrp3XPEGVE1kL0sUH0/J6tDjQrszETr9VOhaGgYi4SaNPZ7gMXO6QZI
zLy9NoABk63hBZnqMQUG3O4/7nltsSv1PYQVZFIDe+cR4pEz7elSfiDL/iuv7gZB
2dn7fkJtMjfjJhOnVY+qisZ9F1wfURKcScHH5wCGyEPbTxivErb+dkqpKM3o7JDX
PUmR3O+1KNDf9a8QqYcohpMV/jUMteuM7UE50t6XZDN3f8iQ4hyPTaZCEPMdAdSp
FjjNLZVj9OS05uiJLcDcALLhxoroFuvctqdFNj6tdyeOr1aiMqKSeMgT6HuJVktj
wtb27LIIu6/ziB2P4euP0eurYK7PfAUTwyfuqFghLWEbu3udQzxZxR2kB2ZXAg1E
VcB/z2kyr/Hzk7wnv9t2A8vJ4gaTkLUSUa/PXfsyfmfGVsa4D/LOtiZ92i9Yll8U
T4hj3LiNyzDzmsGCmzlybMpPD0ayKRh/tJW/64RjtrrN+g3bjHLF0D1uznTnBsNX
mthYrR4lnN24JaytKGWvr9Fiumrsj2S7Qj725xvcffjS07sePMNA8Jb+BIt8Louy
viHogSIN9eay75F0BIem8h73rQM/fgWzp2tt0BCPZO1PXdyQpy1dxi5IMcy+0Uik
jMjcUE0TQUbJKet7ghLsGy8lTzYXeEx0vwmVfDhIZvMXZKfQxj5JUFucOwjyi7QC
Onw+4GAgoKPaodLZHoNYkW2mDlI2kGGafNnpEG+ALlIsY9kzZXofxtaLTyvOrKaJ
NBHARN4KQuQYLN0SQfSZe6QPmtsCsKyuIJPuWJx/ptyZCwj1i6pgkZNEb3NZH1K6
FA+UopdBRnRgHJ9L1RhOHEb/tHEZtrBOKDW6nk2BN6zbcR/TDmBTK95qEsWzZOdm
BtdkD/pYN5ZhtJOwCGbmrzBWiqfjwv21HD5nnj8x2OK8nGJzEoPPemb0DMwt0l3w
SUt/NBu8ooNf/GlljbmyU6avdAUApSrvuNSzyYllq6beqRFd65I82xrBECMHXLGX
LF6XYV+4DTqDGrAKK7bE6OoaCfg4Oqkf6mnQpamNyk54LOSw/xvrWXrrdMgOvMKV
ssJymZlxqyrAbmJF15rhJ1mz5HQFMWZ81FcjoCfY9B/2181Lh0vWWTU6Yi8OkZ+d
ln9JD9ubeYChim39k/x8ksqZ/b/4JRXokw8cjgB9F2m+75RVTHUFC0zVf2nz9qJf
9Z4qG5wn/H76MnjQmb829xg40sUnwKyzjmOIeiBvolwmPafoeKJuifJwY9lPTaRl
3j77DbJJ93kBAV+2C62tJRqt/ERzgto6SA/kagGgBryAjFsxDx9bBLGmw7oTUFZp
tX3uZw6K3fpzm3ZqYuhVS07YXXJB2Exdkr2LObjfmpcnu4ul+epID9TRwZNFSe7U
XIugFMJzOyKYD0qVeJHFYi4vetTbfIvNjlXnM+EMhQpNSd3XeYwLP9CJA59+MNU/
KAbNt2VL90Rv25q0E/ZjnpEWOfTrdZWulf0XUXxNGtZRH1JRHgSR3OGRcDFo+ghf
uxAcVsypu7TUZO3SRUDpDajT+UiLDOED+VREYTBXZN7yrCGWxQx61LEG7SmBM2Mu
jqDMLIJslKbvKOkR9fNSKVUI3ihfGc2Hz+m75b7QqhDQ6GeQA/XUvzY2gkquSxre
frlpv4IVTTp9YTWAzw7+S/5NxHqRlACB4NMmbwfN2qRI5DBlFUjk9s987nPh5uFr
ZnyHK8mjds8ytH1uFmME20SNziGimxWiRIc6s+5Y+9aVxEeQVj/WDMIcMFwIv2NZ
T9Ra9fo3K+H5Hcubm9/0XEGAAn87b+ulfmB2nmQQtYNrfqzfVlbFPh6MOOOnCbW/
bMAOjaR5x6od9LpdzbHs/X6PBthEqnhWJg3eVvliJ4wgrpNj/xIL+G4uFI/dEd9m
Bx+BW3McMZmiwUcCc2feQnaAwi9I5eKUKivYoXGvnA+AmCQ+zgPZ43H4Q5kXAFO+
QJ9oXAO63HV9rLJb1gvOBX4upDfk+gCjIa6R+/DLltyLyE3RfvJd2pE94Fk6LhlA
AzXEaV94/Jw5bi+xJIZmR7vYr7JPgV/cZiykYSGJcUjalES7zM+AOC1JRUangeFT
ZWHZm38Wi2Pt+Pb6loLAd6pXsiYkAtyutkO9D0xpYvgWs6dBMBEULuYDYhfRBu6s
wH+zNlgSYcLUfM8yc3Tl6yBQlHlq6AimwaXgyWPXyKwRgEExuwNuMGaPivROH5kK
fpecH/9nwyoichL+xhwxmoIqGo8KhCPPYra+eruMrwkyZvTpEM+J+sNW2yITB8XP
IzDqPcEyXRT3NW+HzCVWUG/8xAJm6awW8q2RMZ56lA8tfPVWN+sgLF+Xcc+U7WGe
IkOQMf4LrexNtDT63N9lMHFAKfU+shTsctvKy/NfTw+qHVQlBXcMrrtWA09vVHoi
x3xMNFn5PgnCYcBjeX6bFNwUUluZvB6q9DrT6Doqz2MZ2Oa4/iyZ6mQGgdBzNvu0
QDs2QT9mg/q/HPPAz4KXItWlJrOlScD5B4oEUu6DA3Uwg5JJyKdu26aK1VWFqqVp
svv9TyEzq2zKJQVzM8xh3NHmpSugAAfJ0OOb4H4CxnMAaUSIx6aoCurM76+JPHwN
OL1F8I92FFvIAOwVZVpWa24LROZiy9JxfAU3actTpYJq0m6CCQX3HeVOROgOzYBm
0pNu6Tnv9zEI01/V6f7F4DI4Er2jFf8DszULJCu+xnAzAMKnskFlMnfhrFSQhXnk
CG1AxQSpHf7VPubfdQ5tx21SES1tP8FKthFSNBYJzHHENwc3kIri1z5Syi2mqdmJ
2j5xmIkOg7KiAtvdYVMaZf/sCW3/Hgw39vuwmnJ/OR1VbtpOJhGxaZT8xN6QQq+d
Y6IMVT1wAgWuGBUZ9a5EiEN+ntgEe9bux1RPEzLNoejOw1ZajLVN9/52akbrk5oT
4nZpompfzuIinKHFO0Rlx8v7YHyIqB0p97todDK6mT6KKhGcLuqrjpZL1Ikg1qiI
2BTBlYmeiFrr+BfTLfsjazqBL/2dsCumdenBZ8ED/Ypr72VK+diA6ZvowwNgPn/4
bQpyDtC4xKnvDD9wwqJrid5RF46DKTwvWekyMfW95Lf72EFGYXAqihZyKK6hwebc
FOs3tcuR2MX8Zd187ya++UsGIiAyu9LW9UiGVpSzRA1NFUpAQNAE5ZxdW0rZBupO
OzrpmsrgW/zHF5g3x/ajtXTkwVc1Q/nqxyPuyK6dnnbHebnHHmhcp534XMTWg90M
fZ79/N3aZibjNizL6QfJF1JipzUDyLgaZAKb7gNsXaz9E2UJSH5WdaToE8wsyxfg
ngtriroN9LAOlqsU4oVldFT/zGh4SVwxUf56u+TDjv5POXw3NcsIv8S0SV8wG8kz
OEjsSkvhWCQ2/31BwVChkrxTV5gDr+XCUieUoj2ItdqmJ0j2GlLso9NnadSEjkuY
B4zvrI+9BHKeeJ3w+kAsP0fyI+qMNCJeJes7OO8YzImdjClzFvk9XqasJvCnqTuW
n86jxYYnWpYdFDOZ804Tc2aJZdqgV9UIKrgfaYY9nbtUkVmqbKF5rYJ58ZIe216U
IVT/LkBMdiHqcbKLGET10bgibQ1L7IlNwcDoj7RmGkGOONw+j6BItxHKW/HvmTyM
qO3kKbvwB8zmwntxqYt96ew+HZRTcWD2bgOK74kIs+FzBzBXvJGjPwVTLM/PrxJZ
r0SR56Pzx4tnSH3UhUOfSA2V0F3PtsR2lzwQ59C94tnpcL/804dQySs3HwiG7iil
6fHYG+OQ9hR048tQ6rpE4WqfyZAIlHBvmupJiJ0a0PPYKtME7xAygqFqXw6SDzL1
pbnpxoyrpeLnklxiRFstsK0QjgXAu9oQDwV1Ff2mWOLi5fWUS1Rw959QkXy5c2G8
rE24n3fpgHDbmRb3OjpC5MInj196n3yqoq5rqD5c7UxzMFywrpcIqnEb5EQqUmWq
LiWOaWqVMN18la7nw139o9jP53ljzIhQF7Fm9/zRJzmu8BxkmidBbrgoZ9E46oa9
A+K14oG7fl/OgxQD+CqizAWMJK1TWH9xcEdkLCeEYb26d5Y3KkCs6074+NNLstcm
WIqJJPNvKfsFP6OHg282rYJVfw3+e/8NZPfjCG8wCAEj/jJYZFLilD9VZQPEoX8a
2jIf0mEyhsuwXwKlV6NH+mxG5CAhqCSAfctacUB59abVL2vebp+Vbn0y4vNxl1he
99it4Lam3aTCRl//kFVrckZwr3O/uXWptv3W3VUeljn0QXBWnqqyiHO5vEDN16V9
sUVD1fQA42wZrZItWaRlq76qaMt72ejTyggqI1TXoaUKzO7QUUPJ5eR2WaVnUgDo
dsnzojUD8mOk1aqouOE/6dUuNip+jA4IKW+HVN9pn/IbVKD5laAXou/LBxdZh+c5
IibOneCI+yzJ5sP+gBGmEN4DJa6hEg6S1zYaBR262NToHBoFc48q7cAeB2a7/bKV
OHv0Q+w3ewvKxqa6BUD59kl9cBBZhAz1YNaIUOOgnACyii7/NPQ1xxh6D0wk5Zn8
WDeLEB+MXpwwriZwJkeoEmJ6sNPQjrs980FAfXBWktVJJ/YdALJpVfNMZ6836tX7
qrR2Z4jjelUQnHS1/x9cEtxmQSyjQBZG65Nk1QKCMxDnUcHV51F2p0WNkbfsn8cP
ExFYpP1M4RJ3VvJABLifszREpZHMv83879ihW/LQxOejD7pJ03BO6VMpyxrSPk9s
23hFFSk2AxpGpeRRbRBZZ1FddV/KMbG6s/Hc81DQ3JDpB6EUWsoR0NwAg9i/A4DA
i3QQRPScG+IHDySh5XoQxKbDFGIcR8rv6ImS3YNV2yyYXh4EWF1qV/xxMcyOZuCX
6Uh6uPBgGkxhSuRickTKYoAhKlSWk9KWBhou1Wu0J7I/+MqY7zyOZMHycIoKc+5V
R4iQdQSetPH3zrCzDmRgNx/+qsuyZEskX96jianUnXfnipRDdam/xsVqf9G1Y3oL
NEPoxqZeY4tUv8J4pVMYo3JMrvKARGSLmyLKYnW3ybQcx1z25WIPHrOGl0PYa3VQ
tCRhxkeo5RLgmnQGT+YbJ79J21QIxlTzi5BrqTgaQ9wk5IigsfmcuFCN+abzd8g/
g3XgYNWDgq7DxpGzfHl8zkCXbWGGNxaBJnqz9E5gj1xZshARoVlcRV6fhj0h2W8Y
Z1rBPCtcD2OXgn4XeVYosOmklGYdHbXPZVxhCy0mxX6oseH/9pvSGsGVGt+MYI3Y
yQTk1K1T9E1rfFFqfgu8QkcV9Gk6ig/WPLYKdLNVt+paf4n9AAcQpsp/JqG/Rnri
lnGVlj+vvd7EvCQypNnku5pltDddQE8TjaSztl0uTh1m1ug17YKnz1CEkXf+iSc6
BZa4zIFnigQhAciqT6raPQEusng1YsoTr/HQG6F1+hOqk2dJoybjQ8t+c1btaN/4
ILEzui9aWhYrFRPUvlNrDyeP/cCyuAdQ3peMkXM8c4IgifZEzBqA1RwYs+pQKG+I
D8FC8PlHGSypHzT5qgKw0w4Z1iLLHhdG1oQ2NTpHg/zPF3jJhwcZRkgP3PlkFWCp
E/GGOo4u9ruQk7U+YtW37QwqTi8NO3vnEdN/RRG1bmDywb38mWVATaXPRNtFjVGm
iu1d9rimlkg+/Y41LfT8HQoS5lvBaXZfwyvqmZCj2OIFrz70Gr7n7+7RTCbgwFUI
M5Qm2pUmZiC11m6AEsEs6sxGlStCMG9o4qKZaZ2dfxa1arNI+VOyZr0SG32Y1CFY
QMRF1hBNKcOnYI2ALLLCEwOPmi7O5G5csECZmQ/EtMz9l4d8b0yY3VzmiLO1R7ZX
OENswZA7E+LgWlGwLSQXKuINV/aowptvLr45e8FbbU6CfSLHgqfNUpkUcObF/QuI
uWfrpMciR1Zjr8P+eqMRqpDQSStvatbMZsKcZjIFBtjrQBQqaayjjTuoFH77NkD8
1EkRKcENZIQ7ej435HBDw4MF3lup2qfgMMazNbo46HqlOkLxAgqMP+L/mfJKR2jG
XZuTPVBC0FEM3gLy9isXg1nTZT5fngmQuYy1/132t0JdzAMT4EqMW5q3i+ejqsGC
oA86Fq8YhHc0Ht8glZNznzBIQgC+I36CT1jsbNOqFfI5RM0xaPdCwMdWkRJUsWA0
uzMrUl6Kn+l45fOnrp37F0VDw1TQeUEXNl9InScvsW7uEZLxhT0MYf/cMFzCjW8R
Naj0xh9YUJyQWkdGt8mR9elu6LF0NJWQwGbDW4DiBmFAKMBTrAVzs+5cJnWq11vK
mEYe3qs0SEf1kJ+UWHOO51ZlUVYCRyul02ZwagagWkz+7WChPJgvADcswPmjap5p
qsjWGH5rU9s5NQGzmeobOeXITFUoYiXAZz1/RqoZNER1189wMMtlKhhilBucFsPS
+5oxkj/rqQawZ8YfzGCQjp+ogT6cEbZk6wZRCvVxnYA4w7Bix9Y87c70TBrzr+ai
os1qvPaY6/qX72fFYZGtSKhAYIMRIx1XyDApoC9wyqDtU+9nVwdKbuLJs7i/OKkT
xKFXMkQTZ1Redg1IcQqhaXiY4StphspJKV6tgyNX8uaEUaKtH1s/HctfRgXeHlIK
pfrOWHwF2A59yX7MtdJ9GkHee0itxgVnbs+qAT5ME0gW5r1J9MWJnfZprbZnWBX1
qFJBOBrzKoiWIQ1cJGpjTSbHGHoGqT4OyIRkebWp//Ok9PFJ6/6RoexqpZVHEHU8
SBJdGA9lruKBQrNfjsRR0lcYmI5mLthRX2ePq7v++pWIdtT8Nb3eueCh0L4015xS
oNfoqCATTqX4uME+e141CqPuzhxZllbTMezNqgbiWPXr6p1Bv1CvTgrm0nIXXUVW
9+BPSKt5mcUjhC1FGHMfi5V07vUZ2CzIz0IG4LB4qNajS8o6iqB+uOC2+UwSLQtr
2sX7/OlvJ4wbipTIZN8EYAbX5L373Hg5Fr4RQ9Xsn+EQym7v3JbATv3X6q4jPbJX
q1KS+48Z7ucsT2ozr5XSWPvPMjS4Sn9Ky3iD/pXPfCRCKr6E7tcdvXwjK9d+j+mx
5h0Q8U+u3vOvceJWkl6UwUHfbVedQ2i2kSdTgRLEVh8ZrKz4vBsaK+amInwr02W8
ST7PQQB75VSVsPJ+LYSrXOPS8XaREfcAcalPB70huc8I21GPCtuJSqCnLAJpoHvg
DYW0FMFemGhr+lexELw9JTJTCFvn4yb0R6JqZYp6WuUc42T4IzwROy8kU079glUz
lxyN892pwlPs2LUtYhhx2y/QahbaBp8tgvb1/29nqh6VDEj5GqTqWxkLSmnBpRTv
XnVIVexsXBH2aBZ1u+1LNwsdiHILjrM+1iDJ+LFsj/mFcQjHwkeMzb+PJ+16dRFn
jzqsD0GvgYiVbfv4Inil7X2rUNXWeqbLzMMaLMAEO//WDR3lBaUhJNnY3VJnY4Pf
Xz/2/bmUid/KKN8oOG9/kuj+/XV47WrWe+WywZs9WeIaLALB152hJBkqY7i+DFz8
QRbSqcKNlhH71MDddF0QyMNi9bHz0eM1f416EMFKL0Yr2VrrfXMA/hkAFCzPatoB
1OWUPPyrxpBM84yev2GmrA/ynZTbkuATEOe3z/FA8xpam9XHwegD7Swga1qh8GHr
DbRaHdkK25vUU/A6AB80Oc1wnCRUbg4wiG9VpOptkfck4eAFR/K8wviumjse0fEV
D/HQifeP188qYUmGQnKKLy92DTMjbPfyBUynvpEzQkHlhlkIA4MJjXnnZGq7kers
eMvNAR3gassBCFAiMXTDH9va1+eCAT01CaKIaU1cujJ7AA2TpzMDsuOcIBzp9Lah
JjXJJj31Zc3+MHzjC9uuclIBA6bpD2eh62LaZDKEYSCTJRKeskJfKev8jd+iqz6o
ocPA2BcfK4+zOC1PvWvcGzEhx9Gc9zjKomeI31UB6F1E6e0ghkGFPQLiBlNs2LJ+
aKuIj39DtOn6SbHDBbGn5c1y3K9aHH6mCxBbn6CkyfRs/UB9LwwQ62mivaE+cye3
ct5zKQroLeDey62b155wnMAwKdxC7KdHaq7xV8PoH4LLvTYkPMfmpB4RkpPQ47+z
RvTRV6FA2xtsIRz0cJ9oHe+1mPqwC7RkXZWa0RTn9oHxmDPTTgWGRLbj0jmRXPiz
hpb+gPiSfaH/wysQWGM79DEGNmgCNdo8YeRon0K7/21kjlsJnHruoqNukLMbTReL
jB1edNM7qV14aaSN1xHiGQMYehY43PkKP+kaAMXMNVVdKro1txxT5s1D+OjQuEec
b2W4GPJvmYks1Urxtzq3HDqmyFJKv/uGZDcMHlx+8GJj2IXhzVxbjw4jZQVNwUzm
h+jLch3vs5WXSEK1vT3InFoiB2ARMm5hhphXpNoUrGRgXhl3yOQoz8X424GkNELv
g1UOjRR2WfZg0ZQrNVwNsuJKuGrf7mNiAXwalsVJiM4Rcaj9G9oN+gUbBOiO/13/
JWlJJiRoYVphgaKJBKuq7UprhM9RjcD4g9vXAWFLJn80ITK1vtlrQzO1KfR/8t0l
rDI4Qu9eR6YdkF52zcIhHNDEBjiWWIgjbS6wBxG8OXvn8EC5iSiEfLN/tjcQIkD3
YBSdip9d7PXeCzoyr4rzegLq99BOQd/rSd8pCX26b8T7I3AO2RaaaMYKI/ZHffin
XhHUpqAI3jrDhGmZjtaBbIeA5uy0yvknb9v+jR0NseBbAEh9C/jmhsJjQ5nimJS3
KBgRWzR44iFAU7MaU5micaocdYHdVD/nWhZfcCiaUF+GZ6YeD05pA8DkGl3xhBAD
+6wX3IONr8kKDjyZ3t7yCWmGvSa8E6vjcvouofzRdIe4wLG/4ERwirpdzXyO3/Cx
T5p6s2ugE0q841LKixuRf2NNhvN1+wYCuQmCOKpXaWnzOYxV+h4OPT8RB2I9dBe8
2PIU/B4VqoyGw6ePOrJsZ57GSHVAchwAGbo9GW1swpqZqNZV341tp6O0D6iMP1P0
NB/bzSoFpHPDPzXUGTQS9HtcthCisYk5sG7XqwNRfZxFzgHIbnHFT4m2V3OKX9Be
H8jGw1i6EodBuLpsvdyZ7i9ZMYWjZXcELVtFiBoR+ZBFUBugRx2cfC2AiJaI4ncb
CX2CO3lDwMXYIGUjYaZI5nOhTrtGHq7Gx7euKrDaaX3e/Ch7sWC6L8jl/9nPv1xJ
le1rXAi9AdPA/9Vc+wk9fgMX+oqV8rT8/pgh9M7tttUdLppaSJOOoUDcC7nJS3l0
x/GQyYnJfysxjiT/UMYXCxgiKy/KSzagaklcfIWD9KHz6Ky565Oi+midn/n1yOVv
KPWn9zFeRqbviIhoK4+0+o+YsUnF49OO94U2KqbS206I6hgwPt6EKU6ecSzscTLk
/54XUUVJQYKU8Z7wZWRzr9ZkNLpzqeSOfnKewuRTRuqH7CymZhuwCv/uvVI4orbp
4o1zJE5nRoN+VAvCKQ5WlQr/9F+FbyXxPYr2ef1moCCTVl0tAt3IqQamWXyBkl8b
boDchOZOpeicvx3AJs1Rf/F6xy7IpYs1UdyVjnNbkbUa/A3rasqV+YFhz9dyxGtp
OLbcNXSF5zd7AV13H6heokcxxMd959L6oRhHdjFSVywsxEjOU9lccZLUwmr5yGZ3
iSIbeOsxBnoKWXAAZ5UQ4IzKQDMbijMl0ey/RrYQ/AIyKiPcwlyDAyzpHHZJfGq5
HjKhzUGnoz2sUnC6Y9OnBPReOvhieSXTv/qFid8U8F0quYrgUxWwIetYYjsllkOP
zEFL800BKB3pNLhtiCtQwXmhhHHLkm3bA0Si9nYeuqQsn7WiH8fn6xFkyOrgk4Hu
AJcFrHzrqUxiXD2XBnCKDHRmcaIhQ7TMkFbkKjYeth4ak3CmrxQ5FLEnbfbQ5rTV
yiPISVHbm+9NCRTqNzX97ejzPCubc60iwFfzeK0r9WzXU9eJxqVUu3G0qOVBvb7b
aUIt77mg5VjNhSBjjHdrHurCB6wVtfg1Hv5FwvXNfFqkuoW7CkZF3E/oo8fMMjr+
SAGdTQ2hvnr4S3bXEy2UOm+B08z1mYE2ccyRS8FgU5IsZ8ODPbXHAWkEwAVV18eJ
m0j+EIG9RwFUWYXEh7HWe2YtTQv0c+3LVRccumY9XOnCUgjJ2UUqri2r9K27WMZG
wozGSNIAV3o0geCooA9y+58+BLJ8goFPiDzhGl0At4veFBo+WVIf/YCS2y6lcPGR
CFpsrYE88CNamQgndEqqzPr2wqaRgcLF7/5TXWp2Az66lk3zIKJins837ahUqtKT
oBQMN9q1/l1cK/RAGkrP5VsWBN+nWj359CDsOoZm2ZRdQc/mbKiOspZOfLg2aP+i
ctc6GNkXIp4xeMUylyo18qEv3TMYo4xjhkikOOoGlhbmWshSjn2M3GRHaAZBV89c
r1rxLYeRIZmvpfk30OFFI8BRXPjEqqmBQZ0381nCd+/SLnRkFlpLOA2sSwj4Ez5a
V9YvXOsTD8VPGpueIY/b0MTJqhIMAPvjCx+BaQj5fOaM1bx5+oyIH4jrLEHFK2lt
wl68Kgym0FFgRRJbwPXtQjUVLcc2r6j6w53WmKIGkOgWgmqryew/3sffYvS+uZ3c
25G/Qg/U9hJOKA6SzEclNYDEhoD2ZKItGGEC9pGYOUGbMomIqQ1tqTME8oh2X7xN
ThDv6pb5Lb68Jn6Wp9d7uSZD7vHyH0Bw4wknrRacYAdqf8jcGqLvmFdLTnoMj0Zt
FlIA4oHivgucSq1rpgcQwMFArNOMD2IaIOj/zo7yXtUZZSf25yGZPGek13Dfvro3
aFXKT2RfcudYECMxECyRTWEyDlc5eutaKAvd/aA8px2fUt0odlbOcHw2diD2HkwK
9UcNkrw9wYarCiedQWd/GGoHyC+nNyvdSaR59XS4mFdKItYOWWCvQfqt/ywubJ6w
VqwrGT+WC1JUEMTWrUz4c8kMceGJqWCdmuPbIRgRyARUMdnGNyYVszN4+RuKYkJC
GZszrQEt3w/3MxKgWYHaL+FkQ2ShKAs5x5WcUuzsVLkzhv4jkj/4WpuJxJ/MhHda
kDhy3eOKvycl3Wve8xcl1vvlYXBUuI/tMrij8CuwL0g860GQcMo9HfSzuSHlk3PV
rupclAIKc+/tsTCwVQvpIXrdMqOHP7g6fLpjX51iGRAGEF2kcCQIYe6ktVUic+u6
Ph0qkmWRe/GMan9jXsf571UKVWzhaN7l1lN8TygKVfMa/vLg/RM33QqmnuHcYFna
qRtFc4p450rlG6c6FsUeuw4aLhplQTq+8OqpPa2eu2SnAsCHw0nsPzb3VSMTQghs
VTK2NVvRMbk86hFF62AzZGjhJO8OJ254bJx7K41d1CnwvntR3lx9rvbKs5IXWyVz
4aAEpWnZFzzejjewctab8lWdlCh3vsgPczXgxVqTNYshWYjz2bX0z3wnTtPAuyt9
XhLbGKz0MV0Zuv5WlfQ3YEJwjJRX1pk+l0x7HKTjPmDlZZbQFUVTtae+L9SHpUiR
ZOuwKikKMclG0G3TeO1qpL+oPQg856wnAtniWCNRSmpM+jnMLltCZiCb4jlp+Ybk
L711ZITbDytBqcxVf6kT39CovZ0tPGvuR6Am6zhndZBQIYAqvG+UDVby2Tuqw5F1
ANwBuh8H2emM8yYvhP6xq98iGHfoDmXpOxotmmcojE2YXQ1zfep640uCVfR47YGj
9r+oT9vdYHqtw6aPf9mng+J0nQzjpSb7iTAVfcp9haanKNJU72u/vzT7PZUmGhoY
tCBHD1mKANVQNYgoBfbFjKnIt1AcgYBlQUo+TZ+P9qbh1Y0Yiq2oEJC3GmTwT1Hb
9wTKK2/Osk98SwRgGAmLQPkSHt5a4zYXOSJtfgq77/aZ4LMZ1rv+BadJEkJArHjs
NCA6OtoInJPlm9fcsh7fJt/JwVIygxbKoTJxY5L66D0435W3S92ilY4In5qMV6wW
rpMjhZU8qPVIVJFXfEaWTJm/9FBBQ0WRMJ6vXP7jHbJ0TBvycR87oEtc/Wi27ksC
s1NIWPUiFI7uamZR1SiceMA7CfIri1uPr8YSQT8NQvBZrgXAYQ1M+zamaOyUt+La
ozYTXluaANv+qS/yMUGBhiI5sZpoNb6HoG2+etBgLyPuiYvvwWaiPbOSH8uuJLDL
r9uNBgarSgE2sfPFfBVmdCGxE5rnUUPH8p5q50gdkn0ssXiwxa2T3J6G8ykY4dX0
DdgSlwFxQaYjugmDMOYA+IlkywQY1GUsMaIsNzHeHWQjArOq91Kv1fRiBSY+FboZ
vTTyIUWLiBzeIzIVZ4kSw9Jxy3Yt6SfEmS7L/XGkYhg2vl3NphurJKjBSzmdGGRv
yG0EPJF5dM9w0C3k+e62reuq9U7N20eFgUSswzgAlf05Nx/GGesmJRaQmooYMNNb
ge0W9L220W+ZY1Qi/7O/kk+GzxQy6H1iOMsljOZ+Ao5iPLgB3JuouQMpLCGqkp1l
X0vXi1CX5UUFiQvek4j5hIU4k4M3w7Ei25quFDQEl6GQbGGWJ1tcXJYmp4BXqDho
DCHsYw55KyWp8FBRzMpsl0woR3yphyn19eyjaR+ejMcIR9azauXfNus3O5MUFpQr
Kv2Diwef9QI/aziMLvem0BrFkGrYZ2Lxyew3DSqPO7YHbILqd9s9+pizpAmfI+1m
WyfnPPjTsStmhQrS4TC2X7UWPOxgSJZQVFm+DbyS7oDSrTBT4Ggf19sJLFz4eSsf
lIlAW7bAR7T3T8JasnT2nJmlUGiV/HdUsEgMRGEFmFNw0H3Mp616OYsEdyT2WOwh
h6IjqhzMIAOj4jlN5YNyGFvQ8yBHo9LDsaHi7gnvr0SjD6LHgK76WHl4CXQ5cnAd
cnYlXQ4tyVDozM+jg2Q7R6/GQ86yXmmbmqKjFzY8jvX3SqAvpmErTUOco8S4QkOE
zJFsMoT8nuqzFbXlXKJHorXApTtHUz5pyzhGWPgm6bLlkFFYkMp3h1/X29qw+ebt
GeVcimEDs+Tdk9AH1XKMjftZ3SnLU9cNZpVY0WeZ5OL5s1DAv6XR1M+WG0rBi8SN
7KJi1Bax4IiyIu2eF3E929ctunSxdXmwOmc3JmCwC8nFwqA7o/vGkSv4Oeugm5Jx
iTumpFNhtq5w5W7sez5Fw/kaPJJyv1aoIdBNOHnV61F3y8kXNqKgkLc3KBeBWeEy
fQzbjkIUFWtAT8uiT1BW0QAJPbQeWoOS2MzSDIYlV38ATZuWOaOB8BwT3w3Pj4re
92Ba7wePqNFKmvCzXNYtwUHjCUooNXtAaHBQXkZmQccfRKoqXAfFJ/9fQWBr4/XY
bikU6Jn8oJo38NZEUAlQHyMt6OohFve2hALwXxnG1ArwAKU4nya3aG96W5vNXABS
6ozdQGw4NR70fEb3iXQ3bqiTTWP7s69+T9aCjnV8ZIWmZQEtWMUhOSQtjlsuS3sN
44Py8SMEpr9gv3eNDQKTQG+fe8zNuKq8hgvrOvVo9xSqjIfrHgnQ2nInRm1VWtG9
Vkl9640OQHEF0fIAjwcHQ65uhmYFPHw3JWmHWy3X5qluzYBLPs39gt19wKHt9Y0U
Oc7VYTGejZxutEJAhZLRUVU3e4FCFQE2J4N64rspRu04Mt5cBlDIeTMK+JvvOR3Z
B6a+DmQkTLTFBvFRzr4W8fxCTzXwBVQ7o7OkNiQMxHL6wWv3p2If7/xQ+UIPVGSk
MNkJ3OzTIqNqU2oJxTL5CntpoL6pxT0y90WVD9wrIuh012egcDdlWcZ/4R50K1OL
UecKV0HxyqHWvG/0AyN2O5AR2hb5BdNIgVR3m1dX1W95yyRz+w7P3TRnUPQ7Zqww
O+8IvjgxdtHCIp7X3GBJCntk8LQi1QEGR2YMSGb/koYuQJoQUDu7wRvJIx8UiPO2
5LQaBo2WTcUX4D6OKbMNKTYVTuaNVkkcMYzr+C3Hqlm91xXX81SrLOKewD0zhSai
OvGvfdSH2Wiy4kdnUArTFxKS9uixgYn4GJafra2mlsE3ZI26HtAWmIrklmtAiWyx
fKp242jC19WT93fcTWykTeOsTiBR5vLyWzBEORQR0NMd0Em3cAJgdFtQa4xXvYOF
pGlItaq7+7EthOGrNaQWN/ObOA5XD+dvr0NKUE/hcDlTnswQ7Lbf8lbzs2EhfPT6
H8KC9CjzxUCQCcAm/hEqu+dTH8np+w5fZ0TK/ea1g0zRCWm+MaT5Vf6ZfvScWSVJ
eoS0TKBTbNINVTkxKagQlaO+uyAXWk3D9vtTF6gILB53NjJ/yfd6MK53FZ+iAHGb
LlTAWGnmQA5y51ikCsMMzXXS7NUFu7H2lZrAdGoCu6Ecwg62UzkWhF2YdOk+DkX9
ochtcEh94x1TDWF4v3/hVnjj0ssBJOB5k1e+RDPvpGnu4vaLzN1dIZqa7TuJiJh9
+mXFaFMwhe0vzi7eP0/3E9TbWSxzfTmB7Q3WNEtCkVAR+5NuWFbmBCfhJNeakWFA
GEFuEsAN2gAdJ7MUZSD6onwbIPxHFIqKM4fRWFRsmpKVFgOxmey7OMZlpiQrZPQn
XnlRh3LYDSInaEqplK8LYklTXeR79Kc0/mWj22O7j8zhEG1sMY4fuaEX0AZpzLg5
nJs7QSLtyZ7mHsN+PDZBwEByqF9VbEnbsxCyhE4bexZ9YongNdsXKfmavqcAI5G9
vTa74hA06tg1rS0VLpdiAEIW5AC7mU2xYDhe7JDUT3esozbW32rFRQHDf1NT4kZr
X/mmSsTbWeIIBfo2mEguztH42h8Tg8ZJiWq8cJLGV6niERRjrCspPb8/Kt3Nrnhd
gDQj6suZRW+Bcr/SndyySebg2PNVoVAyi1ciLRstJL4MeCC+9DXHvI05as03/vT8
6iGBb6cZlqK8jQnF1ml+bZxnxpxcUCBkoyZ7o6ukQqm6NBGIyomjHpm/NGsnt/6k
5tM1//hQ0ak5SwY97nwvxQ84FQQ04icrThl/cLYisFDReuENN+NXiL/NDWZHwmbb
qq8++f/arSILVNdQt8VT0jxfwOudvEuQzRFpz2g8Li7Gt6RD9IJRJe1sLecRaDai
WKdREi3e0oPOvGL/+BlMMKE99+lfED3Cbk9L45RfKgL01KoZqCBYvRMHU5zQgWos
OgsBFYxR/w7HCfkFimFMAppC4L2ZazRyUWnNQLmdoNepu+kkhmjJrCN5d++zeXDr
Mw4UuODSuxHmO40aqBFIi/Crza5a3TiFzPfd/bU6+KXeNph0SZsyp0J1kqg73d3B
2LiVSUIUmeFm1klmEJQ/hhSKGXON1U2t25eIqsywqbaiOlYlrBQAD8pIyXDLc/Jc
cCAif5gyUriB2Xa7EHMNCFJAFogJnvF82V75rtmlHGDBOYWJI7ewCM33p3C9cPhS
4DJiPQdfuXiNvJHuV9Eh9lmBFGBVJ071gvYdio2qkrRwAu5ikw1f9IChouzDUVlp
CtBfwPqJ9bV8dbNehTQForv4moXYWzkJZoc0Uj83HLGo7IEcP0Scw1SLF/kln+Xt
bXJ98aYPDyymgfCGz1NvX3N9cxba211OjIy7ZZgKxlowQZBBjFm8ap/ys1ypHbfT
k1KJHtCDW7iqRThc3OOq0g1PfpnrCtH7tqE9B/mgAgupUSMMCAF2p37WXlswNowi
X1QkIPNqju0cvaOZTwiqbrB26sh5nhFQq3bKQZVcMP2wwVgNz+xKjwOudgbMjV0z
ndl31K/fyX/PKJGoQ7FI0YW2raEXjJfgdZTBo4YTdubF+mV7fHp00Bwq45s1d7fq
CRLC3oAquxR83sY5iVeWWIXB/iUiFtqLiwRPxcF0d8gXGe1UKc/o6+t0VNpw2+7Z
2xC+HLPEo6i8K1fL1qgGrAk+iXVwHQbflu9QAlqrLeWncNFhoLgVavugbBcinleZ
Xy2SkzosC6Ydm0RnPLQRPfMpH054izMBrIAXW7cd5UtBPB/o/bO85DsSqZrr//ht
pLO30i4PGSRse8XINQr235MtSg9tcEDh0u1eaHcHN+n2m8UENXA7Ujk7aioPPMe8
AsydFduCRmWNHgg3veNX9QNJBX54Cok0GZk+ocymVMOh5aTRayPfNg0Bf0SBPBlu
9ys2b6KKKkACjHQhAJ+jcWZQwnrAzi4/JHpIgp8VKQDGEmdpKutiFgsSYVnjsjj9
rckSZCaV+nxHHQIQaG7y2cMaA16vgMKV7Pbz9hHddGF2X7avBu2MC9avTnwJoCE7
XO+6YG1WZKGc16VaZPT8BlGgIcHm9RBJasMH1k/uU4dR6rgWT6lBtXU49sZkAmOd
kTYUBO7XkDJGYJC1S6llWnBFGq+vJ8evpkj3/iI3aUISLhbTvHHMhouORsTWkbaw
lH8XnCayHl83HfZ9JXXV2Sxk7y/7TLuNpK+KgcyWPyGOUI6uxrtH3TcM24KVgewg
4KrYjqm4yFSkgXpRoVAfVLW9hYJYBZCxw5s6nzHgrGfz+lslXqpQGLfKiL/AFuz6
Fkr9R1TFoh7Bo1XZBchhEbxVbaijjoWYpAR2Z9Mwf6kUsG/4Tv6mDTagaI3Ytczw
jGLQBe4ZoKHWkUQcJhCKir/N4hoKxWZfvKzds+8E5J2OhOjca9w4TZF5A450sCIK
+u9qrKh6KKYbcvk6rEULKVH8WwtpDKyFTvhj6wwSKCpIRv5dY7afbZSXNYZCWDsA
TgvkGZH+FCGlJCoXWvl8HMpRqamqur16Mh3fG6aaKcGA/knltGt5mv+RX7ZNPJ2U
7r58DnwqyKHiiS8rWeLEp3UrSoUuBQKNcxWD8jl62iY15I9vDpBtOUg41QbpuqfD
TIL1NniwEDLh7udfBgQvopGZRdQBPa5qslheXQhvTQXwA4HMrY1wlNi8ArK2OEuA
WnhH34/lvcgEQobaZyLS7/n6blZsHUduL10EGPRGSOYurbWRvO8jUp950Kcxiw7t
GSLldwR2mffCb6aTwjCPAiKOPzbmlwI93N7jgABjGFJHQUsQUP2iWAXT+clfeY1u
7uYNjvyQIUROSi5F6SL24OidjCYPW99PMZnkt3IjDra+ejN9dBFUSjpWeFOlnf7E
qFtmQxTPh9AqzGf17LXhp8Cb1rlOS2/mm8UYreLaGHVXnT2iqtT5vMOrQahQ5LDU
l35F1c9oNIA6hWzjrB/+iFLzVez7c2awS0seDv1Has44xkLO/VsVoUOW/Oydi6yZ
i5RIjwd8Tsg9ovnUYFQJk31ZuSu//bqo+mnC1uFkTfhCFcVB+E9N1m8R2xjNF/Tn
CHikLAq0PBZ7pXuy1iD9KrF//wIxhtmKdH2WktkhKkIt0u26Usvk2Eg0lf4FAk0H
dSQtLh8HitRwqdRLyLQlhn1ozwgkG+2epLJvxt4ry0TZ0pzImAG3QAWZFcHlso63
oc64svWYUMCRv6TcNwJVNxwPhYvoah4TOHG2L2aE8S2eZhW2L6c8wdcO7Sz5CN95
vwwC+kKzBf+vuws5xPrAOoCdKplPYn+bT9FzEFYJemgcyxKkuyem6ZJ800n/5gnt
Zvn7emiracSPLAkZfle11MryLFp2pct900cOlXX22Y85k1kgBVdqsSojPjWcsikv
Q0joDIZEoWHt+lEfeg6wSp35RmQ0vtoYgrdWuMzoO1yyX80iN0sCrgRhReI2Vv6A
AeXlrDKY3NMOGPdBxL3dGiLMpYN+AVkFTo8Q8R4/97BH0w/suQKD6rdzVi+IvRCJ
azZIy3P9IhLLoL/41TEUZ/t0TayR4j/GA+8iOiRHp0wMfSXxsztZ5Fyn2YzjikxQ
6/V5IXDuEwylViG9rRBe6BF1yyyfUUpAkCZ+Md34eg6yHigfOkimtiX+9V5HHBq5
u9GjeMh3NPe1/DiDLFLEdvKBIUqji/Cr5gqHt1UGc2ZF7n8wdcFk5vUA2pv7TH+Y
pVGPf9QHrL3qTaMqG0uVs4KYOUQgAm1WrqwyyLz+FLz/ZPU26OVK6CZultf/+aqw
MUREJQ9z3+b/4Kq5IkkTmer4roMc4ZTldxUobMpFhAazbgHmh+I9xyvqZHbvb0z5
vRAdvErom42u02rLGfNZP0+v1zsWepYPPuEkObNny4gFzxi90hpOVJKxxdeRev9Y
l8tUXOcbC5eC8wB1C7m7Iuuhj1cviSXYZ3/CZqvPNCi2VdpfkDOS60EO0jg9FVH0
ReVCLvxe9xPlbs5u66rEApYwkYjbCr/nJToaeC64v5lttvvo8TFLBPdltCNRwdu9
arz3WeJaAz+NB09GXpmvV3PfxpTk2trVyWU9yBcYGhOnJSzjXMgYmOWRpjVRr5RV
/d7dlynKb3IzLDRLlJfatMWFLLtIpbinngFIQQRNKWeSX8YFC5zyPZa0f25lQwkE
Zu5caNnt6Jw9Y20ytoS7YEaJqVclHNn2omMqHovCCKQucG1QiIGtBTubf3qWb/Of
v6iAW07gL+9TJ2wYxk0voIvkQXrACJ08yK55JC8KDRf8bQ1Ho5yAXKvhxdX3PlIv
GfDm3ofqkMliY+A+EV+nl2Gf36mzXNbK052C+Y8R6B/0mdUYPhbUzbHNJjbyMXka
J9GL4oduLDZyf5/WTKs8WO9VAUFmKgUy8klI1ZL5HVOhqscEgUn+Nm48AckWvZi9
XSeFII81MMzwlqzYd1UcmiN14kq7/W+IbreUVXUxKV1tN2bW3TiO0m3nqSCrZMJn
z2wIkzoWMyaB2CzQzur+kZF1bHdW/QGzQV/TDqWTpoyzFUMSzNkbweDXl0YprLX8
h7o876EamALrjp+Kv+fiejRrhNCrR35dARpAdZPxKwU2J25QfPM8oEX4xCDeuKG9
wU2dpRPbOnFANiMdKn0rSaFoLP6NOEdikwdPu4VXYiDztGG1Oak10ekgQepHO6uv
nbJiPPa4OZvpiswN3vRh1kyGJCu8bPSj2WIG/iw4CSxO8SjCXZ3r9zJEilrxlzMs
Teq+tZkuySA3uJX/TqUp5mOS+Tuyx6ELdjXIpZ/GtTct+iyo+xW+Jv1tgZyuH/e1
SJVuq5U1GXV3YIA7cRNbeVz3ihDH99olClFWN8XOoWzhjb+DLsMisPDGXdvym+Rk
wERRMFex9ijHp8QWMaOB22Wlcoo3c5lWZcynxy4anONBhI+TcaScOjMcH7+AWWD9
aAuSvS+OnGGL5nx9RvzhytlZbYuj4HlJCCGpCkglgnneiYQY5ieFpanihQLHHaYc
FJkRS7mEuuWw5ED5zb5LoBHwCu8GK9gjehSPojcG+TqJ2Lpw7xdTmTbR6tOspeDM
K7D5JgqbV7BiiQGJYPhPBWsSicGMoORJdxLNt27pdbfWSHeR0Lr2gshfdDCMAQaS
kdaqjiCRB0QtKE7/boZFzMv6WST6OhO85G15fwFjvFGJVuab0ZAN+M5Brrn3bzGp
FuyOyXZs+0CFFFpYPCQ+M58S0LeXeCz3ae1BWkGdln94cFzhT6nWaoGYt9alwc9X
yFkPaWBADsXUpblAymU1g7JyZaLTkcCTycPHFYkBoTNLyNs6GKHAFoWKE67QB5Hg
LtrqW2GheWTPvflfrBuXr0mDFP3pbVmi7kJst9LZK8uGNnGz7qE+0YKPbUL3pN2R
Ec0g0H4Dlebo4fhjqrjJUsalYwqippisKlHTNoEc5quf3EoMXSgk7j6DAhW8L7Wf
bRmjNk4XYWvTuY+TP0wwcpxACzEfTdIxgeBvM9hNJoCg3zkHozyjxyRDbHnVaGbI
s5oQMmVoDr5HbwILlqMiExuC1W8+GQp3qpbihB4f2kNW2U1SegU9rv30a99XSMT3
zWEk1xeAv26pdrKV/H+o02hFnkEU2o1X05bmjKMuZWRxGumnNUeHdK880YMj3gRH
E6U4wFFk5Ozs6p71qXF9kqFhEezvxq7EKvgpn3fsWh3K3r2RZ1orEZxsUKXG6T0v
MBYWh+VbxylR4KsJlG3hVzvrprJN8UEx15EaQQ2fJ3fWDLbvwEGoKr9WALZe1vge
yxtME5PdLLAbHklZohhrXRNk4fju0+gu52C8G4HJPwynz/Ib4okI35n7nNJZBRTQ
/FkcStaaS68L91fFOA/xgTaOa+fdPjVkHSDC8AGRdO24p3DRWfiOAz1/KPBdB/c7
rqfOlH90NHoNZwk48mvmm+fntUZ/fbikGZG3Ot33ClQR+vPW40j3XpNzTdJJomm/
qf01/JXKmP6WM8fMkRQqce6BYI0NtV2JGd0fkRV2czRqSXPGXeOtprcySn3CHCKZ
gEhMkQDh2ycVQE87RC4Zc5BZpCT5TasoFpV+4MosShRRrVMJ/G9UyyoqTjNJ2rAp
XGigyVYH6019DqRo+rxyrilWoN8ZHpEIF2T6qPYbUP359YzLiRkcu3DPDstd19r6
w2iT71JkaFRyAVU27ImC4TNccmCAa9tGTza02QeS+GOF0MJzheyAKajVUJr0siye
FfyXNM/yZMms4cVhRkHOwJOnEygXdyDzre/uQ2NDSje8Btw1mrnMVP67X31dAHNS
oMXXuRDqRFBNL7oIsHeNeePPdyYQMN8A/pNh5up0RSr2v+9xXMkJy0Mg0uLYFfvO
UDgGATwwCXHPHrjsB7bzVHJ8rEnDYLgArLz/5YY94oUs5IdFWbihOeeSUuZN3x4w
rsJvSqru7fuyclKTvX9RFxnDoLEjZhU8NyGNI9QxR11e2LTv1brY6Uat2G/jwWCd
Fav9nNx4t0V2TUyBZ0ta2xWJNYcPPcvcVP2aDngjQ5pa79CfN8S+veLjVn7NdSMH
hBs+C72ea8Xdih1s+tlmiPhdUHJqKTJPPcdUNs1mWjPKp2zYr0tKRB1QXcaR+XPk
Nd20QquZa7LYxCpTsaGoj5JhaDdO76BOsq8PkTp4pgRxsttJgbfScrKTstWEpyVa
ONpNTk54a7YhnM3wu8oeUXvjB4MGfJg9e+vPbXMuh2l69Nrjb5Cy0zGsa2V4CMkH
k0so1eptDjG1gJCQ1VDM696tY1g35A4EOeyv0HC2pS7HZwOsvC4HBzlYQ/XK1ltC
RsHVhtbjegBtWlzfItxZNgQXWBIMUKsUWJ2Ov7gi21sJ/ipKq81koUEMK7577t6r
w80hU05CjhGwmWeh94cN4GQhrGITEGp8EbPoHOQX1mIxa2BYK1U2iM67o1UqWchh
dkoE3DcVx3yUE9h3PWqo19YlWIb6QMGrZFAxNAvYOLBkpLp3dt/5I4gvxGwaJ/cM
2aol8wPSqVTaSpsUNq6C6A/gqHedDrl99uImEyTSCf5FNmCPRAlaOtfQFR51hpvE
LgLMB0CWB418Zmw9keKULkWch/Ovr5RWlAfOWiovLuXa5IO8kh5V0BLFBoi39TPj
CAqLWdauR4MXQTtyHKSZMeF1GAwCf7T/G0U3VL3MbSBa6mOd/xMOhZLpJ/Dc/R7l
Rd0YlFhEV1JQ0ZO8SopOQb96jWEMEkptvSiBz1aCkGa3gPuansAIqDXixqCX2bIa
Wdw0s+VkUv+fT5/c5j90aEqCVWt1cH604k3llQTkYcJzbYthnZmQVDxN1OyZgtJz
GQMHSwtedQJXcoz65u9jPZSR7zrEjL0EYn4zoKC4h0FG78wAmyhk0Jft38VgS7va
uvF53x0eLBsgETR1niTseiLRA0XGoHzy9qjJD1BTXjohVxb/0UqCqrSRLBsLHa5N
f3zbhn0X5onKZNlnYDrUVs6XLjmB1cU4sB0gKlPxZkedsjgHdzRb6pbOqXcxlXo4
12INZWHOlWocEaRy1w5DWEAp1692QZRdf8P81nZcbTPkrXZJf02lsCSB5NyFEphP
+JEo5tB5LCXXNe5f46lhxVmuJG6wHCHvrid3rYlCgV8qzQyN2rSqQYd4OMQN5eoA
GTCwN4R+ZHxIDnzqBrUQiNFbPekUrKvc9CMm3CjLyzn7L/oeF5lGee0DKlO0l5nf
gUV6wVEj2xusrNY1x5F2/ht5Ce1G/oJDLK29gVzwlxwzJDc7gzmwb56xXyWejIMd
Nbn2OklF34i2VS8rKE9h4aY1H0eb3OoBnGmOfPZQwotYdsPo/nT4XOWDxQTqx5AS
5lpDUOz+AMHP9Bas0cMmjb/s+nixGrmwTAVCW+fq3w/oAgKSUtiRQmGbrppdtiMh
Akz9A1pT1fwaZ/U1CxmSkcxoObNvdBlephJA9pxdoSOgiqmt4A4d2LH3ZLOJw6At
IVUHOE+TfJc1Sd1z55LFRDhbujnyUJ/dVGwd8YEQ3hNZhjhU0kIEsK4+T1mv0tKc
cRuGAUudPFu6b9TuqyYwDPONSmA4SwtMB66GQj0qJb8mMecH7lMUCQZExDBSU7ji
w6EBrfd4ZDCYtxtGYL4ROF1QmdluD9KPKlqIcKXc93YDNNGYqS/oKtP93/dyq0kR
jKBndRzZ0ldNB65XlpL/5aaQ085qj0x3SXbS9SC0uJSe1HiIDvADCnXDXjTtWbHC
FgyetHwOGjlIDg/uyXJ5jAlNSTWsNWsPxnp8F4OoXrDJxla2zcWQ71l1Ic9/7df6
agg7b41fbAdcG/Z5BWw/wC5zCiYQP3Vyr45b8Lpp8YJ7RiPlYYMNu+wRUeycOUOs
i0K8MsG9pBEeMtrGMiVxGnS7GrXVD3ifmPl5NrtSt9X6KK6bWaW7w7RQxBpTinNc
WjyKVwjSumnE2mOatYHnmSKPBMlHQASJLoTbGg0Dmp1uzo5QRYj+cjw1u7Z7p0Ps
yXFB77wg8MNEgugPwAqxT3v9s/akKFEcEEH80TGyJKbC7fLEUqIelHf/lplzKg83
QqMlvdFdeXEF/YHCwJYpq+DhH6u1HdpHF2A7mvK0g2tmy7+QzYDP2fy4GOnwQG9G
PNYOn7fvviPVFBmZXuNN9frVYlq8u0CXwUi48/zTS4+g+TrMZY9VDLiRHo/Argk8
BTVES6yODMgS/63Qq5voAS3gy+YRCmIiYmlLzhoyQjKFZydoDJs+I+Yr37n199S+
bTqisncZqrF9kdPCPE7mzrENckNQ85jAGHPgm3+SIoMPO1fHAJNpfuoXks2Sgv7/
Wdd7cduDjAsopFerR9M5Q7JmECo0/ATR1CTL8xOIsD53ZU4na4ExQv8wkdrWegtZ
U78fIN2HK9CAmV8rb+CznQZiDS5dk843WFwZXjmXAd7jCLNGMTWTKUXxqPW5KWW1
XjaRemMI0mlLH/3nf9aV3nOgA+i5wymKYdO9Oo4sPI6Og8pKtI0nlGWeQ03x/iIt
Q9ejSADknaeRbiw8LkAtfb+WiDG87fP5sgddXKEao4I68uuJb9bIEHm/9bphMdLI
IxjC7XrOu5iNLHpKyVAe9X3KlmsHYNBICB1+arcx4AqFF4yMIXhybB0JkBjSUvwH
TU4LldO6ugAUbFWTl/K5qdkAURQKozEjUcrgAx2G7qtNze5P+YFRJZACLk+jdLSq
nhaBjUYl6uOyoNEcLuCUKRnCtkDVGDEfkKQB7KVQwALzgCQNfjGF0pt4Ml+ACQeW
oPKmzclkFEGtIaF3ReHv8TYwkqBhIWJL3QjDN4rrZFxdtyham0bcrrobdxhX3ChZ
8K5xRfk8OCrEd618TvSWNPJaAy5J3Oeofmw26SaBz+pg+krZ4VzoEblwJvjMLryr
RfrgqRMnrfXJZ79Nb6iqGI2Hhmpoj/g+fdgP2gUY+V3iCPZaCrQLVcvkw0bP7ZlS
K3pz375EC3Bw7TOGt13+S5DWJHRdfSzlCCZFpXMhco1rgS+Ur8Z2OxG345+vDbqL
p9uKM0kIo8UkgoKZTHsCaxd+ICuE0kAJYS1GTPpY6D5EJOObJFU+o1GJOF9fdsu4
aKpUHpKm6OcrH31guLvZtRlwPcClSPH2dXYoBw9v+oyFtDb32F6+fonGS9QWQkG/
U8udjwHgVWO4+g6EGPU+49oPI6fJ+mrn94bTgmCU6+EpqJOCRQaQgJiCDPOwgv7O
5jiFBD6tF4LXbPOa29p9vXthYqVCyyMS0ySaM8CtR58ZfePptChJwUKmVxGxAdVV
ZlV67xIpK+rYp8ldQjhhfLZqdN7qkklLTRukh9taLlkcNcNJeHNyGODTPZJXwzcE
6sTjkfJbzofBATHE9lJJ9enL6DV5ugDp9Dxvhd6AHxTu8cHXCyV1t4EolVbyNVyF
HnhQeQknySyMne3sCjhPIZbUEGPB+vsHw0pdc0g1dAbidM6bDvEVrEh/7zoNljK1
kClVoibDbYP/zGQcYrCQHiCSR03vTYQp4jRZZNXAxcyRT9bdZTXIeJJBXl/UOIEq
+8g4R0FfJd6qp8p6vi2+vxfithiJqrba6DhpKkrJ4COytEd+fimNPPNe2RKvF2xV
4faomyVgAeQfbXm295QXuxDEFRuXdnMM3xmUOZlx32RZeLKuMLcfSEwy51/Ure7r
qbZIwYbuSKJMOk71a6geQ5++sJBC4iB6M4FGm9o3wA/7VQRT/eTrzzVTsFKy+wBK
UAbCWk9ti5nEfpnFZNJQK3ZTS0PQlUPRWsHukFJRY3g798EskF4xa8WobL35zkOJ
uj0cus+kfOnin4Zb29sn8HIPeLWaW00XqeURSRfHKNZHSbsOKp2rFbVqKD0fkHHd
nJnvk//D2APSpvSNXzq2F/zzvvZJM1t/b0CP8OGkDcntILnd50pbFL3HkbBlcGpW
ah1Flvv8928j9nCZwa7EMg2SVM+J5YBr/Ppa5gF2fo7wCvKYLGNV8EkYT7Ybt/FJ
OX4wQoHkJOBb7p+QIF2dgQcpmKGM2JH5Nc7clNGmFVq+uBcPJuWLJbHbtFauZcCv
FwZvoA/No36Hsj6z8DRlGgrR8+XCkuMAVJhIH9oaM+mKAxAu3BkQ8A5h99KHJTCV
dxniGSM55BYV40WcF/UahSeXwDv44dn+M0TtpQOGIzAe+QNIRnjrvw7i/Jp4x3sX
LEZ8oNuREJqUYtOnHbG5YEfGkVED+Iz1kG900eO0inH7YYS/1oclMH22Mbm7l4kS
64E9KoGXBMAe2CNOtQIX3Idm481RunK2tYLano6lVT3gq6cQuE4lHoGpcpJSJVdM
HPCfMS7a+QPRo5/x8Zyjnbx8Wwy+5TBX4t8wqqloE0xnJlv5luHOf6C6J80VhZmi
wIyoCxOarPxsMoSzOFRXrrUKnrGn1fos6AxdZsnRm5ti52etaRecFln27t7VDYCc
fDY/ggh6MEj4j2bn32aRJ3zMkKmY7vcVLX1asUAgJIo2OgBCf+AFh8H90X8WEnuB
KS5Oah3bQIi5S2wo9pbm1OufLHIkQ2Go58n5e1N6Ut6EgcEnp42b/825C5te5iEK
VC7M1S+XHkvGOqmgLE0eUkARNM3cVBOVjhDmHAc1gG1QOwF0nPtHGjHdHg8YJoyA
6oT72I2v+4spvTdA9qztGO8qu+ukHCHTK8Ko5rs4RMj2mBMoDLUv08Kt5/JVuhSy
jhbytE+FUI1CIGjfU0eYpp84TcugJp+YNvAk+KbLkFujmLpsmPs9OXa325zSWRHf
ps2sYQzM173rB9NLANzHtrKIy3Xn4uOB3qnaIv/2vaSlb3whU5ZZICLCEMc5RSvG
dkrwxDn81FK3jTmtaMuuZvdABvSiWOt4bxH6/a2hOviO6KR58Su6huPMFVpLoVMb
uz290Ps5nNVH0zF3IiaXa6Hm3bgE7rv04xCeqjsAXQ9sU+WiR5H6m9IqVUYxnu2A
FsgSt90TaOvHBLM5vHholjdw7Mq5pfMlba8/ZPy4pKareoEkrs8kJnmupd+adlBt
iWl/5WYETjK88V2wO8cz+hvw6COuRSfwjCn6lDFs5T1iuLZMrdpqx95ScQAr/o5r
WGmPR981I1X3aUhre0ANq3l/3TPsaBq2fsLbBnnOpZ0i0iNxzYcOrtvfsngj8hzd
LLGbPAhv5tqJu+bLP7ASEgVgidFC9ygDXx0Y1OuCm3Q8E4FC7jpCXExoVxkzsmiH
YwNHgCFfgydAT1Dgv6JqJuJMCL0TqC3Nht1kNph4yw557gF7SN7LTU9ynr2m1X+8
KNEAeJOB49iLqbvsDisXgDL5G+bFy3yrHeQ35Fq8gZaCZ8MBDUvvGnrj7MiZdIHj
ITQK0+uE7kvRBQEGZN21U6zP/Mi3ryNyBlu2HjdTldm7qaQu30Il6j1upUbx11kS
7bIMPVueOGGjejpLMxgKE3V/5O3Y17cO/dWyCZB0jlnbfMtUVngzVT3+Ha+nkX0m
qmSjeFWNjxrsjdE8CHGFN2r10Z2MtHQRBboJ9my8smwFcwl5NICjzbG0iFJBIUgq
gLz2UDcrZ0vK3A3M/OTd2MdIkoEPOFM1OMGNx8Ko5YG5CDcZsj+4hBPE8AgoC2AP
s1E+M7O1uIHW/sOeB6SgEGMv6dsvSeZ0NtcguW+U6NiGXvt/3f8sIuPX4XDURByO
jDQv/A9Oxgu4cHFqOalmpD2R1Rh/X1CkVPb5wKn0s2ysUaeD37+PKNcAr0Tr8B4L
wusuMy+GDsOk/HvOkff0Chhe9/xI4+71ciqBfHf634M0zxF+MA5j37XyThceQVew
zJTLlSCItRbaswnJraqSM4ZZWZ5hL0wTvU5K/mWAXk0Ln9/kozTIUv3ZxtY4I7Hd
9EfpFAEWFs1jF0t0GJECpVEt0VHS8eGyk7cZ97T5ExEaINDdDHA3Gy4KJax612DD
BDgfTgynv8v0xlkiiX18T2hwSU0CKPjSGuKrNP+cGuutbcMGmjMyDa1tSAcCRbS9
n7XPURS936ncqRz4+di8ctVES/lwbBOhN0mg6fBhuESjfYN+zOA1XHWrbFORF/TN
rlEBxwpST5CRGBKiNj5S09+dIq7/ZXabVbjTUyrTBTdP2Rz1NHrVl2qs2Lj96DeD
PiY6P//GnPSK2X/STqFHW+J0tokNaD2/Q4MdUEyByJpc40jeaERmjVfz4nItKUTi
S+v8EZIgBqVYFn3i7/4Whcbz6XBei3NHi/tzFkp4yvFD/IKCkU3CiUAC5m0n7Cas
pRnzExJdLQPn94S9Yg0YdeqA3PPTnaKZ9Fb7UI9Y7ppp2qD6lNtgLAE2mohp3Ohs
cYCrf4zWUjLawU2FVGVHvFI9Sfl2E0vzNLtcSDqigmTxJGro5rFzeaBvWf5vQXVM
TdfBvb4eS0jHjLgQjgUB5sARMLO6B6cfokmPU5E0PvoF7zHgzmrvevzY3XmAIS6s
Sho6fyh5MoT5a1/zDASb/Qyf3JFOvMJ5EniB8ck1dxRH2SHLgc8eWZ1657LVOOXg
0Q73Pfjx1Tu354vgVp+u2c9Wx2WGnzBzj+ltJJH5WgDSPJ/pdA5NVZo639gpXOiF
JWz1S1Xhvzw5ZjuEXw7eFKNBocS+ikED15VioYKSVPITcE2Wgf2VXWLc1fMo735R
pq8PIxw0E1w0OUH42j2hzV2npieZKLQO6Xo09rEhAYafNF22vDog32eap3bWq4tC
Wf9mcuR3eQvJHgc+u2tNgMzv8DbkCiBHPi5KS6Uq+AEKsbFgW5HU/B212Tj0f8+D
CcFUsrwNoA7KzQErooKrQfEccEgLRp/08lPBQVDR+SEPTYd7NRliGMRpCa5eVOuK
CacUVGMz+TApm31Jz7IbP/bgmonuF3+zTHsQyerHGgRWedta+i/qLVxeBrpK5UW4
Z98xWMB9sNqL/5QsO/NO3XD8DIdmkT5GmTeV4UnQq8/9a/OiDe/gSbsMj5B4fkkG
tzauKY63gyrjrJVJAkJdDyQMBPgN7Qkdq02FJwT/Rx7ospE6AuDTcyX9Ip1vRkMr
VCeAlvAMeDRZUgK9ituhFmCMHNoYW9rmpypZlOkS/cQeTw8z77v09JAFyb8oO3Oh
bq0Xa1kFOxhYOFSmtB7LGFEAhoiH5SYwuLNrqlcDKQqD6Ded9wDf4v/j/fWHmZA3
ZJEYz159RWhR2DY8VuxYZMXQPrxPhXERkP0LBiJBUuz2Kqs+sjdVl2pFaXJPrRe0
cpuch38ZGgXlNP5IQemS9a9yOVJm8ZF8taELlg3H2ajdMqxgCo20NaSPzA0fCZzW
Qq2TadKKNRMSDPWXujWuRa4lx3KYiMyXgBmPEavG1s4VujCM0N55duxkucUIL3ng
myHrw9zmZKmHSgG8r6leUYJQTw+xWUgG+9mVhHXUVeLW/i4QX42x2gIW/5bstVfq
Z56wkCV/6V8co62afX/FK6/EGxotD7cX3g34a0dcVmshAu4XpPZjD/nTXrwf25Bg
KvxjQM/i9JOsiHNGtSLg3RUw3gJk/6WJ26RlHSH2eXurAJPTaj8UIXa0KFb+W2Hk
/rzGT8hhUhUW5CfKnioEku/K4AE0kmWjBgn14ONSU0mXRKq2ZqGHbTJ2KNw02Dd1
0qVH1HRsNrdYjqmIdNB+dFNrB4p+NIWjciCytcE8HAbQwDalsYj+2BaVb9GdPYMW
4sCJsgIgNiPZbImBiu+QabibtBff/cHrIG0ZvGOsZ84yRIh9EpfGFIci6balnHlG
ILiGOxtxh5fDNpDjGNiJoFY68kSUrTRmi55aA2gjSKa8ICZMWlpVv4oYgC1ZZjso
nc2g4erQqmtajD/wgYZYqWJoKf5q1v5kl4hHFuY/nnTCsEke+ueVxSOQuaFFU6ER
EAh2FsrnjH7mG2/Fhf6g2K//hXp2IbIusk9iiiAeU8lMGk4v8AdYicyqT5dGqwCJ
MNHahSjT0tXFCiRsyM0Zv7PiEAVB2i+eOOIUhzYfYU2nnZ9z95dXi/Q8YE+CRSYt
8YDYAYXQPkZw7BNdkm70TuPebQtz+11FQPV1s6yLfQ1fcSweY7Xf7yMQzQVMWgOz
8fMXWGcrujCrp0kaqKUyWHPgfOnzALj5LIMaaQRCrM3jXQdwA+8mfwrXeMY696yr
su0e9QARcG8iB2gqY71zMTPDSS2qY3mYslSGCTE9sFrg65l4Do0qUYGk5ii1N3YX
jFxrfF0XEBGSGtVOghCrdtf5Fq09gSbQObtFnPWUsDa7Mx/PKFN9MkgbWt0FXkRQ
bnVcOQZnoTAx0M4vOCt36ZyIijgZAaJOkk481UlCzUI1L9KvjMIcfq4WJF14q09q
J1geCCyjP2bQYk5QDdylkGXhrjeDv1lzzdKfMMkK3n0WpFdc6R3MV1FMeMvgfPcx
njz0AYIpvROduivzo3BDhxaX7pBqqa5PA/LhdQCjYHrvimNkL4JtkThW+xYCPSyB
lN+IqsQt3VsONGtRgjQXjEh5Y0eE5swqXY1cQ8z8yFxMcWc8B4ZQj7LfP+D0GI+d
jriMZmwCGXeDuFa5Jm241E2mKzaiF62nE04OfSppZ03DiunZxxzovWBjvBCpLoQn
Zu/fB1cr1oafnUjSku2HFkKdRzKJesQ2W14E3UhHhdUZOWgIH9gAoIttqA4cQ4dt
tibFSyAEIXvayoFVAwYRpKWlXurDOzCYQd0Z4bBKR1qttSi9nvFDTP/EyF5kmaEC
8/+lHv2L9sGWW7pJnFRs7UK6S6BCfF8QqPUfNAYpd+SiVXkcqOyt03d51LUkB3qi
2HfPRP6e5JmJbBLkjdXT/m66upj/ydo0V8OEkTSeVJnVog7vAahtRCEyg8X6J4TT
mnJ5EjkvSdkmFjr7DKIuprSRj+qc8Xh7TE86OHxtzbVOU1Di+/usVhgetnM2i8la
5lOrrMl5CNg03oI4cZELXKMoTY4AN6Soy5JcaogD1sY7JLkdqTeNKR6lCzITmJQA
wnmCBBqgvE+t8IcZsPhQYgEWPAJ/bbu+uD7dsemiIHuNnWp9uTBz3917ujVL14hO
yWjlSKffMIY9HwnFb4atEJIciA/lOmECPo/H+F1hfhODihChc0wRZK5NsOlunRQX
7W1cOlVWybmtWDcWx8yFpvkzvuKWNSP/uZ1WSzXp6I8waimLfjEXNpfo9lk38LQd
w/5V0RldMAANgNQnhl9dGzcDdlWmvnJ04GLh0W+URmmDG1oIsIuNTq/6GpZJZmzx
/UypwZ589q2kCcdwxN2rRP6TDMG0ErLmyDP5TnQK9MupjfBg/M1jv4f5YQrCzebs
ULhyhk4KB1lLpgEwiZGkUcrC04a8sD3P5gLLUjg+lMz1mXyUMDF2l75lBIsImH8+
pszawZNHIslZHDoBa+G594InH5QloQ3z85uqp0tSW8OUW7HUmG+k03iA8q6FFhCQ
nib69w9vVthIJyEM+ZEkcuozFD2hYneR2B/gpvfgyyoq/FQe8DZ94R/jUYiwgUrC
JJkfpCL7jCea8hQLRnFjql4g/3vBqu7p+8dldiAoCJkV3LzMftdEDDaAGLQRMOhY
H661l3QzL2KsyPqP/NdYJ4YWPnJn3Y2Vb87q8vGmQqYZcUBasaLQ9K/uJkrVbV9Z
FIEjMPBHki5XpFIHEINYa4jhMW/ywz9Hv6PENK3PZ81kl4YpWwzpHN7wjeslgjZc
iKZudUssXUi/WNsAAXzmwlPtu1NXptjDgks/GdnTZemYEqJym7Y7l/RIQ+rOK4lI
6vy229HBRzUTPcHOojiSloc+ZxXZzCMFDi4uO/8Ct4+80MTD8463nctlkP+0bM5W
0fdbc5CON5Zh6YToSJOnwxhy/Ase0fv54N+P7WxS37fAUaehANCkEeKqNyWae4LF
45HzBPBZpkzmULjerVoTUTshfUh7GIE5ZFb3C/yTvpz2Xit5A8V1yyktWVBQQwpU
P9RkjzBr3MoASb7Rku48VsAHI7mb1lz8hlSqwAEt1OdtA2hGsiBNRRQtzPhxpuVC
j+noK67PIUh5SJsmSQ5O/MpBTsHV4TwNafzAEeNYecU+pZxjz1vErQnCRcLsahQ4
bStlSdFxTRD+Hb/ceVPTHFVaZJl/7i5BJGZ9hJtiu9+1qDa6LXH4xSWMB9Q6m7w3
c1xUkIYNnzrE7mU+GAiVBsX48XGDXErqrq2xG2zUm+6ZKIurwoaKK/9cxb7xCOBc
P/h5Ms5keU6cX63XKYxJq+O/GF/vxDBsONO+pmaUCJ3mECOWV7S83hRkAQGAU7AO
XvxrbZuuLzPz2XE4dDI+MYRgayunO36aoGt+yXPQRko86EPzhCZapT8Sm3au03dK
qpJ7ZDgqILnlHZT1r1SSU4uMzDpGMgDScEWf3V1nB6BC2pPBrfZ3Pzvd87pMH1ZY
sk76t8YQVTLVfHtbICcVBm0Weo/TVu9OublUZP1xMM4ra/SMFDZVbUzFqLywx5MZ
qhOFlvjS/e0XGtSrH/Gn7YPiESNc4X3GpM9j5gDQbkMkdwlcXoelI/FbS/zaLCPu
A4oWQgTsxhPhU3vbVVFKhNqEXzGP7tyf6NB3uPd0vA3icgelK+eH09cJvkPhVipy
ldsnu2dUb9f4q/qHrn9CXVrEWQ6R702jWrODEzwObKVjAwk0rIBz0istJzU1mpRo
DdDUxgXJcIajtZFVSXukUczfgKjVBZYkyQKrSQ7gtQOvDUt4xz6K6HQv0q1Xin5g
OX5yUlrdKMcQ48pCnk1JqT9MAwkHkXuSjwl4Q13p5aQycXcCGlfNU2CIkScUgG9n
CsQUn96yijKAm/ojT0uOVKaAYEYDZAWJaUgq+PS+sKOa3UmNOLPgGB8TkoqjvdIn
u2HHZA/kZTOf6nexEa6nNpG1vUKFHcOy2HtPXy1yyjqrvbxDqq9IiJScPstrjJJX
ALaaTHrSOZkJg3X9ew8pUpbTq/XejUrwWJP105WQ8qBXLLbxU5JYnElWZGOHCHQ5
7XuX63QWWlYn4WUWrSffaaTf1ZYnVonj9u+SzOofqywvL5KKk5GbwTmpLvyhKJb9
oIiE+BIY6hZyLqGO4NbOqzN09fXbkmcjoiVENFrTCKp8TlfJKOkOJOCnxbnTMLHm
LeC+jYd23B6+RJj+Z5w1Xsh4dk+S2rGfobhXrHYXPEULSwyiZ6jvZ9xwcBvYF4zG
70jlR1O4Pw2SZLgRxqj8dKAB32C7JpuODE9ATicKjuuSqeqEtIUpNNnqxR4vAPmT
l5ixHtQjbRyQ5Cydf6ATmpTc5oXRzuyphd3USS9Ibl2nfzYaWvPWTiylKvrCN3K+
A7q4iQCBs17apnHucfFAlLf2MfqX7vX2oW41m4SEGq8qVJ1p2GNsb5lf8KLnxek0
nKiSsMCQU6DPTqr5KjQasGoEJ81Jaj5qRy4D1o9tAlOrVfvot4b/4Kdkpg+Bv3U8
7RuRkrriIAc0le6ic1swnpBfyYsmYXUlTT/BtetSl7cZ6gRuO9cBOVcpexPeFoMO
8s2M17JMau/DF5FbY+7S6IZkNiYZXz70vSjzs712VmiZlu5XPJMR2VZD9yN8nJT8
DBMJTU/9WX6mIyweL7XUkwEUh6XD0VEDBD277meUOrRQZwwv8ocVh7sj+Mjcd3r7
gdkAT76U45CX8bz23xS3xWrV/aAh0hHdEgGklw5e2p8hd9RgaIE63NTOfIRaLXXq
wwsbCUiLm33FG6tX+obe0Xs5Axezh96PDZIpEcVrRrcjrVDKNPCYhhptLj+Pj1Lc
1kvE+R7yz/EMMtuVyS0CHh2okKv9CSspQZEn/07LCSUKAIAMuVBDb9U9NgKEgp2+
J51oyd19h86gHsfz3/ca8ebAgU1/kmp0QTRyAdc4yUZMx4QrKzLurS6FlSguau6+
ntIK7utHft9GJqx/bCiNFoCkuVXp+RXht4vM10EDgvwzDbuEBzDnP5REAgNtZ36b
ClL1Ca3knIJ3630mmtzRSJv891PGow+GC/ebj5Lb0OQCLtWOBULHTugvQerfOaAE
uuM2bWepYLHU6je4eF6GxgdIfwiD7LfKlojYiERAkn/7mdScwLBSKNzcT9x1yKk3
SeXDE1ckX8oaeUDBwlLYl4zRlvcTVpciewIpSMa6qb4Rz1fLotYz+yrOz7evWyUC
piSjxw7wA1nY5q0i5grhkmcbm86D74dKL0rRvA7VOGHh9LUgBDwuTM9EI0vcVv4U
bbEitoOc4Rc+2a0Wy/Mp0886aXgKYbkrKP+qsmE6tVTVm0WX4Nt7apNgqslomBs4
1B/vArD2hEwcGsgES0ej0S7saYzRvz+F92LqYxkNCRKAq4sOPmNsl6BO8FVI4/jh
ouPjxbzHw+cgUmzuARQz2zlbJoMtk6/GJ8OqaeCr0pulGzXbnkifjTDfpgTJ+E+O
Qd1po6qCow6Lzmse2frqauryABuTZVqEdn4ZIII3fp/TYOe94ZFgVRaPq+zodjKS
6y6U7zyRVi0YNM+XQAZ3sNVkR/G0ffobmrQ5xq69SsELTbuclO6gN56PVOg71BuK
zYFNL5rj/zf/q3+9i1yoXudNRopKIyf0E69Uk+5hH3XwJ1rFQU05NNATlcfuCdGV
zoViNHeJZ2bfm+yN5UKLZhQ7006z0c70zz1T84OPY2alnw44D1Lz1UDSsM4+hpfs
OykpvldaSpnlXYjI6sIoZzpcSLvdqBUvjIOSgQ4uTYaa1cDg/3SCwKl26NfOMBD1
yxytGYSbr1n3FlJ+MFIidwcM7IZPDPp7INXF2ORD4kguOgbyOfD0uGG9jbJ94svW
Xgm3gZdHvatdHFb+zkQ0Y4rnov3fqy1DK0hLz3oqorzcqcbDPQV13e/uECq1Iany
gI5cXqxRbd65iYvxDeTJeLZvSyg8p/+O4llsNqxLBWF1RldHP9XmrDx2VAHIdHFP
aitMbGDc5dEBlr5L2XJUj1WraIOMILIRKZ06CO+wWNYu0PAql5f2p6RpIoGgzMJC
RFU2wOKLtdI1NfySL/xbZh5CQxF0jzklFBwLYFzzKzSBJBDoo0cIz2/OFT/N1ogU
9JG3JI4D9F5OOiuXIYC7fVPD59M3AkRb6x+GElduXfRBzYPR5ipxRxfmlmt9aIhx
9UbPy/Zpw69AwK9a2ULdEInm/7Cz6ZOQeLwGnpwTlGCq7H0pEIceZ8dIIU7ttiBt
xkeDdVEAhfgLU3N09jX+idlKsZy/6xJ6VFEo01YwC0VPWSr6q0U2lG9yvhoanrS/
YrRJH7N96x2IW+UNFT+zVJqsvMSuQ8nmcm03nkeFbYdKNcr5NZaTkBkCEcQh8mCE
3aru+afSA4Mm4stsHmpSmSF/eJ7qAn7jx5M8ySdyHxaAejI47hBp290kb7xybup8
S0i2n2yXw0oyIIHvJL5m48yeMMVHaRPLMKS+7HXnnwPV7rwoEOKiPJvMNKWt7rvy
Rpq+ksIKRXM/XLflqMuY0Q/Wgoms2k9efuAqYknaqTB53tDNCHt9iXhfwNvdYtSw
7G9/oJWhHnsMpPtmbiVnKTDqgx8mSW4TR2WXi9GQJT67cF6XNBvmPK2KhfwXx7YZ
2QYtAA9mXEJdWwhmhHQpnhEht/OteIUsdhK0XEgnmLbkdBwrdYmYTo4QoT2BXoyT
o+dkRkXdVHYaWOs3SoAlllGeZX9UIF7F4Ex1tqslK3PSE3c7iCED51h5QiZ9LXNF
ujDy3T/OL6gZw7G/zoxJtVeIcjIxA1za952Fk4Q3fybHLhLSP6M3hR4sZLgSgClS
19julIGNWC1GenU3oTtV5Kzmes4Imh9OKVTio7uIjdI8EW54JSjcjHYq9XDybaeS
kTNJ3FCaOiEWXVsfbJa1+RmZlIG4wfELIJ6IVWbinDKxUcfmw8QLLQd1W7HmiPex
b23ukQ/ccadcmBv+WeE4cdgHlMjBC0NO/wFJRpErAsGbwS7XUgYzr825JamRXfcI
TTqoShzx+G/kqPj6CCuFTnZMm+3W6IPEFdLSflT6Zbaq0Hla9I28tyoFEIajafvF
dhuqMKxeR731cuuANz0mvG1N7/jmQ4j+wZ/YC7otoHVW8HFBlx10wjgMtdVM5vz+
Rt6rW9XMn9RU8hs1+JocIp6RGDoqEyqDOACUCgHoUNi+uFay2aFMsg+KnQv1PS29
dWba+uQsTmgEJ3sy6Zbcs4iyZkT9RZMD2xqGHHIf0xqtccgolZxNhqz8bR86Ggn/
tD7Mukmc95QVBuPouFpfLzWQONebgTbqAYBI86hqIaL8ZFJS3+vduJi8fL3YNg2Z
9xGGpMFVH+Ypsm4NCTnUOglrfkKZlfEgeFA2ZYthMN5efk5LHxLW53jSNr4ibITV
BE82U2Gsv5jMG6ZtcGy4RYVlSESD1mKbk+nuoEO3XSpUyy3xeebTlj2SdiW2kZF0
PtZP5TleSRi8oxNtDYsyqAy5B3thpNX0L8TvTNfgxTskm4BAIrVGSaiQz5vCGXCH
Ebw18RFtvv61KEptUr04rh+aCK+Osik+dG7FCHLjDY2GTfpTseevYIo1wlDZdn/G
yGmMXwPUg8AJO6w3nKmcnl9Tv2Xjl7R5//ay7ShuaMQ3XXhurB2g1yyXJibBbu67
MXUa1HDt8suyJMeSCxPs1X1JQbJrtuKnCBAgOH73p9kyhjYB3u5Sb8DGwoXTggbI
X+lKZv/yCw+C6Il1oXxIb2Oj5d59G8/JKsIQrMFbu2J3cVAlC3l1n98j01zUrSVw
4wwxOjdNAP7PH+ZROw4dvmcYGy1YhtpZ5+0Z9RJjTAn/LHB1GRcHdGAvhfHCgA8f
H/FOb29cylqOjn793sT4s6Thx8yDhUqIk1pe1IwVTDobdpnlnPqroUWpapkOOiZ+
q6xGTRtXUXi+ptxIWUnW4biSsKVPfxareQFLcLYSDPqYhwSOBcKsSDNxCk9Bzm5s
fMcUUQwrZu5m8UezXipZFmNEgaM+wTeJqBxEJhInT0P6it50vGatuN0KTt7rKRFv
sI5JXakoqu8ll672FAoXYZqbc5F1UZjGvUk78OqX/j+UbZcqQKoSrGK1UewLEpoD
oQqt38VtsO+PDJR0LLhPgqKZE1euPahbk0JPDCq5snisjiR12FcrbaKEyauYBZ0E
Z05Lpzx6GOVhwJ6m5Gab11K83kw2UnKlPnIUUZ9BFffipAJhTwwL4KGAuOssKHOU
dVcq2kQ8gAHGM4HqI6HdNzdImot9opsegYvtn3Wb669KOHvY8VDEJGMMODYbxjp8
rHNPq/swGe4NV75u+ERJdZVPlvFnjr2K7264tG4mYoyrJDfqN365XpwPzrIMwFXc
U0WAaSS0HXpkkCdQTCkx2dFN1v7Ew7LnLyFIVg8xYjfqbE+1Sc1u1tg5/gBnjA8K
C30LHXEd3RXQkVgb8HaFQLH/bEXcEr50Gy1eedwq+we/VyRZ9dLOhgQWR8XxpjkH
YwFajVXzFeSWyHLl826e9ibGI9d0KkxiemTp4fRHxDlOw9pn4EshL5CWCAgUY4LY
nTJpd3E9pwpK22LkTcapdQC8h3jbd5N5sEz6MJ8ojzF6OlHGc7/+f0l5GY6FYVCI
r2hwcMeu8Qj3FpsBxrK6GOOQdDRd1URFgjOERxebgYSYE2M8exvUttKLomdKFO5N
aygvokDJrE7+/qrHApTrpv9YpLNP2czhpILmx3FTyxdhYmIpJ/nXUftfJLA3TtX6
+PdOYoCzPFnmhfnRc9h6x+FAIPdgzEyh1wi8iCKm7xC1YMB05vjhyjhx/98QsS0I
w3KfrF8wWtplRPzzJ7gtjfW8Sr72GGTTx8ZPKJ8FCsyT+QoCQtA1JABDgT3+36Cn
0TuFmZFxFgPzKElsWevGqahR86Xh5GskJRcomSRvcVS/BsfaYSEDTI4ndSu+zDZA
vPZWhe+ZZrawnrla211T+toIA4L7LczhEioGvPsnvrA+g6BsuhzlFX+B5V30/36z
6F7Pri55gZHIlJzZdtAuf10124FaSFqBsuThki0UskFow95htvIKGf7oq89Y1MIa
1g65wQWdf7wdBVzWBN3PfHpVzWjvCSsfZrq4b7Yo74HI9zTu0+pyUSFratS5gFqg
a8TE66II13baQiYkyYlwqc1GWCqpl0RweY0jzqumrsQsppYh7s209p4yQO7SmLpb
wlTsDE84lxkninZHmDg83FXVJkl2pihbgBclM1RUVbOJbd+Fykc82q5smrKHhWWg
hf06DznmiT68zdHIJ5xB1ROuhFFvPdiGnBhQ80sRS7Rc3l9xVOOGSeTwzX7mIkJo
4IF0I77oDBToe4RDvTSTigr7JJvwbHVCYHs7wkW9ky9YXofZva2m30W7P56K5hXJ
tlafmTE9DWGr0h3PPFWdPVWWOMKQHpmwu8aGZZJ1Zj0RdRvxRB+NzjePPMMUEIPj
UAQyg37GIl45Qppp4LLhmGl1F4WetBoBEivbgtcmat2LFFHUYh6ApyjmcFWsSs8d
VqtStn2xY42Chn0R78GrBJGufxH1lMyTGkTV6DaRq/yjl9srAvbZjh7/Bk9bLj0p
K1uoFW5Gi/ZMEd39eZtz/W+kpv4nwgStXSEQd9lPEX2XDhZX47ryfD/Uv3IeTqwM
Yfq37UVTP+mFW5D/voMzi/bSWCZsdKZ6dm1Br7eiJu8Qzq5+191K8F0mZXTAga+D
BpRVi2JQ8/psz57y8sCRaAwqN+3pwPfrzA8zyxfYYZvb7hPlVpY7FMvvhNNhYmYL
s/iCuXdzcQh0q/8oo+8X48mCpbBeZOghQkAXeJ/VUkEUuN9CaJ2O0Z6Oj7yleP/L
5yRQqG6+7Ln/lM6zAZIFswAEFkZDop5JlR7PSzD56niRNcDNfGNNSZvwzY9mge13
mnzTrq0H3oW/8FiYHUhlStVAYXLxhcz3IrhxVQdw1mFgLhMcSXmKhVMaXm4j4D9l
A830J2O632tD12IzKdeWbWZL2E+IL1zj689Xp++TOdEL6I4FV8HgBHyFnfAztFh7
ZIXiau1kjWyh0HAoblMeQPcd5713OiRgye0upz5W30ME9ES21Iuzyrn1B+JAZ81Z
lCHlMXDLjglx9pb+uie1D7996mwTn3TC73aXIJbSjFJGlwveAaTgE//TL6z12A2T
v35PI42MmF4VZt12X67w53Ud5FzdWsMhIjsiRjMVvOdPc/YGbgIOAZk4b1rZ4P6d
5IPRL+Sy9DgnOlORqjRC43KInkr+tdRdJcfVZqeCbn/0R75w6q+LdWJs3OkOQ/sT
iOACzueJKjijURlpt8U9Z+Fhu57U7fXQDdVVrSBjcReTYIyoI16BuO4MvNduOJUP
rBZ4wTyfW8vNWAIEDeawujuYaQV0C2g2M/H+KQQYZlhtNF1MsuZWTtMmkhZMYtEq
Wn9RoIGJq3CwQ41lTrM25bxbxkpPKvLfXKYxNStbOl2/UpYR3w+DbveDvmfe6jp1
SymN6iGklyDz+Jtjvnhtc1RehDMfD8ieY9vcJieb093/sWb5DV9uDc3NX6mq+/JD
eEnr1Sq8sg3XCp8+MjdzbObE3Y1VQmK8GV4LLb4AEFQcl04KnT1tS5BbLNtrvT5Y
HLFJOQU8/u83SiNyvqBN6v4tJsqrhO9/8itosTwQneaZokdknEBYbnc41ExhPMde
YLKNkSZNKFWZJrUo3MpHb8slzG6fdRpyPxo6POjklW3VU2BQQe9iBpdc0z0+BYKY
y0UurB4C8UbQtVZuAxE5g12n5x4WZRP3xdRixvxcDmzxiXD23EvesWL4rZ9jLE78
KfL7t62Jh+C3HanIktSO2TPH6eQDI2ueDDXu08jpS1aArm7QUW85AjxxEiLXo1t+
f3RAFF18jw803lxAYZKHK+TjUnnDylWdm4rWm9Nr+862qFGvAcqNw0fuF3cGlByi
xtEpK2NKtC0DEnCLB46D6qSttD5RP1ypFiUvAmuY4Erlm3A2JoNakWxAe/IJbv4s
xRhsLE08xslpb37fKn7SPXmo2LxhAJ4UGu7SNuyhOP6lUelXQ+ERmLvR7f0+Xwqh
lZ/A6Lh8ZiWSBiFXkT6wYqM7Ez9RcTZUxwmAGaYdYGRcDbG/BMsWOE5532mXEc4I
Z7pTuDFJEDKm3+aCcmczQ02s8XnS4wQkHi+YXxtMUzK0M9/Iv3nHInPZgGK2rRhk
x7VPJkDGJ4SgrunbiQAydrdWO+VtjWMCRBVig1M6ank10aPbLqZ7wzDcu+T9F+zG
rcnfHH6L+oJWbOfStiS0tEUGShTv5H2qj+D4VvPbdx/xPyuMOcRV/wWuQ71r7qkc
Z/qkK82VEEU7Y8ZfobBqK4t9yF+edAGJRRA4vKb8OUx4xni4mXCyWodIlobonTGZ
Wj7FejqlWuUCZaA1O0lRz3PJc76yNjrPNMM8oQmMLD9XD8Aq3YaKQQBnEyzcboI6
J79FpbfWyS1vI8YXUKMVPWZt5UJehKuVY+9P0nI6iFJFgKmfjDbUqSHnQtN8WWr8
nwnaDW8aMkx1/bW/Ltxw9D5VP1gQTQI4IKvxzGRW/ROM6HkhvSHKlwIO//r1+H9D
kSKBHjM6Wj8A1wJQQL3xK6ns0Vb5s+wq7FMU5MVsfv9HvzkgOw5ZrsIedrUJkAQU
A342oe2a2ey/qs7mZD4w9Fgo9+IobrN58ksdM2c4VgW61mX8TwO9Q1qDieeAJuTG
KVZH7Qec+o5RtyB/sWDeB2VkCGP5UultbCWxer2ECe0ByhgNvHzLnG0dfYHBrh99
BrSiUFdvjZbM7WBYmKHnlBFo3D8cDvktgoq7OXhOUYZCOl460/tje1obHMI2n6vc
oKZWuhSZ/+DwIFtJ4Bf0qeoCDG8rIEo7wOo39DFU0X8dMPGx7q1Cz4Eba4QYwAar
pI/YbuVuNzSP1Bhon5IHcmmZR6aIOhL4biEiBRLP5lzqSIEMC4G/cw1+/a/YPfya
fBA/swD+NZd/f4J4Kgd0d+jdM5eR/dFeXu3kzRoICT1nUzBQZBWvPf/ku6PluCvl
Sc1Q7L1ye/7r6I8DoO4B3NGlZ2MS0xkKlwA5Q4EyX7gaAi2nRTupdFG8ul29vurX
kiJ2KwD7PpBIc7gNnCbnulCABB3Bd9w4242byF75AH+M0Uy2qPfccwTE9adaFo2H
jlDoexxxaTKgBVLkKxrDxzkh1CwlyRrJmrODeHePKV1/m2ncTGwVzIDhQyGMqGoM
2MjoxXfLufF42Bxy+Z7OTIIUpeLSt2BBDsxoTi9Z546Prq5szDomyagJmP7GYWpn
agzhaG9zFHHYrwKSd6y1OgN28BxR3lBBPdqjNr4pG1NwTMtliiNuPJAD7ya0V8+m
u6Sn8+mAKbsR4N95pB9TTh+1HKoAID3DP+WcOQe0ERYioZnFsh5PKyFUw9T+Gb/k
h5Qg35EmSJJJGdBXko2ftqWb//uqGNEkKevqGLD+m2ShBmtSW8JaUUuomjBgp5Hp
V1oAJVzp9yPH2en4npHWqdUGDizQFk+oHRT50tNiLmUF9zkjeuE7Be2sktP6DdN4
MR/ZVNtaflp0rZkA61FKTrqQTXPu2Fi8PeYvFK+Rrt+O0yn8ijUfcS8iFRmurbZF
3CYgDxGxaZZWkJMsppuWSggwulO9BDpOkq8ELSM2+MUZSUO9BEI2ufamEr2HNTu4
iWthjH433raLj+OJnW0fTXqNhWx29rCdOg732UNUjYyK8U6mib56nrnDndjSfrif
07BMsx+8Qtw7AaOln30pIDpHkVt5tXlKcooTLogDSS1YIiAfeyfHfq7ssH98VRNz
5C6Nq0le6rqYjxSnFwnYfm8waD9rUj5t/LVgEraRQ4k3fGRrhkThLX+IFII+Hc4r
Meoy5YF1iMiZzPVp9n4YTM92kBimbwTsO06f2WdE22QAaqBc9AhLCqLGAmCHEQ21
6UUreP9Spn3RLxxrg5RtOmP1iwrmhHs/ca5NNkZ9Dm/oOf1lxK63d36z+rWhIJTz
lKcZGq63TOMUn1Zfupy4OelQofausdJbHcNNohf/ZufsW12q6UHbYn3mHNfoAR2H
3kKNyM1kwqsMcZ0NBjNOl/Sx3gCl/3KGyKFI2QcuI3P/OGcQe4rjwzBqJqVtoHyJ
tBn1PmHVRlZ6L+WblFKUYJBdAl1BTt8wZRFas/rRGEDNkY+QD9ThWOGu/B8mNvvK
hMDEg806gAY0ouapPdus4yGnbFa4WUisqXJBsF2Ddv41zasXsW5PA4mu9jPNltFU
CuN4/ENQL27QX4Bprnt04gV3aQ61IoHuDX2fUHlnOX3gyWoLjDhAQmMgXK7szYBv
qqlZei1aDpnVBeHqnFBhE0jSvEgddq0JD7Q07wKu6NqwQfW0uW1KEPurhAbW2MEv
vEyxwFyirZDUxeUj8qP4mA25QXPQuKYehWZ8RvThsUCPIoz6Fm5BQfAIfemq7/c5
NzSk1B6mM5cy+s7vq7EPT46nPDnSwzwG7n0A6C/aBrTPxNwBmmqoYBGJrysiWqUj
H27AJq8Qc8YC5CckfOjeCEAe+q7dmkZ9EmHNNmQuvhtbDgmsOpumuH2esSZj1rS6
UKGYkijOTeOpEzUPAheM/hBh0mBgxwGdoHOzL+vE0RLTDdJ41YR/LlgBwXpmvkM5
KS5iMN7RRXBTsj1+6PG7yDXh/yMS6G7tSVoWULC255TRiqzTCyq0eQc6V7eAWXTp
sv9A0C3bvPuNn1OyVIVYhEX4kowPGprPoBmvdSsm2kyXcpER+/F4qlkAOkiPHKxt
QtH6zlNp6JXJPxIP+8qImr98q4QcJQwBF5aAEE/OXaHUOEPdyAdwLx5zsPpXO5jE
LULNCEKG/d6HiTGDWBrbZkMoeUI1lf9hmVaK5ngViO9Ree635Ay6ulbwXjXjIphC
IUFV2j9fJRCKpMZOhXjtHhnVCI40SW73KxdMTPb8dcq78GxCjmI+jcIEiO3DgoML
3Tq8HZ5r+2e1HY2Frnc4iQkNwJBubWx6viZ/GlmysTzxcSAlH+plVJlek1PvXNjc
rTDCTwOeQ44M6gxezbM2/9lT7d/SDvFxh393Lb4k38PMCIlI81Uz5gAikBMOZRwe
9cxcsfOWxQFc+6MUESsdKOOShsu17Gf8y7s+4F5BLGHYWVtMCxH4XC85SgHfTR9x
yA0kCPFkHptJTMQpXW+iCpq8g2ouBVsGqfle8QW/I+OzdmFLLJ3xci7WXvsPND4S
PHVwtoti3jWcDzPL36RuTMH9SG3VamUjO5ZwHC6B8njWgNNtVtzgix9Fqun/cJbE
JHFMUrIomrOkvRrC73y/A23vOAKobzxPXhVv4EVpJkohakS5IcqlVfiozv8jG3KT
ybmQDZZMlN6nTpb+JNci1kdlFRzUx+KDiettXQjp0NzW1cKbV4EmQ0GPSD4B++d7
QrsA9bKS37xDVQK3NaNCnIgII/Z9Ccir9ZWBsvLIydP8B7q9vC2Fn+AHjUeMfDMd
B7Y3+fLX8y5EQRycuaAznF1FJy4dToE/Zn2l/yHou8zZLgvUESyxbh8y3iSofx+c
AQsU/6X95BsTsxf+6021swqC3oYb5h6Ikb92iTzoIbGoRWIRuekLh/0LR2xaf8Jn
nB3K5HwTeMkLz/kzqsaXnUm/yoNzi6sEX+ocvgomvIPzTf3C+5zMczWCtBW5mdjT
iGzB1JVqI6bhC7PTaVBeHmFFywhkwZXBmNWVQhJaLr7k728ezo6P59elUNnbeDv6
HWwRuHN+heET9qdsqfp2bM2BU10eeURjQL7wuI88ZRwb1afrFPDbCgYkqFRDlPGT
04uiT527yuXuF07rVvG36BNNsd15kGCu3dSodprbwW1zHZpMuWl+ktxT+a3o0qzL
tqnmu2HVzBCzLZZfdWhZavpecXYdmm/wgFtoX8tRp4GlnIEPOkkYdSu4y04j7pff
4kdhobyM7kahmzJXml55LlgLpn5ACZcZe8tU6m3mf0AAK2tYKp13LG3WNV3AeFIq
xKsuLtNDW7n+fHQaeH6g2HYsc3Qz8eQfpGKqgZURHWkgxaT/RGCUhMCaMcNtwtdM
mRmUY7DL6g8i/gxzu85tlD8EziWoWN1WrAi6VcDJFjOq6R2tY0Q9DX6H+RMsE42K
ejgPg4J16abOzL2qWcvuh7tGpWafaflTEw4Vq3xNFbPOla1jqztuMlKWWLxVuHGr
oo9/SXJyN4hvLVQ0BKL0VQ9yGeNOXGBQDH0jAPdNZL5gaI7rwgSrqcRXQ2ESz4y6
p6z84ITBn7TsbNKImOEUFUmxx49Y6KzNqZubqPCrBe5x0gap2wLP5GQ6ZeydytCq
1n5mTSsnnpGa3lUdSm9HOAzDrG9nqqbl7eUfKbs8BEzdH4Ed3NRrvZjdEVe8BR1A
z6KAi+iL/zLpYlvSOyo/PCYPhK5kDsf2+DePxDbQ4scHVW/FH1X1bB9P6TrJSRpY
fSB0a0sVIrOKETnzQ+I7Br1xPFUoapPoQ2HKvSWtBxR75FnciTwibUaBM3cnED30
cX7iPbsNE+ZnsUIhprxsk9C1qn92433iVz2hUphbfkk3Ka0yFFRaAwHMyDjJeEqX
5H1uShzcl6cJ0OoDn8JXZi2I4O+cDspZlhLxxGdYk/hqBWYTysD9z1rY4VGhe3TZ
9NnNH2j2jMKKKvBFvviM4iZODvCaiBWHWLtfjlv5Z0/5Izy7mUhQorakMQ35oMbh
RKHEqRAWBmeKv6EZB1z/khqYspfKmrbOrI6dx9XBpJDjkont0ExsYZ95SUGvbWeQ
wtjddqCKS17zAmwGaF8rKasZ3kXicrAL+8nsregP39pM89xkHD3z1908/CWgDXsK
ukThdSznD4tYJGuZa6gvCgban/hT9lkkh8AYhuy4kCkkwa3+OA61XTKLL5usLW/a
KG1eF20iFIJ845kWLMuc7n7w4RUT8NnAGC7EmoOjvukKRFkTIUUhSZQ2/lcqpv+C
xJdLMyNS2Dsgvqm19zeNqly/35k7EPUVwpChHkzfc0pkBMNAVk2dRQVVEOn51cq0
sdwZzvyEIijBCNRe7lejFw3KXx86fPBSPlqfacryA87PQHGldUTMuaU28jKkDSVu
rXG4hipbGw7F3Sd5HD4d7AGVcBrV8D+gPlWlRtCunPPtGHBeGpcLAbkgSDS3Dsl9
DG1PQtGUBQe6T6nbAQ4dJ3+pzrGzjF6V9X3IjZOqk4H7rRu7FREQ77RCBRCwQp/8
w56dR0aHotCbQIVGoXq9NdOBWq0vmMArIKTOvctXlCTzSvmsY6roDUv56c+FGtse
YVjiSfCqA6hAWqQ0ZQRi0gKc1yoH3E7OyPQ+0zykspKl/O2goclcbWB4+YK6BcCg
sfaynHBX6/5y4vSg+H0Uc6hkNZR+zP/vtBF7Pm6QGB1Zi/SOy3tB8S6O/lVCWanU
GLwWlzPIgp5RhnwR02iVjn/zIvfhtbS43bRgpReA5j+TliAUMxPEnuflzoygBXB9
Hwdfwmjj1dPAViPz4MQSfPKL32R/wfQiLVqMb270lxlAfwdbvPxMGHnR7AMI03ow
NyMtSHV1sKTxAB4KWpwIfpO7ftcYmGICHC/GN17N3rks+ishKTK3aZ7EULwAViAG
uMoMM2udbsNdWMhB1Fvz52pupfYue7BXr5Vvg/POv7DHajDFbbLH9sxZxT2ZWas+
l0JY/duaT7nbxuR8Kvbqx3nPXbE3KAWZ+Ivsn7FhKHU8nmshOApUYxtfTvf0ijjX
7TRqHXTKT5tk36yuo500cxbFdpDTA12t3MFGS25FwTLbxMKb+y8yuBfj87OfPU08
gBjylHggiksqHiwNdd0xY/l29+HjplET/mN5H5aGB3eLL6NqGKFtoMn4KU1dp/l0
H5+dpGfkhZUcS4QaQChqSawgzpHRWAEp3jOceqXOxzTK+5EQ9zv9SZqv/CWYxaGq
ImqKmvOB6ae+ZlzJzqN4mZektqQXR8gBGj3c5KRtqJOIto4ocZLiS8IFqlwyolGN
KkxVc55lP5OHXDlWAb7KNRbnoAYx0LimE/g3CFG/x16KuPTPvYX/YKPvXiMqYqgU
fTniWWmwLJlBjavyxxH7FcRGudKm6/IEqXh1iKcCCfnrynU7BKPY2tTVmVk+fj5z
xDNHR27AsNcS82m9c7lG5F46ujHcRWFdK9OI5825MDcdhr6nNtW8JbyXP024id9z
0z077ijp7iwl2nlN0+Jbn/U2AEcZWuiZtKOQgw+69M98HlJ46T+pu/B06IJYCiJd
wMCQpVd0hgVw7LcPlZ7Be1WHeYRhJREC9vADFy44A17EY+salF7M8L4sZfnpyaxC
IXbgpNKo5erfPP4BWaY1nHJB13KXClOyb+ZnxpfXNdPGmLDR1BdkHrAtanvERt/0
RDq3vIX6M1fJuO4lCaIZRZQi6ZWvoo4uQe0/LcUJDg+77TViJ/i83Gj4pJfDcQhI
VbZ4CWgrE55GMYbAeO6piiireekXNMgk7y18OlcpFF2OyHpfJ3yBhi3Iyd0FzZgB
u+L0cyIxcvDjwF7H3ZPVAweuzAPEllkOjUmJParhMO2EFgZyEjziIiUv74pkq+Ra
872lC10/Ltc2WihrQAHT92eC0syP+MWfFLjD/2Jeq0SbiBI/eD1TVb/xsYsLBS9c
87OQMTpk7DjN8ccoehLPETXMoJkB3CLlzsySKzzL/g9iCNhsosXteWbAfSTcGQ9A
JF4vD+LIZIHwqzRzn90MFi7L1jtzQuEKydlwMC40hXhVKZbhzTZyLT0aGZuMWNUk
Mv8dT6HUfIuEOjF9b8NXrjkUAqY2pp5mQJe078iBvxjudjoyYM204xdX/i1/eu9/
JXbyu1RUPdOk+OfS0H1VZVY6Bx404mQ9hOeF2peNzAaLGzYt5YYnDfrx/tBcOqTC
HrQW0zcbpd3csRLv5i6PhOniBIzllWsGRzHtAniXr+d9JB3xf4ABzWcoYcrayf3I
OZPZLsl4PiVUgfUemMQ1vzO4tLYIZKWKIupaIuwKlUKH55MI5WhKJY+/p/FcJc6T
Wvt/00PwcRP6h86ooueAktx2HXViZLiVH52loOQ3lQGakUthSRucqvDqLuG0PTLQ
cUpT90NoqX/EWYDkEjQkG+VaNHrzn6TIIlS0smH30bjHFTlE4AbdKoC51TgeqdDx
mQXq7UttlwarCm6ipiS+ssWogiMaluu4Id6e5Y3gRNxbkFOCo9jawsJWzCcc0jLR
ED8K/7Pbq+h2aT7l74YDG4ZgenOXCSqMw3iIJe5EiQ6d6gZz9ifQMqB+A2n8xWaW
2J0MXMSjmtYzA996BsnAy/0SSUgWxFpjH7TVHAZkNLWkvY94VQspgBbmwXwgxjzD
o63DAvcFI/5GUx550jJhCZ6BONAJo0SWrAphefJyEVdv31K8y6jgmjqb05ponPpa
PcK/xKN2NkC3b42qo942yGx+4po29yDojP08gWcSg/0wWxH+BDO7eJfeVurUXmCa
LWg4VGvCEdHXj8g3D3CI+G17sb78qLAoZTCjxnfqj3m/GNfbq+oBMraoofImRu8P
/DpWX5EuJRIk3CBFUV65V5IIpvSvsLkZhX6UQuZFC3UIqxdjz80KJ9FLWoPsK/t5
8tTRtqq5YcCxRmQ/EAJHG8UKGI1c+Mbv+9AYBFFV8Y1yRJivmiw8AAg/yuaCnwbv
qsRbsySJnC8HzZ/CAjxkXcCgmXI8mjmm7huARsLYjYPIYPzRoXzSBdQ5g0Fi+RzW
wOrPy7QI0h3jUacqCS7BPxJUqKsCt65AVsNeRYpG3qqiDOnLPYRhAjE0lL/CP5HH
KPMjDI4Gjbd/yesIEs3g+xH2QE1NLvccEeC7RIdPt2nC4yx1EV3iagMOTjRa49OT
Ocm7f72nXKsbkP3m99o0SKOx8t5XL0rjGSLUdE4vNFS/5wGkBQr4MVX2eaFHVzjc
GfkyxwDPdC5IcTADYKqRkjVREpzzixKX1Th/UXk1NNU08FTo3iuXP1whRwruwkfE
dKJwtzdgiGPlqlxC9kgUtib6E2oJCu/0Qy05sSYtDA+HWj/7nbtrr+nEbz0E+a1i
IfTiTA0zZ+aXU/u5SmeVrjpLJ6cVUDHclxEFeMODMdZi/2F8IMj6oxndZA/dkLKw
WD24ZhVC8CmS9bIDJYml/Wmlw+lkjy4AhHIPFpzM0+X3VPnSN1Ff5upmmbDmJLq6
vFNRxjlgyls1n44zjauyTYgGr3tprhCFefyePcfElfiUta1GdLyXCcbRz6O+pLWA
4Su4pTQu0Ju7MvvbMJ1ju0fBq9/2bji+nnfV4l6cONxT2VUJGKUTbnMMxrKvC2yH
v25qEBSYnCai+vp2scNCd1+20pllz164AiurjwzoTSj4mMk441E+ZSKIdJK0mEP3
ddDzNzaEQ8x7GG0EBr0E8mXKqdA1aa+wgOWdzt7xpke4u50fQB0V0LTGy3lhqpeK
1nk6Lt8LkFmyYGC2Aa/QOSpaXr9u2p+XEIgkJQ7XAR5IKqyx7lVOGQy+lFw+A+31
mNzPEF/bSwfVnUATxufivBHA2tj+sALngWMzd8XAj/y2FbkExmcanwyoqNZvXScl
vJPelkZsSXl+xl+v1iV3bV+v5rCamZBvKk3YEbi1aoNsLXAtt3efQD6aRvjGu+wy
7GglD9PVBodxRR++vwf4NxH3k7yPZeegC7Ibdm2YsGpwU9nk8lKAe5zRu30/WA1s
psBM4vUv5AUQ2dk2AQBvdAyLGOHPOui9fJeSd3iMUPB58966j1TaM+wul5K8b4IW
u1rzwPWe0VE/Mfpgj8h+XsTtH4bsnjxCnZ939AlgM5E6gpSqrkK7mnpliACAVUGb
JqLkZ86z9GWr7srxYJG0oVZb0PBffbXIPwK0QB8phyE+0/ApoTzeiSDVh3SV7NGM
CBsAvrf+yOYjK3DIfCOR7C9oqWgz/L0GGPp+9Dr+wf7sOez0pvxh0nwGgRF2KQLd
CINLzNPNJlA7Nj1DzUHibdPXtXweT+4NtvgfF3mqTdhCFxM9LqkChHVhnel5LZ+L
esZfyGT+LZCp6GIeiWLMLmx131bcWePverBiFouJw0CHl8JlUmb4nOldAcVEC+D6
DqI72k7TbpiJROimkkaskDtY65adbgeGKTVSTumn/ABpYIvPzXEwB+FjFQ12UdNs
sfIZYSq6q4TldM7FLTwBJ5xITQDe3w4M6i1LAnay741/S1OHXn9oUhH8Ba/zhJZW
wBqzcP7s7cE2POSy/EZLaAqCYLPJKCEB0WbCwHTpnYEdys1VPPhLb+HwOcSa+/MB
RkUe7GObBuOGfg+2kQUyqKjFOqXYtaj9vyMjb6e/p8vm68jhmEaDtCW02WKCxMNN
vmW6yQ6zBcGxso/Wa/zVfiP3KhKswC0nb5SroRmhujM1B4RI+gCSDfOHfz/uRDmx
YCDShka1QFeLueIk0xZRt4iyjD+PEgCU6Wa5nsUNJ+cyLVbXVvCSmLtoEskI2hQ7
6f6ebIfPTFpKxb3Utc9SdJasMFCYRJ+bQQn+MYw9HQYJ5QLk96sQdEl0+oIIGePM
e306rpudspUfJ0e+nuHfTpDeWj5ctC1bSVQgkdGSTkgApxzNewo8GpbxL/nBa2xD
0grcNw/bPuXtuZWRhtUysyh5pCLFvir7EKEH0p0G6HuspfRK346dHB4Fda2NJUg+
ojihi7WozgG50B3ZIJ51Y0UUgyYsNXZpwPjsrufCb3OaU/yNr1+QQxinNnvw45cQ
FwC3kpkUhVlcGN0UsQBkK/IfF8VralvC9KaBkGM5M6asUbHyExkay+tMMut3MLe5
sBKsU+2Dw+mpJPfM7F134FsYv69ZEZf8pOcgdGGrSIL0F1EYtd6h3DsSZDhyeiOr
Y2clmxKD1oddXeLGfMf7eYObcWXQmAaA0EYAMTmXozMu/3814gfrtqDPPZWv1EN5
CvDREUX/fv9KWaNgGuxgUKTw75lkVozBcg6dSz5zK9wgsGB3VjcX2BXPa1xXCosy
hH00nYLKK+ULLfx05IIkosKkCD1qGZTSN/ueApe5OjxyoYJfUbgCEFnwslnlTtLZ
gEifWAQXuAW/YZIJxvIjVB4mnyNuo0JAPipClnZsQOCLgnIUGVYE3NYUw4O6H4vv
y6Ysblx/gfLfiQUl9Foq8jcsdBeeUOi+ZYB1mEw/LzIazbUJGOmbLH4AbjSTzvt8
W3e1Cx2rv2tnR8q1IYOo9jWHzih3Y4Q/VpDEyh336UD7q2ZStl2NGL83szr8s6Vl
W5MSU0ebecvNSZDXYXEIEafBws9K7+veMarMS/Z+S+7FE1g/dr0XHHHuefYtZUtD
Fvl/8hplAFPU42h6Dy4ofqE6WPk1uM2QIrEONsF6JPZRYtdlL9SczgraSrL4Kojv
BO7b8498pCz9p1VmhsH1MvqrTmQvQKBeTQn3GqPJ4RdUKJFO0ls2AOE8tow1q68Z
C0AAkUbVzD2BRlr/gXdEPYqZxQ4TwEfdAv+8bPzGT6t+HnlNmupz+Cn12iOrmD6n
ZbjwxoaDb6nZTkR7hXQr0ce0/dyLczClme9hA1P7w1zYK7zRjJ9D2MCeNUNLym4d
zejDC7peAm8DfqhK36Dd6eJtfnwbiqccedFrHRRcZ83F/8Kl8Rd+YVphK6R2E2rt
pylaYdoWyiLVVF750qFJ7nbBeWxEfj9ztPAx5zFbwsf4ryrN2I5x6RwPD7lO4HoR
NdJ6C7qTlT8DIIGYY9BQGFj/mxKfKyDWy5CvnKjV68isugvlGZkRC9hUyuKDA+/Y
yI7Yin4GE/KaxkeD4YYlCyhnBvcUxpTgxqlSEnOjo0lgXnuUOGvw9amkyDGOTGos
yg/XxGIrZpWcXn/PPPnL9YmmAc7b+5/PXho16Dh/Fy+k8+C1XGo9TpnX9kOOXsC2
j82UrkNd8BCZPpS+eM41V+QNsRFhWi8yoSB/EWkrnOlxJ33Y9b12IyPwvxae3Oe4
2EZaFWJAUamT2ug8b2sA2RtWPxlLq3PJZLxNSNDAcuyUBYvgpuQUPjiFjNqpm+a2
8E/TX0xQK57Ik+yMpkxfdI2Kv6FSWUDCbpJl42pQcV/n+hLNA4Xl4NMtHLf5eHzx
rCt1WrdfdT1i9xDSzb4cpVdZ7OyQUiaJlm5t6c0vMxyNxYw6hANNSN9v/fvecUdg
HYZpFLZmAVGjObkd8vHd8h7lW4kU24EhYz2VBqsVmYkOTn6A875wOQng2dQ1GV4l
vCizAONewmy4zal6uMzihCFoF7kXVWXk8cKojYVPbXaZ5hV+1jUOF/iuHBPQy5eF
fV+lf5p0scyhmJ86kB4WrUTK+iO7b1CIMiDZAcVd8t4952nv2hXxDexLqzer+zVc
NgIhpfK1/0If6dz6zILZUNjAnWVUgMvSqE4uNqXWY1eMI6yNwMATWYI7JQOsDTWx
bBpH/jeZ18EVLqEJal5ppuol2VzmQw3IcIwSgShO2ayFB1pTQvwN9kadwxWVyyji
7F1+NhsM6NX8jK1wR+694FOdzMOGI8+6goO8ERhcLv69E/hMjtyf0Ikrt4Zc90oe
myvonSYkEjyeJUBaRSLBeF8irzD56axJdRzfzH94oFA/zYg74Ypl41WJ6h3P0XHW
CNPX1JG+dnu8HP+AcdNq/AOjSVOjA+WxuhH51ZwDKZU9LX0UVskVmV3uXBn+bVIh
GORY4icdWiCb/xq/VIALMY3N/m/+WpPdwYQ54cOwmsBeoVn8d/CqxByjhKoz5UL7
NDXGDIABSWqLVOGpZFuj+nNVOFNQtlFmeHzWFX/bpZBZNXyMAipKOYVoW+G6NpU9
O7KgcuVJeFQK3RW5XaF6v2mWRmb4ihsfuGms/KiaXODuL+vUPYzj2wShPJITgDKX
+it44ww/aa7/obWC1oh+8rJSgXNFQbh/3IayzyFAumrOehaFFUH7UV8j6dLmWXGw
aZTpqr4zPmPgsOPaudYs86Cx2xLe0V6oFqSFAAr/1cXfe7tiLSMAjvrJkJerABTt
dUmnPXQLGQsltIV8IgsXAFWJ6ddtXHLJjFXyaJUwpgRV9ZJyZXNIl/y8ajZ4x2Ye
s1HeUnLT9MP55ZALENjmEMUzGFJBeHUUFweQtGIjlu8XJr4GUPQ2h3UBJm1nWchQ
ZI7qd4Z8fE8lHziJ7at5OezOa8QljwjhyDcfoSOpgKz2kbcV8NMohUKUL1/JbsdT
W4csvf3xjLvzJ0AV6i1l0cGelokaprZ89w7NI/uj8/MpAzBby3wOzn0lAnQ1sQxK
pByxQiE5emqx8m69Vozemme0qdbnvAo3o+v6rvkmeVEfHwYtGxC0SlrwgUbPjrns
AoUqstLAAAfl8EleGkPQczxN0Ctq5e9SIXWO+uMzyOmUj8z1NIIgGMm3nYKuNuEG
B/JqyadhojYCgGs/H/GJOqQBzWOYqbselUYMV2N2jCBAUvc+bbpPUdP6xSbu7X1j
3fmjgy2rF9jEPLCfCB2S6xs1fDmnHe6aNf2Kif1wm+jVau3e12yM4LPNWgJyR1Ok
fOgvkOZ+BGGjeRVuCbdvxw0YHyl6ZgC84ORhKFXx5WmwmcRvRtOEjjM7jj7PnQCY
KP+KE6xkMYxBrd5P+yfucfbqo3l9PsRi/QAwYNf4p0I8Wf5URoAv3P7bVZ9xxWIb
+Mo6meA/LZW73TzJgFcstRSYgIPsFCoYOAuZplP7HNmLvPXXdSTTdia/LGtR9pZ5
6tH7vcgGN0HnXSa+DfDkcDLTVLZWUrjSv4pOOFGI+vsM+SKIhEErpr0h7dVBG6Dq
Y9/oC2ersdZJhEAuPIbJaF7ew3lM39CaZtmEz/7t/jzOb/BTBNM/vP6FVkKmb9uW
iLb1PUgtp726mrB8OVQ0pCmDyetaYPie45X+pZfRmMjQ1sc5Mr1RaDf8wsgaY1Cs
3Fjd//Je+oGMKCEEyQXTgumARmTFzCXObaKdb/62sH/ZLMNxTTgIlUtrLLruuJpw
6AysJmbLeoK4m6iYroAhpnovfean/StVklpimrOpY196lkUezqpe+1TnMo8Kw69y
UZrbM5xdynOfdTl4kGKBO9ZTUslM2EZLe6PiDSv696Nb8xjzCSOhPmQpznE7ffZa
x/ZIXSmqEtfIRTBSOJjN/NDfr4FGnfgHQZPLxGrzjEXyIgj8WIToNYIAGnNA7IH2
B8OQQV/p8zJbEwjs2Z5Zm6oydA4ahpyBPDAGas91B3IcnOq7t5YwVrYuycDzYMnV
SwEA8Rk7RRkrSeVjowyajMa6LEm+1BS2nK9503wHE0DyzMY/ceSBSod+vV6BIngU
gUvBuqWMQ4Nd2GigCqm7lAeVKXNzgxEIjs/jE2Uu19VZ9FTOkPwP7uq720jXA3fc
udSC+Mn1MhXPLVfeSy+eQPOaIc6ByOKL40jKQQvgm25fJv//ZNUnbAjZNB18MYR+
cbJf66olBJHZpypqxA7n7lYy9iQU/apmfMbW2DwxN0NswaIbe1q/mpVn1T4VQPEx
4nrt1GZXF+nenKhUEuBJYLpWBchhZNTvMeOmPuSG/V/ZYNSulMwYacC0qu6LpQdK
ji0is3XIrLyaXEp7/Wl8nfiHD9TxR4IkpMknYiJYHHALtMtWuDWlwL6isBKymsgi
6DHH66IFQZ/sCSzDDEeQQ2lmX33g9NCVcB3xUFjAybZNALcGerxzVR4P+sdfIJ0l
AoqAhSlj9ccm8VBizWdYDSBovTQnwrxw1RSXwdkY2inLZirFUQkDIf8IWzcwU/UG
8S+a88lgqvhiLuzH0i00ikES/Ju6O9If34fy3NoQLw9+pM2QXguIqqNM18FixM+D
2XglBzMn0dq9IiXkeW07IjSRBuCXcOiEBEOsms2B+RWmoT/cb1anBHedhsDrcB5b
h2wRQFlx5rPoijCwN76MpUd3pF4HOolcSp3w0MPzEFC1HEoxwC8ZNEkD8EThLjX2
iVcEh4sf8BJy1gAR4BXyCmAZD1/exazzAxaXd5ecGZn+I99V1PQQ1jWSbU/i5hwU
JEkFwshE0M+42wf4swO+GbHEmolcTcwsA+968FsoDWOj7oX1JPYC8faMRtB41kWm
w8xxUn5Qs/W5R7gD+L0prByMS3f2UIWax7ZJkV6PgAJ9QVKQkX45Edvb4SrElsAl
cEnEjVV7n7KSWipAjwTDMvCgkJ1W9gZEFXblJMp2TB4VCK5xXvVOyXMJl3X3r/UZ
l/X4VZhZ+SQHtU5u+HE07e8xo3F1bGCc0JPUXsz16kd3EpWI8Aprw6RFSqo4kqRg
z9Ytxk7AoLkHcleHs3KLUymJkgEEdNd/MPIhNAV6ElEYJU/xvr3B+x/xvdYLyI0y
Uk/Kxck3TtDPZAikt464LfbJOQrn0dA0Gw7/oswmjfzeL0C9AwtCvGp2hZmSUhKp
uVnqrkCfkVasbeG1V4W/W8r+Y9ASJbfb84oxvWhJPeFaexj4ZAamYL06Ij1Dbvy1
e0Iy3X2n/kVGSabZEOoRiICHkLCzmlhQ3pn8tr/7PxORp0QDVRoCjonlei6L8FeG
2IrUuQh4GwDW68O3pFtFgpQ46HtcMp2wUVRxAvRFfXEl2sTmMNUXS3HPL1pMgrbE
5N+hFd3MvVsiF62Z07FJno6RB0OSKnnGNKmOJ1X1YFvcKIuT/lItb6jJhN2pGJov
4s8IOEQF0SU/jOWUtsnSDkemoEl2zW0ljKTg3r8LF+Wu2G2K/vqVaha9AyMkLity
WeDOnG7dXqr38ytFiS0GyciwvSkDKXf5IXE+pEqmBojD1PjyknonIjVueMFb/lyi
Ki/bJ1ABlNmkfxmrUAgahPXi3HU8FZttNVFPXn0RkrY9FKi+6JV9AZUhMI5xuFeZ
l4meFhDb7Zi2SEoKxMMAey1GSzvHVDlDtvO4+QAP+BkX1EFh3nFTrVKulUQrHuaG
orhD6epLtmULz4yAE3iX6wlOsbyebJtV4Y2fQuAzHLUhOveuZOKMeDRQnBGoG/0l
AreQpTzjphDrwML+0lYJ8x8DwpdftwaRv8rnA+nn9vYq180XGM78p4Eu0tSQ3wGf
6hrPPXKS7RCQVFR7NrJCMi+ayQEYqFZKwt3wQvw+FcpxZRInVZQXNG89TGMCLTN6
c1XM3iTnJOqdWzHtsexZ3Ls0Bl3g7pdUFRmR8DM6IH7RVYnz6fkEvb7KFqbtKtsK
IMfjdkr/jBP84yFVtjz1LbAgkPTmjtVM3tRE4OsV2mhBp5/FIbj57EJDRCLfWIR0
hb4LLphIIeFQeldvfJ5Hcfy4dnPHwccwnMzNWlGf1N3i1rHaWaOBVeyFdKbHwXfn
5jq5Ut1WbZe1/W98Ingonzm2casRBowUYaKej+6iz5Hnsxt4aWrSa+M4YXboWiGN
qlGCFBhb4Z8alWbpR3IGygXeJeFgaLLiOOj6V1RH5hqjSTUddRXhvDrgcKZO5lkU
NNzDnRNbyb97wCfF1AdIVkksNrInSIP6d2h8sJpIkf5JF1nYZaDw1BiVcShsCf/R
TqMi1dbnRL6NDUedvNK9dCt3BgRUcfuhHnxuybTj0pRdFomsw79cXgDvFeQo+EuC
oueFNBsARHs/IOl/fbZZ5SEuIr8n3Dtsos9plplvYHEptMLuoP/qphI3gcFr4320
U11wQmXybfmasKXMfHM4TsLS/e7jxriOTC1Ooyj33hOTI+RtsoKEdy+2YTIzs4tB
ku1Rzt0ZDfMU3OCRz/irlos2sVvvp6Qwj2AAlk9qz5D5V3/xKWDkKBS0Cdc0BiF4
Ufn7BGZJwh46AveW4jxZXxh0vyM30GoU0CGNKcVNgv5m3qVy+PwYSrkLAEyqPulq
JImW6v3z/sLEwxk5WiWp9E+vpOzXvS8RoGFldjDYPyCNBYPmEEuBvPAExH156COm
Cm1dDLMg0q/lPUrIbVTk4stfPpzugwhsg4CLBarllZXdsThHTFrvdJ3FvbvpS1t+
bz+QfNxCFqBWO+fCOm/VVIo6hffG6SmlYt7f1gJDOGmQA6LGi/6fQem/mnZ2vDnI
FNB1VrtbEjGtwhYBhfOGt+uXkkg3DlYGAynomekM8sSA8lnJOxLXb0Bw3zNOjVMC
kIe18KVGc8R2lgtH/We3Y0V4UhoawokQf8lCQGSK8p0NKkxSI8ghWoSFzWZNcPKo
WcQVb9E+yc5+mJDj8iG44oLsQQPvrZaN6G9GlVSozq0vSZc04/j1S41rgfAO3Vme
sVZEZ0JMX84W4Dvcb4wG91JrhJuhmb55uaZOf8N1DxWMRkYvjS6GII+M9l1gLdvo
ZRUuOLjrC62WV5MlFP97Zv/xPv1eAleHGZL9Y/fx3DtUDZUVIzByZdTyqtcyS5wi
IFK0kxTwes2kAe8LYukpQitXp0AtBmK4n+54XOBdDi9IlWxWVQRVf5Kvuta5Wnu1
yUUGerP4jBxN6O4+eU6oKxtpP4tCyLi+aHzLAJCe1q+eZyVsVODfd+5lbCLh7176
il3vRX/tHWnjC/LeklAJHLvXA9HVolcPGN1e83e9hll3owrVM6empN9ClQzNGdMJ
P63PELa+G9EkHDT5ZJOskq0xlEOf7+sPHl2ekVuuhDZ8JxvvrjljAfus6AjVJfiF
d1uwBnLqGLqQFO5fJ+k2rfccykfxH613e2z6q6WExImUyvTWtijaP58/L5S0ebX5
RtGDPaOS/9xS4Y9pLrelIkCnts3AodUGNE8NFRQIoZNBC3OYFm7w4Tuehbo1NW/R
18qPpZlSoksk/IawBb3M+iIUPKyEEYK63GExoE1Ak8mrgvRl7i7dPWd2cczyVxQh
Afcf7GYIoDWtyFTy/k+YqGagMEJf34tkEmDR0KloB6jkL9+fGcegEjOzle4G50Wf
R6Z+2jvgwdlR+/sR+dOZhwKXZ08RtgCjAIibI/TBK0jaTRf+FmjieppvTlRVKYgM
FOIZRcAwVvkP3C7TVB4mwhavDIuPTTJwAXs9zJgVbY6RkwVxvBP0fX5ue+ZxjMnc
m0QVXTwgmKHLVUOblRJ5rIFQP1OQBA9FDwP42Rd/9SaD88yujGW3kn6SnG/wCthp
Uq2nRyoGezaNeJABKCMxbI51QVxODt1Edb/IMEzCp235CpKI1XiBsD/ONFog9p4k
wnII8Xl1Pwx6k6/yR+JLoH4FH9ilZ9JuAskS1SVN2Z2eZG8yuposCTYV+M6RQugU
Qz0Y11k2bKhyHcbL4RGr8uLLeKNS9cCR7rVb2GwE2vUoq3QoebUA0yqp4bjYhwki
yrn61rjH7Z4aFa/3KMx96zFwp6Ir4VW31hFqc7YHadhtiL/14sFPnnk7ls/kHN9d
fCLv64xOLHJzAvsH1yljgA+GBxsgmRX7YSj9mUUFClu52DQIRr1D+61j5IluBMrH
ZkYRWfNjO7PYrcqvJzSbPLRpascE8zpDxIQT7pr6auu5ORfM8+E3sZtkZ29HjkJ+
8oArDLFwNKO7z/7mxN0CLRjKdZFUMup1P/+KiqDQZXasrDTF6jKrSWhz+g22Qc8J
PuvY5HvQ6mLCRVIbpboCtnOBRNLEVI2HkD7X1zLr2WYA7lSWP9c8XSQrr5ExC5MZ
LWnHpShOIAiSspKeyE2lWfE1KfHXftLynRmGbREtD8ttkMAqf/KtdzTl1dOf9RpL
jRbq7WohV8oe2f1+LpWKo39ApkMKhzBXk9lbZC8W73eLjkdu7ccVVCdqa//E+Hw3
71WkFOC+gp+g9Q+wvP04sJ1pqNIqqZF2ZYumO2ScZYlEVCGk1EY1c5Juxc5CfDKv
XwlCyd/1zo0SMghvPVRDOCNnzjtnHvyoWtDnJalBp5leOY2CcJsSjduES/t8Kdv0
uH+YHrJjmPf2o9N5DfrwbFwgyxmAeZlR1C2zxiJ8aJz7E2tDGer8mknyS3RqOs2m
zRkZ8gzctjRU3JVR3CqeEvWNU3bckmMuoP8P4PSR1ZMcyNLzGVizN1DzMi2phNHF
ZJelom+8ghXofPBKIQdJXYbCUXESUQsmClXEf/B/KZBmRIOGRluA7II4sPjLZR+A
aeIkraYaMCok5PsdBVTsYWnPLv4mMEiU/8M0RTe8gmpkGvyEagIs0p6x77mGuKTj
PJJ94ov89cNT7Uoi+EEuZ4F8xNHVUzD49zRwTIkCxFYALRfMRsiFr1QyuJUi4q3X
zVDA5AQwCbY1d3wDeMi4DMN50QpguAAoAycymwN18Ka33H6sOAdzzneYNHxvW4Kb
4YH4lAU6DAKFPidqb3HXMtL4T+F/DkZqZBnOz8gV2wUHHloyCkd2yQujR6p9J/Fo
TkxzASdQE9GbPrxR+4MZ5TsfIuPDJJneSRf7RCmbedRGge8PhBUKEFCb/yAMqY6z
eaxFmlrfWys+njaoiC1En95S0rai2rNe/o5imO0zVTdXG5mfvozDjxcWvtfM21se
JBbpK72v35jF/RS05G2QGuh0jLFJ9cgHMUa9bAPM+YoCpRdPjI0osAHVJpqoBS06
jrR9NJFMCkLCnyj5PAQNgJ9yJolnD4SEAm7NEMGf7pHrShDW5N4jurDr8NG9prJh
DImjtfOZETJFJWC64fNRTkBa/jexMJifM1fMKCVkKmHnEaoofXRM76fdpkp50oi5
LzDiF7IXF9GXBVrq9RkVrmdVetYpITChjxQPd2fEPS8BREW5GWxWb0CHQdA6pmW3
pR1buAE09n+7UtKRuEtlJfWbuQSATShHx0LmlldeFe7+o3Gl9OY/Ne75EnL2AK13
LxSkWmGhnJmO7uA8C6P3zj9ixoTz5haYBqMnnXVyYJUHmXljVU+QBI7lxRs0O3G7
nNXWdyYyH2UA1GubhIGsRbnYBFjefDqvhfa4FANGl4u5ju4u5ZWBnbyyq6npVTfe
8LYsawuaDpj0rjIltv1mdSrgeJoWRrvTyT+12FPnxAHJtyYjzg1dBdHztZmIx5mn
y2UWJfgw1dyDjlg4iVCUsWeafNEGk9wDK/8Sr6VGtPjJwfdxo0WZ8VhTgb1J6546
9p5pOWaLEstWElOTrIEBJh9OblCBl/ByOJ7Pa6FOA12nIG++94GLl0NqrnaLmWpR
EqNH+x2+z8D7Ulv/xXH4B0e28IhQRShuGwNNazL9VrXWPEdXzDYY33vFIeTPbm8M
O5cC6flqWHHJVipf9fBHwI9rS+sXPzrWm0vWBvdGEIbYBwia0APOQDGFoqf31zWB
nsSiK6KMB2tS967O/tQ4Wt3333J163mpiud3/c0FSZe1MDvPg/d3/KC6VVUzqVVL
9hsKCqCa1eqADIoqbrp8ogqgC+CwMIaTFJxIgTayHEr2FnmUanNp4pu6Fz/bEqkd
HqLyhqHwOZANhRAUXm/ez+7CCXS8J7bpPJBEAnd6rZ34x6bTCzgIpLGdk/6OpiH2
81gAER0vMEQVeKaUX4ZCTVFpPXaI4VXe9je5iYHvu6TCYQqJa24FPfIAePEZFjtc
eQnNeq94UPuy6XxuVKTGyCdRaYo8TorFbMQcrZ2AX7LozH6DAu7FS6u9CVt+H4gk
UtWxOdvSFT8rW+0LG5PlWVvou0zHVvdJbETbd9BDz+dX+Ixe+KjPEVNjdzWsphsI
CmqIAwis1BHtN0LjA8MHk/poza0vC4aj96gakVoophTQL/u9frcMtPctSvY2Mawc
8MjQUGjoUk62daDglYxSLOFFDlSIY+vV7ngMdJqcyIxOaJsDCeO+m3+MMkxuy4c/
ephKu4ku1Z5L6QKbKlqALGhsIAVrdcpyGC9d9rk5CBm1c+zKSc/3qafss6EAl+Jl
UtLRtSUFuCOVoMqfgEqDmiO8hLMODYIDISh3iakoskcRKXEAw32Ch1dLpZvc+y3j
V72EDFdFUbIZoUn6gkzJHTXJFJgX8tk6hV8lO/nPVBoY6+f6loP44VcqiqbVaBmy
v61c2rZIdlBmwVgUsSPICpHqe2DBi0epbJvuOaasi5W4mQGmN1sF2UxynYEFOpRw
nVs4j1Vns0tL14NKZZ9pSntUkkM+3zi2xcmlqKQLv5z+KdVuOQvnqbhyG1GYjcnd
Q0bOSDxRFlK1vHbo5TJArZPpBxKoYNiVi2Hx+fCssjWZMpVLGQKycQVZoKqoANwl
7NJLw6VLyZVPkweehkK6U648TeFzONVSuAuUKxg7DXTc04uvuGQb0DWOB3WNjoFt
BkzlkWLJaqmGQboKqdxOS5dHHhtC2lT8046AmIO7ehRRbYZeij54vo2/+H9flaQ7
LEZHPk4P4ugle8FqDgmah5gtKaxr/S0JCEqvbkASk5YeX46m8iSB/EGChrzAIvRI
bLmyAOXCCZM9vxrqpqiph3KH9soLKEPHDBRXAb7W0E1SpjWkzR3G3jnI85I/OU7g
IBVmGTIqZq1wzLoic+HxrEfcde52o0uivqUdbCr8DhhtLDs2m+k+fwiiTdBJ8utn
NbYi8qIOrA996vtHHKx2HVZp409NV6BoI4d6r5Nw7XbTTUpLHpF3BAdB6V7f3Xb0
Yg0fVa77i29pap2a8p0lWrVpHGs2OGqX12opITUA7pEmJSPqiHWExh1g6CSHL8kq
sEmG8V18KXfyUqeMz8f4NStBr/rR6Php39pU1nf7hyCCo9aFDPdybOX5ZaiuDvxM
odi2Ualv6lwiQQQ7ofxL3+FmXYDX3VvAZDDibW/F1WbCttURDuThRQoCtlvbPz6C
TJYi55KNXaVJC781iPEVvycntSpqXidPyoCy5ZqYp94VGXrm6b5t/8XUQEKp4sFI
GqpVmHo24TV65/4nYQL0vowC6Z8aWQN7yv74+5LZcMqVwnF4QSDJQN5joZcqEXD0
U9F3WP2iZideqihCt7K6KjOUjEu10XZmV4LpQGbU6lO18q/nDUjVK++tdfYjL9ja
1CvfQaHuSCMpSLGCm+UGu3uXqKeuZGKS8Z3ziUQQfeBjS6hilZkz//5NvdEb1kKM
DadswufQIHVsQmtuTbzdoX6HXDF5cw97Psgv8n0oc5vYH+lwLBVzD8ybuz4RLrLO
7E/MqLdbZHyNFyC7UGgsH/jiUKSmCGXH8L/OHkN96N3T+VJNWWVjTo4NCzSutZuK
BfMuIMSFLzHalPT+vJMaVKvzDrxWxMA6L+T6zxjpQwm2XBWAvGIr7u5lhag8JpW3
6MZbH+LrC5gFC8JvHN7zzL0vEtFuRSsS1qREM77mv+6keBJXu17V7Iv4LMpClapm
O1HM+g+i8pCKmPsBEbQnWXdaETJSLWx/nSpIH8PGMzv5pjiC8HC0vkw1TpS+Ewc+
0HUOUdAXzM3zEBdR9gG0ZkVuRMO1PqcmQ0H1XQjhoe3LKZM218aFyW5v+QK4Klzj
mwapmBSkpe4MlPwPbOwVq0vxwyU5atxWM5jqXzY9AZom/MT9CNV5z8+iF1O57Fo/
Bf+4Fns4Pa4Uq0zRBWoTonZPE469MqVBM/6XHTm8ESRe/x5hnn6Yh9xULdlA5uo3
RPP9EqCyveu/yec1KP98WJchyOUEn5dGIujOcwqiW7FM4V224KaYHc13nA0Z+Qwu
IZlQN35fKPi6dF2BtfI30+kg4vUwtP7C1u8JqPHPSskUMstT3VCaVwTM0tg+viBd
5tqlIcK6FUqWZVLBwIjtyxjEqmuapPeX4QyfmYo7hkt0fg9dAlZZVb9g5aGlvXUH
3vhGlth9RAncjVWPiTUPIcxbVM584JW/HsdSE3D/9D0iLfj6I33w1RH5evuIvai7
hxOr62yAAbmhmVapbTZmiclL03f0717dmt6G4nSiRrDAqu45VsfqJn75aBSL5ly9
/SMjsIhGQ1B0NRp8qE70bAb+f9Ttu3DrFBwSvPILSaBTWmZd6HnIU/LZPJB/NRpJ
zZ9cWgQvcTqsZ+IsGJt2yIyQC44OlZ1nzm6vJpV0ZSZ8KLjQ8RUWFen1ShRaI4oW
rC0vL+RQS/dL12u92MIr6XpmH5PmGtUNa5wlD95/3+c+dMF1ObW7UuB3y7MSHGZo
UnGHMRZRlX6sISTtURcgS+QkZrfSHGx6igqJ73f5J11EGkP9jhgv5bOa0WtBOF3V
3y5O6/wag75xK9UH7X4p04GY99HkV/BvrecTnCKDfrJ+2lCwIdMfc28tA6g1q+YP
vacciCEsQI5b0KEdc8EngyPdsQvzRmNinXYM1sH3xTNGtFkHvTLlo2+DCC7kOoB9
gbd1DSUNqoSQNr76kD75xzosTbMWR9NbCrW7cuXA/Yq2pIlfvo5E18v65g8WRTbx
2vAQ/5hpyh2JmebeqeFcY3cjaVuVksWOaXRDlP3l9QqdY9JrJRCsjSKEqlrQFI+6
Lg9pXnEXt/3TwU0kTWH3sq5Oypnk8wPLGm7MdYqDdJgRbzPqYaKitOsR8sWnGOye
xv3PdG8u2RJdTzNj0HZhCEzF1/MA/70paOZIxK5ZvmpdPa05a4+XlepfciPxqjbz
dp7l8miNhfmtIB8KoUnZFSzJPk683vQi7yfpc9OEgL1KxMMyqv9gwykwRw5hXrKS
EKqUgeNZyGyNX5iQn+c3MwWy3efA1pAUiTWMsCv+1nCskJZOG7ZuixycniZYEV66
STVGmTreVmNE3MtEQZYKoyGrOrvcR5/cPBvkiUWbWAh8HINnyM+tDkCY9kyYYEJy
6RXmjX/jEQZqxLFdqsU9JWHTDOFx9U3DGJVMTEl/uaITj+ICZeFMmyOI2yFhPi1w
J6aQrL2reeloqBnwypWOZnbtYX5/h4U40+QUPkInk/8FqGRJy78aSDm4tJjBlIn1
1Fp0jWw3MaVi5XQNq0RdFpqHBN80frZ+lrFDlp+up5DXfU3HHvoyGEGut29GWR2X
SQSI6qA4dwjnIVeW2p8fFiNcUflqW7fiSj2vimmIZRikYeupb25h5kpMSdjM3Jfy
RjUh2QHb2VQsZeJF/tebYnJ1m7QiwychGXkH2cFaKmxDdHD3cu3syI54bLw9DMPW
8FU2ueLLkcd0TSIZ7T8Z37GdyGmkXPFfHgYhlvSoK/Cc6xGv/lEyK90yX+S5EcSY
rMHlsg/JcUM7oei0/LZACEzc9/bkVYAZ5Uit7wfkVZOL7g2tfFcqGDNmntPAu2i2
aaUGVNenTWug228dufWP52CKL0c5JPdifOWnpOS+a7AoeCKrVDF7SQw5EndEtJ2w
fa6FQ1QSpzy18f8WfZ2BJcWJIdydFErV3O8/O1eSRfJOYpExoynqE/mvSfyg6ywJ
9091arZGIsgz39/xIsKk15Qo2lwnilJpnQvs+ltxayH6UGmmji1uMfTlfSctEK3u
Rk7MxRRpO+AF9m452ro957H1hpmFBOuoPropSuX4+erdemBJquC78Qs5vQEdeqHw
qsYZIvR+UiY45NWuzQLBCrleqEDjq3UmRUXR8Os3gUheQvigd9ldeI0txV8kTwas
pt8U4QwmcLD+5jz+Tj3PCU9On8OrxnCN+7MpuFyDcEr6mPVc9oPbMO3J4Qlr2Hr0
fCL3bBflch3fNUu3ZqGpBM8RmnsRBw2KB2weqYUZh0kasi+zcHQ40yEOujJ0LrwP
vwHY7Ukc0WwrAHGmyTibnoYQcPKhQb38q7PmuMHD6WlTpVWotyZQe04hlbZlvhk+
vO5ljOemTvkRLdFrgyr8oKqCfLlwdeIzHsfq4J0gAIDs8Zn74QFc72XjE6mkgP3P
xyfdixnCCyo9v726gIVlLJRRKOn5mQfHGvRWOrzFMD03dqNMzDqAB55QxjblXaDG
bJX0c4eKywnBSAOxp2YDZM1ScQf2zeVMnrK8DhckWpYoX/bJn5UJpL8HPXA3xsx+
sHRq/NhSoTmYNAfuN06ljnqV0C6J5ljyTHD4GLCzhoSjLnqTwFzRCYXSC6UTA0gA
Koknk2kEWQsM55XR+oAlkOPDG2tJKC7u+Jfld1xQ9XsK9e+opvwgwyeCB41DuTjQ
4CgB2i53l9AaEcDzSQHMZVRzaGBZ2ExyvRokmSriNKSKfhOiISZ5BjDLz3oTbXmo
hd83Abp9ufNMaOeuh/HDSUwa6YE1na3rhwZdhv8a2NZndVFEviPCUJMFdI4IC53u
0sEHTtQ86dLto9oyCN5J6I/iZxj5lQvVx0Ej1Im06JochqGNB20bE/bYpZp+rMKp
sck7JVwn9ttO5TA+Uva4H/ZSMydkaiD16396TI9PjcoIqjd9a+C8rx2yYDjmd+od
oGjZ3kid+7OD0CnW7G6eDED8PkKKw9bB0cbiaskyE9G00L0av3VLTCzSXOy2tQTg
xl8XaAlP68B5RXPhdFU6RWgrFZ/oewX3k2etmP5lK5QA67AisiEPR3EZFgqkkHy2
ylsVtfNB+WMi0cYpIII229Qn/7GjJ5cRu+JUsQ78mVMKdC8R6MKSV9DqUuepz4Wg
B9KlXcbxvaacFjNzIaZC0M6cKf+VGKlO0zsZY1ikX6auDxsAd1iWuS7MY7FA42/T
+Syc+Phsf/e3AAiFcfSwAptFVMqsjdxxYXzOh5ifFEx0I3wCUDOtSnvAbpUO4DtO
lnegMzXBQ88YcOzyRKYzNx6N4UJW0l90meUOIAEEh5auCnUFWRnJHoHOVDnynbjF
Jq0vUNHEi7TmFkagWSo5vthCGDkHjMHKZBC16K3l7hlg+S40RdmvKj473eEZdkQj
5W33uX8x2zP4QmBhLOAppAfidODhrJ+fVAGcQdFWecOjczs1zooHciOkbfWCY0Ce
4i9TIJQGakdB2S8GpFPz7cIFo/hzGrfurErPC8akoRDltGRAdKTcctqlbR29EiE/
hwhUKoCWNPkTUJFginWcWoI54AQSsUNuImabIwqBeuMXDjNp2/4eCdwIIGyK8cfO
ioZ+wdv5E+LjwqyJV3aWjEqigqtMttz/7IIlen1Kwt1FAt/PNgulHc/yhbkzjaBH
OkioF7WOkAJLmOUFSAXmvF6GPGyRDXKxaxRzu73mtYgOyMDkOv5OdnK1+XxDEaHs
iq+vddI5fZKsYffvVZfyGqYUAfRvcQWhcZdioORewLEcsgzI2TNvaskgx0oUShA9
rlV1FT75oE6LKeSxPp/AI8JoelJM0000FMBXm+1yln8DauJxpY3iRHXanyXn1dNM
Tg8sLhDW2r6gec1DKdFzVRsavdcCjQQybJegGLwITqCbnTL+tyRhrA35Alhkovao
4+3hXEJRMZ8K6JbMk8KyCnFol/zO6Q/MyXcXiYTKx8T/FCQmrh86JLIM2D2LjIGi
1dqNEIjeJbL5AqxGIh3X459co1l/L2Z46cOg8+Um9c0IUNTR+W6wQ/a3/8S8vs+G
zhcN2rwY34d3mRs3p2lhJR1lW8/zfRdh0O6S1YFgr19nrzmHht0uvRe/jI2fdVsW
YT3HjPapCL6pmbcoo1jbMjeezY5/THy17Vdnrz1AnVn1BY8P7lK21kJrAFlt5P10
IslKJ5yKFfwzIbe5mAGVsEuZjIOV5BHYPd6Lw9CzXrkWfabRVA2Fpe9hSzg533tx
x/h35CYn7YwZovrSHChO+qMoH8YXDRZXcaezw665iv9pWVwYHKPq8BPIJkI8Jz+s
IRulRgliZLupniKSt+j/HsF55lVOVJ+vGZZK7/OQkCB7qzw5xSXNt4CzPyt3Ijm+
Ln6LZXksckkjz3wcgy0qAIF3ps9DhaXGtuXfwdp47DPjAVNLwClqihzpPRjznBna
OCf5kKdltAkfUaE5k0qvcglnwj4Ib0PFw1WtNeQZKlDxVqKTL9CQ+FpCTIFhIS/t
G3vmu8kAOiVQdw1QEl6s40+VEgJJ/hSsrVsAprfsrG9EmUgEYcFq8xu/tc93zmZ/
gVQSGvD+ATzy3vI6DnK4nkgjIHUVkek0mGF0EmDQ2yvJukN18ZDYxA0cUhQNYVfN
4Gj8yzREkqFRvYDgKrE+L4q88HInq6uLgfMWQ1J8VCpOZGrZcUN826RN/lv5jIqf
e1bX1CrwZ6VYnAgCN74mie3fq+W4HI1eSApPNp4PvrVIEMJJDkDm5Q9gkfeta5EO
HY6j2DUeGgIrdujJ0zximpCVa3e+7uIM51bAm/LdJxLyhDf4XYP8Z1pJthCucXa5
mgriVEkYuAs+778h4R1IlVhs4+JYgxcMVYl2qJHxWTcCq9RRMoaAYODZ1Wr31DHl
U0lG3UviK2NKsSjESpsl1asoXiI/PRsGOcpcsiRHf4dXJU7PUwox3k9qLYVhlFP1
VLrFtF1BYNf06tK3rd4Pu/BHIowLckqJ7FaokTKnC2bT6r5dnCBO/U5QYwKJ+s3q
EouOWwCHYTZtU3QU8ifAlZxzi9fkswLwJFux1j6a0SYMOEyc7eTc2NVQQfc3Iau4
L4SZZsfqCnZNqUG+PMDbZHqvM//14yWdYpglOx5XzQJQwzanMsjERm0XSKq16m80
ry8p4mdhZcUxsr6l3ZmCfPnGw0lbucuUW6YgvREuEB10ptzu4soKciqliKYkkpv6
5gBGVIjTUmT44yrNVLz8GcOL5f5ii2++Dn4zRugR6SXcaPlc0owomcZzB1CSPI2m
W+uFsGz8ecFm6qXnRl3Z3tjY4UJkEmlF/tOihihU+49rZBo+8+ZQCYqrXP45MLlM
xvfhmGzdWMUtnsVXPKSEynqPhYoTd/0ddNoIxTTVZwVW7U1l9Z8aMqwp3/QJH6oY
dD0oKlHkBhV6MqMrRBE8dI2CUrow4MZ6ezRodEvQ7TwOu50aNQ+PBrawfWOJmKl5
XRIE0hk+wiOXBXdAn6CfPyh9Kh+wEco4HfC3m3YsYlS/IdRLu1SVhI8SY80S97I9
jSDh/E7BhCcLW/bf++rjgJZyAD+SVvhYgsixdhH49YiHvj+X0z4mrtmhFYbV+3uI
KDKNmWIxovzDHLyaJj9Wlz/C0v6S1eKBPjHvZlxBz8tHvMhTI22I77CYOYN14EHc
9ovue/KDkSnn6h77Y0xihUw7H+qnNRGH8KjMkoim+2h01yFS35ISG9LErIoGWFxU
pRGH7ZDbpkCv/Pn7tGW+b9QI2g3dTOfBgJyOekTra3G0SjnQKEKs92xzvWz0K4j8
OO7sfeEuq0VREHPaIVX4DgDJXVAvc+QOPHztcMqDd4WpcaETSPbwpMFoR8aH8Aif
lsW3GZG/zUFT8YNmG1Hx/vPRpoH769G/tsSrjr4eUIdwMxjeAFbHNv9QUbKvTk4/
FL8xtv4mFQY0zB2/ts/X4mdbGfuxFrvYYWimvah+IiZd2ThieQKHQP99EfuRLDSc
MLgN2RUbf7IZ9JjFmd/i07jXZsD/CeYvcJYjVKFYb9ihwa+6SPzR1k/0BLs5+0eX
PVEbSMLcUYigQlToGGymGyffTPbwGjx/TAFplsqbH0JS3lwMF4HA82ix4A92ks1M
/VYpYo8pyFwUJD4NIA8gcLZW+szQ1A/uUKQsqWzojySNkPk6+O11ycqYZGSCE11p
lv17cPz99Ea9zrLRbL6JtBJhk9zecC1bqUcKPo/IryPjeTn/XDBlPBG2DUcuGEpF
xPkXQ98VtpQ//bV3rrdwrXMbKMdaLWEbYM7LfF95uufG49l5g77legtgQazrThpB
+LeMVIs5KrjrtuOfm4zYGrlIB2GOFBGnefjs6HSD55sdb8VSjglu5s+glRWTsEHl
9PhYa/uMz5zVTN9iLcavChOjD+vXDqKD44XcMW9aKIXIpd3s9WSqzatumyg53kwz
8KEAhCiaq0lWzEw3BQm0eH7dmhj4Eim+eGEAboshqpF+8TLPv/Ay8bEV2ya4el+S
dfo0CSCXG4tZWY9v9YXeGRYeiersd/wXTobjF+XWt8tpOl1FTThUsaBVBZau+xtB
VK/jZnqNeFaLl920enjGWhvJ0IHvC5PlEJ27fdcDBy7Txkypn6XdRapUIMrvkPSi
PE4SZCg88f+XtbKgHvvXVMRwfkJWdeIclDtt/BUsccQfxiEU7XyXZ8AFkbDa764j
BziuefSr7cKHQfW+j/EHfXfKRtnHAxGbjs+iY+gx/9+t06M2UxvTCCAa45PQK7ZX
F/4ObgFVF3YhsB+YMMIFcBt+XgrO89aIW5qjeA0LL3df1kT7mBkWW80fq3etlgU6
tzVGgHRErUTiVVr+j5M0D1eCEo1eF72jtK/zmbspfVaQgPxVSdqHSnfja6byEOvO
JgxZcXoQoYubcovlwCICDwrQwZiVT/u5RB/DSqRorTVK+6nxYCL7kgDgwOTLmJ1k
Pcl9faEbGiz48+YBHNNKa8dqrLqD6DacRMLwDlupXnMa79xoKtcaoAJoHPkblHSM
4lnFO2IHExY3Sxnfy9/Mo8HTxgHTVfhk1yjXpNOJhLBoWfG1+PUbXsrDUIiJ6XaM
CLE3Xk7hiVPSA8S0lv/9P8uM338muxIyb5r5A27noRT07y/UOCUcGUUsL60/uXrk
HGhXj2nwf9tRPOKfjXsRoIUu9lfNWKTySIGN6WdxogaiKiJaIVJa9/H05fADfj8P
CK8G0RJew6iU9t9Yn4mifG8LoSpWZXPFjwvu6urLOHkLr9VFBdkJ5bYsQuPWnRbw
Hf8N+7AaRe2WCcEbIfsuMyzsWjxMKqE/3QsNA4cLlZ2rkFI5Idx7Xz8XSzzYlUKa
ygLqGBSb4uqIBt2ek35zJ60wbHlwuqusZVe3oo0WLq4ty89H1BEXA5R1uuhJFUEE
lMZsxu3098SbfYM5hTsoDUN3CwtW921ynPYsYpStD0Gc93KmaL6HD7fSjlPLAZ6o
FdhA7Lgqhb5lpq8e7bSWpZ8qN4PkqgmljyzUaH8eGTJkquyxZNOQMkM4QY6/U9dA
NjALiIYcQI2BJoDlgn+cuEH2We/+BsrQFol4H8SSOomSbuyr+hWAXxOen2UCTg0A
eprbY/7Lw86tQnkknKSnR+WmOr51m0kKjXOmuVGJitOXwJBfWfozB6QL8cWIapwc
lauCShir2GMb5zE9F9ZYrqTN+zQ8SeWhxAyntf1VazKLsXO2eo00ggTShu868sXa
r7F+7eh2J9TE2Q1gU+SItEM66l8y+tFFJn7gyOVyEbUJfjx8Qtg7gDgfnG7gznea
9LhCcgCdHdRoQrl/YVEhqLNkCOlmiYT3bYo9rIW++q94RO2D3ElYJVKId2GLL/RD
lVFUwJ35G8nCocKy7thtBtyygS/1C2+yqiYNgxEHFxZGFi58xtm6Lo5gBv6b/fuJ
ikfkmYIx8mDg+cU4EvF+Ja2iBC0SHFja9XT1MgZwmlLBdwhpQA7k+XdAkoXl06g6
bWznSVu9Bn7A6Xby6paZ66LziGk05Lms2lwRwBAsjCIqlh9Jmlh/5p5AhNlUrPOZ
Wx2b1oEdNTMPMgScKXXROjytjK4AqraOkt88/2iIW3N5ggaFx3npGYflPseVu0Lr
B/i/H1UXiNj+fgd9eAyfzU38vhXdjFdOQmQ4k2H7fYFbEg1AZe3Mu+bHcwo8bFUj
l2ZT+pB831LT3pSWjKWrm9Bj2Apwn156uIJJhtVQygYAxIrbhUZ0Et4S4/dNrleD
Sx2YXBrVOrmsKk77aUjU7Q3xG7Al8XbEWaBXotjCtX40k1bG6Iwotc3pmAjSkN5t
c7sKtglUIGYRGYwmhGYvc1Ps1PkUf0IA7y5P2LoghGbBT0QAvpqYaoqVQzVWtgzY
o3n7D3fe9GtZrIZhgGQzg/SvlMlcxC4vTzhG3pyZjuqNAYrkI5Ugerf8ogWTlokt
kXaysYdYWpgbWxiUYq8EZg8Vd2ZWQGnL4cYntaQgBHxHamkSpeiR3QWwhrjpvhKn
4T8ET92MLSsxe+3j2TT5EAWtHOPUCVXcCnU0oGtvgMGQrZQpXFJ2t/DgjHJIKRF3
TsI0pe0zZDosBCb6GfIn683sDR2F+387wubd/E37dnnmI7RYbaIehcJiSZ26Yyyr
6+bZZTxwruLe2U1h7XVARkO8N1Msaz/qUDUR3Cs3l51kycJn1WRHOrPUM50OMpqi
IxHIf/lTYjgLyvkXk/iEOUpYvRpwwZ3JNtyIlu5jy/4gvA3xIgV6O6bF0Ic8etwR
3bLc0FvXaX91zsob3phGUEckTNIGI99TKIZ9z0zugKgq5SjB1CCAxVAPw97kRpCo
DtSe4IWMd6cQuFb8ynz6tz6bRA41ugiH92G0uCG+8fPp4yze5pRVjXni7ap44kJa
23iX5V1djFJN/a7P4vcV0kQyVQJkpVCisOWjlplo2t5TFGLgt/BEyLxP5cQYTOwz
r3mBZIH91/cz04TqDkv9y/xYwr+oAto/MX1FfE0wXH1fjXq/vs80bmzc1+ki4WEQ
KNxRHQiHB6v0ZNNK/IQvHEAOkMUxRKA/mUm4ZLsh9Tc2dvBX++XPxezXKH1Ne7cS
BbG2Hg+b4KwukrMa3CzKF5zhYqIgGUJIu+OX/vWIvZHohMz795hjdi4VApfC8T2W
p0oXAl8mpAeYlgrC1fUbFh055F2B5O02YCwY+iHZt39ciRaXhhxM9frqvpnR9Q4i
bVlP1YcZSdz+7vWc8lmlKp/xvAydTZHi/il0xKUcYmqWEyO5ED9B5iHDV85YdkHL
3f3xSD3hWRYntcjMCdME6Lytyp/lJFrQzeO8oLdihts1M29EwbDcZqj3kmuoAkLF
R8+b9H8uZcFb03crNkdqq8uWy+Hj3Jm+iAADupgxNQfFlIEDw30kgW8JsMjmtDaZ
FDXEtK3Xg0bAkUKBsEIdjzj+rGsN1Y2PVx9hjlqGUb32QTSlavIsYxlmod0cdak7
4ZROLQNlYFXlSfcCk2kA5BoUqXBV0ihLHUYfJ+kHC0ba4xCo2CQhGDQBz9Rf08dP
kwFalpYpDt4daWTf59gFSzCZZLqhUZkczCBhzZRHSbl/MlEPcM8vAMKD84gsZkol
Yd2LfXYU2BkUMWs5op1aGzJOwUmt8o+RsaPe7ijpArP5c2dLii/vU/pRpSxuw1St
hi6f3mE03WjndZO29gWC1Tmxken471Y+xSOkbs4gQONcPi4PdCiaCm8LLLD7mzEd
H3PAuw0HZ+yokPFV4gNawDmlY4qkp11qJcNYH5NLfkOERKJDBn0LrSk4cZUDAxNu
R3HbLEAF9a9ZN/maWbRkvChlHB2EHCzpkzkWpUq72GtrSqyiNBtugZgrf7BP/jwJ
LfyhlDDakfu4LwKG8rtehNMLpB2cR3I9EflG1kDiLPF5RALJ+z7qcFRjIUbgnOdG
+e16AnqfVzERolFk4QOTRIIoMsMiCYFbuVzSA9Y3GPR3ZmGBYUGPc4VgZAY+++H2
5XDe5Zuq5CTEK2W6ZoIS/fmqz0Nu8WW91QmaXvK+4vQK/cU02HHo5yNzC1ZUdNwV
9b6rBNKAjqdxUmqDAiRBW8ivNyGZnq2mEWk+TPJMmcOGXALxqqBEJNSeItlhzNkM
N+dhb6cyZp4Ww6Daf40nqVji1UXJWO8MysjQboFZlfuJuXIVvo+4NUMYn8obtYR8
KB3kPvXbBzUa8SlbpDhABm6V1G/aOw8hY5Vr8716ACmX7RmVHAoUN3FITF42Oj1X
84/MiPlHjOJyXoWpBG6KWzaWxoQCcxOi7qQX2J5ENqWrpXc3TJcSeUPjAyEQTJtZ
rP3sXOW8MMWiuLRyjf91lH6gPfON7qZkJYVcSdcVQ7lKOQSxUjVZkLOcmvWgRNkE
yMBLyb5Qmby+h6ZEdPN9LxB4Lfd84CT6FnTGeSMcWRizTcOup5FrEp52k/0r34zh
NIxomvxCkCeoOFMW/Y0gHiJu1e3s8yk6QcqlYEEfM4CIxCIk1Jv07Jc2J2bZgomv
6KO1Uz8ucGPMoO+vXVO3mZWR8hcW898BOyfZRAeYvkWirYAH/oyVFmD9BdqO0BuS
eSwTOqkpTJDQDvDH/JDVmBAYhpT8ipSojtUEHVHhSLEEY2U96yb4d2BJtJ2Naldn
pFkkRnNMRkeOfGmwTWyClqy9h0YuVNAjLXP64462dRFd5q+gLXixMw5NgJgRuAqN
GK+8cx147yZXd+mnNFioIYiApfXKtXWboTwF4cPcf6IEUoxon0Sa/TLbTc4bvxtq
TFNdLk+bp8InBdZQdOkAseG0TEiTImQleN3NCqN4dR36lSS7XdKcqJzKxUxPq7b/
edNzuuZIjZLtW4E1NhAV0i/F6GdRcvb5P2v7KJ4cQeVmr7DpgN1APlpWOK/7kkh3
6G60oEf6Gf+acINfLel7pgBG+rWttULXTvZV93+cL3pD/SfvCOwcsL0+TTWQ3OHt
uOVhcpesUNa7xTWjb39Uywu6UczS2GmFAjT56aidhKv4bIte51eCrA1BzNqMrU24
TL7wCo/uY1l7nkKsMEzLrhrQHHJU6I2IRthnhZsSv0dePsFBxf66Bxh7lpQHhLY5
qd/EPej7d68BhTnfekpeFJoUe2Ybo3bn8k7VlnY5qfZRBDlxdrD2vNjXiIsBgOn3
ZNLJHHoAAZFo1lGhrMo6w3UR2duClsv/U7ILai2C6rnJJErTO9yvJHQUmsgmLbBl
C2SX+Q/sJjk8wJ0Dzl1Cq2i/QtolzbVmToiRmiUoeRfD6yw/D6s9Chb0QUTeoL+8
ZEKQjjkj4WSjzZmCqCaG2YxM8y2s3j2qtZKEEssQMEHmjL8I+FlXD9BedP4Okuft
TG4OKa8LQYYTcgN29vUNwpkaXbD7dvzcCEVgnjLQnSVf1YGvzgiTCSHmhXKeRLy+
Aoxtk2c+uFF6C1kt3zRn7zLmB7xyQh424i3SLI0Nxt3036+1tDN5LRq+YRBsHEvi
PubUr+D02SlcKy9aB2maDVnUpeVQ8cVa0PrJp4QL1P/NWQPtU3HjqwkXeGX8Lz/T
DbXcQnypbwvsnhBQ6EfZdsaBMzu8cjZ6kMNNtn1Kbl2NUot8rF1anfUbDMLK0/EM
lNtv/sO7GCVPOJ1grfpFBOQftiy3h8dkO2BPhq0W7pzY+MbmhS8dX4HmGQaQNDwo
JpRBGp8s2UxkhEiwDsqlntsU+hnFxJ9FZ9WGdgLIwUoIjqDprS+GNbt3tyoWlzAk
Cd/Hk8DT6xmskMw9TRf6N2ymStdTvA12MHlSvivnayJdXN0I5buJs4stJRh1P0Zs
f0Gi3K6yDgdnrdpFlaD2qc8ClF8uo96D0EMJxLn1ruzKJ+KIrsZsnSwL8mkBobGW
D9hSdCe2dz167VZHXpHraOaS/mi03IzHegLTd8UM/I7YeJhjVqy0uIZA43PZIuKQ
/AQMetEC/qbRkC/kVoBcklrbxt4FhrN83FcDKUe/FpiRK83Hnh56+gOpzseJuzXP
A5vFqERG2KnGfzv1Amlj6qIXOL8LGr0rnH//6Qg6O5efFLHvbx7kN+bM8F8B/DBI
uu/DW3fNgQC4O/6NZHnCCg6qzwiZp+5OZR0cyYOr4NEaTAqxJb4vk4Nkjd+M7sVO
/C0MCyDShp8e98pJ+Owha9OroKaLaH+G28A5/RbA7C7PVct3Jn0yamKJIfmj1sNG
81meHqn9plS/waY8WyWDz1/NBqdCDJ10P3pIRqnp/2drHKzgIuRc7ycCFlcL/9sM
ZnWOMtADPPbZ4hrZUIencAYOE0tpCUONv5WwQaciaFc12ishp7qbA8q9YldQGVDH
0xxpXWqFRS6amcI4mf7vkcfElbkLonjgIjJgNY5jf+1L4049dAvoqSu5UqiIDnyS
zeUojATUrBcmqaL0CqmGiVYi0ygXBdiCG0apm+Un7tbcSCdtk/QQLksjOUeHests
mbRbb32Fm1oOqI1yH9IFP+Dp1ddWE4Xl9bxnsKu5n4ByiUpnrX1JhjZ4BSljiLFf
oc96RH2SyhkyU74Nj8KnamoxSlRzWQ5bgGctLHp/d/3do7Rj3ZgBckvHO2IoobEr
3FPQwXytUwP+fUBRfwjiZCE5/vWcTPBXzSlAcNDTskQ1K6nfQ9cgMRqutJcQcSa9
siH9l7lqpI/hDoRdGSDYQi/Jq5OwwNbNrlPNDPkTR5/TorwGMHOUgKgEcw0DejZa
z5TRmdvNdoVCv0qHPZBidlgr3yITZkB24cU2eVy72BtEn8f9DbvJloF3BG0F6mVc
BgUxYt/nOPEyRwkzYj2iZ7Otf271X6StMzKCgFp2VEB34jt9QJpVeGeK9f/U/XrJ
B4J3lHPbTFurX6X9PGv/aJr8lpAPnKWdSYviSqvimVpMovRNr8RzbveUwsVB2oUo
SZJT29FxOImjA9mrP37TpSS3SG9Eh2FZb3HXsQyyPdUq8XjX8AsHAQy5T9+y1x3w
r66XUOKSgGnVniG8BEXfxW9NZkFPpWKsRUgVU4LqaEuFHibIcZdzME9vx6owidD+
higuGB8n3QLkVcXjUt2QxgqtlNexGU/6leIukyv47Ckt9flYyoLjgSkTHeeLUxSK
XFm3C4DMVNBiqDwYzSutg6QYYqT0qTlDzMaAR15HHEMdhV8r4KGo1q1Hq1pC+44O
fguz6d4yEkuCq3H50Hj6yiQuzs6KYpOFKecGcfSTpd4eAod95yWZJnxsnMLemRE4
PhdMbjwDadeTMT/IZrvjE1NgpPHtU9BHQivPZUPbQqr2WGEg/PnLA9AT5uRlBkWw
L7CFNnkI7ScdFUgBCMM2W5kPAVhBV4CWdQx0xAGFdVgkvg2Zz0dAoZ2bzdLQOKpH
qdEQNp7+o0dKEQ3HWCrXhqjKsvoazE3GJ9fBUEiBddtHECip5Mxz+CYw7UNgCtr1
ffI8bvS8GG3Lk9GBMzpgRlyp7OoYLdidHueWvqfjFKhCs53WshY6VKqxm0EqR5P0
1O7MRG0zwkTs59yyVa38FdN9UQ2HelkMFDn1kKOgub/N0ilXGcdpcYZG077esXv2
sjH7wXcI9Qz1NV/BzlbaG0P2PvAAjD7OlgYEJuCinplyDQO3aQdnPAup68HYkLwM
cA+hp/W4YjdkrAIYj+Byc29gNHpvdPKjyC05sSj61HzsVrEFVASS6AcytiheEENa
iVlR/LxOcvZ65Q/FUgSoqJKSXiaBJ7hLabZptYFt1atHnD74h75Ng2vhmlGqnsqH
ZUbEKifAzMHkaIkuD3e0YeXwP1+8jDC68eHzgt2MHFJBQ4l1Yd4n94Q57FbbF9Cf
cW+0Rhuz3yYWff8P8lWd6NVtKGtvDfFsxfF1FRL2SxmcRyWS9pRIAxS3hCUN3cki
Yvf9Mbd4JYPbLADe/I8agZpEvPFGSdd+ItcjQWplv+CqdsHC4ZqSmC1SW0219qxg
yr5vZbBPXUIZM6A+aujoOGsLz353TSQWLfLZqpFwjIZtlTGByTVwpM4VG2l6dZQE
YcmEK9vTJg9EQc852TsQMLiPB1BrT1obNTaJwxlFHNBQbl1cRYHr4umb5VgGhZgM
LYIH438CQqYx3z/qxrf/fL6mTKxhSKUbAI8buSMKDZJp5ZjY78rCm49ipNFWtlbr
zVGksgGfWevthV3gYsjJrHOZ6ZCHcJSo0kGovjaoefPpf4EZ5Rt4T+E4wAcI0wSv
lUcBjfmI1jjN9ap4XylMSHT3T1nkhgh2sQrASw976aWBOGXUhnsDQZcA4LU9S1d3
PU2EMtVA/WMcIweMZeTbRcAOOPGm1E2t7G8m9FM3zoMuqiVT/1D3/gg6ZLsOzkBM
tUULGe4vj5lIjuMxE1AUs0Od7ne4kODpvYW8nVEAVBVseftYpnpcuLdU8H/eVlxQ
sqCPWPN5QdFV66kOyM0+VO1p3tv1S4jA5Xjp4k3G+vBVLtCOKsGsOzkNL/LAZyEh
G9FO6z7YLkUBNOeQQ7xw5JHDqyJaI7CTw1w8K4jnDk482OHJe4yQNj/ThXAQm4KB
f3bCj8aNY6aS54HhvNAc+COTIFpAgsnbxRie2V42JlNcUZKpZn3PrTqG2jmdfhdw
z5t/QBRmQgqOwil+PpMP4JUPfauTLHC9zPn7FSKTitZOlEwgo36Hokush2gthccQ
zVnmmvFRXls8lU6+YNiIGFCxvMY77RwYT7kPRIp80RE6jSeKp2KXtMmunESfm6FE
j4W2FW2DqchzsQISW4qXvDy/rxrVXBRVcJrw7tWKdijedenF/32rLjA96jiKpuW+
hBket+WNaOyQYyn0bLakVog+UTPs7kCyCp4rEVMbQ4oU1S0VjCCjBCVe2A7aBsDB
7V8i6PoPe4H2r2KqwUGv2yOYjh5iRs3iTcbzJHhy1CH+IFhHYMpnMH9lF7a96ewA
Fh8ckR1qkhUv3NSpnsaYex6c/q670OkubqHkzFgOMQvJVgN1cuLYX9zu+B0vrnZF
ZA5puNhfnfucYcPWrqyyTstpMHQN3XzIAU9l/9LeLEtjmYpBos/OFTq68x79ydke
bg7ZrrB3CBq3c3cMoASul0f/3oeP2nni/X2OYsYP0yydLu8bwephFMrA+xMrX4AB
xSV0Vgv6U2TLkeq7hYQnsxQMY6pahQp+M5t/w3/6AD7Eq0ORV0WwBwG6XgNTnP5e
R5f+74HRvAT2YQ0yvvPre/OPLIXD0qE17JsXGMWPU/sTgDM4mnrFimAYzGtzYQDb
YFx6md40vSmVzeIqchU7taMb3uuJAiakBVx8lZWKtJ/wFTO6pts1kMY1Flmfhl7G
RrseHOu6/cbbQmOTMINDiK3XPr0XMHkwIpvarv1XkseFIq1UoJNnUHM/5DKrW6Mq
x4lmd9seH2VsDEG8qbAzdsl/IB9dqY7i9RcDXj1xOP5d05QF3xvOpGT8GthuYIJJ
KhiZSMxjQXFC+aUzxR8Yx/vm/b0BNmmMydbg4gDjL7ikqgBC3ICiHGzTf28HvfA3
a92eYnQi6lYSOEcxc7rD+ejT+SnzU5E2A/iFfDoOjIh/GQ+VDiVJj1OD5hrLY7Kq
B6P9Ye1dLa4Yq8W9WTKcnCFal1fE78RKUz+4GkUbkcB8mKXnyUmsiOUdvCoAVdb/
t0NkPTMxnKS9DHtwLQHOG1w6jrgkMs4ULdFl5zzDuTgKQc2sZh4THLTBfuOnsTWY
Jvku2joNhboS1HggUyZeasDT83nVUhnMqcKS8K/a2t7ILPdrb0WYauOkXIoq7cl4
n+Lj2SPMEpMxJE8qsL6E1zfeTTSu2pv4QsoNqCKYZxvHIVG5qqSesDYzptXvT0DR
AGipNtODQU7CrNY534jxEEF/YdY/vRlxEM8B7wJWslK0SlLYo65bD+85IQfsfkJq
su8auup2oaCjLNuODADfbCraXCEhO/x/5AZigjpr6LYMvgvvf35Jf0MOXT0aXxNb
WSZx35cywYjO20m9jrJ/zoU94wriXeQEpPUxb4Bbi99LfEGXigl43j/iJz0RL1gk
MwDDUJ6SMSrNXCIQ1BCp3lv1hDtSfUEE1UKaOyTiHrPjuZTNTvL7rfF3tmpSA3LI
Z9f2RkuoS+f8cG1FnWjoiAXISSuQI3JUjsnThSs0Gte2pFGjrLuvg4gQzHVCbDQj
S8wXVROuW849ZU4WkIOD6oymerlEhXqns2Z/xs+wZv4VEaxc5EGA89PtlH7UUDSW
pepWc6PN1YH4mOUJPwJYOMAtxdwQFlGb8mSrjID38xXEQsAgxsA84yEWmtLnnxYR
Rzo61bnHiy/pZtmZzDXU62FZj8Fiy5dbQtOxzz3yWdCGJTUUOKZov3iZJr7zGf1E
UHB9ZXNt76coC06G0UL1vJU8vj8u3uv2UAeuqKF6u191CJN1HW483Io5QyhSgWnB
pl6MAhD6ChMVq8NJMI5xygJ8cY4AP6VgQ6iabQJRLHpBpXKcpLoHAg99OIuHYIbS
s2ynX6pWViQGJO0i9fSr727ZHNV/yHLsJVV6tEzLlJ2jvO56+TJmSFLmXya9csD5
+AQHE7+PNya/miPDy6CB7K5jXj8WfX5PDHQCuJcKEa+RV2k3V9Nh+Yq9MBXZhPYD
Ebg19C+iA7rcK7nM953H0Rrv8EP4C63Q0IojRAQzJ7X10nAXnYXFvWGyadcnUI7U
mOIOUtWbTQPReLHqtjUKjB857d4+BcGYF9GGFGQ4vhNerRU2Zq0Z8PxXIM/jbZ14
IH6T4Zn6otSvH55J4RWYkW1/+Tm1Sd1g553l5HlsQ9yFLaynORGrmFMUC4bla5zX
IgbNIc+ZRxa00/FKIVHEKl7UvNPHt4gBVPYl0rp5rLyq2yH8IHglANwKyj/PRm0r
EdFCLaaiGUAy9miTZLKuuUXJlPf9SBp21gW7FwDHhzEPEgWcotIHzrumbzn6T8Di
BXyy73bbC6NJJAPTNojykp1O6WpVKJ47rYPIwFWJPpeUGNg9HJ4UFZ38r8Gysne2
XgB2f9NGO1M9uZGe5TAqOZSIKGjMcXv5aE+Lc3PNSYelEQSpx4Oolow9WX4JWSGO
fmQ7o1oTdRVEuEiPakMJ1QKbMpXr10L4SVMFOqnXdIxUZfl7/t6IJEjNytMkLKmd
UuD6I2LGbkAoh73UDTzSQ5bPZGTvL4y0s8u7+Vjt2TbfE5LeSDAmvJQ1B0vaaCk6
uJBFbOvkbCrfTFHNG4VgWLcc0H80Uq2ok1Qq+AM1y9iPTI7a9EDPbiu7n5e3I1XT
cfQzwm2ft8wW4vggZSG+NhQ1gR+NWYjhRFCHPcn8d+9M3+zuSOof7szekzjGXcCn
U1FBNzFTPLriWAuLIMeUi53+bhg2r96at0JSPSg4MccjExIJ48dGRQYOlw7aXBo7
q+7zWX7h+SL3Y/LgmX65jL7KX6hT9tOzpKlYK+W+VbxEBpkhIao4549EBmQCdUYP
U6twAVyEJYJcgmuVhA+vq/jIDUyTRNDH9VzS1trIch0tgccObJ0DHVwAC20coja8
dYnIkI5c8rscWR3ltONaqR0j2ibFhCGQUWCGFlOdx8Mpbh1SYW/idDSbQMqk1M4b
27qR1NIZABON15S1QAHAivK8twkKcPlYwBGJAjC0yNLVU7Ef2MkTC1R7be/FZuCP
wBtGL/QNVVhTDuh7212Hv4eHZwX/aOrYhwcX3haBc2QKGxub+Iq/TGAwQujVJqNt
Oa2RrXFrScY5fCcg9mvzGYOSqgeENb+CRknw6K5TeJarf5KylEymzt+2pBeIzy4b
VygKTbv77Xa+mB0zNmGQwgTjlRIuxoDEktcdakpU4gv9LrgstRLEI+W2g4BQFyN3
kNV8YJvM7KPLgd9e4baeOQ6h0FSM1JoM2MgmYIdnqx3pSkPwTqDbokP9roPaA0PX
ZdMCHQt3hMQt5m8JtSxgfM7/J1CJfASaam/eCPakEWzImLGYUHwzIT1AY7Mb5uGD
ampRIiW7ykBr1yz2hHIrjVCOeYqnAUD8PEmoCoeEh3xBO3eQj11Oyad0yYHtb2lS
8v92i+x9CcEaQgc+12Qhkp59Vzwu5k8/3w4jSFBjXSifi9kCCwoFkAtDhhmCLYnj
/UzFuOi9G7cgL2Lw7lqdTD28TwVPbiv6FCJPPoj+BQcTL7bzut1zrTr3QUake9vk
2EOXPuLZB7F1oWSJY+78c1FSCP8FbNjgQaCOEYy3qGm+73Mdu5COuWxM9wloJmZ8
MSqHW83Zzp0hbTTUZB8YVe1H0jDh2pFrRHSF/bM/ZZiz2kMlE0bA4N9wUq4j6JYb
qC58WYkUQti3JBLcV24YNbFT5TiN0m6mYNMiveUrPjBBniirHeJiL+ZisAKIttg0
WOfrRDx1sFo/I3wEfuE4a5EZn1smejqvYzuqzJMjuXDIzn9KgeuTqRxOnCntj8lf
4MEqxDtW4efgu+RNB05hKoQhQGd5fNXrB7RKhJkRFc8dbEmDIHsrJtNWF0X4no29
duLvQLX5GfCvwZ0VBe5MZ4z02TgxcQJRu26E0KzQP14Oi20neLBYrBqCdGpnM67a
58Yq+vnf46MW6UUzV8UsiHS1oageEGdY3LtYBC1MN1244vPH+J7kxeL6Ya3IJdNC
3RJYBJmOVcf786F27d/p5T+nGCYKa3K80FQqskUvX6YXfNTqaL6OYKc76uYR/bJ4
uxCfzAMkkLW4ZQRC47YWEM8mtLmoXlrA5dpS1bpgiRPK6lwCuqEgA8xdvDJ5Qye4
NkvlXCDpoA3x0gpus3gk59JKiaI+9kRsmPTcL1ofjrJ4OE9gaRRSKWdZidYG79Gp
lEu07GatGXSmXdEvYCMr5Q/SdRB6mzsLD8GByvFq3riCEpScFkE5WBGi3ZTJlZ8g
oignNOsL97pv1a4KdIYvXFU6KI8GbVtPlSba+QVzM/KetPQ/MC2lvgGCDVE7udRX
1zRC/K3kkoJqrYZBkEKpyWAgeV70KYqC8pKf3ePDvKMMVa7vTRDbvn0T1d3Qz2pt
D7VJmQEOUO1MAdnOp7Xf3wHIfm2HMK2k71Jlx69h1tJu4O7e929FJ+rNEwvQs3m6
8kDzMUNaUnDHEzdqDVAVqoxVYxdRMxHFabZcTvGRjQpn+XjJdFwOlxLoRR/jqwfv
zwk/1OyXX/BLCjMArKt7N/6/gzjfMYRETELGJm+lE3U64WJ02uvvftbECadrhpgr
NWxS8nsQ0VZB98MHyHJkOAuAS1Dlg9S+j1Kuk490CN+RQ88XC0tLYp1lXFWaMMjU
+88qDdGAlYh1WBvrQQQEZ3GwTjwmQbQ5nRpOcO7PaOIBQq/XWuboVsGYbhMVauR8
VDCC6in9AZn6/1xtbkQ0QGX0XUi4NekZe03VlWJ4zjjGaeM4K0/PnML6aiHs4CSG
O/vi0OU6cXXYpDGpSStTXSv81tM4MrSTWLBvam5cIkYLPZpHZUBO4RFWsBWjtcnC
VHHKrMtWVHd5eqwRL/MVDSAdQcjZZFbImuyqB4TB1oR0n64bLe4nUlu5wtbOZq4H
ilMyOP0TaPrZM/jlAmo2cK93eBp2r7Ooh/0nj9B+Z07tCNY906nAboBenR7h4yfb
MqQvSCQ16rOfXkv4aKxwfUfjECwwjUE/DSVUPnaOYk5eJIkOka3tOYgOTsqr5DAL
pec+fZcHE2y81Tra6nezCYhWDNjsQPEB1A6DIQ7GirK+PBT9iAaty8nIb8py07pF
Wn18k+ZWY9tt8ReB6c5+mWiPXALHcmfEkJPzYg3qQv7Ev9bJeAAzzdlKMP4RjuVD
6oQqRlVfZXZnhSlnoeVwre79Rz4UxY6LHBQQSBzRU5eKA/xDdCkvqV8PM+bt0qdb
zxm5nvtl6zZapPIgooJkEPmY6UjJoasDOzMYhjg3sYhDNxNNZr7E8ucgWVKbtqU/
LoaSR9bFb9mwknhDAMQLxKMshO2mxnQ733gNxmErYmap3UpzDRR/YHS0g6ROmqeb
nx2nJjj1LgLfqpiao93btTnwuqIgPfWYrPjjmVKPBLLQ8fynTaZA0CEMCbPLoguh
uZ3nU7M+bswwJvHdXNBEdS3rEfkGCzrBcQHuNn9KBAZIrX+xHQlLEkQwJwACexdB
K9jNjmBIsuZVePLYyOJRwA1HlN6Hm6lEp+R1kNrL9oGZt2OIDcTrob2bVkY+GFXX
yK7iDcbAOTL7dq7jiYpiU/aeFBDhjQ19lx1uPLkzaqunBwruZBS4JImbr3Z3X0rB
gtmZRE91T8HXLv84MFxA/5M06q6l0ETY2lWRxnAA2a3L+D8suaqcUhtALuFqCoLV
YVhPxWExt2Ab5hWuMbAoDm14Q38coLZJ0oAorSyRgS6crRwHFdD/ajHo7YRhVuNv
/PJNEPsUxKfhS6WMApVcMmy47YUGf6yxmG1Q0lsvjgVhGuHSFde9JehufqbTqxjb
8/8KSg3yn8gpoBpDPgkfhn6CiqkseXRxd8/90JS1E7PTkc3b1ZrhTDNB0qAm4CcI
EbriaPzXLCGMpUV++SNGj5ZwUn3qJ485AybpmeKd7bCFunPL9oYnV8ci3RUlUA77
ZGQ5LgjVhzgGDhRpBUPN9XCiJrGuevh84ZPvu60cDDh45IQ4nZXlLnzpfr1hiGvg
JedmrTHnmvRGTrXkEz6vaBWZFiSvtyosc1ecAEOIY5bKRuPTE0tUVfuAVAFujpDl
5P3VQLekAR8nNBooviWF7EQ6PM6MLuuThvSpv13CghPA13Zkx7P25W08y2rAarbb
BD0QDPhe6jJRVieH2OhT5bAsro28Jf6MuadOXMLszcpP0tx7oHpstSFh9QS6deVp
9TKFyu6OFjj2SNw1uXhGrGO16eXYf49m9710pmKcgXZ2ZS9+oxtTH7PFvYC/azoX
vGSRjZsxd53Q4rLndE6VjqsLaVsqfdRw6ga4Q0TKpVl8hCS3bkcQHiU8M7hAQVff
+S+X/21yI5/3gfStf1/FlwZS9qC/HuDxRb7Hq5mRonEVgDotnnnSsHf23PpSBJV6
qiiYZr1GKLyfngJlVXOQZlAN04fOd5nXKXQHaPnMa180GR6CgQwBuYjmy8/lQe0b
iDtysxyi/MqqpHmCD5f8N88l2BcpjlMGU31AvWFmjhEzecWxWrVZ2mdHSJpAjrpF
d97iMOQjyRDA6b7FnjJv+xeQGy0qQJmoA+amEvPITD3AEA+GDPhyryaSa2H+t3w6
0oMmvMiVSD/JySR2/PoYMgACnvjUBpyPvAJBfyTsJnEXf5QdDplcMtH5Jp7t+tcC
74O3UjL/3lVGerg9pm8SRFD5ZAjHUtPYMoUfSrq5X8wpAVF9zGceAC03HMnINJaS
Z2ifIefoVUIARA8EqStzHXazJJsjQ90HoTQzGdN0IXpUYQsNXgk1A3aknFLG92zB
b/bmg+k6QDimSaaIlcj8M9RFTpw0Jhmvmfg0j/fReE+H4qCLb+RygYi/2duECFsn
hVDK+Hr0tsoIKkTeRkEGugUudDVQzbKs3ON5uBFHHx00wQh5ToXNB5K0QWPN3BFb
+Km+FV71+04F1UNIaAJSxRnkm/2RJXMtqeVGeHGXmJ5/aCswgDyjlLN6JyTzT5j0
mi17fC/4QwVBtoqOyIgvRkbUYNEDJmzpS9Ny6yw01IsyFeGoo7MmD8lY0iZXFLp+
kx5yUWTDtmxUOhQyBzXrPoJdzS9hfGNgJbV1NyTA8PQKjXIeazD9r69QadwIbkcf
4r0s77WdqpjAHWNSG6LkOtGLs4ZITNiEYjlzp+1mY3fInJ4vUp2SKbl80uUWBzj8
nU8xgCHIMbouTsza1kbSlhFqEF6U0KN2F1X4anCzvV9TO+PpzuXHczEHSSp3BndY
zW4wSyj1Zxe2zHhB6DyhqPRJosrPR7UHvQ/05TF/HXlVQeZlYV++nt7cXRDcsQA9
l4IHMMlbFmQSrYyS0V7f2o+pAmOqddffmZDCk+9NrlnhPO+U6iaPx/I+E5MUaCek
jK6jQfWcA0zPaoY1BsFsYzcC5RI8jj//98VZU3erUcJ2ieODdUmnunbJ6B3eT8kT
4HBcRXHy4p0qDDJdzNKlRjZvyuRSifgV+0t0SyBaco7ZdBPg00vENG/5hxQX6W2B
e4NYtBNabk0Z2Ofmpv+uGlXIrCPrSMB4/Fx037/BsI36g8A2wYT8pSsxVgLfxtFJ
htmVMHMIS92GPOg60nSY9GeClQEieO18rt/l0egNRlJvPihgGaNNbf1xpe9Ustjc
QtyBiX4KGuQxPmYo9/5zGHHhgsuUM8SijLI06q9ckWp4J34hEwL/GOcxVIpYd+mV
2ynyFmMlJoOapczKYL9RS57AdMU/rdZuTGyVrNuYhe6SmfgunpstkGVDjN1EvFXf
JdFzxV3iZVLcb/2y4qMt/M6GIu8WSn9fZN8YkecZDpKKiIqy8z17opxK1KaqU/Bl
XKn5But4saEEiwR0EITGzjmM4lvce5y1yxar/kht+o/wqqqCh+nWIL01iWIH/gwE
8USW/X/aPTit8zZv7vF+a9SpW6GbJMfwGh5+uRXkjUgyoE26QvliorR4qoSkNV8r
JOxCp5dYQ5qBaABsgH0QKSHl3BpupFcIMPNleQyODvpymwIQ1rhy59NFKG0zKxDm
xErWdWWqOVQA16QVctWEixjCmxF8LlYPAszHILxrd6zHytYJ7a3y9sFOYkdOQK41
E0AXlHtlKAcB3SYHm8oeU/Au3XPKHv81+mRx+Movo7QW4wDoM4+fUzs6GGxG8+MX
2JEl8iHES0s5I0DXwjLVNvUXEc1P0MnoxsUK2YB2XVvE1Ba/0I1/iKTt1GSlg2Ux
rGtUVpMKBEx3zSWaYL+KgkF2tNSnHf1wFZmfTzKDAyh6PWsm1fBnR4H1+AuenLDH
Y4Jq5xaL0eUsKjmPnUtQYDrl+YxLotrc6y5koVjAlMpOdYeW2bBMxdubUfQeJzeg
+eP/iV3HTfdKIOaOViMVJR0rSHBowty2lAkefKUv2VnyBVj2jebqps4G7sYf6boQ
dllHU9t5OAzq3Pn79J9xfGkUx7XFWvedFw82SdOxTESZv1P/ZihEoyw8zKS2PQds
mIjZLh7ZQRF3DPnJZq3YQaHJsEKSRYZXEbYL/0mkDZXwv06eLXVODqqBLRD330Bq
jd3bKf8dFeI9sXtaKtzRIDh9jz275Q2sjvLtmGbfxRqoEh6omx36aXW18MtLEGyI
RjKsACzYQHTIr5I2WKfpa5TqjYxfiLfog7KTWRU5wghruaZM8pZLmB2ZixiC/Jqy
Apb7McD0Cf0x4iax3FIJhmokjjt1MbtFYl7/XTMiZADCjTWDUdsx2e5FuVtqQ1HN
GSGOW6KJhjuGkdmP3XDqopFzToiraLDKpyWqVlWk+grDC+N+dGqf0gOn4K3xbxxc
ROF2R5iWUU1qhwAeJgIbBHRro3TePojgLyTza0n+qXGlXdmCMfOBBcgqiywFECCz
MW2tmdghnB+Xq3N/W8u91SkEFczAuZJdmoVqLrpmlw8b6ikQoeePoQ/fKtbtaY7w
It/Qi0mvKjMmI8iCWiOieQg0Sg20Vm+s4CETezvloKC1RCURzF1spLDhKA3jtqJd
Mi4rYjdFOyk9RgjLC6BrzWGR91G+wj+XDlH0dZrcqA+mkcdSoluYk1AWzE5Vn/m/
yS3G2u3Rt2ZDuST2Q5CaOgk0Nm50GFWqznTMqkKCYLAvq0+TXBiOLDU73TBUNhUD
Z2XihGjQP+bc2v/RzK5VWoGoR+61bMYudmKwSoDl1aj/3Pk6rzUhm63ZSN8+JWJ3
UUC8te4EET0+roYlCycCsHCiv5Zm3h3QD7Du3zgb+rio8HUNXmid75heB9NHvfJs
4t7jhqMx487J4GCn+Gz7CYFZgvHKSWZhmVVwOTrovpyFA2AWP7PME/faJ9oOCvWn
dzhBE6w+lD1To7YVvwtvM7IALoupyR9+BmpUFyGdZMgg6kwoiIsacMKrzOUSXQEz
B1a51xSYuDcLPq/FAM25SFGiClIEM4Weox6WdXQGUOiF3c3//168i0/Gj0tG+Agk
KsJMiLjqFUR2SBnDIBCAul5rHO59GFY76tvkx13lMEFl9POT/L90/weP3s4hbLiv
+HsYiVq9EYyOnAFGQ3YWb4oXULKhWnsd2SGLiqeEsqIi51Cz2hGSbCwJ8+g+T1FA
4ZOM35gWvfGrAUITP7BgkizxofLBXFjY92vSA/WC6AhcMMGfzXWi5xo3kGm21AXc
9sOG+UlMhb87i1j2a2XZW/xMe4Hm78m0OEROjQQ8EuIIh2VFmSRz8hWOwxDi9SO/
sADGKsI23/8v1m4S5ABauM3vsvu//r5lYWNjUmxql8C3UMVhkuKPoLhLO1l/rz30
GxsiZJM1hQp+/AR4S5MGcdsGCxJ0EQxCYNAY9lQqQ74D26DYpgqHJCBJj4nsQFew
wlGYGNQ1ZVDGbNGs2n8CxUKneASoHowCRA1LWYAegPoGGZKWr7ecCyeIQ5j8XXqu
SKcdBVkZNKEsO3Dcb9MfT57G+M5OJrc+2G6PTZag/FZCm/mkW6ky1103O3XBgVBS
MaC8JL/Q2YAKSldgMvT/wROF9pQSMLs7ThAPu1tyzEIYm+sHslQ4vN+l2ZwzYYSy
iju/UdlRLpYs6xNkcGP/1ULRNNxpeQ/n8b2MQJNexSn4fIT5Ea9hGIzVI6Uh81DM
qkCk8dPRlLAVBaqOAkRhadr6tDlk7TR6wGFJB3nouICQHoy+ISxxOR8RdQxoaiBN
znaCW3QMiUyYpynWXDWyFgIOeoEi8cp/flHc3Id8HQhsEdm0OFv6/MyXIMB46A+e
cVUaWG6j9eFTR4KzeLDQ/w0Tu3g8iYc0Q9Rbc2DqYxz6TrXPdtkhlR3omUth9sXZ
BLsjqCaiIOflO4MryOPp1JESO/xkaqSCnFmk8YR5UaF2rNdOm8dG+UgFnlB8JSnR
tB2qyeq+/SWfyrVOE26N8V1yIcVrqpV2yMtOf7IhyQ+jM5gpwEuOqOZ1OwVZ4Vsm
FEBT9dYsSTyISj6NDkESz+dXUMAxaceHxZyH9bDWYD5tVA190FMBW/9B0Ymr/hdB
ksY3U8mh8W0dZ470eCgmT302Qusf+gaGMa2qD/LPt6czNe/UHX2CNBZUrpwQCH1z
T3bgQJZxZeOFs0nNK9g5fVpz6L0SlV4o3quW0OnM/JTKbL/ph4h7PhUDYN8tvgnO
cgxuEuN82xN2jZrrL8xWZLXnhIq+Qz4qQ2KYIvYeBTKPoIjlYLRt82Y3ZMmNmF+P
U/hSUFtnXo0s7Q6K/MT/Oh4aka6h1iHnCNmftrD73ValwNPYbo6mPGWUN2gBW44b
KGf7e9K4uHXuztpRQAnQr8ep/DcrEwE36nB11Lurm+gXFTNBZPWinomXMCiNZm3B
Nnuqcn5huOG6MRFbN7H/IixpuShJ8Swu1vIvVdERq7W68ppZ6YUgWjirQunBT9k8
foBxUKLYjJqoQXlMP5nF/9yBv2MzSmFD6rQZAd7nVEIFq+xw+V8N477lVESIUbEC
hcqNSvUwtlHpfeHB6LF3FD02HrIJbXm4JGu/MU2G+fvmrfy6l4f5AfHaickWZRHD
ztAa8a9jr7VvXzua1ZNV9TQLwUthUUy6j86lsYZ/UP4b1hR65yzkNb9yMTOG1/wv
AIBnec6OgbvKeTtSiNLOmhZVMClPNB2p8muq6W8hELkaHOa1XV965LZiVMMHesE+
r+qIpGLDMS5iQkwfi/0tG2xWrN9bzyFqAqjUZw8L+uk5pXIvxIzul0lj0gA/kwFb
XW3aVRBp2n3VoJf9TK09a3KfOWfAlazBIAHXTQXH/KkKO3UQ7gzkMkfL3rErot38
o0rdrnaDYjCecPE1jChZld4rjT7E6J6iHk9dWEM2DKczmCnyXdq+gtT5nc4DUNrJ
HrWMvvLdfeHA28cCZTqKgjPeP6dtqPz9SA88TbGRCRXaZbN+JjNmol1u5ssKbAa8
4DtrwB9vRjVvxYCfTviUpyWkV94ATwEZrLcGnjlEo5ibEmtkkPhFa7ddH3a0TZts
LbmN2VbkLUvqKCC3crfqdVxEyAkM7LRdSGqjy/TOkUXvPiptHWIpVfLwFXadnw/1
A2qBP03mqCgR51cbGdo5uvxRsiP/JCrqBYzaqIg+KvUTT7aLmOaWtDNW/ZNTP62D
vxQ3YFdTtCBZ9qJs3wSt3uJpRaqeDc+PTadvoe8Bd0FdJCYqk0PvHtnnn4BjHM+2
3jT7A+VF6n7l8kQenWi+8e6J0Eg4TAMpQhNIHLI1wGNK7Qzpvi9gk2x0YjM5UDyz
gZ6OrFVsfjoSXhzh3g57Zntk3WpmPlAwTzvshTdedEnfSX5nmBy0l4O4Q7Gi6RgL
Z48Ta3y6rSM0O+WFb8jg0V1QUYqgea86jbPJvgN31LQCB1IBGV3lxhTJMKnAdHsn
OqRDuENn9WaP0u4y3R+s03tTuX5uouYW6PS2zRLfTbtsSSz8K+hn1H0Devr4Hvud
cF/TsHqno4tspq/jqmv+Klsx7+NZPX66sr8i2x/w+hluW4bJoafzjxFOhAORbjpG
x4a6HShD8PDm+eudezo55ZcPOBABYLG6KRxIRm386JDRXieGr7iezaXb7fUkOSML
yKkbA6PkeFIK8FkeQAvrmCMMz6KGh9cudgYsUtEjDR+ZRFIgalnpx6J4FhvrqN9N
Fynx8pB2kweMn3nzcADdY5+QpLRUv9oDIbis4rzBoHHczxjJRXxnh9ZQs9G+K4Jz
6/+Wxdg6XzryOZjc78+mxjRJXxNGdt5GOaEgUePnCroEp58YYx2KaPSnM3YfnQch
lK1kVDByguwSFI3ohtkNrPeYhIdNiNIUVjJIsEVTIX8Dx7lDhj+TQ/9DjiSMYIIR
ncD2LBWg4+QhoKvFCaKsIzZpMsSGv2FZCnoz+XWxEHFFr41mitH++st5JngrqkRx
x3WvYI1QnUJLWwSNNxdVYQA43q9UkN9650kIBochEpZESjpRSIQRrylsIzKTXRU6
figVJiVV+OfTBtHk7pbZv2b/v7zyEYyFd5NFw2FvrgTfwVPVaNRVSrR2ycXDYD9b
ujQhtstl0GzpIC50CaGJbmRptuGqzz/Xb4HQvuXaXDEF8L2RWDlm3RuVuQHW8ejG
rlIvTd8WM1+oukxSVNVG6+w+X4HHaBQgMxiNZgil6p6l86D3NLi91ebAR0TW1LaS
dyWx9HG9iYleW1oT8pH7hU+g1GtUp8zk3M6IyR69KmmiFS8lvUleAm993/sqprX1
IYv/fhRwIYxpNZyaQ6fWZlW5sKmPYT+6Xtbb/s7GQUQF7bYWqt6jn3sy0tYFK5y3
PwQJqiZF2hIke7R6+MOe+Vum0v5xoO3/UEuJ5Y2qgAcGcuR8wBNAKWc6H1XZUh8B
seEhBK6VXLhCh6cpJk0RByj7tv/HfU/lDfufTotFB37LJGFOuHFAtPiXs5+6rjEJ
pqj3NRz97LIos871QDtmx9OcR4nbevDJ4hR44XqMXd9EYkjmRlLh9SKxH5ZmX23D
46ec6JDLHkXLYZ2SmYdCyxtjT5UEoRFNnnX0oNSSbEiGloX8LA8eQEpxNEKjp0fL
HPF8e0rG7MP6Cm+ufGr8G+YRrXUmbEFg/zj/G7O1gncmo2TWt5Tz1cvvwJy/2BWU
KwhriNHQIRoTcofFA0xJsfACOwIMfyJ1wfoPIHQvw/LLBKQHS36dr/9Kt4JB4OZB
oSxbJiwKPgk7soJLfvlryUvuxR+fdVyZ+HYi0+D9qD0vg8lpWpzmU/8d2m4y/Ri3
Pfdqi4cUCJ8NePXoh9iW24dr2te6cfmj8/HEM8GV7wCngViSpfEaLxy8Dgsj9cR+
LSBhkJNh7If31HvHsRhQvXXL+6yUZLZ0O2hKbi5nnv0cGSWGFFkbk3fDWlnEaEZD
vwCZE2j1/vzyP/39h0BUN/2l7zvw/IiCqZnGVWm/4WloD0hKVtK1CmVS8QXIZg79
kL1V9Bl+teW7wUnr3pwhfB8QgykAU88VHZ9FiJ0tt/wCCOM9Yp55+mLehKOg4IZq
H3Gi8fpPHSvybseJSK6qilqWom5R6D2EvYykY8hvNyzZOhRToqGXv1+EGcOMOyii
92RoBwW7fCEsL1ll0he2hZu5pEj7VAZM3yJusCNx+y0Q7AnZF2ggLDTT3/GrIXPb
HUPCBkLPhhF8VYevKIjxuCAKrk2D89GCpj5mZDMSPMafIn4G3l+OOr35zZkkBcHw
jZeE02Gg36lLaSN5dMKsaiyJrGWd6RyU3seIAu5SafFH8O358Q1/GLyGCdMAUz87
xt4rsqNfuo9opVahDvqevOjHVP5gyUh3qOvSdZuCqiOm42FRpODQDWC7cbzkXZMI
Nlnb80apOtB0oGk2kCyBlvjLn7L5QhOcRMzrc076IdYiiao3hfO7j9vvorpNEJ7C
9kJ3AZKVkQM9jJiyhJy92IOEZFaozK0FZASP66a3LJdIeYE6USccPZ5YzrtQI1I3
sC+kl5+xber3jogl78ljcqR3IbBx8HyihMh0cSLdcS8yXXosp5FWtsScxo0dPk3b
18nGCQnLh/z5lOmuN/+6fXHpbwvCoyRv5j9NCZQuXNy0P3DqrBV40D9tdX9J8Qrh
tCEoiN7XYCvNMT3kWkdNqjJGc66JN0TkGE6KQgl+3p9FD+5G4+/WhanevB/NkC9q
qc7zXTetwIrhwMadoa4ZfIHdyJrNGK5P4U6HUQbLbUwiOty8QC37RgECivqtusvt
SGxIzAsq6mQE8Im1yNESRG4cb0Vhy4O/y0YcRaHu01A0j0WpxTsbg2/9QVbuJxhJ
iy32kuLh4yNMPmB4SL+ZCajmcaVSQMup25v7ZDD/Os2JeWD3J+gkeB3NKswdEzB3
tOW7VDTPmmDajNDdfGx4PdiLsgll5XdocH03yQVad4gCxoF12Oh0KDIEYuLoS5TI
Ba7H13CRXiuTolkUsZt+HkmCbJtYOGJndB57tNEGVHoyaRZbGI/m4XcH6b/kbATI
xgqZ4GaUZxhcaTkEZv8NJVRc30IkRmeOINdjicoUWfqtgaW3nTsTKkVPpqOub3K0
Fn9WXFJZl9lAyPB/LMpv3FdwvGgllmNc99+EkkpNGEPpyJ91y388IJ5c4A8JqNmz
KO4oBEEXcJkZeKM+Jl/CiNcwwgkQ2nRbphWMiWXlBonRR9H/7yitOsC0Dwdk5sxB
J3eS4voxLwXDDwssRN6+UCwo09quhirT+wxfhcLumxJcYP87+RjDE3mSExh4ubqX
MPKxX2Pm5sI4YXxrzkj+9hnU8Kgj9yrgoDShYb6osszDD4MKpOwJvn9FLpsXj89k
iZsuzolLbGCVmf5m0vY8JWKrbdrSQQbQTykyPJpSLmwBteiBOBUIW1V/l1AWiG26
mJ+dJSf8IeHaVAM2iWn7WOXLP3nx4kmgttaj5s7FCsEey7aFwCO4rEZ5IFaIMZtD
9X1K/2tp7wh3s6m+r5kp+zsz1MjT0/66GJBZV4ZKsKJqFk2D4/F4A5JG8C58dBaR
FTyzo3bZDNXlYheGdnRD7cx36GtsSjpf7mFSbyTe0IX/jnFdi7QrCj2nv+r7szbg
z8viN0rGC49DvauVB4zhSDmFRwSFsRw5+gpyJ/1TcM3MNW2eBPb36cuQr5qL5CVf
F7KBDdAlqYSZvvsWqPEVijAnKnZz8yDeMl7hT3LxoWksz4iF7k017pPy6Z6ddkqc
fnLXmi9Yvbt6+BEFoDWfsrZj4eMVMkaha4YzgBgJ96jWvm9Vm4Qu9zy3MXhq6/gL
q3y2JEa6CC46BhiDR063boGZjEA5FjnMc7iin2dUWiSlufaRnVxAd8doFIaBLp+h
Nqy59/rkywMU5Rtyi9PyS6f6CqTB1FFrKJDB7lpbj5azbtc10QE6GfvoyzIsljtz
qIDcZD+hf7MlFPo4CU6Hvtu3MeuRQAoqsBtCIt9pbG6vW5TWXfHhB09Qe0Gy/Emt
lgb9Q91KD3bU8N6KZ7BnhLU03V39/UNSvi6hIcda1DShAUdrGJ74HZq4TO5UyS4V
Gnrbh+KHCldJP7OwU1d4krEmn4/KYweLTw+2IQeIOoF2+Ccb7itER+OZpd8+grMM
nmK90ZNYHC0ZmBM1Yi6bLFBIu/qWm3O/8r0SodSpMIWBvCIL35xjP6QdioJJEN31
a6kDUNKR75b8Tqxd3DH6b+KSyTNpsRzVJw0kVHgRJs16hJosajPJBqPO0x1ZBwtp
urbvSqRiqlx8Z7ce1QhWmfl8XieZtkLnb6OP6+ksyOxH6ERm/qOXbSkNSdKVp/wZ
ag3oi0TKOrBXMs1tJEawH7rDSHFzD3b3nCjh90BMFU0vVV5QXUKdoOhp2xQ+JqM3
srtsBmS3GBGQLvejMJPAM5nisH+PUSG4f4NSrshGOUGy48PgS1EB0jmJO/6S1fii
60dM+7AbvDL/ZfuH8EByvhZfZolMwR+HvlZVGB2kMc7w/Ai6zGYR6AzRdjcO/eeN
Js24x5VarRhBhw9XZYPhGWRba2eXQ0kPE/6j2pESiJUG9/oFPVqb7RP08i1MpyVO
rET+BYXYiDYw8e1f2Ql1++eTUe0pCFeTiPr3NUQnTbUPsaNsb0IROLKT4VCztTwr
/Cu4bNoCCLMk+VmDDk7rO7hWOE3SEy3fQe2XL4Y9dJ/DlQc22fZ6s0EpYdVJJ1iv
nzm35ZzWF91mJx3uG9FmmQznlICt1atK05oni9zW60Mcyl7wlUARqP3BV5epXNj4
y9zXtg2dsD5xzeQFC1JA4nlm485AjAmXtepG7B5zy0NIdG0RpcltRutx4BzibF8x
x8oLBFeXn+3e/yltvA3ikFPpADM07aaAmUXcpK6y6KWVy8tFcBL9ARQt5eULAS06
1zkQVExvh5uIBmEgNxBigeYS923lZ7cNTpBpVR7QPXcmlPv1X9spTG2hzvWTb57F
Efumor/tHWzt0cr+QHvLzFQgu2N4YuibKiIv6HdL2cjVDpr/C3vblNiwqfviRfai
qpWPdv877oilrwsCJ3L+lom1Wwa9D6cRqZdks5XW0NDnyRCOV6hemMGuTj69yPqm
AGsTnMKzEQnq1ue5lcejnSB0Y04ANFOQO5mQy9d4aUKSA+WyhqmG+1K1WWXqNPux
hbJbw15UKS+RKGUHJWIKHmv+71Pt1vOrjuQBhj0EFu3UK2FxneWIJ2NYUfVjsbQ0
oPg1xS9wRFOIi5R8uAXttDwAx+7CxETg3Fr3xXxdIg5p5h7yEUX0uPWEMVI7U0OR
8jAW95UpP41Iip2wMFZC1y4VzUwVSHxF29haMXrY6R2veRHXVBIENZ6mXdcpIr/b
1zcmhD8O2s/tD2iBng3Dg6MYKqi979ETKWmt73OlImLIkK9GjSmbusMf0nVnsdrh
pWnuQl7ZQaozi6ZnkMUsMFDc2fA+i7t6oqyocE5rQtnwgvcseWdnAJSjhD4LMALb
QN+d1NT96SvAXQlpYIoQta3DWECfBmi3KxquJhKRuUBtvCcmg6Cq1cuAJK0fHkh5
JbhjJw5JL+IiaGs90fqvMrR3t5YzgYnHd01abvBrkhnbIa5Wotq16s9z3i9kiIgY
jGTxubJwCI13GlFL8ehUNwI62UTtXb2FG5AwOCUbtYB3LT8Svm7FxgCPuNbekOFo
VsYexRhFqVjlSLiymYfMLnk3WjBK7wOFhHXQY/RQZi86XQuksFN8T+MkJ0Rm0pUo
TELZ9UbQsN19BPLQUzuvncZI78qAKpuBtDlQp8Q+5/OAqlfUrVD/InY0oKaRWXGZ
3810HZfPmzTCHW0i60oHHjBkg4+PLc0XVpm0q0PJRMI7m4tsmhb27SZ+60HCo3Ia
zihmcACojjnrUwzzGyPVY1AVcGwhVULlsYSdcGKdd/UJURtYtdO+8r1BAOTkrAA7
k2A6kuoHbAwrwBuhk7J96VPaQgny+fGbZSEUUuzIrTWTOpuCTuzVV8zFzvlmBYXO
yCZhDk71OjAa3SZQNMoT3NX5Jf8kJ0+5FJCFB2hvDFVzr9RACeAx2MftFEnX+NL4
Nh+VAfqYhJb+vo69ALgWVaw1nyMs0xqhcBVd7KiGCjBIZXkxs5vWalP2/b/VjzZk
Sn679T4kd3ezigQMZpLOsQ0NKmeSfqfLwquBc45RxY6cWblf1ai7kgdQSHWALNm2
lK3MbLUbgKQSNyTeBoM6iCE0/yhBGzt40Pk2Sw4Zlw7blsQR3QrBEwenQeKjFoKa
n3I2SqL8f+H/ag7HDmNrr5UWOat+M3HuWz7bJYJYxbGCxLp6ZiLi7zbsDDzQYOmM
JAHxtKklWATMM33VsSpPck64jYplRrSifHFW3nkC1jao1qXFXNrah8vJPLf+2KH9
occWsTrv7LJ8qHTxZEpgbySP1P5JGe4J/j2lNk8gyZaKpLSrvmIVdkVjGZlv2HVH
EHQphL0g9HQdluTnmAB6rasKkDdgd8F7CaqOIestp0HUupJ4kDXICJuofGl2nH4Q
rDVLKf8xPhNSHDBbgxuza7SgaMwNBnYJPL0ZcIaYH98Fz/nJS5NU8EfPAB6/YL1h
5VymufBYHuL7QBdbDI8nAVKHs6yjHscKtmKeSaMgfvqr6KEylu3rl3xkOKH3i7Ps
J48DLwkH8As+ohn/39pjnFKTlVhBIIXPPRYGb5iRaXu7kWKpWlakRwF+HVaSdA4g
qNjkdQlaKkN/ZSoKeGf3R/ZsUEUCKCg+khIrq5zweyLPrCg1y58Lgb/XXOCo1rA0
yQRIHB8iqd2Y7zc4YP6FX1L4451dR6BHEPrCOMiwt8Jb67rSFN8B9SFVsBlYlPev
nsKc9F0OqlPOcwDKVEl54NDLeOtd22VWna8LcpJqBUB2FDAqRL7eqlVyq/DYENQY
342yF9lYmFsroYJr8AxeG/P+9e4zc6HpvVtwIhbR9qvKhkevFY+vpglybMC1n5I0
TFinYPdAeLPst8+X1MUrHQi+NW4GrVWCue40jRw/CPtbCdfIS5yadO7IxHmASgdH
p2TEHOlASAkqyFY01HSxkXv4CT7+UNRGXGK+t+k0om8WIlNhV2ijChFMflnZv+2q
8qDarcdLscriXQCaI2/v45beiDRhmDRffE1z4TfPjFuDlYVcTgHL6UJAAiJsvpAU
oW1+k4LaWiorhOmQH/5LWZvuzH6EH1QBxiJAlb31hKGxVpQVsQ8iCUXbOuZd9JCm
jfebneM1lJnKnhq8D+RhxKErGrVMRzseCjbf3inqNpI3pcji526IJjvXN9x27pRm
WsprsRXvgKQL7U/IRb168fTXraJJR9+hfBdnd2+MXMzvfsz7gdL7od9RsdBijO+C
VyE8BFkl5MlWkDaFOC1sPGmJW4yQZ0dbgbHKATo9v4eLFTB2L4dVPLowzi3t00Qe
w+7vw396UW43jyxrH1Zhxf+GJ616ZtLvkCjXLxbmpGp01R7Eu4atXjHAH6hO4Wvv
PXQLSxx3+/Obq7eO9Wqq0E/hX1fQymQWbU9Ns/atVNmRA2bsxIX8ZgJe3s3hvtxp
MHk/egTdel0BiRDWaoSscyXddokQHw8oqdzD0Z5I/MytZdO7F+VDD5hj7PI9OmEL
4u6WtxBnzkTEc+S0G2pa5BfDAMMqv87ZcaAH4hot52yIQvQMppLWWXmvpYAbBrOE
LQAvRkATfJX6GSlH6AnLOlhtM7QrJxCl6dwiYUOqcvkOvMyIeJySC+eWStCF9Sqx
WDTRS4EGZdIzlsCcnm4rAPLQ25n/XKT67YcLpPDawYM1X2VIeLC0pAh2l76MIzq1
IsdLzggxR4DkA7rSXGzXGlHiQPVojbCZ/5AzqEsHmBSQ9gfXe7WhSzOjpaqGLIb6
ddtUGQdH/tvtB+KamOPonnVcPpGGAWO38J/Z/T6PeY6vCN5GRyaXjUyAHPAcU80A
hZRH0m/sp6Hm7t+iN8pAlxMSIytx6OCHJthKUQThhvShwise8dXmuYYaTDVsZdwL
H4QsoVGbDjvbvig+LNGNMl760OE89TLmqqx5St/zQ2lanRhiKlhbohJ45wP+ijtd
ujlRtu1JzCnWIUXdlmqLuwwfn8aVLya7y8lo/kSXlIGy6nm5KUx1ZYiP6uUBRLD5
6A5PzkyphPEO6wzLAYNM3uQyMGeX3ycfW+f0+Xp4N8p/vB58CMI1J7KkjaT/+3cK
JO+/JnKxinpKNrBlpzbfOH9rLpeI9WWMGmhJ0ZhuaF8nXemL9adnb0cXsGvDIIyr
HvQoU82if4/rpsps3icmn8N42D5H+LtPFSduMKhp6KbjCA4vNA3QvMrgem610+HB
RQmEb7P4GUJbw//cOE3m/imvLjpjz+9uWS7A9WcIEDyOvLCttUPFxL86jHzTAocc
f5uVYswiYa0f3wjF8vFgwOoAO1+wQ9R5sIMfCl4pgo7DVQgUVxhfWcGd740qwf6C
gK13mF8bbgux/cz4womlFZ0zHTKgD7bVyLFT89vpO6cizQHknbybJcZpG/VF1QCZ
8Si41/xyi/NbsbTy3ZkTjySleCkpxch758x//5x0p5Pj/J/+OsLjCAEZxQ4HulEF
TDRyOwqgeaJZTvazHiTaMFLBiHhPOd7atXAEe4U16MJKfRuklePThdiX+w8xXYPS
hmmFIaDtWv0EAIKHc2M9Wv0MO8AyIMHbR1PnIfrh5Mz2Cx+LQiw02XZ5piMjf23O
sKZPlY5RvzdSKlXjGBxuStKDwHTSrc1tg52t4tQFnu7UX8LTkRnOJkeB27vrlki3
RJhJKwtUnjAv18j72OW9ORUlOpMrV1cpIhUX6/yS9+tDWjG49ORom/bA0lzvM1JJ
RrmrF/rFkbSp/gTMbl7NfXLGazTAoNSuXYjDpqKu5Xf34A2Shh+Ehh7AEwjKE37d
PgXJV+w/+z8U2Rf3zktU7eS1MIFJcDKmFS34JYQGE3IovgMTXvwLEb3UnyG/TFRK
wAl5DH1ezW9ANmiNZmw7tkSUUf3aN827oQsVba8E0YCgef7OiPN8kLg8r1ejVqSa
OvUt75K1dbjjgLqHQimteUAQgR7t17UWvgdc7rqo5vSG28iG+mUChU4h1PIAVKeL
K0V2iErmLYOt3HBfB97jz1kK5hU8recSGcBjebvO4potsB6zAkTkKzy5bZxwiDYE
vMkmsVsJp4dPRP4e7kIfH55CIJSnfsGHDl6VWshLbIFrdzERd8AJV5LlMzSwRqXL
VyD6FakEscmyPuvSJVtjcU3n+e+yOm8dTeBsQ9sFXHim9qGV8ml1N3yzGLBiTS7q
UhfOKZQa0NQEtsOk/t8uqXaTFU5UMP9TfN9U6kapsgBoasAuypKppGHEMQ70eLVP
X3u9A4cO4ufU70trZvSM3Ago9cDGw8DYi9X/iCD6bsammZrmbp6QQ5mrl3bL8Ojh
cuyQ7pIVspg+G/GrKFGQJkVj8mTH1qORB69QNWNKxUNKW7vkn4UdK7Cusi4CL6Ne
DX+j5um3KqmgXx8QJiMUin1rEeUGSp0/lfbK95omTzIAgpXJbf12F6I90/G5U6ud
V5TXFtjQUB2d+oc0+ixZZv/DEbiPEcd6vSu7fleWW1UymJD+gcqEkWlvppGzedRj
QNis5BW0fuKNpqhZ+jvMXNN5M482mRxtBurURkeyYqeOaGHvZl+dhntXrXPJVwzv
ab2Syfhrafv9hFVf16xynz+4K5qHj8OWCN5vlYMrt5aopk7oylcNodFNapELxM2Q
IUp9Gw9rTgRWCYQWCKBEVpkDdHOcE7E3PxndkSHaIf8/UwKZydFeKAjHFoNad/Rg
UPMzTt81liLZN2LWJQWVWvvpDP5n6sx1C0bigZB2jUNqjmQPXzwCQqP+XdABroVY
v9sH3bxQ0cUdF0m37O9JcKf0ZmKLhsK3hHSjv24udfr7Ud80YBd8j32n1VViZZn7
pxjg6e+HZajX+NyRwULZigamDUp6HLBmBq5YhsOH4r5zI+1+FxZDApUNWCZC2Yml
+Oj52ZSEu6CuaFjotigJFlKGj1ki8vi/zKFXXRWqk90rAfeiWXTHXflaAS3x0Vs8
xpDDVvSfYYTGYlrOhS6qNZZz81k8Y/Oe7dztl8EGf1KE0k9skEbuw+3LOVIjrISk
MmL0/UoCv0sjlY9E+qfgbMqno8a0ph/ZNQp7ZJAFcR3w+oPq1oPzAvVddgSJdWX8
v0eiHdOtDf03AJ+tkXNZLdYr2D0Yp1uKa0WfGIxrZ80t6x9MgoXU85gVxkTooLNG
ZrcC8H+EuBBEfp6/BxESy+Ncjo5Fqt9BXi71seEqWZI9ajSJ629hwCv6juZLSIPU
skjyS5Cko285CMW25k1QNNE3j/HpHNP8i7sGiCU8xtVeHm9nwvltEk2Ks2ttewO4
oZdOixjc27Gt/xbJMi0G1+z/kMtaXDazsrTBtJfhaPxqBWPxsae11aK+yCa4+eTI
STDR2BRWy+bv+k8UO1eXqgQujpMeCgIiHoYNmpa3dXk3xP/WHFh3KkJAlFS/nSMz
UJa4WJGaRQDTklhsnHvxOjyKAHbhIeMF80z4Gi9FKHcN0kk18BqzZEXAm5s0uj3Y
jfWGHunuwdzaCQGEuB1EvUGVqCxX8TPzvApndh2OxzAT9ISo4JMagFhfqVTM4ZGY
NYLKKgUuBFWBtghi8fwuDIhkwTI1phiVjNzIc4uwh/J++icu+bK00VFcpXQdeLyo
ItyZiQqgV4DGHFHZL0NxNPs5AjLdRXdXgylkx/o5ONcYpE84w1V/FFCWDky+gxCV
NTgDWLXDuRns0C93pX1IxpoGVKz2aJPeRdnlf43A6RDQxA2YeJBK7YWt806JOjP9
Q1/ATy/lXDK+/l8oFT8OAXB/L+IhK1wqj73yaI8CQf9leepsf4w+75J2lInM6p3K
c/KOBIKXONDBotbhhbD8Wh1O8A0dWM5dPzC57bePq2fSC+oW6bPfBp17J+NLa+Yb
E+5U0kaYp8/39uIrhKs7KAtJpBex1y3rYMPgv6AERGWzPpdLF3FK+IXnBiiWO35D
aEnYOwT6kKbCLpT+Idx8KuRuL7BJAnAGD3k58WBHFM0W9Ae+jOjDUpVoIPvSZ5Jg
VAxRx3ScpNBbqO8JIxzPY+rMZNX5v7cR56SeJ7oXKIiNVZGKAdrAu/RFWnvA3elT
UMrh+9FZ3oa1FPYKNxKqbmXjZtk99Dw1qvwHHleNPayVisVwtrcCXaoRb0WENLDT
tkxhzhtu8PpyUapTvXWXCAzB0wb6uJolcLTmcSv7M+JQbB/PrezwpYOyNPYN7Z+h
BIB2PRT5agftVq58EjzHj8B+ho5MLNfMg/HiRAae27qGF6O9HAWgv1F9xy19E38D
C9/snEgrQ1YSgYICz0uZftUu+9hwwA+St/oHtzRxwNrku1NzoRbk8y5pCYXADTP8
6iBA5mDXdD7R4yhzDra8jrULg6zO4u39PlT/4SdQgmqIqJ4m/d/0WqZ0mErQ5sTz
DU5hXUI4k6WQiZUSvIVe9A6furLz/+kE3ZnyQLMSrGqGB+EsjFXbFwVVPCcsYzkJ
bDJsGPyd68k9DaNg/7NibZ5M/uMlb00UG9oUhQjecKbJCX7raI1wzSz5JgxJ7zWS
g2BVcEBcJv5rXg+7BnTzcf1DBEqNTFwQ8Jv22ShbV2OyJryiy/ufIKBzDaITgoy9
f49rogxVLqc1ynliKDoQibZYx/KLrr1rwNDhBs196Qnv4LYxSzoZuWn4xrhVuLj7
Fjc8Zur3vpDDZygYE18T4nDWXdYr56ApXi7JQOTCXS9WF4n7NEcQF0A5LofZPcYB
Em+wQUeVPNdTBrGuAgIDELhhqNHHVuIrzRiVq+RYgxBNQ314v6L2LF9wN/BAWcny
0H8A7na/zg6Dwq7GsAuMDoPJyvE9D5a/NuicrYqDOhcqcxeYYJxgcirJItAzoSqB
Xt+SZOQK2sFd1C3lIZtIRsyxeYYx5uLHQA38XJHyCrXJRceW9mxPoEQoZJmsGCcm
OvqY7PyGoUVZ+Ch1D3tJpyWZB/PhJ8zwnD2Kocfyu548zqVmZgW79Xl1CIziJeVg
GJ5Vu+gWbUgG1ZJVq3Q/e+5G0xbz8ykSjgavrO+YcypzmliKdjiMScuBO8tGkgL4
bdPnOWXCx4pETZ3uaErvz6JAakMcxjFRTLXlcpoJeR19pkJAVu2YtGTydFmF4UgP
OeL5ZnaRh6dlZfaPnechvtXji064HHHrYXqO42lRawIH8/ttvcLe6jkNKVb0iwAi
5ScaoS2w5SThpylgfxMn36ocETagVoS9/VB1JJCBswlGn0S01p68DWj40CsQ8Bcg
8t8vQroJf8GAoN5YKnvJcgG4YAxE8Ohp7NsI3kEu6f5po3g5a/DhLaeNdhT4KAmc
2FTY+tmN3cOCWfrYOIjoMW1+GNxOJBAbI2KpB2bQ1AQMIqDkQnoEOUjUfczE2vgQ
KgGiAWitwf1RzlV5i3LHqanwi6oGILGmi4DV43ukFMv5+2SkxdQLg1og8b62o/l2
c+M/HMAb/B5Y7ff5nbDgidxR9Nj2zblsO8GuZoyY2iXjDB1rklTpA9X2DnmjPCGS
+6qrLvzcJCaEmhWcGl5EutdkpyjxoXrxz4RgeY20fen0Daf+LlEux3wG7BHbMMkI
Uev0YN8kyodkPcW77zW0lL0M3y945xO+mkSx4KWjs5nIu33O+nfdi9xiuIIzaK3Q
/HCmUv8WVjiCqEPDKRn7zDeY8XcUZTKjnYPHrOgkBAsiTQ/dcD+xoX0LBlCpWmKr
NlyEYPXDdy99abopXdBUenrxdd78VbKqZH+9z3VEaUiJZs2LhGCLOKDvmn6E5dnx
KGLwl6Qu+XeE0tdDYo8cF9x46Se2kKaKDqiMB/3YaPZkp2/yc5ll+Jbt2HfQSOBB
OEr3gkXjyGxBfPUr+jX7IgW1G3jybKDKJHmwndSNHeqpYgxhCwRRJ57XGIWncf9H
R8mbBghP+OqkU9DpJUed5JjVEvvGmYg8fxZcTCHJT7uk8osf7k+nDjW4tQG1pdQW
C72MknRIZF1LkhGqIf0EsZUtwgKs6Ex2tbgNQXJ1NQeikd535gRPakbj80/XUwn0
bFAE2cCOVKuy7NABalHhrPPIy4Vu0bskg+FSgiL5UR4H5HKm9wWne6Idz9IgmFn5
2uXbPkQ3u5YN1MKdHrdSG4KNfGWvqZ4UGHJAz2SFNs1U+CRssE/Ojbni84ifYt3A
7tIeOuKiRRiwc3pkkSJu8DpPyqXB/vgiVhZSbtY52CJn9DwPgayMvdEQDpKXVjn0
qVTPr3PmOmfnPrM5oAboMWMZuAUopEr1FapPt3+55SRstEI+KfjqdHTGE0AzwbMz
UsQiYspsslJo+AXi5rPhkuyn+4t14tMWsWinMNgNMWwDrojErfv5HAHiehqFKiI4
eu7V0DEfKBLtIlbnDSIXI2wMUB+d1yqdMx2bL98veMTMuFxGLRlwIFRF8GJuDdF0
TZHGMPRPRcwEbBFHlQqxD7Spbi+yIJDYPdt+wLVGh1iEPS4K211ZhCXLBLpaIWuK
AEiB+ZjiIlWW6Kao/kNsQ6VNyfqMIV3IiedHdoW22foD8QpitFCMnZutePDtyItd
qap7zWVQdhWhWAzOP3JdOa0pmqJefPhEKdPidmBrgEkq7Zhc8VH4eew+VFSlLrOL
E2eFUbjRNAwa063BzQSS4/bu3irct8GGzN6qksoXAnWpu8r45Hpg2akQJfVmiXfy
bdHdob8cSFAueySco9kHeoXxT+EEYrpjjwCJP/FzFOEyeLie/gPMAcXw2GEAdoHX
Wd9Z4DCrS/F6WIINCBJONAFEKYjdj7wmAjFereJDY3eTOEOAMBgF4ecx998udVXf
Cz2zyUGCb1l1f14TXl0IYzCtFj3OijhXshPbzTmA5Mw6tdgcFOdQpLdXKbnBczu9
LQdBsB34yZu73cWgPlbsv7/ImtvafS4p8SRWrghuL+VQq5vKwSkyCj3JuDnf2rnN
LU3mX0VYUzhbdFVi8FU4ZRDvnFtxUKFj9p8uoIdTBj5PdBY7C+josUZTmI2hT6TG
NaEgni7vGQbfv0XHnznOuohAyN7hhWkM0wsgBkFVuia4WTkeq/sop6UBl7/IkF40
KY/W0ziVDwzF8Dd82jV60yOSFc4zsgUF/PdTPIC+OPUMArxAtkwOCh0eiVyCrwfr
quqOMPLXi/4z07k6NoVH9onbMEmA3Xn/28KWLNaZz4E43n3P63vkgXDAxCZ9xZl/
dQ9Dttbze5XcSPDdlgitekj0ug0zWdEN8CnOwHMjGddDqzM9s5NqDG0LpMkC8MbR
6LoNXggudSdgc6H1YGviAa+dZX328h/LwVtXmnnQMXd5ek4zHXExnkFPzZehrQ+G
RhPiH9EGFJIIVPHqO9ToELWOh6h3Rc5Y4dsB3eoJ4e6uTKYVDLSMHunUPhJNs/cF
hfKeTjWw4S4+wtWE9VlMOFDTtd6tBmcvI+Ml4jbdjJ7dJDw+0aCOMAybN78m4/Up
4sPdsL6ZkBDbADomxJ2RBKZwxx/eW7/Jsxh1SydCrIMJ42Oun1R5ZNCteeMdSB0/
vWbldFn79ZP5vskYzevinVxuh1ioRwM8klf+WaJQqC3TILPfz4uN/cz9/Aa8jWBO
ENLWe0W+fRZKrClp3l+I3X4fyEbtUrXDv3Km5FvtptRHZMyxxNGBa/nwP+eR7i/+
qGOIPhXzyDd42YFOOy3aZbZTyct2ZYHIF4SXqX3CqzsqqgCh4Se4bGFzRl2Kfi9i
LIIrgprCODF/g3xDDt7ShEpRBwp0/5lmUT88X93Jq1seAk/WZNI67PxkqmHS6Yzt
iTsi/z/fiH4Gym8H3Tax5NM5xeodfkDgeeaacZCO1DwvmdsXLK7VnSEceZX3VDGQ
lINIC6xJ3wWjK+qss1E2rXXbyG83B9jlcj0AgkX/iO5nGQ10JbNgGRFWY0n8Z/X9
oiLznftKY14bT9DKjcsJX9cHHjAlIHkgwWvRmFVHpsxL9m8DMnxzBivkPOMEgnpP
ieBSGpSXLndhRi34WpfJitv2j3pMQRteB4h0FALSIPvlFVI7Jh4HMPSLOvsSGLyr
igyTXGRJjhQ0uh5vY47eB5CKrbD3Timrk67YZugpXhClJ4hOCagcN4RiRPNra36m
cyPEa088FBzUVCkXbtn81P7h+oD4/8MeS8JpowuUmr44Oj2gt62cYe2w12cJLwsN
Pll4MxTTY5NSee3YwG4bvnlY5xjUapVolVzs5uub2eUotyFur0jUcAOXM3UGZ/vq
i3akkCyjJ7ux09yoT7Mf+UDwBnrFwPj2F+DDHvk+336f4mCQNfLaVwOmUH2QSdOQ
+cWllgOsaVqQczb2Yot7nkvYMsKypC5zi4wSVYI1eD24vGDUCHMt7f9izhO63/lc
hKwcvB6Er/LlQMOB1WHXrt1QF0CFKd4fzl2JzOi8/z2PGx/MkGywWoye/wWdvDRE
99NsJdo+wQoUTzOhcyBkTIuHAeCfYuJXbRHca3rBCaNy4o7uLUzXFfJV6IVDBO8q
N2qMvxggTXd5H+U2zFyHny52LWTGvtO1s1kL/BagQu5H5Vuz6F50aSgY6aTw2Kd4
2m2h82719Zz/AoR/hJsqHg/AZMFkPwNeDbkq9ymjFmwY5Lr3yTuUXh1xgKy1qPCa
oXVtt/Ffh8efgjcq1p2cdr2GUoA1o+bqY9Z3sOLIsWlePl9adG+QaiUp+Z/LWmcC
9rj5gYSqfoehNPFI15Wq5VH+N80MFKPNJ+uM2XHFffpywbJq6A50FNZXWZ63lTYz
8+t5L07k2cWvLw+QxGVLd0p1NTRZ89m7J3i2Iul8ZPj0MfDLqiCPsS5rbQZ6ivLp
0m6mkP5thGTN2wdwrAabsuumOcCj+/e0ifT5USkzq4avrNcvsaG/R+UejjaYcjIV
afTiZh0guzXzYegXYWpr2V/9ehOSmQDF43oinqE9abcHxMsCEd048akDw4OtdXYC
IDKbRUKYrPrm+PN70fsk2ezk0T/9/j/Mz1/bw5aYeqtY0xWaRWREsLP/JRJ1U09F
Wdfo2K2gyE+ffdsm1dDj6sTu9v5uYhlxOF0L6Jk02kdmTDwD81TvTVCWPlzKjgKC
xU6K/f/b5pX3+ab2Xp5Gk9Kg4+Wrc+aagYcScHLk5o8lTq5P3fcEA06ZNtoTG0qZ
vAnC/FwFtq/uymduEzbz2HqOhMt0fcmnb2O1ZALuB7tKC9moB+TA1E9Ltjd/Lo9o
bnVi7v0ORcCLtGNb1EJopcARIg+n+zydPlu2jSyO99RqH1t8qqG/rpT8SlnC/d90
bojehmqU66CKW2riDXz2Nsm5wxAC27aTiBfkxTUNq80aGZ/4Rg1AUOFS7xuBw6fg
aaplK8XOTCcOo45uqYvIkKxC86m60lU/2EBBj8rjAZlySej69+uuw/C3EPB7q7ti
G9dBeh44ZvQO8/04xRVw5rU0owA9Aa+pI/AiM2tef6TRcAnMUESsc5s5j/czy6EQ
q7VHu2vNu5vuD8HMlMb947KH9UUxqPKJ/noywKylqLmHBnRTuSSYlUeALdmzO3xS
aFvGT79nedrYG/2pxDR3rYoo1y1XxIkwPKNyTaA+7xTLDlZUUgIMhCcm2WPyvh69
7fqEY/NJAAkv/9m/Hyd0t8rF3R2wuy3w2xH7F4Vqv6KxhboFOvJnECbcAFkkZyaZ
MJtXNEW3/D6lDqI7XH+98dfBmJa/jyK1hCiLzzzHkfa3dtV2dUrjZz12vgQyV9jf
ptzNaqHnH57D2z5cGGFCo+QRNdkMDsu3HfBwPbElO/hhM9RhtYrjm1CNSRJGlk/3
ofum/jjcZ9N8xQfTZNZ+vQmQiaHMwc0Afhj7SlLqWCBaM8Oz/+TLE9UJmcd4eE80
j6lwdxhqoHo9mvteZsiODWpx+Owtt8845yuPo39/H/ZxnVKD/vNo6pr7vcxK4lS7
V/qlgcVnztQsUk4xvZra/kEW5QE1gv9gKTpqMavZ2oyYJyh36lTyAJ4oJkW6kuXC
FKtCnz4Shm92iaBWYf+nl904qfmiDqMfSmWgJzZjgQiguZNBou67kW9JgjZo94gZ
0/5VuD4tZeSdTQDyD1xmTsaX96Lr6yblOT+BU90Ihj+/n0qk6svfJiAVtV2orSkQ
BeG6nE3UrsiZevYRel1HBC2qb03VnzoHLth2OjAHvZOdxShYyRmJQkv/osL3/MYa
mWg8HdJfQ3i8JcQ+V7ddkWrJO4d6cg80mn8iXq9f03Sfi65miKCvs063iOHYdxnq
+61LahoXl1XpQxQv8uWBgpYr3op3pT74aQI8tKuIT6rMBoz5EgjCmzDfGQP9cGG6
cK5N9tvwDw6e9AG8rbXHqgCY+uNJzgD5sa/1qQoHVFxcb3df60+GsFsp8NniPIDq
E9Zz7NVi+ZB7qDIn9a7Sw6gi6lxMzFMA5JF57nqcRyuKm9Iff6fDZvQbTReA8N8v
FrSIz9fbnES7fxi0iTd8gxVtOtOYYwIgOy8ck1LDf5xm1CsJSEH8CM0EIscYA/W4
qvaZe94RIrfMHiwNTKrkQjfVgX8/sFmAIUDcnFZpTEaNUhASv+iJ6O2rw4gWwtP2
rWQ320h6rAXemVELIoiRmOsnBv4EwQzhcsLBKkr8iwFzqKiFgltR/31FFl1Qok4H
2Iej1SyuwYLKccZWR3HPNE8+YVl+AGsK9Ceb4FPYwckK8Yqsl8tjWisQC6clvRym
h1KhIPDlk7KGUSTTg46aYCjFSiDNEDcpPswRPwOaKy4ZKq2jvsYlEFLrP5LPQ+ID
wDZVYVXZxyLZXFL/HSAQnZem5l1dCAoe0mZdvH8B6GUpRjv70YkPMsHilZUm1uqw
lJg5TgtEZguYG9/gsojZzU54ZRGDzMY5DNWBEE+D7NTQLwqnfZlWTwr2cFJePKza
g6ALJKi3V/ZUDOVLR06quapajG7Ecgm1bhgTpHRWhxl9YRQKbHrRetRZMTtBw93x
S6j3kg7mTLIy2JDcl5oj8Kc8O8F0zkbE68xtcCOW74kffWQzhElfTaj9miCIkxaw
i/1DboNvsyRoK7/Zujdu8rMxkCF0M1z3AkUfy/yMl6nqEAC77EYFqkPq4TyIWbo5
37P1/ior3jtW/jRgUU8nDKl2/QNeO8dRbQ1rAUdiMcjXn9k7uAj+xtrCKQsssS22
TQk4ThYpN1xbFtjq3XEvq2sZW5ga3Lulh2YYX4kanmipjk067yw/x2x7bikvqTxQ
R/2SRuRI2+Es/7Wh423kDevqNn7VIIwIHJGeudobxiOVR8pd/dBqZEgC3EL+HopS
hZ5lGi8f/BBBxPjmkzhSd9wxyenXQHwwiioQwrL8DGoTv2B2kkHbLMxBb5tyxz4r
115wTob0HUsDOJEYTIKSW6sNSINi+ThkQnpBOLYFiJ07Rjd57eA6TCHq3t50JGVJ
Tn5vzZm91wKiS/x15guV3uraayYT9587xMCoYqHiTETywsQc+t+lUZ5SyBg3mWrq
JjADi2xT9bcIen/227pZhx7KKED+R9c/fwZUIgxFPM/vQel0pygeSzeI7Sg+FB6M
z/DWtjQaTza2Dlx/YW/Nf6aWfMHiImEuzIW/6svKKkuMwXzypF8B9fCc8kHnamW9
471nOd3Tf8Guz6GMF1J+Up2byoLp828FevVuwEXSmWInT/EDm0q7wUC6qClBaJiH
5cWeuHiGhftOfuVmK20VjF98MPvdJFs8i3V4joO4MiONJY+SAC9KwgKsRwV5x/G/
8GXocmbdGeKB0AOS3sc7gVTs04o6KfGuN2bsMnqucPbqb47GvzU/Sv9U49tsjA2X
e/hp2yT0YmXrabHIC679VD2KVX5tXsZ3ISPJpzaZJ9KKhVEFHfk6J1D1LVuRraXH
GmlNkYLvs3S4OV9m1HTyNtvCgnkjq4Qw5AX1ZxwaW9Rh9RILISw9G7iSFflkUTsK
bIYdIRdabTJxpQP4ZUtWpY2yHor69m7NEptt0MxtrjtIBxz2uZzfZRd1/qWjRqLP
+TH1w7Bq3iVzXcRYAAun1tgruPK5mLi6za/TloLsjk7iO4lFFX3RWkv7RthKA/2H
PfvWqNbniwWsDk30Nis//nRRFAQ5hOBfiZXR2tVYFCyHIHWPPzVFt+yj284pf6uE
K/SQdOGfc5GvVpXPpcQ+hATDucu4H3aVBkOLbg/TrwFd83SvLu0Ee7aHw8vxm8+T
BnwpLm1Iw8ozlx0hmZ4lgNRWRbci3ucjEPEVSuyjRZpZo5IMwPM/YmLVmx4/zr3r
Lx/yXVfQY/4qeCgqOEF57qZ+EsP+tt0DaHnCBEOND5eGRwPky4/+9fORETwZlMTF
Dfzu/S/8VGO4eIzYSrFRFLV9uSxyA3cJypzbBYZXyTVEAYzlUd7ou02nMyrq7Tjj
YiJ1PufBVWrV5oH8zfvo76qFuq1WMCaReFPRQPkuUxedciEhiK1jiDD/6QuNUyho
p1cDtV+c5yqvxNiM+I7VY2MzHKz2bkmL4p7v4OF1q4UXkAokrqDWaNwJcO+WVZKb
kUKorQlwu58n4l+PGWw+7JPMz7nimVAOcbFzfFfEHKEs8uiMX819ue8EWWB3DHyj
FauuKXb46rx2QLKCcSU471jrLLzNZzdMkCvD7h+DbxQqMu5kIW7NhwZXBGA0p/bq
QVctokS/rsBKeO52afseaCJJbqkGkJFP+POyf6w9LqF6rRhyWYaEo51LK/0ZLVan
PsndBosMdCksfiaz4fedQsMcVrmxu0EalmnOw1sSSWKAYZ9vaZ3L8rJZIf47lqjH
aaXBz7qvukIWxCFJKWqCsm9kmvLtCSO0wnSTBSictqBu115sHB8PRkSGuQwvXOiS
E7/SkmiY2+N+HW9HMeWB9va79h2Drc9kSJ0zhleh1s6WzbvsDQ6mihGhoy4yCaWo
QqWK4i8pz6ui2f8P4IygAdqySXq0lNY8RAuV/y7RDBri0L3HVjzW9z3iFnjJhp8F
pfDGoKmOYaRLtp9uSGDJZUBaVj5mzRzMjOrLfQS2Ngv9fK0HOh3ZTdufyIhWzRfr
zOarFNCi4/XMivPB3iS9bIqBl68TnsLifwsAVF7VttJKHl627RZhX5L1IctQeYbl
9LhJprl8U9XuelqrRYjq5bINg9bFBHJXcOq0jrRSg7JgDD8EfwlzfEP/8qLWiMCo
rXeT0z4PmG76Ug4vDj7wFcdLLj3gdsjZNXyme/D0V7EzghuzjYIsK30eWOOmdj4t
VzkgaPuS2IThMIwa2TnmECuHpaPW/J6SFZQXTS59IYsXqSFuQDiyWBAYIaaWtL/B
Faw4L9aHcEP55xI3HqgmgqYL/oIFZGh4QyOwWYpzcHl4g2cqaO3PbsX3y/rUl/oH
KgD0+wNZyDFiBbYMCNKFK5fYJz8K88bFWXqPhmZ1yx71YgdxnxJH938aVvzskx0h
AJMzr4IKymB3O/CBJ4szpwXnntGMqjcfqt0zal7aLviGxE6DAdH/RY1yE1Kx/42a
yJLleG/2yUpejKeb2ClMD8eVRUShLTLgllG2yrgBPEUl276GMj3R7Lt4ikDWmDS6
t3m8yN/Ak3Vb8EJ9bIRYMrRnItdrNquSoBHw4mKYbfA927yOm5flWJcUGPbfLNjz
xNFkGe3MhO68/XYfvKOJvVGDbQqlpXNOWZoLjbQCeHyThzNEmu4gXaCU27ZhBuUE
oB1oVr++k2hqNo9xjND8LliWTKYlZkwMA8hEyxYBNQqLKaYX1idqtLOZQUQEQLcA
BHE4jTP3G+HHQJeAG4Jsilks96ewkaneUQ79dckywaUfMhj/7Nm+Vgc/uskfk/cX
EwporyB0W35ZXXhwy6qARuGjTjH2grdV3RU+Egj1RKFF8U04i0gIEmYawXNw8IWm
u2WjzmL09nCY+MC+U8dgsntvd7oflqsQgIWF9aQzRxuLF1oOeiR9nkbs+cxcSg98
Fwx7JZnYiNnw6sqcSSu6KIb1ylPFhg9X4HKzDzWAJwxXA6CV6M6FJeYhz5+hi6ee
MoxcVrQac8rqrJAbldtZdXsMpi7UpMtJJW/W6l0MYyMlmwhybKfY3xLJpHpc15SZ
LAuHRUMmDMc9mFw9O2umVScmUjbNbAH8ekuz1AtgqZhjpscWOYb9SRQLrRIRsbc1
h4PPYsKJilMife5y9xC9o6pQSA3r394cE6ggVtHHwnyLjjnOtaoxQKcD9cWcdTGB
KFW8hNVtQlSBZrk5gJH7gTLrXq5sY7uWKUrbXNxHFjg5hbEvI/Mdpk0bCpDKH74N
oqciz6lUMMZOiPAVaEnwBhNRl/bQg2pdVGkh/xGZ898k/0v8HjT65d2h3utuBdq5
ikf/1Q3ovNj1s9jBjSmLMxkz6cYVAkvNWhH7AHPPdEU2Uuvfd90qgjdb8FndhCX9
JJttCTKOkkFCihCQ1oPQgrMpJw3WJqB5BKD7Xr6tyZ0cU6PQZkVak1fhCqB5k/qb
hyOsgHUovoxlel0DDNZAlU8SB/Bi2QB7pwjyay5Vdstp2ydyWHtbPsrFy+btj8aM
YPtDxlRurJnigJZwSVbPx8reO/9Qkpe3JBAG1uSQlbFh3/nSvk3GcrFirNIGBBS3
02M31flgeQsQo4g2teax/lNRjeomeCjdVWYir0Eg3ch5RmjmgvXuXEDVDZT/eIgn
VK0Rz5FDpXk34HhnDPvWy+sVgjUJObRvuG1PN2yGYMARn7WWiQzI4A8slkYJVxpN
nvx/8m/j8iI3k2qTjmm7HuO0ICUKXujBdGTbUUSViw1lnG8G4uTZQsXckU0NJrPm
AXCi5AKqg+k0CTwSBORuzGmVu1mFdSEQWPnGQLc3FBxlGjQYvlKta4c6oO3l6IsR
YRJOu7WOlsgZKxJRgEIZTdIFdk7Qln+F9vs/1+RRW0zUf/wcg1jjMHArab5bgDUb
vrikLje26MkOv/trYg0KmD1vBy1F38itzHJjDH0W0zLJM8CaJ4c6phdaILPvURWS
DSDpTeQSc7lsi0h63tIZ5gxQM4vatUxOoUlSwCMpdqE+VnNy1mXSObpTHRG1fyeD
I+zcY1jxSr7fY1omzwxy+piRdIV+WEKFyEts9uw0/tH3TPzUIeEfPVJh31yeh0oR
THUmuPnukzjSxPI0G9cxGREdZpro3ln8oLnCWInxaQryU41/YX0jwFSNLtiesv1w
4zEbiiyJt+hrU6MNB8HGSEQdpCxbRibHKQNJk7PNmUCh7Am83HaSJWqtZvRAo0VL
VWaNvJjDjWQT+xmVEFqQ5MokH+dg4S+MF0kEl4OZNpFWPIF/WxHzKZQwKEraaxu4
my8JtIPvtaRkPJlDlNudMgfBuL6q01KsABy19MgGL0Vc95FOpPZ9z2BRNVDLUPvC
iLD2wIKTyx6dl1e4ESGHSPgHiwBAM452nAGndZzsNEhxzbfUn32N4tT3+vFBWwgs
m/IjrIjg5OIcALvgIjHNPPs52WnMAY/pV7NnU2L9oD04wR/lYmO015XAZmBhLQfh
2kFy6UsvYJtZ7/xbSVEWYu5ZxYsNFy3x1BRaYzJvlPZKAXvFMxvG+/+YjEsKWdGH
tF5n7BOIItQH1BRKdvdC2oxbHKldKLfm8kEs0SfqpIRYZwhjdn6XR/m6gNoI40bt
ZNDhaRUKICVrimYwLYvnebJZZfrPol4gLx4OOZF1j1RTEbvXeum+pnuoQqxiQ4v1
5T835IN4XhYznAZcOsl6LuZnDlXheCogEKjOpk/OS233zVIhspSxPsOO2ohS3bOT
p4uagKXuUAAZ+q876/VRiptvBjAoTAivx52zo7WaeEW+lJTXakpf/s1vYqhBInTz
nDEDO7oCkrVe4D/iCV6LUSttqtEosYNBg6HGYE8YmIBj4Y5+vdhgX1Xs6F0F9WEa
V0VRHlR/qbMWOhZoDXIooopgA7SYOXrrbAsVS9U57GGdhdKj8O0ME8tgu1+tbXer
sq0L9OfhUN5EdjeXSpVwOtbcTukRQk2RElkjdQp9of7pVOOcgC+FuXLNpzzmpRJX
KBxJWL1dDMXX+NVyu40UXhDU8OcCs8VKn7+WNFWXIy2tMfmAONQQO//NUpw/kZq3
J3YSl3n7DJ9PD9DutB2a9E3GoS6ukbflnjLGkSeQdtngFXaqRoIPrLkImhj7E63+
f/ejcVwNJkVKhB85NFfsQPT8IKDx5gR1pMeBQQlcFQv3okEWiLJMx/i1+2ePEYeZ
5k7tMEC5qlm101UAxQoBvNrjv/2ixHgOGFb1O9lpxyZHJKOMvJfDy0buIHtJ/F6o
ciIEYSvLFAs4xyI7IwNoEzq9qp0ckLUfUhfkydYnQnLNGa9l0D9SQ/+dsmLqk/kf
JXssqyk4QntyqenaHxlZRe/U626G5ViIV/Px/cwmyBjeaEoUPhjGJRo5GN2hVMRF
TXkyRPE2s8i2i95Nm7nAi6P+2tjnXPbCo0qsCXmRZqsoy/ly6Qk1q+eIN5dVq2M0
Nz3ZXHwB5tCZJqmaJSEI8m2QSubCNRTr5vjkxBUvDL8iw/YmzjCfZwumFqkl2ThY
FksYdIXZWqIjSLG1HRwcNdTJVa4uWZkc46huKt7wdNvr4FduOlhgWMCklRPN2jHU
9idL3iE/6W/JPCS/Q+mTRQwk9C+HQICXKzPOGozMnviOeYI5R5EvNXnyFu80GyXm
7p2sF/pPeYtxAHCItMgzL/NnxdHEkWd57rQlhfrEALv8Ynk/8x/2SuMHexFaSaGb
rFLSpIvh6s6z8LD6VDeURUXof2HJXyCt53FktGTMNy3wRkhddUCKkzDyOjzOAruQ
+cDXYYFUoemHIGyriEt7bXGmbJe9amYZI24YWCbAQ70UmEOadq+zukHxsgefFyjJ
rvILKqsSP6534YObZ7Z98+PaYGA17l9d0D9I2fudD4BkzES6Pq9NKIyCL5+lS4Kz
mJY91ulw50Rowu8Ggv2nn1wwMaYConqLXgbSVqyRi0WkMD4rzyiDI9nETSgLnqC5
Rx+sg9Lvb919wRL341oQk/PQ3tTSL/e7lWfh1oi0Azp3QpgCv7GLaRZixOhHDdxg
i9rnbAIkXFDPGg8OoIFBh6IDUyvATYEVhPGQVlU7H8F+kHK0Eu9ri0nSVEJ1egsa
Argwsip91FPIEBhlLsd78H9by2bzEISNAkp88K7AIs+VpRSrww9zzX6X6J5kQRC+
AkjmuDnsBJtmQfNDamrGkzD9JGME29T3XTJ0rRVZZK2KPEwV+rPlAUTRKlHjcqzv
p9b5TliuN4ySeqlh0mlU4Fvhm7R9jmdrQqgEIt51NMnd04auKWXO7oS7uFhEZ6dL
OJjaqoqOQaE0QKxqIWj5GEApSkpjLqiFlrz6o/C9FoD1nzZVVH2nKO1fZLS4rRoh
wE0WGPS+B9J9FDJenOkGq/wsVStOnzUuKZ876qx7O2+hHkcq4ijyHqJWzLfiwsxm
toasHN1KgIPjh/XWssTzrIvf8/HPRo6LOLFCXIAMmCFDMhycrW5TNkntjXGuhOmQ
d1CUGldz23kk1C7hpxvTuyhEptS5OOkXcRjTgcAcNPYj3+cghwmfwww5YkDzuUNR
+LUagfaWsnNbsRyUR74g/og/T/kz0o3XkAOkvPqCZ8RcvhBzT1D+UKnWkF4a5rl1
bKU2dEEc1YWCyRJL9ZyGkQOJ9oscopGJ/lI8Rve4LWnZix7LFFw14BKvh5qZpKTA
cEPywyXr9nHHPNI9L6CHzbDALdK3AVbp/t2QuE4qe62lpDRPBoO2ix0ZcvkKI8uY
++agTay2/+Mu//Rj0VBJyYCqsEY96s4xpYyDbKr8v/4WbNiDLtbIpb2E4iTK3w7y
6a2rZEw5Gr6bgTfflfKATVKjw5GVqjNZdYzHq2AexMYaZr056BfZ1EPWZmGHcyFe
Msjtj8QrKsFoWbsE6PzoYuUK8BBdxOYLvvMVFpZrqOvzhTVwwAp6sHUL4XiZy2HS
lbw9Iz4cHe+wlJtBntPRx7/weS9AiWAKLcg/w9xb8TLKgPrj1oc6zzWy86klCohA
vQ5HWmo974stsz56u6Tk99082EnN41VapbdVOohIaz4C/8l4CLMx+DmtamjydUv/
dK9jqv39EJHU7vqHaPMQs7IXKM1V+Rby6OPcDfvnIVv5OHHgzpfqF2dp5Ri5AFJW
hYFRcv0hvIi/8FHHXQGT+SVDR7gmr8gXxKoP4bzYvAZeZknKPUJUQ7aakQy5NWoL
lFeLtdpJbXXywRWvzB2fxstEOJeH2w/5BIKOlWRdBAEYhAaP53kJH2qfCNs5jGOY
vAL/lDBmR5VJX7iV7DJy8TUMHP2irsgxlziBhwEBfPNmX120NYamaK6lt/y8ctRH
TdXiKftBxjucLlPEMB2p1t887iQiyN5wtkm9Hq3PhlI78DPbKWqaiq6elx67UbYW
T9bwKHRpghxUu+58lzBqz+1WTABMXD0wvSI0e3RFf2Xu+7o0r2jqbl6MUAoEWNBd
3sz6xP9bu878mZgzNI4+vPRWyEIIs6cvrdStukGFxT2yxI+y3kWfmXZWndELMPBA
GqWQx9WFYlRqQE7kLchiRMl5DCYIiJL/Q+BfSBqnIAHLcS+vuNl3TYAUeH0WhT7W
hKIfsqN9KDFIPS5cR46uU8i/ESSiaTbw0cEfAmUSazTBFNB78txsqo/DAs3hfLpv
/mRCLOE0FJ7NBMmGIEuluDq9eaJYbI1T/S9dyYSWg2FUP+kBBLTjvKdIzjGzvMZU
GxObHE0kFIFnk8ACwH9NiST3KikX0lQzj141bDFRaKfIGkK6iEjJXbgz1Judd2wd
zK8hHqgdc1pLm67hXExnbylJDNl183w6aHf9yEryQofcwg36V+ShhFppztmbqjAE
IaVltUyO680sErEKuc8sRJpoi+b1uQngwEBS71U2SGV6hhbZldIhtG42196Ik/kv
BaKKulXgGVSODbu88lRWGe2Y59OP83wrUM0PAIeE4dS7tycNOWEymJimIGVO7JJn
K8zbftSPB3b5yfTZNZFWWLc3PcjOkZFyY/puxGg2eS9lXdvo1rbaGJIoUWaH+asA
HuxRpOt04Kv0431jY3P0H8Jb1j0SM0P+piRtXT+a4AKZTwPgEnIpb3i5XdMtNT3M
Xy3Z5I93GhpPlzQjmxIwpYcagCMVw2AMxTA3P1MDmgYRWIBokNJ2X4FgJXY0/Dr+
AivYNtngxOTlDKb3sdUleT+zMfzR0j34W7sInbesHOqHJjadLToDtL506Ns4ZhDz
PWo/XL5qfjDtAJ02sPCQ1EftR8LrZmR2i/GWp664gQOX75yUHXQnaknxpYaZJLo/
kjBHRUWxSgLafFlVt/s2Pf4EPWC5iL7x4u5VghyjQvmwL9yD8fBwKNELUcB7OWoM
CcigTMAIthkyApi7QwRDqQvJ4F8P/Gh0fO+EdKwHoVp2EZ1E749P0Uwe1MK28zFK
g+0vPEfhOpZoPVHbH9mAMxr6W8DJeBiPDA1/MKnK/mTRP3Yq1J4tZqOJG05Yof5j
rNv+JxTR+Q0BIXN3vcy/1/0CDGl1XCFm6eYr27pgO5c+AHQ+6IK37WXecSCDjpiQ
AE3aY7DwYt1Apf8THk+9+I+skwaRAKcjVSNvhlaB7SZZvyWpxTmuzsir+nKR/l56
qv9gsBsVmXW7mzbqt523lGDI88QjoC7BuIJ0Wo9sCE4ZA8QjH9+jIyjINxA4s6Ri
OtbrSQPlCXQFGNqsx/dZo543kGu/PoZLQp/oZ+4aRfOh4djXyXH7moi2NWupQeAx
37gek3Jf0o3K4qPxmhTIuhj6NgqUjSJaTmw86fdvlyoOB8mwUCU2gqE5f1gOWqno
YFpQ2BkRGzb2FC4ntBpHFPKyKcQjTBjk730oKFfJtu624td+12fBc8fh7KgxdsEv
bkbaBtqyBi3fP/6lWwt/SqKaqL6+WZyi1zoOFbL2Jp8iwbs2VcGuVe4bCKx3aPIR
5xqpeI5tomSoILBnFEdWuwLAMnm0/6z0yvGLKTNj6zz4Stn3GS2/0PCPUSjufW5P
u7ctEs9jL8LcCgbEutWlHfiQfNdcBSBxhz9C2DSEMAEHuQwCwPEffx1FTvHFU2AF
Qn2aSb1Ca6TIMeEJ1Sw3qlwVf9j4bATiBoUVHtba7aDzjvCvD0fZGQATGvazOLH6
MuBYhyu1TVawkUs8taYxNDVN4sTOR8jJhiWtePOzoWnOsBkvHim3JdayBN1lfUQF
hKNdysYMPVYl/Ipz/Bb07jSIbi8qdIAAF30cFkPQETGQVDsJrvrvv6oNY3pF3i4x
i1wIsT3SX1nsfp2yJ1OJVl1kFbIRKFc6IbuOGN03DY3hRkbumZVJmPWmjDhXMKI7
78qxHtBrQvJdaOi2vFe6nKhKOJpXQbqxiZZOO3NSoo+/lp4QOhsPsqXlZZ3fSlfq
T/CYqAqqwOZVgNoojdkzR930/qsr2amnnpzpLqC2N8LIlwlHFZxp8dv6fpy8OEW1
OFY0TUZL8PegcNUO0i2DGe7m5MFDvbaRP7cmW/dHQ1zf+yCHWlkpwUiRNxsZb9nm
9fIwqLtJZ2555Wevlunxo9Gc16knhyHhIZI9O88Y9BkX3Z2dIPyhtpQklMC8f99r
6iyrXzTBBM4IHoKo2em5ZnW2AXn3fRtbfiLQYSq4OI0xfo9dOIO6dpx/sJ8TVUz9
6hhRTmSYBG/K2IV0wNUyk9aZBrmwTbJz1IBMyf66Rdzr8QiyYgDEcRZeskdotVPN
EtdTX4sqLuKx89dqAAGyUFoB18+wNc0EDQGAyVvvbhQTemv8ju5CIRGwwlL2dEYZ
fPuoJbaqCuLVq2CCtRX/cnVL0YzA+HI1Hve4JQYg7QkbzwtoIX/IxkKKPP6p7ZS2
Fh8DjGbgxkyH/XjnjMF17u5W+WruPgzQ+HRCQfnmqiWHFkuL/XylJWfeeaEFOAWA
eX85YhquO5BxgcjO8+ZE4n9p2YZE8Y0mW0bzLArjE7lcY2uq3LfG2fwg4GEwfBcf
Klj/aXq4o9WDAf3C7lXKK1qORB5yYicX+IldQT5PK9NHIvLlDN5aJPNd9jIV71+D
zvADGlBbwoZBdRCgTT8neVMjVR0ahWkIRkpzSl8bG0FZjbnWW5Ug5Ff44LCHxYEi
2ntoKiomwTV26l9zQGa0zQYlUio/PAq2tSVK1NTORphZ9/3/XOZjrvXEniMUXPwi
Y6cWJUSqlT+eJVKpGMdMe83D6FZKmek6wWhGO+Veh6x6dWjvwsypeeNrBmuT/gMA
JojvdtO7IEwbKVt0cRWW9yh9uNKXcZVBZIizl/xQL4HnUO42+G4dCCO56Ul382ye
NRibFOyawQKtYkx3XciwFxN+wQpiAbuQFITasIJoFmfiq0Sb8kcM9vmZpEFZaJPX
fuJMZgueem1QQwf5VBYxAjkDalrlTRKxLYg9Eg28n2P8Xk0QMgVUx7OakmIUEEdA
gi5VfIM5FLQ0hJGYxCy9PNOuX3N0iI656ir9dOxdM5Kz3vfbN1kP4vt6VM1YiACr
ttMLzRrUgfewOGBqLUZr2pNsVQppa8pz3tvSeoHKb8/3Ne9cIhnQ38/2iV5gUquI
aeQp8ViuWC4+qMiovAJjyzQkgsvfn0c8W1/DbnESkndiZPdxOX0kYRuDPzWWHYXm
zUStT1V7FidKMFrsPUtP+hBm/e4p3Pm+uP7PIdZXQKM/s2ww6jEsTl053I0xusAP
eaaKVu0Me6UuX4XXhTeoBiiBN5D9C9mpfLIogpAPn/ue/pNXPUDhyF/ACXh6bDZX
ylZRrhaoTVvhMsZWTjfzFHphFKiCU9SB1tsOmJIlaqQgRmoFQsd6iwGsPkmxLaFf
qcMIxeb9YJDdugepCRCfLjXy3gnSEfCBH2QFPO1vcKnMVXq0SvEIKXVHYpPiswMp
Y3nFXCvnlEWs0ThOL+cCXTAzZW68RV9q5X5nqUKQ6Rrv+VlrNyTOH0Ozs1Op9esd
smEsdF/2olX7/EHt/bbbl86dWqUzpGv9NBfVDYv0Cl9yi0AziSD++XWMSLDVLi8m
w1UXxZXhUAAjjKmFdh6cIEXx6wmefjZCXIs4rTbkjrLsysXHeCTbSDMOOKqhpLJr
uuN3dKt7PWXEhqnii2r+3ObqS1TxJ4oSAZ4do9rtHKBk2bmSday1UKuzEBIgEfxc
j3wRxH7Cj1hcvwrNJiLhNh72Znm8xWHkYn+ALnIC2s7iCO4LH0ryd6zb94Mw1tao
0JEA6DnU5J+VGj8D4D4tcr/CqOZKCS0do+/JZjTPlU4/yPretzFJ9GNdx30JYO4B
zkH9DHTIL3HlNmCSopTGhQlqYb4Tdl4qPUEBMGpPXHw7+0vsyegxKi/aPN204afc
F+wX5qr58009aA8D7jhMwPEkN91DaAeLt69lrwLC+j4sS9beNhje6G4XKQ3yI2IZ
7rPHtn79SLNvSt2A79o7OuTuD7XOhooNDdz1cTWLjUMhVh4B6OgfZY89ifcudhMb
IXxhZ+wP+T9j50rh/uxiDmiSU33GjHAg9K86NlnR9s6CxEt6N3E1OK0ihWN/R5fE
bp+IT/yMPG/KxrkrUrNG6M4NSjqXmLVP155FRVuEp3s4g7hQKEzlPwTXjpBsiVUN
bl054lkxKp2KLHs+9Aiwozffzhqi+v/B2GwojqAt0siYy1KAi9ds0/6HYcEAjobu
GV0OlaGMBW6oVhiyolpxDrGcvlGDeou3qBdqVLAT6ZYeNTevb50sq/PJsMy9Bhrh
nqitMoVBHnyfIwgrtk6IvQSJ4Qj+86U6dOuBvtP7nq7lYpBYR74MaOJ+JC06lWxB
wcqg7PSX/XM96VdlttAsqWAIFHvBZ8iAkYb0rvSajWQFVB1j7A8JVMquoOytCN2s
nH5wYq84F1QO3jbNEERuY9zZhDXEQ2C2HEKM/LE+sxEXCPxFR1wgad3B22k3BclW
dw+nnTDskxUNBy+aaZh0q5BomXuYt/dpv/70dez4pV8jin3YMT7Y60CRC9mt8JUH
mBOZuBB2JDA49Gp1D4nboTtDQyOTfLJ0AhHD/rVSKcaUptQVrZWxUe6cqnlRyhD4
iS62NU8CbkKggZgGddMVg3RFbpNvqKwVuU84/BL9Rlv6rokgYX0KIbM6QZUXH3S1
tr5mQB59tp+L3pwTO+LPsXclhNgtLKvHDOim9rSYoiFNTxZMhKyQfwDrxk65vmB6
UwHp7GOzbYTc4P5U/A74cJOzqyEygImp4zJqqKWNoSaeG2Wuoq5vqfj43K+1Ydr7
8gip/OSzjhGyZh0lAWsUGC2RjhyOWp1s0OayrurSNrXjbsLB2+ZdUxZlI4WtF7pk
ykiYta24vPHl8sq8nuh4cYZQ3PYJ0TKtUPX794FMAGOOESnGbF4iKMkIm/Aw5KsF
yXUybW60+dVeQndovMw3hOXjt6i9b+EWG5OOqXuL60ocFjbiK1cP4NrPWqF2yfEL
UD94At/UWycFKb/jAz7EMJqr/BQciIL/oY0G/SzrwP2DDCkW3iTb93qfLT/jZs4A
AYZ9DbwvOotVNGhho9yRDHbO+l2jjKOspo3gpsCUVwEWBMDretThn9SC2XFFAeyz
t0sFbz+uR82reiaCFRRZ/JPjHy2RwzU8mgBSA2lVMpmaa7d8wawUZMyAVT5T+Qvi
tiLOuV2EwGCg4d1FbIujHFeMa8Wn4texazDXh8msqyDBDCsqX36FQr4qesUR5t4U
qxPY/RmNVs1yba6+nh6ly3rIUseKOZ8ZZ/pWaz0EBwAUlohg/bdmA/Qg6Z91diug
6XDY9e4gJoAPr+or3eU6WEdvI3hke9+pN0E0ZTCCj5fOoq1sPfuPG9No7Lr2IOCV
WvWxlVWcciM7EpTfDBUCe0yXCQ6i3rfIsV0QPxcgDusY3xbZjDBvcv0wp1lHm7F6
RDtd+PIZwFOvX62nvbuN67M8uv6mnZwPUo4lZFuDUW8KXvZixhqHQpl0WmEf0JLU
dvamVFbxlvpw0Z7uf75+Zo9JhO65hHPrZaTqOi+1SkKZTohAsicLf2LFkDufikqz
x+xgDafDn1Rz23IbTlUph/+eJZBvujtabJFlCzH8j1VaH7D9A4UDHI52/0MWLJ4Y
eLufftoIoUB5Mnkl6QT9pHzxUsz2BNtLMokmjmBs7Vpc9Yp8WQry/OPfNrrYq5sX
edfKEUNLWFkzL/4Zbf+FUxxe5YPzxVqHMWsBhVQYqQrwIjzGH4j3C8TCKr3ODcNk
WFOXdxKeIwDWZn3Ptj4mmeO8O3obdT5LRPZdy1x1ERjYFRt0f/y8LtWgRNQgH/u/
2hAOmCMWs9Mqpjzp37nXK7HUyNL1JoLf3W+fWjoaqJxNhXOG3WFs9Z8v1uKSopJX
NK+4AMciNCSEoiTT1Ib1mvaRlYDLgDaQQygW7aA7/jvRHpMjV9WnzxjLvvmck0aX
QLBFD72oL2s68LukZITJl87JAQeNfC8ZVWIbNIyq+ZqK6UhfM7tUhx39J3UvrPJQ
GzvaxBshnwP2UVw5Ir9GZ8eQ5Uy4bDtEfEGuDFj5KfgW8jMiaksjhfxMpRt1plNI
D/A6JTOyawhSVIiiBkYzSpHCFbIHE0SyPnA79kPmJtyiTHtx3uqXkjK0d61goY49
kvrKW5/NuVKIOZUxjL3jvthZMMvICyuYrggJyFXeRI/YKcpdjW/RyVguqF470y5i
hVzHhwcLwzCPY1tFbgD0xbcfW0J2zMDLakqFUeYZZBln6i0xpeF9F+KpjDI0kfPI
duyReOZVwk/Z2KfzDmdTan0Dt6ZzMgwZmjvp3wNizQnHE6qil7DGyXGPyqTH3boC
kYPBPsLnVUYNGZQs2nt6++DBY50Nnvf6VQIKHL6DRNR1ViX0PPIR/eMCbwd5WgrB
xsKNil+O+5HsCwpYuyWAyRtlsFRtwOB0HpD/x5GK8XK33RrZ+PWbcqfOcRhzlgV9
n2uwuHrKN7LP7El4RLCgeybBN2pacaMC8r6McySYz9OVMccLcX9oicjUrFUMEFGB
Jkn6ewuGIAaIB+tdFF+b6DX/yQLZ+kVKzz0CvUK8Cnr+SNe+NVfreZmWzzyKIZFH
hZ7DUNpZlCPRP99glO46wOqdHogg0gPAVy7q52dGyP6QcU4D4A8AEFDrhSo1X+Aj
iY8KfJa5pGyJ2Zf1mhCELKCFglWjkhKDRq8qwtA8YlJ0bE3nO+oVVvdtvYy7wEA9
OXgl1nIzjF6VDFfO3DvofUn/NuftXmR2HKGrt9X7NJT6srsZ2SOZdcAYrKDD4YIo
NzPK8Ch1V+R6NtC3CWLNtuBHdwmqbbn18gWja3iZ9hKl9TVw4OJgyHPwahmWvain
YGq2k3KxxRDrWRHoioi8RrvWX7rA/wcuKUeCWhsq/b4uLG7WR9023IsCrQ9Bj8pJ
niZkVs4XPNLLyC/4LubCopDLqvnwAJb5IaK3ASEaKs6UW/6gr9UJAI3X+WvNYRaQ
0rJgUul76MwFpqmDq4wJDWyyAKTuQMb08kPLQTJlYVwR8fOQ4JTqVvT4PnLrUh/l
1VeQl7UxIEQzbr8g4IVxYyE+BULi6HH37n/HN90ufk/wXHbuIY1xrvtf65fAOWrk
uCZXjQsLifhEUVdie7eyyA1HE9LADPRVPXUvNtmpp6TQPtp82dBlcYQzHyOM75I7
d4KvSJ5Ngcdro+XZVO6mLJ6oMAIXT3p7m2EXXhOWEyw+tpLykugP12TzN0PpEC1E
cDbOlzwx5XJgOLNZLAzsYR0r1k5BDHtZiw4x8RjlvpZUfRfe//keLNgeATgzoXxT
jJJqAQ5AJZq9ZY9EE0v1ZJ7+Kn1zWGhOWhKRaC/Qs7k7i9fSIDcDNwjB4euBz8yd
vJh8LXs4odo8iDcQsY/X6kw8tC7XNufsZeFE12fD5OJHqsfLEt0Bet1wv45DdURz
oR3g7WTBBwNjJdi48kpH81OhXdgy/e8UUt5nr3ewt3O22xidqV20/xDySbrlOskw
9O6q8U9usFcOHaJmEJ2RS3fFFoaLI6kX8/d1wvzB7BqbL/qQZor3iGjsdfF2MKVH
kYJIFeIxF1OXWarxUWnt50XYvp7/yS6l2lymEjoOzcf2DBeXi38OuC/PGx0gS4S/
270iSh+q5riA0SdvavJMSP9sMxW0sYS6t31+Wh02GAaSwoZZi9AD1Q928SPA8Knw
vQ9cZvhRpR8EmxIVVCJEL05lPK5A/U0rtGkq+iI7AhT1+dHnQR9rxcyZL22FJ9NR
oWCKO9hGmmzAPdUjZCn03pO/6bwuwVoI4YsWIS1DP4QkLqv6CMVMCm9nPlU6ifzv
QrPnQih9qZUPyzoo/90v4vhjzI7fvvZbZbxjiAWv+mbYnxKlXueu2Zqay8QKg3hI
4Dp3ITJQ/BIVVA/aUIy2HCaBtmWvqNA1nXJYp9XLMXDg1QOcE247CRrcWe/LXR9n
QHjy7Kql9KWK+QmLhLdk6J1+K8fQTk4pXHI6LxyZXX2T8J0RpObfN/ZAdJ/5ZAap
AyCpfE2yeLo3x0guoc85kjN/nyN+T2/wX27ZZijYC1H0vmdA3gMV8CB4ZieQ12Bo
N3I1p3cpl6+5fiKsxoX9Ico4ULjdQYzfdmMzIHAFycnHS2+nbKIRgyMtrJpUn9OT
Dz/b7iNcvdPQI9wRt64nXC/L78RoNcPu+aRS5gbDupfY6h0V/rUuiGPCQ6O3URHb
KntjomltZWmMLCbyNri3bil0d71AVQCGlcbV6kx9IaU6V6YI03w+kyig+odsWk02
g5J5KHIPGhsCtW6gu585DFXYz1e9lA4YatAZuYetLmhtwKehW90Cxu/nFeqzvJfl
TP/FMI85lYQc7myOH/fjPQ8VuhmBSXLZSyr+WZtWDutg1l4wFYSQ/lc4mjtwL1ES
DIpSgb3IgZW1rHtmqF3GlUfKlq1vZJMCFm3xWtUQdEXkhQ5g/+h3+WAT3CsmLvl3
nU3IgY59PCGsHaatD+zV2sruuIe/47vDmzQTu/3+QNNH0H/0bcS1hcYMELZI0XRK
cQ3PZ0POTjTZUNxh95t3zJ1Qx3ANAXzDEs8TVp0ishP25Ai6QZxW20q2RIMT4dZp
8ZCF5kv4WXRU/wVwTi/fO+V5uSCCwC8FlxbOTUZRSMAV4JvtGlwCNJYQT+pYbSDR
j9Ff9SUozt3nuo+Bc3gEOZ9IfLEo1gAc/5EXj/RsF+YE4wCU3HOdLEYjkB9hDiYr
tI3naTQgrROqj0KVppFc8Kv+Xux4EUn9YwlswlyU/Pe31gxl9a6t/0ilgH+oIu2P
rqFWiIaCl5R/kH5UReojlVfGQXllhDpsUdWz3Ba9nIS0dtgb0OKDPbwrh70NrtD4
kFcaxYLv5bN8Ge5fJLm9UY3df8+FEqKW6nexBS2Os2lJrLwKAV3X5u17WNdaGY8N
r4BQRBUhJMXLeoreIKMG9NQHPbw8YSKYQnUiOlyf3ls22FFnpCGXJnFbiACcC4XT
FOGuWj3b7xkSM4ImUAbIBxEl498cnOztjvvGU9BWF8uJ2LxLqrG/AbnwIwRmKM7/
gwxMOk5GUp/LrK1UoV44bCKqis0jwKQl7of6+DGSCX/FVcIw9CcK4Vg9pXYYFemS
T+tX2YJouQFq9b46xedN3C/1VJa1r5DyTtSvvjhA696mBKUeHmEUvjHwBI2MIqT/
IRMTDmXpASZFd9PxtFu6ax2Obnumf/6EY3ePdLAlnI/aZrzTZWmGz0boBIu/3hnY
8qvx41ZWh63gy/0q/ZKTpmjZN0Gf9EHAiH5FTh2i87/CAPDcNIbdKPjPIM64Pijj
nFmlIKt3FO5j6gkB6dZCTAvgItRj3PMNflSzCuzlmySSEdWAh6WWuJIyCSN/wx5s
jlHL6HbxqQUyfKVUEMZzfSLkrprWYDahwsNAkUXZ855laqp9IKp59Vohe1eLbz5y
KNGHSUkihSmCJqaMyBTvhmZ5/dQCfGgr/hei8YyhGFdT9Pi4KXl9zE4F4Ci+Tka5
YbqFQsKd1eOOs5dJX3C0RIIMsWC9IoSQcX3dtexFjd6DvYah1gB2Vxgtqp5GzU++
SukLYGUOHQ46T5Pd8gsQGLll4cttRbAAUW0rFlKx4OkCCGCgbd4Ch5BK4IwYMhfI
1mFyLPgVb6aNmY77YBcWDLFbNUnoytQ1HlGAdsKzzSzm4Sk+5N6AMIt/6GGzttwT
pDOXpOl+c6sKwgWJBO8qD+KFFWvg6wMtzqLoFGPmC7PHwrae/vyoL7eE/qNnLRn2
h9GtiiieY7FhOGl9MCHu6DEYbnXrcuONofINWoHIElRRdwpEjSxdYtCXFGLzIMRh
COrCFaHCiDnKrya6PTbsgL28QpAn0Ymjb998kJoJ0oUsSFq88FxbEquPozi9g3/T
CBXkzYSL6i2HsQA8SLXTSsLlXbMV0G30G4+cAHI8SsZvnwUXqtag6ASUlMpxF8hc
h27+rwVkJelEhhGeTtYb01C7ygKWZnuhHr6FkAcSIPFHMRC3tQ0i7a9iOBJ63j1A
xqLQve6R152lup0eN61SQz0jWkBWaTzOIIeSegwqffV27PEQYWQWMdkl1MuafY5P
fmrghjCViRFq+GjHEiQZWLixVjbYmu0Oy0x2LW696vuSJ0Kcez0f0Cm+Ha2zwtOA
nVZnhS25t7+pZJKeDU3Voa0hCIlidRoOYcrfVrRzM0emgjx+v3lL3uM4WfmzGBL7
JDeK43DVSgXdev6Wo5D/ifRCoHOKfHumvWP2+f6Y5W357rXpsdO4WRixO5gn5I8U
BSMn55dgJhG+L2J4TEXyCCV7p2f9mzAH1nMTSdMhuH3fIXzsTFo3DB2HdHOp8bCy
6CBlq+waTUE3Fu8qf9yqxFiNlAlpSUwS5PmVXTxmzVvJzgeRi7E5xika1AcT3rH0
eQxxqA4X2o36EmZ8zBRYlNaGdXr3dTg/lEOfNyARopVI8n/yeUQxdIBI0aK5tutX
MWEsOFN0lt54Wr97DfKOggE2nAZS/BWHXfL3wdRk40xzptEWFxkESi5JcORkff7m
l3mk7jCCX3o4Dj7kAyuIFxnoqLdT5VJTI5ttAyhahoe5ZMwjt5z5wmJZftR0vN3c
o1lfF2DUj2l32ibpDbllX0I+77rjjr1IZw4k3Y9lh1Ca8sAhw00Ey+HAlwFU4LUp
Bjkb43cckBDo5eakTbvxWAWDAQgb9/UffSPuL9PLQSJ5f/dSujwYE0YJF87YWrqr
mRm/vwaEhc92cFZgS60BIoefGlSIog0Txgz+mEpQwD/k/kZsY3qqHnXB1E29/AQj
GAfSyp8tnaDujwPz+TxoHTcRvyL1UHscT98wIY23QYkYWFxu0gE4OrhIt5/EFprb
2r56ONmQY0rlil+7kw2GKaWQAgRllgv4UHL7PUTJdaFrbzUVSgouy2DkY+EG3JW9
KjpKVupzOXK4o0R4cvFruyPrYVL+ynwxiKwYkseNqT/ZsQlKRCH6Ntd2inwk9D9A
B2zYlO7EfxTjC41eSUraW4lybbN4rUOjLqb05y0ywBe3V0B8u/W94dx0AXKEXJI0
boK0i3npVTm09Rsgn07eMCsQ3mPPPl0WdYT9o07i6lalKIOBN8H5RK5YeeP0Jxy2
wcsT9Y2/04CGzLye9z/OUtg3aM+UDuwJ8nCbnHJeCfbYnPq1UkIocgwfSbSElTio
0YITNIr19jKVgL7j5VTk1PHiE6daH7wU7ZnFKlD/pJXRqIYkMoRA2+OG4cNh7puh
fGO0dPBDKHURUJA5b3q1tXo3ocsvpqMtPEH2WGby7bIjWAdVY4NFI1hxr1gVw0Ok
5lJjPlGujM7dELEDJj3py3PTx6OTTAXAGjchJBhrF6Wu2LiVnLYM5B6J1+BbmXx2
FB7pGOUIePrTvvj3VbpvwLp0HrNWLbGUPk7ls8Ufl+gnklvVT7Mk8JlKl4VvzGMK
+TyFpH3/ZJAnt9E7EG+u5Aui8B4ed+i+eqlGafY+Z6ZX7lhagZ5utpKw1ekLqw8A
Tz/34aUu5ufOD8oEg+tQdl93UpBlPMKzmUyQZYgijXiRmYrw3MdUjnVq51bDGUG0
1udz/mkaeUIkzcn1qYFhoXlcoAFi70/D8eVYQOVQ9fukwa4RgCe3bKBvhtudRYqG
C8Cz6bxIYb/qu2zGbIIGTKRHCOI9t99rRsvHV+Wlo77BTlTS2UyDuLnvXMYt7UQb
Vhgp1jtMldr2/0Ii7L7uFq2St/3RtkdcxQdGTFIYAuygIdZlCWLehR8RB0C9j7lh
/CZDs8BbpegC9U720w47UwtQDcYu6x3PLzsTtvtLSGglKiOMeVvf1T0ubV0m8wOp
X/XB4hEnKOcfA0emgEdgqW7YQj4/Qjw17i7Xnr5Lt+8zEGrgzYg3u8KsX6GOllZp
olQBzJAd9vE7z8XtfW2eatGCfpcqLE3lvadNnhOuoN/e4QHkl97vIuN8XQEMzC1n
EEvdLK2SLwrDlsGoqqjGsEYofeljCWhbixn7/9yIO5c80GI/XyQfiVle3B4S27VB
hmQkqbYtqx0dXyt3O3OE7yMqGdCw1ipdKBqORC3x8eiqYSJJqVtN4mmozndMJYuB
F1+QOk/5uYvBx4ZFxN1Yn3/MmNd2QKi7343YLvpjEd6DPg6vS97FFQcOVF4YKVRN
7g/+67akXqvfvHW8v8Kl3hEuUraRWnG6L/O9cZSj7VX4LFu2EDV44+jkL00AUgZL
MoDVzZhkal7YX9MYJ89mg9Lz9EY4qNAVY5hIh3ivpSOpLKPQNyp4CKWBbmhcsGp4
CBVMmVlAfxPQEwOuYN6+GgBPNX+ueeCNavahVUrp9C2PTGoEfcZS6zLg7UbdtK4o
nZhM8VTleUvdFb62WNOHY9WLKkWn/em91TzcaCk8kMpI/MEMHPWp+qQQgRV9IfQa
uc8Sffoc1C6naYQgac8aDnKS0eEziYz1BrZQVfcP5+acCEta7T2XqkvddO9n/0Hb
A6w+igRNbzOKHW9X5LH2T8jS74I3vuQNi4IHsseSQSgXLdj5xJhSgNZD2Ung3TTw
50dAqDl1dHVKnBdgmdaFVXtFiozRs9JclIiLW1iv1JQxRkXMhL4xkwlYZVzkDjeq
VfXTXpM6jy+sysmJt6oKT3j//otx/VIhnE0VHrq9F1lyVw7has0R+qGOX7e8wCrB
mHAdOmZlRSu3rKmE4g3dtS5K4eIjZDByLja5USs16AqEjZ6fakJbaJehFEXNxokQ
E/XVgkav3/aRfUq+cRUc5RCXTrXjnp1vBoymdX3T5pzGGfviZiF7FccWSkY3R+s+
rKSayZLRbSZByVJ7ub6u3EExIasNa96PhTwa0MTUDLU9m0XkxTk+8THxNIVhyE9z
6Vd228tO+j8m26lQwrXJahxF9T7LxNN1rnAWAZ+E++5eoWZJEdszhRRBH8KTMt+w
Rat2+mErDy/yuZ3SD4YRTQ5Os6OHODOqwG4l91eIMHcuImIl2HhJEgxP3c4amhni
i1wv3BfC/v5iRvV5LuK9vP73jQNsZiXi6ZpLWV9hfz1eUkcvyrXI3oKdJd3Fe7r9
g8wGbgg/oPzqUKUEzTQRUQ+c34UpMOlvGbcqtl+2s66ZJFVdJ8DhmLnuj2Zu4ynO
JpXwMVvVCazeBXowjosbUVOmKGgsooCFGrWHpThQroMDgp1Lb3CpS2nd+GsMWqtE
c19YOMJPd1rOhDalrVZHvfx9eqApuNLiyajQtjLc9t3FPp/P4zJXZZikaGue5ZVc
gVBLd8f9hlytgmkhNrjyirnu0e5rzGNaObqmiJDdBwKrHVXmDEtvm89mnyWRZdrc
ZKdOFMeRd+3ZILuYogiRkI/8oj77bXUPFTWZQE1VteQh3aHyp4MCe7AtB6rRraNd
ZCMW5m+/zB6FYU+EP2Co4LIv4eFPnb5TWvePPJ2gu1Dt21tyb0Yu7QHO1euk17+o
URnWCj71ME6fnDXbtm5VIg9Syx3NUx2Kme8brf4dSVY/rBX//d4u+Nv4ZqR5UyN8
oButba4oDXO6vTSHtik4z4S03hPQ6dlTffYtzO3OXTGNGjWmKs4zmgwVli9pMfAi
LZ9QvSAzTHZaN+fZCiQ5ZC7gUQFOM3XGgxvfR+LKpoEAGqiB7oVCxIoETklxQw8x
vbHVEIx8oRsf8CwZuRz+oZ4fOwGrHUlKfWwJJu0nJchwFu95Xno37W7w9EL6xHoQ
JAlFbTE6uZOxUrFh8wRRkeq/19V4Ph50ryuIPszQ39hUiz8Po3s0SV66dUJATzRb
4siYew16O7jU8OI7AQO1ltembz9kImP61JVmBjbZIn6qxFbUtxMa4EXV+dYcXbo4
DGXSGTd43wf6llYNFpvEjXWNEDaZBibW0Wgv9lli4h5bDbTJ9CjetIKhcrQp1Bw9
yo6XTrAoSshuorGca7W9mrAmnYQH/tTF+ETJbSLqNl9gwW/2k8E1fqZ9NX75H96J
kEvRM4VurxaX3S0q9sccqaQIAB3AFwR0vhjDaCUvnvuQurOTeP4DEzkk1yFUIvi/
TjOue8LXCRv3HkM32lO3Q9iqllaXG/EkyjYOQT4sJYQ5kdFuq/4OPxdnZJyy+KEt
dmb3k5ErbXyMY/0ra1CsixD0fjoKSEcOcT0UoZJvG1t4A5gqWp5zTQ/Q9w8hr84Y
D2aUG2+/LCPOg43HU5/Ek+mJ2ym3oy0xOT4UUaTWktptrxX+NL4StzCVnGMacwzr
1Wua766IjP0RYEyixwSQxMp1tmoH7X4I9/Z6JVJEo9I/sAfbEyf6vxecDy9YSzkE
2vNECXY/IdnAcebvJoe2iF03nVlHrAxYuKkL1pU+Pr8fstoT0z9TC1iCKuEOKTIO
u3FHL67xmZ5Xm2pCDM/KT8zAQ6CCfzfomSvhW6syMMRdXR7qA6lXBsnn/CUYu8Be
fKq/5bUARi9FlqZ001Q7TVUQign40h6xR52kC1wgFv9qlXereODwyyk8EmauXNlo
Ed8HxbuLmHW6J4/ocG1EujojGb0PoSwQVRjbO7DNn4+ZJYlBQL5MxiTUCWzRCgqE
CLTUF6cNBA7Gdr0c+2mzg6BD08gofFUPrtPyglIg2hbUcnKXG5d0ghCSChdZSBNl
ogFrnUQfpYgnAmnPtHvvqKHRWtTKXVb46fnkxtEGh1TJe+coeorRJV7xJIASBwL5
HtjB1IkhVN+1baX6sscroqY2dNXIEUb2bJxtSskisq00op1jUPLzp/Piq+vkGcSU
wrBxycJEuREfwTNKPjvL4+s8Qw0ZzXguA/FkDV/HuLAjuEgJcO+F84p0bUrJ3pnA
sm6mEYZwk2qLiWNbH3EE9CXpEWhk6l9DDBhX4AVNWZNTgu2oGsRKFvxDVToHr9UD
Ku7T8dRIIxdLBpKOUGKtxO6igoiRj8Dgsp0I8HByVS8ZhyqqhwCCWLBEpZsoZlqu
biwpDZxkSdi+1JFmHeKuf6WAU0HbbG5l+nFOioR83CetZT2APxRsaO/aQ9kbD+Od
yYaCGaz9p4QMiypfQkFOwHfg5ib1/sLTLvuNHR20csIYFVFag+KRIHL3Inu5OFAo
tuPD83XMkrhHY5r0EBLr5f2v3O8wx3MSP+RHjX6QuAIaYo8QZlT7JICp+UwH+l6N
awbhHSIpR8J/n0LhwktlgavEjx86IIGeWBdSB20NnKJtuw0Vutc3nMDqhGnrOPUx
sRimp0MLeHq2odrQWr1VWVB1jBfBBFO0uZ9Uf9UBVp+IglYoT8KMDMzxKq58WWx3
9mIX4UjRHKOsAkXGC0HwzOa5Wc55/DABywiS1Co3O9Xnv6AT0f8pPOtJweUIqMVG
B7eIZSp9PSEgyguIUFXvALatmtmCFK/D5s+GmYLd3Zbb4P6HPgYj6jL1ZLPWIdx5
3wJOM+KULmBAmtslGYYj+UnLMzL3EtISc0nCE23XK2MTRanpKpnfdgA1lNiIW7hm
arUIiFjzfAagFEvDF3zujHSK9XbUvoLlfaLawq72cEilccQgtr5lOBIzCZ9+jBEk
JFEa+jpUTYFshZiSGskrywpQZg3UqxaXGinIL6sxp7ygmZ0srSpKIrCStGpmA04N
vg8fvqtLhir5/Panvrcammxkqn3ARVsfgb7PFATZljmeNQm4hET1+/OiLNa20Naj
JlwB8viV9xTmUk88TdXcb9emk7rfUKNIqckgwFgl++yv+m3EH9xuGOYgIY3zmqhf
7zETH8sVcPjuFx8Bnfgwj+8xRipA2bps9PMURSyALjybZmgdGNAPNbvif2emyVeT
plbEC8YwdBIUus0VDw92UjmnzWIxrQA+CpwNwohqXxloAO34Wpp67XtPRolWLOAk
88oDzj2d3blT0UsDWoDqZHjpKP2h48rrU+PcZDAe3caUPwbiU/wrCPSfAzr3tKPe
hCvw10a0JG8opcROONwhzy3xHTNxLrJSjxjymnPevOvoHmO5dpxtQwLRSfsDKFPf
X6uwaCrkBK6YnLBSzeO1uIKFm/FGAwuQsQcZHwN/cQkTlBzz0cw/mPhWSWOfyItn
kYh2DKBbIoZLhHAKeuTtWrIOgWYN54D/WUh9r32TJJlU0RZE4h4O1nFMFua06yWX
MlPWgGe7VXOwqxAI4ZOYaC+QC4eih2+Wc4lfWBhdKeBFq+J9m2oCk+9AlBcQ2eUv
66dgRTS7Gyle62czWl93XUWX4mdyqgHJYPg1JbVngaYbXwCKus92D+irVZ22FToV
axisnH6q5aTNid+Qe+mqu+m3u6c9jAKbIjG69mvzpUVSs2zTicNHfVzYHucNl2fN
Pi6jHEwSK7ShNgVjHnaW/+SBarEQipMBCT9kbFXWrIWfGZREXPPMJqrjOhtb3I1g
ilPfAvcQRvVGwchB/j7xnL8/D6NiGeP/+E4Y4uqVV//3xY2qetUDb6loQniYfja/
PxhYwBeRQhS1hjtkXy6CizermvzYcRGMKHbmV3Fqd+oagUrfkT4pmuPoh1r9eNoJ
KBzPLF7nC2M+khxxXJRhCmJmvjtv3N6OwoD5IcUtShenT9kxge220ezNhhSkQnOw
N8hJN2oarfhjvb8/ODCLGtbTJ/vpBfX14MC55prQ5KgQ5jUO/NwVlfS+hDn2u2c7
bakX3CcIP5La6bGRoMpDWtymJPM15iC58dIXftNruRfpQnJIb4KME4WWHm0Snm+k
Sc0o8E4Bbpjxh31pGHV8wCO1u44JrWmyxnEE7CaShsx1FB1BvNhm5hUuYp9cJeL7
nipX4AT7E+KQanPazMvzyNRRgDUWV5m9thCsohN4FDTPGdk6KNu9qo/ZlscDzOBo
xUsF8RU1A7jgnZMwitNKb7NIaeFZVC7ehsfATcd7F8+D54EA6Aph0NJnXauC2C+5
8MdzRCzSqWPQvAt5hmoh2DwlqPAk84kfZPn9xwcTmvpMUJnqtXk2nil7JjCglXju
vpnftxyd/mGQL0dnKoxmzKXLl+IgDh7BVKiJk0mKtJDw2DcsU2bwbGSIjZSL4YJ5
Wo9mM4aomhL0vGYAG3WFay/9ldzcei+WEvpzicVGi3LNKXMJXdnr4khc3ITCNwhi
p/QTIOW1MsNgM4YBjSMn04TCXyoPEVP/zvOWrWBODDkNa/ZDV2iwxgqFnq2bYuOY
JrWLyMZsuyr1Xlu6zyzhERx9EzFCfTEfkjk3dvURmLBIMd29uX6lPj01JTZgmjqz
YqmDuA0lcHDN1Aa0a1Ww1J3wp/kJNNYMRbkNCMpz+LsbUV4Fn898qEEKqb+pUElM
51MBk8zyO7H2kVQGnfRrnJalWtTptLlcHaVmWejlQEGMhMXlHtRtK53WVN/ehPzz
YLqC3DQTKHAyKGkA3R50bwviMpuPH/ZC6W9R3Bng4X1EXuQkbnz2cD/RZXUlYS44
H4AuUseHlemuCOpU7ka1bjfUUJFs4bYcyjsqIYkElt4/NHTXLKWB+7lXzZsPgIXH
bqvDTzYmJUfiMmxsVpIFY3CwriQNZ+oYCcFiCkUQFY9Eg2kFYQbsLhoR5ZGsS252
R/73ZeWdL8Ftoy1fslrubGPG3lTZfRleydidcSveUEI2ARz5eVRSZFNPW/8LjvkW
Y96p/bd6hVUMr85h2xofoe96tWPQfCPRzIg3+gedI7jwSKjcfXyFUL2SLTeuvYuB
AXuh/ykxXZVzZ6XKDvHUvWMT4+b4ah0znJmFAHYMwrAnQCiy42YOmeId6F4EKOWi
//H0JEqzdUvzheq/+tRcyAXkG5fWuCGS66xHXL6KvDGWwfPnzfrp4wunSJeSyvHs
3OLuI/6fbR8Uulf1Le9F+Ir+ei5xBOmmEqjtLh3RYWht1RHJoW14nFisKheZ/Ipk
K73SDHReta+ZINB7J8OrZU+xoVGLPqI1rg6cXjMPws0X9TicVyL9kwXys+o5Nlw7
rXOdC18yKuKK0r6A62d6210x+LEpoNJ+d+Cn8eCZ7yZJQXtb6D2npK6Hu3V2108t
RkPilY3USwcMtq/rKJxWAxT41fH5lByYy0B+nlwzIhzbuj7BsvwoVy9JdptKA+uG
bna+aJhy5txTrmya5gl3RMnbnKl2dSemhGlnavkGf1mBPOGdUpY3ma0qBGdlXgSq
jOlJUyh9yZrGpeagdK9BLGSgFF/mfxTUZI2vV5+E7PCzPDTkKxwUkMnpyAJD7tfd
cxo8F6L5SRYQc5k01ipdX1JaT95xMJoFDgaY1OgmeSfTSmFfBO8X03usOndb6X/D
BUKhDPPsVekRgvePJh3TJBCW/FXTRPJ7uJGe0JZ/OXac+U+s8HmYcvf2qstwbyVy
glO6xb4EXMe/MYwz6a3jFpFSwEq+eRfYUh1hScMDYmjawt1bcFPg02XawP2t0g9/
UcXHTo5nW4hc4PMwl0nWsL0FH+JrpJcOsx5boyW3zs1aLMssuYGj/0ROfoQf5XGW
zUAURap0a02MAK7JdfFYKPpADrMwQTE2O+sp7vYCqtPp/M+hJ75pvfliC/HKjcw1
YwqMwUDdlvYgiSpwQcCTowjbLrVSm4LiJx9kJ1YoxGsIoGPpp3sxjuvolfBrJAqf
29VRiUDrKZQEUj53TCqwpE/FsxAt5Z6z4AgJ23HHxmwi9dqPG1hUYzHE2sD0O41A
9TR6CtAt7IHeqy44Aeud2vdck9cuK9iubKiPEb8CA7fIy0SQoBNoQmu9ehLhyY6F
kK0SuIILaSrKi9/FBpEqFxnY6y6MzYz9E1YlaDuU/H1L1NeYj8yp9B0SIxvMMzLQ
ADDjkURJTOW5SDVHvtfeKh02YB0miKXPDMZ8nVQg0OqRnN2fVJ/VgvihIBzuES/a
l4SgrNpClXOyDZwhQIQMHEmFFlOtMxvmY03Z/k3To2UJqqlv5q/DC/nIpy66lVg4
We1xHBvCT8Eo6z0Tl9iRh/RsRhh09x0YjG07mMoYjzMem2IYKOT/IORjjUGgHmYg
+5HL6y8IBYMTRAWYxqu05QwMtZeK3D2lk5hlxgnkoZD6/fdUPr78TkXpebr5MiXN
FNt0eVUkD5yk4Vyadg3XMwn03AxuUeATZ1fNp8nbXPVslAHuxAjSrCW4Ux6CqGa1
Y8yxy1sxr1D7Uj/BfsfhqUaInxJsipLfz1b38ytqNsgDIvQhLfnVf66/Tt5UOlue
GkosuXjEeR5AON1Rcdhv0G/O27maWug9wynh1WkHEWDBocPWhIalrFYRUJLV4nCz
+2HMibM89BeMsfvuiRiIjWQOU3Fb2YbTxVwBq1tAjqotAKv8NYp8DuAUukn3z0OF
CZ0r8q3WiGcboHve6qBFPIqYCMaGKJ0rv1xfo4x7/E341olumNdFnzwj61env9Xb
bCMZlMuEO+N1SR5vbx+CyztToUxNmBk/gnppTEJavb4h1TX6vl6ut/DA4b+Imri2
cAAW0SxhNwOJebvSWWyZhKNfmN7+rhFQ66sQssUmFF5uubaMFpab+eRcvex6PijS
2HRv5pLgDpYqplLk/1F+l9Gr8YpgTqxj+QRH3ATeWP2nxyqYh7p+of96yY8iWk8d
eH/tMCYr+gG+EOxHBdkGnN9C1e41sT10cWcZLNMj3eN7BsKO4+zEQ/QHllWo8kM8
oi1tYOWbN2fiW6NvypkuUxvGnObcKfMt+77AVBBnLngfa2NUgHrUPcW7NnwWQ9PE
ulbQmBL+7NTQYbG8+x84DGUZhljCiYloe/xrjV2LFQ5WG/m4rB4bjnignt3IqnYU
0DN71mfBxzG8ZAA9IW21QxBNhDJ0hiRdrOUGzgMPXJq31zKZ4y5RDAcJUzu50scP
4nWwOlUqCBKs3Lq1fi19TYPl2o0uXxEHxZ4tf0ZCMHYz4DKIQwBby5KAOEd5AyB0
oqszJ31VV7tHLkbs1XN1ZuMlH+U21Kh3GOOO378B+zDQxGxG32eSwNxeG1vVcBUs
J2eZ4sHkCc6KYqzzWDSWXxlk1rS/aP61sLX0FXPdTnWHCXq2q1lGiY0s3YZKfhmd
FsaUnPtHp2Z2AcGjoDT5GyqTTaGRlAfUkJfceABMFRImMKqic606ZcdphbepbXDI
R+8nqHeRcx+N+vhj8nSAxRsGeYtMKilLymPb9NR4SUlnTpMwzCAwQDnkICsaEkXi
TGl74kYTI+Ile2rs+w5lVfqPITU8HjoknDrp6nS/faeDUJuSvECo25nmHlXG2e3H
W1FNm+naysy8f05eQcaMdVGSwjbi8V+PTN8XL4HURhUuvbSeo612Bk2kQs0nQ9de
S/d/ip5aciQcqXonr3yvlCsE+HpZebIUZZ34nPu4WI7IorCt1KxZXhgeHaJERA1x
3CTKoWLaQ1Fl0SgpcHNzkb/av/aH0n5VFDo0gZiWbgap0ZwgZ9naxQduL9qeYnKI
HVnHMj0B5SfvMaQ+TaxuszYuVSvht8YVBjlHZrJ+ZCouljDiS69aM+sKhZDCY1bg
WczLQ5OnGjPhNSQnsP7h2YY/jHd/sZ9W0emiVmVeH0QzPz4XovbXWaCxMpq6Ee8Q
7eawbGOoAuoM3sV8250cnzflWX59xXe4OtGh3/E6ia5VYKmaxHDo9Fkx91wc9LBQ
WUlQflCO29VYvgHVJWaWivHHPSawH2aPpyZCsF3Y7gIIOzbVOzhwQBywbb6rhNkf
KRqJS5LvueaDWxg4K7Rqv4pa9F1DfqTPykkkfh7DZ5m4FANzyC0bhADbT60ut74e
N5YHUVr6kRew8yJrzKpHS8zFTk/uzawC6qPlcU7nkwCCllbe1ri9oKKFwq98cF8v
Otv06TQwnildmdT7Fa2Y7YDRI91D5K1GqdOPAMl0knoliCa6tWrv5z5z6I2LMlVh
3JlV7BwdnVDbxEc/0aAuMkncyW8rxveeQ0NwL+ZDTbOQl54NLBuszaDn2+feMplf
uolJBwW+0jhAiAU8peyBTt9lYG/0JR3V1s9ke1U0bhJVRTnl4dAjQ7DruqOVTfOg
Fclt5k4t+O5rhmkMpfjty4hA+8q0J+WESJl1lA2MMqkAib3MohAPpLNAMdFDI4tN
jPMyTJQRYPqwHoYeRu3UrfKehHRgBVKVVh6MrCBpywk6/qX+9s2IKefCW7DTEvl3
IRXTmV5pE16w8gWD/cPM5T0BdM1kM8qftBXZwOmei1lkgr3xw43cbYzLsyGNXvC6
8kqo+cOPBwPpIYofGW0qDmVOumSQynEf2kOvxL1CxY4neezWH0GHYO50uFPJ48eK
lRms0bbnX7d4hPPrQAVhK7Ud1tMHSst+SyPvBACGRw8dufXkzg5fHtpcURQ49taR
rG7yWZ15OIfMt5SYIcmn79GKgU+/gURUmEFijNGNQH2HUNdcH5uxd3Uzwipdih6A
5MnUaxugNqveiwfqFd1Lva62j7uiQ+4IqMhDK646M4XKpNeIJ6fsQIjwnAZxYJz8
YyW2cyBis/r7rIt9bgfvtuFF8MNKJ76jNr4S7EFYQw0NZBCyJKT5NNvv5urG5hyX
+h1xdGStleIk5BnlXEEd1b8/5+kMWMI121R3fnl/usT72Vx1EzERn/4pt5SkllRg
f1ojP6O7YJSC98N7qMjUexjSj67JrAjqLMH/7xTYqyihxip2kYrDQMs6m5oMDpgS
pL1M+fDiZmcuQV3B2eJ4HQ4bNVyTrJLJ/kTsXKUKiLuD/mG9KI+kV/DASp6EYmrE
4KbcgjDyqBlJhGHPg10BxUQTcd6grqcezcq7CmM+X6KSY+mX5xKTGuif0nsnJ+Zw
ZG8e1CRDofo2ThB8rMTUUSioS7vrz4dPICietEN8CgOauq3atUHKnFIzDxb15dqj
dXznt2AAMRbZMEu9Tyo0QtrjbRoWw9MdAwqBOrbvxxvUjnm66cFQDLjo7Maijfl9
EF5J5/5nHakLDRMje1HrbO+1YpbYXdKofGIQskK92sb4p7H69MrYhyvKG4V0uGGy
xAN1kIid6cbUO2nJ/ejqwhVYKNaO/RDOVuVu/FDq4Fu7jTuLiVIhqCRK4N+fl05T
lANG0j16V+tnaVXp1dpqmhxL9WklLweo5D9SXNue0DXNrum13QpUae4EBA2tSy7F
de9vW04vYtTyR5oBcD9gohM6wX75Wol+FAGtqafoorYE9hGLBjzupSibOl/aD78a
PHFs1yI5oaoJHPxpnyv5XX8yzJIZJDcSG682ScQaz+bgIpLEx/5JWmv4mtJPbTdn
LZNAmcV6XDR0WMRNRtMe33a9KSKFEEZyjGmzIUb8VfatE21d0lADcIKmBrySJJVI
ySvm+YLNjVycIWGaDF57k8cCSv7bHwrdgEwRM4tODQE5jPEP7+Po+o/tCXIGqqQv
i3UoBFJdXCIGr/iWjxfqWsSmXtxdK8MQg0HdYRTNvkzOZBrguRRFs8XKVOA4ECSL
AuwbzPuU8amzV/1e7iEtubQmMojhN3fq0SdtfSgDurScAN127SNvTKp8OK3cJu4c
rbo2zBD2B+41no2+9FczDEK1gK76DgZEa2rRbSKiM9EInrMvij1H8v9K277FHMlB
F2KKtjS1SsvxQGdMXNZ14eslcd2WCs8B5hM4xXG5vjJggXT36RyyaNuk2h/u4RzI
0C5zpBoRvHIgO4oSlr6wmayRo05M9vn55N/2rKlPvdH+Oekhwia8ebnETX9vdy8s
7dP+KMR6JXjDz7C84Q6pdWHBBIgwAUB5nUThEX2H7JSeupPsJWLrSM4k57LAQ70p
6GTRKhjb+xviKMfMExMpbIvBqJzuqSCMhn+rK2gYaDHSj/RtWKhOd8Pp25VYC1bS
VYkkvMw+/8XqvHh5GN9SH9EdMfUBcOUJt5nI0Ue6CeeZEtLRxYK2JJ5T/6NrGds7
izZONoCD+HcuaCUy8ib3a4Kx+P1ul7DevAfpDm29+PVabVEpCDIH9Kxe2fUZLmcX
9Jalw4gFfaKB+lD+ojt2mp5euOBhgOgS8IhNg6H80A1Ng+KtjUL5ZVsEyTw/bPzy
ZS1U3zurXCVIm3eQjmct6SkMPP8JG8WPxMrCRIoXCqUJzVlg/rciunijVzPaZill
ayDtbjnYN6pcHnFqa1AhMmSYg+GdZLeIqy4Ff0IGwRDWH2yczOstTyb0JonGbnGr
ld80b8GX02GXAAGt4lt6erNBbNxyDkLONAv/khbC4mkeJi72jEimoA6gr6ki97E5
43t16C4ViueudoWb5DcpOj+/oW4K7a8OgpCFHHV7/P1go2TSKCfxutaOdYFJsNWd
/qeqBfxwG0NpiYMXCvEPQmukgMYU6kjiKIpTk46OalMwwfot5TbY2sipWRr6TD4S
0dAjDkoeyHef004hc/hbqSEtEiJ/EfDNXVIQyieRUbZti2NdBVmqD2i39unQvUJI
slbMgHDbtCcw82p9KiL9uxZylE3iUKlxRl09KKgWpVHGsrKwS2/545b5jl22nXFf
KaEnQLflGldNZWRJxg5QEqwa4c0qa+fKRGV9Ei8kOygpXx60siPm+/kebf9uJ4mo
/Q7dS3Z7YrtHGk+qAfqC4i0sI4/984cjUnZhHrUEOL3XoLNIER99Jqhibk9JJ1NT
nPUTP489w7iJ5ZpsBVtOrmfMZpDuFkSLFeTZPZOOL1Q9XOZZSdsHOyqes5hoes7F
EuGfPQIbYfTNafATmW+SrVR2T7dgDBOcTU0Gvy55bs6yvlGcBbJpqUe5rWsjEhUr
kXgmGQ9xKvf8Ar1HpKqTZqF4tl+6qI/w7ODx7CaWqaOSCwfRhSeoRQPm/uXtE27M
rwLBTGKbNmhQ+W1qraErf/CPFkN3OsnKhBbzGQ6au8Ai7e2WXlqjqyHyIoeJm8ii
VS6717KhTujUmpZiXbFknbtm0XF6s2vM39Apsc1oWrzq0cKSSuTGOUiI1Q0AuO9q
RfI9USDs1kXI/H+Ln2xqsUsf57vt+5uvq5zt/cQNzYeBRCLs4KeuoJJ4ewxgk+hh
rSVME0o3nmmODintRvL3IPFh5LeuWPRbtmORN24yeunjOTt/TBfNdmCSq0jbWlfC
gTg5TrEm7q6m9UlH77gSNMWY2tZRH17zncHckIn1vo4E/We2GUbPHX1TXPsMmvuI
ABEsHAk997L55vOoUWIwmhYxHdtmtI5GyZIk6h1u2C8HW5hm0a+xaDqVQLFFYg4z
LiEq/y4kN37ro/R2p4gUanKCLwgNXgV7vcuFiGq8+/6+nXiD+8Jp4CbOoB5vLiMh
KIMQ5yaoxzqoCWAmwGXZnC0/6XcmAFfBH+CwuF9sGhue6Wk74xtrl49n4cbkgSXD
uedz93vC2pIp/T4LSfaG6IkksfOhjGlaWf4XDkbZ4BDtStEj4LzkOdCFkoaF7NIr
oPLqYsgaYiwvZS0oWyCWQpo99gBBFcjbYq/3sb+TI/F/eM27ug6q54avry2UqyvB
11mFCWmYXZwEHaCLbMqQ+4ZRXuQ9A/g1mFM6AFQQGBau6iIKjWIuOVcFrWYbJT85
o967gXq2zErUeHnWmF27ldImQJOdo+BvkIFmVqY5xDbwgZKBr2sYvD5uKsyHjSxc
+MIn0XZcZtamKDRCSfULa2WaoRkhkLaJMBDsew3XUSCYDoygePOqAJ2/6bopMLRo
aA30pyXOLH9GkzoMQP6jho/VvLLPJH4aSQ24K+xR5WZ8oSy3VAR9EU9K+L926p4U
QckKWl7uUfxlm6asOzc1XDj543NgWHtSWJjF6a2cX/y910rr37Cn0POgHNycXY+t
1wuOnfgVbVGE0RtTe4AgJop3kjUfQDaP916hf5dGWy3RlrrE6ZZhL8Q8WwDfk0xC
1XVLVjr6k7z9+SDs8UX5aIXq+IrsvAGMLOFwbeNqGJxZcMk5hcLD8O9wl90FTsvG
YhiTCA6uzFO/pXnWUmd4HcPkgcxPiAn9U+xyO9wRAK+krSC5xBqOsCXbM7nRIhlG
9JFjX1aWQrxoopXfRNWgvQl/MhWGOxqCuMwfNRB0k8Rrp7NmEuhEzRJ3KwoTzhg/
YGcUA4G0eNZlekp6y2l8dTk8c872xLdq6AUDtZqrQ25hHNuKxNAeQpXQcIej5N9R
cCiBcZgJMwQPFFHRWsp4Tl0asJEDzu4d0fCW/kIrV6EPV7Skj7u0CgiKVUbYUXuM
PRFA2PN/1T4Y9MkKFZg+J6B1kNsSwBbI2GCORM4anyBKRhLHImmb9jCLFQh+cgOf
X5CiYu65sknmn487M4pS97R0npCUgAgjiETU8WUnpChIcRaIwMFbG+VRRKBAVeAX
zBed7QujAnwRIG0deTEGtiX2wPUAszo+wGgAOC4JEAphoYFw0+FW1iv1yFIsA6AX
X8vOL/A8/z5wodgKjdtU/APOym1ikqlyW/WFEtQpUgwFksGmioiX6Y42ETFLewQA
GGmwXm5c4U8ekI4hFKnltyIrpONRtvhQZGjBzC3VhsI6TAe4FjjHzwND2n7UcT3z
zLO0kUcyMfNEFVZstRBiwYF+IksXmHuRuuZk6vrOEGrozUkdYJvICKtKqH+NsFC2
d0r6cfRfWjlAJ43S0/jGBiHU/BFHDHFzSnPy2mPjwJi3lcoLfSvKC0mlBJlcJcNh
zNNApRE50nNn++oHpaxbIfJodSab1CvCLpKPfU1oRzdB5VO3Py7aQcAwCRq80Un4
zh5mpvafb/C3eD7fowsL1IE3hS4ssycOzbIh9E+EplU4ulOSGCI8gSq/zFNXrShw
A/h+bWOJnAf7tVeXqLuX5c+lIkAm3cOvLF+6x8Hawong9jbs/K06LRF6Af0CTZDP
r5BduAQ0MnDrNtEyjeRSCtjtuBA/vpl++BhCREqRofNgVs2wRiPc7JYhwo7VaUv2
VqmsflsAlI6ne0Pa0jGtqeuoT19BqWR6JMTRrYXUJ8n4q2TZXL72SfpagC/xNql7
TaQpSjL3akyB19tSAw5ZeTnmAhZOB2HZtEPy1j9vi+VEflcCm/JpIKJ6njPabMTc
zei6niluy7JVCMx/ZdieoHv2GcQamEWzmOLpX1ftJqnVBFTLP/Wbm8EZdel8RSb/
uzqgbXijlfzpnRXALo0iEmHn1KXIuTZrIqvcGoZWN+21391QIjfpK6rSAJQo4puP
z0KZFMyvhI1bhVxgOwOpDtMdT5NMXng9AJ4Pz4zxiSs5Y7Gl6yRl26FyfdyDg0nL
yTjewjdvmm5eT9oc2ZYBQHnpy/1LETH9wTlFlwfrIr3lw4C6SDcn5VgwjdbPXcG/
G2ThfIw+xgNFImlXN28giwkSvCEzG4VI2NDJmMXa8D7GL0g+hcdqc59lcFj2z/vH
HuTl4h7OkogjoZO2utOSrB5XLMsSaaF1N32PHgBnJXXCQkJL70I2eFmZP7h9V7Ds
8azXDEAHp3hmJ3Vpi4uV4Rsfeq/5xAII5aGx/Zg4mCLTpyeEaEDyXQWpJss0jN4U
b2Wm3iTxFR+nMtAIN5N+7RMvXBasfdC7LgL1KwALExUC0x8tVOjoy4eqwspkGW/h
rMAhPyI5v1ZljzcG7Wa/mCzosFJIHl/sAXLYxOpxT/lC3mXU209Z6lIglYyTd6bx
WbEnYCPLTEzbjmm5eGvJvZWh3DPWLp/T6hsffAWvQNn3pE7coUF4ecxSSEjV3mq6
wVQk2d7Ft86Et5DzqQOPKGzxrfFuZU7yRb5AVKJeCALOaRP2oGYG6i2RDCjrruCI
r3KVUOkQI4kC8TrxlzqFD440+WWmVkZtCPm/XwCB9lmmS2sszsZzDX1XikwMheMS
2xUvb+jKOtClfojFbvuyWcDnVWQfHeETdw0MG5aHveR3az//3klLaFoUkd5P5q1u
caymlDwax7XxkcvzvX0XEKTAM/tz69RaStLW1BwR3t2sgFlICMtrLn9jFeKw4RfZ
xLX1wGYtKgq1oleeqkFVJ/zUi1OMa+YZIHIA5+ACtIT7CepEmqzWgMuivbufh2d9
sqEYg2C928SwSM5qxHTSWKC4MW9ediiuCI5yXqjlBOryvJkYyikjB3R2YGFjSTB2
drZ7W6m7/Rt0FKxU+ALTqMCMvoRGAtc9dUCUunvNs3EUdb1/CF8TUBvPBEXAU0JK
B9r7Y/6rHDkt6/3asVkYZ1LSjnkeFaA5Zbg0YHNRVqCu5HnKAFNwkIYu+k8eBeXh
xevdfoVMpDFe2tLqEcHj+82fZuqJr5qXM8hQOgBfzJ1NoRYIUTGygLSiQ3D2XleP
BZidDSNPDRT6yNMcDTeaalTH21Wj6t73qWWhPOkoAWTdDlVbAECkpC4pWnADd2os
m+islEEsFA0OVaAllcOzBNLkIiHLKKUAH8e3fF4OmZxJxVY2iDsdKwCQjk2DYjlO
wNm+jIN5rv77BS5hLCfoqkMKEQWcmfbPJs3kE+VQrYf9SMR3d36xRxW1VsA9rIen
Xl8u03iclXXOYGYiZ1E6+KvuTc3VFC+/i60q1mD/M4b6+u+/XrG4Ti4HPLPlHVDz
YCZkzjoCbRuRIkkBDsx2D2Z8jJSfv/J3+IOAH6VjES5y4TOH0WeQQAawgzYSaZO7
0fOZJ35/dqcbBjUpWS29dZIVIKMf8mIed7aC46mwXe9edHHNHwvqvtwBudSjTJwa
yHJOp02LWRbwTn8Fm7iStK/1BQ+3KU/h95h5pTqp+c0InMq5Y9hXsrva3MWh+ic+
wvaApAkrKtpoDxItX5eyZS7KNnxjGHE4mZ37yfCNAbnjYaH2FyoCrC+SR6alEknn
mG8lRvcBDUYNmQYnII6Q54BKL0I1E1wbVUM9nSCaZ/Kfc5litmd5+7OPPN20Nxz+
5AT6CJ7TkZWnFeuNy8ocHDwgG/6L+m7k3SYMe6aPSd0ZdI81M/Yk3wDYuOH+ATeV
uuFQyIJIhYenLDw3ezhhoz5nnkhmBVb6/aUeIWTLBNG1dyJomC9/WKCOoaDG08au
crwrrJmTqOj+5sLIFfxJ1qKZh7tGmGl8cQkhYAaC8y9Vcqaj/KC12Gr4HYzyLEZZ
CZjxeQl1j+OaX91Rpg/iCWSlkyouJCctORUtiGFaPbDB9HJJVK34Sblx/TJEXC/Q
4LGpEi6jhiyhk+gaCbwe4X17czzzGqvwnhF2CGSGY4CclOPv67xyC1M5DnliC+DI
761HzLUHUA2dM3q32Bp9OprlKRLzKfKpQVM5xci4qioLXCLIoUKXQukqQV+LspBb
pYq0/jJbXKlXumv2OxKUuDMynZdfLqRdc+L1EvufxQlMs3ZgduOKAbSgoJYnxLrI
SFoSIew63frCaYLUItNbbvY8cbtN6USLquby/6zMOo+DMR7clDd1B01n8mN0KBXT
AhKF3rRytjeXWYfzjTXsI1sQ8Iznso/7QnklFjfSBSv0UiofqoHet68NXAhCDM+5
/allUOVJTGHtMRO8t8r31UFuIZMuYoJaUqDJHONYc7c5UHhklBWUbpge3+7jp/EI
s08Z8ERklErR6G51sPazHptP4gS95ONAOksPl2A4HsixJQfo0Tsp6heFk64rDMas
80yfaGsBl4KTszZuQr35MTy1iUGF9VZTpstPa267WkQFuXthiWCDf9Njg6MyuWKu
Jg958E3clVoj8aTnrI62D7eWNvUbvlu4JpGgRc97jD2U1lu6HPz7KSxKFxqy2/J9
J1NmsuFw2J52yL0W0wOyghJiS2bqqITFvXKozX3/mvBrRwyBsOyV6pZjbaCt+ga3
0lD3v6FeRDWJfGQ/y1B0XUqrPO46GrkVhEj0//MT2fvOB31aLYHK7YSEv7cE+yrw
mtZLPefTZeGxgSq9oLD+iGT3FNz7WvD0xjlbrdAStlS8baWri9wO251E/Wy6eyvi
uNzh0g6El/PixfLiR9cM22v360Q9BAD65FJGc+D4ue5Q5OrJEw/wxgI2y5dWPseW
o1Wsb0c+y7BHHbLuz0yKwFU6BwKkqM1s1NskcOrBXeencHQFtoVuIpv1+x6879/j
Qs1K41D3ztTmabyWc6v8yHOAVhcJKlFxXuMAiSWWaToN0h4NS7VecRBVA92/4wLC
ZW/TZGurJXxz3D9PmPADI82UKlgwItAr7UGHrQ+pwmK7QdIzZXG3h9kxrH3n6rnx
EqJ/0gPNX/eBWv1ItGARqh3zGC85ect4KcPpdN7RTgP9gOlLMP/SeQasP4R4gjpw
U1/rX6fKkD+Y1GMTQE3vaPZkynlq+utU0bJmm/Ng/YIYwGz3dd5xt0i6kVFSSIY/
TksRj7EsYCPUDIWwN+bo7TZeDn/9ccwDtArZMp77SCQ4IG8jpZC+hwU4Ebs14Kjc
Jq27htJuf1pFUBXs1vQVk5lakWTJ8heMl7IScrPsc2NF2bQDsJPQqQrpklk9ExO9
ttCdHzun8t3YfYswHAmO4pP8VI5ebRtQHv8Mgy+2Nl2v9XKSBko0HnhZ81HSR86y
mxC6RF3cJkipkWhpx1XZbhkfE4+DPzl56jxx4GtzIjeqvfjgsP4UO6Grhw7lz8Fq
ZEBTNn2rKXsT0vXeD0BWdJYOS7nAkQuywuS23vkwkGadx7tK0D/a4P00CWWanOqy
NRqCX/WaJ4zYKD0VdKjbFV+c0XMSJpQ0Q0RdMHHlSJJ4LP1BU+V4zeY80WIffKAi
ekuX4No03cMNpJcHZxFf5gVe62XOJulIQzwrJrhqJPsuozAnWoVwxkeWCA6Oc7Q+
zLpLSQcyjH+3Qt56JkNDzL/yI8QwkxfaoKn95N/igxer3z7mrqFxLQSg9sFZ3Mc6
FeIinHJR1ZvQY4s0wWsczMPryU1MK4KT/TCF5UeiscDBxTIiR+UWVNjRWx9UHLh/
oQs4vi0XCsIPirsHdvnDuZmLED79MKedRZyBUqa2DDCG/qt5eHmRtClUf4xeDQ41
oJ3/Zbg89GuUUrW9UsWqsUYWlIsJwtP7OQoqgX7uBWEGm8pMxBCpWOx7e/jsnezx
I0d1RxqInevOaQHS1F/DrDZr67ozknjTbkVr7e/9bizOyC6t1wMi/90N0BN8roKx
//cFAgliFc1A8GPemzmceXTCXl5+gXLY6+5PEbyIKF52Dou9g/bRuZa1cS573atE
MDYf3I7cyVZAGxwN9fUqP0W2CHGAz6H4pXtpHdpOqRxbsNlRhdkXyHf095Enc5dF
DzEoHI8ONrQNzxwakkyhooOkKxlGVBk2QVl/Rm5KR6a2z4NR6btohRfMBqTN/eu7
cwBEyMJ5FlCwVBexNJSbQmUYVripBmX502I7LUII6iGBg7LhU75ox3McOeNJXVam
XA0AAGhHyO2lNG/1/oEwiaYKqeceth79qxZGTooqC21VE4j+vqdvvnZxbsSQcb2p
PjUWKOqHjAVsjzvJbMcKezQ2Q4B+wefxc3veUDr2KFKscxCO7XSXgw7ktLEcPMi4
GWHBF/p5V1N4WoJWCffb84qazuF1G4ljn2bc36AvyQFXNE5oH/4V17xiRg0WvtF1
GsR/W2NAhmnXEo/lJlvYzl4NYhWzWYSxoFSZ7aLqLxeLcoD8A0jopwXxhunKeUZR
HTzvrDqwdJMqvOrR0DesZ3vXAXRUv1VJQbfo4eYPD7WavpBz0mOWzFBCFmWLumfh
A6Pwzpq0PdKEzBVm1S/0ENXOxBiJJHnX1nr/kvmMu3lhhXLQ+KAHRxItNpTOwia4
Xr/4l+bks0OA/irKa20YbieGGfDK07aWdMG/MtvFzRDF3lLFwFBSKzs0geRSCPXR
XwiKVKiY1JnvfbwuwhER6MzUU5T6AtQZNVJK8W+EJhbWtH4o9vM2lzTE59WFh5y5
8RC8DVeKYgD2Tc3svcdJaLTF+ghP1sg/er2zlXoFxj1fTc9M6RbBqnlr2dlZKyDV
bBM5gVg8XLvf12B3A0jHhsb0rT10w4r1MwPdTFvqlMY0QvqHBpUa85iijKLz16sM
g3UkWAs/Tcm9rp6UssWjaFzuqV5FzUS2vC9rBF4RDqQKPn6SKOabnjV3ZpmpoD5U
haC01ttsUOT/vNmElmtMVpvEdVybLUfS0o1VDBVJJnGKTgegs5wtWpP2/2pNh9DT
yeH9W6zl2yYrnSJutk1nvOvJpW5gvGWDed1oq6jAiOYQFj8OepmqZzWXNyC8Sy2b
KIxt3OHWGdxiGrzllfjSiBKWEqNfzb/NLKxhHIbL21BjYtTWmAwPbUlcS5nuK1rf
RvAGRft5nNSuwHgrraGgq62hsQ65M6ZlrHetau747+ub+KG6udUJxoPfqa9DeMkl
EsfzZmo/Lxyy/hEUR57iL3d4BQ897cxLvna15Uv85K2e7vweXOQuSHFdymRcoKa+
q5hYuiinLTZguN2B8EGQkTdQCCxGpP0Qv63KGcxZvNCJXKxIcQY1TqTkVEZVelt5
N6Yiu01H5v/FMGJb9qfTY4TeqjB1eFXzT2OT5shlrNhBw8mkXfu0de66h/nEWDA2
SwJfTSWzpTcx5uqFIB0wjIrk7ovFjDCF6se9Dc6ZImSxlXyNUVWQpprq2Uibngz/
J4YVbrTu+ZIfVHD5lbaiDES4/ZOiSgvWlle2kFx4WT3NMYbQJp//OVi864Ot6pOe
Fa9SIRqP48kTUckEIGNC2YiLf9bpZNkkHl1J0N9SwIJgyOsA1xrzJJhPiAb4vhCG
cqLvTVYx1a/onf1yHjrxvAg34NesVm9kjuIoFtSgofSNwsUq4heTu4PG5YuKAGKU
OM8VbohdZDx2q3rNRxePpQNkQdEkiLjUx+BAbQEFjBtIRScSNBI7ds5VV6JoZ9AR
eo/KkRdourn86XoiQCLmIweqrM9fkefFMOrqztHCvYciSgR6URJ7n2tuHwm6WpSj
5dOghCpPwwrF1LR0f0ZyemlpDBRszqgWG8nLtyu2vnLXRm9fva3Cg0rApt3fSAus
Vz+hBWsPK2N3MCxRocODIm8h1CJqhvQL0BuASPtkobC5NRo26CsdgYIAWNfSdgAr
K5/QXn3u72RsDX+Pr6Isiap5bhayGALB6brwAitXunlnFuCYCcIkNodUt1SY9EmG
WJo91wTwOQXhuZ/MT+3aThshkL2Kcf9Vp/9InkfICrEItTROqLxZinGw26VWqdwe
f0pYKmOOobtFF1kZ7BBaRz32RW3gQpStpVhy6RML8rzCOv9VKst4gDWnVWCw5R3P
9UCBmEKD84axfkigPcnmJhjDEpcb1eOAnblijLf93HCGPtS31A9+Ic9Wy5U4kFBk
eG3WSciiHfSb38RMsZW+wmYIodlAABtA4L4eABNcIxmUUB/OSOMnzU5Y5tU4I41N
5Pet8hgLYJiQrF1QjB5N7eMQYTYpfz8fJCs0lan4eK46jh5dRIfLQy3aLKEr6KZF
2gjsGWA6Yr/ou53dd63KagDPDy7OVRUXnoas30ZA4f6svwUhEKnjhl8WfJNtk8gS
YbAvNpf1+aJQkg4UU70RE59D6fMrv1bp6qUkg40E5dCE8FHZ7XoVEMBF/UkrUlF3
8iqy2P0G1nYcFp+8LKxHKIFacJb8/Okypr3euZgzacrBZhpRpXvEPK4i3JwSixEx
J/5hfo4IMoyZ/YDkTfsUlkIg4ONaVGSPjQcOkOqy3SkQpwBG4p/fzKN1QTy8s9fn
HJRU+fzmVIVKrkiTcFS1Y+7OcAnnO97DwuwAyukCkTCxBHr0+jj6bAHoznDFUhID
mxkJRJfeLE7z/x9tsiTiAa84kDw2H51CHBSc/DFLi2EJ72uoTqg1wRVDcTy3zQRJ
bAACvMg1zjjcnOuFE2N+orZzMf4rr+2tnMNwIPGEw9fP5QK0rDPS+ImfoTkZjZC7
PZxwDTIE0uxCm8Z4z9J0pI+P9Fy1rNloN1yTsk0IdAYp6DU0BDwDwHRwXD31rO3a
f1uKzgeCZ/033kfhgDxUDcUz/IjQGZzx7GYx2s0Q4n9VbMjA1F0hNZLVKsMe/NIc
BmLjdEfVxRos+X/NPYUGnftgjIrNYTMOrcmd/rYdodZQeJZRaQGVg5WeOf1X4VWR
AAQ3/59N7cqU1c2RfkalZCXUEQD+PS458aRr0Bc+/fr5b0/DR8GVUQ+i2Eyicg3F
Y74958buQbaJZY0GhvJYB8n6erpOMtKd6xLGg20Jb1vW7rClmuCHEU3/ZNyFQMC5
OsU2cMeu7VMeNBu3BmgF/G4rdCOQyRq1TPo/Vygh+BCQdDSTM32eFMRH4yvz9Ta8
c9ct9boIqXF4biwpv+liTQshJ2IRIamGmKzlKA+yllcUmZD9TXa36R8gxwECBz9/
HUirypcaNl6miblODq4Mq0ZbKrsbY+kZ6wz3jDuq0Ih2/BZX2bAle7Q7y6K2WFY2
A3IkUMqSMQwF133Iyk72COaWkJcYRbJ7Zawnnq9oUN/cZSYe5sT3dOFubvio5aUZ
+xCeiSjVIskpTfOwOdJzpV+eT4z6G0ebl+ZncOHFCB/75vVow7wYhb6dacUo9vB9
G2b1hUQYpLS23dciGFloBSQ2U3jz9QpbmwpycYSo9VJ82kJ4yjNg6/osDyEwtANO
tQ+NyS33kGl8jc8cv5ZSQTFg36pe+1if7cAL++QHjqo5IGjaMRKjk9Dtw8N1eT7v
Vru6/n7WoUru03Lo3CuQB16+zrddJeJNc4CaWzBbzLsQMsgBJV0eDOKEaQVSFSZt
mvYJRlJpsjJmd/EPQJfPct1ab4ZiN9y+XOnaiX5kJ7SySFpNzV72ug0PGNUyKvB0
ezyk6NVUT3OHVssPoyqgufly4xF4Hwsa9xlzyJG4TIjLIloF3Hcxu4LxYV3xD3Y5
pTnpPDusJN+RhWF8XW6Pcf//jUpc3iiWVqvUya7lGGjVzfdRiwRTI9yeN1RDwt/K
uimcw2+WrQHll10/YZTPPoL9mymSTQYa8E+/QCM5zHiZOrS+WKZZx1aB6UUC6RdC
YqQoIwOLZOuW44ZdnmUcfWNN+BbHaidUZxU9oABvk1DuDq9YSzKJowvuSn7R2Suw
Br29bH78MEeFI9B3+MxUHk4uoR+PQIo2Ys+Jo4W9N61m8+gIfF+DwdENyjrhJw+z
0Ug/tOO1jSYU0BLjGyguzrGT8zgZQs7VedENE623Bd/kl1DUTNmMaQyVQjaVz21F
R7rjWYjW39mslgp0wFRkSQsWcJHf1G20fBiPLObe2u2bOxwX6ytmZDqJBzhMD/yy
wweS2xsjW3oySiKL+hxUSsw6Vnlb6nnr5/DtvAEwfxQUg7ByrIzNSKzEmzfxnsFc
pac/1uhMyeLPrL4IPnhuIz0D41IPQt3EmK2v2iwA1ZYB0YKNAHPjMSG32mcaJqQe
3ERXwOya8txKtn7E/CEUpTVclPYQGj7KoAj8BaeAXTIm3LoxXdGn4eAGYVEYloY8
X719GFS2Db9BMlXX6smRXbX+ocF2osB/TQCVsXB2AVDQhWWaTBATxIej3R2Tlzo7
PYxtf5zM+I79Wc5TrTEwMN4YHUQ0z2wUT8sNBePHl1MuyU2RvQULOxt7RZveCcwm
r+eBK8/USvYf+c083y8yMvQMkhSnucm813Pa+tX2K2KC1MsiS8Xptv8cQgDvkHMy
f617+8Tr0oloj8S+SqtlTIEnuWPc3IPqW0FvOEM6D9LjHz84ZswVErv0ZBQcmWUj
4P1ktXSp9hKR5syeor079ysfmYCvCSQOCDqafyc8+rl1SvHjHGLV/o1tcEkFgQ9h
GNfrSfLK5UcudkpMvB8J310W4O+1AUCLcIF1UZQPoeqqkEHuNqphXIy2Lb1Q+/S/
pXpxmrvkX7Re7oAjkqN14wf7EshWQftyajFR7OKGmtHst96C/iGBUF/Smo1fXYTB
aEkdEOafycmWl0GXxEZGgm3gy4mCyG7cVPhH/0sjzf0giCp2HrDhX9eHrTO90Nqg
qHkS2O9c45FdWNC1jbkcjLGb9SwetJyIz7bj5sN484E79UqmqUmDK7NZn4yygE9n
uMKImdg4KJs6T4MAMm/ZfOGdniLtxIlWHmEqQLyNexUFbrH2B/6ZNwCkUPx4ouBt
LgtxaOZ2kgE5nnK/+qU/OAhSaa49/KyjubnXC8xxsqXgiXWH6PASqb3/2dDGQEHE
hsuPP85DxlgsUy5ZyFwDtug8TTuRujyupCitNiINpLXC9rReo1Lj0ranPME6fDXc
3S5dgYJPCJgejWlMA0yXQKFEcBjwKBNRJYepF2JCvjAQbilYQt2gxrm4JlfDgf8C
VocXlT7I/+A+VkVvE7hgeM6g/vmcpANA6r3VKF01AWmEoT94PJUwvKVsYi0MNOWB
eSaNLvFHNceMUX1U5v7trBH2HCJD6sEQSQ+Ei3KDiJ5A2MwoyWVkwj+Xg8qcwgxv
QXhf/8EDInqccTENUMzk6jaz8MDzoWnoRGBnzatVIMIBDsAn4JRHgr9N+qRG0cYa
2Nu7oqJrn4wAhOxS3MNVine9la8/HopoccaV5EJFwpCPKtYJZMMSWkZbfsIeQowx
YqcbfE1jGerkzOaEWRQGKyRcRBcdlsGcjmM88E56oOLvgrZsGoFG7UQvN1C+usl8
hoTcAGPbS2uf3vFPHCTIG0KqQbzTkXq2Zb82WTK/7pvt+SvkyXkjWrWETK9w946C
4VeA8x1av1p4LjX/smv92CalIR4qg2mTDU8mEfCCr81BafnMjqlHyNIltPb3lenQ
/w7W0lvnS5yUyvO71H3cv4fs3/woG1LqKt7RFlislSEOFZsXd9glltV4hUmsI2tl
n+9ghUHCNRlTzgECamV4XC7q/uBXSk5p6k4aYipMiVjfjkXURJlZ9soDYA9SLE3c
QfhQ4LDMcIviJJQXm3yUeba1cGU09VfX9ASGqBShZKeZd5gwndOVtyo63PMkS3RB
v1Q/XyY70LAryVjO1j6Vxoka3PHvCmzNXgMhH9iXSGYH6tZ15Dxd6DYklThrMKKQ
IjJuTglP2EO9GK8LX0bfJVmHU6cDYCGFw62aG/UgxUy7fLPSDJiYY/Nw1SE8eLp1
TS1W7m68WQj70EpSnaqmsTVr9mDm4WfBK1os9MwMDRMapoVptIAW7rtfxQXl5L7w
zM1Ryq5K6UKkjG19wDCOlCj718+XtBqlzPjPEPEXjeiRdvzEcE0zGGK/dOgQQUyJ
G6gEg2WLoJyhC35Im6epNpT50NUgYTYOjeUIUNqzhYuUMBs9PqHWJJXQRp+ozLEn
gHEStQm7TxGjhkF6OFl7Eik2Qz6Y5L7BiMsHTfEBGuLsRD47DqqNHoMD3IIdsZlW
uwR3h5G4GAj64yY/lvTDbfvu9S+6xz7i8SVY4ioTrW6eVYneXnLNTqtkRm8YqvVH
zjRQEbcMeaTSDiWuBMLcgkZgqgdE8KW9raw2ovJrvaCGTegdndQXPR4JhKcB1k7t
u1m1vIGXgrBHRVU41GijbufNeEF0x5dyA0LbE1GPySwbgKEbe7gchjWdQVgKk4/O
u5MNnqfkO7akFG0oSanLpRrf0qrTKSueOl1KRBa9ouaZaZLLfE/sONkBlo7iJ41W
QMYm/m2Svw9jDi+GjamiHbK2cFXXxODI/5gt9Ej4ojfkRHhbT1l4TG8fUrL3zmah
ZzDsZXdJbJylIteH6avJU6KxISpLLC05pb2TVs0SgucW5B5fFY6Rs+gDg9W/0nhG
5fRp0YHqXwqJ6odDI22P7hLh0LS3VIoy77ro6RjeGgHdeIPiUyCg5yW/IyX/Yz4h
/jfQJGZIrXMoM3WTHIr3bKVVzZrNGGBaLj5CheHLnqmZpoZnbrzynakIde/IN33t
Kko6lMSwamSEcwKLag1OAcO7Atgi8dG+JcqC/Z0lhoAV8+jpsnFKH2cK5ikahCPP
ONDlUqN8Yj6xIVmMHHco8M7L/DKROA/uP/CMeP3OpRiV4GwNwy+uU/XLilVBaoFY
hZ1RYUvXjX1rJBCqNtitXh5s2O1Vn6zarO+h4G4IBrpiMrhgqpfo61qBkDqsciFV
y22Az2NfTJfz0ns+nRRX3vCnjKrojcMS2oxASL2ISQFrerQog+VHI/Zg1DJMzjPp
vKtnzZ8i1RwRks/IfTa/1U1WSmz70JqBsxwNskwiAGoropeb/URsFL0KVNs0El6d
4YqzfkD7HUQ3TLszmTsPKDgOkDxqwniCVQaZ/kpkk+WyVqP/b841Qz6+RA8BIow/
9BXTxNKdXZo+dRhQYqLKFPS0ONN841C4ywnPWVqyJQ0fWHBnZetRpYu0xgEIyZQ5
PPXd3HCpYb8doJj/ud/4qpeK2tOT5U/nxRavimQ3ewiktRx4NGWxbV9hwiEdahMW
AuO8x/miWUD+otxvomZ2p5CDxYPTXNbSdNYtfCwUe9zpkk5RasxgiBQK1AE6HWvH
fwQnLrf27RFBSh7iBRCtAksDUWAPXXDedg0ephIff1hCYf3P0cR+7c0ilg0CYSai
6twgJkveCj8zFHE40q+1qAx5WoQQs1XAawlfo2cechKpEHooSV8j8i/WWllcS+Ac
gJtHVOMsEdi3z5UMzy615yVlMTrB27h3Ajbwt9wG20XlabaGdGKun5vTCtOP6pM5
IlNFbojYgFn+x/8rH5CI2rQ62StOe56PicmqvjO5aDL8B9EjizW08IZM5CVHXbTs
8Sg0W4NHxfRHfpwi9PZ4S74B0mIw4ExFBEftDR6DNpqY9xLVeae6rcSkhUEg6hkC
MYM9T/HwwLFroZiN9z+yNloqiLpkb6Y7TZHlv9n9cP/ldvpFuYXqKFDKlf/dNtAq
5vpMixrWWsNhgcamrUDVy34qTTZHop7NYQpAFiCvuT/VYBjfJE/WEtiGiiGxmwD0
l9fBMCxZhKjrABzEd8TKWh7JnKCuIMRhQfetxQMzGzCJOPBCAB+UuW/QN/Kf2vNU
SYTFFerU56UqGDDvJmYM5BCmgBkDnP578tjjUk3mgtBZWQoFcb2hgazMOLuuhwcl
eXOpB34y2eqRat87Z9OeuW0ygGM/Pn3UE5RLNfSehzq9Cr0TcK1tkmdIARe3Dex2
tBzC4sQ/j90fVuxWfdRe9nrlgDetRV5xzlWOqO2bdiD3DxtQdjQfPKKdSdGq0rgy
gr+Jnol/XaeEj1zznN54k9Ueyoj3y3zYZ3u98Z+HGt3xK3uEIJukkMafUcH4H7Jk
6lGs5+eQeFckqKA66qTG5V0B6laHRpQ6fNwxv77HbCBq+vMoYHOk0/TmkrL1hOg+
vnbSjy+rk8swBubmemP1d0Hvn3tvXEwnaxyZ7Kzz2HqJBmUby+6R1iJ5uTbdUssh
Nm4zULkhhmVNOlTtJKo1zvIQgjwfwYdU3oeE45NYzi185Pa3EJLkVnsY3vsXoHVF
ZAhyMmkdL8IqtjLeU7Rg3z3su9Kaies3wpR3+DV50Aubp3jYXPhJKTn7kFskKiRX
OEPNm70ksQsEpPoXaBYvOdeb9QsLPtwH0iYuimqTl7EeFyCOIfF/5i41DdHYqMG6
lQN8z/sxfiBHifHVDn+Z2ymJGJksW7YCKWcIAz++2b3SQWIOBrT+9xPRo4Y+BaBU
1agP/dBdhwLj6Z8pNkS5VAFR6iuDPm36UeQDdrLLRK6ubLqWNTRRzFfHQ3vheqRY
yx+8L/+HzyXd6NQpvLLwLFYLpv2aktPwBj+SxSl+IVqcJ6md+1PZ3eB/C/XFfNk7
R6AYp4CF5vCV1X2n2LzAl+xWYJGt5ivv9kP2E5p72eDOLJQgb+kzBXb2f8o307rE
2WjbNa7010eG9FF2eIzpY0GeAr6KliTk9kHevlNO3DdBAeh6K2MX1lkgUEMx1hAU
PkOjwNlhgrCOEUulGT+SY662zM+zudEYfvBldZiSvpz7yUeRjcSpmI4OcgvHEhtP
j3YU8v5YZfEDI1+HkBRtaww/2/xrRady+kR8bSbsPj6Wda3nDWi1F+qhBu8HXmnv
USOMIn73Tp8DSTT6rMTH0h7tbB1FXANzVTUfCkbZH0WUIp2SCTuQOhUCKwqa5zuv
oruqjE0HyJbIuck03AthipVAf/qzlc58mOV81xi6aeuIm5PZon++vILcyEAdDC3Q
Spp55UKzW2X4fYz+wFWVbcJ0Oz5g4oRmmIWoTzoix1X28eoNUp/6u0nD+GYiaO57
Ag41ItL4nKDf11tcbQVCtWaqfj2qQxL736nkxWmiyvPc4o/3XEWZOQWQUyMvMUlQ
hlPmRsBNlmEO8G2EDSPqfDYJKi+Z8nwgN3hbySAZbe60FJbKc3ArieGO/m81Sa2o
qM/WP49iiDg8p3sOSSPbBJlfT4fcQLzRsdnjkw2Isu9FpuBBzYdtT8GH0Fjfr1TX
m1mjgyBT77CNOgd6B9U2dW6uaXFDPv4lqEy3FZ/z1pX+qof3aovELRiVlN9Oj2q1
PgpHj9zMDhCEyQ+e2infEXx6SbLpFQ31dxvBS/x7xANQKHZVhh20gampKois8QjP
2nX8WmQqBL3xFUMIO4chEaEKFiYgmvb7Zlk1VhMsGgKgq/e1WiGrkMCukaVk1+rd
TaOo4DVdbZu0xZcEQjXiKsnmsYXoOke83svYSyIumzIx08nTChCwTzIbBtBPtsLG
7mOSNMWZTyriySn7dY4F51qFwzfsRg95bT85D24XqrzLxE0QC7bUYMN8j8KCFjfO
hKfpIopMoTfw3J/Yz76jCJLgZAQbyFp1gge1d01jiX8HU/xOP8xG1r/8CunUwwJ8
aZrmhA4Yw59wmmDwMWkpWCjRuoTrP6Jmaww7X/Xcx5FjfKMBNVmqNjvLIcYZkN06
fGNZogZgqcxoXgA8PmdUlrCrSFHCB/hEJPjDLCRG1QADkvE/zfgQu+ejiPICBpXc
xSJRV4lry6wKaWLt7ZsZqkEF4zuonsnkTgtdvLNT5Wx9/tssHWFJW1ERUDAWu1ye
q2/SDSGrM5JYAG1bjyBt9MfC+qMQpuvDfIKFpP5+VH6UzZ7iQR4wT1yFnfvIfcbW
ocnChlG5TQTTayMnB/TRVLrT5zkAk55/wLhHHpmEWKuhXnur/UN/0pCEkjQ2CYjs
KtYInS6HMEriysn0O4G4lW0ayWIitrs24sxRdNO3n+C29wzhBWQIcaJ+9WEjcTgm
r1Sf+Oes1AOvCM/f6N88KzdOfu/Mo20FmHE/diTVx4qwJHhXxK/El4gfh8DDPiAy
F47tbZM2Rt96l34jHImKwZle1+SWQ4D0hfK+NrnaByNDWy9Ivh+Nt2fPbammRGjj
gOzIzvxnpuKS1DZiAXbcBnhfR02hFs3uyqKC7OqmzWRO9LdF1iKJI3znMPZC4u55
yicpHknevsnYaI/Evz+3vHSrn8H6WTa0lpQUqLhieGVaxXdglD+5qk9OTByvmBzu
u2fdjI1+E8cFIMgQk+pYGw8Q0yJ9ICblUOos7j3kiKcWDhmN5yOR9O6FK+DahOBz
bVYoKHPAR8G2iwGhcqkDIwAAVH9BdG5O4BYx+jLHioygQGlZSFi1WieCnGZgLMbN
//6IFuhxXaeuIH+80gnOC5qYfpODM+mVFViHmVFOi2J5orVFJNtGFM8vPxk1SFzr
4b6xVPnDma95SUW80Hn832+vIoKLFLLDpqUwxxpuEd8cJpL5XMezeVSRq4RjAaPQ
cSDoyLupfjGGBM37EkNten3KDglVwa2245FACZ3k/O4AwW5zNdfcmYeHQ4U0iu5C
v5hENRuzTwtw6pCtZb6sxQ3oiB/MGhZAmQmsHAjGQIl6dhB3uUhQeKaiBmvbrFUa
3bSIBKQKxL6q9O2Q5GaaFphoORHltGN4HFb0VVr1fOVAoL/YSnVJuCQ2VrnmpMxO
sMG19qNazeZ9CS3ReG+7WKbcEkJ7yXUKKoMUkiICye3/K3vz+c4p8pI8hgU0jPFl
Sw/M9IpMK/e4za5NsQNcmjYGqRLrmR5EaOkupHZbveTnTIQASBIYvX5E10aryz1a
/Aim9aWswHreSpsY8O9Wwi00OCmjnh8jIrdKFLd6eypWjTQ+xzHNqlqYZA+Av5BN
xtjP7c6b6PAuzqbJ5jRUYCKQeofmVfjbMOLPT62D3H1CbKbFWI1DGegb5X5DJQr0
uE8T9FEyxxKNyuOrmd3izHAuk9zhU6dKzCBVWG00dbbtrVEexV6FFGB6BEL22Q7M
KgGs5eSq4XjcRaBkpt05ZVg//8Adx6Srv5HWnqm5IqLOuHX9JWdeb83l4mx2FS67
nBeSrzeO3irQ3lyQMfPlU9swO/eZXrAB7iMaX56PgvT8pYnh6UdXXzjsXXYgRM7j
5HqD9uvml7q9mCG5b1C3Tnw1CtRpdkMHl4GZ/rWAKxJtUw4x7ZYKIbpp6Uy3uQYD
gxmMu6RqAFlCpP4DeZm7jteumOZjVdnvZIxDmkF5T7lY5qxvkSWyCLk/S5wsaOo5
nb6IAsg2iH4+Gee8HKH+ZLXdaDfgNghFjG5id0Y1ZyEzBIWvJajzw0CcP21JEPvK
+sf13tpqY/Cnsbb+wF/Igt1E4zxEggEjhwAfXy/he9940Um+ZP4U+w6wZRONCCS0
fozgPajrztSSnpXeS9o07kbFR7m8oRXcUS4iGVCJfz0rgqDf4S1W/SRWcT9zGkiJ
r43+Fhp5EvFcuFbRJSuP+Rm//YM1dKVgW4yyYcoJs49FlNrRspJ+59GB2RfuypGc
a6mFo/u/1BhZyre9De71NrkekFIZLxnWbpeOfH0+OWcyfzRDREHrlJCtbzvABH3H
9JkCA9shNlWl1DQgwIIQNzFTQ6+7ivm0n9P92vtS0iP+E9ThBDDv+3d8TXK0vTq9
sIbof67uFpHmpfggLuoVtfwIXIFGHS4VM4waVN8WPS+mFqVduj2FQkjCRmRa972z
7tVWTd8wluDtixSdel/E5ZnE2xrYRSMBVv+N0uH6JDDXOTrxM1HDWi/4AXnVHej7
gtp5Fz9tAJmyYatr+Kzz2b6oCEpF0//falBuGO4WvqJMdah0a+E+SnCZrOqpfgX7
66O0TfFcfX5ABeOUw4/PkY4JcAn7wp3ws801OnaWv6fW2v8ma5bmVGFXM8Whm8gC
b5/hHod3yRI7spEXgDcPy6oUKHnXZibmEwPtJfIUlLXzpImvIaik9h/IbqBY1Scs
xydJL3GOo48/rzlMlI5wJRXVEFsgM3x0oJ0YVgyM5eWT6kO9Yggmyxi8yFmNSzXl
vimUCqe2iPNYAjjLlQ3Kdhm5kvI+pI7FEpAl0w9rJY0uPL6Sh9U6fcaPAIXa5ZmR
8Scsky7YRSD18DYKnzdzYsP/o6HmmGbcocNrpyCpOP62j5k8v/Xr1N4/17nWMdHS
RT6Sce0SnAqoaPWyXtB00twskIpEFPiZb6t3nDcyqeX0994Ku2pnO/vo+PL/hspx
MR2bgCVsqMO34UfMvzQAwmG48w1JZGO4ZNiCVojsSWCT0xb3xgQr+GMHXTMOwyTj
ImiRbE3nf3TsBrk3Y+TWdeTbBOPzk0AXff1Q6V81d1Hvd6BAfy5UiQ6neYaJ9aEc
akyWY7a+z0UcDl3XPjLStZJISDLKBZc/OdNct1yKUdhAb5LgVUeF6QwTbKIsg5Jv
hDtdqpgi8T4dncqIvkUctv5ZAqu5Q4OrKNwS4KnDj1qlwelzSfYIlk29EXIw8R57
N8+CNtQFx0tpfIBNUvYbbmXtjPQX4wyB9yv0pzkWvblJN33F92tMf4m3mzU5Kw2q
lVTi0kd8QIORDRE6fF+Lw476SFOccDit+cc6+IIcXa++JJylxFz2WNPiCVTNKVqe
HGDRuFtq7dkfy9T/kSo4DOp0OQ4HPMSN2SuCaMfVkf2N+lRMiKalCKZDN87IaUcT
SN67/v3PTvcL+l7BgZJyryGU/xcI+kpIS0Q47FOqrarTjVQyZJdWfr3sCix6taE1
8DhyBC8XheLZa/DucQ9rvRuCFpI72oiDpQ+ugRoKXOzzvRx/DngHbsFIom/jVEv5
jytvNJq7ZDoB9qSDdC7Oi+MTdvqzmDQO1Ypw9mhBwVEvKFfoeTFPrcvep2Ux66iW
MXlgF7KydUwYrwsDclO6Ygkg1Y+/Mt1yAxLxEIox1YV/vtDfWqSqUvUzSxhfeR3y
Q/3gAXjQ8Sz8zWnx/UWzddRWkd6rYHqZHRFl2FbhGGK8kAyX87MFf1mgYLwq3You
zAH0w9aW1DqAGUmBoWZ/+gWvbMKi1fgwb2uuFXL021xJRHsu0ipa/ROPdqA0yGhA
x3C/h7b4wYXAWL/AQ/DkX0c/prpMtultU8eIPF3zYLuqY8JYQShl+Mht/x4lm+bK
YyT8z+h7Dibkx5JHwwiOkiZgMvhuVfyk1X0iWTBdGYtz3FtU/OjZVz5Q1cEOSvQB
LwlW+T1OCAlFBhGTIV35KgcYU6Wmonh7gqffb2vKZ2dQ8wCz+L7NqBggdz82W40G
K7SoGwCSpEDHHLHo/nsqa3DkLo9092Yc5wj9djKiTKk5WlKw7Kf3zvZPC2wMd/O0
c23qcTqeIpSFvwXPL4JUhRlLqYxR/YDy2gQ/5MkZS69k/sGeI3oIJbExMsEkSDQU
cQnoNdurLepBd2qK2/mKkempHZjaNxnOyKo2yxdnvm+HZ0dv64+BCnfn22GOIYyk
VkRtRzyKNqA9Wp+SszfcFRKIpVGu6jN24I4lFN/aBXbudD0X3le9dLQwe3Ix+GKj
pxaaJPyCeeDhLJZyu5k7vEwQqnuZ5MmzNVr8COV6eSYYjw6fF+l60xYwDEtCVjhd
Qdq4U4ta2jHt2wkZt/zjaKhLnzvd2kOzFtulXPkEBM3s3JlrEcH204A/up0yAn3E
WIcMfp8qg0fQQEjSivEtFqFxmnOdoQV+hPb9UYAk7DEndVJ/Ngt3BENez1YX/TDE
wPIzrpHS4WP91TvdKJ9IXpKDei/6W75EKzjhja+uUefT/6XVB1tQYmzoVLYyaEho
FUNjKaAOLmqBL4NXDHbIhAqCXZe04vLmv5pO59Tz19JB5vr22SmOq9lprqXFD6kw
BTmq21k2IsbXhdSv3dRqaBlf3r9K4LUGmwOi4nab7qH5PfmYL4NqMsF90lXXrFNF
lDxbhNQyaHf0OFgcZJdm0562zHRrDF1ybDHPrmBmT0+yM5A2AwHqFyJNpISLz8Up
o6OVUaterxw1xi+Dh464urIjmxehlxSY+wzKGsErm1KGkJZrXuTRtib+kU0MwGMk
IjsurGTwqgDQe0fjh7cvqp+rBYVob6qk0hck7oypRb6tj3/SHXHSyXD9Fkb9OGwh
JeLpaAWSce4aDKrwwZ5AK00RiWO4seUMZkrC0So5Ow7qypuQkzXC6e07WdTUYDX2
Fc0uo18AKgzEU4xaicBdbK+gxerMgHFLCME8gvtgYpAxWpReyKXbS/a4mzkNlp7V
a0BjlTIH8DV33ULoV0hGHpe/gDT0tpae+svRVXDa0pB6YbIArHOc070m2tzrkuoJ
sZynOhJuLb1IR+jkzaL+PWGuaWkKESXHsmBHsCcexXeOeye1RutTcMNYFOBfxMsR
Kl5/+5FSeIdcDeTiohBBaac3yu5mj+vP+WsEpSqS+2saeCkgXKfvL0b4ZutgfZ81
L76ROyQ82YyMwfkbJgx1DDsdUHKLWnfjtFvjk1DNzDY4fde8HeDWY/0jAMfeBZMQ
Js93u88iV8wjhC2tOx93gqOjUWO/WcJy70KSiTx3Rdri2Q6rqUC4qM6rccAV7AnT
uHSgnSCQtJpPEFK7lph1G1MnPomin6JHHGT/X5gwqvtWnCRL8HzQFVoXsQ2gOBmf
0xeGLqZTIZaxuF1DgdExKMpkH6pWv9J2ll79zGst9RtTfQBYSqUpY/leRU21fvKN
42L995fGEex6Fbj3S66mQb8Sgc0EcdR3x7JOdClxaLVh6ptjJqdirSEnAFQ/oLjS
mHagcjaSHF6T2/CHv8F0x+Cos+dA0tWQYFIKO6B1Heh1aL0AgpSRQn+uJpI8vSMB
4Wfew7JBLWspZmb9RvrDu34tuEKuILmoCb7nl36ASEC3X1LMP+qoP2A5cGMqIsHS
l9OlZ8HhUG/LIqaSDDCsT33U0qEXVo0YJh1ora2FAN6BH5Y0vsDVBQXFI4HPtO/f
PdBrn6q2i+NgL8LCCq5hJSyEuyAoq3LSWIt/SZ00xn3E/JHY4Ab5EaunU7WxDYXm
fyvvScjVuwoMofMT2LHbCyV1RNgspF0LZtjTxjF+6iP7NiIE7m1pRhzLY47KJlQ3
sWmfsrec2u8JOyitPFcsFzZVyg8TIKfEkGgVeVNjex6pxOjde8syB9yzrY+GW357
MbWMvxG0L3N0czF9XUfkkuhZePqzT3A2z9nkhVDIv045xPgKqruo/3sRqNik+x4s
AFm1d593ftVH7BEKey23SvP7Q1ilVng7WTVBMhIezMV9dh2+JK7Vhd6/NwjTd8S0
RTOK+tnltpXNl3nDAHH6nuqoTCF3fiwbKwp1KOhq9B9wHBV/iGStbjCpTpIoKQ7s
jnAn8qTw+R8mHZXlM5izuhEgu++ew20LmilFVry+5q2gQcRy2TbzHhjoa8CVlZrR
mNCWLDlygGGo8oPqN1tcNaRsUB79g/b/uJ1P9GOujeqwC9/RnnVNOXTaBtoTGtqW
zuJaHXCxK2ZOngFOm4/+7c9Usys1uKQ65B9bQUGRbAZaNIO7a9Ryo2iw4vaaGrNP
HNptLgl+ua1qupSpu6Jb/yu14RAMhg0XIlCvsrZcQprA633D6WuHygoCr6MYPIfX
6JTgGGYIbQta9m8a1J1CjAPkUSG0hLxylUWrvJkZMNMVQ4qwq1KRpgzE8CKYy4du
10P0c8BZvIHKwpSonaFFbA+Im4NZSLzuuuJt6l5Bs+gO+L4NxUZvXF59zErR/V0n
kT09wM7rAt1Yjvp9T/mo8waBBsrJbzxphRIbT8EZUJB463cvAu1MEWOZKJT739AT
6sbBnMEKND4z/yxH4QsXt8RLLnfC5UwqKRMjYtEdH2DkTZXLmwqHM511LzlR1mVI
B/PCjelyqQIW7liFPAwnhgmTFV9rqFj2yVAj7t7nJLI2K9ofdTJg4mlPWGr19/pn
tra5VXooOBkozqL2Nhdi/nRbhK5MLlbVE6gaqFXAhCSCAcADrtXgfcARr7PGCSp8
Qay0giL1bzjNeArS+5WbTgmrdjyCoTtNUeYO7nIP5BFgb3OcvsjhP/SV+JtuarNn
R44aASTcSSs7xgIX0LdtnFskeJnTArh8wvbfVES7vao/z8pcI8QzYgsvSfjQ12kY
JQm2QXQepgK/Wie2PTgdq7XIG9Xcv3eTDxEf/1ugtenu29ILAXMzm9GlpGkGjrnL
hzzPlWKrVXKBKl/iwUT6CjUnumTVWLo3RCGwc5Neo84JnzZCuIV0NeF/j7DV29rR
c2RnL7REGzi3Yo6mttaDVYrnoHL0ULZCrOkP4swyd8dWKHXLvij/oBfQlKUgXdyd
VuGJd47nZeq5TlKlsN5/uX0eMq14+tsRSSauT2Y5rT3ErF1k1xM1ZwM2OFMaJHNC
8Ifhrm4Fe3wEenNRWGybuzpP8HlZhe+PkaL4FeVrFAhBOfF/jaxLQV5MUeJLAI4M
IszScCea0q5zlbk66k/vR+Z5SdZDWvzZjHh4sPtwTn+kyos0AaSS5P4BjG7YpEdC
9ZDfwV4dJsKIzgCZqrrqIyyvKKXAl5Ip8kbLDCblD80IVGMV+aF1ru6KAHZ4iW2a
BK4hnbKtDh+qJockRXyc3tcG/gCFpb9b8cshcMESfeo1yzUZEh5tG8aorGKJDSMR
2rIDM3Rja5l+uTZ5xDaRIolZYrwModAfs0MApWacQB8cx1Auk6mcm2yC8cPhJzuC
nu1Vgaxqpbbc4Nz7xuSsZpxU26zmEMRieV4ZY2MCknivhSByOQrmOpZt9MkVs8Nl
t2f4meZNye00MjrinA/uW0NuwHFZNxQJ6QL2ZHdRGLoWMpQJHL2XrzI4JHmhKIfL
JkBwZWnQq6tSxBFbSI3VHLPrBSeK5odo2RobwNFzvgASXeP0R5nC+EH6od3W4Vyy
KQDgebDbH8UNONznSNWFAHhglUuAEwO/C0BQNc4OSou97byT7B7QqoVRAahVW29+
rz1eY8I769PZhadERwEgvvGbBSvuG/xqpMTv6Er9zQVS3wU6VcXZvOo4e7xZaaBd
DIt/oj8TFQ5zbB5nTKTgFYIQo2u5aVQrLa5XLJ5m/1TTNS28iJyDMWs9zwFxqjkl
+/G/MdqwXbl90OOzETnLcvmJ8le04DumiqJiofw4kH994y523zgjFW0Qq2zsj6JL
z3xBS1fy9O20PM5SElTpG3I/P9WrhPKKFzsvvez0sSxLtvBtO8ugoMFH7ioQEML9
R5nqZTLMSmeRdQu2sfmWFv7wmKelunBj1c+gq3yVgnT1AEboXxSwksC3KU7WCIc0
XLo5QQQpsuj4O5/NG0vkzlU3YHt4+5mN1J0+dV/uwGTIeQGZXqwAQXYpm1syKfhy
o99CndkfetjUS6hKFaJvv/YN58iL2RvwxsVxC5uDaiE7uMGw2vlTy8ytfGw/hhhK
8ZAFDUyDX9g0Zk8exflaUyLWXuK28CId35TfkPRNfQr1bnniyGyXh9UaHHgHqobm
2yUiGkwnt+3DuMB//x/OgvtIISIFERheM1+y+1fsh1st3ZKqHDWk+AUmjJH8oRrK
cz0kkDMvFk9L/pMZRXvd+SJnbedEIBw+pCCXaGgMpBBvFBL1jwFZHd4gnlo/rbgX
uj3RoOMXHr4YE23hoo9xGT6U9uqDavr6Zj5BwhIBG6inb6zpq7H8YI4FslWpuEQh
bTDiqm/sCvGTDV5UKESl6kX/thzOBxbEkxdinv9fsBcFfhnHGXWMIm//s+VhMU0P
lrnvLV9eN951pReRb004gl/MbWDJ9vJbjyb2RTpW4HTsLZZjzRCEG//0N4ENQcwb
8DVgPrHWsxrTeowZScZgpJcBYv96ha+8vkLhB4+fe+OV0auPp4s9oFksASuRaznk
kUpsgn2DWjsYNzgPY0Ynh4BSbArjoDvd3LTbBWGmWofxgB9XOqXrJmSsf5AwP7xZ
AGliIxVTw9uJgCQrKjWFmIgVZHgze1pB94FK+oiyGhIEKbYnAxbZkl1FUhaWW2gi
LOgUGFF6VRT9bBeYPBsdjmu0PfD61kDRS1+pSfKwxMf1zEH6WgTSGNImzYGQ1qwn
q3s6MmO8j3OzDrQZc5Oct3EpLxwEw6matTz1AFuCywNnu5SakVtQE2X7PZHWTDpw
nVHOBPKdgI8Rz9yDgr6GXHk6X9J4JMiiN7PlmdhwLegr5tpn1DB9fZms99YY7Xzg
cfvFeUwThE1iZFniopKZUBKnjLT39Gjish0tbQLCUX1oxldKmJiTlp3pBDkoleU+
CODJmRcmfv5ZDK5+pVJtq/JVFnqPE1Fs4dDKu1437Gn9J/Bq5XmblPJ/gF/wS2rF
xZGR3VzCqIZ0ptRJ83+rZrduqqePM/9TaPkphMZz9dmu2RtJqZ4lE4t1Krp7fga8
0s540e0pqwA0wH8VaAQwq8hajTBhQuI+867qW+27hwYviiQywl/ssRvsUttNJRx9
5BWJxNAUZ/cNuDOUXiQR+ZUV32d5IIZ0XyJQ7JWH852FkCbzJzSzeKspaDIqWp0A
UE0LH1hPp/MhXlBBtljMZqeVr/hY4ya1hN5B9jWpYD2+NmOOID6mP5Z2TewXnZLv
viMusWugd8ewYDSuy4KKJheDaT6m/y9IUnBZS8HfZCTrrBtam4n1OZn3ZX7GxVHD
sIJafZ21+e4S+VIoEY64mXdoX6VPqsml6irqnCBjkjcSUG0Mf79lbZxOhE5SL/in
JmY1tY7tC+fknavF0yqC+0I1Sl0HN28dxotIH4epgy2ylMVIdVsTV6o3+n95WMAq
zSPDpyMcA+9JhIWT4BoNXaud8LXmjc4pNX9FJXdPk0NaCg08fKB/BQylIIfSZ64V
LknyviGhryzGcXlWh0012rMYV8D2gaSaRD+SjJVPcY01unTXa2vKHOPdEAGcV2r0
4FHiyvtN6XRrOs3xFDXbE5CUzq4xmaztyBPGajRerqOr541zf4Iu5ASTXg5XbCzc
fGhlqtccbEHxpuLLNhPFxaN2dJI7W05+uVSgNYSwR1ptW//grJwQqmE2AsljGlfY
9Pm2M2dGCevQ+RhyyQDk9d5rB6S7yyAjaGjONhhszhnmTuTzkO/k7VYR+Mxcm6hu
3gN2fDFIinO3ctbbJVRjQ6+MzX1QGLeScdmg2S6HEyzDNncIKBA+e3SjIC/AEa7P
QREvBXg3JIyjufUFmz8z8+S5J3Utlt6wHzlZtGFWalRPHOjx2eRbKGCuq6Ui8sez
5HXMH22kI8PANAtXH0G8MrHUis/xEGWPqnjdpNV2WraHveuu5wlGMlVR9WY39grb
79txq/saMquPvlx3XG6hFzLFWLgmgu7zWAIDlv9ln5mI8elx74Ry03fE9GDtL5O+
nVRyg9Mf7H8JipFRnuyd2OupMuEl88ljR0C9e51baU2UTDhwUTk174pkjYKMJK/r
jGrf4nfELu98q5qX6Wygwk49+XzG1vVISsj5GA0f+Bt/+X3VxGuwngYE7fdLygE7
/01XLhV/hXJ1i7eSHvJxoOOz27d5WPPSVnzGgTi4VbZYPF25Ao7Mw6+1IOhvsuYo
jUkAror4D0tG3tCFzw+KLp182+2Y6FRy+JoACzkfpvbGh7e6/3QRRbcDSDzzFh1T
v7M4paBhYK+0lLPec1xhfQRpsIugIgA3ciCUI6KSWSEPIVCCPXQMkldbC5nalrpG
B7zD/Cykq4caFMrQqEmYtusTwUjG/zNyMcPiRlhehqN31NT3nHPizcwmRXBShKw9
m93vlFpoZEYYuf27F/E740eSBccGq+lIDNOIH6a/R3LOwWGMNNOa7ytj4XcPoAfV
1Ui2HKz/gMaVEoF7neqG5MsuTZeEKo5PyBJNNM5O3zMFSTy/7AbrBZ38PJBvjI6E
P8/1bpUq711mVaurSbFMQEOTxfV4pVthN7LYJ3KUlx6Wtjnuh9Eb0MGOOTf0WNJ3
YIrL4BiMnRng3GUF902QDAv/mBRUps2Kn2bVubZ3K5OSNJvqa4tebbtcz8C2iv32
1e0CkMgPyGY8CephDtDvo7EBDJwmQx2Ej6/zOI9BS/KnA87789ObBxp5QLEz3CEK
N6yMry3MFKZ85PDQN/Vr5O8jqU6RMSYLE54fEbGDQ7GC7Zq9cCv+s5/KLDXbWLxi
o3vANOtg4WnWK3y8PsgS0+dsfuE6IE2vo3B4XaZRUac3vnME87ZwgIJtYXj8M86F
r5AAx/9DZQOUyrl7Gz2MhIiqL0m61pV2dKG6sKtc0HkKww8XsP47UnfO1I6OE4L4
5B/UPHag/msfTjBZgaXd0wM/XEsiR1xNCBHjnZJt0TaKY61sapomG5gh6FdNCYuU
d4FhbS2Yk+sgbhBKMD55fPCaFJGII9OummjHlR0TTpMjR5hMuJ7tk0rEIJmo2pDk
A/HOnqd4YKMW2F0z7GmHGDDLZuNE5QJ4svAAooRAU27W/4Hsfb4gcZhpR5nhcLRF
NvsW2onIgMjg3nY/P40o3SMm7A9QyIpGq1kZz0fkJZfwNb+9WMuglQz1c0UagXWA
wUWfClyCagMWV3PDREp4p350Anjtgc9OQWEjWJMAjDiSfQxUm9+W18rAYy9nR2NG
+s0xCkb68nxtl/NB6WiZJW6sibl7yH5MwBdkOfEVWulV2SpCW8rUDOao5AHWwbIq
U8yp42LnKxozxJ26YaxGRgrgxyUh1+mLC92lMduZMGG/KHzdjrovXdJZVxAiobuD
FOfnp4H6U7QZq3yT9ktW8J8a0dWmhgAZDLDF2+5NvPJ3Yo+3YfLlejY3F2j1HwHH
2CZkbpYw8kLY2OWK/VaRYZQeZWvyASh+2RvNfhMef2oxnipexP7zmzj1KupladZl
8vBFrAMF1Dk6QkKdXKgHq2Ax/usQLicIviSSNPhWamWdv3tcLRth9cqDBZysUUb0
OCRLak4RdV4YVRyVBUluOtAo0kJs5q2AB2xxP7RF/IK2VX/U/9+as4B6Bm551pXN
daFaezkdg4EB4DgIuN1mXxp8Bp4/g0xo14pdBjWYsixa4TYDQ9dJkiAE9zLgiOVk
UPApw7oL3uZRGLEbMf6pF2PyVXPWydM0gLNnlxqRazG4QfsCtBEeQmv/A3DL/hsu
PnTUsXuWNG9lmWL85rFsUXkrioqgk9cEBn02DTouwVuZuehQX9e7W9JsPAAzVsKH
wB7mPCjJgMzbZjA9TIe46OpT58qT49EDrT0SvCwxDNDwBpNzyPFZvpiEfLiql6ee
Au+0AoR5Qwsv3JDNF/zd+ZqrL30l7WmoMx4EuBHRFEtg7LdOn+Pgq+ticxoqrXcv
gm842aR91fFPaWCOn2jvk2VdQON/AUfKw0L75URTrlV/p80m7ou2gvt6Xc0O9CrV
sK85R4d7diBhG0vxL2GXR6lvONU2yowkLotdAOJ1CBxU8FwoP858njHWD2ODhkHr
9aDNG1CBVRIgjc9QktXiLVGFfVXLZrTVEvUskCtjoKMJ4G0aQgmnIqKlqKDPWnNN
07flsaXXu89tJDmqdaGa3Jy5uYzVtud0naYikm3SBu5mIVCq0XIzZ7TJT7d1Xph0
+gFGNJ2PUjmenvCLQngdHk7eiV0/p0AGtfwBXB+3D21+1TZt65lXZ0fWHoWBLC9f
sHBWD2CDp6lZK4wmdQh8k5cotb99LikFQyNG5n9EyY74VluRt7LdxUqBFjbJPRiP
C+k8UYXfBOnecdQmwlHySFagqmvPy7g2BLbrDCRmqBZIHiheUhHXjmDGgHJ8zwEk
OXhU64BCV+EEoPkqQYpF3tlKF/XxBBEazR6te9+kXZegdsl1Ypi7O10/0M7Hf1iw
HoiArcyprT50+1D+pO0xI80oF4HbcCoV1SHQIKfkg/2lEgbEOA5P1VZnYI8pHPfA
wmcjrCCgQdJQVDv4iXtF0A/ImiXXPwadJShTN9bC+vcyj2CZsMxCpKAyYZtSiJUm
XkFbzHflAnzDhs8ewFY+mwTV2KlOlg82kBOksNximVTccS5+DlKKUGATI2kjsZLh
HzhQcM+wy02JLNtefkOmLKj3YacH6tovZQhID1SsFyCRY5nvQTDvACVCAaysISnO
BUForcteJK+F+BRdvW9WGjXKZvWm/L0CJu2eaasi5PUhXbqxavQPrWzgpZDU5OkS
EJVYYi1l9PpnpH3yBxCbuXFJz7l3SNLQG2jfdKocryaxo7VkWxh6i5N3DdgthmN7
M4M8lSKksRVzW5jYnhmgMQVlp72W4vu6OIiMQf50nQU0wGqY6lBpmsx/MxIcZegb
eRHRVsIdVQXmRITs9wIytNg06oYpT04cMJejTfa5GeRBdyHy+YzG16dRNuU2Wj7g
CIAOuIhy9orIt6CAADbzSN3pIp1AgHkqvkmridkLoSo9iMl/OoyCxTppz9cE4+3P
/CQVO242ym7Z6RuKnkyiL+oXyaS37SzFcpKjGNT9UVZ5G+wsznf8WjCpsqXGcQhT
P5Iger4xBx2GG+JLlaQ4zTb7RrwYsJYJtXhTJ3JwYxY4r86LPwaSiHYt79+nOv4c
YRF6vJHARBjUorwTDHz7oQIvH6oOccCYlCfRSXOwg8g6rXz3j3gPRoSWczCKMYC2
N3V8V6Bj7t7sgJ1Q1E0jcq2NUPNQq61z/oGhiq/41ibsth80Y0/vL9BsaCYjt/yh
BcGPQaQDBxdRkSV7sU5RqzQor1IM6+HXQtXBGVm1yVKEUUk4kkGn1LZnyxC3fG5Q
YcGXRXstyo2Ts4UP5/eyK3CGBWIvmbzPTSQZJGqdRGymt5g0JwUw9v8h9XWpT4Lm
W3zL+S56ai3+m4/dzwyXQzruBIAd4HwaCP3koTJ99ypYxJQRUGS4RqjWsyxUCRsk
bbNBpVhRRwdqkz3wLmd893Wh+KKJ7PIOdqn64/oweIi7gC4oEMNntIGX1+obesEN
I9pfGMzxpgmuqPgBz1f9AAOht4zJR15WXVv3Rek5Of5Q8p7U/6jxOpf4WitNvzpo
mPosbN01/0NbxZbSRGtehFO133Zr4Kjj47SltKDxaoWyV/85f1ZmiKc/r/KTKvbh
/dg4JGhzcYjGLl+xPKCmDY9F9jDK0JcZGEdVAt+E+mNylLILtD2hl/jV6ZThZ2cM
uHKiom2r4upeBDw2rY6e8iAcOO/yw4cgw7smlPB6TRFG/wuM5hWQH3v4k5ACxqCf
UKYmxM4mkjBGIPTGGNQ1MT4UtNueO9ltm2c/FhTHKT1c47WbAaDPYgAf82UEKPj+
Czf2v4YepU9k898e8/01e+eQGYjpPg6wmp956PKWAINcKbMVvsOh3Qwu83ko8T5B
MUQ/hbjcCv1KJchOkXKjyRLYYsitNajVMfEEldFr7w+GGHmOFUnvzvvtCpZwJIAb
LmKUQZQDgKaQNwt0ziG2ztEilqwQ7y6d8V1LXGBF3UgpieWvpLr7zz718hq/Q3DO
xd3TkD+5UCTHN7EbgQimS7QRXWQ4X+95Epiwer+BQ1E2o9d5akBi9Bba941bLYt1
1L4CvolR8ywnhSej7jBEhukzpVUtPcIVyI0GO+ZsxlFWaWEtsPFFywObyY542aR9
0Lp/Flsin7h/41HtMJdq3/esjI6XinlQH9duflspnGIKFpkVlIzqhY0QPUlBV6K/
7d8JUpW0ZDQAaLhPFRxZaZ4JYk+Lp/KJBm8yDoAaiM0N7jBblofwz0Q6lxoPFpTn
gcG4Q7VCt2F6r+eVXH9j6V2zKGsurcw2Hc/P/jKTMXFpZOTWer9B1ze0eEhETpdr
FG/YjFHH4j6VCn4GVpQiOB/cneUUNTnvioJ80iJjr1DTZ5A/wpUhuqSkeoBe6b8z
CmxSNn1KV3Zep1PCf/CoYbRZCMm9VJPFwNcf+RWud+2A7B0oX3d6e9ZQFCh0fFSv
7U3L5Y3Ndt/KULPKq21nPj7KQBJ7UZO31GnJddovMtMja8oTXlru8Ad1o+eLOOZe
00ya7KwR0Ke6VSIfohz5WTcRDNno9dqtuPeY6wYmMB3zwIZXbu9LM4+UR7s0+nOn
27hoxOJPO8h02ZjBedLRfeGHXAWdQe9T7LbBq3Wx1r6cJ0akyET2Vz99cSVkG7m2
Ib03/cI+PWc3PVFh9hb5Nc2po57DPS9/qVC+PXoGpMemDdJAEp0UvnEgdcIo1r2n
Sk99FVOSLFRBgoRgRVIG2zA5UICybtnyKnwFoNAotiuLBDGRVr6pAOj4JMgwIbJ6
8BNF5EcOSVRgL5r1kHpCqvJ7nIGil7dNRD7lj8mEp47DmO+4GjRbjkCupX4qUVyS
yGfvq72IeZUcOdkS//Naq6t1+tHFQ8SqHIe3VXsPVodfd3EG3P8zLeMrxE8puWTH
0WCaka/0dZvgSzIWxdkQO9L7trDTrN+kJ8WHhOAM9ACR+ohIImJrnig1/1DdmMDZ
ud8ykHKgAYF7UHXoj4jmm19TU/GlMpxsWNeUqUf3uyjFQZPk8SNSL9LhQWJA/X7X
NRT/yGU3QTOasX00g4u/+2WE6Rtx8z1Jb2pDYJpZ0IYHO2Y0jmYRV3hNFwKIRr3X
mdqiLYtky9TM6f+6h70r3qmzRA5L4iBfhLH4zplgayHQMTM/GZGx5sVG2yt9O0oy
0obBuIxaJxXiOrCOMpjYIB26+51Ux4ZS5063oyDvdFjC4gSka/mhK+Qho13WrOZX
d/NUq65Z4vDFPf4FiVvuwuTCNqkdEVBLWsgJ2cEk1ahrZhzuV9sOKdU+ESkOMGX0
xqvUvIExYAnzQNowmVfTnyRwqEoXjjZVtp3qcHjPwJ7BotVqdrxfa1MigyGcrPBZ
UysNk279XnNnt8IzJp4ZJ2opOBuSjszfTpdsmNYuKJhXGe3jegbDRHsonntMDrBb
meFyy14mQs3yE37D6dqa4gRmbpGpOJStUoJ9fna1tWM4jm0WDapKFPod5SszUsI1
N6644uUVjf+wiCWOkvSnv3OZ3vVujapvVzit6XyxqaqDsDp1mRWJJ0hCHa39Nyua
KTnjh4NkAqz/Zoyw7yG7O7d3+2UmPfmxvB9eGymiJ26C3QfuB/0QVi0RE9WRu81s
IeyE90zqY5gQIvoE4FmT8ffxE/gstoXDm5vDbh5wrTwncqbtFMcq3M3Ft/Cbi6Z5
k3vnP/hFhFxA6Qe8ojDioqsMojK4M6JFMyRXORJMbzMVs/pv8n+qlbdibJxgrE7u
SlnBYxbrutEGz0+DWtNoZTYi9e96Hq4O0bUZeTKaTRiYgs2/3FQIqzSJL940a22z
sjaW2QUOb5QwJQXDo40lYhuTWMF7KsIhzfl3lXymf6VKYVvISwFYsEBQYg7fCscZ
U2JYejhVVYTckhyykyPqyoiCeOnnHTleCFv1FNzkFVXVh/khbjrEmNqarP85PR6Y
ctp6YqPXF1pdd3NiS3hzfLw+F+5tJeOr2Gqvhea8HeeVMZ106l3OjoMjJM9LH4WB
FWPG1it5xzDCangjk6N25MUzmkahkb+NnM831WtHC2dfVWnyTo1T5IcXoongg1IP
0DRpD1dhOlf172kGdvU6ErqQojeN/Xvl84zzxrTs6Q1CORCMGE4XWku1DU5sNxGD
2Svv7myfnFKMGVg0h+kWdWJI6DPkilqC4pbzYYHS1R1Dt2lBTXOH1q5fw8dMW9yN
tvRexxWJsBbhHC31fuHYHsZ8Rne5V9ta0WzHs8HPIlRSTFwes9dF6thA8tlVNYcf
18jfXPkJcsx9/dQPfiY5KQspC3zE0LmZ+tA0qSBtXIAI96skM3hpaULZkmIQFlvF
prodqil4JKfGiNldbBE7wurYYX2mUWE+EUW6iP7IaUHPkxvGYuZtNQtyoYjaJLBv
hl0fGPlZutHQZVxGuY9Tg3onOrAbBXK7JKy36cegEhtAeiIbylYR2uXmtOvFR6kQ
qsTIy1yq+mCnLvnDUkdhIXRDL/U+QvSbBPw2En7RSKKFGRPezOc59B6jyhifayDj
l1jHNGJtS3t+hlDxWdIlkIlamI9Cb8Q1yedXcN5kffOp3mfb3eXlhZ7T6wcEDnrE
OHoMhEG8Imh2CrjZ1q57DB1dZSceI1FYYBGPiVUhvM+4Vd867jDNr9b4DAJ1H/li
FpxOqKdvMPW18b1f+5Hs9n7WD6UuABOrpqhr7SoqHYZL0r8TcBT9uoR7behlRS5I
FZWlO5TWG0maHRhn/CZk2B80bUQMsMdPoqQmQ0MlHEJR+lSsqCBRMY7pyl8xvWvT
lW5KnSH1TVYALN5LJPG7AlTsTcnu1585HNCygWKdUI/JOzwwQ+ZvC3QTU7dHC61w
PvKYS61IB9I73hZ1em1KItfmOku1+nApY9MBahXw1wc2r/HEZW3bVUA9fTBl9hQR
fBNhkCt6q750OjZvRLVxLzs8Al7MoWXpiqPo+iXntdwGLxREeHiS/zU2C5ExdQqI
jV6CBJ9lARX4o/3yF3ymAXKCcRR3k/zt6q8HzKkqKGUzzR4MSiTWJpnU01MryF9p
DXfnZYfxpHHga7pIkc5J7ji0CPVg+OEkB5QpV6w/YCZYvjPtWwTGOg8YO0q13cAK
APdp3bKUQJ0nxIWHyjmVJr2nB3c2cfbypkX7Rzg4Zrd5e5gsNS+m7bPTAeFBONOn
Tg6FIeXgw3nXOAafCT4Rx0PkBdZKjV1J3Hm8FVtghK0Xsr9+FVafTjc6QaV/WUfE
ZqOEcUPW7ipMJQQX0hxWc2gyq2PWWDX83nn1oCD2jXTxhavayqMWwW8O2LvWf8JD
2PMWbWgXoSRfF3/P+vymnwLBENOmNlvTOBzp0qrp46JY1ge+Tp0m+AiuWoisdSe7
iLXvSEZ+Dz1h+tkEW9M7c9bgcyeZKru5ojMQfsH74M1F47DusxYBPYdaOleTEzao
Bi8keLGuXN3Qp/U9PkXf1+/adPS3mvD4YlLgBCjpMcjc5nEkGVBWVmZueM9ti81G
gkt07gasE4p5XqYjz4C0adVEAY9b4HxZVeUMH3HSINQX7gFu7zQOU86m/mZj7TLx
3sRGtsUrUo98y1cQuD/jf+8ntmX61Tg/9RWpcyj35ybzjv0BT9YwcvzVPIrp0ymc
UsO/UkwQ9gKCZBWcG6Em00Ypw1AE+UpD9adcqMtnP+e1eQvu7UVdjR7VzCUDD9Wu
LQaru+BYXVIHNHNVfmeq6RAYXULF7h+OwHNSMzrRhWL1yF+8yD5ehSELb5IGNXKf
2o8ZS6gr0z3mxVfGe6dfDmi04SdWxs0NhJiA8WUde9KDccVfoQSkhPDJosfOG1Fc
qsLaOwJUb7YxpcLm+xuqttzUEX/jr3th0BYJGyIfLNdI77Rav3Td20fy20eO8vEg
gaEbH9u8NfmKZum9/yN4kVzEsQ4uJG1YQgn8qkrFo/Lon15vcdGwMGn/0dA0Hcqc
Wy/bCDTH1kUEoEUf99mVk19YVgsy4tl0UxwR4Py6GM0lBwcC8clqHZTL5WB1zLel
res+JZsVLpC8RUIqFHo65wm6ioV4jw6FN/Cl07d8s9Zd8kDzQNVAUeJgE4IXnxQx
S+P1c1ea+fLDiv/rIJPRsMaAA1LxZwlTpnQJc0FGyDu4qOHvoIbCeOl19eTIpyd4
4qlEGIjU0AzKp86WEENT2mOXLiexinrFbMqclnChWEQZcrixuusp2nCPOmpMhnwN
fnR+iCUl/24F2/5vkLoQtGASgl4p09muiPq0bKzrfCI/lT/t7j1mC9z+h/wM88lH
8PPlrXYWsV++lts4nRFzI7W9LI+vpdQ3DItCEncm9gE6Iwav4HThtQadnDoR/z0D
+WHJiT4qriMuO2mriD2GBi8zwmmTeqKeeXEBJKBjZMhrS0b1BRC394iZzcRD4Qh+
BObGnoyVBTbbToAcmADltgA+YWEWhi9fvC7MyOmiEOwBLiLyF0j04Po40F8EBAi8
JVZczaVTyduJAtdfhjBB59uqRo9K5os6/jKQvlq15AjY7qanz6+lXjAKaAt1RnXS
zlHHZ/orx44aEV1wNQImx6Edi/ZswixVz6y2jwbWzgF7Q74hf5wD5to2iDOSSsz0
a/EN290Er5vXGhZbC+n7YP7i2XJ9xaHq4SfSlLDZFeVfGjmX5Al0WCSjj5OMtEr+
GCwTxBWCldmhF8jGdDSYuj49rySq3pwpdfeir0WGFLISJRHybzxHzS0Ixxs36SYF
+dr56dPS/1PbXhy1WxMwJdAcRIe4UimaMDWYqud2SW2CW6ztNoALGU3eV2J/Hy3j
FQ7r5VU/MCypuEN2WGRmThJjvFBeNImAcCPYFrw8qK5YX1tsvL0K2uBYJh+oPNoF
ygtgAOyHF6KS74HsNLAJxSj1oLxOpVVJnJmvZIBPqV4kShozkv9ZJnYbmvWB50eK
DRvdNi6+yrQH53eQiX+r4cK36AZxXAYHAkFOi5FsN6OT7vI/PLj2dDmjhO2VNLOs
ondJdYiq3NxTK9qS1eKOLw172BTrpW6xWHZmVsFROT6ttHlwxXzIg7znLDgCEGRV
8nMCfYfXUhmLhmrMzqAu2t6AAYPeAaKG6UrOARjH7gisjlkZkeEjvHthf1rqtW0v
/wf+xFSMqKMPbw+Z7KeQrCnhmAmFP4jcCp6i+yEakDnhi6Iiq2jLeiCCwrPG/fqh
AqVgJ6kh38mD1UaDdVgQ4uGekdFBrPPlKkdNF2wQbQ+jlzVVtTjTrmuKQZ9+Ue35
e9pJtLDoH5GoY8eTDkq+0fNGEuLH9GNbaBeltgsZ5dUHUzmFfcpVnkR95oN5VDy6
x+wQ4pp9Z28n1wpOVC1HmPpMHpJFAgIJpoyCAiMa/ykoXIDca+DmJS5zlsBdRpQe
TZiCP402dgCvT2Z39yxSql0Juf+og4gCYrd5tP+NFv8ZpnlQvyupegrpUJUbBAwn
ZWAg2EGxDnE6VJhfBfKwWqrNfMhpTvFdrT532NvBkeofHh3kIo4PPeyPYQN3Lcas
uJO7m3ocCLKn0xXDslMJyoVljYJypP2LBJIuOfATdnDGcgrnXjYhhccEbv0amQos
SJK0TC/N38eFRS6HNcRu2GEXC02Bdm9jcQmQ/fbHPY/PmkAjOMbVCuhMq8+2NSt6
QGgI4BYfwiu1+7CTX+UIP1E1/SYdZylhQbDhN3yadBv+okNknX8hqyAWQ8H2F9SI
P7JGVIVhozfITFHg5ZplLWmoNdsMMErJ69GcMA4d8izdJijlp3yOrzQunatrYHRB
bOoRPf6kWHov/CQtwYlKG1dqTQ1kBagCIdNEnkGinsb+M8MGpXiCFrVfIQoBVmht
eHe/ugBhsAN6r5HY1tclKXMarBnktyv1Z2bq2N/omfDgpugsKyleLGBJBSYKovUI
JOYDsUY1q75vYHozyeepqJdhofXQBlIOtbNS3KqYlIpYOhfLq/I2Osx9CX2qZsSR
u+Wqhq+/XbTMevsl7YS8Ncv9CDNyvExpq816rlDQ8MrIylmzLoee2BRk+0ok3/sj
huJtjrgYcD+n0jAxIKOo4SCDs772iyoo+iWgAJOhMzomKLQNCbXp/ZQ1T1/34YlO
Mz8n54+QuPVlIBEUx1jEbjkMrXVj4VwfVkGhrD7dYzVeNFmgo2vlTf9lEDX1xa/b
18zerwKdaTs/nDjWVEtaPYXPkoXC9nBAeTYWytjzRSwGVYp4JE/1hFCu/CtRtoJk
HwISkZig1fzaOMRaoVzte1GeBfrNOG3oW/p0XkUva5gPYS149T+iKJVx7F0hNmLL
qn3HHBaKFQRbMzxtkPAOj5FZPAHhjqSo6FLM1tY0o0VZJqKwS60Z5bKlbBADlRvV
TPDsqZL4Q8DeGusHLz6lmCGyU7Fb8NWOLvXKUmFiOaaf/LH6WJPplaNJBRyLcdgN
NqYn8onwUShvLKxMmasF0uX5o8Ce85wK3H8Jg+6MRUK+BhmTUOpM6vq3MIiyRzT6
E4LLNO4yF5tnw1mt9/cAqZhzJZjBTJuGlF+Pf4hKNySqlRrV5mIkp0ueFJc4u+l8
CHB/BUO/+hV6Y5dd0D9t8acFIj10SQ/6upsrWQX59FZXPETeQBXyfVVWopeaSJz5
fpcAxmhfGDikiWs1nXGGGnKbH9ct9EjJKDd1zHPQ6nc4SPIwhkwsxajyX6wUspC0
3cPSnP8DfYmWi0i4N0U6bhEZldr5q/DLWD/RyxkVYrTJ/DQHHXBMEUTOqkcNPB6V
mpdxCEmRQI+cIyBPUNVzCw1rXT7Mv/BlEX8Ll+xAxgIHcrBKEIMJjnXhQudwN379
KwyMsHECQGi9TmwpYCWumJJEA7phsxTJ/gPt6H/xxvyuQ2kgULuHz+spTvnEcLjM
orj2SWTj9svcJGISv1TXE/P1EMKd7Ncd9ReH8iIDWCIWiKYevihIqdXO1RPcd8g/
B2fWa3dXO5kyJshqMqyD18EOLC0xAbXIAHtLYaOEp5gCAOBBr2dYNj4c1r5ce/Re
RbCcNP7paJE9PX8UiL+/MM7JJ6pJXG+h3f2zy6CKKjWYVM6gXFFgpixzkagJeL2L
Z5iKsh6CBM17zDyrCng+euqq9aSJD/RrQHr42W6rNT0dMD01bME7Rrtnu241q3Kk
Htc+hbJZjgvNTIguISpK/jPb9FnQtTUbSQs1f0T7A/Xbxw0nCIR/CfUHmPOuEi0F
radITp1HaF2LjgnYwJl/2rrGgI1J/SNUDQBQSlPQGZDFNwlkreeAudolrH3q1L3r
QGVsMZVk9wrR9Mby6CzXTzDsxhcjypMALo5I8+MdiYtiaKzvBaGbecv4tGelNrE9
ZeHmXjpfmjHSt1Ew1V88fz2conLkbIVi2tBj1/iIfxP51DegRV1BAjkAz1gm6upA
CrdXk6tpLLKG6X83EzRJhHI1WBgVca7wUxwuqJHXkKFPUj/wjGDuPchi5np/dKN7
xoDXByxLPoJqFqTViAENyiov/YTnne8vV4qGSASC54UFSkmKTOERTsQBYq/t0AJJ
OaxJOXxIjxzZKQTM+SUF1H9K1LheRXcqv77iWYXyCmuW8VDZsTZnctKU+FTb711e
UIsnIRNXit0MV+KTkoMgAOgG/zBIdkokejHN6YONLQvzFz8AV85begZakKfJdGK0
IA/thCbg+xsayxszLCSfU0vSTrLKqZDONvA8nhF0RFZzyjMoLqyoGgPisGC5i7PA
tm8TsKuUYUMa1gfYRu4FE/PraDhkjd0KcbfbMCkVkXZpNOIbhecMRx+Dnl3xwDu9
JCi9UB3MkoCesfio7O8b4JNWI9xtLZ9RZyC+8gUXqNPKRFB01/A8vbuJWHdaaZVa
/SzzC2TBzIMhut60NRkkOOcSSmjpQmO0Sh65QQCMvPB84UbtBO273oYs0xh0nZrH
6FCtW2C+ix9XqovetoXIbqrGN356RqiB7JjjiXm3HXc6D8OD5RgLlwJx0ichp57q
nc6CSmhKmjRKubgw7WujcfHrjq8rVTx+XAi2YPjyOI9yxd116TxTZ0JadVxSprMS
fuoFN0nCQEMkHCXGpLU1bwv41Y8s4xyZminilWN6PW5/kTO1n9NIQaTCWabixHMn
0Wun7m8JR7wA20MtTLfTvkRha/4NgOnGvL4zrxiIX7V4dIoHhRnCVm+ec5rmHTax
r9rl7+pyYiW1O2PhSqYABFzrS/b89xroJkIEoTd8zc3p1eTE5Ud6RPLeANdxQUM8
R/rG1P4zQdxuwTYZkoesplvwoEE2BUzT3tOz1AGXihHmd7hgENnCzD3+FIBz7pck
qFnqBRBxkBulEJGyqbnDtY7rjEf/wGufTRJuyvEkGb0GeVnx/V3q4NLDD+krewlA
9sLKby7KMI7sAXARuVkn8A99atXeb7dmSDnghEwnAyiCSLFC2yNIGCeW2D2HylxW
072CRtZWthY7ZuD01AJYJK6LwAbmLbdhVbbpQ8mzDnWvmv1K3cnho1k6o2d3lp/W
9+o+e4oNqCAybIzY1fq36tJsZ8bNHIyIxuZy7IcywdtdQIS6RSssAgsvfABzCarV
Ml4TwaEcx27t3PoSKSfJVc+3Q+Z/MNg6OXDpi+Yl4Y3uY2s62wT1E7wsGqZADkoT
LwW/ZxYnSBS9eQT97cc1c+RHQG5ZpQiyTPW7E4AafFry/tIVsxSeB87SHwokYlhk
YbTUNfkE6Do5T1R8XUirXKyx2riPteRtooXkAhxxkmN3Sb9Wys/ACCnYJdLuzizc
SHSfHfPrtlqMm26M311Y5DnGh+O1HNP+jp4SpfeN16khk1IqSnx5RG4lkV2ZZxA3
KhwOV7lBjg0PaD2mA70UulsyJhMsaeSvwwKUdEYPulvoXgGfgOB/A56N88m4dr8m
nOT1rXrj5qrdA0NeD9NOODrGCCMi36FrXx7NFvjtd/4F/szV5rgaDBhFOjQz4VDs
SL6TZrRKUahyTey1YqETu5V/tijU9/W+jPn2xnm6fFzOvQi0R5p6j5mLsyTZRQ8/
utfeJu6TNoycdJPpCja7zWp4qGnICQdJlUG5HmTXbYvADSzznNs5bY6M3lnZKLai
onblr4RFxPLAvjf/CEQGts8LDCLI+p914KItiCouLwZSzo8pifV8PGcEC0gp6Pui
Rr6gX0ELML7IkJkKb+s/mvox5nqUuDUDsfdIchYw6kNjdbXrkdEdjGIhtBqkgKEt
9N3QFyy9f7dc3OFROUmRSSZIx3cqpuNkZuYG4LYFKJTwJYtCrzy7R+8jgrHuuIig
mvXRrO0b5B7kZBpH+8Piir1mTZKpF/vB4tAN5x7WOrDJsZ0JIZ2kE5sizLamuA31
5/mAauF5qxJwze7iKx+Idy+9RswuwFCEsKSrHc+YhYCxHmtqeIBkNVJJM1yHnyGm
ep2tnB1TRm26TaYlDtZNBB3S4Zvd3uejyX2RkmFdqkmylg4ytyEZPoULZZmJp1RT
4+Ff/J0r+kIjxQ6lSETixCRPOu6QDSMzrkGFK3Azkq3D69pJ70jKfz1B5dawxIIq
TwHDis8q3ySTpmNXgKrw0e1mdVDD1Pl5KZk36ER/F2etTElo7sYs4Bpi66n9evhe
+Ut5eyf28QjgueA0bxgEIrxHg8aef0Fn4ruwxvezXb6PxL4AE52kdT7XUMqg+2Ys
pgPv4sOYvxgCLQZErLUkNyPlOowvmKKsSbDwJJ823u9f0DbL3VaA2+Yv9AKKiOGM
41F/mxVDLRdUTsaBetlA5DkCiqhoabn37fWDKlWVnhRWjQETudS30Xwafi/Z7qV2
IjkSykYEaIovbdGiRXY51nN9CJEfP18cj6OzRWiN8gFTvxNaXxfh+FUkcmQwYrfH
kf41VkWM+jIoPMHDtMuOy2MhgxkCfUIFpI5LgeiCxzKZ6/a2wuY6E9tRUopd7ScB
GJbwaLK6jSHYl5MtZO65CCsiI+gNquEk3OmGD1eI/LfMkhBvYST1vKk9f2N9TfO7
/BMAOre1l8jQ8wV4Wmh5V4MeRfwdNOKN7FaR5m6gcZ0LUxzMDSoiOH7CnaHRrcRR
eM+RWmgGGXjm1PDC2AxLj/vb2fMajKp7AJGTPsxVQADgUHS3TDOEh/kOHAfbKqIL
hWOXZUbjaNofo0uQxqpCayM5gMtz9rWip0crsnjkHoYEPWxZXTr1sxErl9apHl/d
lEkATAWT5wfJYgQowq518Pfon3Wn41WsQfvDjv2NM8VvB4e94Dpsv+JXhrxm4G1b
yPNPj3bCib69PmsdAcNblwXWoBl37top38bw4g8sYaIqv5vmpnLXceOeNaabzR5E
3QXMTPqBxCqWpJhgsKKqGDcDPSendkNhvWjlJ9BUN1vlKzgG+UkG0z4zow5J/+of
9+Wc/yVZ+bkooMW9H5nDPxw5FWvuuU5WQX+bQ3zh91F9ofSNzcrROOBYMtFV7lF1
2gQ43YzYcANK98+kdiKY6wUCN+lfSvdtFtTQazHk4A9/+0D8OgpOtEiP04scAM5f
GGbVnEJnBLMIu3qtIjjI6t691ny9GOts6YzUfxiSrZpb2kpuShef6NdK35hmNQjb
kp65yZDVZjqe9J/jzfCz928geyfLavDNxZDkOnbOPoFQEKWK0mztv1mrQiy242aT
rZmbDMC2GUuVCQNXDAWUsGGSnYLr2m91fqmgaoSejT+S5yzd7O/lztvA4g8NL3uh
2aK0kZx1p5NG8MxvJFSuRVNLKdeDaVbGXV0m6DuMx33fZ9sEnguqxsN42jIWn5M9
MOEHGyekTnSQqIn12Rp72/td/HCH0EqmljnryvTM8Bx079Y17+N+0VqA93L+nrdk
IQ/h3hihzJqQwF8AMTHs2cxEtAsWGBO2TViRAbwaN0OrLVP6/Y51CUsjGFBmClNd
RBdlECkmkzH7aCAi1E86kTyB/jFHfHQ4p5xWRYP88tyYw/q02SD6G6fuOe8euTXq
I7ZD4gnwM8l7sY5Q6zsBcioV6+prY/ecjapstXJGLdsxjIssaL8taA1ne3JD4vo6
r/6uwBjV3wzDUNI8w62+v/k/Z026Wt1G7rGwzD4M4U2S5WoxGUhG6HFTyiT1VLJW
1xRr5UTnyzjP3DbTH0nWOxcETI//OAsqsk0u6kfh/kKKmm9+i5yWFPSuC9RVbHrt
zPePEtiUJ0LumaYxe1L1QoKbu4RQHZQMVx51TG+izZuRsc9Ch4DnTXdOINTU2zHP
RWmwUrljIonIxinqQxxaEX+ffYcB/S6wrhverLl96PCxBZv0V6bwjnTDvNzy1TFV
VguNWlQFyPiWLz2xqhigkucmA9s12P227tXVXjf+/S7WHzDuVyRFf59b9ZD55hQ1
r23d0DByIVI2Tl/snKqtSa40nrmbcXrE6z/+4K1MqeS1v1VpdbW5n3UO8P+8t2lt
n0FxIqaK+ge+KVvdg2AYYoRtU9qeb1aBNLtYNnp3868QgmT5gPS2P4vwQeAPjqab
zYxxTnVIeRht1zeN2Xwem3PF8l+tpPZG+APGRhnRBwAv32Lu/zjJDKnrddQ3RZoP
+HA+YoNU/TJSrTOhAHQr+hVOm2kro3nam/7zgJNWtQj0g3BMiMnsi6Z68iepwRt0
qL3i/IbAMjVRNBAiKBRH6TA14MermSU7upZ9KWpW5RN+I5WeLUIZLnudc6DunrB/
PA+vI0p6zqi443LoocT+aPBY/SJr212QRSQbL5Xnis6zwwT8bwLLJLxzhAQNUrpD
tWyg7bzhOPw9ZFuN0+Bez6kVpc1x3bZOEmS06TkaA5CiViBZm/9vicxMIWJ0Xi03
DBlZi24asTN7LIBHRuOoEQI3+3ZxTD8jveymlQ0A/4L8pU+yIGYu9ghfR+aV6IoE
ENp/K6ehrtjBd9lG+FlNn8sHrh1olJfkLvoH3MqCT9zUWyHCYjNXpno50qDA8+ug
iwW8fGvaP6v1Qyf0y5gcQMNLtEmOl19+aCqvg+pcG+PjQCjg2VFS/CfyLxhTay2p
um3/cHMEPz5mB/CShZ7eVrR7I7px7rEmZcGlayYkFWGWs4lHQyyztIFWyDJI3ZaG
fHrHqAX3ZiwmCOEkFyV1zYSI6WbMnjL5M5ca5xXfF+HztgN8FVb0twhqLWPcKpGa
1nbUaAxpTbnWguJ02qYzMwwyM+t6axgUwbDyuvS2qoYTtmSmTLOPIuw6SI6LWFmH
xIJcBWaNU1sGWc+Gglj6ScToKQDJc93R2GPOHLWTn6zQdm1X4ja6PReu43dmqGYM
roibJTfXwXRbP7Jlhty/GYB6QexcWRVOe+txsRxTViy11oMyw0DI6wC7COy+mrgM
vi/k17+uqqZpkBkQuXelUEovSH/2YSOBBnH2LJ6hLQ+jxMfWMHcshLh6rdD7wSZ+
W2eEFqw/9BmLxyKFjajCsCf5fJKfCXHtzCzheKHMCBT2q0gIcKU+6sU9IudwQ7cH
r5B5cAKatjcv4CHJE4hH24FjH0iakaFfsIXywrKk6GT1zk5jOCHLqxWL7WzyXHJh
6OMHMjEUZ7LKhqlL0iCVx1wPlybKajd5qKdHQqlJyVQ64oEoVCu1aXfd4dG8yG/c
4eVFr7OL2ucgMtlBFBZ2N9ycs4oK/HMNcjiA9bP8Btqx0i/KhZIfn25hmMRzBMsi
/flwNJ1+xUipTLeKv8YIoRXMI3fCoG5CRnbuIyWDCo79N/krJ1Ibx8xCdyAnVdm+
C5Nq7Mq2yynIqz0DvFuJvDpdEAO2NlkLci0FAYyiWXcC6JmjPcbK1xcq/lMdQDXO
ddZtrIW+hEdAZNUNxrrhTuFelxEYOtSLurImrNG3nDwYz9/eI53oBSch8zUIrYbs
zJ9vMUVo5WyvcGlTJFlXW8dmR6XaflXjO8NGc2iS3NSFMr8mX/1zdo2gcmGOHuVV
wVyEe/Sg0AOX3B+QtoC/OxG9SQKHtAwgqoJIERoVTWjDHjpIfLKasQgh1V4aOpK6
tYVLu18jtyfWHkw8+RSsmAcj91WOpbTXnUHWNgIF87bdPjipPEIrbTcEhTWa4tVe
XWg1nLRBkjx+2ddHCgHcXQJCVeb3X9u8Abjl7EIGfciITs+3arI+V6e2mSi48wzt
/dHgSzWnwIE4MI61VC9TTSc3PFfZ2t0tIBd/dKgM2EwcA3ehVmA8f5VDkhB9i2PR
LWrLgeJlqO4anNmaDmNhLuigMqZ1EtrCU2q3sxdone25CP9ZBZQJ1cIn/y57MNrr
HftcZsElE9Gy8A8ka568YwRvanvq2CR+uzdbb9AW6YZpicN8vCnyc8ccQGZ9GVMV
pUKUTY3oPO0tR/l/njyhWY5Cciz3tiuPzJMA8I/TQQSf0TSs+MirnBmSWZLbhWBK
5T156fPRM2933zhTh3vyg/2Q2nNn2IPB7UR7MWHAOIq3hTjNbhTvsz0QfUtJ9h7v
1I2XYHU9YyAn5I56TC4t+NmsrcwfW/iduZvunj6bMIDhhEcaYmlLhXDVI4hiJb9J
kzR6dQYIVKFFM7PKI8jZAMmsCROQe6MFRxpWVwdtn1BIwhHmz52N+BZmlTPY5zwn
yK3wdHql8o6XWJwuLQBggdv+Owg/h2HO6/yWon5tfYTa0Ni2MhomyWnYODfwKOP9
hyrHj8Gi/I6i51XR7XlUNdI6Ua2KTff110xg0xQnzbd1CYvdyrwuBc7v/Mz5xsEA
RgHS9HqDXeCUyKS3zn8iFUiAhDVXdnKVVTjPQy5EzJIUHcAVO6MxleufreNql3M0
/Px28Jy8KSn/7fP9YfMxLR8sGTvuSXiqUjtAqcxDBzKDB8v/aODAqBL5SN4ORaC+
D65UaA5krSYebSe8K90uJI9PAa93FrwEpf4n82FoVna+CZ4EyJOeOmzARp8czR1J
GeXXUIXNkJxQWQmKPj6jZJTO55FPIk22HqZgftBNVBBbCRYhD/RCFm8gbmfpKPIo
PpvlR89gfSAbG66jSaEZoyJRe9C4cDh2WsX3vGTtuwL8utUkc6CJfnb0O2raiFV3
L0y679Odq+ci2oOxRhEBKu+2jA9SlnUZdnlsKzikYjBkxo3D3n8f/Z+PCuc6efg4
NxdVHspZOGUmIICiU96PelDQryQguvF8Xi+8qjrSip314LJaBKOicRyDhnXaOE4g
86M0Hgq3waOgqF4NL+MCjsWSpyfOm+TiYHUEWFlEKzcYL8C/6o2PfGPrnWIm1DhM
2WtFHckpRJeFeOsreDZSM5JlbyApiPlTbNU1PR/xXCmAp7C6HOWZ7OOft9rlvWlT
JhS8jsBGQupWr7jL9uzxgvmCssETf13ODH9TZV81Jzz4Oor+ap1g/WVivHsh3wS/
Hy97BE69asPW5WYCRmN2S75RJt/NaqP2/dcCduo7woSTy164vty2+RAFqUeyyI/Y
457DIKk2furJ5ArdNHatTmBhpczYXJLo/49la9ncnw9/L40Nb4PdzTtLuKzuPw32
VVbRShTFUCROTPpQsStfdT3KecSF1ajv91OZuDyueEEaEqEVWT5JQr3jVSgL2WfD
IKYHQq/iaHV1MfedTFz/TGoWwDuM55GbiwTYuxRdi4QNBT1jMQtoZ8Yb9sxlvCAc
2d4y+NbtdForV/ZB7r08evIDIWNzyMccp/Upbu6SCCOyry6Z8DerEpNgPWO3qlnK
CL1SrXSXRb9/OEukMrM3o/g2Dh7Gw6eQpGl6/1SB154NZ3/cp/o1WWcn5uUdn0A5
WjpCOrsotNpuLFM0KzNLULWLrI1xaOGZ9Pd+NHykoosmAaMBRjpPB3uPDqLqFtDy
Q+NK2IAiqObHybEDgJsgQDcNju/ejhd5wLDP9XohwEODGiRp1dNCgvF0kEey4Q5z
Cr/VsYzGLD5pzFdBUMd7EwU9wm0DsjBFIDGoDCgL3+z0LOyFw4PWYVT6hf0v8Urb
GojgysU5OfZ2S/nEbDLDi+jYSKfP7/0sczNPI4vnagESYv9OzvbpdOgLxgiqTXux
hiYjqxypxvzx0Ct78CcIfBrFbXzetnIPAnTENEFoeKr107qEVohq/Un3DYJdE3Z/
I2i8wU45wg86f3THQoFoi4tcHYd58SVR+abRU7z/xHo55D3Luq+mRMC7BoWSJfLm
HDCj1f/o15rkCiIAgLHW734eE70kdS8rQrhira0TvD8wDTcRNsV4FlLFFRWDvRHj
Q/vEzw8MhQccgGxQZaaJIRVB1H/hwRuVCOb8KUzh4SqhVXxzpM+napLkHE7mw8Ea
YMll82bfI71+uW+78dAFXgXbyfF4rsJdrRMXLwdtZpqH2U4E1JEHImoGi8GKP51Q
nhN8Km7tNc7vD4kMnU1C2h7eHuq2ng5JsVHBM9NX1A52lCBXIJO3A+h4oUd/Dm1Z
WxjINzYiPvYwFwmAp+OR4acnWo+2d4RmggSUyJqH3FiCPhaYlIZIz0D3AhTsJHNE
4+O4Q6mAeUHgCpGAHwSM2ovQrNjltHOHjFey/EvRJoTyV6OWScjhxkxOMYs75ODI
8yH23wAEYuma1ImahkQyrRPoxqjsM8VZkmMbgTPyj1X22jSMNaY042WNvNmXJlwF
I+UYzcDomGLiynDuv28R42bD4YyzGh8rmIaAMH9GvV4d9lzEzltKuWYbEChuSuqS
FUljEbOfejvr4YND6Mj8imZw+n75k/yiGQnL17mEfjm0mQmA8a3gv6By4VAUK/P2
/1HrgEWdaaXgx4xkd51kb78ROqZhA7HoO8RkiuBsn7La1dAPIPDHPb6YUglotdGW
shBGVLlIovtLmVGE65+cHR7jT3Uoswv5Mhbz7eW1u/W5XmFRmqSXXW+i+KoEiec1
SdzQdMQKURiUb2Hpvf9CfOf13Jz+UHy7tC3MVa85Di8r3o4To26se5aDv3h5M5Qq
Nrp5ZFNZEcaCYZvBPPmbJadpqrZUhSaSSzehiimfg0wsuarZndwDixb0FfOy9Qfo
qJf0MH2J/Gqn0prtFRroiofXOh4cwggpb+nJOg9+IEjbC9JJw9x5SyDe8bPPXWTR
tM1Q4xDZ0ABwhz0l+kcM49UCz7okcAfncKWeci+EOMzMbJNVbhvE/+ea54PUe1ZK
cC/O0HTL9zb+Jc3Ivq7D3y6lDxYgIAjENZxflYlBEMlIbJ2ClPGypDK+jbdZJMRN
6SMd3ZHUh0evt6Wqt9n8NWdfFC86yZZIIHG5R9p66yrlXB8PiKC5y9q4AyVWz6XF
HK8bTVeIw3pT7vlO++NnSHWWETrV6GzLC6a8ne53kGXwmRkYoHwgZgtD7uJcZydz
g8F05dpGh/o4jk7S7JkfWOLj7KofUNFOaF0gVn5y2DsfFEvGqKEwtknMKe6IWGI4
iNNklCCE1YsalnAYw4LzBmkWTPX1gfUnHPmAGnZU5wC8SEdfmqUgcVMYrrpBt9L8
2p6CtDDJivX1VNaOWwtnORTe3t+M6lN0BUehc4qqiThbbHfg3pvXL2MuqfvmW4ga
Qfn37WB1UJC6BQ9aiZv42/Temx4xXoqrHnnPpK5CMGsD3v+U8hKkXkA3uXB5YM9J
/cN/1jr951ThvcX3tZHvqJqa8ytUNW7tjhT8N5I0/x08YR/1PxCFn+0OThyfZfYv
jO1PfMZ3TDqxN7PDNOQJFfjQv17r78kn/R38aj4rZrUV3icAwPJ3fXUfYj2j1Y2V
jOZZralkYBtPJoc5OcL1dFDU0ID7aNkjSOcaXEIXaSfBVR7egIGBdsqrKGN5a0a7
lxDRkb8CwDqpUFnJUsQOOnzcEa0L/xWcB8AMYxsjobyTcIW4ID9TId47Jld9wZs9
VLxSPXLcPLqIvwn8KGF1/4C3R8eEtBz5w18syY352fQK4hZ9mHjhiUfozQj1lMq9
NC4riy+ZJoc7M0iUOg6EkGr8dnuo2Fg8dLUadNnaspfHPoKVztIvuMDqpEuKip6w
uKB1hJn/Shosxl3C9PN3mudhDGX3SyhpdoMqjd+xx3ql0hniq1TRQa60DlGmTCKK
yHnZW2gvmeczMxy0VaUsoBDWH9P/M9RhrtrwHV4lhz4NKknvXG7/gu/OXXpswhYT
RsOvq5LGI0RBYmD5Kri6ha4mn2INxWUw7iKu1q5a70CHVoFxluP3QiG7fWIcnbMv
YnsD2QZm1Bkmp7EVENc4N3oAcJ2tbNMd07kX9YAXw2munNDdgYI0ngxII7fMou67
d0G2Au78pC3AYPoW4H/ILCulvbXPw+QFPE6mofALmuaTf5qy+rcRLLA1AND9z7Kv
Nivv+A2trt038b06FHlZJoJJceNmZgg1Ehk/bFalV0BvznjU/tJKyahkWD7dZPF/
WO9M1Kqix5IfprkznsWrnyh0wJe8XN8ql+EfdwOXpNx04Fq8tMo/YRWYqi6uk6zf
2yT0BxsFCF80BTC8M70JGexivnEt41Z9PUrYpN/eOBL1i7AxDjO1RABnWzxRC2Xd
bAKFkQ/qnXLcjuluNAXP0EHKt7OIAMIVEL1bYzGpXsAmzT4aAi0OWsQrXZ7zW2Mh
ntRzo4xGvzQFy2EqMmvqBXqYmspy4jaGmgUKdwtl7lmjoJzHund3XDW0Wr1aDU/H
/iWbGVBdtoVc0m+51sqEFnkPtYzwKfT05Bpn9RX64iAQxWEHYuHGL1VgsKJFOho3
W4Aq5fmCXfTRbqn7kFpAsSCLK8nhpO22NEJFK57YYTwJwD0bjYU+u6+2RGJYn/wm
vStqvBuaM9vpKnfpB4AvzX2RLWemv3vl2umFUVbZ4gFzMWSByvlmVEiK6bD8jBj/
YJZ2cMEF/YvS/niHM4Rnh5DkXdlPmeL5rhJQJU2qgMKkyHI1F4pDOZQ7/1tq4ecY
okty4EWFyERMVQxeaJRgALXjnjhfj8ja5bPoUSu93FmxK57IGsjxXKVn2Qy1Msan
Ub30LAla4ZSDpMD6pwvt6+uEBgZ9Lfnw0eS0eqhTZdQtnm7Fok1BzQ8t4nGeqn4Y
cdA70BBnxVm4miuWKw0C3q6/DeaJtwMnjhU0kBUce7oyc14iSAkSDL+dS/HLKfSl
jiUy5rv4/U5cKQnDn+Iw7w3orjfRWNFtlGnq499/OmeH9vrEXKfETQx0D8O6qsR3
kuQTovt7KUt58JgYtDFmL6fajJ04VD9JuLLMbS7nY628PzW46YRwjdH+UtZvecrZ
Rfcet5k49TDKCJiuSguMJZ+hzQbh6qP19w1b4IS2DYT3P3eNqaOzGGPO9GzOeVU/
1ZiErJ/OLs643akVLbi4zypK2yPrNeime4Ms6qQJIUGaRZ8DTl9hkl4yQibuw4Ny
aOeFpIp0AVsBGySPmNCgIxdFG9ssRw30p81jcasGf+4Fvmab5FlgnEO+cuNk3hCy
dBHbz3j+k859KdlDmqj4ox1lxEyAzzuWMH8PYSJWQL07W8nwu8R26UxDdWmJAbn7
SU6RCDh6GrPUIx+gHk0O9y6H+HrrvDDlfvrA6jVs6SyyReFir6c49byrxn8PvX5J
DgDUmjFoFvIXh2kMWqdfSuYaV9O839mo9gpeLSp1XF61xlwGnFckLjxghN3wtNjJ
LWGjOhE9Pzf0WrQwy9jbSn56vJ9akhWb11LcxQyDEB3fjK9p0htLZ2lu3DR6jPT7
xhOf9pvMm2YDKijC/xyLhKF+4za0aymTyvYtUlt/s0BOFnYuA95OqmDHqD2bDzsN
iAs9v75FX2vSCErgn5egFs5KkeDLdgFMsK9f60ooFTRQKKZeY2X5Fd6cdQPlB4Tz
YdxkHbrplhWtSgjgXefpm8/yACMzDs7m6Hff7ylAAPANGg29uiYhocHibVxL41Qi
618xLekOl9i49hb6X+QR3qHvOEKrwN5I6AZ5vKCkEgR7WJfF+zUdBYwP7EbaAD7+
cJ7V90XDUi+x2CjzCaBYnmf9p3fUxBUsZ/j9UnwbcMhMLTQvSJvizOjVNqPVJoWa
6hb2PjJekn6Ocml+w3T1UjMbWBjSaIptmTiZvrtmlNk+M/+FGZysvquT70gy/mhg
0kIjkTsvt2Tny+j7klfjx1R92ox8XA1VZjPyAKNsycDCy6NEVWBjp5YG9tOtPORk
WOCy4J/gqd+mfFi4EjpolVK7xC+Ih94FQN8HdbT5x00zpEcJyPpsTaJsbkePXegO
P9D4gJH72rdqcMUbzTtoaB8VAuAJgEnH2D7LfGn3IVNAvWaUmhC7EXMY3rw7YreK
klVLiwIGWRnYlfMDsE+wI0WZ8CV+e9CpFHfaIAoPcFFKSkdjGAts5kLxDnY4y1/K
y05SzI3RKUZziMoLL1vR6kLkoUkqUzY+vy2HgOR8xFqHXF46RZTeN9H5TXiGyfuw
jEoeqj373UGJjafgJvWjoHwUg4yB/yMmDuepGFLpRyCwSzlFMgpMk1MP3jquv/2A
QWMrLAGLlgXapb2e+byBBdzrXSJ71a83ynjV56jPGOf+zbZt8yvDRIexE+BntE4t
+xh++MdyLjvRNpRAwHcTvOOD9kNRTJ2ZEGI1SusRS4lPFHfWMXx3qWsnZ0agMW5j
9R/93AhVn0IsYDiIf4YgzSku5EmR/HAriSc8Xh0EgSwwGIcXOVma65MlL6eXPWU3
BXkfZh7rSFOrHl5blj8F2EzCcrNoysXVIsIORbK9MDzUwoZzutlcvD+lM5VGU4RD
3Gu4kBYcTfWdkYLNlUQeIOsF0AXZeUkZ+5VQVXP3N98yOkWNhC8mgZzv+RiUmCcs
nsZ+gUXO9VAbaJGK5K2pAKURftq7Gl1lmVQCdDV1flECGtclhBVjqjR+yzK3XmQv
1D9qBZMPWsVLd3b1NigL2YadsbHEf30v/r4QYcCJTOpCdArwiNzNxou2AkWfge+j
TjFQ8uF/zwjbdvtRNGhAaig8VCxvG7adauyzlXCGrtzW4R2eyA6SuzURh3rKeHwH
YWqU9vwXivbKJRvK2b17XVOcxOrGq70EQMy4FA7CYKj5Dja9lOJ53kchLiSUFV7y
Z061kxhxav0FqjqcDa1Ht+Qa9AfymgJnnAzGZqUTCkMGME5vUvuN02M3izajiuqT
FRdJVBVkd+cU6QGI/b6r44tUT5/3weKWI2FS0+0TSybfmGs6D/pckF65cY4Nwcm9
Xe3CgJ+PHlFAtdolD0NtHeMNMs73SWHsbVkPq8cSHXCt0Sm34eAnJFJcSwQY+RzI
MdIWseUNFxRXvCcuWNLJh0SQyxS405J4Ak0iK6fr9AUqEAqOTSK9jMPihqtpP9SD
yqat+TrBt0zuVwQOFtCzJbN8nnfAEJwK39qxnmuxpY5k6M9zlpmwT9f9Avg3K/A+
WXKDwrB0abLvYXW6X1wSCFdIoEc1PWs7Jzc7z4KbOY+CnsUlXjIINtbziuUoY2pP
FT1/VCh+D8Zhe4BhDxgwzoO7sv+H0MCjMrTM26pb+y+Ij+2qWn6dUqA/TAkiqVJr
mfWpniWpCUeYTQiKWF7iy8sfdZlICEOTpn3hobgHjOtwMPBZNxJ/u7JvedPtWGIC
UbD2mxW0de0yjk9cEo1c+lLkB7ThQy+OcCgAWABnm8/Sdfcu1jQGP5RiuFj0V2aM
YBcEOxS6OdMLJ896WtV8nKYmM1X+GkOxFBftUCPjpS8wIopIYWcuVQhIxUJauP0D
AfCr8kYFsw6HSNhQzWprtfPK5oRRxWQH3kPxW626jVjhE4S6msiZPe6qOV/NqooI
M5jlYI7eM0//i2iKu85UST3HwkwDRT7oTkJxvZUNRbqhHaKxLw4E4jB5z+hGTAbJ
66sDG66Tx0SJbZIClQ0Q1gJRFK5iwGeSRRuLBH5iMu90PydQxXSxz3Dcg765zv+y
TYMwbGzRrgOCMydeP+iwGNGVXk/duggihV3aIZb/P3w3JXn5bJLJDyUnijtICtYv
bfkBX76jTCqA+98Ry8HoTZZ29adxX3XaBUBRZNOMn1TNjfQGxhHiT0B2H3X/+K96
pAJkdGsBPFw32hDz1c0T+gk4PdY+z8IBqbNpWt6Bbyc7aMKr4r3Ct4xgJ8ORxksj
eHrRJ0kKTuOfeWPLVWdc5Tq+Wdm6Sf4blaPEFdAwZ/44WgGotYr/KceVeJpaHHK4
2JyDvzWDO1gbHGcJXzWyAGFAPv5qQYrc1omloqBqnynUsFDYv/eMjopPK/q/W9ZD
BZIeErO0D+yC34dqyOqKOD1ZzCreEJeTYXIc4WxlOEZV1xPxIWJBAgDzwFqYNziu
a/H3OOGG9GR8tUbhdC+FLO2dZJy0UclmgubCkUNvvRvzENiYE7BiJJgWncHb1JGo
c46z4gB4R7oFzdijELcT1INHGYu8l2uw5fi3NM9BDeIvOHwYZTYt1Rqu8S21qr0o
HaDgzGzG9WAzWBr8B+uArSnsFZhhaj8J7SDR9zXJdhJjOlQWo3Q7fhLf/n86rLE5
yEVN1OY/8O5jj8gwtFIf37+iI/Q64FJaoo+KNWfoYUBT/2LTPLfR0MsP0FK8yAFr
Cc/T75Xbs7jrnuq7EivxOF30JT/7bk8hB/DOxSG5BkYSupQPDyHZ8dckR5a3sQhb
yNBfwQHDsLitBHlnbjSBgGTWRoYqaKdMq1GcIyeTVQq66P81G8yVYj9vARZV5GuJ
bBLqUrGwX+HL+Yyb/8YnzRwWFAzPJ3KcnEHBADQ4lcR7GhFkrgkAil1MWr6FnV0u
UX+3qzCwzawwDNogU0ZVMlUTwpjpZWlmzy+v4LILqh9jKCpleEzyrn/IC/wdV/u9
OMJeMLGAq+YXJoGewet81y6nQdM7osc+c1TICLYzrGRf1Ck4Q729K38OiUc3rjK9
48HCAskvCSVjQ5923gFMZn/40t04s5caErSnirVMaost+MQTh9UHpxG4gCcnHzUQ
QxfoCPjvj6MQdDMDcq/GQRpYxR1GEauusj5YS5Rh6l0anApNurjhaiS7Q54cPYsJ
5rjQlRKgrLV2Chucb/QR9ZZ4lUGptZbSZzvONk8mIQ7WYF7Qp8+C+xm/5FoGzb1v
mSuT2e4JH7giBLy/TyBr5L9Vt4St54JDdMueX0EGJ9zZkmcWOt+3/YPQJdCxuoEV
VuIWY3H0/1hjly4dvl3I6iib0nKuSgIwv7N3x1zjNOSdzs1mgu0eLAytCE3QKw56
AzJlTBUvk1CWElqrRBfpC51yXxQ/W+F1PJMYlTLk0bbSvVOoAVJc9hUCmLRq2KNK
ipg3uwN9zDCXH5BfAhIGHUjWQfs5FKiTXYkwQEgeHbyWSUHByp5Dy4Gi1jhIR2XZ
VM7WsN5YuRQ6XwCMKlGB8b9rQ56b3r39yTGl6cfe1QctCPxk7LXluDFFnysEWmOk
LGtxQr6CDpPd6VVHFcCxV4g37cd5Xs86m1ADKzlAUFtUxPMBQqQRBKqihxf/Ojvo
DPxttvHgPIBbwmLAK47/SYuUjl1+T/U29qQdWFrd4C2MgyqE5a6gZ4yvjG+xjSjE
vkmveViQ74zZVY5Nn0K5/U9KOb1a9ncAW61untYyyM/3x5Gmy0tUwexpfQR6Zpk8
gYivAdDD9oWYNXXRbJ3Q1J5J/Jmq2v3bhz0C1xtiHCuzWEExa3+p3ZpwVQ6Aje1J
t1f6gpY5O1Fqin9WW+khXxwm0LgwG6sHpaO2no6h6/t8Jo/z//xQSM29FF6SSgyD
78BsxYhQowR35Ny7Cw4Oo9ksNMHdmR+ts1bwExFe+cu3R2BmXttFfFBg+QBA2HfN
Piamul4r4+JRTm+aEwisYVoUCy46fA4bOP3Kfb0dVRud9ojN/qJTZ+qWS3Kd1sHD
b9iIyZ8pjX2ayLHbTyp1NwNhW/ltZUmzHeUckKd5v3eP0wSttA24DDEkRUswYrox
wDj9k+7LTVb3vpKMrC2YJTHfZUaf6ZlsdW0VvmU8InNj9I4aCX6IZqyWWvlIlBPu
2FiqvPbUeRbTtsBiy/GL6dC0EIQ1IJrH1RAFvXFKKSzTAxrtNKnJkcju6iw3sxi5
rx9YvGyvZhumEEdDtx0+5SZe5hYpUFdLVgrJTAw68BneCL7JvcpFnGgPIj7oCxav
nQxjDmzLQy+N97wO7l8ESpbv6jzHyUMCRvdvjdFhZyppkFTLkuWvst5mGEp/Dh+8
jkPNNTNR7OvxsIk/SYDrqwhbUzr4MclSHN9ugs3XfvKjlMn0p8HEFRwaXcbHE+6A
dgZSasjULL/1BA/vwUwcnxNSTzgUm3h1Lj//3MKT/K6nLkf2jcjWYAApzJSaoWc+
y93vHvG/3isLHQeZjHpAkW8DZhmla/jZgO44AY3e6qBkSrmQ78uVXRMqrO4wId3G
shjaf3EakIolnvcZ83DA7gk7TvltAc6bkS/WHOXUj38LAn8NP6KGgBIfQF/NRwpM
2I/1MDeKF/zdjt+RP4xkOo+xTlrLeYoV5gLrMa7oTPNlp5uDgw9pcEas11r+Cun2
q0hlVesPtc/0n3mWTg9vhOYu4W1mGdX7J5Q1F0H3TFe91OGnkdwoQGyO9QAcss+Y
SzRuqsiYj5CcydVVOt+VyIDiahJRzotmdCIffagOrTI7FEHi0Ls3zOlf6KNKVn5E
LQzlI5YlLRoj78TNqKEyOC6B6jEz+3utaZw/v5Slfdn92PDFKrwuLdhYua7BgQmI
y9h+ayd7coOfpg14pD9XRSFbhr3VmdUl8drFvVSWRedyyy6D/zDATeMI4Ixn4mna
bxw+C24vWDQEOd4UyZWT24JkbNDl1emfdKMxt289lBtoTVeKXmBnMLZCfB8vq68N
rvVDgPgpxi5Z9aLqco7aZ4tzDLBpT6ge0L5j0EPPZ/GynoDLb2sE6eT36Cgr9Dmx
kgrO18XklxQ9D2p/FkgHGp7ERl78meW7SqRd4LszMJI2UYgtwnyLmuJaGyocQnHP
MdZuza406nJgCRfhqbZx+XgoNnwgidqK/rMhd5lzihrD9kQUxBJyj/BitCXI5Utx
Jx07fFTtWihL43wrdtwoctRWnNyoBmvbzWieritWUbbjDu1gK70IN3go46VqHxCB
fvAoSRpLIzkbCaZzyXl91BsduPQtEEvLCS7VYaHUBk3rx+y19sl42OiC2Bo4+0MR
iRWY8KnHpUWb+iaWf1y1K/2grySZcZPXWATD2A7RyFBUJakaPGL3OxM5gbs4kVqd
csmswTLPL5Ba3cm/PaTEebzVid4E3I/XUp6BotPfn0DuZA+IVA7rH+Ht3EwfAjBL
DFy2uNoRgZ8Pter90TXHxOSezyCg7pjZBfFyLVrp92s3sR4O1oVPSJH3QT8ciuQR
adcd/vnwzNM/SkCEfMRub2ELPwW0fR/3Su7zJD6AGmVY2SYnN6IejFRXTU/MlGHn
D4yzMEDU6vmyE0cgae/Z65rXTsORcPPWxfC3ncFijbS320sdVDdXSjhiHvzQLV2x
RZn5gv9I+u9jDUjLR7I/8g0JKNyWgtNT8Zn+oiooFUn6CkXYNJ6rTEFEjVSf3N6E
L7wPNBABcoLViUglu9214wJmM5wRzIPymFR6Iro8yWQ2eWFjrlIiRxZUzinv9r6u
4tbYAogSdZNU21HJMxGVNwy9N1+qsBZqt07b6CkB4hYXFC/6Wa0cgyAC4lkWebcx
T3u/6gqDFq8yqk/5y4DXioMd2tdtZ2IrJjpww4jrmSUTe3E1+HyhXW1qS0IOlcay
zmHhXtp0218qaUU8D7nSjK77b4gx12eC8rE3asK5Dv+zZszAPKVE/A7j/ppnet8S
+/F03PhDT1GsoM1POOtWaMXfJ/L604GBykLPJjkv4dH7pcqmRBMcWH2iNhxIJg83
2qFpntYIjTBDGXSPFnffN6et71R876cTzpM4VJ4um0gmtSZYBona60K6QksEC07L
uD7PXP7Q75aA7J+tT+Ero1mfjP1rM4qw133xASV+X6s8LCntdM4hKvds4+GDJ6Ni
Gu1ZKbrxwKqqvwL4oXYQXAcK1v6VhpRsl2i7qoc6bsMhG1BT5NHaNlbYJpNwn4Cj
AU0D+DtIUzP1DJTwKgPN8j9i914cmUJgHDR8AYj6NVbLzDdEhgBXTX7rsWmKhcFA
L9ula+WYH2bpoHXIAKKOnQaN4OUrBrMxWkEkTuuEThEkh/cmpNOKLBVEyCljtsac
NteSZY4fA1A4c0VR5BzmITcSDci1DXZLYfLoZmhVIuOgu0SMqZRuAxjrGiKQyPOl
YAJWOYqrfYA9PzDzo/sb7KXAb53UhHj6JTav3d3xHY5hDTRpS2X6US2BymPwrnx0
iTK64bUXZcQewXkQ2qNWO9itoUPrq5LW3SWcPp7CneRYPoXwPPlO6WV350WfhX1Y
CDV1GEm3AL+S00tPZQ+KVJrhRt966Zoa0DV2VWuuR+4PiuH2AXyDSKQ2y1WCwP3/
u6nCe6pU0HhcJ2uKFwVyV80pWZ1I6tMUTU3HY7mhLyzpRZDno00vKCe3hshyn7VV
XSv6js6WZJVSUgDvbGL0GXydy5Vi+KcyKc8XqLTwjK7AiFEoA2dO7Z4+y1r2C9Z/
giVg6IdNdHGeUWkYM9COew5vAkpGogsSMPe2kBvAGWZteXhg/XPoZh0laoeC94rY
r2q2V1h2hoyPCQVEuLlqH+q9FVCc60T/9nw47eLTy4zF7+MtZEGfAFUpHrla+47W
0t3ESQYTyrt38wLzXKxCLSjM1btStFkCafqx14c7A5qSUJAZURyEjEF+w/ttIlnj
a0zhuwAxIMx+IP3OxJh4d/yaTqHQjVua7pDjYbmd98BfntT9hJZkE6qlSPb4562r
QHaSMBOFB/SGk80YHTpRlSCsa9rJrrzZ8K/496SJh8Jjavqn0zvC+LdJPuO24y1b
YU4oA3veowRJIiIgnq5CWg4vbFkEtiAx3HaglLaHLGAgVnCrnDDV6SLiJp7i4GwF
S1Kn0rmNJTarHdaLBmQxlBV924dZdWUoSzN9QmqloTMGwbse2ojKbzHR4QK2x473
K51mkOMRaWXGSsDcBuBasVlJ1nt5UhQhbZLKMX6MI0x6Y/OyQJWenyrKu8n21XJb
UrXoYmwW1KdXT+dKAWLP6DUHX3w5wTj9JkbS7hxurhKRdoqRjbKSlSvp2FEBdN6I
51A2zMhW4VvKK+bM2bK1eBGjCAlKVrVaTcv4lBhpE21MSoymuShHbNq9UXuHJjAz
54Q5vu5rPcnoFxkhye4xuWeU0GeI3rxULGHdwCPnprUq63mA5Cmy+SiZMdu7i7Ru
MhzW5gI/K+1LOajTwNrPeeUEGZ73jQMvR2Cb0NjtTWWPIdoZASWISDNSktVADm9S
XdbxeWFpkqptwqauNVDWmE8dSroIR3f2+srseOW1gYaQCteCU30NLjLhYoB6VALc
G/9l+dErMsYBV6NU5kq67TL1hnP6/aqso/FqH2LJrvsL4d3+PVzvOC1oCMPsRMNn
EXiNS37Fv1SNB07xX24Esj7C2hBTNRYope/w+ax+CR/NZ+JjbKnA6+qYSVMLGK8P
eUQlbxHXdAY+GZelxe9m9sEnRr+VfY5Zt5HGwYzNsv6sJ5WhNDnIgZz8nNLKA9YY
hl9uQzRSLqr9U8yPBzSwsgdumbrXXbOeKhRRGIZwpJ3FacbxrUi4cUXeWEbuqb6T
tNAjgU+yHbEZWqeZB/hSBp1mduwbukKbOqFUW2gZUm2mIquLaq5BD6vFmAyvMKUM
Ycudw1KaTWSQtIuf1fHN/TlZCTpsHmWZcpgxkebc8AOBcI3YrnhL9dPNt3c2xjMz
FyquRBfET+KCc4UWIflsv0ZGeBM/7b2xIKvCwImB+J2cjn6FdeL13zm+lZ+RFPbK
y2fekNOJCPvb84aWznbr2BAvuihALDhX/J4LCRCrEdDeUTa4k4HEgaUjokiaK8Ai
34cHHk6ZtQYxk8ez/lqDXVGOIsNjH1yNlU0JDskFyFG/24f2PUUWZIJpLuNX+0Sw
RJUEIhdogZoR71NSlTj+XF5dD9eDGONix39130hBEBouZ/uHJYnSPcm8uv3qxNAH
La7mn+yxWvosC7Cx2bJ0MQuqD08quH5TXq/QEs8C9jgrLv+tbMQ0tJOl1xt71FNM
TpyjGKGqMBBoyDTBtCp5MDT+oDhnMK/Qvr4gTusJCV1pEyH7A+TTeBPVi1fnbxrS
9GgHr58Pr9pYv6THOmrSZcW1y/T7KJLobrXKY9GpcK19ynmlkyFXJt5JzdWkiKHz
fziRuuWjB9BEeGZmnTtSjCCUgF1eloUVmgLHy7vOiA+ej/2gKtG2hxT7PxtRbhQi
M8Vv+Z40/1bsr5A6OxCE7QTpg/3xUDLR4OlegT3ufLNeAEfjurfEymcXtQ73MdlN
qSbv3Xh4v64qHO+ntiL7dg9kO+lKwk0pXV0DWYJx+D+t1+b62BiTnE8+i+GbxyqM
+H6GZmbQlR1DpZ1qcuJ8riTuAH4g8+uWww5svJFJp8eixJBuiPTDBUEe957O9NeF
D7ycOSTZ15W/FWD/8+oNC1mKYj/fbV2RzOWZWLDMlbRy+YBUBaYiXnOlUIShhss0
kkWzKx9rcrPZA32agOCPXVlG7TgmLnJVFqUEX259/v6pAK8ev675gSWnGFdlnZws
/DNDHa6yoaG2fraRvIPgtH3LNIAwJWzBytrTqySUSMT6wtri9gRW6FTvANwfd3hj
Iw75PhqtyuXXJZVmgA8AWHfoWlqBASMEixyn8U0oYkDmZ2CaIVhdUedX1rufUKcI
tsotv0D0N7IshvwYCgc1zkVGZQJkq0I4y5BUL2Z1cUFxU+ce0bBdfkK0lKfb21tS
Pc6GJtwRdoSw2G6kBnc+iUlzeR0UbWHrEieKkLcJXkflvoHbEAf4D3bBePu/GkCM
UisjmM0a/SXRPAiMdlacD9VgWrRUSO0W8Ck4+pkMJJXhlNuU4aEbmXTDyJzPgvqq
0IiSRsS3IfVe6Vx+DdPziTR/HEENmewP+hOT1l6gM749KZeGri8CNH/T9qfZXRUO
fOCVlFgJ80qnvfkrTc4t+R0Nc8Wyur9+EhMzE/GIqQAZWD/4ysWcnlKwaRFY8S+h
JHzrzlQKYzvCGXrH8I75hISSya9/osRKG/yqRgz3huzQw8m0jPktHqGCfw+g7Mk6
SLdOmlqK2JKh2Y//JCUfXXNzhc+11FHmEB19LpGd2YL/Yk96c+wM6D4rOknz/taC
0ny2HsAGPcsjVwVyW41VF2/Qi11/ebH5dredy+TCuptmh9vKM7Tp6IEJ0TdT6cim
xAY5yJY8QvcVXXipHGBiM7pOSpaakLlGPIO+xvgRKU3fdLxgtsNePVxU+ijwKm6L
ozKcGiKivWq6cyybQYiFgOKb70B3XZXXCajueKGY+dfWvyFqeapo7+/ktj3sA0lE
Dn0ggDqVOALUyIP5Eg3XZwuDPNxSD37rFqRZQ6KSimaX3pdToHwLURIfy1eAMYQd
aCdhOogKAbrnTXiIALrOf212YboEIHO8HYe8sGjyRC+PaBa96hdWOL7/qtldFbRh
eMJafFzWYuXYARmnrA62jZ2Q79JO6DmwhsOhrvbAdCmcNqZq8aAXKdNxeLRA15Yw
p8sXSWKTlYw1SjD47Ffj4BwVyFoU/6Fn28kU2SA74+SKnSJXArFtpwatsqvpvI2Q
39ZSGJ7wKGwppKxAt+O+0ULps+o9BrEdQ+Agtu17zCxbVDr1e8DjW+AD3UJ2IgQU
FZMnvc7HOhXSbt2DrnIy0Co1ln+wCLae5Ijf/OhbL2AxrekipytzPH5LAX3CTKJA
qiGHAPt2p7tsbgTJP63XwQCuRgZ0JnEma6skNFE2qug80bC81tv3Pfaa7w+abIst
X9Ay0HxAwuwXcL/RBcR61roDIW9RTfPyQd4J3XeJijUpC37nC/GecchmO346WXWz
rKETEf+Tki9lCpxEdYY3i69+l69cYjJKCx0cFySnSSNHFnNindLwJq8YE1jxLA1V
x3YpJjgmAoJfLx3g0IHtFdSlszdhDHMDO8/n1MgsEvbPxZfq0itUSNb+eCiLLGX+
VLICvNWktUAQv9Blovn6ypi+q5qW9LcyIOr5cA/KZPL4liW2CPgZBYw3lG+uAcMc
jqNkJ1A2GOcQuzTXLqF+G6EoqoHgvoWrK3FuvjNSOOOs263WdyTeQhnp87aoTBNv
+8vBS+Hs6Z2abvku9RHGm3EsrxIFH+tugeegzywzxBwa5afICzXF6ZPTLTJy/N4P
3znVJqmh3Njzel8AzJUw4AzIj0gWvP73LWiceKg8/zsrxXg7ZoEDJQZ7GhBRDuC6
OfvQjbpqj6+r1fi2+c4CFs/BZZTHLg45vePSa4pdTylXrV6o/uryG1+GErNWZ0mC
997ZgtteL47FZ+fvvXOYrc4tk7LUVf0SJUfn9xno4d7RU09gqPiuCx+/JSGOWPbe
u2WWacF6fbqBCWM+t8NXWjOwVbUYilBmLA3ahlMxBawogJO6VD3W9mWHGE183xGs
yCKLpo9qfZpvdxIdTG0uyHcQzVMu4ALgaiZziVKpm6ZaQgqiTUn0uzwbnthEBAer
ynDV6KnIrjNcEOj8NZJt6IShufjKLdStVWRTcGVXW/nrMN96ExU+U46C5hjEvhzV
/wkzYYtDh3PlWKTmpYnSLnEbpKGobA9WHZAfmQ+0ed/ImHdv0MuOu0/pfGSXQAUP
NU9IaRbOi2usQ1rCibYjLP/teXVUeOYsAYYPOeMMHPGx2CVHFspMAKnQMavlqsC4
CQrjM1MSnvnlstr2AauyVsrtXvBJ+P5xhD+V88hl0gNj6tsGEo33SEDsWpSAwVRP
WDqJHVAtg3qev8dseOejCh21Fk+hcCpBOTN6QIJbhk3RkCNOv05efS4jWcwDr1rk
Jh/eFi967rlrAnsb/OGxL0q7ocatAujNmNprHd4DbAeqvlIZFglA08a9T5bPyptt
brdfOh9/B0zigDWCQfj3ROADQ/Pdo6xOGmF9vDKnK7sQt9ipN9qg2NeLfnYTXMvE
GAy9/qcNKrYo0KYTVmoOv90XXBIOQK7EuJdt0y/vH+rHz5P5NcUGhLMUdgnyaYNV
jn5iQ/CT9ZVNBuH5Qs770GD/rpUyqWM8XATZ2WgzTWwsfK1j+J8zjyeD6VPdfY/D
5v4mQF6d/wACZC+SFqwQ4MuboZnXNLxYhq5ayOPFeqExgR0VUAC3LU2zllY7Zawl
hHxkZdq94mB7a/NkC+fhyPw1fRsLiF9pJMZobaqXhhILAEnJoqvpAWIwNahnocVA
LVEM/PG6HEDVK9xzY0knrexjwE3NG6Bk8WPMIkTELb7BzUhWoiAOuBTfvkvispLK
sj4af7gUApj/ulm9rTrZL0g+9DswDyta7vg3maQg25c6PLA8ONs0LiwOyL8IMpL1
I3RVxgl0LkaZ4TP/Y1yB1OGGSKoDz7EC2ogJQP+6P5Xj+HNw8tGQDPPZ1TZeOTzo
y9ZwmTLIrkZHedzpwWkVSSBfCsU9f5j2KzsgQv6IetpsttCpZdfU7oRIdRigy+ZO
kadAzEb/F6QhbQJ474lTOzRL6tnREQQzq901Spo/R6RRDjXVK5aLokqsgMoKm8qS
XGi8jjWY21upWOvnLIOpVqndkRo0DKkLATgkVxZxNDDk/v8cFUxRgzvXgdb2ZmkG
+MZbtaKQCDOjaiiTLj0M6v5X06jJlTCbBj/Q0n3FmPeYtNfSEUaEavxcQT5l0fuJ
QqlBvFhqRm4MXOdFsJbhIk0jhQUNerTP1+Sp3s0rKuZosWsPCdSHpv18U/eO3iVV
5PDixaBj5O+KOtduWBu0densxy6ta5IezDQweZkBtwgWykOmPelTONxfjo7TGni5
c6cujZpEHRrbQdrJbuR3i7Fli5Omy7bVxeaax3UHscXnBDBCpTUZ2K2CBECgCtv2
NxUCeLqNv8XQNTkvEddaor/NfHK+TMVsqmbLPtcXrh8wrtmJAVYq6ZO+beJAseXK
5qzqjUNY72s5Si8h8p/tsoo0CUa1HUAqQpHLd14VJE1gYNZrhuAeA1HdD+G0aO2/
yPc8q65uX7ffwK+5OyP3x92Yi8uKSJ9TZhCNJdALjsMbnF0FQlL33syaceLNxHGF
Mor6donAEllmgQpmNmJbOR9HBJnCQXlw3ulyI7aNGNeOlh6dRmUmxH7Y8rqUSvxH
LZvtOW1jeKZWNBFJRiWjzEsC4tEurJDPGyHI23dbud3XCvrv9J42CjwcYxW7Yx/Y
/gTKQdE9X8/qwpl36iH/a2UJt0g072zZTnIkS8SXdw7ao9U591HXzz6auXKs37+D
Cn1mr2bvbhum47DU6XOAiYbz2+J7mKxKTMvOBJ3zEy5CGRFBZw4TOJV1iYVoHiNL
9ikWTrGlLh9FTiTY8tbscIumEn93K+KP/TGMWD6fMkHG/gXUusShvy8W586CouA1
suwiSME5kee1Wz0vf9jf6q4iwv5lwRLOpsG6qlpHhPCi78c73k7HLYSb5WQpWrIF
/CzRSsB5Ty/6KdhTZ1nDSqIYDkqcvgDm4ECSeTfvz2UyHCLErryRuBYdTYpY+JT+
Kbubwps1/fvLfHQuRyHTHcmNnydmxa5XtKxnjK6H1hFFH72k59MOtDu1Bdd1L/wt
GvvaqgQBAQB0AL+pc8fORsGQjc/lyvTbcI1FerBfQ4AfXSAlazPI5C5mG6eOdh3V
hB70/n49uUGjZSqO6wDg9Y2u5U2PWNsikenDcdg9Y3ghZq06q2BQTF1tJhp10qAn
BDDhhULW2T3FTspd/IBW/uo22+NgtMGO0tX31B9q6hhjxPZGL/R4vukRPpczV+oY
9U5RILSM+tWSD//iJf7qEoTdgC7+4SwX2z/Lg/IWD3esuNUTjQ8c+FdrQ16iJv2E
JjHydemuaX0WQuzyjaTmV2xfBqE5r7PcQOjHyLic/50k1Sf6VuArwGtOTPxciaCD
2xteELkIQ+a7t5zpJMUbluhT8mqF2Jp5+Vvn3sWDtl4YBYJOxs9YXfHOph3jov9D
yP0uAx2rTXAGesMChtAE0AQdjGcPvroXLEubByKQBXqs9W60At5dDG6P4sPPpqd2
uUfstqQU5YQ2n/DpfOiafLWgXwbv0wGCKv/iJH+GT1V+fCUy6LTFiclD8MPgnNJe
fniAqnMypXTSYevwsHbNWVET94d/XzzJtPMidBDc0MjuKKTsNAqrk0UqSD5Ueia1
SnMEI0XNjCC5keKS026vIt8PLC7jsqKMaQTduFMa6jHuhpwYuobX4rqH5NGigj7h
xxs7fWxaQmTuH1GgRQX9rKTwPmUjlrRcESV6vHtlrW5WLpYRKpt8SkZ2zxqsp2P3
KPBecla1Lun9nHoWir0RJ0F+JXwYul4nr12uM1GtE0BvL5Cdgx2epMs/VOncCm/x
GB2gC/NWuQw9DnIESHcckwotsjaXeDx5H/g6nBaNSsmxaZK+z+H0xh/nKmT8LVwD
ORIr7MYFDoRtKDw9+x1hLJGtkECCkxA1BxbADkkP3T7HrzEQJFaQnXrZEvwKjVw7
3+sTi7S/THC8Rc4PmS9Ks9YcmoPEBsbkWmxGgWrd186LrII8dyVWo+/9G27BhsVW
vzrN/fS1/UPD/4+EmJDbcCADbOVkwGR67YlPY3rI7gAcTNNx2OnKkJjuPERVpv3l
o+zhXVEht15QYoKAVdnUNjDiNQfPrY6ZWL40ZlSzBQPplg/c/SlMwjkeTECCqBAa
rpv1DTDf9qru3Phcm/O2TR+YAnY7JH50rSBO3luXwvWH+SKO2dp3ujbwNjBwZHXy
pert7WFj5gBrxo4CGpFer26+f5WuAl/jL5oGeDoLPl5qNG6hAym6b8zSKVh6l4Z6
vp0vGF950Jx0cwkKj32qXY3yMXjz8gMSfwvyXL2bTmc0Mc+L5woAhb4Pr2SVZ7Yg
8Tz0+KZvXsH7pKUZ0Cda+t8HwyTfnjD785eXw2Zgzb93UNNPk9HvGZvD4Fkr4JbL
z7RE90OQCiXY/zXJp4P74EbT3WRjyFTZXVqP9L0hKQB4a/sZUwWvh7ABzbAee5OZ
0Zcuqz+V8W+hbkTBnxmCR37mPUcMj4ezQ6eCKro6ZdBUTFxMzugHYLGPXQbh1jvX
00o0mXwk3RPgEmk5+rRNA7eedBXYyg3iNJOE/E8XtbLd165CJTBP9m6gRfudNKR6
nWrLPJK/5/TdCorxisVldn856roF2NP2aUI99BOX1GLroFJiramw4ZXyxirO4X/7
VtVQl93WbTNZsYL2ztGtG21E9pkdw2icshFfn+m404KNB6UyVSao/r2SKEnzelU3
KSsXiYx89lhHOGOgAf8CfwdcGvQ0hRTP9wdqyEhbya1x1GtoUWbZmGJKVp7t8Y/P
2HCm4dejvIt6veY3oYxGcwZwRZkRRXp04/i1kq1crRfcBC4mZEShvV1ge9vRG3Xo
M1l959RsXtW6pX618Q+jjh7sLnRfj781ztlWN1csLYr3gpJx6zcIVyujMw727vap
eTz/vCxmkiHlQnfaHvkjtmeO1WICBXPwZ2YXHzJnK08O4AQJwh5lC3TIJVbTAb9H
cg9mBsa8NoEVkVoBfxQiSkp80TvEybZdAczntcBn4ERFB7EPOdkiL5f7mJTCPrzF
nrmclm1GQz60iaXCbtcLt8Wyb2au24N5wKEgnT3zDrY3RxSKba0MTPKHBEoMclgW
PtzvPDMS037oUorS+qN9U5pDyiq/d4LB4JGJbl43yKGeFoadu8Uwsbw3dW3GNdvz
54Zh2TeYQ5oKNaYjuNOCutw25Q0uzjbRQ51ggzBb9zMEQSETnovTs1v6PNUiMMxS
KUKu20jFLNPjpWT36xn6hgqT8AKl5rvfk6ccSZAWSXd7Mp2YqguNLVGEJ6s610ns
5YvctWg0GJCSOOvr9RSxuR24Cm6BMWhVGo64Oqp5Uu6D5O/GLGLbTOwzLkTvizjr
a3gcwUSwl83uGTadXTbEsgC2kjaHmvQztMP1t+Xjg3ZVvvLRza+zhYDhu86e+RZB
sD0yIhTSyKQLSiUq8bo7C6+9JYo1Xn+zFlPAt4c/qVlWv31/FPMp0YVAGgZM9oD/
LLTRRK9VY3B4BgIm1cvDwmEPvtHrWze6AUUWOXMFn87CWyWZmF7Qhsr3D7nAD9HJ
jj6MF1/E7DWjK6/zkYAEyALK6TrVEIivbHoYvNlgao/02Lu6JJMUQ0aDHTiKM4ap
z52lC3+QBrSotl4ao9qmuKMYl3AUGmkdQeqtRwfg1grsufTE9wJxvlC+VpD5ln1Z
DjZ7gWwBLekjX8aNbTFn+9xOlGxMn89gJKF99n9a7kx0/fCOrs4N4/y0vU/jAJTE
8KrZHOJmVo1ETTmZ6rp/RUboscNSxpCSjKz8VAtXRR3hH5r1vfef5t7lHKW5ynHq
zyksQWoF8kDrXjbR04//97WbbG7FboHlGUEJGYuJbLbEd8iY5KBOj/CPIR1DXa8a
dXgKPQkKLWb1hHZRROfvoiT0B3mgom/VBDZzvkVLGMHt+UVGTqZBlumoMtcFXD8g
9nFqk7FeoIi8njQ24PefPn/s6ZLMphb0p1STh7Va49HemGyZ26PLye4pv8BTnjja
oas+GI5UlMMSjypJ8iW+YvQ7RwsXKmbAFgRetS+VIwgrG8kZ11YSGeloT8FP0GN5
n2HbEIYIpSvXGTVpmVPMEGBi+BLKCRgMEq21WMWwhctxVklwA4CBkRc4GI4+AOw3
K04+5RY+drBlqaPnrsV+D8oT5WRsHJwIrWe3pbQRv1VmBfkWOOzC1P7r94y1hqTS
LMhW8M9gcse+OzyNIegSMSDZlMyi+jdb5GhobDFTpwYkRhW6u9gC08DWFkgZMnXr
jP1QzY1qN9kQ9q7HLJS8MF2sA4GabM0okXQL0PxRwiKuh1apomMaFLCuCv6tNLpm
2Vk7cp2L4O3PTAWgE9rXe/SXJp82kTBN4tEoSAs9MbQzrs3yzm3UNhvm9DPrykme
gI7aIbqZ+0NMSE3ohvKtznwewBJy9BtQLBfJ+mePSjfahYq0b4poho1SawBNVtkD
9GdYXmU14Tjyc1Pw5N45qZd8s9S02oVmCRw2Ck71z1+nnq0V1BUVMt9+o5JP57mT
V9sx12rxrsmnXFOizfeWJZ3gUF3mNLaAsjxYHiLtc2s5SpJzavHwbkcOXUd4Tg5Y
1liSLky3Dr51jOQZHNZsMoDNoSIcC7NwmEMiNcZyxRE86IJUz1IYf227LpuJTAQo
hwA1UxnbvY5/8niois/DpBYaTXHWFkKgL6ySFwkoor8th4/S+Lp6976mXKg+9nPv
9fDVm9Ezbi58eBXw3PsMroV/cRm9wvJKRxU3wsld3VSH3uisoig5CAH88pD/MhEw
VORtFeqSD1tC2CkPLtzfTflhaZndLIFH+5xZbe9CfD6G4Ueclw5jZ0JjcmOctHBl
zWRowz9kYxgdnxW6dcxDGXM+7/kDHdD7bZafwsDI4QYnrqu8c0b98LPr0J9Gbvx+
Pc/kZi2BBlC6iTfYfkCi6koCqFK2UhTbsjqvbgpM2e/iVdHjrlX9B1HgmwOHUP9w
nA14cqn7zrK/6IYAtIWCQrA9xB2fJGhj5lU0V1b6n+aj8zjr1N6f4MYZPdk63Uqq
W+I0GVCwT+P3l7NVkx8WS451p+CjYWoIQXrLDvvKi1zUuLmSAO3240cSn9rU7tYR
cChO6eauWlYGBhVlUP+14DUB9T+y/E5lxX0pp1jDumUTyr73vhQdDR1O6WYYJvLu
Tjur5bJB3qZ1JW3kCwwHdAGd1THQX79b3f8SXe/g+JhJUVMCaShn5bNG1d+RVIGK
RmAzDxXHA66dSzX8lTE6PR6+OgSsf5OZAKer6Z5jw+05bA2g3b08tYfGmw6qtbGw
eMRvNIiEdEgbh9GkF3xj7WMAKgky6NHPkD7MdUHtl4DFlk7ZVCOdZ/YcMIzheOp7
UPzMJqDSfK+Zu2MOiLfACDYxUogcWAm+RvNWeOJpSzNvfgvCs57MdkWwtKTUYQPJ
cZDEarN4Xd7p8FHfDBjm+fA0QEp+etSmo6+tawqsXdyz7JjhD41e32sbJzOmt7cQ
NTWa7/OjoSvC138VzFhltQKU2uG15MbSIDa8uv9eYSWaUQB3SLsaZa9jeFhDnvFw
pMELXE6C9W24biflnaIEWm131bkbHpIvgGhTyvm+zM+RlFXY7aNM/DgUsVm8Iph2
sZOtJ5os9VZ46hfm66vmZ0391lvuYU5DV0zEZcZ6KsGYdER8j3NDEGBKDqJDv3Jo
Gi2Z3S4qYFkg3178Sx3u+ax9jjd8XrdftUQQSWFPfs+L4Dgr2AUXevM6jqPeQEiU
E/UiIiFAMRcbG62AHkjHDLK1mjczXHnky4smH+/hVHq5OJMMK+d6DTtZebsPYMLD
tZY/dpxLzEplKJaO2fi8I1xn/pUDrFQ4PBkvkGTM//RCT2OVQAoriP7P2Ncia2GC
I6tn1/RkIT6RH5kQ/TyIQqbw4+BKGD8xpWnFikAYGVF3HvVpNtdr35ioRVEWLq5S
qoIJmFG+PLalKj7CectHlurNRuaEwK+/z2iCKWXpLUOUA3ebsUbBCmV/PlVZMt1j
LgsdszX91lyC8lf57PnNVmyhVtoWKLkDCHud1RnQhQRV3MNvSo88+nTjK8IdiDK7
WQQzLcrp9iYyr+cDk0ORxKeU0WDnfIjoxCs3qS7eo+jK1bU/uSUwYvdGV7F3bbSt
0K5HVK2v0Flfmxq2nJUZa1wZvIsp+cKzCTKao/FObzZXEwHEAESEXVq1797Q2YXf
x93/Nsc13uCc2B8iAJ/2rOSlQXY9ghoWuHhWHbk9AfUxSMq7rRQ/MQwiHm0bSQBv
iDeMlUS4txRrsxq4+i2C4UTTObCUIPvihjfKPMgGXaTK8Jvd5VZBzHiLWxqGIccs
6e4RX8K5jIBd0a3PsvmhgN/uldQKrB7V2OP7lyGsdyZc3YgQfOh1lxuY3QhT7d+C
FyuzDb8mn0sNpVXl1i9nH7ZYLY2t/igttCSJL/jArhfBpKu+jV6YoEiKSnHKoZ8b
9q1wrVV77xh8FP4okXIQWlG3MjaY3vedjxeuIGeNXWeU8cP+FjmVMR4OXXe13nHS
nwuONgXCpVCaN3Em2s9LWzQS/TCS4YydNZAj2G9Yy/+tTW7HUvabvGFNp18BDqLB
TFUet6DPrDo1UZmPDk4vKIUN4DKkPFLV+i8qTVy+dcK17zsuESIwXK6QjZgQX5ZN
SL1y1sOhLgyBFIkEjQ9oQAYXvKSIidtD31LVkuWN8rHQ5MNxht6U9J4b75/Zztpg
mdaKqXv3j/HoRhv3jZbrfH2lIt5RD5f8hM1tl61xBOfZ5qDUDLXNgxhOBnLTOn+J
iV6So2cqd2JoOc1plP9GuDNPvR+0DY+/x1qiCb1sto8oXuSZlXpcuFvkF/r407x7
Ceyfx60mml6m7gXUGgd5nUgWBR1thrzARrJOIVKqBShwPyUtHVUpg+QKZbjscQKp
RCAQLyK+eo+Y9baWQThNER9rHSDzLMLPrQibYgmIoF3CIWimy7zDfaLqrW0X21lg
UxtHwAMGQSHbOfFwiIZ0IgRtOMfXGYH8hxx+VtP8saZjdGR4kdH3AQJ/fp31EWSg
BuDaCStCRg8QehZPUu1RB3PtZcFQRet7kGY+wBWoFGhbSXTbCt9KOvmmIpHqA+KE
FRAtzfwkL6AGuU3AMd4Tw7GO0NM3hqhOUgw6xZOsfYqNVUiKYAsHyg2eA5q0fX5P
Cu3hOWj+yYBRmvr9QH3IXSA4gEFdmtmgHvKFNmHHy7G2A+acgtvJzh13H6ovwCZC
01K9YhDX7C7umLdiZ1Q2so+FkCrAEP249mbwZJKWywROk2mkwe9xra/TKUJg8SSD
zrJKV0KdeyFZhmT3lTPCkk9MIu8h39/qFUOSiXFJBcBRm3/fjIQ/3pocbq52Kyii
kh6OKSY/LpfRIQ2LtRsuMdWnGvbWkIgeAvahvsjyM8d7yPBgAMvgQ5Od33uwjfnf
mkdC0EJGh78DiAHtjUN4Na1ywkBPYUdsro0fIbbNNzN+IE4tqdayJGXUQRAtITUP
ZWUWJc1/oopZjulYowgFJViajZoUQxtxSIZlTdrDAQ76CUYMHWVZwVBIAQdCbuqS
Cy2UCZHpaZyjJqFLGLWnrKj3rq6HJi/1qFBWYeACxdEqpuOlGomeWHfwzbPh93RN
DQWq0dPq6t/lnNMMmcuzSJ866fjYmk7wE5w76VHzKrzrQEuaZWZJihdpjm2UzYlY
rhZzPG1W1UJbxvMXD8+2t6VgH5c9Y1260ynCYehyiJ7oIBhczva2OsQfcWhfOudC
SMDmSjmhbZoBnVMO+eWt8iLRpiq0pvHhWLA05x/SeBw9fgfTiYOIoYyUWtVqV9JO
NuHgZQaQrcYryM0bLfhcqCfQ1Hg/OIVGJB4h9BIVx9rh9Wfcq+vThxmjbm0KNsm8
xKiwNOisSxtEJsjgGhDkDjGXrXAhU/uoaYv/49YB+8wvJmph7AqyT9n5nWt5IRkO
GhdAkSySZVGCz4XGexihw5F9cQ3VPZUYpKj8+K61JVo8Ou8965TvRdfsGNtUskyf
JGEEp/cy3JcXxBlFiTZB0MTyc8vOUHDlaxdXBQqnIndrZS3G6HhUssgT/o3QYVx+
w0aRM8ZyHannrb8d1LRHIxDCU/jWbap5Uv6uiB7R49WKajH6kXvR3XdLHFbm5hFt
dJAX+Up+8HMQJEY75l9Ld/O4uFdQaJMnOu2Fj6dlN2rRSOkgxbcV3tPyoqHIJtct
AjDukf1gvE5KqCVJ/gzaV+qifGzP9keJp0P5UDhuyvOMiOn2M3rJhOFwGEVefxw0
odQGVq5H2hVYhqsajMGABbUi7rxKORAmd5YOnD41u3hD+JWXHCNcvbd6AZun9Iif
+pn79eis+5OjoTzZk4MPSvtxDjbS7vQPjxg7gtvk7/MZ7NXxSw2yRWpm8xfV1/7q
5U5nEd4Ypwzir4rXr/9J4BkmyGz1sRUT8ESscHk/lbZn4ecxFOSG+4HXkHOEtZFn
LSthusuT7wRp193BWHCWW9HXZZKVzF3RQe0QIfzW9uzY8VsMYCqUsJEFy5CrWQyO
t7yyw7CP6wy04YCuiHwJ29kwzPcpNxSJz+aTFGdnvyzaxVlF1TtEK18eTA/7jDhO
hmlCEpovV/sARGE5zS0nKU3tNWVkeq48A7kpsr3oD6yM5HVNtoVr99TXFNbZPe5V
EGzlnMQbyE3+LTptCPtv1G8FLJlVmCJsqII4X3H5eelKTFvceEW1lwUeXjWSr/Qv
rLT1Jlo5WTiXCkec6N0OG3bMkVYX4oui4pkGnPLU1J46NBTzwmaUJ+dKOrjmVkYt
NquRYii8DvCxhem8OrUXpKxt4lHACKw6gt0k6PXv9fRuRVhAWEqHKwn77bvUDNWI
8NMwwoZK3hGP1VO1+cPvfCpsupgknVZLQnVN2XJzDkHaDEgpwGLkWT7sl1OuQku2
OhbVO95cn3i8aOUz1baBZTwzQtOy9BNt5T0+rbnpdHVYLM3EfaEDJ8Af+Cr4P2Dd
E17xI+HVz797eaUQEPiZYgEwMpsgupBnQ/3qXbuKskSo+ZwG9r+rFOsF9keyEbkM
0W4IgBrskberP8UzuRmCc9IWe4IBKz6YlWX/zsKWuJ7CriiZRJriR7HGM9QOSUtO
ZJkOV0yHYNosUvLhyy0HDXOAOV17gy31jR650CU2/YKsutuDbREaGRkGA4jlyZGu
VIchDtRebkbaeL9zwXnQ0aeSm/SSFD8xNrb19xHVRL5j0LiqtXQtBs1sxLlYa+bd
YGV616Q8GNkeFG4XRNUTUaW/hw6GOtnzHq3r5xMiamxsWLbIFXUOSTmSk8qMwXN4
fcdnleClRa0YE00HmodlaoezOxbZzxiIETuj3mI4cFRmFvkYLqJe6nc7y9RAE+8l
heLx85FBANuPnq4+LK4zKHzhSKjfDtnkx7UicwEcyvahgwivPFVhdk3A+Q8iPCt0
U1U+cH9XEmkcx/+bXFt250weF37xwIXwFBk42CHL9a7XfZf1jjSIpM/STWg739W6
0ii4w5ZU9/jkCC8++XiorCNHHNBj+tc8ldmtj+tG77f8vOSGmzVbw35yS0WlESmA
hFG7vKWpJtZtqwCKFfnBmuawFuOVr2MwPL9xURCU0r/5XZd6Vf8twwn3SHnRh5IO
unD4rvmJAUN5EdZvU1BOqT7Rkstsyb+DzTH79C8Mh193sehz0doX2YI7oNt1LnjM
XKqiAFEj3X6cr0jnNoCDzDeUlbQ6JsGSdWOVhKJuqFQfVkAssYp6qaP/byrNP0QC
Z6oaD1QtNm5mPQGlesexZ6+Zq+XoMSE6WJZrZ1aFmK/sHCBdw/ZY+EiyDEu8NShO
JdRdpmpquH1O4avxJzehjrbrH7W608ZepnGpxu6VPwFkng9LozbHd/w1anSD8pKT
lsLZSWYLbnyBnXDigEXFSk3Ac0nCueAGhoZFGnhQVIJev8diKFD79buT8MW1rVkl
gVtcm9gVzJTcYIoeirFB7W2ZVtM2ZyQbT6p1ySQK97oOb1HG+JQplcMr8holYfUG
tW8UlfZxGn/ujfqrqr2n/L6diQp3TBHCTA2KVf5/KQcO5g7MdXd5E2qSoBi7/r6N
Y6BeymPXZdKi4CG37cOEOO4dYueHHeC9iOG36KlSXoazI37leeTU/XrCN74CUnrH
jYjFrZFyj/epxr3PLXil4YQf8b8xWeCqfV6KyepoCeLNWD0iNSo/ls8seRq3+kp8
SWQY9stA6/mLFCoGq0FXrLFkhfV4+jd2EbnMsm5MSnG4OYa8i2WFcTE3v6hntLqU
1fXo4ZsYg3TdGf3bb38+OAXUEvDEIUYli8Qin92FvezdExpDl8WmjsgfUxmCJFuE
aqo10sIdjvpHBdDJgoLykPgDp/u9UsCaVKyKNoxPhRmRt+mQTXSM9ZbXOxqHOywX
Sy/CoIrcExWkWnv8Q6Pa3NICJe0iTkuKsbCNQHLIC46HYXsXjKtLoOUEJOGYGt3R
s2uim59b+WgXARFZstw6cBRj3bZv4P2ls0OJebEG3XudLW/MSlXQkJAzc/voBJfJ
7I1XpnDz75dsuQM1fGKUO3cPqJ07yY5+BIfQByCHUQeYTgViRXAfjAxbSBqUNlFg
GBy5irofq9jC9rBoIvFPEaDO52Oun9jVM+8UY/QxgUUXsW8sIDSfQ1cAI26WbP6W
PNrTvZDYjLpe4g8uLpRqMIN9xpJAELlr/p6JzanOWpTILAQAZ+29fQeMiDRjXgP7
WjHe9ZD1XhqTWUtrpphRooS0FViKh/Ta2XXCeCEpDJwLjMeUkriztITrpw5AMFjg
qEoh7yO6Tbgx61Gxv6PEHi4+4q1VYi1pwNS1Hr5l5BBd8jbM2BObf3aTCj0hUf3d
b95UCL3jv6fuhIqB6TZ8q5THQ16nKnvVybW71RMBa1rMxuBsfYrU3b+H7If8Wave
/a9o2FgqwHleEvw57+SCGJEhGJLIOjM1cXq+DPOzmxGuOr+E4OaorEYZnxv4ObSY
4qQhp2LH/NTy/zRmcnK32S9vW8tIjcKcQEQl35OpON8Fkwwe+nh3xzT4OluQpYYh
dM+kZZ7irojSH5Qe1J1VCQPkYkalvhpHLalP/XNZ6UaMshmNcargCrjvG2+UoQns
dDknlnwtYZKaqj6sL+OsIekUmWIr0UT0ULHHRQLkPYDt5QJ3lycbZEyxi+M8+fV9
1HoEk/M5glLi0jBCOpba09tu6By5RPEMTvcaZeY9gcpPEOd0zFzYueicXqw1tyu3
LDU8KeXaD8VW5AHsCouVMov9ueO5Olp7dRjkL8LEKePzYGTlL+3W9sZPX3uJ56UQ
pQz5+EEJJa5NWiOYCIMLJNY+XJ9dsrezv8N2m4kFRQ07lZn8es0Ur0T3P8XGRt2I
WeFNIiE0hUQvQ2WiKSyw5iZHOc4v9vteaOp0X8hefMbeXXUvAjaXKmY/1X5qyaeN
4aKXFCsVoviSMx4FA2B+KTdA+Iqc1tdpZSGXsaDDsbRi7ZtgYkwdc/AzM9eSvecr
aA30RsLiX/KB/m/hA1evKcUUfGVYB3DXDouD/Hm/f0p/T5cLpRh5aD9ELJqNzipC
pl1MV3NfNujiQy5vBnUTtHScu1TJKVc1cufOaTD2/uflJU4Y0Knw0evKFR2Rk/wq
9eVHWSyQFqfkEWbLd0VazuijxO8S/p7q8TCu2mPWJ/wqSoUM777nP4ZS/IECzMBf
MxB7FZtk70SZj/XkjBPh/C9aVJ+h/0ilLehnHD98C+ijaj58HxDW73iFuRd5CApu
+OmOB+nMvbXUNtlvJ4uzYmx71hP/u3tmjOYPzymtgjzxqLjsdPw11dtymP0/damq
XB/ZYILg46CnvJRC54hgCtYSB6t1Eoj0YuT/OgPNRlsPCilC/jsiEVSc4Ec++uL8
slcMHOqeeRrQug1+b5elaBdmYl60yPKyZwSnEwEHzXviLWXzfhOTouLReCQ9uvkc
RhK7GOlhKRyJVfkLW1TTB8x46qNLtGAOdhWNV+YTWCCiwzyfkbahicht48mPKMY1
1V0VnpFH1T7toX7uu/J6nHGijwvh9cirMZWTj6uWu24eju5gM7JDdeIPbUNhgpTu
DeX6Gu5Kw8/khKo8GxFOH6TfD/k7aOU3wbmdRfzASQZubBPtqfjGFe2MzKU1yYyb
BC2+xozIYp2J318BjRnZiUMqbs/4kAE1L4V+tQsxm46NmUHRntZjVJWVtcr55F0N
Zc4YTQQrsLN6HMXN6fZyN8nHRQIpp/zoNkUhXXIdlynG33uk83+XLhEZtM3r2OMn
SKLJRMmF7253BsWk4hYnTkfPxjqX5vcM1wzboa5IWdI2G/qhD1dZjnxh/RTVDDRw
gMufgRqwtoZWw5092HFj18TAZA9kqFaaa6HAlccZfxa6jHP6nNviC2+FZCzB2ZJj
Xq//JqzazENogHE/oHjmiiJd4YX8QU6fCNNFaDZcnwJ+MHq+oPZ8ZJgPwKX4b0jY
JxXqJHO9xTn/xRyJn/K4KhVjaG29NrqTK42r5DnAs7hkwZF95h46ZfuZaSw311wp
fNQooIYtBVjKudvuuTuU3xUQ2RMIVBBpgr3V974OaH6ROe95RGdlCSA247HNJVWn
joW8g1ok7Zqb6nGH+3um0hC0dfEkkNoBPV41XFmFTHY27eM0jKLOdIpCSgg6BYVk
7LRt6lVO0/ZiujsEx9CrLEDR1HX5Wa8nubuOgQyju+gCOGtZNPCKOikS3f3SIokc
emyEy+pZq2ktXngHz+ePDBemQMY5x+8FrS2ZuDW7NbEdyjPRDCokuDF2wT2MQ7tq
J04ZckqYUcwSKC4SKt8XZsKY1etZKLvUx4eBB3YvrBVL5fMzOsoKDYJd89mCQspL
WijPqzw8rWt0CIw/ZqQWmNLVXRt1XJ9U+FO7DWtPYy209NarWRjW+wisw/znleUw
tIoPTr9fJL4B3WGoMAe51vPuxholZjTzQDK/h4AJQzk1Fu8t2BujCBjFv66Rkp9i
2PWi0v/G2UpMFsA/IMhQcZb0FfdL57ot17h6/l15Uu7t0qhFPbZSS4PqICSjTAn8
oUOoFCVQ/SDr0hNRnWY27/fWeFFvEAjmUlj328BkJY1TUPEPnfKYchrhM1ZNt1eG
9pO6Z+xJDmUpUbIs9uNr92tSkuJJNuuhZWmjnYVlbVQXh7ZGW//FtMdGghdVYa8+
o0bqIR/OXqPYyRKGJw2n1FGzBtIvfIB4P4xZ21DM/Q02ajaHRi4tnEwBx8A9AKZA
cnloE9HDnT0lq8Z7C3r+3PRP5HbIGB/fwOiRL6P6lRNxquZtP4uMvEmuFkXvo9o5
6JJkbvKT2r6Ac9RQNynkRguC5Vw4H2Csi7PIhOh1uKPJYuazTe9r72MiFI6/w9xw
mckN2eXkrlmnpdVkYzm2QZSwi6ArAxD6EZWJBT1jDtIIOSo69no8BgLJ+48vRQNK
OHhkULVxlrZvPTbK3PoHKWBeUVqR+BDhIl7MEW9JHQi+cyXV9AsHCy8zg/BU0+IS
18o/p1NxKP4T7gMvF2OP9f2WIN0pq1LEIhzJr3IXjGSijJIzgG6R/waQAb8iGPln
ayG77dX81TGhFTTmklmMearODtqC0StxhSzNnL0f8XxTZeCVmeJ9zfgHmfZmMw23
HCYwKVCg37NFv31ql5gqRmsUWKvwvR07g8lyhqZ/QRAVvGC53jkr0B/pMoROJpKD
WRWTvsd6SJoMf2agJZo+DRDO/c3PQGgf+epKBeCOF83Y9rLH8yQcA/gN0GHhQGYX
Cv/ehaamZR1TUb6uLcaR7wK+eID43rSw8Y/R/kVw7UXS8HeTtPo3Eg0/xz1Irjlu
TETtKkE8M0ykJFN931Kxy1Ue0mKNzZLJTbrhM0BGxIzmIWjRaQQg4hK+M8s2vsDi
hNKv4kLvpCuXbJajKYVWC6diCg70bcKjKADQH8pyFoRrEsYP1Fcle11uGuEpN5oW
ugNpOZYhJ6u3fNF73xHdG8NttEj/LK8iJM4CktGhIT68mMTejZdfi1geCItewpZJ
hIpH+0UFBmlqKi26+Pknnz6vlRvkFxZrfeYUE/Tp5JQQUMd+MkReTisldY6wilbq
gsPnjIJEPkMTeJI3++q3GYUxhJ+T+VRqzBKDM7ziIB3p8en4taMRW6Hx8uX0+zGE
vrESAiJYCkmt8EbkGw20pmYfeSPis0yjeuJBux768I/sGuegnHKNfFEoYUfvdVej
AE4K9DedpeuU+94zWlLYItuacVOgB+UcZSLPz1Rb54Z84G6a/4LzYy4Gn/gPKJPP
gbIHtO/EgnfBRgMj78fK+I1n24FEDzB42orCnWik68ccm7OKy2L2EpLi2m3xDPM9
AOoqleT5B+1rwB0CD1PprM/014WgzL29FjIUNoHwR287dI9+8GLIoSZ/Sgrr0hlW
z9UpW4dNXCDo4Ljh2/ikpbPf7QxA2itpKrB3cJUpfQp8cvzOt3nZtoydb534dmKR
02bn+rcIgbWxLLxjcgB/oCcS1MAWp02T5PKBaFsy5weWTtH6iMLepCmRxq9mxsu+
EnshXl0QKg+YEvr/MKKnEcjRwbHjVYgaBdW9cFYZkG4huaV9GRcto3337662h28I
lw+p1FZm9QoxUR8u++jbwr9nPxWjp20WjQ6Z+7w3z8F2ttazPWCblUGOhQH3KhRE
Kkl/94Sv9oXOBAR48Hk0so3m+kX+4HEfQXSPOZZYOOpqmeprRueQ6An/t0fW61Nz
mArxLl4u129VaP9nbMSHGL0xcHiLabkC/IokdpJ7Ummxt//d4ZxICkhHSJ8lEbIC
uG5cKUMlY346a4w6V/FJkw5hsy7scPlQrt2hFtdD5XHimZJDOPJjOCKNKirmJlXp
BuV8VrdVLiV25J7NMw+JcQvSSkr6cCz90Vw+mTXCO8UBWs0mLTPLmmC4K1Ibxd1s
jZV8gMGMcGqEU7I8lG1XLgriFo9VWVY+aFYumVOYEzZLQ9lW4e4ZxqSTfhg5U80M
PIrBDQV2cW3kNWA4fgsGYBjYakg/ACvFvXkBvxjEIVD+G5Dn+MneHoRIvQiMhhnF
1i6oYtw6LoJsac+7Vu3eOqpL8F66eIR3T8jam5RuD+t7hun+IRyNeHy0c8RGYZ06
eYvDPk70eLoGdsumJcVB9gGCs9jjqI/zRdcuh7aHU1E5ku3HZHNpZy4YGELQ6UV2
Rnh4wr4oE+8KPE7kG5NxwJIANGBtqqI22uI6I5K6wgAqIVvbq4mWMATFNbRlUO7b
bgkde+bpvA76KUqndYL6+aUbbZtjtGo2rOBf5Dp/tMr+004TWvFkebqywpzSTSkT
FjbJ1KTIhvoxb4U82+mSFWg7pmmF2vNZBZbbeq2rgfRWdZUKGMYQOkkKsB/Pynr/
R0kLo7Fq1Q9+08j4sOc5Yvz0MBXHO43Orgwh0KR+DGiEyq0V+1NTPXMpe4Ww3TIj
X5A6tnMHG8Lp3H0J5JmkJNezacFwKILr46xdDEvOcwxdHQTxa6Vr4UlqvN0WFa5p
1/784cXkUrpb5D05luql/E+ISHdT0hpMzQAN0c95gTNSGsrtoLxhrVyG+iqdWNsn
zOdlK1eZfep5AZT5sFJ2lznT2hIEZzv+Hgl0VjmbTmRxXHSuyhQlM4hpGSMRgv31
9FpqwDfwqUojIGt/nsOXsl+H0zH4+uZY4tiprw2PveKjIbUfmt+EKCY7j0XeE2RS
Eu1NBCt3kXGuCNFgYArb4MzdmjD7zHMgardJdNqvj69s07ElP/WjxKFSzq9TXTM2
XvaDS6Tc1q5oUdCovLqu50TZpCT5tgAKdAvaPDESCJYIWhZXmuoHrpZ9xx0PqscL
j0QHYRlsufvgONPyYMSZIveGHZJ74EcXVfCtL5cuMdt7X1kPLD6VBykjbWxjzukC
IZx4skDZUloa6lvpmZqHp2cQPb1Ki7Njv0F+uB+SFdtBgNuHA01+LzZgmxeRpFxL
BDEfR2s7o5k7z5ngMQP2LrIf94Vzhu577Fl85pZRIOUD5v4y6xDR+1CdPKXnb0Zs
REF84eQOzA8Ht7jn0H38itmKE62Aj7RoNRCnA2/YvtZffe/9dToGH+bR166K/Y9M
wwE3k778KRvhKQcNhareOrC/5tR5RdTE3b05OVzhb62rCjk9qxulckESS8ns5BIv
UZbfJLscoZSiRZGxNFX/HVrkhBvYX2tLDiJp7hfB0ZjwO/bwcubS0CycTh0NMmLC
J/VI+1WqFiAv+St81eZos986L/9D7mB30TShyPchcYaA3cB6+yVHKrccsA1l2+2u
6STSsreXZzC+z70+5cxyhPsAiS7M7iAYobuB7EB9PedolRicPloUnhRzjkG5Wb3I
UXFa0zDOeu9XgFc4dHv9On6SikANm28HiSE9EduvUI5ETMO0O0PdHThrhe7kGqSo
12C8Fb9ZwWPMB2IIZ2lcqGUcfo6WZJEUyJvcxtWyemm7S4jiWo/q+Q66PPXq9VfX
V3bxc1Osz5l2rI8H4YvQY3MZCi0gqj934axw1vjpaLrbXXJWaGwOJWCmEXA+dnVK
RYnO9Im3M7oUa7n9b/3lbvgb440qrVpcJsaFrabRS5ve3xNH8fOvKGh7uQpRVDvr
Kp8DvjENyIHG9jHuRgjqD0sXZ8KhN1jIdsPoc8x9Ku8aDAyeWiimHyAS9UKrU0vl
TyD72I3XM2cWKIsoXIHd2ycL4+zWlIzkU5ZjltbroFULD86dbm3Rm201IXtySPR8
RVgDPgYLsLcLrGlVun1KOM09y95rHyrDVwyJDjtH/hd6SZ5OsKoedC4eZdQEnrRx
FcCUjCJjiyGaV6Tr0wPpUUlqha4PGWWjP8+R4aZ+0kekm0Lq8L/xn7CoTlqhPz8C
zcFhhphdwRjxKlVyOO7KIpb5cH1HDdykz7ogCgXO3lGDGO8zjZhbo5bjgxi7Zl45
jufK9wwzPEhjtMETuU1feewg222zIO0u9JVMpmrqHNxjF1QEqzV7PSHbKOAoyjJu
AfHCZWJAEPaHGwf9mJPKkmhvIV4zeJMXO3Y4w2z5bN/wqth+uJc4Q+fy1Y4jZO2I
8f5MNOP91iep+BnYOHj6wDOeC5rqd80ycgZSO/EMJrUKTPfbcHFWGlVpcDwZ0ZHt
lar3WKZ1/9aOA01/j74dMXwoC0KnUtADhgPP9L/G14fRPIaxGiRmhe9qqzXUzHZs
H6GOAIo4e+/qHdQ+LyEKtGC9l+ljePFfhrAtAHMdOK85MCpUq8RF1AhZopPyvVU+
2qhac4BwVmINu2wZlU9ceskJBdIHvRqJ5BXOwu2di3RgMEoWnziJmLpHqnksLcAb
ecdcDTijJBakZ/fKG5TKCxFDbQEnQsTIFEg5m5cmEenDidyfWOwa0JVVqFKJhXra
u+AwsVTGQpdFv/ChGJKRzHkEdyKla9yi1USTM2Cn+WEGGAh+lxokuydgzTKaRnyG
20wLSriiM62H8/3yhuMLsboLVaJQqCSPWf4o6zEZVo/w8L+wQuOPscdZRq96s0+n
vgKQWC5fhqY9rNhlbAGqFyn4vlfc0NpM/0HwCVklV86sr/W8xfV4JEAAOGRc4g5H
b/VUY3Atf4f5ehnMMLGohL1fEkoLk4v+TW1PhtTZQqpV4O2CIavIGnKvwf8LWagw
GERGk3un3EATs+USqRNaBiMOkYMB0TR85BAqtqO1BN/TNMg3QwYDQnsQUFxWqysT
Lq+dcFp/KGVsY5DtzM/DfRcVbeW24MYCDU3jmCCYQ49hqpeDvMB9LY26t0jtinrb
sqJns9uPXTcd4lX0j2Gx1qTHAQ88lXi6SwpPjZD/mIj2yP78lQ2o/IAyo/MPwOVQ
o+VNyl1moFwJbdz+51UjhFheWgonhVFp9NPRTcuzC0ieVknJXGe9KiEM0BAj2UhP
0W/ZCTPgaDJBT0MWF50UBBCMUj4DnT92uv/6eER6WQYziyGnxro8wwlr/mtpaY18
xMShzYQ1zE1AMO9KlFf8nekr1wPsawbZrRWHZgo1pII+63MMTOcbw/dKCdAz5SNO
tiaqllqzvA+gY4uQs0xsT9HYxVQ2SE7obsMNdfa0aHUYMr4S4HKH6kW9+HxLqOJ5
Vny+cLJQK7RzUITPAyU2mGxRbG98fwIFQm7ojFjgRJt+r91xXJz88hBLwBsUuBF6
YxUdD9xXPw/klkbyhrsD7k4v6kRR7i/K6q4BCX/JggRQIKPJn+l6cRc7IRadnvRT
+g/X+bCtiLgwy0i1XoFah7ybmUxdfyuyQbYhutoI9gkn+r5iE9KEQsehvVqEDfXv
pFiNizY6Qo51OpqnekjEBKYTQPkhxAEl3eHaCKZwb6AFbyWp8H1WEA1PZTlVHoQX
hvzQOZx4GzfJqiDF5uEk/3VxKTLjguunrnW8HmKn6+Ltr5rwGQRfh0asAkJrZoF2
piw+x+9WtwNUu9616O7DnAo8BrmY0WixjZRigYXB/gocMWZPp8RW1AvKhX1pBuUE
+wN65VcrVvrKWri5X2TLQxXK3Oi8yIRt8dczC7gBGTK8+LRF+Sxzjfrckhr75ejG
axwy9PXhwT1USYmgWRvJPT0H/p29VnCEXLzSg5rSF71yBdSnp7rGuUmBfFyM7KCK
uMEKSZ7IvOJoigBFlfVuWQQ2Zkuz19w1J5p7qhn8+79ztnfDcx2UicRzRRXUlqLb
/rU4iov9QNrwknu0IEaB3gyMUgPBdx8T0Fwls+/hrq2APywc9RzOOQ3+LTByLXnH
vd1R+kGFwwsM72ly/VNOmyI1xQstdsEqpF7fUHcCvGsQMs043+t2cKhAtyySx/md
fBDFl76u08bMinvynq4mU15kIeZfRpnGmC+gLY4GLZh7lSLbOu6xUQRlS3qd8AZy
9BSw9g/TTlRq+mNQrprDn2lrDcZcqLZ3ZMCYBhHEI1anin85C6G3s7atjY33sRv0
JKJKVNNiSPOVMoT5URRh/vFPsMIM4bofGhwK/qJUvQew2OCEffXYUf6IQB0BrGlN
4F6uW3MMj+Q3ctxcVrJnwo3V86Z4+p4Enfox58ffGwVdfjD1YNa6ibvhk7fZJ5iU
ZC4x+HzwBSYuFg0h4mAbmBdAan5JAv8DH7Ys+PqbpfKnIs/uCISBDezfTeXFoKjj
l5bnOPO1ErTjeJtRSMnROQBlKMzV5WRWvbTvk707t7pMfl1/1P99OSSN44n6M2j+
AZByvcbsarzug5bYYTJDnCRA15eDpp6B2Di0Pn3AL+Gn7eB6OA3tVm2arUgqrXgQ
nSoHfWus/ZaiFjEZVz+ai6hb6EMvF8iSAZDQGuAO/FfPuxCpOi3pV+S0k89TKn6t
1sVemXb7DAwE6AkHy3IeHjGqExGbG1xivpAjfMKTlaZnP3XZAW3weS2nH8ZKXfHP
S52KinYp8hQPK/z9/i2lwh6uGDm/xlFNgdTwSl4/mb0CCyi+lKRq790RscA/e23e
U4NaaD/E3M7XSzfz63ZuvP1WecuMSAyp587sy8ZoVQw74Z75R5YJqdFwN+XeiNjp
MWgfi884qo5EMwaP+fzGQLS01zig1jNjyGID432PV1nHNvL+2zG+oD7N2bOBQcu9
U62c9FI5+LDR7c2weLgkNnNxgkUHEvHV7/9nLy5/jvf/FjVJGoLFosRZ/tjOTPmP
B9MJB5z3+BjGxfHmCnKpdAcCFBDXXZSwAdItIfli/uIgoZep1fY1Ui2c/3B95VTW
bt1Qsch5tj8Et7vhLcQUnea1uX40fvmFSVnIcZHj9bsdUQMVXQpTbojfDSEBTMt3
OD6FzHDHzbiIuXO6PUiq6f3vIp+x+j1o4/hskzRwZZ1I4xDj12V+/eokPEvbsbhY
3hOPo3ps/tFYQkBNWjCyAlWv4r3uCdX6l+gDuNIdO7J8XpVMcw/MsrfNWVQTKEH7
jLoZB4DKnQemFzyKe1RXqRzvrwf8jZfiucpARyOL62HYO5ORCmyrYPma9TbueGpH
JGcf9K7jeZHio2yHSFPxPSL472qLoz7hXYbxk7ME5/o6vYeR3d0xK8ojRvSqvSD4
OlhaEpdLlbGi3rVv9MxYLy4N7UF0GS62s2+4ylskgfdKGfo6kBhN2ZzTmLTq5sU8
T0Le4wG1v9F13cJrKg12dI19/itewoXW//Uresg4p8MWyPHv1Q9JPRROB1oAAski
8hG4gJgdhqxw/fQkwGAcF5Ld0bCCjhr8MsZa4RTPVIFbvh4Qz93WgWfHS4Tofy2q
hYU2h4ygvYt9T4KjKka3GRNf6hDgTGOtE8Eb2Xma7i4ETlaDiCr+bkxVvASnGXpm
AIZDfyBMlfHpARtSf+pw1LT3JYpi9RJWhaKaAWzJUCprGo50bTAq7+ScIdNZY7Tj
x+wpU2UzY9e2uNywxQ2jmlHvsKx93cDf75xSrPm0z1vzSy0eyzvsAFp0+Ye/N6EC
azAr19xPX8YPQL+fmDD2RnAxOjQcZE2KZos9u6fI5tevvscaTSF4CqDrFt0Po17K
ZdRnoBmKLXI1f9KiqqFWqJVYl66CyzyK/X93KG2yHdV6GV9vbNAhwveGC1X1t+Xd
fyC7NM75w53FlUClqnNgUdAU2k/mTV1++eeo2AriFN5QFeXgLk+49GUU1xhYtkmq
i2smh7NXcd2a5m8n+VmIH2oFLlYCwWhIyYT7H7EWc2kTQ5sPm4Bu0TNcmCYGzzod
x2FI/CI9VuMiWMgzVZCwqKgBv+Bgg0q57Wx3ufcnY5vmZ5yW3FvYSKSzHo8CqHa2
irqR4/7NXHdf98nef95g+diBDZaaEoLn+M/6kQteiArgdDbueAxl0FrqkwxbXZco
5/9fWWJhWz0nVMC4ygZ41vZfjRI+Kh1FZhhxTC2Og6sKo4wyzf4ZMyxzr9hU9SHM
ypYpH+GMVU4bCkqjrDlRuthQz7/gwxx/MmG6rc6pKOLV1Hqif9lsjnD5RErd/yiG
F9+4lx0bthQRJxWeEWD0cp1Y6uaa3UlOfQBXi2shuAUoVxKTE0BfvKEHajdPkbWP
rCs8+edowI4V3B7d/7AMCjMiEmLjEi5zGQUJvaLSQCrKJHoowO1sSJL+3dfESNDf
5jfEtK1bS8DzcoiVawc5MQkbFNz25YP2ZDCL63qau6cudmf2yNLUd8f0xlGXbYca
Tmo3m5sCql3gkP+7zo8eaTpcbIdGgFodcjnkfLz9Y16LyC75J9XHTu2ZarBPLypq
dL2Nd11QT83dyz50KHoAVIjESxVmTJ/6NjaSIkVHyNRiJMgP/j1jKg4bW6qNoT/i
HRjQKVhjZqQhI4y4PyuQP1/9Czrvv99z51xLeo40R7+jw826QrqIX41Hy8P5qz1Z
hvUOCxBb6BeHBoEh5ucE8HDbFBZNzHz5OKAV0Ay/7UaAzvcnsOYVci5U6OnN0LQW
0QiC3UPpFtZ3K3avATUTYKvMGgocjvz+glazl7Xe1cmS8SQy+m4CaoaECTm8QVZP
DcZSKu8iE0s89Rew+1oKK9gK1ncNbUW1KlGZZSGBDwAvnXvdT0En9cHzMVX96T2I
muaIgdz6XpcD5TtIBqB3u7bGuyr/dmcYx7pS1Bq9euhZgRq12vYluix4l84s+WDp
RKgvRi3Zr4av54dzsXehszp1oWk+KpJ8l5rLoW4T4ZpiWEJHWQRssJPH3WvySRRX
tU/V7QtpIAbOKifaMzby1MqrGrxO+fhKqeiUtriHCT2e/XvvpZkBL8P/zkUzvee4
QKO5EjTszeBG10u9FIgOZmpxvS23R2UsfXoqB39Ptoy3pRHDlWM5XxuKuMRdeOY9
O0w2Rn+kw6+upLXdBKMTB58y756Zp90/x7XEspJ4rw4H/yrnKC6xDdn+agkZDuRq
kPgUt+i2eBobS+YT9mcVMkxIptaf01VjQ18q8D3rpnBulLB2Q0jAMwd/xqvIxSne
TgGy7fplkZCcBWulivT3Za67gLz3CKfRYRboUDXIeZfD+OD4LLUt2/6QzaUzDXf4
xOhaRm7kOyss10dycAjWxJOOy93nOT54pd8ub58h5RLEtPxb/x6LC94e2SNLab4b
N6bQIwJvlq4P0lqr+fsVNyH39gjP8zhtYEdCKXM4vgQHKtwFHA/oD2wHtWrB/FgF
dsW35xI8dQLAx8Vp1bxJVZdT2NiUC63sgQL3/YwFjfw6pOoDJ8+4pUvtHKUefBrO
yrOHLE799FU1tRL9NaYpeedPRXzdVFgDEMdD2O3nR/N56G/ElkBJ77Y7sM/8F0vs
55HkPF+TGpxFTuQVImh79LPbfXAWL98SpPs9+BVPS2PTKMlewa21YjhFUIu2l7SI
dhQtysUBDuckPsywqaYCvAfsn+GVEcDdPXiKZjEnij6Ss/1OoWZ0X0jdGkLb/V19
zfWZZVyineMzOH1TNligztw/0oKrgA/i/fTjbDNu66PjJw+ResZxhq8wDZB8wFpq
6UP5B8r7F/mH3A7UkxxMVBU3Z5zigdJP3xyZ+caBzdz7HCNtL3mHCYqPt79XM69u
yAXDgI/wxKev41773XxM9Uq3DNi1MXuYUszn7W7kvQEnwBA/2Qa9VqXk4rsggMwu
9hmxxz9ikYYAdoO7fHAoRh7YL9yAHd/WqXjsxbKdvTBj8Ct9yfnxKtuQP1WbQ7wV
NUOkUgcMJLWlWg1Fw5gRUg13rJl4jNnLgspHy6XnD98X3Zk6vgWeQXbfFrrZbzK+
lKhIyKiyf7tomwaGILz230LgGH5yBIDe/yDPD8L/IQVOC/7RiSgecyvxqAe0oq0e
3UWm4fNR/kNwhgl188e91HQxt6jm17TIaezfzr1dzEUG+hRr28EKhuewk7lSTXvr
eYMsCh7keghsHA4KcBOFMMsppwyH3p/ymH0WGfP1M+wEFtgFq9L3ln6yzlBLhYHH
gFUNnsoPT0NOX8K1WTgOXr4PCHCHzlqyFO5/ROvaTFNFtbwmKZ4NWHHz+ApaBf/b
Fd3WYevCjJQ+VGOLnhVFo/Q0D89DbeB8U5TG6M7eJRDLvxBfD32Ns82WmFpKfY+b
0q/stX6AncchhphrOvrUN5a38ZuujImquNjk3GRoGtVjkMGZGgpdAeqVq0zljz0z
BeluXiSN/7PgixkW7oNtPz7Os/SFLIAjoaqzxibaE3JAsVUkqKh38kFFlQCEB7PB
bjBqVeb8IJuNsTiZmDC9D0udbWrxIGVKToiVXuhHQ+SbOHXNk7LuPpFDwMet3Il4
Zk6FJYCsbHYUeGsiDf6Envxx8wEENjBvjBE1HUVBRE07xtrP8CRuk2Ilhi1ylCP/
fCyZ+6OHGqW0WvXqyDiegWro+JasrTi9Bsm346IG5Qk76JNppOzihaiDQd/0N5vC
IOF86lFS+bKTe0HNgGIj2eF3WBGyHxVcaXjJEMRJHNO8pb3ORq6Tv1RGPBEKDDeX
JG/+oCAOtZls0fEK48cgJoJViJSKk5d1ZDv6CNWc/wOBwhX3DGLJ7IgpQsX4QggO
k6IVBncVjZNG7LYJCqLK9lLoyIi+8SIBrxU5FAIWyvrNbYHwvWSvMA7GdFbAwb5D
in2DEH3VyQPd2YFsNe7QXmGWSWY3Z6ROGELSq9FKux9ZdcsNtPjW6sVkE7DvoRWn
SRqZhnUWtBRnJRxq61dKPBQOtUk5s/XV/xesJnIOitYypKdFBUGnw1mXd2ooftqY
eY3qcphuJ+KH9xFy1FHdhMlhd7P3Ke7P+PI/L3OqXa3VI/rYyf/lvpnWHWt3/cxE
JbnExrV6aH3cSWN5Bij70gl8RZhJclHKnYnzvIHgkqS41el/Q9rbqOM4VVzipz2q
VbLuO83SnsDaOKGmiGef6WzeL85c8xjx/A4ugAQ9xzvNltIBehh49wq66mRcyokP
Y0xl6oTV191/HntdkoBfwaerbEKUkIUS/nGJhoOl/wY3YdxcXv5JvIIpi+FEftUg
mkrJHufxUDvDcuZigAz0AcjWIaxYeT6fvD40Bi6BdaJkjumVcOhrbGXynyDb3Ene
auXOazeOpKyDAwAlEElPcu0GT2YllVHqWmE3BPMPYQioTRjydnGo+rQEtsBoOyWI
wKqwq5JOgTY6jVA9CAD/7EYZUD6fssmAl3mK9WNpIMTCuPhk+COoCVUvw/mwMrua
CZYDSP5Zmhvw5JkPGwFMyeaMfbY4gEUJhH9QiDozj81nTFOSpo/ZsM3p9RR4s2TO
Qh5X9sbrGAyERxH6lIXe82hCjWVgW/N9Ar4i5zZ2a36VqJc0/i3kkM9klYMknJ0N
wj/O2qKRu5pj95dK9xn86qO2822VGzrlr4Pzi2Z7KCGhT3XT7iX3BWyXw5cC6G1b
wbiteyLqtRXjb4rqOhoJjIVOHoYQYNks02gfjT26/Z3ZrPJzbPktaq3HD8n8SiYr
aGe0cTu7Sr0hePzo/kOqkPeur9iHYAXMWN8C5Wf4OhCIpyn+c5ISttw8HqTJS0Cr
DMxJ3ZWu2TquW/9ggQP3QsO/KK02alSToCcvCszj8BPlOOmCMhDoo+GTwRbsF/qB
1qooEXGUfxaW1NikXzbp9l6ife5ghKy0wUiXmGxiEP0lnYCseFiSql+J0TQqsQyp
nH3EgbCCtjP+TUA9u2EckViUOELjGIvlPwPa9AEUhLJ731d+8Z52GILvuKsLYVJT
d1yV5W5VCFfkaD4xgxC+fcLVyYrOo4LtdTDqK8jj0W0tUGINVqDfRPfHy83QUusJ
ODDnxp/3wekF7A+v+x8ff3XkBtFG/W+Cb88WDAYfVQeDELcgvLJ3kjLos7WFihQo
FDOTlcOm7WB63JQPdW70JuogAX4dEOmFIdGMa8H65K5mYuc/tsl/eMCoNBa81Lpm
A+BiScSH3MQlnK0L5/KCeICRc3Nu00QjqEQ3xtfOgqhfNPHoZPzSpMtu6n/1TE+S
7S/ORmoUAfzcKX8z+2gzibeP/8jKBX0ldPBat7172nx6wC97KBZElq1lRuu4m4nC
9UaAZDmFLwH+8IEnzHSVHK2YYSvZ4B+/TUpHZJBbaFxrWKavma1EqYHKIcQEdjks
Pol6kec7GaNyh8VX2wzqnR11BK6TPzUjUgqfI9SrvD72F67mZEnpC1Og1cG8SS7P
KfMic0d7f1FmMFRqz6HjSqZUfIcCJRjC4IxhPFFH454fToKVe7J6IR2IJfAanGco
oyDvRQVCfEC3RJqksMy8JlpStW1+jpxsUb5rcIxNT9VU8qyyLjdIU+WhL3du4wjR
emAKGWWwiqIcXPvi6iXbUa2VlXVn7fkOkeHfPHZBceFk6h86v6Kc3zomiSOb8HbC
e6L/blz6hO0KEIACFnU+mMQh2Q9cIyvoQxad6/3qaA0hwRO7fzIYlyxs6Bw8khNw
b4tq0XxiCgnL65DgsoZlyQUHtOhlbVcItszLTiVvlCej7qz4SAo3zDmY5lEcjxgf
2jh4vPS/1VCYK9YeNELqWbUgVZsb3bZv9Ec0ZE0p1xN26T8YRw26X4IdvIn+RH/H
uPeUypZ1UbkAPI8CTYJa0sHGdIN3/VJNtaWmxkBpG92+qzRMfYJ0HeIUfcjkniBQ
GofsxKIgIRHfzDlpnBTsplTgYxXy/vryCC0SRRFJhlATcJx0PT6HNzD0hKOQAa6k
JhXUw+i+8lNm5AWf2mGzB18p8RJJAfqzMyXzl4QJDSAOhgIqbCpzS1fi5W4n1a7r
dNhpa2Yda0ArGUjYUUXsLBYqqNJEjw71WDPvjqHqlfGvJ+bnCmc/hts8l0BgynD9
C19V87nj+SgfV9v1N9jLh3/8FVrjKTA100V3BE7iEbmQzoF8zrWgDYRLBgWdq9kb
SBdC4a9Kq0UJETrAsTxp7KD/pu6HoM2ZmVapnEuuS9Xes3Pw1n+NQE2hKz2ceN0s
EYhV5HzcRtdljpq3koPGqlmIjPtqeg14HDecdGNFtZBZFHY0WzIhLCEO0Ej52RuZ
lqMSbPh5oheezk+6JAxVMlLsZlArv22UTv2YrWgEEPbDzgcruDBWNSVuufOpzKj2
hh5u83rZQcixYEeTebw//4LDFEIWSIw2WDj4mFzEBoXmx2w9CFB6NCDegDRDTZwk
rquEK2yXmEUF9ncU5l8r6MXMHNdm/nl8ZEPVc0oOKVHZKZfhB/x2PsaHgKSRb2Q1
2tGq0DpLDyGwGTpak4jPm/MoZcbgh7eHUcVtdiBrlGH2lXkjWNQRR6AGhBabnCFP
nlIiH/Nf5Rhc2DAWnPRU3a9sbjbunQ+sjezoBtS/QbnNfRggreZzEBY9vuAsxwqm
eqfkMeSiLjYGouKWe7fWoBa4QhyxSpRhK8Bm3qiUxl/wGc6/Ns/QNrPKzzo/n0RH
5oxmZQwEOefrJzZr6iWepH5BqVuruDQj2eh83UArV7gShFddVICht1Fu9XeShMY+
vPNKcgjg59TqWKIpji1dYpHQYFcnn9ly2Ne1AoFDMm/XWLGwZZ61Q6qUU7DMyY6q
YsQ9smckqWwqC3gUIJr+hbLdsqtHGX71V4JOlmLrC+5dtf8fzO8zwFRODB7IY2lR
pxw2imfJpZS/z57X6KQg1zPyjT5hFoFD5Wd1jjmmWyEKWEdCFxQ1h3DC4Dr/qwaE
QC0PXhQ58D65pP0087IwFPHip34tAnNOrJjxVBDmQJ6JAOHWFSBpvCCazdiA+xC2
/JCl5Rt5GbKv/qVVsfZxWKWI5Pj3I1A6rwo7gKyKUBfHwdtbnaCF55aDk3/Eyox0
IjyZpYOPps/8Hm89yuwjwn/iOkX10vPw9EG2aQnSls61oLjuBg486TWPBomJkLPu
49j3cmy1/PdvdH+gBpMSUdPsdaLNcIIOQV2/lu8Hktg9dkmq41hTP2NdaGj9ufki
CLyDtMZUfJ7H8OKI7JVrgDuu5+JTc53pCtI32YjcAgNR64akC2ZfMO+c+JrTTCIc
xkkVs7OApV22s2ExzFzqr6Yb8TbWSjjWhdq9/LwWuub+FhYxv9+yCO1W5vVfwMKb
JxeHv7zHzjTWKaA8ODlDYMEWMAEIlYJnVLMMlcu8wyZNNakCILDo4ytMEgvdpI5k
pmMXOvayo3g4UrulYwFPf5AgcTAVcowJQcsyjWp2tp437j4k05QrzJEeSR2qCCU3
LjULrAl3/u6M3vSQQ8dVvqYbyuCLxiDRecYcr2sZry90MB14Eec8VD5yj/+Wndtk
i3VRYuPi8zJXhdXk1GqTP+ZBAFxlOCrn9+rJyapxVkAaEuPgteXjKiCRrWG4hJCi
rVZw3aCxR01QNL0Fk2sXT08KDYavQmGCmeJ0U24dm/Of2n+8/EnChtmqlFfa9ZKw
o2gIdWPDZNkSuE4eOvo8uhjGKDU9uMOSPaHJICEKc4+1YM5z5m2rMZkORXLLfBfK
gmxXEnVgiIP578L7bJyD020duzCuPjmLBAhv+S73+1NPK61q+ruW7JkCrkfbTqzs
4f0nFWJ95O+MhIqrek5TKTJ9DSILYLe5B+rfOs+L9fGPi6JAnVSlJHD0jVPtkfam
X8I/SL2DxJDMu7z+ZFjV6/YjhmQU5yq+BMCuVDkkorfKc3EK3FbNQSdVBlksBM3c
CNJjFFXaHRYSjVFsLcn1fXgEYUi0Ir76bl6I4Dmbx7XVnm1i2cwDCAVKQHgGrS7c
3hrazRgMG9C8S6pmLm86Qx1TVVRRKZ8rb5lZjE4hhuOg9q/D0K3fO0QBuyJ9vdjq
TfQk16SevF3xwHFNc56z5d7h+jnBsDIKO87Hb2+1ss9NuS5f9to2LmfmvFjJs4WY
9rqsceF3PDvH99xQgy+jGtLiTWfDm3iP73AmVQe1vU2U3tUBj16FU1niQ3XGQ3Cg
Nq79H//yugotwEBM1u1ue1j9orDAXd0DJIffck4OS5s3pVJrKKPBUiPOHQxXyZZD
11lyM40D9HHzzNr4nz2wCef4f+hb2DxtiOKCKw9VDtboib09TnGXZNDl00fK6lpv
m3b6oWeTD0JKvYZ2mh4gI7oHEe6BJRoXXjm8AaKQf5k/qrhxFMxfz1xry5ZF6PfB
o/XbFOI644oRjvn7DQkthjddYW8EKrcBTC7PT1BNEvVI2yEXK9gkJnGS+2E/MkGM
+eYg8F2KVD8lrrUEjGDMC6jl/NKMqYx0AnNWeWrJyhC4EIm+9q/6BjzLb5Ea3Gbp
2AQgOhZPvgaDk7SizodKQ9FJ5zQrOMbA326T2yBc+nLdrNz/E95rc4LsINvtsgQf
Cdc/8DwymMKRhRqc48pQWQulhgu2V8edTj5ZzKd3z3hBtYBHsJTGZ0MVj0u91+fi
k60OHrzsXNhgoWS2/pE+TZhMasZzza4RPieclWe9mDaovoNWWeqy2t0nuNpoGRwD
hSV/XpDlOkTkgNJtNloFq8r3A1BETfXNbZBCjmzjk0lJS3rm0zf7E5Vr9ZKsRCQg
mabAa2r8gGWZHB0OGBwvmjX5fopLyPcr9KCe3bQxgyFg4wgxEQU16FkH8lkrsrBJ
J9KVx3AuA4T7EXEVEyqTBDN3rTdiHUJjmiEEm1knn9dDhp3+FVAzCJnP0rVcXPWq
hLQ+bDreiEqfCOZiPPPgrnAzDazPuq96dms795RKpDDa3o/EDrjmExmsByoC2MoR
Hb/u53tFf1+cmTg4qYb96j7vDIOjesylgx7yXc3O04MFU2Ypv+DGis3U7AdsDS0H
ASy3SMIxzMqrvLUz03p64o3/F+lcLy6R5UmcXUFKzjiQ99zPQ7i+RN6H0eCow63t
dFn8+9QKQzp2DznsSt1JV4/OO+xZdrXY17gK6e6zVAM/0COeTgX9phOJdiIIh6rP
QZ1AqLJiTMz3+cEOuNmyn+306rsgIkEcVFsu7T6+kMD4xX4W1s6qwu7Isa4ofS7u
GNpQWqQWdqwwz4T/j3UtzONCztsXUFhATrpneZpOyJN3SD8WRpSPoINbHFmDg0KP
BVXWf3cglQ+5FEpZeY84at4jelmAPRoqocsEBXilkyR9jiZZOtb3W0ooYo+uBSPL
nIWr/rMq6AcL09BmxrZBWayll0/lRAjWuLgc/SL25c4ZpD/QhbpIFskyr2VL/9Fa
UzZOAhuKw4DiNr8/Hx5xbKqEkb7JabL8diRB6fGy6YG+e+5WujL0AVDVYsXACN1z
3lqUTZkWwDrvnj9AC9vR+BdkNmDhyBwbrUAuqw+rpr9UnWhtrsDVK426BAJ0r9bH
9ZyHcSujy+qa1FpAIih0T/1HDEtLTnau5JnDQDxlOvkKlfSFtFhh+P0bdiibMYvp
uqTYsWUNrY80s8yBYz9mK6kXpLJYwezQzan6GXLE21v4C32FcfovM5ImCvVB+FMg
G6sdW3s8SEhwVMfiKiOJxXYEKYaJ2npePG9uTu4xRjt9I+DuAN8fF9R8nebQWINp
jYG08kVVJ+0DNeD5hl10cRVHBPuDLKmkHf/UMaO0y5ykKg82rOrdYiNHP9lXAR5q
7IzVefnH2IogyUViAZR46xIyFjKhBxE9TY0sdKak/1fwEcGKy85BmDJdEFlvW89Q
ArloouXB9jTOqUPHuEhHHT0f5P28UmEletcVHa33XykkSZJ0QliGdOKd5zc+hQrb
xnG5VFeEDbaVOw3vmivXrPrl4e3W7khsW91+ERxX7Y8bQUE9P8onvKOOT7W+eOY2
zLYuDNtVQDK7t87lCyp4e/4QYZB04/TPsWg9C0MfKlg6VeBkW5zjBM6GxYVKYpmv
+yUELJNKKEgI+TYB0xhIEr6aRuF9tjFJj2D/knZhMEdZXcFIjw0xo1HT/NVLRKzZ
f7WTq9BjaOwQtCUXd2SJFsCR3n50q65hbSQrkt1pnqjyxv1fD8Nb7cOFXNpurLnp
iP2EE3V0wFTQme4ij6NMg2i0j1uvpuSsKwHevcdp7NCnFhVlScvebLb7yn1qOrg+
fgEDrCl0rHx+0wPV8Z/z72DeDB3qBjlltylmx/OhT703qkyQtU3AcaOOLVQyR+dY
UUiWvjGRDzgaYp2xPLeUuxrwJ0FTym+viRZnW5YOIK507KGIZidkVYuMeg0NZHlv
uw8C1Oz+lX2sFAWhqm9VL57ZvptOrD483BkyHxfpdN7olaXuHforWsKSxlpGu53x
DnIA8uWj4O6ggfMEqLz5ye4qYFDVfNsRU2FZ0fYLD0q1zTNTdQHUxx2DgcETR0G2
5dqV+MnXjuCQZRtu4MLIz/QtjTAqHVkDT5eoK4ERn/PK0FFEtfPjPpEEtR3mANCx
Ut//kQRS7uPMWdPY07mli4m1kVrLxukqD6Nltwx0MrqAGWCYjGDRX8GndooZ0ag4
gJvr1QX33jmt8JSSZjqWqIB4rGQRLvS2Jj7iDbBS9kbCs5J4Cs79Djv9TCj4yCpu
mxFDCV5ieV2mnYVo0n6mewq3V6YLC/Jbh1cN+jI1Ol/1BNIKSth8C/hxTrsoF0wx
H3+YLtDGfUvpxqly2yVKJOUZZkI3WvH3c5D7My2Uv9iTMzukqPPk7duxpI2wqbmq
Ft/rBWag5l7XX7xu0Q18zID86cZLPr+Pd1ib1CNX6HnnWqcx4MijAnrZBKqK3RJO
Q8EIBXuR755bE+6bGIusy8eSgWYu7s7p5Qn5mpeOpWxxPenIR/D9hyZn+oH0akGb
gfXT2kmK8+m/fvc0oAa39sA++1CVvxAwa+cKcV1n7V0WjpFmJlowqeJZWsaezfdx
QJZhoWvWZBRyglP9+A6Yi5O1YdouxEDKurJco5o6b7SPEZ4NmlMeXylBrJhiOJRq
enEw2NzVdF8WDYhdJF4Lx5AxWkR8ecR5SBcSS3ZaZf59RHHzwDol57CuO7mOloo9
cu02g8W8QZUoE10O2mRUk/N3vwW4jUA0fUS4ZcuQSj5Uhix9aYt1QEOV0KcS5bPn
aTCNFU01M424bbztahjVOMTVrQ60sI2GdhSKumjbU2dHSBdYmHfdAuJ47AWB8i+O
Yv0RNRvhsFzYf9yx8lxnBBjJlwCu0N7j2FOFBc3RA0PeNhZqQ+/LKWECUNJzlYtU
Krl2yNVUepw4pUCC7ID/34E6UgOjgpMlZVU0yxDLB1fQUdnDNcgotYp+fYeX37MN
5ODhQkmPnt6LfscZ5A9EJ2YlToTbQkUcnKwBq18FVhKyswlciNiM8O30XHbyU+bP
j0dzpcV39nkzEQI3JaWOoO4O0QqhYoRMDxQrvJanrGrcuSQ31f03G9TK2YDIOR2I
GnBj58p4RSezFcdz+n5ww8q0g36vsCdvd68ImkCOp62xbdWGfEYhQgoEmiIh/ggy
KHJkasdIfLGWE2i3gVKYjJ+uPIxGug4FtMBb4P6Aa8M4gE1vzMVM1IhJ43W/V8dQ
CmBiNfYpwIdNBNApUy25kNIDvilYEiQTwesTUZRZHCd+nX1gs+wVEc/n2j0+TNZq
5q/9doRX5UrrTUX1YjD5gfX5ipK6X6ZrzucMqAL9IMEBW4pFqqKiHJd8emCdA8Uw
KxWIoWCjmn0ARlY0dcxKBPmMJJxuxGE72awuOzaFlj/JBqNg15r2hqyCrPGm4aJW
F3OYxT54vKR1AIzhO27ozyf9ny/mxzVccSnfKW8Lk+MSdh05J9u+GF4a+nKsNb28
A/xdzXYpfbyVn4Z62AAX0lUEj2zyYrkxa61YHEs51s3vikmG+UGzPKd74MTlT6Jn
MHwp2nlE/YUDEwAhtQu/nED2d55KzFKj9D4Th++5fzxgFnL9b0khvcIpvc+cXh71
AtJVAqCXm54YPVM9V/95gX1VPH14ue2EHIlT00dAlxUccc2Ng8E6esyyNRWIMWMD
t1y+lalU1puj2rRFNv1r7eR9YPWkBwkuBkwAVqrEze5gA/YRLgVaOwWAnmMAl4sC
1agcPaP3IyHiDFUhBRNWwTaQwcciRS47q1gHgdPo62MsKdNIXNNGkZ7TIHl3+W7R
dNVUR/B3TbDIAvpgwec/TAuhUW+NAzmhYaZLB/uUmAjfreyy5D7nn8Pjd8aGvpSh
cFrkARbAuff0OqO7K/2DVE5b8/gvuRoI9tRQRJyAeNtxJa8NbILAP9osQqVg8xIe
53LlgXeCbEZNkn2n4lng49C+SOfY3lJlWAL7gnkC1pF6rpGbzj8UC3f5LIg2fXUY
qpK+Yu2oXwxRKLQvE5odTtXNSZwRRS6GwCA2fxbrnNpbJ4X6ta1RkloltyWhxMIe
Y38GXAMNthfvSat48OU46S9sAxXyKDwMS4E+oewgOt5ApkXGf5mC8GOarIy7ACw6
EDXOzjZ/89/XaBSlq/BuFxtq44keiP60irW4sN1Y7ySGdskTphhzQm7UgbEH3Pat
kVu4GkPvrx3z0DWaEfMzeYIkyIEYzMBRkgABZZhV4mdPbckipKOxieScUSHMshEA
FDCAJxzRjts5LtMQBkLmyxMtKGOZeo9ZfH+GHe16p/kmeDuL8ZbbQC1jdjDJsB5i
/EKP8jtpkY2pOb7cntXxqSgJ5nCDf/H2Rc3NGR/JuL+92AR8oAoAsSNSALVm8Wsv
lpT/lvGLH7e8LMjVGALcdeaqRUqlN+9S5K0zoq5kf7LKgWSrwd0KUcFnBuxTOp7f
XE6toEUT7N8xCbpazu6z5vutKKqIZxdYyjKSbrTCs9vPB5zGV9YAwcPZn3NqXira
ALU0qjOY4mumusGjdsAbeM4dNzN8fOphoLwYkHY+Lfw1244PLRCTDu3J013P3zZu
RW1UoLyO7BLzHGiUWHpPpxISgDE3eoHGvS3Y72rigvhA9pVWc1tyAVelMh1NA4xq
DxaHAhwWdfVRqDPGfCgqoW4GoF5soCTNgXWxe+GSG7M/vMgn/a0G8cs2GsNgzPAw
NNvupz9uZ/7oD+NCJdDlW+SejHWR5gL5L5WBsdgwCDjCc5htQZw2WLKGonpn6IVJ
MKosTHZx+Guh5IiQNnfrBvO1J9OH1WLdCx5nTUZny+RWuI4sozgVXNOBgqQiQ1vW
pJDc+gWw4BhBxqsg/qx8v56oydvd7ZRgIkVlIbMa9VGaRTkrKZowwyHE62e5/xBN
BzNDSYqItVj45j8LKeduVn7HlMdPzPIyR77e0ShBTk26UJmqZcwN8/Fz/k+NcaYz
5/NwuLz/uCzwrvjKNQ4ow9DdGCE/0qPJYKLDSp0j4jkpC501ClX8FZIaBSRgghdk
VNpmmLSu4uqjZPoYXoUHT4+7NdeJ4tXqUV70C1w/U2D0qxOtG9ZHC2U5A23Fum9f
QTcIvI7H/ScentlhGAKsUWb6lF0iOFxkfZgUPwCqkpBKxuEdvED2uDBLC+fr7NFZ
ixmN6BLSQ9VMMc4mWX1o0WQHRiamkOGPjJ8A5nEtRq81A/NusZQe1i/umFXVJmE8
38WA3E4oWWJO+ZH8/BnlSM5pqYeqkm1+sPhAXmHz5XIZWOpnNj3vFDYsahlRbJDh
pX17Ln9ir2joBHedLcq3SAkOPxC7BSzK3FVW36DgLdemw5ArUZxIspG6JThibe7+
YQ+zR1hrajM0P76ctlcov6O4jil1oM96cBpNcm7XT+2InJndmMy+BWlOUy7Dp+Pr
ow79vtZlfnzz5MCPs5Y6ha9Vw5jmwxpH22//BtLLbgWOf9V8U1FsER5WplD8Hz7S
M21Y+MvZR+qWdW/YZ3OJig6GmZQxnBk7yOF7gSO80pVF1uFsfpoYAwTqNxOpPcnc
tyhrzaKC28nZv6eqzmL3zpAWOZP5aQrEytw7o5bDP8JWmnSMXkzxJbdGhpWTESQH
NfF/RRI0+sTsYeQZIWW15bV6XhvB6/6Mvl4XZ+Eq9N8uBFeYlC4dK42iVANq0nu8
BnwdBsVYKyGD7oRqvlImeMVyhPbxJiKljFoxUVJh73itxU4TzIH1ArlJRf+C51tX
P/oFCxlbS9kOqpPZ6Y/B5bX7nBybOMoMC/oL53janDCSzbUECW8PCPEp1FuT+mCC
JQdIuZbie5osHpAa5pGPAdv7zinHfXQA0z6V1p5PE1kOzzY1dAkXjq9+KHHGIgEI
QTrEJZH8uO3tII9Zs7DuxoAnJXGiKNBWbw8DDuHppqNIxviaZ8+G1TCA8ZWg3LXO
Qu6v8XWUhebb6KfahIIOBctOLLf1i6bXvWTlZaQKo1jlE0bIrWyYxL6UOcCg/8SH
g8bHRAFwuhGiTwxcuY63RvhIJctPw2v2ftHGma8BVz0GcB5DpcPZwB1BF0A8VBE/
y9tHNS2pYJ2qbakxM285Toeu5o+tTsY5FZ7//S1Ls/W+E/SVbrzle57AUszlemM1
JxqELq3XTGmmB8eoMZYfj+BmDXHzadi2k4kAvGTpyppbQmSANrMpbsZsD+xKM4ju
4pIkXXP084sG2X9FEhzSJ8ZEUk1MCGNN9XnxmqIAwz7E0DgX+K+ojMkY/kaqtSYp
D7YXP2Zvvkh++VNmmpI/nV+0XbmTaSxFopqx7hRBjyI3sreeB8oTr3VG+iiGNWGo
4rLdGCOoFCNgmeRKYkRIZxbZb1gN++DAvhgkQCvQNhSNM2uDujiVMspp9EMAPDyR
ntXPERUk6rkoSdLuw6j+a6Htk5O+gLcywJ2qbbMyPHzqLFjAtwwpN/ZQ1Kkxqq63
obbD+fXD/liolCjoEs1O8w4uj6xDUBLYvPibny/D57stmrButY3NmS9Qi+snoIot
f9QEWZoStjGPEuW9JMlxFCvhcGOj58w3VnSFcg+I4HJXNLqKPMyfSEXSPS0FnfJ4
INGxjv0CtFJpiZxMloSCCybunawwzKWbCklf6vEeEsd7+p2H3CISdl7lTPozeZiJ
ZENCjHy1sa/7RQhE1mwDW8GzaNaTGLCMiujfICLl0j6Q+j9Mvn2yD8K7CqQVCy/w
HI/KYPDNunczzje1/KWFVODBKyLROklbavST7NAhT7Y7T66sDw3SKVZJWPJ/O59l
2IDJIAXCbRu8OcsgTf0L3YrqhNymtn9P/odcRmlCxkMzW39f/KHr7MGD1fJtZvSM
Bzc1UVXUS3iEL4OXied57u6HyRP76VT1PSIZ6wMOOfmptKWNKUoTImSyOpoChaAD
UJhQUwN6xxKKwDTxJhFqKeoIp6ISpzC+w9Y0pCkhcxxMlXJ3esMpnsJLRsWd0IDU
Cd96eAO/YcLdKGmHQhsW7gcg0V9Qt6NPFwOguD9yHiS6Z0N0EN8itoYV7/q0ceGc
4MmGPoSm7JG9aks7rD9veRGB1Sed0+Ub9DiJ6tZcm3IwNnxSksBCAw1CwfJLKKQ1
/V7V/hlY5j/tgsa0HKyiFDffHHdY5Z+X+YjXDqYjt4pzwQmhDmOQ3KYYfPdhAC8f
Yw99N2Z55nWfr+3qT+UbO5d5NaXlaSVwrsxPtuLeMAsokf6b8+5JMt15yW3bUuwj
umeZPyKBYrCtW78/q3V0AtUcfr1WzEXsUZBEneJy7YmqnfiAw6I3JvbT/YslwTzq
xavDF7Z6XlTN82aqVqQ+JVW0HuKwXU3TXiKgxMy0Q1XGTvliNwxhMTu3dQNU5nIv
Bg+6AoIv1t1zhkxvR7ZyloxC9C3cK2TkgC6GpIyrc7n6JLCfkSZ9L5DdmojncnS9
vjFF2NzMErbyVfhWl2+9VsAfx6+A8J2VuoCm0VC0CGjW7uoK+sy7COnTqZJRhf5F
zR2po58CUdKBJOnDgFQ3y1Bet/8MxpLgrF/A0ObiSzoreQTMnyPK1QR0XasP6jr/
8rcebJ1ohTWjN0y3GW4PvtN9xBGlmvIK96/pL9AAnCgDBxIEyrTda4Fypq99fWN1
CWBgcV9OqozMXCc2vQL1FW9OHw5/xK6aFmXjesklUKvBSZEZYSbVpnm4JJPiIfqi
bc3yADJEvNaknXrVva41FKaTQjYJ/dolpJvDAZ5sHrPZQJSMZjzCGUoFo+UbZtt1
KueJvrjJWyRdntsJBEseij+wFQbf4hENV3yAJbSTXX/tDga8E3Wkf55V6nLnI6vv
oibq5QmLy1nAEvdJUciEP+1ggMA3TQr3d5y4JDUFlr721R/XH/0sAmlt5/uxuq6T
5s1AVaw6fkrRW3/xBsUEAd7iKUvD5UW3ZZATsPQAWQqy/7+4ZMY+5YZCG+rkpuCr
kbRfwmKcqiqgegx/i/Mj41YvKaIIWCjCFsHvJihf68uswqYi5IIdXOcLsaUeSvda
QUldoiXjtKZSjGOwGmEBa3Mo+syISZgidqJ8mN06vB5VYFikeg8VjPeeluLhOqnZ
WYCLSw57TadihEBBQQWu3SjbSmvDox4kuDBRmORf1IWUJcVAfaYcH8L3yGu0gmhi
CdTLS2UHjPhzaFriBs0STFc3X8QJqBtdbpIHKDsgHK1iE3gQYIxphrfR6CaEuEJ6
pefB0QZI3MUZtjBErCGc6VJmvvlOMPeJzFNBP/OqIEI/PcfybP7kkYDwkWd6yOHB
0bvZiYTuF3gBL2LPePHB6MtjBTW9CDxAaS9M4Ad7WlLlwaXg/ksLNoakHaFREaYg
QL39YLFHhiFPIp5FJx4X1tMotF8ap1x8fI2NDZjM3wO6Gyc65HGmiqQh5oI+c7gw
OHC92zvM7U1/h/yZHFawV4m87uXXi7K0Z6t/XaVNxNVCjxSqCp053PW0iu/1JB7X
KNqBFEEL4fKf4mtOCGrjVEpiCX7CTHnG1c0waHGBCI7MbWZBdy1318eQ/Mg8bhBB
4hTPBgS4bEU0yvSQcV2WXhK30zTihHrRmILyE61ab4PkBPDgOY/70BHB4l3lRg1R
EaEt4HMW6/LRvfZqsnl+zF2M3zi64bsBDcJIQyZjQDXD5EZ0jiU0dozQJsQvai4H
nQb99DjIshZWGxaTpF+jY+OOnOuKg7Y645URr20ZMAmMjt7GCWQQvWjHQi81kKT5
oH50++OmMgyQMhHVovQQJf4THYq5tXh20uG92jEtS2S2AuxWQPsPK3xFUhSXE6ye
k6WVEvPVuF+UZojvKcfaJLfGc46Q+iwWD57pTx7sKVSFT0B2le7nLjR5HK9dE1cO
V2DSNpv0O8Eu/Cpbvl7VvtG0HuEOsKuFJVkRFlR5mqH7ltHK+lhXtVvYHuovW44D
/IXQ3L/SqaN2Hf/q1OmB8/V6/QeY8eYTu2KXo5E3FDpU/CLXUFbNTiByOgVm7nDH
3qHR0nithFrf6Fbo4IqjXmDDr3jhQm0IsEAUIcMgq66dRowal73ACVauhcJT9DVh
eEoq42dIm68GSkBhEME7Tew+m+YcC6l1G5W36n3g6fI4mh2FHnX3bXSCDq1pgvyA
JcDVLrl2r5acCVcH6F8Je/8MvqW2G/YxhRyq8E8stGUykd7vl/WRatUrX6DvrN02
7M95VggvFAMpPJe9EsAwHOyjqOMsKYHrMW/iCtSu9cr4E07uq3F2lZsrrh0htPKF
U+dAqTSw2Bnr7/BW61p8bVEyjXSrfGkOMJLRXpnUA59larmFHl4iVXAV3iHIAuAD
vPKCLRActSeKUI+Ap3rGK7DBWVOsr3Qo4tS+kyAUGR/bqt4z7tvuRHIQz7zUvIBo
WSC0D7LbYrEgW+7UjPl0H6sm9lvKNlW/aN+BMT9P9Z2b+vk3Jp+bx//aqAHJQIeu
cu5FhvuwmaZQmpvg6PqzBQrKKIVkcYPNox+EQPFJdIAguAKGeCjjyAFeAQ0I6xJq
EWN25nKpcphtSyLWcXom8c/gEd+ebtIF8ezEogeW70sQ2pstluXRT3gPwDQV/DIw
5uSzigUy9OunPQLGRq/s/cAalbVzawcNLfg8A0EiD5WrHF8G9YyvalG6TPWe7D2P
fsJxjgg3kWMRkvAAKuHX7g20Z2TuRuZ6SZxueYI4gofODe7Hyu1ucVio92XljDzs
67DdryruyLTEuS8BPp6UwhISnntZtHWH1mCRzZDQTMqCes06PNITYDeSjaAO7R5t
PJBa8p6bDB9ssqC0F50QLzh3G0VXDuh4YaQI9bO8StMQdH+I38+zgIXmuSrZVNWq
HFSzb/XX8Zm1NTZv9TJPUYSIQiTo7oJzg1xT7aDMEFdA5kyivzO03Qgmhu+E1YH7
8m6QhWfqtAix/P3vTPb1bK55gTFe22ctPcakKMuFQBGrohawAJYS/BW5J7fcpTGv
vEDU51A/aCV/oRoginQIbWAEktL3dMb4o5I0+K68XHg7qpbSvb0cnZ2gidDpwKB3
EF4kfNM9ZnjOn8pE43rQAWqr5A9rNVgc8CjWVfa7ErCtthn+0wLZeAqz4NjefzVF
5D6LQvJ14JjOYY1ikkezq5WuxRYcmGxg8lZ38KJ8jhp80Vb0qVxPrQIy2BS6kHFk
trag7V3+78mZGC/J5iOf7lNb5EiskoZkWKuP2NIlNShC2s2bSwI4jsbxdz1XncGb
pBSKaPy/EovbxqiuC6Ov9WJ8RjhEcYmEa7+Lqo/8CLTdrMxzUYXYAf5zc8Ay9QtM
cJCF6HYX4SJtfwuJwcJBd/DoCKPm6TIUfk0XbO3wJL+OarLc+LqknuseY+pG4wNe
qw2rfdKNZQt17FnyX6O0LS4RpPuhY78A0S2q95BwbTKbzZXKXwe8+Zx23XmakXYJ
rvVXxSHeweTGfo2KABXG3qWzM4+gLuy/KxZsR6oK68J/6zpJyLbuvasrywQPstod
lI752HjNIqZ//6vWiqCdY3WFBTIgRdCxPwajodX/DMhukunVHV+PKDoRVbhbg2k7
0QdCil9NjlwbVSy6vq3qVPx4XJs8x+wVRWcdBteC12KBmZZVJ/YHiGm/L4f4ezC+
QY9yXFMQY3ZLvEKbofqYuS+3bFMVgGuhPYm+tqilICKbyjDqTeruiZiFyBuXskNn
L6ZT5raQ/H4FK/YPxfvbBEBQdfjYNwWVASGkwGkFlYR/qbLSvXFu3+ltmALNa9yC
d80d2UwEzwub+2QMeS+vnZjK+svvjmmT9QkvEZdnfWF1b3gQaDUwwUAK1An9oLtD
kSzSAhAm2Sbb8S5kjs4M+viOfpR5jVZyFNOLp9PDy4WksFLYcLI5Wm1qrPfMfKPN
kjGilfQ1RSlsF4eJ9kzmPcTEorrcXmLeURweariwEFGwj3PRrpVFT0CvXgiNAJsu
I8r50RLe159ZV9O8bh1mZz9X7fZtAOvQSEwsMyHJSoe7RuhTMSZt5s9aFWY2lpuh
abho+mshwToPyNB0UhPO7ws2HppUIxTV7Z5SsWXJLoocMBrVJKGHPlOnn57XJ8I/
sm6A0ibOGNLJldQmHjGZfb8aJ911S6ntn3B2QSr0njGkD5meuuyhW4CSVtPcMoAm
V31oxCTdYnNj5gwT7nGq8dwqSaU0nvE6Hgc4ElJxF+f0bOZXekkKvzgpCOWW5Qg5
kT2PDUynuHoeqXpHDxSlTWbSDZCMhA5cXGSPceIPMWz4iSe96fgEzVuVwB+Txp5K
Sdg+hVqeKR34aJlekcd0W11Mp+IGjfSi75TQPMKcbQnQmvPN0x6v2tWZrxX5RAT2
Nwqfjbo4YZ53bkY67/lrzjqh+r0feB+WTkEpQ72cLJ9XxrCUBpAGkkQ5ZTQVcY33
jZsxaKGlaJBTU0zEKSWEGLIW4nI+mk9ZdZidJOjL2pc63V+ZmIvLTPdRnTF+NKIx
0Wed5wLopGdUDmu7AkusiGmyd32AyMmGW6wDRV51Rsm55GEusxUTsku4dCDhjQxZ
/2Lnwo4Y6/DTD14E5TQZPP0GSQsTy6ZbT+qTroCm6v0hTJ286AfjQbsH2eJot0RW
JBSC9kN0h/DvwlIO6gtMiogUkAx68NFgRCKTyWCIsSM0JZYMXbgs/kGKcKEC86jU
D3OS4+2hjNKugyNf1jobbGbDqPP+myjodknpTiiyjbezPNY3aA3blmt9/YH/I1Uz
mrNJX+5VyU27DomcdzcZC50Te3wDgYugmg1UmX3kbQdEUcx90/ulGjhaC2GZApts
mCPmPbvx7gmBAajI99jl9gCp4ku0pBzXG9sxIkUqLz2BrcbxYgYCVqbL8JonNqjE
xvZ4I3Mau4px1ovEaSIRamuLLuFt4NgAS0frrNXiQIeZK0bESiuNCaeolwZf8CjN
yO4cgLKIHlSpwSOV/7z0KuRwwhABVmF6CCvyhy+7cFr6DTHTcBh1GqI76MeUGxYs
D2c4N2mo7z1KLQvPjTEhiOR1WYlgseZ+1iOfq8B7ZN+ADVklF6ojetL+h3JqYPC5
Gb4eNEDIC6B+M7fExWjahASKtH2PEu4UjJ8fQ8U4s8kl+mDGRiPHqVRlO934oU3s
Gi/gRCavYIssqbE4zm3Bz5yb1OG8VtlCCvyzHBLv/pGJXetDLiN9Objko7Fa4YYs
JKhiEptHJ9BdQ11rrgKvRXud85Ovy+OqTh/TjU876p0eDaENiZhw6mld19V/Z2j5
VZGU8FknXTsys2cPWk0TaOiHpE6hF6cAsOtvfEsr7wJnY1oIGfLyd5hyStgh+EKt
QIp38boSPsNlsk3Fi9f8i1QK0M0cZaoFyrrJeTVnaqCSOM/gV8li7USTh5+obCpP
eO14PyqHi/vd1mwx7JopsrCEVpXXbF1JpBD4R1O1mmk2luYi1PU2/CaAeWPfZTcW
8Ta64AiWmaKGp8Y3BwpD7uiBf5n7hOhzhxDpdmYvgKWGVmngVBSy1IBnkspRZLgh
/9RdowvWa5ARV34HN8grbpTlnNRmzP8vTt8/2f+m7hLr6pHca3K9yZ/0Yhy0AEsf
xIWlIP9GW7R5jXOXUiE0VqpRo5QutOEhwuCHZAibnjpw+18DNIp5vyqLYKoDTMHT
j6J5oNGocseE1fiVAiqJ2Jw0nYM619dwhAguA6rA6PqtNk3FyjZY/ExOeYjMsTLT
XkYvHlaUaaN7HuHdwqRSEjkxuWRHFLLRtwH29ywqYb8YgAVhRLM3wSdQjYzSGlTG
ajhIADE8KVGZ4CFEeU/zMz5rXp+KfnPVnYGtZShcmsJ0qJwHr+GpGImumJs8BRD2
0fvKaDSXtu7QRbHxBmkVHtfptGxXcbELquszOZ4HTqHXWD6Gl3MG6MQenAK1VU6D
ZRF2boEm08J4vBpb/kEqAPeNi1VCBKQyi3s3xGQmpRMaYUSORWBes4rri881kH8P
AXZEiI9Mq2fmaTALl2ay65tyH9gcIsFjkKnSIV/gPJvLH/6G08rkDvQwKFo7M7Tu
l0QnrGrc+//ZY2O7qrjnofGsyhFqEfLy2SXIJRu97iq9MR9ENaGa9UgIa7l3zV5z
0tmvkaXYILtT3JoQaHjqI+lbKKMuPg/IitHgp26KGNDPbrLV6UKJmoNZaqdDjNAj
GYxImlilKAKDuAkUWH3RT+8yojf4X0wXPGzEkZqYTS0m+81/+DOlUY7GBWGLYNZi
aUMKgOuBYKCOMosQhGtQcTsppZdL6T1YTjk2icwEjUHYYm9lKNQqHf4Q1wBy+O9e
PHyEn2rn3R8RLtOIFnvNtNp77Xc8P9NmEJziRBDgA9HsOPB6tBYO/vD7kcwWowwJ
mSVJYGCp5eIxjb5LdpXSVKygUVlgKIfvA+CGxJ1nBxn0VvgfjCOqInbe+Jws5vsD
Wg4VBuk71mhfr2UoP3U9ZhJNB40h6ftfKOj5if3pwIS4hRVs2Kdc/d3/qwljfvgq
0dXV+5/7MPziqRQANe9BRzSj7doSsXliwfa8grz7OwbiP26vaMecYAdIfHrYyUTO
uUiiLtV4Y02ZGFRD5hJwVvyGOkuamVekUtonUBHqgivWtBm6IbQeNVb5CjgfpoWY
143VWpuy9CZDHZY91Aq4l0GvvXiCcVHZ6pwk+JXAiaTNMM0T6yGOHglc7ISrl8vu
Hkd8X/H/mE0mXm0ylWdV19AiHD0UWp4WqnmY+Ue/LTrMnLz7IScVcBsYL6Puk1i1
8pu7kn23Q2/KVPbeQ07p4zrFSk68wfzyJJfH152i7JS5wRTcJUNmTIA+Va226EwA
6vQnmFF9FHqP2wg/tqX4KpCfPTPYzD6PRNYuZDTSvFRruCxd6pe5l7NrAsxkbV0z
40JvuUyadYlc+4iBcABf+NNGg0ee7UWx1pLaAyjm9NSeGF1afk6CpfaOmTNTvHBt
eIIgqdcBgV8DRcr+jSUMgEOr4oPd5hKAiybq1E4OuzC9Ds3tijGzxr0yQgxo0H5H
KsNFbHqPGS2iDdDehqp+8NcJPf5X6VTqx8XEce/incUSBtCSxqxLMwV4D/yzXEUO
jz2fewqQp71uvs3nooOXu84tdGUk4zfAiJrgDCgcT+7V6hPhuYT+rwOo3osT6p1C
gzh9574Qyg7dyWNqtGDpw7CLwM+UY1DwhzhIJxVax4GctD+JHXLiPqOex7pTlWvB
uP9lSGsmHIqFhJd1vS8YibnqXzbsfJXwHRUptlmnoNnupEcL5hr7VX5K4kynckmA
e+JoVdTL9CpF8PogwLIHdH9IYDCKFLwtNPni+B03Bul5mr2b7zYBimujyctM9p4C
5d+NGWq0ZrcDSrxsFWGexH41RfwosZjT7GuLaJyFq4Stdsai2dNQpJzA8lNXy0eK
RGAONpw51ZxWe1f77bMIK5Dvs4l69TvyypLdPuTSb89ULqGC42Top7/N6Tdy7mgE
Kkc7gjink2n99pJ1AtjnnxzFxEfU0Y8s1ZzR1KJyclg095x9vPYctngnhgJ2moEN
vgl9z09MnYSXrdK325mpYuQZkBt2yR1g6HZIAidr7Q1Z86DKwocaac4fo/QZaicc
YA3QdtOYcx+2gxLbNQV5dMRhx1envIVTEjqqoizYwFHfUe8sMp0cpw74bJ7b2jl/
S8nSp2wQnkHZjiCaU5BGfMzMribI1wIhMP3L64VrlMJLMBSUBL8qmMwdrP/k1bsm
rLVFtCuOlCv6xE7IKz5BoUVDcNaXWbf5Wz4Y+7a3SgGyWV6cHtg3jYIMK4EguFS6
tL7JQeEJiswaKKJ3Gk9cg+S648b+lUgICd/Nc4Ki+lntwK+peXh71gCP3ScLz/K+
gn88Tsj3jQuNTxi3RoVv22ao7P1iDDha6+3s0sixxPisZ31+vLTPTli1ZrR1eEK5
Fw0KCCDuTuuZRAqJoIYsM8ggmullYpWlM+6PLiie8C7QFa+MGDxCOoZgfCihBAPk
0PP/5iCWUHfpVtWxauR5NtNB9a4T847rnsBJefJZUZdSma+6LBz/YjWApTYS82bH
vkjGK9hWYzAZzRgqTqUWrNq2wAHjuq0uzlk6vV5/mbc8NA+gw3q8OzG2tGjDATuO
B+NPcx0MW5VPvDKUMlmHYEMA29WVMz9s70ZCROHswW5VzB6eDB+Kk18j2C2oWYX8
KgdkBe2lVPnoQ/mIWCod4il7y+k2tTYR+J73RWBYyUI9ocNU4N+YDhejER8uTuJs
w3fnogKeHpflB40x+aOVncvF8RTN7pcuBluNfb23IfmLL0Gd8HPLR/QPjTf2Xp8s
815QT6lCeXcEiCQZ1eiWpU8xoPP6SW8C5LvueItgV3h5P76cDDOUWGvK5Npn78To
MQgxkrtfZ2doFGLn/TgsV6yzVMUlXvVHTpBhpr0z43Xr6Mic1TLJbqNv4BRIsisp
OsKZC6Rc6CRUZT726gkv541q9fphWi/HPUqF/paKTV63XXbI6PB69UQl82ADM8C2
c39I7dw87ORJ7VsJsiwpDJQOOeP3W69xxBfBTtzge3yW2Qr2ALRsSQ9K5d+aRaZJ
QuELBSoo2RjhS/QWnlBnLkqCM0CaISgjgoTPEfDg5F+Y9f6VNRoZ+ZoH2CXVIEPp
zvdtmDx6e2M5SW6Q/JH4Oya721T3pjCOzWwx2gtALXfltEQoaRS9otBbIcOSitCz
2+JCoW1HVn7JTpyWdpijF9RTBWgYCcjnKBL237EFNBiG4wK6gWDSbfFtRI0rREP+
IlFsxloaWxO3VUAyCJCHlQ/SKT39P8PSEizmg3BmOeZ1SG1vLAhXtaXkxQFiZltJ
CxsDdYOaADK5pfupNbuS/1nuug0jtgYxZlXISMBTa30QJl7kRK850J1SRrvpzWTU
fC4Pbu7YQz4FXdgumpkPCiAeSARoZRICvlHp3K3551Qn/HgdQ+2CJK8p4Qpvj8Gc
U6/pCvZu99dfOcSqY5k6Mry1QEOCANlGyeT9z2r3CtiKFwqBzgwMRZybb7uPHpWp
I/iEq+k227CkKZTLdaTpqlaJdVleavclxmdXHzx6CMEq0eGll9GUu0dDuZZk38Pq
01c4FhzeQOik6Jv/eKMAHcndNGvFofJN3AtVI4DFEQPHfQyiQre8/ES6gPR5zN0+
+noDBXG8PEUPgmnghf41airK9PB+tYOCzO84dw/HaBgDlhAhufuw1CKpNFVZXtMy
k+zpGuRP1m2+Z6gxbfpqqSuEmVgGxKEkB5S/NwjoNBTseR6s1puJsrO5yGKkyRuN
Q1MtwYrVhcwfzOWApBEyV3qtAqKTeYQeZHaZEE70AQv6zvQKEyDyWUtqTBRj+o20
q1/4O4BvXPDeiKG0yoSMB6B7OGP50cPWruxktMb6rESCtlTIA0FGRm01/WY2UxGi
S6SJ6TA3IPu7sHa3tnSasul1MyJOEw5YPXpeKUoNkV7oEFPAf312Vb1za8W9X+Km
OR5PzQUERvOpfbReU4VRBBAQhokhKgyQsn1FLucLUzfp+iaFzFAxul8jS7TaHBv8
EEbnsBR4tm8W6AAhqOoFE4hLNIAwzTiDyWurVJSRVRZPCmoi8tjZvhxc8gXPbCJe
dQAoabStp8Tf5u3WyBkWofZAWTF7bDWJiMfCS0IRgcfk0sBtFm503VhqK3o9u287
nYaLAMkuEk85zVueX6MbdRq4cNWARVCNGxSPF4JEIobfsUoTR/cU3WXBUQcQyg08
E1ASyYiNXAzEWG5yUo2U7xhJNsI1DLYj2OdDBzJbb/ROfCe0+zCCG+BQk0y4vTL6
+dsGbaGP1+O6njHo9y7qqFWUwy5fJLec9dvbyacdYyZv7St0ClfPfJu6kU33LvzM
X2Qdieco2cOp0qy41exfUmYQ+MNNNrvKRITT0pRWJjfH+P0Q2gXFHqhTRDhZcqo5
qSucl5mHv9o6d9O1xAglamdnma6IM0OYRG6ZpEbzgOHkDH6R8mTb3pl+EWIgOAC8
sTttRYyyX64MvBkrEy5Vk4Qe3pXVMzLZhKf78X2bLqFC4RHcTGMcrH/LtgmDMWAH
qVYSxp7hNpB9PHkPI7lnKWZYp7r7z+DJbzfg/epTw7YFkbAG+nOq1hazR78hmbj/
3PElw4rVt1audjmNn9wtIXyHGInoJUiRIGfIyG40y56EoCrAWHkepm10C8cyNGjC
/tzMp50mTH8Bf++KcXgYm+L0zWowgfwqzxtD/n7+hOVSymGFWtvQwJFIqB9PwWD/
kApzWCOMENNX7ngqCrxYdhTZZLKWCQsXbZ4fE3q5J5KAHRyXQLjV4+eEZwp1udio
fRRUDzyXVX+lPPjagfJ12woF2eLiIm+PiRHJsSgdVq8gyvRtJCYTKFWxv+TNaoGQ
Oz6+TcK+71WZbtS0le+KwJpAWZSmNEApk3JqJs1kvpCy0k1aiBTZBbujwHUJqqDt
vpBSw1etWHJg5UdlJ/7doXRTQKxqydxCWCID2sb4GFSzMX7TaWBkcRuV9S4UBUqV
kLkmYHpZmOjje8hjkjAUFYqB66X2mdACLhib30mevV2cQi4vs5LnImQD3eOB9TMA
8BTyZtbYo8Dobjtp9osjmcQXDVYsz373Nm+dPhd1PE+joWpPu8QYCS0abcAaLj+p
FlYe7Wz66/M3Z8GAfX0I7zy4mSttS+wmlH4Ggb14VgUbkKwKmvL0i6Wam4wfFdnn
lf3btd96kR6+oDYjJ7W+bkOwjoyXRZtYbPQmgYoKh+mzmAAb14xauDiYuXXFbxLY
bCf9cvuKomYC5aSEtRvorEzmRrjqVo7fPx0hVcAqPWN/bk1NQeZvZL9UJqt5zh7T
HeNqfK6qr+uJpM0qcJB8IzkLln5VTmh8+iDKLh4BIW4NQOllodDji4sNHNAYkdMJ
exKjfafgvKhAezV7e04csgsyF6crrZYqFLcLKYyrHmk+e/OWmzx1FKkHz2zq7D97
CL+zOFAWk7UNh13gOMUz+9rfwwLeINtTmi+qLEpQtRZRW5C0ndbocfj6e5gwl3qo
Q4kiEb/6FRahgW5Gj7r2UoYNEB2RYpWLK1g2sBRS/VMWwvFMLbEdwka7G+w5CWCT
ZO1jMfFmekVT3VvxrgPNQ9qxL/ovlQqgmqQ4QQx2zP6U2rRo+o4fcYf1o7a6/SXK
aT35y3Bax+/aZQwhKMkgJKJQCO+FfFH9ls9xudhfp2gI/om8/vtGRoOXqlDrMy3X
xXdgGheTV3ZiAxFX1x4xCw6Pzh2w+eNguGnzqDi14nLdacZeTZfbzYIO7tNu+uz5
dCQSgpEbUkpytemeA2p7EQzYE6WX7BASEX8daCAvMdyF9RmG3yUXoTTrh53e/FG/
g+BJAqK0A2KeG4yVksORTeGJB3p52K8Ylwp9nmKhvy690TLv6fNKtzaFBQMrpqUk
44TEq0L/2v3/49+ggXGzEUMFVsV8aX6C7u3hosI5oOiANkS4q4qqK7xQApc6TStW
pcqg7X5xjmOlv3aQdkc4XPfTXV7byREAfkLi25xa7POT5DjYw95VKEmKBqNk+g18
40Kx+AkwiTHlnuJDyrkILrl3ofPVLowCZRRtaj7aGNUVbRzkjZVEe5uffXc9mDkx
wagPA3FG1mQyRbTCsEu0MXOIg+yE58WdqoB2Co/SPhPQQ0C2mUirSOJWrt89Yyih
tmQk9nfN2f1rcLL2Ff8WiqNAW+/sGxhI5itZuj5Og6TFl3qKKXeqLzCXO8eXQ6c5
e/4yCVqCXqW+5vaYoTeQCdAMnyG+eLv76diwP0kgIsn2lWeSqSJjjJXS2F8IA8n0
aV5efkxY2Zev0flIH/rlU0UxC9u/Bv6+onuvfXY6WHJL3fX7D4BlcvFQuR9bVhgt
ucfbYm+eeBByG1sUp0w6ICkGpU4cK9uhjLBeS+lnc8oUB8u+x54wVpg0Tp8ysfUM
c/FwQe076Iioalay+B6QlOGLZH0fDh2FptUnk5skxdcL53soGxCjxqW00REPsyUg
1jU73tvm7EBp0iA8NqbWQG4AQnf5pFCssyoHw5jhS75D6vm57Yem92cxA4JdM2Zt
OIGlrAPRKSn7BmeKlZdSS936vH86vOIYBsZKeRxYA336RuQcMIiZ8ZO97/fe6WDR
zpAl3Am+EvHvtQMOLj/9zlveWuPX04Nh0y2oDqsWAtNAxu8L9DHTZD53WUyzarI2
CSHxyzpRG17XFt0AV4LhjLYN9FGjmoHUFgVmO3cuGlBle4KKtfCae1FJzazJKSN4
y9uetjgURXuIBgl2WPFTZcah2UZK+leZNCaiyi94UreW2Sw4fypm9iS9ImbY/wX9
+KxYrT/Ki+Pm5DbCXAYR5t1Zqq4dYfaDr3qc78FB5ywaQBU81S16Z5GXy+7ZjrEN
M2S3FpHeUYb9cUWryrDv/tP6gynY5hwxyxZKwmKh2f+qZ3E2HLDkDDaIGp+aJW4g
jmk0LSS6fSGncfA8yPYoZ6rRpbpyUWcxzyzY7VHt2cmROZ1Y180lB6UMjAk7oYxG
H+b2UDZdPm0LKvMvZgEZn9U8EBdjdBcwcl3Pxh4Wltmp+WLW9DTk2U97oMpddOIF
eah56KCIaHuV/j3cVz4ga6DvV4t7yY1bCGUVBhyUwMjMkr6wsdjJ/ix+nKbDoiqH
5amb0XGqwwPFjGmcGFhei9f7lwJfd7q63bo7y1i2qikSIlVxK6w5Wuh5Ijfw2nqe
jHuJbGIA77/jA39xDKcTzZJeRhb5+vG1xrZ37U8yggxNMIenCUOf+JHsHCpa/Nff
+G22zcENA62mDM7a8dN8q12zbHMERmPQRwDiOfxWUcznDqbp7+6toA0V7wKbNUki
o9BxgzOtnM7vcamC1cwDZ+QhqukrC4moeTmm3dv9MKQLd5tThGCPlqNOBr+LeKGW
Nbw8DHNrLE5gJiMNFUGJgEw79YF5xQazbe6reQMqJxYYm9feNZ0TgDAa1IAxtK/y
PFayuqH3rW3U15HHlNvZUMZvGL8dmisA8ZgXHm8hszg5PxymhJJLVKJNfmXYn8AF
o9ASMkEoQdZJ++lUFaeYJVubpZGRLuI2rk3UKbPidzU7m5Dzm+HwvQPySnbVoY57
uWQU3NBm6EKSUHcI7ah7ceYhLXHJbi094BmyWvrUercybXKZc/Q+vV2m7DrkYCGY
JCeWzhclaWuzaGfSL+/PNXzk+LPzWHFbjg19+bjG4M7DjN8/CrVnSA/yMWLbdv6+
7OJ4RRs6lRfd0cVsuMS7T5RcxUpMQyyRNCaqezubDJOvbhe57o9pFRDF/5MwSEVr
pL5gqtWOdKH0QOv7ia+QIH5SK96HF78HP9erxgXSYgqXyKCSOXmQ2kkkslGB4uJz
3pLPzRYxptDexOJtTu2VkUs1h1QIVut7uHQ4/K9WjmMXO/6JnVI5Mqjapi1Qz/xQ
Ibwenz5Xjk5hwqtHTKpPj73+FRDs8Bdzv703snlvFl3PN9cZluWjNm+nfxcy/EgK
GxH6FImG9v3hju2qA2gx4xP/XPonaUnkNFDX7wgXnta1TxscDV2sWlanrAek+rua
Lux94oHXAEYZ+ugnZ/Ta5kHzRKJ2gicKRlFMH/+i41OAfA2U54l/yK3G4Ysp9wtm
4vuzg/RR4TzQ+wH34f1E0K6KvfDrS19JpkYfYFc7uxnE0Y3Ek7fgeFStrS0MYbEK
FQ+cPvifSzc892+VCNsBiu1cxHj6pABK6nrABN99G1brsPf/GPcAP+GwNSLlt1fu
4X1x59ohOiHXnXOt27PqQpDwxI89kkgTVy1NIuFpQnBgs8jcTU7Avzo03ibMNRZr
J7v2kLLS8iNnRonatDp7Y2dP1T1179TlV80Lk8ESWojoX0bpA+r4TXNi5cvZvFw6
6IXJRo8rTUslUwqLBjqAnCqwXl3WWEyjige4iSIkU9W6j4V4YvmgWVkEr/qOMt+x
Nm5JPTOly0YBcgi5LnDBqKZqesL6KJlSWfAetystrQ0l4yv4Fgaf9f0a3Qeg7xDj
e3NH8+q9MAzw8bBeRT/yjqiv+kkFJzWq5dy8hIe2nV5a4EG2DRrcOQZn+4fkFjJy
Nh2+07UmNeF6HJwjNA9VmUL1PK0SXQy2bv4NAE579e2r/IBuPVmkqFtZ63iSWahN
t67B+fweW84nMBZKaj0Jatd4hAROxttFtQRJuKkCUBJtOtxTRCeRjJ0Hg/jcEnrM
2JxGsghK/sg3R6BwMjXoPUCIDIOaoEtz90e5Fy/Y9tvFDcga6/siY3UBgu9vu34H
fW6YpSuGHygtKJtYkEdNMK4wxBVvlkFacSsd7nFkntSGQoI0XcTf4vqXcUJuFrYq
NMUfLXQgRUVwUsgZ/VerLjaZs2sfcC7PDLW7i2VRfTOw1bQQfAoebF7stfTfd+8i
gXw7hQ7B/PF5SNqV2SrNt8dvBOgSy9FGzDbGCUItuw3XtUOg+b0ooMNnTRGkc1QC
Wpp8xGJX39KnYgUvwXQVbteeyxERD3oqJLliCsx6iqZ8bKzXNRqXlVWgZlnMet/j
rseyPdViRFp9Q1OiTe2u2Fky41ReFF45mZMPOxID7ruqskkxUVCwIL11zTpO74lA
keFwRQTApb45x7pCZRAZDL2QqSZZVPMRHkj+uhfWY5mwiKLoKJw/8HKBlntLnOrd
TZ9zCExJWu2uEv8qboMeNjVG32qpLMZQqPkpkDbOo0U25Ipz7u39QD0c511HWWJX
ux7ascbzuhxyP52rwoyF84RTt7yFk0incxd74fM6RwBjX2UHjSFhvobTy+9G4n/l
7AuxkMcBh8WEadNU+U1BKrAUqBntqMDInrTsJsNWYlX+PYvFo1vnYcviceUx7abx
IWJQ6zGIhEywGwT3Y8bVFVHckqOBFP9Ql0LQP0lxO/cWLxUISmYIZMheiagJ91zW
q1gCpUBQ9xD1//uUFX1KMQPdrLZaI9HtWCTGxG5EMOZfw0Yo4bIItJ91SXbXZHtJ
bP7CiQh1OcTGa0CRIQikz5Ky18icjSgdeu0CNV5FJpbERMbYML2EpzSP5G0iAWF1
PCKiCnCqoV5gGky3AbRXmMYFnkrowYpegcp9xIBlpVu9kYpLwEf86OBPaUN+Sc5k
Zz1pf9Wrx6IuEX+ZWdIcxl0pIIJcBdh1VA9qP5upc7viuwh+owx9t7BreA+ZPkne
JQgBxbv+oQ3exv8X2jo3OfqI/2PO54Fvh9zlUw4OehB76XjkzbZIJjxihcjjIrj2
JYAPZO7a2uMEoKJlfF13FeoY2IR0kvuKa3E5y7qYYFitxFaMUVWqbTTmAfEOW14y
eZj3lI9m/ER7RIEsDPV7RmstmBm1dcJkk4Z5kdOBYd8JG/WoSjwpu5DYOEZ9UmgC
w2oOa5gRrOE+8o9IAIArWpEXzQjigfShpLb5iJGvBKs9cYc9ntHt0aGG4hPucOKs
qksxr1W9W0x4hMnsv37MqM1VncA+g2G+jBOpolmQABLMXHmEvrfwJoP//NdRHi5R
xAN8nC7TyP6G8ktj76nkpyXr3AlyutaxMcl12zp9oX4eUVCDj+soNCTJ2cZLy97D
wAxt9FFiTQJwKWqMEaRX0giOqY0Hiuyhse0PoFATzDqelGrNWMnGGnhV+Cvggw62
zVR8A8F3svIezRQ9G1hA9/t3qCJ4ArVh6nrTVnEWWyFQ3XAhWDDBEiYFEzrD15/l
Tfaoh+fN5fI016p/D8VL0H66QvZzzwtTni5VAOExbE+2t1ZlTJWuRykp5ngpp4Zr
2HRd7YwbNtVqDGFg+ryzg+FQAOzgsyGZ7TQ+04LMCNZ9DydkD7eeXnw3pb9SbG0v
Fcisb9YkyJ33UjvbZB5MCmmQyxoX1UB8WrUlgu9QtMZbnegN2wWrr99Cf3mwc/Fe
lG5HVt0PimsWNxC7yD0uC/zuohlGKnQbbWDotOxdNdvVd8+k7LAJIFZ9B1HYXyzW
VJUzZRdv1fSomIKEicEpV2TVS6MBnFjpr5LjTPBO8JQ7+Gx31kTYhzKDuwfWVKeS
S1Jhn1mn8ZhYhrUcfBCqAotZN6DZaUKG2N6CQ/W8k5Z/KaXpo2zgZSBXzLI8ESqy
gbXC29YSHW4BYq6mL8ZUB9b1OrCoOjHSL2wtOoJQiLIPa7jh8/ySIsB6pPmhkpFz
udY7HmMebI2x5b4fSOSsVEQOdIacJc9PK45ysUIJKt0L9J/oQ2F8G24EEu8gD+Nb
YxyarkWcw+OcnWrLcIdZXqOhH+YZvnR1hltki2sjjVWfUcCf/wCEh/j7E7+QzBVR
cRelaVZ8mMWRqLeuVGlANW1yVk4d4ApyZllpW/kRpmjjyzW6XcqoGfWS9QQspu2r
G9v9Y6QtTdwWDS/IuWzLRIZdO/kFPN+s/QS6aPYTyGwdXhI+jJHRkxxNnCd+yyqm
+ZtIczmYdBn1Ak6rEQ00QA9hioZCKf6vTO+sevYkvZB8uwj2Ow3lQmE559eQdGwh
IVoOxmsYFUcF5d01ecNEtKB+uovwDnZScSz78lp4ABD+M9mbLayU7QMmm23N+n5q
CQ/Xe+ZoNpc4oyile7QX7PiNV8Wt3KD6UjUQkwmiWp2zpf/aLXrTca1nOmna9ldY
6VoJ73+w9zg5XlWALnBaBselKx9+Qk2LtoJbQoPwfBCnvU6M/DcNFnmgF6ObtWBg
Y65DRVAXxTNRliBEETlffynZ9ZaizPg3/cOgLiBBrjO+EZWipiliu8gybZcWixbs
dovZVE7vsiXA5JoElFNA02gym5r339MY517syCJxWkqfKFYhGuqHA5K+F4bnIyVk
ttHG3/3+G1DRqwttNcEXqHHtTbsSUu5Xp4iQ4GNZmYTDLQj+OxLJQHKq5rnflihc
ii3kEoSjBrpC4NDPIMKbHyBwPoiZSAl+hv7TmO8wrgwQHTXCVot9hVFjmJExybEI
YWOBW3fjl1FUWalPeImt26PkHEkBps81zN3RdnEQ5Ee7RbksRX0O6wHofagzyDtk
/iSDMKeh5EptC/baC1FjRjMUd8ncXRl9AYerZcId0QPB1wnjOqlSChSTHAoQq4Z+
mD412Ey0sAOInI8RXf20Qd7s7G7pUOvzack1PVsz6ZAy3maDAxfQ1S4dR672CPRw
jZwZFsRExPxKqx6Zc0yZggH6Km0ytBFkK6hi21DHRgIo4Szbnno7Gp+/98uTMXB4
Qx/L9o0c3Jg60gRnzQwr1W7B6Gd9JLEBKkGJg3dZRDU7gmhmZrzhJXsOMeKDNSmY
2smUC7Rhf4lhIpKvkE88NpDIGJUlTF0RmVWNXMad4D9dSfuJ2Ct3xBX24RGBZXpC
WtSaS548fe1XLIAQmU0a3FU8/QmQWDeZd2tVwvc/3qEs0ljioYyE0ObyH8EKalBg
8CaCUuVco83cae02Qz/21tENmS3IKfQtD/T7HtIyap9BPp3/pveL9X8w7VIa3DBB
gNICxSCHwgAX56RKDOQZHzypyOL6nY1qVEqmR1X0C5dLSymTW/+Y6Hq/WEG1b1i2
PgEvTnij2/xc+bVrm74HngwxWfecwvwst8PBDfolucpZji48MPZu56SYTeM63kJ/
oKrJVg6ANvCBf+zl1tG2oVSbCJHc5sS0yhyh4CwSz9CRNASIDkYx8A2eXvCHAOwb
eJkCA480sTi70Q3gLBsTmVTfwegzBjgcgb833CzV4iVxDN+tC1ROb+b53c5HCwbn
+MZvwvzMPFSKkk4LTQsYDqouxIBjAvH0r4yJJIfztNuynxKN/ydLtVNfUTOsS8RA
bFxK2DbC4nOptdfsj76pbwCI+LBYXBls3qW8azciPr/5nfIkHMivEVDHs9bzgg0W
r46UTZLYP3mMeQk0bvqJDnH07M1K0MQYTf7k8+IUJq1U6WQyvu7jM8pR1Db4bC93
UkFUBzam5deQ/lZBJm/2pHJNckyUONEr7w4C2XxxMbBT7dUGwJ0bnPmUiQd/JBVG
OFT1VptMi6Ino3CyWRqOQq8USrcJpN0JoKEvX2n3su42F0X6Gg/xZDfKaGa3hliX
BP6676vcIpbC3dPg2j3n74ASe6Bi9x1inVCqu9ypM1Dyr8uNYxZJuJQk/6+uxZrK
YAGr9+v5nlNRAtYnG00IKW0LwPc9q2bcnh8Gx1GGrtb2E2+gX4c3j6Yafx6xhrl6
7IR8DTN507eqKrQeppcWdHw6cRQ68vf2HwlPR89cH0uh4mR75x0sVaG4KmwdJDMS
wrvNn9U8tkGAR2kS+RhbjGVRb8V+vST7TxqvQzFSVilXYb3gzJdG54HYOKP7tRqZ
v1ZdhBGqzwVLBKdP88A0iNymkzf662IqJxmygH1XK4Z2mNFkYue+MJObwQl3sCh7
+U+/aCVy4rikR8U72CTLrIel1KMNXMVWQxofZtsL/ICEpminac4PxTUICeraJ7CP
c+KTBfxN+vKRsGT62dsg5V5eQrRpBoWKl4KqWB3rWs6ovSss4XIX466veKShl7nw
9yDSVSH7agJjhjkuqcsNOrYmHq/WL43TMR2jpgZfnOA5toI0BTJmHDELYhp61Uzw
M22c0TuI+F06sL+WHryR99FiYovnLdPyTtswUsgkFlwlw7+JdXxGeqpQoTUdPerq
PmmUIvcOy+y8SIRRq5STN3+3heUuKS9h22HQ1D5zySSa7WyeZ/pmJxosw8f4Y6mE
51r5Lq//qjcBZ/QcoSBsspMN9MzzquRlGTbi1Esu5eMlCWRAmi8P89yk2UKlK6Q9
2WeOJ6huXv7+7io9TC+P37rV4Q/+vq0G7wWoL/KBAyQ1Bjdkdp46DZ5LZnIXylc9
ER0w/yS/bqzRRSMpu9BE5YBrH3Cut0ppnQfB/5b8kGuYH0ttol3qVN2cw34Mw5wO
tU0SzO4xBZf2wCvr+TMMuV2GlqRZxa+cwuuo8s8lXT5WPxXjY3egX60sH6B4GGki
gebrP75eSmfNkPG3ST3VIk9J2rETBvJP89lyq7UFjsPtmSXgfMFsRQjrcr5NA6ck
MewgpDM0yAMjTu6hybm0YzMBz4BuEjf2JfdtD10qLSC6WVm2CNFuZkVbMiKkoqij
avKLKbn+ETHYkMPRdMs62YvRMODiYdkSQrORKF97MIU8ksnYTQ8kPzHqWsjBgXCe
MHZ5VjvbelSk2IZ8Od5W3VI+3EImZkE7KBV3XlHHLuPUHnvE8xIVflRtc2Tpd6HT
6cinGzM2OZW3BqZPhp0Otn7515GgBAmCjAWndd/KHtElcIbHeS2nnGS+eRmkBgu/
wMrbZbwRepmWw8bcywwAjNodA0bTpn3u2G8lN3SYo6G8jLJx+SSxhQVjj3EI/ont
dAkE8TiEGag5sclSJMDwzeAs+eKzZmjIXaGtPzdrcJptkIFruQ3lB4hYq+Vl0L0f
5eUpED8XtI4t/vTP1rnA6zdBGgdY8QThOq6zzL++t+AKXOjKcMOasRUjx+/L/Qqn
n1lOqCRmUYc3mpRkROvm4bzljB75u2UbOkI4xr2dHg5nUl6pPFZzGE8aLu1kUwVG
5PhjJAeZq08UOhPq4+6niyCBCMI6p9LaAmR9St671FJpCAWvDcdqhZ34Ontt+gAw
i1a/pVPqdQKd4SvKE0jRrh39Z1vdR47qLz2I0sOVDXocg2xtx3HmMC0EI6BPzteN
iUYhBsl/MUWJu+qTiAM7n0SjleYCmvSJmS4Zp8rbTIGY+fwHUDA2F92Wq6lcJWL2
0nhzP/7MtiOmyE5Q3MGLpCJsNaiZZ13sZs/fed9WGcvI3ETK2KrN4p+5Tnat8m2E
0C19eYA5utkNtv6gvydwpVqu5b/AHfb46AgKozMi+706If/zzCg5Hm2nHjavT6IO
TRmOrkI+Ftk85Rtvms/9SyktQkSOkmdUbTgmN2YWacREr8vx5R6wYZjZ46L7Va3U
GbfXRvmwmRxDZVHL1x7pu5jo/rx5+Rdv2lx3+2ZKqOIGEWvxPaizISRJv/ivozr7
c3NJDqgISJZTYLMzFnZgQwYRtDgXfyuO5jQmRR7FlFWab9BJGHWlipZ0iHOKg1VK
0TAOFFIjbPHJkqB4hcesN/ABFhAH+zCZFpc9OI2jrH/V4Qcti//DsQ6lOUQVcp7a
xtfMYpERfcW2XZBFInEVepTqPjpKF656L3ZamjNAhgZtY+5q8ga+mR6vVptKGdNw
s6yqMwir0G5F1S84Nt3UAscJvMqRmofWz46EplU/KOyXkjTAeC/zsqI/20FVih+9
HKSs2UvN/f2HMqBcHqGuF5wQ471gLx4UnnF9DfqdAnjmNQ2YbvBupZs9SfrQtAgs
odKwkWKephXKXMLqHZ6VXqdAFnL8azbj7qO1OW566sIl6qbWzVGEEf+s7jP2DomA
PO4/T8X9psNE6UeuiNCMZlhNK7DwiPy+cQO7h2B+LvH98pZjhgrVgEZm1LKqVS26
ZD9SoATCIkbbp1s+o6hG7LRUKJmiQC2sR42J5tF16Qhi2aoI9k2QWJupWZWCeo1o
VPMHUtCewcxyIu3UisdYpDGyn/3bECT9DOM037Qp/BUURTmtcuW7YhwJoqvcNVzC
oJ/39ZVLqsoy81rdSi+9OfJBkCTk909+y0L6lTfXJ67nwwwDu+LHPdwPkS+n54dO
viq5WclfWVMhqxMaDJzNkuV6XddpyPMAOIRQY6zAcL6RcT5MsVnclwmpm5+/T/Qu
3VNIV0KAbBVWIlRl0CpPSqei89yfofTZd5FQjMNUMxT4pqFMRJsfzy15/VaaWxBy
rOWO1kelBJno+vJXpt0JKtubhG/VAUXMLKINGCYDNYXjnrCQvIYKdqXyvHaH1YyV
PdFQLU1HeJvfsyfS4kSSZsTK/YAO0lZuIWGlJ7VTnIH+qF4Vr/zrGO8oydDd8h71
eOe+TDEMI9lV7SfkrX8U4AaZ5lDRtfIym8C1lPuslkqFBPm3YZ3USXbnVp6LUeuS
Ohwdhz4P/R9EEAViLD1Cqb6I7jKllDTRPe6L9fKpOJ/vt3a40yBnTI28l70Dk+tK
EQk8Ux8v49NXUtWyX+r/qVuXwR2Yp3hVH14n80PgiWYKP/o1r9fC5OwWvLeBLT1n
T5sBX03TxSYLSbNOnGEGD3QjkB0y0ynv0E4GMLeAyOBmByvOwjCcPFMRaV6+J/we
6zwrYkomxtQNYsH5rTe8EvpDw1CuHaacPQ8MF1G0fjTqOitJbQ4E3ItMYfYKfOdR
C8rqX7m8baetwdSOtGo2IIn19LvJXhXyIhas6KZQjpH9RpxXkbQWOnQJ6sPLPMlf
avpyCspqfZidYSfFQgUMlJSzRadUgNy1zALTkI0M4K31AJim+0GJbRYuXiQ6dAWx
rbaJ8HTNBCDnTMs6/URkBuJ0X4dmJXUFOPR+7sr27RywNwXeqzcgs3fqC1TP7q/N
cLuOkwSpfRl7x3SDV/1D8NTkajS6BnUdNSg1SrHsqP4A+dMZwBfZAJlbbgcr6/a7
cCEdsjZQXPAQhUfegycfHV3huSC8VCzaN+TEQ9673IgCJVqGKmVi2FuvwyQiwnoT
t7I9FvBRkVdV943ETrNM8lo7kwxtPv1dGxYMAlh77715OekM+1TS88mFhmMyVURe
8zrAg4z+ld5nPk1qZuOUe2VXsIfYW+GehIH1qLyHCJSp8lOIkpueOD/BQpf1+eiZ
HvQ6AbV6h8RbMwH9x7r+Unb8Y7XSVKTT2yPIH1Aqq1ntSz45pkJ9nlHJhnV3KQEn
lKvXj8qxEkC+euNGtb1VqoPKz+W7HGSTC/uIYMjd1dr4iPs6H67Oe2FA6hjfLYqR
MpF6Zt6ZLU65DxOen+/+FyxOwgkHB+PM/OmDK3mC2AHHFrqc4gZ1JnBnVKX9QZxS
GR//2ceNgTXN+zooOGzwj6h1Go34wjZlGDYE+yK3Ttm4Prw/k1Bby1BHhLbygFud
Js50JTBhT15V0uBkpJEaKZoZL1VepOm8iVmeDSmcXfL3hJF5QIcJY9/KXKv4HRi8
0/xoyVjs1uu+lTuU4BLzUAf8I0LnQB+5kMzblcc3n98Hm7bAVCgNOz3f+HIOq6IO
emVykNCaqXlB1zaMeEB2HtoXPw7f6QUQsq3JFE9hmSD85cKg23X9mUJGnsPVD3Jk
rpwPoEfhxomqiD170ftVE86E7l42Ss8/ss7OHAOfy5FhJPlsJ5JE9T66HklGFJ+A
gOysQBfkx8SKqzvMuGc5Rl3e0rkaD/P4v1OfwUxqJYQ5w8/V96dYJhOIA5lZ9ZGe
cG55VXaWfl7D/4y7pvNgU+AwS7o489PmH05E+lehvBChE0VNLEnpC1hCM3D11rWf
M5O03a7by6y78PXCBgMWmsKtqfudxIPungMRS+Gy8tyz1CIb1H04ul/kLLEIJ6fQ
ihZIumVTAdyeSg5k69xREtAow7POeKgTwWIuYDClu/KMRmprQYMgH6R31nVNfkOG
/M4huW/U9bHODY3lt3xqA04BvbKsOFZWWadrrXqGs7RSoNFc2ucaKBR+KjPws3Mc
KFgJCWlG95HLvgigd1yOQEAzV5gjmckg/YSq+20G0neL/RkhXW9+bsTCgMk8GKc8
GdTly3Gxr2hoZ4MVBjOx+R0qbWKHd0a6PKUFmnw9Rq4QUUf3GhY7vhVDFtVaGXX2
FBbI3Qym1QncEIAEj35Td34IJ8UHI90Qni/5kw3pWtKpl0uiyvCu48HDMRixgr5u
nzNkMmRz81+AHjprMO6xzh7iM5yNW30c8gyk9vHZuH9LMT75ZsKzKC3w5eRkpO9y
PcJa+qQy1/6YNLtaKKNgbzcpacGnnzAGctluNgsAWOLG0X0eVCMHmILUgzvCaHQH
1LShYqy8YMF5S5yYeEj96YS2Y70t0tRpIW7uo3IGpSk+SIMrH35JvQTtGIYjksPe
nqe6ctLQGN98YyZvesSP7+68C0fVo770k1CG5cwgVzTIMHCIyTUGVoJesRok49vX
tqvI8CGxRUCP8khprWBp08TkCWWJFqgK4seJ6MXhPR8Me2WW1LralJRLSqg1yA9J
FYHHbFJ4rbb2P/pgINXEI/THi81FRvlbSnDhMz4beZ08o7/qamMRokiIscWqqBrL
BLbbueva2FQrLz/knP6AUsfQGYHKcy4H+cDisNXE7r8m0fz2Oy+HH69gg1Betuyl
dKH7iqvC3a9lk0e7kucOFRJPcS78GCP0Sjucpdzcup4Z7VoHVUevbcsnOWjQKoGx
WTc6drDvN3LdavfN32vjo2s88aZXBI7iF6BHs2Yd5Uq+KwbAJKDU113IdOak0CQT
2t4H440Z5LLiH12d3SLfJOqZnIwI8wdAADWxy7N31bF8vka3Z0uCj1tc+WhcjBGf
wkiWWuuy2402NMf6pUZc31vLDXP13fC0+TRMtnQMXAfR2dW+OOFCAu9TNQhQL6Fz
Pg6FGSx0B/tNRMCJTIbug8E4m2U0pWv7bM6whW9HKP49F5J62rDsl4eu0aFSH3Jv
eKcRhzawi6ClSMQutcccCaYq3uWf30HjhZL09ibLf8Qa3hQ89M/mqizIlsHRfHlJ
sQ7o9MpvPxIUszDN9HoD7qn5a+WLnU5u6XT48fueLYdlXZXodVqjIlbJ+VLAwXoN
+/5GddRVJH67c6eCJbu+g1fq58I5ylxVS5aN9imbmNiHyqJClf6owKlo/jUdQpTu
pbUumsb+ZYSjzCSBy+590KnItpQd706KwCQAX8WznZSDvvVq+vanWuXL/fpl0a7b
uvVedyb9wk9y43KTRUk4AogFr9xuko4r3kyOxa354nfs2wIx2isZznUM08zUjgob
nnff+0MOB51roQIofvHoxVtLavIzolnexmHb980roZ8djGuSGFq4VTmT2IfqbnYL
tnEQlWzocTp7p/cxL1bkJpB9r/FMexB3Ge/nO6+80lpEOggVX6dS9HYp0HJN5zMj
0uVjlTcllwzRPBTmlicYDM3V4h384/KZxLYIxInS1ZpFZ3vogDUq+i/u/EuAmm9a
iHkvyoX8dNExo58/j4GUt+pCVIVH5w1w1/dEG0zkfK9GMJZ/GRbG5JCw43upF2O1
oRGyXib5RIWeXeCx7dLLLbI8K0z7PP/ft96fJfRVmrb6+LF2C9PPQbUpOq33xa4f
/gcGD63n722X8t958v6frt+iJL/345bEfsmE8z7B2rTjfMRrCOwHVnQFdCvPyBJk
pxCbrjrz5HreSxP+JWODmABayb8ZU6qoTMhipFtyeqLH2eGo3em6uOpIlJB/NJ+p
4PZcNNibF/m1lZO/7SL+LECo0Tarv96oSokikQ6+PI2xMqIgSR8Q34HFafoSPwRw
b1MlmOLcpH5j+VlS3X7nunfmJBgLoDXRvnxxecHJQBxuXhjSQTIKPS1uIb2Yu2ka
SCLnFELyUqjjYEI/a8y4B2Ewdor73/Plb8T3BCEZsU7j8vJtkdxP93TWy4TCNxTZ
WUsg7Mf2jAGEqt0+kuDxoonmPecQ+BbXaVJrc9LatnWUD/+iOiRh0YvrUD0FvlCs
8LmKF9JldOLib8095n1mfR8sfJhq89NTvlhzGPMQ5qjJx1Tn99M1zECbMxVuJe0Y
aMRKZbGM/O5G5ytXfwtaJMz8Wx0ayqaGU1nKk3sgQf0IRNmLMqDhgKUEzA+CEwUd
Yx270h6LOxXcMCSKpqIqS9kTvVHbsn0ePjr3UsLRa2tTvH83XQxTrWcQBexmvVJc
XouExpDeRDGO/XvJ1f3q0Oc3+ylLEO/MF+ZCNwNy6KWNeLtBcs+yJxOv8W7+oo47
SRen9LZb28W5VVJuoBPYI50oF+RrTF9vViC/HVt4xky2UK69Xr8h8KQHn08fBcks
q5mBTnaRgU1VwhwtABVczO736o1ZBJgWZj3vzvVPgHuQQ1GpfzMKE7cRqoKip8OM
YRillL03GupqFSW690CRirBkSUwItVjkdcuhCKN1zNo2L4VXA0KzGTVzfjr8KZGg
0A1C6x6LprI2ztTUbcYKcBBNyiUAnVxy5C2PY8hLDg4AYOn+flx6GtQ5lRvUkAxW
MmVLvPAKVUSqq3DjYSI+V/q2xzkdY+yHgN/8sgMO6DPIs3gHS25NvNxBj1CgFKGF
6ViYRv1HXpP93VS9m/K9dSGEi+D+UlNPXTPV84FPTSeqi/C9I2AjUl5lYfXsNPvg
mMyfZ3re05k7fKrrlbUBKzp46PThL67t4Drqo5s413uJwQdct7jFdSdGIZXv8o47
WhE19i3mAefzuNG9hlRF3jiX59/wyVkTGNeTHK2VZhzsA5RIWwmP/n+goE8zwkw8
N+7gSEGuRV4bwWu1fS1IXljOmLUD1+FXiAW8diCQrSNXMBOE284cm2nl4bOAHDt5
i7nnvmxqQqn3ukSPlt/rDLRBarlW2sPOth1nL+JeIcqXGbVyDXEBT71rqpNGNQnQ
G8f9xcHe17G2nTWphRIVScdoC27CPpf0CloZgKTv+9ZD4dSVQHXB7uftI1IkeS3S
XoP/062cWQMRakKLH4uC3aGyyQON5XnYeq2vAunKB5lN1BXaZeR53Mv92/kA/WPe
qFRB/e7M7AmYVyj/rRExmWfTsQnO3EAozwlA9PaxS8M7OaHNlMyp+gggg39WI9g5
LOFoI0k9WkoCowDaQ22l3NK9OxpQJ2IIpwFlcvDzHDth+BCiACQAS9MIn1AZxVDl
IRx0m7P5gdy9NDtuDGC8yyoRok+VKWkGfcHtlalxbMMX7dpJu+4lj15fvD1TfRG4
3qqnbophbfdzn6Y79EDELTI75OuvZACYsIx41SQlWUaORZ35wUROlwOs+PYpzwb7
vbUuF6h45lICRGz3rPzL9aB+liG2ZWIUSKP3KeQBqsle6Ac/lSnXyfYtB3nY2Gkl
dzDesuwmkqqjIEQOPGnPFhhHvAn6MNeyVoB1SKCa42lKb2UbkNuOhUZke529xhO1
k3OMKxjezHClSe//Jq/Zdkf4iOR0a1OcGRi9akL+OVJcv0p+NwBr6HLwEZLZ4U3z
ZQAAFFy+JGejhCSHHUo3t631fcRrrOhGC3dagRYnOMYggVes/WpRsjlNP5B7jvYr
EB5ToBPOWqGkHpGD5eBEqKPTgvrvK3O/lJy5FNyzf4cQZIAKPIDopoRfBpuRjt9i
MAK00lJOnjCw3JHsNTlaI5oYHziqW+tr9im0P7HvXZhOL3QhWm/znUkvAuxDkcWo
tnQpK5thhMxZXsBFi3L9oYNay0e5c23VsmtwlhY8MrKcVzbc0cWsckS7Nk/p29sT
JUlzXOgjtl4ePrX2sPlEfL3mXRlJ00/QmCTy1LwhVeDkYVu/ej7UhyK7txnJajli
meLAPh2BCuFwN1yBJIIAEAmsBfNQ6oYukgyFSgvCVt64yV3S5t7FuWzha94jIBLa
vYiNJs0/XmgzEKg73udkHbu0rnWJ4r6ZHl+mznYVZDKzBIecqd4ymTMGyufi5kfH
ZfQsVE84eSnW4XI/Fi5h5ZlGqTm9H360uEWX1dYY/5S6CvU9WmNeFoTVQTBbx5UU
FazwGnRdVvQjg/AeycTjhzCpbDAfibNmoOxYVkczt0sBRacCaFG9o98O3SZg43si
Q+Zp3XW3IhoG6XgQdI6i6W1BF8W+wVxrRu/G5L4lQFivsAJdn9/eOTY7BF1kHAnp
EEWyyr9m7RafWFnitQP8J0aqvb0rRy/YPSwIN4JqJSvvflVPGrbsFziHc62vwSzV
VIpTqtm7A8TYIzVtmAobmIa/++P9kjeV4PwPkDk62fnsrhMHjXIG+ZGgwn/whIgj
SFpRoyFwSEOOr6PwNFyKXXQaCtepBJbxFQoAsgzRH40m5q//usDIamM6JUKIWDKv
a5NY34EhGfYWLPge1RsstIkpSs+y82daTZ2ZjGtWvFjWd9LtOMGBUCx6R8qe8gqf
dpUHkgtJKN163NGUTLO/UdE3uMqZgmliT7LcK66d+RpMLzCdVbrh6PGJENZ2GAha
NmZrSlIC596+NlkGZq+2+kQJ9+bLddag1fBBMcYao1gONsKUUzJN8CyfzSasM/Po
lZGQuFFxbnrwMvTzE/hBFp+hg5FBdg8MmDziBTogqWsBtoAWIz/Dz5t6bB4sCa46
IhJGE6rxJ9DtRWZYh7OgY2Um9XhtKr3VswT6i5hW3qS7c5QtbfSdteeAV+Hy1p0L
xZ8R/qy0X2/OUOHljrIy+09YswSWJP5q7jx52ZSPEbtctMl6DB1JkHgVWrqLjhRZ
6zf0V0D0ULqGXLrO1uFm46aRiG39aIFIehHuG5tuJFuefV/BI5U40P7d95VFhiFQ
b9O78Lz1yiJwlCDjfMIpPAHFvjq3/LdkmbTCjugV5pwPlMrJaiHhgnWbG1Cebc6C
Dy0jQKuTRSjT54jVzgLX7x+SINNs0n55OZJwpEilBrHylJ0Z23vGqJ2XfMtoqg1+
QggMlKxC9/Bg2N36JgSSmIJByJMu0q9qDPUteu/uE+dxJlzCWy+JCVFdz4+yQlf/
DSIh/qpsAt45tS5Pyx7ilRKfKTCdtxcOs1SIKVqUHAInXD4xmeCdQ06ZXb/ZCin1
xyRbuKFJIBk4a5EWhhj2An1Btznjt/y5WoyHh/khco1M+gp+jK9aqKR936b3DLuy
dA/GWec9A/eIb3wQpZl3D8R+8EzoRJBksLhwZKB3hIwLRryLo3IweuZtKUC2xS06
TXlYxaLngEy3YodFu2LyEuil3zcOID+LIt3HRO0lh2jRiakmYznz3YKtS9Aqvt5I
sd7NaJMy0XzILcuKo3UMkDcnexap8wvKmgXbEvMk0JlvSNKGwysbG8J5EZ5Xej2+
nddKFUblvqhQhBuvu+E2V1h7yoCihdDo9+o+tVC4ZTIdqxIRg6pkbTUBWzti0yVE
cGbgPDKzfjoU5t0b2O2hpNb3yxpWTlzG10ydpA/oFKG5brrH6Rk0jaFBau6CP0Fl
MaHS+whfV8i0pBLNn/knIL8Ravm71X9Pb+UCdBPpDC8LQamIAU2sFOMpNvNP7rLw
r69Y/dVaZUDqCJsP9A7CkfsPDBJmdV5yRDY2Dks9+o3vWMWwXdCmWI6mFlBXbpvd
LHvZuv9Cj58KjnIr1wivVWcg/pI5WCdTF7HFRCUmjqLfPPSYoehpfVMZvjk/D3nn
LNq7hR2zEq5Pn5vjDn57jX9T2eMPDUbKjogeJO4TWgIp9rbthymzasbI+SSQqlts
9+42bioMmJIDpuou1HdkgjIsl0RsnXKDYFniaq/YAT5WljgUk2zluB5mwQ3WJ3SO
HFTwiyFHy5x8cIp+fIddrMvJwfakf4abWEmd96q0V3RQCVTmLxN7TRUx3l1bF5nO
gxvdsjId6mN9w2NnTp/j/PMacaCLpREA7wGUjl/316/ynZtaero1Wm8RXWh17PfN
6IJ1Li01o/zsAvngsJKTOaax8PrhASp8+Q//UmAwaJYaUyqViey2nUQx7+IG66d0
jeUwFPI2ZOW8mbSQw5I6ypFbMoqwOqxVvP1M1/au/UTR5C1g25qy13gmCQDjNCmV
MKiwshuj/pfnvka6Su1YMLZo+1qleacpGOaFp4gGbPAJMJsTdtkCHOsKwqVJWmZr
58UjpmNRW5fj+nEf9hg+VbQ7c5+kTlGmxc3GeljOCTVLAYsCe1tERMHUaB/LBY7U
HUeOiOG7dXnyWVW7WuBPk36EJg4qWpmr64Q61KUQ0zRRzFIvqUPHDKp/4NGaPjsM
FCiNdB0AX+dAQfLtnP0GDynYjT7W0R+eeVvv4T2qidJtCS3aaENbXAqKahAxrgPH
6ZFe3PVU075oDczioPZa/dTXsLPDpZPRhHsAk3aAFuSzencUhILWN6WY9Y1s1mAm
ZUzwPcfUl0/X5IihznZSWuktbGxWQuPgVxdxRuFM9PFehNS+kX5Zlj7yGgEF7wfm
A5rLcqosWSR6WjTCOjLt0b+Gid8liAkdZKnAKLdKowDVhLYdXq2ZkkK1aGHuVdeB
yKRhAoIEOyizepvZH4LdUXbtWcn+pen40BAwwNEzB5r5Hv7e7W1NVX7zrn9RXOwP
PPNOkhtKgEP6yJt2AlejJ5eUum7kCwjox6ma3jdxyJepbVWYwuqQxrhGF3tFxdDy
Ix0VWZ/avJwqeSOMAGbVDA/qsYoJ/SXcnQw85QbBe7nsyNaNcDoNGuv+MYtCfzNG
FYViY/8w/+ZsZ7jiFu7asz7ojW/LzYY98RrRKVyI4WYrtbr+LHXlb59jULZkVHFj
CQspRJMIwGygJdOSZPkIrZzCetB+41amRCyCwHTzQR9eVhwUm21tZKjZXX5Q6MUI
2MMElQIXXp++XADzUguPofTdh/0Wvr6qjfvOQ/bcDREf8HMH5vv4RX4UCazTv5ez
VWTYR3j6my3hovIFcXy0mDUtWJE8STsSnYW4vj3iQ27uU3475L7pxBoUo44fCvMn
RdSVz49QQek9DNhrZvDn0oiPKVmAlOBa9Ce5Q6cdjx9Fvw13sU3pE4xGcYKoKUrJ
XrFOiYKKA2/7k/1+HmLoA8LzXDIw1bksrJmhZNopruXJasn3zuNsMyXg4goVEMlp
5g6iVcMtBXIwamrHMxwSyky7zz6pDfHNuJCpskEkzsFNxTOhKW4QVrnOa6QwGtDD
DpHc5liO3AeQAVHM5TmyrNM+AKmqj8VLzWAFMmYB5hBIEjMznceKWc3ZUYbtX8Un
r8A6lGXHlfczOLyAXGt6js3qHivaJWkv7eeYq4TNsGgVwu8rTCTqjk6vA+c4UWx6
FwwCw0ryd4deZGA3E91CJy5sh4eecpxsrY4brFdjHm7ACqsvePNg77PnHLh9tIlY
VgVLw7s7n2opeXBQCugviMZVveyoJcMzZ5cB5gzTpb70nAUXC/bKIyQzu/86d0XF
gNsMAMHANZkZZ0i+Q7JHiwfa+RMksc6YuA7HnEGu+VujZcxyczrGGas5/+sMFeUk
QLQDvfcgESPKGGYOPooyMfjYlL5uiLZeY+f07tldNGaqvb5OZyxleUxuEaGnFJwJ
NlmeATR8wfgvgqKdzVVS8O4bFdTKzKqqxlKsE6Edes6yhoOVNZzJsMLa2OR42FtK
FmtuF+TE83nUtSCTF2oHrbotoCx27ox5Yx290v3MHrOd/s3LCJq37TTnG/vCUJf8
kRNx6qXHhyHhr7Tdne/yB4pxknGjkB0XZIYnu2SRxtOQT7LgxDBivItSpXm6m58P
drApLJ8M8DCoY9BolRFySDAru9JRvrkcYFV0uAB0t8916JWogNIpN1+8cOHpqp4n
N35Fxb0CDPBn9gogmuBZaURgdCcXFMqUdwCV01hPZA1SQhbMQkFoY446Bc8X0sxD
0CAaeUtni/sOCkRk0sELLM4+1Zk1e1CFgjYrnYAy94dcqXPHN3EZJFZ6VGDYRZAc
NnG2ym0/XYuJxEb8OqWdonWLX0WXmZu9DJQ1Oq1PXcTCSG/E0UVoor9tnzkaJ67H
2HV4AiII/k1zIcaDLO8nW072xJrVfLa4qmlGrp7qmsSdZ2cnD5BjMZvnt8CBfaVe
8i9AeDlx9vUleGbDcLIrGNTsenwC0arskyVGz1i4oIoV/8QuZWeov4YPgjevAUlX
SLon1huSUDnHDzrsC8jS1tP/IE54dl4roIhAsL1cB9nz281Ikwj+qyQTjGLvzpA8
Kl/IgD305ycUHpsOxgVWfj2Qqj2v2x+a7s6vCFywI3QY89uyVcVhX9mic0AoKVx0
RCNCfTlk4cb2iBCHY9H/PfOVob7ErQIjXGwP+hnGR8PN2yTfrW9yF0eZv4nKUP7f
TDCeMlUNXv4LWM/dDBhHQ8b7aVH6pEsJs/RN5HsXJsviwNltaFKKJIGAJfSkGjRH
L7vNfbHkrkt55oRKjTvvBIC5ji7nNgxpqAQSH03tEOPeEgQCAiPZe/1A2JUgUQPc
myYL71FJQY2GncnnpyaCXeY0xiXktKMzJZsOzuubDFr9YI6JCEnSbiwdz5Wg64PZ
c2eyiOyyPIG0EW+AcsBZOZJan1YR1IKBudvQVH2i653cjCoiPev2lCtqSRD894RV
AcIt9mo0zSvttTIWxF8Ey1WuFZsmd64uLigbM4MuQRKkpf98g7LpeGjr36ObHQL+
Unb0KXGY7Z7x8h8s/OeigaXVGGuq6aAXv+6Lylkro28RA0W7AY/KGyT2oIAzohnf
/fGVOA1SQyyYwejJZCtINUmLdJV/zA2QmDxb0lhyDqk5i8dQs9V6Jr8xB0LF/h4e
uC1zsJlqLozEFysX8CX5TImzTLfGIs1pIkK/+FJqXVvjW/GzNHz/4P2xkpdsaEp+
CbtTqGFCn/jvIEY1nbH9NTriei95+L9VmanDRWMMN/ysVMuYWpzmS9pXqWIhDZiy
WznlWdNObjyuxHlqgPZrYE3h9+LBX34pNdW8bQsZDTEw9CbqrPWz9Vg4O5KvjQQB
GKFnv5uPV0r80c7BlUvQ9to3ejXdVHbL5mClEShxkK1abWFKqjP1Q+Z+nAMCij3U
hkM+1eW7QdOISPtIV4qEEa9hMCtUt77MW+WjeKEdaxaEMHDv5bW6eFtdJk+TRZ71
AMdqR+smW5CfYRKisZYCdAcIyuidvghehSmh5DyXlKGstUBs/G6EH1Mz9u8LDc9C
5kN+sg9yGPV2U501hxOBcgZ1IPKN3W63Vp3bHCQxnvuTPdq+bp7mMTXe9MM93s38
hhmCZ5+QSDiUmpcTwq6/V/dv4ObHWrErqU9UiyRYELl5i2DwtejqfTet42HtWPxZ
NuwdWi9OTYyUENNbUtP9AyFTuDB+3H5eAf4lQ0lvg/PtmuLVz+yhNwA9QDWoyFig
t/n62jZHX79U47UundUpXKFQJ1GcD9wSTCR4xel4knvKdydXdXr9yT1x54BvKzCx
77rd7iyOPiPtPzw+I3L3mb4JCON7yNL1CtqZufmufRKOt14dPMT7Dtgj4YicIHgr
7reXj+BGspoSl6uAK+b3V/9aW71A5Y0vFKPEZt2MWi+I1LssqpXHP99gizDA61Tn
+U1rO4mS4Ke6EL4SaGTGT1zzSzZm3YS5CfH/8O5UqJbYQkR1WKKeABI8eXJuOO8Y
VtzJD3HUeVrbPS8roE8MAQWhPtHvhJpFtD6Dn82rXmFcPb0XO775TGNLJO2Ph/ww
qhNbSOObM6Q3qc5xq4wTDjYvPnZV2fd6m4Q2fPToZTOBJqjz6NYToejBKcJaRbnJ
KueSEZaTr3MkGSlZLxJS3WQPNc8N5EFQss3W/gq/xWwAyyIh8bm5dOj4/Q+pciTi
h21uH8orrXiqJ+KL7NxNH/SFqaoammgH7iFISw9JnLyDOMMZzVjXW/2uy8xe0ZME
Sfmqpmd1QvMVsfB4mQfEKKR7PdJUhYOdpXdf8enV0L85fRilZ77nSKCBWxP4iQX0
3naFXd0vFQRnkjApBNnbd/ua5sOz1y+bVAXBEouk9FWsNCdxVw8Pz35jDV9Kp29e
+OQVBBqJ9aTHBzseNX9DaWJF6kgzbXtZyzSMZNWcSbMgKFUdOgYBwQVA30MFGlr1
StCDg96H7tMSbGGR9fDbcV6cAe8dGKhsrOjIEtdq3OyKj7EbfD2h5OzgdyAqG7tn
Yu9Dbkmqg458+p8FFPfGVtyYClkLP1keU9xZ4xpVnWTrAfeRK7CX/oGU1eJar8TW
WFCKtVvQBW02NVWW6XspGDbhoaB/6Jv5htUMpcnoPal0i6Lf7RSuEuQll0dpqxQr
cER4IxKpKrz3pKCDn3ihLRfAYU3amJJaouJ6wM7w11+4r78o7zAL5Dsa8IfgyxO4
nOLnIaQI8RJTyT4D4uSfON+lEUutUnPcWv6TT3XPrhZqHPMBLD2vW9DRiqE9p3cz
LGkD62x4ogg7Lza/fhcVt1eT/stqRJ978RhN4sKyBfTrrUkJCcRpqxyKq5HC1XUv
LaVTqiRP1LaPBYYty7FQVfzWiqqypsJRdiJwBncid27A3pmsXt7Sf+tBnI8sJuuD
nxeqx+PdVeNlX5RPi2GPAUHgm5g6fGE4TJq4bNtzA/Sy1u4NT5gECuQBgVlM22WV
djXj3BuE4Ou7Vdrol6cl9FEYEFK2LNKBbNEc6vyATO0KnH4PbfVx1WMYo92gNrfo
FqcQR6RsfnBaJimeGvKd9o3YwVyDMViVXx6DIviBHxAJo2lB7KhrWfD3HHp/F7eL
WrDM3SeEI4KDKw8lAlJELyz0EViUYYLlUzA/kNlgSq0lRy0BpamB5xij1kkRuyXd
MV1LHhePKfdxlwSI73XGPH9o6chKPu1W7aAv7dNQigrOC3nruOdWTbJ4nz7uNQWA
1ZIFQclE5TwuWzsNZotKNTfrLQocFdSYP3X6ejGHrK1kwylE3I494usnKDBLKcBt
VvJ8xYLfEq1VDAEnff7OWG3HldOOH5S7kHqZwbg5BZ5An8ZW5gvrxTwCed4TZqUJ
HOSZdm+4a+5XwfuJdOE9UHo/XhgflmfQzMFS4y5R/+tWFhAuxFQ3sG20ldDX/fRe
7k9UjKnSdEEnsrisJLvFfCs3TRU1XrG3fHZUUCsU9xNuQcfGNMl/VECdLGNjmyEY
hwcsruxjasQBEhWp/OkmsPDdw5CJdmGGi1foWfngfuyEw1KDPf6/t5Uq3eUcwT1A
Mq3wL73MjWznp4Q06czAqlMVN0tsGuRzhe0TELIEUrWyskBU0Xhsjgzvw9bvlpnp
YbEMhsTox6IZDOy7nvuls2cKXQB8gJLP5+MzRWtSchFGrZOqtCzCvAax8RA5toKt
LILCI3fBpsDKYw8aTxhz9t5p6I2/POXr0svalvX8DGojkB96R5OoQtRDMls/eqjU
QsX8qGx3RIm9II1mRm3k1tZM5e8uN91cD9afrjKTXihkPouBth72Qc3DY3g9URdN
EcrdWZBamGMPID3m3B2pa5lSiM5yuXGQoposD8IvD6wUCSv74Ofde8CBKdg9NVUj
kjR0+OmETA8AUWz3lu99AJ8fMG+1scoJF1SVfS7pnPpYTkPw4d2euZeRG6KDfEYT
R4/9xPqzvM2qq705yalp0w/Ux/ZSoPslaZn59dEtpHcnpetUSJEOClMcEV5POuBN
D+arpnwyX405Mzn/vebbNuEMISudVa2+YnZQp+1JatmDhwVoma10mBt7Pjo4YdTP
WqHM69qtkYCk2ApES/8QJRIPKLVFNFepDWGBtY4wmEAIU8RiGS07nVxolySA99gZ
J+nx+N2QqDqu3On4okruszs4wG7GXBQEc0RhQcz2fZM+T8WOHovJyR0A6TdPBIFW
MGs5dIlkuBcWKVTWpvB63KcDZ4QKnriBF/6JsZMCCcxqMolz+fJG/LUuST4bKlP+
1yjxYsAZJYKn/gQiJ8YxtpvA2VxANip84FV8e+pMSIB43Rh8aF+R8FKnBu4Ps+Mf
e3F3z3RfDih7i9nwGJEusCMQWo18cNuGNr5ydDKIrbpdoTL9Bt2CBMwhN7jKBoCH
l6QObzABMwowoDi2ZIg+74xUmmeUia4+BXO8AS6FMJUAlnNNt2gmeDHgXPcUMNnP
ib+zh+bj4pKJBFaykBdedYuygvw1IjTzMfM9CA+e+jaFcq0tUcwFv0UvtX1NoY3c
NfgPopW2N8LuLFbq9tooaAf+VnyTnrUngQjckAago50f9iNWf8u7A+SSHkn58zqq
WRfLrvs5zuHyHF2TGKTnuPih33Q+57rUee8hV/sqxXSy/xG2EHw+nqF/9K0Y0Cmg
i9OnalAsTHTqzVRpwZNZnPfT+rcTRuwqe/15s8sj/y6fIOdbHT+itbb42f2aDH6e
9iSX+Ed2gaP9E1sIgvHbNdqWec/oCZn9J/1w6NDSm+sFqrzgAYa1NPag+ifaY39t
A9dw9ZzaIaalEow3aoUmdjEFW1Y0swBUbtIgG9e23hdEOgDx0nkquLQRfxce40Qg
XPLm2f1S+eupiXlshmZjQc6FYbZ4QJk9JHqBzXWHyW9UsOWI+pEstpPhx5kjuy6O
q//vUgmtrdReITc1TPc550OWQqsM8HrySIa9HrTVFbOC/A6Jftc/yPtGBvMn/spk
gETYXNBGF2YPWOr6qzHEcL936OwKu6MvtrN02uFnYfaWlcak1d473ozoo1TRqsRE
dfFBwI/Ni0yjwQI2NB1SmnLDiuT4Tewr8+stiAQXtLrbH173SSSz2CWf48ACIKGW
WY/E5KGKh6FszGqsA+jD7Js3FR2uQc2YnaBDnE+wubY7oxTlpCLvsYFBUZ6cSkOJ
Xyz8FfyioPAoPWtWiDxAIvnW/fu1DMP91jKkxSDj2w1R7jVU5UHF4W1rPkej2V4K
73/3xh8dz8aRMQmK8mqFRhBuI35QQnRWIEqDvL2l8CemXo/DzFAOSUmKo373mBCN
7RT0oA48osO8kwfHofU38LY/y7NSdmDvNiTvvnPvTCNZLFaCXhuPXF6SIWib11qs
E55Fq4bvueh6Nvod+eFaOPYkvnPy9gLsLricND8fZ1HUBr7Pk0R31nJKk0Q3Jk9q
jwLDZbnUDt/hVDhbZkT46Qp674TTxJx14LwvWaYnUNxX40VT9dzkWfsCwcoSTmvh
baRn4BXOCEdG2i65Alb67jIVx4KAyE0GFk9TdYDJeZ4c9UOT8VjLwVozZcmQkBbn
16vPliJhUX8BY4uSFawZFYdqX4svP4b1sdg2miltTENxjUd+DTnk9tz1DKKRExIQ
Z/kp+7HBXNn/O78vxbW+z1AQXoGRU87F5kFu9fhiGfLf2stURrAk2HuoHx0uPpos
qC4PiLYjIom/B293ka75yHGBqbcAV2s9fm/JqFZVCw8EAk8Cs3G3YjUIlHl9B16M
0ocjNnbEMmpPpf+0RMx168CiL66QGWDGwhtgEjp89a0+0s7bLJwJgAsaksUBzBmx
EWEDlCyP+4rs93xms+K7Qazc24CELlTJaP3NK6fZ2lntSoe3Suuh3v4xeDfvPZV8
ZQWDtc840zzbu4AechaZ/kJpRlgTTqkpCnK9UQpKRZ6jzMD2QQjNBZYbtLXw9nLF
BHNRKr8SLDXvDpk76DHNXDPAcxrd5SsKA63umuuIZ6Vp+dkNmvry2odk9T/FHE5A
36djTYWoSIIzMjY1Zt9mWfkYx+AeTvmnnqarb9KvT2RjPp87DdFgp9lSILX7ImHj
AndkoQ3A/OousZEnSlGDpxGHDnaXhquo4VlPll/2RuUa7O8Y3LZ/fQny0t9XDB8V
O6JH9lj5S/RiQ6ZyNTnasAn2tmHu6+44+AiCx5YjAEf+35r3MUOkxJCuKYnhcqxl
z7K2I2UUevbmQt3YsNocJfiVOgQqSRpsd8FDTq8pvy9dIh7n0hFhLwUc8moDvVeQ
BKNtwhgm/m3Ss0/5H7ZpLUKUSM1RXHsNlBaZ+oL7Bea+uNc+nqrbyt1zldAUVCYZ
ZHx9R/WFIrrTWFC6BHi+U5IY6WZLKlCNHhfKdLGhe1Op5+RCtgCBzc1rJkHJbzUS
bp5VUNm8mHeTW2RD3C476Ac9bgj5MRcckaQdp2xP6LKCVet/GSlqfGWdnYpXZRke
6tysyHOgw3P6Xj3vhSaaGkbQH1zO4tTg32zeuWS89cZHVCUq2eiOsE5vjEaWYIdF
2b6/Rf+8ClrgVw4MX9CxbBYUob9Nc6idtMrm4WCnTy1hvSuda7KjdtT5+Wb5e3vT
PElvIRYcZczxNbXJ8MqRna95nDVYWrKW9UdyCs1W09j6iza65TosS47MMayFu+xa
dD1ATkPqHl0rocqNRSalWEIn5ZFgA9qbtgjQhszF0XJz6nOig1x+6agx5Yd+0f3Y
+e3b2ty0Tyqh8XZiA+91KyyUJepoJ6rx0tkNeY7kB706dKF0nQdLqEz4a/X+CEHM
lCPyMMhft/rMHtdVWp0GMFa3E3525kst4o8dVLZw7CpS4sS6DsvQb+quGfrVL8Ot
XtCc1FpYjTwA1zD39EfAkeUppAkP9GPd1VWc8qBIIM97IwVEtkFI40nJJcPGkhhe
g2xYhBS+YAowaF/YPDjRgXSOwE+YZDgiLXPlMOxFmJVbfZ/Che/1al91rOiyuw2O
fRgarukpABqqYncvTqpp+t4+MZCZImd9FSSoY1Z5yWVU8tKqCzztfPkjFaby++K1
p8Ckdo0Udp5uSy2cOJBZ0dXoZiZgwSIUyCtpd9ZCyHDCiFaX4gUQkJI5hA+cQzxx
ILF04q0kREwRmeyGoka8ClAtzq2D7PsrePt2GlLWqXaUwb5iXKFSuysueA6vw2dj
Fkm1pIEU0F0mXbwnmYhM5nNKShNJHLQN741LjWWM4NplzXOS8LxNVv4sHYQq4KA6
Kak3Iyb/CWPumzCmvp351VRI0pyH30C8bbZXEhYY+E6zmuYELR/orvLNzQnEHEUj
gwnPwiEjYEyi82lqZk05QcB28VVJPTZbDUhIo6UIKDJJZE+ItU3p50z8L7X5/qjU
pTKVHN81W51LdNXtuE6/vYSoOFgPXqbqTBhWJhsMlIRxVvWHqan+mXq3MkmdwAPa
Lp73/56q9YOhlx93Nl2mDpdajeGVe+MxIZxAu/6uzA14PJNW5A7dyqJa0Q5sVSyI
PLA93IfDXtBh3mSih2ojdSl8z7jhPVdTZ0AVDhLjrfaOirYKQwAqFB7n5I8g/HRL
FqAotMHCxGQfsqGET96JWrObPqTApyXb6vKRbFnzL4SDN9oL7aDSepzvdiJ5/ozo
STS7PsgBvfVl3KEF4p4mtP+pXHcq+7VovTFM1p7mKTrKu9Lg0vgNIYE8hXjrsvk1
TKy33E1BFgcGljzoIb9pzL2CRUvWjN9zecWWS6BfPL84IYjtsaBFJ1hQroltBC+W
78pcgGv5MG0evCwiy2VteBoMHx63jbq2NwAqPCM6CP8W0FCHOH3uqnNptvxbe8DQ
0jyR/uJLPqZBVYJDe2MWUKwS7AxyHYVTkr6pUTnzlbo/tm31Gss3Rkdix9i/7+Je
pNXfedRNaley3k+c3DxthmqOPQUZryzp7BS9GNTsVQ3TKnQ0XYsP3q7MXNmtuGb5
5Ikt61vSOfVw0+/XB5TJbRhELgLrWZID9+dezoyG3QYrsqyQ9z+qaosUJtYtNBv+
UgXuOiGVr8k+V3av2qky0muSibcsCkbCI7lNBZD3cW8tixiPgtAetTiSUkzRsdUz
7c97oMLuLYckmtu63GaIlmj89L3+FwOVuiu+pLrzVwRLpLaWByQqlRZ81pI99M+P
0T78V77GpD5xo7FdrjciXhXHxMlXVnDmvMwHxVkmZ2EMVkhxuTFZtki9n0WtLKKw
Z1PDz692YdY7E5vT/sqTLu1eoUrEBv5SILT4NfA1VEAvqr5+BTvAlK2ZaeEn741H
vgXT3rz0apcRB/dOs66s+7eRNFMyoIemNGy9jr7k1mPBMfJr19lkrzIHzSh+R4qd
MV0KfPHVGOH3k8tyj780R7SAdHYs2SCwu30YdF81+j3gWQGO1oIWgkRHfyaIGwJT
2sU6dNof0kXOWxyVA60hGCvMCAELX2DtkssFcAaCiMNP7Yw1euXJDK5iP/wXk0zp
pdEiGwp6VCHs3vXIm8msBpCVBbynC/Zm0Egl7XpXTQvnsPOAoaYb42377cWXSgPJ
KEvMwNGcFAM8zlHTR5S6Y1WzNujhVkBMpRYipTGQDOvtgWmVV++BUiv262SZUagh
Z1ZZwt7HALLZv2/8LksTlbpkKIgAKPVK+9FzTTWX2J2ZxI9h3IpQlB5Quz+M28BV
F4/L/+Hc2Zm9mG3jhz+80TLAuqdLGnyZICk2HjAYLSvJlPN1H2cimNHLecbMRt2k
LFS/bV39sinMEtXHFWjtvLRSnITfwMsy6tQgeypy8GiOxAHaTMVH93Qixaxz8akW
k2YSivFq1oWX/fv72EDG7j2uxIc5mQNfifCmIi5ALE8RMwYkUyXPRQiIykIcsGH3
cEvZSw/FMOW7vLR++lxjo5ZhUcUg6Fv7wViCuDqjdbbM8JVa2bRwyKLWhiFAfFc0
KTw+jLhEP0JRRV7TI6YSl4gRBtyNd2PGUTgjV2KE31DHOgGbJ0c9/VSXaNd29lV6
qnn8PzUOi8IDkyTjBvGJaNTn7UrUDdw8gaYOWj5mK9rdYARekzblPYRu6g2cLLs+
g4nZnBnanLSd2UJfA2pr0/HksEvPZ/g75pJiTYLIKnW80U7kov6Ld5H5f6oPkKxD
lVVDXY27gLIC+N8cJwNmBJKXD9gdzP5QNzY6d/X0F5RQQJuHqQRcYmxmh8z5cGFh
ZaOXK0IONQYMlrRNHUTrySpsXyOGGOOZg8FabOxpURlROhHPqGZPbayaGlM2WT1+
IFgCVNjxiSJ7U6yCIUoCTG4/AzGXqUYjM2PIHEHYFFo0UV2qkNL//MhAr4kdyLht
pyupm5LcL0t1FkSx1CyP9FHRFGR4N+/r9QZNoOXBxtAeF7qUjHz+Ldcshy85U6Cu
x20CaXGv+EAyobb8jnxouMPIzDscx/XpiLh4MnIEz+vhAQEdun7xs4nVpYVk5Hsc
9LcB2y068SQhVX4fOREwtESoPtWjlMnjFvXZd8Qzhbetpqj2vIpq6l1v9+p8aDGY
qwGcXSBQRqfVrjvMZ7qc3biMvadnGsk7GFUtqwNB0NoTdj2ylRZC8yNcnzRUW8Fd
ztq7uu4UEAFAPNeahVezxo50CzEglyXwXHD+jacGonhXJ5hvUtnAX+Q4Z2/qyC0d
PTRv3EHmvaz3OEAmTqvxY1yBOukpFWsz7sBNiMwdGX9kMPfU0W1mX2FIWGH9LzuS
5Sx1wBOHVkym9KKCuZxcDW1qnFQgvLBHovP0diPtN8DIKFUlmctIxtK9ZuerHwYv
Zdn4DwrFwhHVPUtTQaIZCCanIBO5MpQ29uli98kO0JBlHotXg0j+3Rid9u3oyvFI
khnfV82xcZh7AEkhOxTfVeMzw7LUIuHYXgJh8+I8NBYU0hWLG/6R7rNnFhYI+nfE
M7vazy1rDZRFyUU7q7Ptbcbx8uoUjKHdGbflsZoc3YlvhHYZU8yQoOgEljNsdM1H
3J4hYCf1DQfILcmp3Nf01vl1BiNhS2sEoJyGFPVXu5B2LCHpb5rAOQ9nzU6C70a9
lJ1yf5cK6uvQnzSBTGhvm60VPh6/qZdztqGhro9DQXL/oKPIznc1UrB8Nv8HfrSD
elYsOaxonwT/q0aBo2ujm3S6mCn3d5dM2sQjFUW1i99oJDw4SHKpplcX+wjwWzO5
MDE49Te3DvzkKubH66xUROipJ6I8+vxCfhKKm5VZBOEnxcc/jyIRMme0xAmDFzt8
jIZUT2w8fw8azFaJvskJM5f8Y2e1ObC5vOq/LpyAzREIIQ6hlPvgGNn0twx8uh1J
BhaPOm7ixbnEmPqgJ0fIi6Tl46KYUD1+OCVDcS/WfGGrtbzVYVokCFMn/z1tdwH2
FCaYHjfXtrrXigxhrYAr6g2O+7RV6271xwkWXHQg3i5SQZuh/ci+NF4V9AhPG9dg
d5wzlKZP1Wvef6Cpb0rgLt4+7UUJGSQhC/Ydejr8uOt7HOwm4QNWRSZcgdXgNkr5
/wcaa4B5ag7Cp4FcA9uI7psvrGzvcpQ1wlee/OMgByKOPq22FJyHsvEmR4HNlm7H
Rsx21dGjOVPlCxuigAQ8I/z3/xUpwQZAPFa5JsBAffZmZzICxTJuHxwYxxIunBDv
4OS/b+wlsoLfwWEoEVPD9XIaK76PGcFb546MlPg6DQzgf6NyboMnB0ClmP778LOp
b08mn306VWKcIPDlEWtNN01WNRtu4ylFZU9hOyXGyYdDeiLHnXFp1NYx0v7DxyAW
pi4XjybO3O02jSl6MPm4iWxl0lvr/Pz72MAiXRLBHe6YLd2kZ6WWhYkmugcbvV1l
bkJSLuS4Gyuaqg8j8UgSTTNyIb6hl156fMZ+j440fP/PXpGQ2GXTRaiZ/rFG3E5E
x6Gnu+dtk6Ob49UsOA+LhWx5yKHt7rK7lQk72Itn8vWbZ53CAjb5/CPqAvKiRL3p
VctfQuZiPJgrxB6MhAqk3rMhPjsyMGuEysIP4fE5xrcenOJdJ4dvtRb8IbrciAJ5
nFuZ2djneqLFuIAR6RybZgv3M6rEuj5o73fj0A033rozFYPUzCHp318n9+N9rpWn
LKEHDenIUlM7pktsqjwWTap2gci1LyhF1tSHeiQGBjWu6xtG20PQ5YW7e+tioFyX
5Up+jeJb6v/a6k11xgtR5HM990hWLhPrAIxBc/dlW3baLKDwadACet+EZIdciVHF
kpJkjVbRpbm0xHE/p4WZ0ftzF9ByY19/vaKtYGdzvbsTbeKKP+sD8d7CyWzpc15H
iufs/n3uMzKZSIUV57sWaym/9yuvgnm2vdanh6eeTIcbz/3kZhfn7xX1oQOuLZu2
uYu5Ab4LvxUgYPJ/DIcUrJg2HAL1pwGuihftW1et7sstkaouhhfL+e0G1gLOlp8X
mKTvk8KmYtEQ4pm0b2QvcuC5ze0eLU/H3y3d4pAEDu259OjAnUtOAZEoLlPjLiuL
88/LGp7cKIO4zaMmf0bFywRg1PA18beZrWzqAvTS7E8y4Xo4pLAq9Coc/cmXCoQ7
kcUhQ7tpoE6dFMWv3IHhIe2pDf5dHCYh2114E+BW0n1i0owxozWfuvH4o32Dxxgt
03S4J1WRwJapR1gQhrfO6rXw/DLANPIPTGjsvxnAXEmI8aDkGJ+G7L0SExjwSWyc
dNhYMxqlkXkqE2W3qlHvIm0kRl7HeDaBNGSDl2WvpNlEPQhrk71SGjIVG60ptNd4
HLwsOWsDYEHGAMIKCeG8OVBAMaz+x3U3UE531F+RMm26C1n6PVP39VPdRSrbujQf
iA/UTG6gQzQooKPZ266mqDUUBPPcN2cMgmUu/xXQimk9E2kyuxLEn8OJuTQDUTVS
G3JYDVIaqlXvwhnw2ssriFfJByzujM//D6vqgY1a5NJZwER5I6r+xH4HGgYyHfEX
AUXgAQQ53Acvn3FZ2OuSgOOz9uWlU/C5sfcnoPJ/f8WMAVOdlPUV6IC0Rc/TMmnM
OkPsebndyNgBOQLrttUnwxVhQP8BfOBGZ03oeL6/NTfsEMGPPX5s6cI0waK/vgak
lB/L60lhayY1HKDpK/YCe9rZRi2zqRFvLpwYSVBOis4SToRK18sQx8MxNnSXYx1J
ya4DlwzRlEbESoS7T1gS9RYy+Dhg5TANRKJvh+FXybxKV2zN/rWpl2QDFw+Z5LT5
5BLF/mp2dTfTnxLF+ab+kuHdu1J4pQg5YNmKsNfcTNlWg1yQwYm/ELNJmCvMov1Q
QRcRXMva8Wh2rQ0p2fXFreYf+8LzjMo5AgaRTC9ehb83T7ioijWMBV+jwcyVtLzY
3eg/ngvIdE4O2Vfv41cjFKTJQh3E8EjGBibK/68frefzv/89b8tAoe1+ugwSGipk
nK1r7js9p9XlxULhqp4cRiLRv/gc+Cmxs8PNyrgc/8E2pSv62XJn8Vn2YSR8MeCg
Ps28PYykomuDIRUPZ4tFSp+ta5IRQtXxX3JfOFssBnRkkt8dFZQqxq+tL86yGIKV
b/zUD90wjQhVzlPt+QmPSx5+hQhwoFgHgCmuIUvBu/1ZQJ8GeemW6eDsKmVLrX7U
LB/T4CRAllYHwC7gam/CMoe/QiU83bUImjxykld09ibbrgqxssAB6vwUMsLqDQTe
N7iLbox3OhdPOMHj/VynVugtla8TUPsyKy+6sHuZijOUSENAgUCVT+Q3j8jYrSFW
Y1AIf8KiIeI9HyEClzDFOESsz4ztwPiwo0vZL5ueZ7PeKc3HzU7IzCbIGx+8M2s7
9It+0vT3HhbJhFOVrC8UYLblqha7BAb4mUR0qu+An2xTaAMRIX9m9k4YP1Dm4WWZ
GRKao3MMBbeeKT/+n8pOnnAPdknR90vx6cPqRmD9UwmXWVYUUl0YI/0vhsPB5TG3
sYrpgaGi5WG/v2QDd4xFTV7ANRPP/QZURGaqaRai6A1GVwdxUq+GM7Bs4fEFzG5v
QGiyekI4Wk7fPcVSSImNa4PBAmEGjJm2gwXC1K0DVtoNheC6+BzqYMLK1MuMSqou
G5+dz0yc0fN63rZIjIib5xFU3YSWFztXVmiyg78yTiKGo8QZhIGOqwdgm5mQA+q9
/XjFYLiXkabWJ6vAU9PZ/OcAa8PtRsLtCEEs8f6JnsJECpbwuMqAEf8UoXFKe8zW
r+wfip+ScVZEKC/zgwWBWRbDa3ggTZP9Lotp+8tfYqVilcys+bdwyMFWJx0ruDQI
cVG6Kq2k6O/gsBVf9wzq69sEYhT74Q8AIp7e/KiewT5TPupN4X08RVxIUh+MgVlc
gadH/BvlBZXvBpeBSFRTsUsNe3uWZGza2sE6ejxuZyb07gRaUwW12ygKMTCUMMYl
eis0CSCF2Z3GL4V3HeqEGZKgcjz+571DdBbXO6epUa/cIB4IwfeDFZsJzwj32xPn
MIZxAJMGMps93aK9HYAUN9FSb2hgDi07VTlllPCSRYCLlrVYt30Gr7bO92cE4usD
RgWJB8QK0Cr/SH73HlBDY5sY9dPiryK1qk4PgWuTuVn//o2TpmLwobFRbR3umdBU
8pRAVdkTLkHfGcsRYdx+g87xT1nqZyRcKRobcKx9BsGkfmiziva+EII1npKZOKCv
L77DiU5zqmzDdoKTRnW6ROr/G+PSgmiaTvg6zR3BZHh9+yx+uyMuWHLwzi9Ne/9C
6MR5fZJapGpzedRqggr262sj7w/FYnVV2xiI8Hqh6rJFIy9MIPonIvkIGojvu+wC
iQ3kXGxDrF+aZoM4CjQTwtakwxyLcYrMiewTh/W0kL86V430kFt8qW8UQ7oFO7mN
kYAlu2WUSV8NRmWzdh0OVybIOIkLZ6EaBfJhj/SlRoebCUZ/iXD8j1q/znvPu5WB
LhRBoghR62HNUzRePjHLbXJKTpBaLHOJROPUj+dNHmQsV7/nDUWX6e4pXIp9dg9R
CE0/claOet20M3vhdceyG4n3kp95W7M56NvCNru2Z+WCCkIum4Ao9p4ys3zkOhF8
RPbKlucIz2ueS+Mx13j1QaanrB2KoBUe0GlvIBjeJeIytE7/2eiVAMGdbltZ5nxa
fZAQwJqBQ1VjmBc9zx/ZBE8u6Hc89a9e5eXNByPwUfYtIz5st0ce4vwfDBy/aReE
DjV8dHvJVWJa+A+gtwQCHz9OoQVaqFZwI5J+EAnS3s5Jp+xtgeeAUm1ShXZWJRh6
x2Xq6+9HLgwNOrr0i+aelyxsJ42i8CD4X2Ll3s4ReHRw9CYoliL19mbP5MFxBxQS
26BYizApitJQoizkwL+2oeG3z3a87f8FoWsGm1e1o7vd+23UDiEVYBSzkwSPijW6
AHayCipZRt9jXPrw1kAkE2Wu8BJIrIc1hMGYTcfCPNfha1eJm/M9IxQaQXHXoRsO
SYB/LPhD8Qf5YHyoEaKjhfUAu26hUs0CXzkVgZwiHLzxx59iwWsOrr6YbcIeUxU+
3e9QkTsT3MaRnSVTCKjdCByxN/2+jOGFbo+PF5jtDo58P8Klfxg8fYFSb2tiHZBd
JHa8zEOirfJDfpiTLgHNauO72tMdN7AHisjWWoHTtXb8DItqXs9tx/f3mO3X5AQi
RipPjgdeQTQ1JRcZOU3J/jj4HXxrak3hRqjftTioz2LjLJcmCaEQ2AJRiyjS/drR
X19Krr7BGXz/EROx+/RYij47zryDJ2qZuKBkJyfmZ8fZ9+FCzR1AlT6nnMvOp8AC
qmy5A5Yw6ihBN3egIuPPJIcsTAg9mzyGJhbd4HAeWjNjtRWhJRXFW1ptLDnkWXYK
glSHZOwfYbHINL34swhCf6QV1Vl5ZHfp6lk5rcMEGdTWN4sWeuTMSMlCeq0GzR9n
G1dOHsWD6lPP+1uo6D2HAWAtBCKMBodQHJBQKAIekxNd6WGv3YHdFDYdEgHSZN7Z
JVVvxn+AWT/JFxx0CufafUKH6OuQkHjfTM8HsE1sLGyvqxNCybq+H9B/s3ltLHuF
Ds3gpaKkjHjKkiZTmLt6bVv7rqkCaXecVzx7kP6uVPRwljqWi94h1kSRLtCq1uQz
IKHHqbZEXd8TbI8tfoUOz/DT406VoKtyTOIWQKZm4F0D7R8sY79vfX0x2R30TTdA
YlUyczeo1KH9Vzb9+2bTfMIsiRIbier3pvJj/oC2LuPxGC7K0NQj4M4Qnw++FQe/
0En2iA+pAHmNPyq7ZAd4iOtSqnAGqlt5155tP+/ddvJjcPqcOr+kaW3psdW+eKe8
PMUIgSSipRWw4xUn+G6Wj2vSjPSxcLKxy8Q3E6wjfwmNshmsEsx8byczqhk9nZ8o
CBtjn5+l6dChUSWzdNlp9ZlDv/MCEbp5oUnSmHZ1MVcfqLADUohwgNzmzUDWN07k
4XFyNUYIZabEglkvAGlUpXKxh0w53dZMYjCATNnoLLjOKIEO2UWSsJNVW1YVl55Z
3+E0rhqRuN0/rKQD1mUeDhgcJ76PfRxMYd0y8HfF+JlJu006FFHVffXpHxTkkAaP
ANHorfNHmfZgiads461PhlJ8niH9FqsgmsMOnT9kuznW+LaElqqY195fQgWX6CZT
Fnn3bemYS7hP9vkQOUtlExlF7Gme/Qe7TFN0ZN1Uk65wjH/WGmvZ2EICLuWfMtNI
t81PxJW3yoKf2m1o6ZRuETLVLU6xPHMOTEGY16/cOoTNFsxuwIm9n+KJ+6VmyNKl
jcOLBrvR4xCsRrQMmt7YJVdmkB4jeEDyVt+B7Hrx3v5o70+M294hCqKE4UlWnjBq
0kd+KCKzM1JBtfOzyBv88eS/nhYdXgWcMeRIt6W6BszVYfnz76vhNCHrXlazOY3h
3sHxu5a7EBmix+XinAevf0TLRawz8WsTvwqYCQ2HMVrmP5pnMdQ0lkjYGK0A7txs
wfpwLIcSVEX217S0r1tA0MKIxgCf1E5o0h5cyxQo/2Q/sJ8KrAvHdk46kMloGk0X
eAZMMDnsUtQkYOpCggmWFPb3YdCBfL+Uo/rppxuCJqtVLiF8yz3bbLK67eYopy1Z
vTqZ2A585sjzav5vyS19D13iqxWgbh+fSQoevI9lbrTd/H7znphpvrXONcCL3oaV
czIO1pN+M3zip/TzH6JFpRq3E310o7uukUDQlh/M/1V8PfMgQR/AjMpXu7XWHitJ
0glEZiuQm+ojImrHpmJeiKkfs3wJkelxISTTCm/URP5qXvcpD44Ykj+EOxB57WcQ
vzXwfOCLac0HFtivZgbQ7XU6hfLilDVZaRAgUuFyGGsFe41lCMMMVppqdGNgJAGe
kyW8Ar6yEt+YwY79kusj8lDyXeOmoPdxFXAxG0Yl1pR/cSI1qEFV8VSRLXmP8KKR
UIpwJExPtrIRZq3Jyh9I7hfI5EWfNDzEdHqRf2vz2pVysgwR0IXtmG3B4RZmKOzS
GoC4YHvF5TQxfmEXcmo6DqZmz7KMPeN3hL3gY9Ca1CSTezM010DO6P0i+YZK8bNn
zvkhlrTbe6qbNn1dYgNaBjT0bU3qx4PsssKgM4HFzsTpw7STLYMw7m0IyfyF+Siw
qzbVG8tmYQFqJ0KUAy9PIxbTq4x5W1rp+H5hhSgRJohDDJlJAPFEwjY4+PDPaoNB
7+N4pN9ujhbIZR1bbCPsVtKJjfcVQAIU4rPVgyf2vm4oLoF0tI+6Hu5zodaApEAR
det23k46ZJ+FTtNVcEVUKLTCxUNwJO65EuaKpyjvjfN/DkEzUj8Lnm5ccBvNxkyC
cV4HKlisVOL0W7NsrzAlKRrYcsqzBeCJpIGcl5eE+cai91uBtHqLGozP5DJa52dk
zm8D+UpEqH1b579ISooDBHER7hSnrkUrPX4vSjuSG8PVjhR6OPpGm9K/GeA048Hk
7Xf1EuKJkavnL4ttfw0wdrPyzgH5P64fyBhukucoai355ATDeM3bgBU05+/DWTUx
wWhvWeVLZ0DLqH7avmR5K+ji2eZodTzbXGadpcNnk8dxYj9S0hbATfBfRFv9xUld
jG06Wm+X76WjMmHqD6viZzP6+iDHF9GExSS4a34ItpvPIOc+srChfKCbewEaxN+0
CwA7i8K+jt8zYSZGhN8mFdC1wxWSWCcWZiNmDC7AJ+ObaL6iJ+e/3Dm++4YoPjEb
fmcZdHu09EnXV72gWuo1P6Ncypf2IbNCPtO2LzJ5u2/yfQPwaaZfi0ViMu1oEYWO
yyYJiWJ6LE6CFg+YCzwXVitu6KXHwVH9FscEwZ+hI+1VDZ4vBBLoRDT9UKbvJRtr
CUgKRLZRL99VgafImemABB99GTo4d2AqInSRUWRnGeYNEtTo37D0EGzRWOCdOUHt
kGkYbKMDrrfZxJGCknZC52ogVsEwQM4ptOpSEowBvzypj3YfahhroiB+yu4FLA86
ywk5vSmkjhmgtBmXgH/AIkEqc2PUYVoKi1x+1qAUb7p+zIISLHfPvuf9/FvkE7nY
gmIdDBCcjp+akXbLzN0tGElngb5vIqJ43xca1iwVJcczN3pFBQ6wQz3N+yfK6oNN
l8YYhoLyRYG71bblO3MxVPpL1aow6KzNWJGzZKNHIS0K8nE7Q6chqMbh0iVQeNHz
f0ZXVdAj3cDRXF+BjfAkNAC01KuuNLohFAkir5vc9xla0RkqUOuvVeLjfErz9tdE
F01aW90Ei8YFF1yhCxVLbcNJb+874H8gLgod1bYEb5Y1i/Mx7C2NtLs679lx4LQm
E2RRBBhYYiaRuUv/sOJxDUH1PicKhrturl6hOjFvIGWfFqiXnXErPbyCMcsg9+5R
TkQ+DS68zxHxMl0kckFbZwTKitQQIf4ChzYSGIWyf/BuFXsT/u341GKjSFtrQHY4
URrtKbE3XJplZIXI/dhg51n0d1k9xLdVjFZyzwJec55FLEJq8yq9arr2t4+WZYv4
7DXN8A3ZtugDuNNkhOx2lSmCh8n8DkU1rg6sW440W/Ulvxa/orvVT+l13TxIcom/
CqHYRHQwGrkoRpBOR62tUrXMIiOdtaS+t2ljabZVsjTM4yWF9qbWGS9r1axTxJdy
SPBmHYDgdM0Oy9W2zuztz3UUyeyt6Ywh9jvGofP6CzyMB362ZCkxBnsGIB2kjijv
jLZPuPPUwc7USGWOfWpzXENpb0Y7iU3MZtrbXyT2Kf5lKwEKvGRkwx17dJCiL7bQ
64Kinov0VfXsJ5xT4bdYUBRfcqBTBE66SqozKmiSoyNV2YxVvQ5wshETpf8ca+27
MnjSnqDOgxrHxFWb8cHFksqqfjhM9QIXAnxVYRu6FtOSeWoRB67OJUtdIvtipL0a
OqUGcpvCFp2IkECZOJqN+FYJXfATH8mzbqqXA7MqqIx0PG0ZuGy47ddzpcXR80wt
+6YVyzaxmwQZfzsTSWZVslSIM9cmsDW8Owxzrt9eUatU8HK7F6rox0pzFuXyrzjr
RhCYNIWxzoyXWxInI5plYdj51yVgUraJ/vrDgLm/ZlftDrivGfu/iZ7BZAiXFB5O
2wm7gV9Lz4d1GMl/QOQdoqWF/sbMPRueeypy8s6EZhE4CNsgoETpWFUgeWtmEiEk
dj3KvKLDpB7D7rL2oySexSZIcVhZ4jZPG3HHgZ8ko2p8xnc937DswTKCaI04iVJx
l3V3E9jWGKuMQD2DfmN+ruDOD6+h0NHiDVKA+YdWD02WAFByqnWle79atSwzl3D8
nOel1ZuToA9gS/IoWOFPhBxJfxLUStjmCAc3dOvssKcOZoFEyT8R+58Yn6StBHZ2
oxPJLqThL9fuXi7FQPea55XkmiYPgCBy+jKRg5Yg4uXT8yT/ACKulKu4p+j8E/ru
9NX8Jf13gX1FFZXeAv101ag5zygBkNmuGyUDrtl5uRrN52PnPfylKAeFypceLJav
aKFzHLX//m2asaubhEp7+qQaGg1bfogELsY+gIdTrHudHb7DmhWLqN2JElrRl9Y4
k+2TLjgGE14ezYlTZOZIp0unlhyTc6gbvpil5S6joJMTWACO9g7IXck1PhthgYry
ELqtub0W+hTZRetgjDzIJA8f1N7LuWZoRkiqbzYT0Qdb5UsSZeoGFPCr3ZN7CPS9
DDqnmCOajRQIkMXRnGDxE4VxO5rtMMCPh6ouRIa//jYqBqkX0hm3Bt9CAGsERC7h
1n5v2Ii+nyFnWo88pviCag2dXRe6lHlCB0RgCmDwzeIN5zM4C5gUwKdUiyDELBpT
8OYPBQY7qRvBy5emxjhYc1DOHkAnoQr0iabRQhZjpbBSK3+hQITC1KehHA7R9/TU
DmI4LluxAac7IYHhVmeVZ2UMhOfYm/KKD4TlPHzKKyALrO7Aakm1IkWZnHBe3RxP
2JrMNJ1eOO5olwplw6d84YYyubCTR3TtzgiE4ktZofjNYRHzAFpDkz71fEGnKj8l
BSVUBpA9/ksXh7rE9Loym5m+H6fblHSS00VOCXQGbqhzy03RuUqlrHumwDXaXpzW
QeXvy0sOxkp9Utz+ut7nbpk98B0aRoCtjsHF09xe2hTEdqYFe+kzrvkl1giHYoPn
RZZ4ABt2QTxD5xBTQsvzHP85Tf0aojbBbkFQ+xiAS7dESXYM74iIxm/omzv7iLK1
fJ7NhbdExpSma3L6++hNgUJm0i8kZ9JXelCH8XoiVZ6mA8+1+zSG9kNDGn+yiSF5
vpYjtbel+93m1iwfB2SR9WvCNDmfs0T/rfgH9oF2dEUE4NcCidG2vjPVFPLobjDo
N6LPit3EbeJOSNOs6HQqMNmfbxMGhVPJzX6owMjmWHpwyihSr4vODMGBhMrSsyCr
6dt8mji6pA++v221057KtcettA5zuQ4Uyvxd4J+dQUABauiE/UVy2cZ8KJjeB5O4
i6xnlOuoudSUUnGtX9qb4YNq7dP3AK9Gl4cRBQrM5ZPe0P6/4UsxJjo69Ab/EJp+
9LPJqGnlG9zyAo2ep07jtD37tm3aPfFaC4dUfbkF8q+S+rw3wZbjGZRqDJiNfw01
o1JMT1xyQwG9u+opdZLn6NacLz2QsOo3ACpcEL76zf76gLM+WOWLbrOxtAc+Vfpf
6Alf9jHCBxO2gDj2nGViZapgWuhSiAG2LlNI5WByQgaBU89J77BLMMA/S4kw66aF
B5hzjnQ7MPw1z+kRIWNapmmMuZMWsu58HbY1u9cEnmsDIFiK0TIoYm1k3OZ9SamD
OY0PhkrnnWW9HGwgi62rzVoQsl2tlvRPlhfKC4SwHbh0d/71fWJR9IgpdgRunaFq
VKdxP0tdtABUHX3oCJOu9uDokSPSaDt76dX1/BgBl8DUMvMIRvRCQZESErvs126O
YLWwafH+4Y1MviRYT28BxVvkbP7UjPNBv8VphYEQlp/8wb9JkaLr+o5lwbeasqTe
VinYuVqBJNRoY+fEWHaSIWxEBEKJvXrUIyAN/gHX+nP93VCtJsDMaoGg0ItUdpmm
1ZZ2GzOZ+34SegRNc4ActX/BS6Rq0/WQ2ZTyrMF1RyE9FpPFHCKjOIgRgDXRbHoq
Xg3+xbqMWlYibmDmzqUPx9pvifhwNe1g4APXQmGPYww1e+SyguqZuD0GeFPCXuMu
oQxvjpy5jD9zv2IO84tQvGbOTNoxdWxTXrxqK8Kon+30lYaf7L4XEymUylFiQjfO
z+A2DA2TCYQtKG0NHM4VnC+Cr6c77q78Kr66x5ZZBdcwFso/1/Vpxwxo18GZHlEl
7cqFIVPhx3zQpzJBK0D3nJQ8VOs9wSR15kyHOHxLiEhfeGgcwwA+TXxXbdSkJL73
mWRxaVT4kbzzwbZ2taVxUQu47ihnNSF6W8/ZNJmwifhrn9k+mkMwuZNBpj35/wVx
2PawkcSI65QkRw43x5khbZgvvKu0+DyW77JVjawhuRR52VLlp/QeWEJbIi9FBZBL
oqPs1MksXTdd4foWfmNlJ73m2PkzHL1dF4MEkupTNjwl5gdRU2a7gbDNOQZWEa3A
8TFk2SPAu9IpSDNaXARWia0rLXOsNmmoJ7xRmDpKZzZZD5BibBZ9Tw7IIvL5Pzb8
4ucHwhIXVWkGd06dEYSYtyMkufvaEstfHLf8iY4ItPCGkPONGt9tu2U2OTO/GVqC
DabjODdusfIeCq+Ce7aUP4wn2ID2/0ypxrKnu5p3nTXQHe28ZGIIB1YLjvuL+xSj
P068DI0ExVNjCCCM7qdaF/ZkgjFaa/Roj5j4l75cePkfOchjnbaLDioAnyQTT1SO
xnMJpWT0VfEJBjtKi+ma0rtjF/Duy/+jDg/lD1zs6LWlmKQrQdaSfV7LDpqNANeG
LRSGXQlndaiQYV5sdIoc/QB8Rxx7YzKvO+lnNL+wDAHed6Vf9ytG+yihO0aa2CAa
d0I3wPa2dyonWMyatKhZlEzftR8l4w7JEMJuckdG0BNoJDPwBeiIS1lkanfRx7oS
Ez8VZmnbA8+/vRCLqSQJxohAXgIhzwJAoQqb12Eks4wJDa0Ye8R+sCEMxyAhV/9S
hfWJBfawsnZIH0Rph0a+2tNJq95UfMANkpxMPFugSdgIr86nIRzzzNYEdKPb4QU9
WeLi5dCLIHtiMr/lwQV+9PB1oewwUiBvP2Yb5MsdblZRIn7JBScPPPVH9J5vDh48
R0NSdM+DQfJY22eb64t49nypeqpnt/F5w7IRylMit7ixuQJFhAw/pH/pXLnvpTb5
ChkZ0KC/PzRhh8dLAl9hru2DjMQvBGJyL25Ek+7ARr1g7PSSBzJAu33OsMa5M49G
Ds72ZbuV4zyPcB4446zJwfAajBDWmduVSyGW7PlJWRhD7kfw50q31KFbODFUAoWh
CsMp3NQk4z+aUk/sOtEJmuEUMakbjg7tSMlQ1OgBMcOmsvI/TgrV8ytU3bGavLsu
Uk7NqNZ2KxlcXN+Pavu3FAJMRnCTy0dkPKbqsv0NN63L3D582bL9HKkUL9hgkzaH
Aioa6bb9UDQa05yk96yF3C9lALmds2Z65qooOxtteCGBzMKVGGbW2hzmjsWcRJmY
+R4LLrGgqwovcUvqpk1Te3j8N+DFGO8/OM1qjsaJNcLnLHhwkHnBbq6qWtB276p1
L4IkHDlNsNVKVEcmaJ/yGCntMCqzvVuu/fm8bicPkN1TWIoyJfJt5eR3W27ymlAV
BveBOdvOd3c6APwzVD1HPCN9FfKumQXaYciwiN1lFnjue46vFDl3SVxTlJcI32v9
pk9E2LQkfagjMjhSxY774SUnJfe5DtAb8uL6ep/dQw1WL4ySimqBU6/QFgbVjsTi
uyFR/wlY2gFVeT1A73OrxDNyiBeJDPP7gg3uf2H4AwDueeMpPvcYfyAE6ejD9ejI
Aa6TjLVKTNVeTtcs90XTwBGHYiMRI8eGqaS2tPXM8qUHBq6EYK8Hq+Kzjd5nA0X3
lA2SnLh1SBsMyPLHG9sYJiRyNksvZEvDffn9oyvFsANaT0LyN2osb39QWpv9flj8
P4tv5ektWyOD46B/PWqe4hKP+vdyjtt+ADys05J4PjMqXPnF47fVR8SFOB61b/4O
su2DGCTMRb12yIX13V8LLTfvd1U/g/VeRerIEQ4i7VBbXm0VJI4l1t1jIm+aTgXV
XdSvq6Q4Jzr9lIqHSCBjwA8nSFmuihFl+3lVM2egY9P7AiAehMCiet1uGPXPTsro
WWf8/g9biOr8sLl1/tu+Jrq8WF7FByENF2wuFF2ZmzHRKFusNZXoasoUHrprP4u0
Tc3O/R6rknbSgXyp5RB5M9LSGZnKbY+Pc+91Pppz1ZzyZEN6fYBr6be2ikvcJf27
XUbXqrHNnhCIKPD/jjAcsN2gFLi4XcFRy8Ob+eh/nSsQLOdbcwyDr0YkMfy1mLa9
GH86EhLMd9O8yHjMkHpWlqUrVi30S9bpbfoTT/hMiUqRCoRm9+nUGiQLpqql+5jB
ZC0/L33fzk6g7oX68aimHF5jmNFNeRB28XwsxNd5AcEnpvuoGYlE5ZDpJRQpolIR
ZuPKlcoFzumm3sZwCoNL3EthnTSN7Tc6/iNZFhPf4vkEVEDglGqbLiUBxuXgXr9h
/Xph8wcp07Yult0EJuS1yYFStRZhEvsf/U0cgTTk72sPEki/08kXRPCnQPfuaIQ9
T3tWcbjfxB4YLeBLTukhMLFnCkfE6s+xJnpkuaXOGOrDUJDUL5vjggzvAlFBY676
MVC67CT4RmeJszD0J/Ad2Yaz1QbrJCPll1xOjnBUwwR1EOqmigF7+L2PkFefYL1q
kTvjgplBMzIlid9g2movz7sD76llXny/oO/AKAZ7fEGn7efzGPN5bYPdO50S/q/h
TDjF7Eu+Zce6P/Zi908Tm8+TEXi3FzN7dFE/eVud5nk7U/nQhTFWH9slradRvqOm
awA0oZ6bsptMKqvkAzs7/rJC9gxm48wLrd43EOt3lWqBHGCT5Y/KB1tMkrYoMGz2
EOxGlBigSdPOdFgY4WlKJbujRUwU/FvHLOy8RGmPQbmiEtRhnk6YmHEIUPPVN79g
HsXb/Kq2LoGUfDfpXyBPDpQZ2bteR+WR9tLWCkOt3upaYAjaIhmYvOW8bPh0f7A5
7wwV2A7h2iPqOekB53bdb5TpXBWzw9BKe1RcIudmksIBk3oX2ZYXG+zQhMS0HTF8
++kGt5y8lI2Vh6Y0U/avCekEh90hg4V9v8jY/YsRvfB34+U2ZXsHV1OwgRd2bRuk
YtNyjsMRY7t4MP3N5U0Ga7JaBVD1He85dzM+aKjNR58ZKZQ3ZzsFoWwtbqr9xKEq
X3lNCxItMQ63lqhr3xW6Y/38Z9UHsZPUf6m+bnJg+Sqw5XlqVy/UrQoV0WGolZAp
OgF+Q5bLrIPcrazZa1rleHOOHwZePoYMfKiOoLRXmGQx3xrwYWpFTGJpyj9nPkuZ
GXb4F8w/mKbr2+AYE6NvwNZAi66isGDSL2fXN4exWf68Cyo+6b0uqHEnuyjTBJnd
Ij7hXlNoUS8xK+ImcxJDDrYm2sBJet5jZKUljD42wk65q5rHMPvGLcIaGX6sL3DD
Fv+U0qxhe62KwU1k2KFR0M+uYqMPTG1IA8v4xuDfS6paE0r7OGVXZP8tLo+gyrU0
ReL5Si3wexA7ZiiyhZRMv0gHK5oD9a9791j17pDjOexklhRmPuVwct4Hcm2mDwcg
0KIlvM4gDjvv/7emkfKsqRaXw4CtVgmVShW4XzQmaL7aeTVNC+GfKxnKhWVXvYYT
4hwY4tJ0XvVPWLd3utJvvI86fTVIOIVXcJ+0mORYdKw5skSsdypzcZKMkmob5BPi
u/vQ2TWKfSTp+oGgY58N+gZdLJZ0lw49tFUQb5VVAQGu9hc6Ft6bopdqYOJX4wWW
meg59+ZCIwq4uOPeII/kgzJZASthHpUci7TbcUWxTifBlltcD/cphJAKjyECen+E
Bs8HlHeaOpdHZy8nNrZwqhZhlkRyI8w44t4GqNS3L36z0I6aC05vMZVFw9pJIYMG
d2mO1MoTPaORdeM2/yHI6YNMdP3O6/QMsd01A3HoPVUOJhij3/xEedcGPyUxry9D
B5uZ34dZEx6dIyxU1U4LxlkV/8MzqdG7Rh56lrtRt3tzHyfpOmpI5HBdsphNcs4j
pznyeUayk7Wes+K+RRC+t4YfegLzZQBrk16YDC5z3gsg6TnGbgDhrENjIP5NCXAE
gAYGUv+vvaPFgWvkLci2zxME8H+f+c8/wYXU8B+ET2pMTLpR/9q6ULusH0spr1tm
NyDTzhG4bt3MZyDkt89/PvhyCyaRpSbc1vjpr68WhIJkZr8JBu4dgvEMXaEqVKmi
NU4KTAm+I+H3t27+VNJdeZ2m2pzZizNJNoNBZK91W++aBheBvjK8u0AuVtow9Ciw
uGqHkVmuhKxAkMkcO6PqpTdRKCVLxT/US3O5OfX7gZFduZb3eJhHc8+CJx+JfvkA
g4o1Tyi6bnBtDQzGibrIT09OMYaSBsPGXmQhJ0hXFHBPJZLhcHk/Am3t2q1fnYpV
+d6Sfir77o+FxAZ118ODrV3KSLHDnfy5AJk+litd3PosE7t74gVLjMBoJwsZVry6
JwNVec7aN0+mIBqQL1BWdCI9BWBdn/HgM1tUjmBlsUtAWol52bcgpcXV/6yDXccU
id4ZBnEvtso9nQhTXlVwlEyqPKYgLiDwFb0HiLS7ewPM95WU6wE35j51FZEh668W
Nz0rvnVY/74SQGeKx7T+iB4/Yn3RCPvvWuVsQqGOPQUIWL9P39q7f24JLR1kucZJ
AgnnrcujqhyLtAmZoSwGPdw05B5M6422kzop9Bg+PUAZi50xmkKLAvj796hpvVPt
TR1s8jgQpEmOpD6S/hAcyzfgm9BCspeT5aB1AsY0EQVDxxh0LnQR45mTeG/o2Y7f
hx3cfOF3QASqZGbdHvxcTrX3ZZ8oJ9FUbLWRnKEvl7Zbx0sxnPIPyTkLTCPWiXnK
OLSZ/Tj/Ss5GuPrxANK7Zgori/93C5KvE4HfzLWCZy3F3CT38HWuS2icwbFSmVet
MMZiHp/KjV7+g/sDWOVbF6ipFixSSwlISNtbrQLF2zP6hrs66lcggHhPSVZyQKHo
p+zyBMLTOl8hJIUlrPJTOUaVt80HvRpcZcnVZ2KFxyxceCi3ELeUcGkKXomM0REs
/Yt+wOrhaQVKxMD42wKn2awIMyzh3HpiWRGwF/6N+Q6rOW9nLtUpmzxjOE9U/R00
B+5HD6Y/IIN1kk4CJ1TTEYFhVuc1+C8zv2OCLdc7RlGoJlHCX959213Z8JfkCUxg
lfFx/wQoTMfzeEmheMEuSMH2LSHZ8VKGd51mDv6GWFB6iJoQFt143vA3QN19MXWN
ERZ+WX60qGatzAQu7QQ5dGSOSuuiFdrRqcHyYtTmbNJnDQOPvkI845hNbXlY7ewX
CiX4jCZMqv4uNrS75QlXx2+0QAI8OHOvbCanO5+0fPTW+Io6L8hrDahTqWkchOLW
Yg/3BNmjiajXJ+18KwJAFNu76WlglGpF10eesLf6gpxOgsFyrULB1iB/E/UnmF0K
MuIseccqRjqtJaAM7sigV5CsrbQa+PYhip5b6M7VnuZjYJVsrbkl7zb0Z9u0sc3e
34zXSjpfSsW7qSXQ6q/G/WJ4S61JIldTecr8L1mHBIEUQLhPZwPj7Et2WmNki7w0
yvDlC0Zu/8islTgujikc/ni+f7iDsOhx/3AFvz2Sl9eIRLA1Nbi+HO6HvPk8gjBk
wg2sJraymoPKBO7LAmRhwFU024GIW3enGiYJ+meUairsIBnCqRFKHcflWa9qYBPP
XpiHEAKOkAwN0uIl6ZJMh6mGUhRiv0hen7OOUW8aoZQWlQ/tnKuQ1CV+A7bI2vFz
jFrnM4WHE8OmM91KfRuD1RZSApLxR2DqzQYMTx0Vmk6cNN/VaxyeybNeMfAQa5Xv
9woDtdn/VD8UKbQUCAqp40aG/Z2FD+myD4A0JZBQtRPf427Qrk2Bp4SIbM/9qSco
CqPVf87tF07gagVux0pmVSosxZIsVLfQoxdqHF6sNKNw0dXoyvVrABjDxmVqvRoo
oDRxOt8zSm//eV9KPaJLby2+okJfIBbe6An3vUiE5M/RE6DabhdF7sZmUZ2d9x4a
uKrG6mDnVeSQurYXTstAdWu5Rrf3KOXbh6NkcB9GzhSdDHpBl2FVsMnobr/V0DzS
bItDBt/borbks19yvGXr1nkOZrPxA8YucC/4AsmAF3omAi7nEKlpTQrnuGJ3HewD
WuXxmP1lKhWhmJbNfaAG7cbjiF6N6myGXVoFyc2mB3gO/mGymOtiCNsDogIOdXtm
b5cUDRx9W17Z17qC1DvHgZHm7CQ4HLDMviawjDijw+xOzt+UL7J6htDARQtZVIVo
IqjbwS/Ai5eLMsQkU0LoAs8JiaixhEe3VdW4MFZqUrZKwW+6WXP+BTlzoJ32/8gs
ictVvpmENFe4ilBQXfyd+0rPA8kd0/U3BDKnsRCnEh5PRp4v6hZdO3FzvrmRSvd+
1DOvHwtGLaQdJUnZjZyYuAuV189KNnLatht53fENnm+x4OiJGyNwgnS7r3HMPEaQ
hAXeWvq4mrBLbQI6gagGyU+RGqE9GNzSquKX6sv4FCrlcoR/bqo1F05y4WHoDXet
qkIeX08qMv1JSEStglFHkkuPCM8frIkuMP1PWlZXOk/btILqpgYIiVaFAhb1x1xk
28F8yKyDImubADnNiAcX1UPmFlMcTX5/8shGPs46OA0ykDAHv5tzDukCcDByaQIu
J8f7wlOC4VVrte6YzZ47SZU57u5uC/v237AY1nCLs4C0RzFXdYGssTM5oCFI/4c2
ZtnJdBihzQ9BqQRJB20ii0xJ4JBkoOw0HyGO7pUcki2gN1lPu5wT3xOGZwEEVZT4
LHFZwOb9Eceom2JtCVMoVFto7QsTXhR1KWeV9jShupMqu/xIQJBI78WlVC3Fb5hW
4I4nuL08PG4m5MIhHd3HUt1olEW7/QftMNQSjp0kG78RG/2mxhIT6ZnvXSOv5FPn
wVB3ksEn5l3zMdnsSJbnsefw+NlXZygvgNGJ6AJGn/7RtbpXSHm+DAlhIAxTlj/k
np367nXj1aOe0snW4DNgVvDmfIQ80xUOr83sZHGWSeA02Ao0T3JKsX1P2FrVUI5+
C+4joHVZFQ3pfCIZDlzjK1XObafbUpHUu4FZw6rXCjBc/nk1+8EnZO2a2AxRncnW
WYDxeA6srD4vWgi/vzFi2XCHOSXlCqSl18zO7opUVfoQCWTdmlB7WWW95dt6mgm/
kKED0zyGBPXyC8X/vcFtzbhff8AxMooijL0JoYWQ4+WIkda4+NcBEKPr5Hz19ug2
kGsozv59bkaJ3oSjgTpWrjKhTU0i6Kx310y64TODDD3DSGUErMHscQ5xjx64d3t/
fc2MllrYZ/PMHCLJ1rDV99wPMbE46AdnjyY6hD+IIxY0itrt7rJolCCCjT+bU68a
FdTCBH/md7huFhZUuua7hObkEV+6DAVW3FRk6bgnSZrWQnzWqr4reepVjj88nfae
URktT+3CujiorOnJqK4OK1i29Qsa2ulQlV8vXgTN7kkCDkWFKPkKMVD6Nv3TBiCa
MRdXGLwVE+aT0GqBToRXVMQs6N34CPmllOVu68ueehQMgzE57UlWBCmJY3HothkE
XUKIN6vVMECLSUV+HPfFyXe4hqLMOEScZP2U+Yiv2qaMQkMUGSa9892RbrKjp9hh
smg9S342r3dwYdVfeTex0TYsLwqxwCZjGBlwQV3LCngX66lKRce7KR3tJPtAuC6A
1OCUDXaDd64S17wfuuEOoorvADwNWL66AWzYa2gkCntbOKcJyN3WAvQMGtLSxkey
AmcWEYNSQOHqwmV2E/cCWtvFCuSoGH6en7M/cu3+zO07cNyUDzwjSEKhqfwhHP4/
eA0IgBCHyfSpglhwERZdTIFJFGNDcmzYOyNrNbzdDH24PUV3oIkbevOwmQ8GhdxH
I177AmgtTeJq9oK3MttvY+9xX62ED2RkaTF6GM84xkgA90HzTqxcYuws+sbsgCFU
pwGTy8KkH2whcbGEpDNEtZy+sSavuSAhei6Hq2+tb/QyLBaY0+GhwQhXWbpsCf6y
6Xvq9g74uCsQhydbx+gI/TOpWu97j/Ge4vLxLvpR3n74124jLT34haZHH2HJr1Qe
2k02LgE5MJdXXXN9ojla2w5BRZrmdDkj/yeWg27wAL8RLF35apa+jqniNoSRBlYZ
M7e5UfLQSZ5cfV8ERtQNvevXalxX0G5Un/S8LE+3ZkNOn81eQUosFJIagO0HkrzG
hsZCtOgftExAyJSU3kwG6R3D8wall3jH6PCZo/mvfNFQIjI5gn0jnMw2SISuk2Nm
K1mMoAiS+vnp4sXdls+wdHo/KTb53cI8fkSKQQ0aecT4FodAUCM7/nP23JQUAxAX
bz0482OM7+Dh7We4RkpOQ/IXAJRb+Cxw2mJHgZc7tAQuAB7AHOpS5iH4SPZk5ze3
/8ie5fwqbu3JuafQLs42KeRsaZSBhaBRbsaejSnuiNq008oG3T7FJRajOfcm7VCp
Rjqtv8rDuS37artY+nGwx0Q+UWENQLxsOJo9Y7RTR5EDpGOZBg56uyGHI6HRyZqS
ViYLd07z3+tI9iBAE7gCk3k5pxrKaih7KhsECjrsMK2inESZM8ThoV5Sma1p3YE4
sqfcJ8rXjHDtlHMhchYFWNm6VGDmknuMnVMdc+XmSiqnq89xZYLqBftqL/XGcBd0
RJhD5XbmaHh8S9n+oJaH1++KAQXGmtCagrtKPGev5o8jso3FjaHtOY/lW1wP5avH
ijQySyBpGlVHAO41vj8czlk9WHXO5CzUg8hu7pbitOdCDRq0i8gahEvQSy0pyIep
6Gn+s3NCKCzyLPaKFCH0VdA/6yC5uM3PrBj13tEtb37OFoUQxVvNGUhkvBWiniA4
WAWVwWViRVlYtf0U+PbvUVvtDEJzp5D6cSeVXrKpmpK8zcCyZiddGVbXekj4qo/o
9pSPE/rPH7jf9Y7/CmZIFnP8xc7exLWxv7gL6ZJIu8n2gjOyGuD3ojgNOjsNNQEf
eDWLyr5HFC9js7h9tWCNMjxCGLHlKC/tOqnEb/LhICFBp+uwXzKRu/WanK95uRaW
xwrv7QQ26Mdoty8Yhn0uiwCHbPUSwFIZxcWZYLnjhSKHB8HE5meoW/j10jbLX4FC
dBmUaSLXhHLLsWS0wUx0b+fKsY0EoY1urtfVLWG2uRlbQVotJfIfKAq/OiG/CNsL
AejAIIdk65Cn+xI0GreeYjPD9/V8RhgDmbVWrH4tlrd8U9cpgIDbH0TRHx/iSEcZ
jlq21GQVfAHk/wI0KFDVBldIv4TtfKBrBSpwHErnUfXyDZbt8qmwim9vW1wx1XhH
VrRv1RGhqoSX/RjbzLvl7QdbQDBxZqczIzzkUdISWN72fPOUz6D4hSH25XvtDxl9
DYWbQ2o8nUF61RIOEof478FzTM8aGJ2rqY1Mc7bEnQmZz8XqLaY8cqLlArSb7evg
J2JWhTP3w5xnops27K/7TcSBGrVh4JMXhkbthQgo1EXemfllo/LDpg7G30uYd+7H
NEItQtz2+2gmRVDwmQHuJzkR2DuuLyHso8Cn5n2AMMg6E/9jA7T+emsQFZvFqOsT
a3nV7oR8/W9yUiprIu9R9X449ypVISM781TkMcVwGv2m2ptxHZCucyBq6UCIjOv0
J/L6+nswfc/xi+zJVGkOkZ77lkUw9JhGWAo8t2vTo7p8JKSQzSrBgdn2mkDw1UYQ
qm+RjFO4OTaiTzOfn2/78mUWPNZz67xkR3rkU8pI997ADr0aoLRz1HmFrJsDopun
SVjG1f98GYag47tow4KxLVky5Fl4FpnIrFwA1xbNu4ST2et02QWuuMSe4qI2XZQa
gT80fAlHEtUBATeOVUxg/ka6K7lhDZja4oBIzeQP0B4vHVI1RYDGDIMmKEL0QMLb
2LY7ADgxfUiLmsiQPvICwGBlLOiVxjh88iTsdo5iLg3w25vvX5HUjI4rEBqAu8Cr
+b1nV0cAwx58mJszU7XyPRdW+7+vWwbLtBL3TAFu0IwjJH8LpalTVlOcCJegQVYw
TURvUw0Ihxpknn511k0ZZhwHcsx4ndJ0uapLBcJfh5o40ILmCj7g5g5dpQ5xLfYN
3ycbftIdy6ddB70aEqp84oisjfx/FyWG/Jb4uWjRPM5n7PACu4hKWPGuBqpnl6ug
L+yGJWeLxATzQmohVJ9ZAxzlkg3/RIrGTT9guhSRRxRTDtHZyryx9Ln1mzBPn3ei
w6nfGzWpY36m8QHbnt4nF58w4uUs2MMBJPaA26LhHnqr7vQMy1DxXfbBrppz6lDR
CiVURYOVM2o4icbSkQ3iYpQutkRQlZdNP72jkWrjbJjXra9Mtb52+baBm5ZCRWw+
UvT+sQ6LBN98wnq6CVJoBCXmJ7YQvhgoCaBaiBpCuEs3zmDA1mXJt8+1KE4bx9w5
I2/8Sq9u/LKZgJDPLtcNFGiOVkynsZNEwAzNIcnZGsJsJKAaBTApgI1Q6KLI4RbT
J4wf0JcVSaIKg4c/FcIp1NlhDm93jUv675Epuz7IPEVu/c57MelxOsis8cpETSBT
ygoj0HdMKdO+cVETy8Ncy+VqVM3ImASZjK6FihnIJJI/fSbPQ+5sd1MxW6uy1VMX
jwirsKlI6S6DzZicOrEi0UjKxRa3Am4Ls+Cfr+c5wSsaWDFXK4FTaIMrgAZsyEB0
rt3Q2NlZMDS9aMm7vFX31S0yA1uDa981NnyjgRaUwZqzgjSbAafEDvhsd8DoO2RK
NjxDfsG+ZXKbyo5mLQpcvMq1geEXTNnwYGr8PoycK2y5u0kHIDT72QlgqbbUbais
Z+GZ72uOMqlSvA8QYPmEVOHYX5r+fSav9ZjXALrCKGAfqqDql0jmWUA+NkAVti8+
GupabXigoThYO//Blgca/WpRrpWZKlNoZEE4jQw6wHayrE85wmvZaSpn1/GSAYSt
0MMP6TO49nKp4jMURdS0BZ4WNNcqGUVY2gyjir24fSzL610ux2+7j6pjIa0lbrv/
ja5KjhzLTPYtdMiu2fenk/3Z0zFD6FGMYfhQzJPKZPxzGMfdr2FAh9b8e266bgdK
FfuBK6OPm5tqhT1qrABRrw5fwkmCGQVYcul3CNZpU3DkN++gEabSqqkt7LNoF12z
wYVNSKP2IIDtZSRyov+fcBUTMgeb0Xeb2R7pVB0vtdNI/OjHovVIoJW33G/SoHmr
YHGaguaLjaSuDQkuRAPDMce/BFDKXRU5qZedevgFAfJUZbbXKNvPjtZpBuK8AQfY
SNBIuwqIa8XBnRb4nS3XWjGJ883+Dtrn1KuKz71IrApcolpMAJHMLh3rFG0s4YYZ
yDF/sJtH5KUw6Fr6KUe/6U14Y5hDHJNCGkYOkYDJUhgsndRVdlNFRUCF/qYoaE1E
rHp5P4j3c6iH8JTHNQ3mKaKM9JHvred98qF4SaolNxTE8q9tZfZ3b2uN5b6DnKWw
1Way95PvfRzhf0xReUXFC8Jp2YFWpiQqlw/6Ms22+wUoLxQd1qkySho6QDvyIDvl
s6EVHiU41n1x3R8JEgUjcIHoPGrjKD+Z/tivhCBB45cMjKmxMbB7xF6ReIxS/9ZI
8IClwn4xM3EWI2FKD+dFntAjoEkVkKGabvw3/bG2n/3PBDkavuHoG91EFqlDeraS
Fi2b1akSP+djo+8uHr6dU02f7OkXvRIkmaForpa1CZIspmOatHfjdpbrLgbQPjy1
bU9pjJ3Dcu7XtDjG+itD6CehJ0DindRCde0uZ+1kK5OVW5bjtXRHWNZky5J4ilbe
qaplQvb+9+UGQnjSUaCUC3YgyW5YHVlS3lqtREbCBwnBjh9Y/FuaBeNobTaABUdZ
pVQlcQweLJOGkCMnjSacbhwTl4TUpXh1b5G+1f/VIW2MWI3OEWnBZs1qokFTIpfu
v8b54jGI1sUUoBz4amFPZEWRwMXiJdvKa9Cw6jkEPW/kbx4puForg7NzgS8QD9RF
f487EEMKVK6wVVt8vN5jelmqHe2oEHknZ/gb++q66bnczQON9nBOqZ7Hb0e1iZ78
Tuy5gz1732h9Jte0V2BYJ3KnJy1WFJW2HxR7tNet49T0jT1p1Pq8LnaPaGuqJnO+
scs8GhnRJJqbdq5zvxGNwrMO7REXKYSXhpmC7A+8V3IMgEvumcjjbKnlQSWvIvKG
Um2UtBwhkIGLFsDmOPSo9ZYbPXRqCJCdyJhxvqSUaL9Hg3N/P1gRxVrxcQqh8xsa
hn/ksdQ4VDYczmjZeYMbgQIpiQDIAlHuCoSdrTVe+p1eFtT4eZS4vRqwrhFg+FGj
VS3UJmPjR8ClnXEFbJq/XcaTRuV230d1rNh5HAtdf/wlB20MgLnfyPK+t1H31sgw
P9EV0h+HhmapHxl9QooqhlSAuIBvr0PMEwLQ08ZrxIZ6JcdTTRvXGCEzY2QSekew
MfxfjfEiC0nL+2OC0dYlJLYunDhZ757rePcwtxk8xNKnLzgcXlASQKVIByedelDQ
fVv5NIQlx28Q1PaBiSnTDoB5wK6DIIWJfkbbpSpFjWe2zDgwQsEDWFuwraYFHLuO
aZYEkWI24ff3SHiRZboY4rgrfl3RdJo7oX9jzE123iVKwzQO2LvbfYDDUD00A14V
3TmdLcvBVEg+MEu/V4cnNJbjBNflvKOeqDaVFnqCkmOabjiNMq7BGOQ1dbUsr6LB
nCjsPxZg5YFArQ+KY8ylkWTUjQWTmPwpYvl/uw37bWKf0lc3biMC0RgpSSw50pbH
4iT+yu34dRaNOyjqP2XYM+qgHnFV3kyU6P+mH1RY0SKewMwFUomF5ltPxhpeLhta
W43vlhAp07m04X79riDVrwGih6hVkNbKkvjhP34EJ4UC1SEzPlTd+EPaeMj+oIfY
GpcdwqkFOHBy3CJ4Ufe4eyjNQOTBq2hCefK8aAjthMQGsyKDotYTMmEP2urBivJU
0y+aNiFS89XCChE+MD1hNMOOKNsoM7w09ZOSAaVk310TGZXL5Dbi4Q8//l+hCABV
hMtYTjHcP2my8bK3v0iNjffBGRCknfVS0L91bAVmX7/j7+/7TgwO9Mw83lDZZCPj
1aT4XECibVWOlVE9rB83Ei+4BgTk63LsTl45h54fjyduu09rXKeB1/2rU0LGfJ/0
uXDKSgL08UmUO/2p7ZO+4iLTr6oPZnmRTWVnwc2+7KiUQRNIvuKKzg4+EfEM9lS8
nOgUuRIpAG9Nr4uZ/CfGxUkr/7waTs8b2MH8f3dZKqJXo/hKaq9FBgSacCnHNo2N
ZsvjC1CLyvfU10BjntpKuuVbQ4KOPynL/IMmsdk4rF2ikhj4R2JlC798paY4ueow
pxRsCUMpgIZJenh6bGJEeUqQgTCxxT138wkUgNYyNZ5U9GmrzliDHzhkVX7q4wPC
8BYwhDBLxZEuqeTk3zQSeQedtY+t0//cZ5xRChS5ewAZLb9u+WRBBu0x6sXvYbgy
2cP6iAd49dL8jd1C/93+xhoErfcEf5bp2gZc+L0GYkK2J0ZDkV9s57cKaa5hZGKo
+WU1XmZkb+tO7sZ0SyilSZda7fn8HUz3WUxnwgHWjrBDwuLu08BhV5GFBb7hcezw
OU0lJzZ5ckjtAnCItEuG+9/m42pMdvRRg3puy1z236ecUhZge2nEvU6O2HNQ5Fi7
3cccnxmHcfvE17Fpk2DekWMSOwbYucRZimGRhp9Vgdmw0p84SGNiTu/M3FafIV/W
UxuyCzWW7XWeIrCBiQhOesBD/QeaikXvhJSh9Fi7EsPMJP1z30wilv4tflRJ+36C
WxXA1ZmG8gkutlKle7NWmYCwZiXJMtMY0Ckjixe0gzDnhowielUUXj8AptfTGM4x
X72kRCQG+EEAV9UvF5TE/bsfkVxRmaajKkLC4DWcJKKjBfvBnXUgm0yUeR0DtF9B
yjtdU95N7JkKeMBGuUUx9dgYqYswjmqS7vZtg5c1oTZs6TYXV1nUTL9tpnQnORrL
mmm1JdK/EHIMGpCkDIcc2ldP0W89qJq77fLFVT7SAqm2cRcrKaMhOPJVVhEvnICY
b4S37l/vfy5l7apYxYlGGLfVmyBN4k2CojtqnElNrflO2abQNB4iUcCVpoPblN22
fZmG8ThP+tm5PlIXZQmYO8LDbpr2+GG+GohF2YOvHVbt6XHZJ7/xFp2OB6w51nUG
4OgAbMAFK6Wgo0nZNZ8rHfmGG3t1Rh9C2uNF2Z+HekJJOpfPaXBVOOYl0Nrsd8Q2
7qZ3ZT8zhUZPYviyFP3OEYqogeJXQ2UMClXPkPI+I+mT2aRp/6qV8JKFvu4wOjwe
HISpFsvMPLNp0ABWhuDdO6VMk9RnqQndZTK24OWupMsMSTJ4teKWf7/ODv3mD8SK
IFhZoIBHDHc0eNwGZIwrjQq/CJeBrSpyhTkSbqeDwKtamcprw+fXqy9nmUF3FFJk
MUyAuPDr3r/kE25sj7FPItGTnX2ui2vdSrFo6/9KhPyHx4ZM+4OystOi7RaM8B+9
jrI8AqLMzimDpT55vbcPgM390q5ZaW8yITtFBjlvvQPmfjexJ5Kh9Jb67plL1ijk
7w+kvBbdiNpdEWD8eHqmwFas+LQnrOsQnKzRC3iFGp5SlIq2SIln0K5FFXudbnRs
boWm3HiSipnuQ2JbLvvv2GDClZNkx/M40dWOuDWXyhsYYIREArslb5vU/b3MbVxR
kR8s1264O378WBNki16QjKbNPkg1pKPyzzwu7lPORo9Z+z9ux60KJEmfFFFL39Tg
uQtDIE3dlwPGUQnVWp+yNSGQ54UyPBQw4Sqc+UJWE5E4KaNergvj7n9d9CmwZS4R
lHOLZSC4ye/4daWqmppoGXiPDaN7OzGSVxkDJ0UPuYZlf7gxy7y2/WO0TnqFNj/L
LFKieL/cOsuTXidQM/UvqycHXLlKsnBXvUwHx+9gRPGcf1eCX5i/2/bYOIBSz8bc
+f/pp5Qmt6Q4yIEgolnTNSLnUrTjsp8A3+Pm+Y/hrIvMmLSGkNM2HtQKYeJXyydc
U9eyTgPRfqDFr7slPDuw0TMZcor6tEKjWCrcIBhnP+RAFhXyBjUDiv84Zan7QsA/
8D8K33iwqE54DUXDNGxcMVdUGNHBMBIiptbQWn2SaCDJh0NtS339sEGSx25NtqQ/
JCAvPz61qtNRkhkEkTkOz4nPRzLkc9vUC4q2WIrKHbp0GbznsyFOJoeBb/aPPGCZ
vRvhL/wMF11NGNzXBp2XSoGvrpR4vChBo1yTXUBX36uB2Pt3rME8n3AJ2RnQu3+o
P+mr+GQ1M9bdm5SDwcvm9BAPulhVStn+c8UYOKtvU2XPWRwbBxsqLqm2/Vdmj2YK
mnicOEj82aocQu7cXJRASh6tQ1YO52YJ1oC+wSrVVxWsyDi7GL7Gx1HfEoVvv16G
+kyKWVuq1N2z4ItiwsU9DTniRelIkhTV1IG1gqqyDVtXleQoqS/DdqDzKfks7pu6
sbjoznfd2DKzRJNGuvruVFbj/HE7ejx0RTLL5O5Y+wpYpiW35Oc8kcegFajXVytA
6V1LHZrzfRpiQuDqEwPyIqL4+SuH7wKKU5ngsJB9uB2BRJsw9gmQl03hXNcMFHP9
jy6EGrFcDcQ/Figkx7ulPzURMCSeVg2rhwZt4GKgrHdDp3lDr5hQGYab1qZocPZa
RKnYzFr1X4+sOwyg4quo3N0E2cYZIW1LtT8QMm4k3ing03nN649zW1QRtc0l2ZPf
wbgmKRgnZr4D6Q7e7oj7OJQHDqqZ2kxxpikRvTSWptCR22exgZNOvZNGcoAmeM8i
D5HGCBmv5hTmonJVxcQ+4QCNOxCu2S9e+gn1YOjrOZufpiBNPjP9syZiigzNgRN7
4gIioZx01IqHfhTKTZ198xGTK0B2OZ9+is43cJyTbFHv9gaUA/7gsniFFjSDLlzj
Dko3r6LqpJK/ar+l3ZvTMd9As3hihUW06Zp8ITGST7io9ypN6fucf6VornLl/N9U
bbAJv0JSwc8HnieHdKqxGAlXgTuyPPGN8XRQUK8TT8hP3O2ToFlI7GrWW1KcNDjS
u70MJj2BDMCjj+LYD8bZ/D0g6SzXi+rhVzNMEmRyCKupfReZzglGR6DHZGdvj8zX
o+GxL3k9G05SibIWY16FwCFG2al4d55r66FLUe2rq6ONWUt5iSRZdc3OODNSgCPJ
sCovy1DETwAdTxwtN+x4blROf0ydmb8s63zVmJpoOZoTrFMQmkGpZOGDR5bnAFrY
yyVUeYDpCLFdE+zFHs4xrksBFrHVRuHf8/gZ/HcrxcAW4lZ1gIdTZDFukgdZk8It
P/K6x/xPbWMNzaxiIEZjAewGsEcTsNkPsHzZFqClb2b7YCQuR/KTF5LZhKcQOHaz
IHfQzBnFG0T0DChG/8Dl9dq2a7kP62ViDBp6QXb0jQ4dRKxKD12wUMRKwXqREd7w
DTg0E6+c2P93hnp3aZIpIfAAWvpQIE0zZGpiyMg3I+GBpR8iPpdP8bs4LrS54pZi
4fp2UUMdhbOrzv7xivsM7kWCKvp3UicVk6FMp8E+oEDvox61rp/YdAzXKkSL7WuH
1D1Y41ZRQsqJdN1wJHDeapoD+kkPD0W34gm/iBKdCOizdkxFDohE5x7t8bGsmbJt
zr1RDmYMYu17zLy50K+zIAwsk6O3iRRiFl3rPjU6P0D/6VzpOJwgaN1w3GZfYmMq
M1IZEGOH2AOJZfeW1lZDr/0EAg7nZwP3emYVclqooegcQxQOJouG7kDi9drnKefu
/qq1H1SROX+m1CBuHQmEAGz4D82IIDvZ/yHA07G+Vunk3fg1cS5k44C9bpvmy9bg
8W43RGTtEkDffxZTw5GOUDBoVPZ4kCw7X0bcSPaJ1fGaGUf81CKFobAlhjZ5GhEi
CED47+yRctAxU7LnwZaWByZMvKdrIi6HbzCXuIutay7q98uzEdMMhXMxUiuctKPP
iSUhCV8djNcO+7tUTqAQIP7Wn2EJK5vNzp4rNjHltZzvKN3M/5pLy9mkfbkhkhLK
V2iVn3kxWvHo1p05hlRgabfeOtf0gb/xxdVaPKEBVWaDSDnqFNFlQqrErgvc0FFq
Tmp9xKs+ZUidKFWwhhmn8X+Jp0EqNcsVkzMZ/oRdIs7klkPPrgJEB7iygUpAcUpU
s6K4hLsFWMdIzAnBjbutq7SeZ/Zt/E2IGWyeHBf5o7j+vQTprsNeUfK5HkuMth21
4G5v8dlYQhm2xTVhnNXg9AcVch4g1VBj988KxIuFAiJOvjeHPILyJGCKW84egDeT
yFKhw/7w7fJjrHC/kFIQq6ZMaBRv0GeOgTZuHn1mrqvAR7p5CbIr5Be0KQu37WnA
n5t4pG67+i3FA6UKF1cPCPuVOWguuzEmTzPaceCdnmYXy77sKExpUd/kdUXy7UlH
8XD/z4XzLaNxzhQVaY+7bQsjjOabDNo+VhFIfHu2bdUfC9fNYi3wysiJjph+yQy7
ue/Db/Wohzwih6DwnQEsNtEoS4ShxBfUqtAvQIpFk9/8wz9sl17gwQda+8yy4Hnb
5DvKD67ZU4cNo7SXMohzwNTE4rzFe8uZBVyqAUkC0QzXUv0Xa+fEO/5vHdiL1JFx
7AmJMyE7c3YUWQOLMa0uz0yj2mqVxLggR70KOWBS8cZOAL34Aw/jjQOEcVEAm12V
aNdkQ0r81nGINC9ofq/rlc/EO+A2cvljEVxbtv2aJ1wD5+gugZUkylrVyw82x/s4
pLZUsotB2ps8qopLuO8VYqUD9qlsRQw4IxMyqU6e+hWq9qf/uETjCwHdH0GgFw2E
xvtoiGCCn4Bgc7Db82fPHodvMb43WWmxFNM0V2M6XNbO8O99DuxHhEqIlnFAT4bM
YksIEmFIabTGnmNK210x5JTr/xUBpCyl+75oUWl8FZRQWFUEBOXR2KaA6QqCUs0M
LnXbYQKJbdEcJRS9LaaIZpYUFiLS9jceBJN2wF0yHrShZfkPvs7AKAYC4rUtDRuU
Mml6EWo+dRx3h+IIxOenoUnGvSXO7L6Mg38hMwVIevMoYHUKWxC5C/rHgvsTyt8h
6zTv2UDiqrIT1p1vr+jMs/YLSTIQtWelas+4IF18jrWRFCvrW4q8jUlyH80g3/Eo
r3m0h1vJsiInv/+JjzFQYvBflpgOQz2fe8BVdYKlpuY9SL734p8mN1roF14BXmkb
8CUhotbiAxijesxeNhneKAiJJsJqxVvz9Cg0FXvP3SeK5CyPnqI9wth+nBToaXJ8
EFJCSukqVkqdXYBRnNC/NpSxU/1VFfTHECIqpLr85WSrTGhXRS8zcF1tqt3bBFOi
EEUvClTnc6/fav0bu8ybc4/+TmDTLPMD/5u4reL9YI7Lqht/j3HoEY4O91EueV65
hylbPhpN9jf3KTPCpGZKVLdLNuIitEZ9R9PrID/dFPmjXVBMl2yu6s/ngp+u15Cl
rDW9Uk7lEWG01WU9jx8VGOOA7Vp8umLocmiqQyx2lNj51DgY71RBGjY8iXFcE+tc
umKTLBP+ej9LrblgDR5HTVyNo3+h8v/YRUC5pShvjDz/VwfgMwJ1ORYvF7+KDOZm
40/RIzsrXs7AxQJ65wSKNSj5pBoLR2lfXDxAAGnZgEV/V8r2sbAfNwI+BJaKODes
WLw/KFratANkxIJOwMVA28W6kezR006sI37lbQZN3yfOzN+xcbFPRNI9PyHMkZPb
7/DMe5IwdVYgFl8bBBOwNwcYOYyr4tI4/doFQtwwLiv4xjYXkYOejuRdT59KGwxG
OyVJF8MgNZNquYGSTaATNPHYBZqWTywa1YIiZT5l2Sl56ujTy2MjDZTh8hlpaE4H
+TMvzDZg/o3AXrojJgs/zj6QamvlrZRigwqnRbF3oU8A7yD+HS4+hPkM7r1cojXU
CcM3lQyLRRPPljPW7+wh8Jm5MIG4FMjStH45wsYQKsKjF1J2cEVDXTSIdwGEkXTQ
t8c5dcWwB5P2iUPmiEcVUt/t8xnT7tgK7HFbZK0jVFNYiOdIfnKAt7zKs5t3ULIt
4PgvI2G/TzVQu/Y81O33cWCkLGMQ5M9FRM8bDSr1EkyrfLvWHnfUAUlQU4vrDiqn
kvEmDNCOoHzoY8h53d2pe2kimdfIO75yGhhAYzzm4ZBXdj/0OuTAS4rhRaBbhXGJ
M7OxDo2RVsl3V63YSgAwTXs8ef9/d5tlmGqqC5LVkze6RlY6XgEhve9N3RKj3Ao1
2oGXmrmmMdH4Nq79oOdFB6UEI1ahJLL5XnWVhZzEzekua2mokvp/KwBO1QiZ9rel
jw9pPIL+DC4o/cUxqduNAdggPnQh7tHtR/k+4owzbxGnxtYxVrWm9fWAmcVP4LZu
XJbW2IRHCBR/VrIEBUxmB7Li2hcRt7Cj6VsYRRGhQzsQHAiqW56Ebk3kAXTEsabd
+9Q8ZwqzI4fHoujimugcXJfq4thBFmUW6eWIWr/geOluhdz0atHI1F7TuNb7ec83
5+xTOaMhn3MSQpERlvHETh6EGy7Gcr1v6NkMDOk/dQbVOKLp49Hynhj+JUzJsj4x
d2eSZGDxcrv3s+6ioPbOTOnVJ3mubZckZTd0HReFKjjlv3IIZiTnsFgfx/GOMjcj
wPOzBBqN6/bkiuefvX6fPiKndHF4Q9DEeLeNAaYp6rcq8SwN0gCkfO15foFtzqb7
31orhNWNGIEcJ+i2ZD/gx4toviF7sXluu9hjS2D7jx/wy32eEvpFM5nXagZ6jvaw
fiCah/oVO3322lCeA4jtWvf3i1ft2O9OKFllhRu6n3c3pR15RRMxCz63AbHuj5Vk
ise8DupDeMIQTQVCiooVES5rUfYpGktVKbMJkdCMrNm1KBwWBh+u5PTakqQJ1HzA
EoX3xkmkBerKx6v1weEzUcX+QTZn1GpJD7If/SofLcZ2/7H2NDdus0KbgOXk08Q3
tjdBEn/315+1ahvC16gsYNVgYqDi9PrjfQjukLXQg5Rfp0qdgPUG54KaC/dOQwja
zVZ2crBAv/FbpRyLI+5rbtasWOh13g89fXbraIdVWoLVMhCXebyoOhfx2N8qQk+d
CDcNNY46hUDXgMz8UTp9iyjnxcmH1LCLKyWBignw1vv08ZplQmP4yi4junDzzaLk
DrqctRR1B7AWxX8P2Edq2dl36Xgle1nNqxvRrRPOAm5S/T2H1ZWA6b/1a4isH6+9
vfGk/xJE7/4jW+Vqd6734bh0sMlzdrCPOWmhn+vPGCP+G5ivzDkgaU5KTFshGFFa
2TtkisTKbPge2tQZl4wHErcnSTyCA1KXCcreTdk75C/Xw8lQTsPHmVClZpfyCJNP
heChizD/OO6+aIbjat+IIh85ilYBchjMogdB35SfgfLDAsc8kkokopHZrG+KKjNo
ECMneKvWYZbHmYVnsInr7us8BqV/t8O6wWHaOBh9Gfx31c9u8sma9jnA+ugPLDLy
PEpQL5UbwVJA+sBK4CKAByxF3J7BkbBkdBRIxr2Qk4rmk71lgAkcFKTKFiGe6Tct
puLLB0tgtiDBvo5gqS9x6JrRvajUEWYISjF+8BvBZAyisd/LUPTbneM7yOaUEZBZ
QGo+QhSAUURBjng7p745JrJ6w0I+0i+qDMWPlrjLB7feW4dtMLoi3P8k5YQ1cg60
DNfHufSblxg1nX0URqYCE+bfPgaES59PSsNCkAmMUKS+LEBQwJihMv87FL7M2Ywr
zntlx6QJZlfowFH6b/EkNv/OjOSvyPUkwGTxZ4FI+/qd2BZmYwg6WjUfE/Es+N1x
o+5FT1achwWD5DW4mV22vtJfbdK9/chzkWqtV0532mYh8tX0Uz5n0HrkJaPOhbmG
xZuQBI+lGsU3iYmPDPoSQplxkIbWAFdcYzAxE0igeME2Mbn36gBbICmtW7Bx0Oux
3N/Q+swW48bnFJo/z16L9j4Apdyi1yu1E/DuJwFp1TV3+YshnGaM+jmdpkEwgqXD
6qZlCpqr9YHBQNI93UstGassZ+0XK5RpQ1mza6qi45Yig1lu6+4JYOiDNimmGjly
7Ua3BLoG4wib/QfTAlmqC+IhibEohfdeblnDKldFDaXmZqxFvuwJmnWpn9LQ2syv
a5w0wMI22ViJ1RxIWNe2A6QOLAFdBHjWQ5wonX6D5AWxM+z9Nn2P8xVjUp27zcik
VliSEqMYYimXoYw6+ZV4gTt3PAZTnc2FIyF/qk564yioG1xV25b2H6+aeGJxj53s
1qc6C0iD46OlIOIThwEV2VNOeidqBN8UDqgTZ+kUMbT8PemKK1Q5wfH4tHvLImBF
n5J9SStamGuwvQb9FoOokTqudnhWVMFtOc4uatujGbkkGOKX14ekxp5N+IIyS3xe
5bFNqkx/78EUiucZn9YppHY2ATkZvxq26pSVNr4yfu/aypie8YMZOQ1bdLeArKsd
l2jdNEOgGgeJCSNjMqCuiynoVQp3C3jEDAF9OAdj3kCIDnMj/2OnNxb2i1c115UI
CZt12HqLMiG+j6thjajYzlnGVtBa07RNRR7jTtKh1NJ5gFdg7ZsisT+eRZJhfQ0u
GVUJys+Dd5i+RfCkQDWMFgZxYiQ9q/ybEau+dDf39Rt76efA14DDrz4bgwYunsDJ
wZBixpldDMEd4DrhNShyIZeEil+xN/0r4I+LG7aN7g8r0Xj4kU6SP9Wq43wwARCQ
PwPavoPbZ/fs3V1uXcKTguBkHEsgxZsjXexjwgCAcm7m8cjW81NORm0oKZIJ/bwX
Og2EXv0j7n1CynfX11h4CxQCb3jRy6MpjsbedReqXHKGlE3Ir22+qXboS5G6ciFO
IKug2Vi5e8Y6XZPdJ5PIpOzUIU07w7G6aqldbMNMZyoUg1PQVHDSeOehXw4+G2aR
6lKjUfM0yU/Fuy/SI1t+BZh/4qX8fyEx7eHQP7g/YbKCL18yBTTJttIhTCpVCD0t
32pHu+ZeAoO+wdSonPYBHA0a82dtrCTod72qdRLAMEubsGZp3nA4EV0cwfM5dEfE
1fCFiVOqt5CdlwRyPs/juO09kaaLefFeg0IdKbd7iZQ09nvDd1gQUQjjfh6klBLk
A6cEwJgz7f8CQVnCBHaqPoTmmtV8Q/5louq/a9q7wwb0+F7BhSJqInNZvclpc8AZ
sxtrmLlASeAWO6aMgXVAQokV6s5GugHA5G6QFk6sEjW49YvYYR4E/b7/qVamX8OB
VSXGoUMCaJMfBXYeZB6egZCyGNkNHuYISwcZJhsveJ3AA5TbfmRrGe2S+gAIB6fS
ja4F4HahcwPlWDclPiCzqqxZ0Qkcb7grTnekfQj+1s2NPpcb6/tPsNDrxNsPzvVc
rSb7KG/LrskHsGMR2lpnlifPUzAPVKvbbTvFFVOLw4EhsA97bfXWT7ltHbMSINp4
uTEIT3/80ckMfuGee9JBIK0FcRcUWKdbnv0wlRBW/bKVXr6EerCoAyX9FKpnoDXP
VJE0vlf+dc2ncXj6ZZWzykCO4jnqa470a22yhee05brdWUmaiGLkKq0cVh82lv0C
36pSSlJE/hmPtbSnG83Xk0Lon9tlB1mMPUdLCMrOIsv9VgY81mn5TF4WFOScxzCg
RCsQ/YTzVpmMfFxS1NdeH+vB4Hq5aijFKVyUccxrMBTFXqrO8iik8x3La+gOcR4N
KO/kigVjMz2f/7zAlJCxlcBsvxQbAwxMMn6JcZlbe2iekr/TGKMvMwi9A5evs7Mx
PXPBTrkmF2bAPhjM/qDcIrjR18fEnqKJthkbOO79+GCaxTgO28p7xeJK2pb27RBs
lZdV5by+SI1UZb3uRuYw1fOq4fe7m7l4z4dK6IcT3K1Zy3pzbdGuqAGzkoUjJXO2
lFUrOzarxzgJXuoApFimNKZQKRtdq1AYBnzu1mnXflqG87jVY4ub02KWO9+4i1dg
uzmUwQgCRupFW+QNRpcTY5cfX37H3xSDiYmQnOXi15UlgWAvl4XwgWSZRHXlKo1o
3gCniplBDTn7XwDPO8s+1VZzfEn8FLk0YP9toC0VsYqLI7xB7lWLUs1bL3aIcUqc
tz7aDghsuYmEUJCglOIdYv3zk/zlcrtCBg34RW24DirZ9DObqfPhB3c0vZWJPI4Z
8w92u9pOybFiKjHG2JD9f857xME01xxzPvkQcaJO4zjaF9uWKcPme9l0Rrvw95Ic
a4o7pzJiv1CIwg09DMbF6oywnAVsVRZouPw4I8XTss8BKCPMwnAOB30byFclwYeD
cmbqKI6ofuxVrFars368XPk2U7h52+jtAvdND/LwqWgICyOigZCr1H5UUPHzvr+F
ip422EV4AQ1xII8vLR1nldOkatYie6fCivskZgViU33HYpXyGG6uqMz1TS40DgbC
yW5kVS20Tmc5ww6gBScxt8wnxhxB0fK2LzEkiseOuWU7zVMXnXQkR5mF7+a7HL+M
DF/BcvqxBqnWhn+o868gMzpj5QFMIIyhPiff9xBw00f5GqTt56mIwmVUoOccP7oP
oOx8LjqbUKLpM5Etoh/SPZQQV9RQzI9NyCAuS8/wAaY9N1KUlnVhcS7dgpYNSTA9
c2KsqeFZZTZsBPQXabBPOktZXN1ge3PfMaZFJPZdaYZ5P0GCoFfTLsDS1ACaJe7o
xrW05d9UJvviFbg0cHqmTnOY6d8g8gcmxBBCQW70L/0Gwsh+nlfLIieHXuZpVGQZ
Vi9/NMblK6GgmB6fMR5LMizAL907x8zTrvqCgbHv3k3ePK6Mp2z5qe0noK8ZnWC2
oFhtrx464nAUGUYh2BxbgEPwtp8SBWjPXiNaw7Pj4SdunS3oXePdQe1FSROuuciZ
geVz5YzJEAlXXHVNYl5ouHlkGv4NeZiK3DRhonJk1yIbPrmK+dRpI6XaRmayns3U
EYOgcrHwlIp+QeUCZA42M934QHMABfQ4IGoF9ePH3c7ygAzQpcSPZyXpPgSjSr0L
x2KeNwuERu+mDMZ6+lJXLAqmcxyy/ngalZX70zsfeDe36iYICvbc0iruJU/2y8Rm
pgLsTxGJKHjAL5mU/ftXvcEkFFQof2y+IB2rH+pcGGTWks6wBoeyYW9/c+qo7rrV
gTu7L+/VZ4yz3hNWfOZSCA/Rtzy0ZhD6BZY3HT7EhkLYIP9CjBIn4zSPlvtK/zpB
Tv3E4snjF+rTbjodL0W+s1mKWaoyhLZUovloYmoLi7+/3ENIDdQRzD335RLDsrgZ
51TLHQEGqBAo+PpgNyGcBlB0NCNKudCArv6g3kh3ETCfrIVVkKRnyoCDvYb2oRji
Bd9LWL0x8W1QSuUuyJIsPUa+tQxZJTLqSBusHHtrPc94FpTckTXuCH9TQBoEh1le
m32vv//VwTbp+BBBHC9y+jPKor249PWl0opz4jpdQmcwDuxtz3VsSK6npTucER97
FQ8qwGFMq75nAwHIauLcVJb+oITo2Zm1PERyib48NR/swXCPZErTARXdkp9Y2dEZ
JoO36ZhdOitN8rUY3v4oOvOhO5lacpTsGEJUq3piuoQ7d6usOFQXB5xRUyLNtDDJ
kzC6n+RId29cVozUYFhvyRrs+zoDYojo5cDi3+fg2D7PUvDQG8eOFgBR3kzu+iFj
R6ysbx4XxXd6zj5UfH2t+JnHVODvBcQL9xYtVfkmnyFHEVlKibVi5CcEZkOzApEE
jCCI+VhpBBQ/az5uQSgcnsEdZescXWw8MeCQs9M2G7mt7gSv9MtEvccZhfKCtOTA
imDGcxXQuKbAgGPxXHW1jmxpztaUBvwAi1iLCeLVT1Yu5zg48nNmdZTYXgTPpFFH
BHlQALMCa2G9mVh1c0k65jjGNRgUv/ETHxsJUR0MozpDXdnzkVISRYUQb0u9xSB0
iXCjAJABR60g7J/4H+aQ4KtrTlqF9z42afGkYNOyE2ZUHqPisuqffOjV6OlhRd1a
Z+m83yUSJrHWMOYG6MwXkBa/jbxpcxhK/C+4yjnDLsxkbv+U+FfGtb80CDsJCGsj
HLHtyfApQryao8x4UPbtOdIumh3K7nHCe31cyMLKk2sWP40TgbcOfPFdf0fiz7yS
55tJ2wFDSkv6Ft4JFY9PVPWvah/UXAhqV/ZH6zT1kP1zIHZJXdqVzLQ4EYdAMn5n
2I3NeQgXDMvSc1zS3kI3MJmYYbbLCmBfGntbKJ1H7QcAZj3AXRW9Z3+RMCvhzTKq
j5JltyihE1wPUFtvEMvbbRvRcAUkJB4QlAAjcOH609GDeI9FcIMKp1ynU42wiCip
6rsCTV2nqdpri6YLGBDOZNSYY6QS4faJkoOVNTEjSnmTiOyrGqc7A4H10+8Ru93D
EGySsHZ01Xv8OptNm84NFIWYAE+STlK+osjqgUCo36RwTafN4zo+mAT0y2TZKgY3
daAvDtb9BBaQHC9EnYw4a/JKVy64sdVjWzKhpSrUJ4FB9a3Qt4rH9c7MLew3S+75
mGibJptJ9f537oEcXWmiGdAPB0HFWWgSvtxPMpeM70cromCMcjJ/srpG0Mpu1PQJ
Xc4xHGZALxAATByXQINfufyzYZdFYEuP2JKlXG4jER7NpfnFv+a5bDzz5mVzSF4M
Kz/JYUrVc7ZlBoqST3xYQSsevDpey8/gftJ8zF8LWmmosvtAK8DKpPIIVv+AZnlZ
k3yrYDLYkYTEHq0YaBkYKlZq0gdgtGn+xB2E3R9R1CnYtpXA3mjO8k7+1h9ZEVjk
fzWRKN9cf6VaSSMYhGRLeMcgWJ688GAy2OiT4AMruWz0/sB51qzg3ZPgVVGvYMvX
25JRzLYZnDMwg+BWbl6FBw8fMD2wl3B+1G79mvZL+jj46LSZrMLq+6LNClK6T4Xe
WJNJzSpAx+qkTHJoSzowig7NAR3SbnVK5+z2zKxlfzqddYBXBZPdCFjQOJF9UH7H
1Efe4YRTXhhfEGf5cK9bT1YXcdQGhEg8MmCBl4Eka4AmmFZ+yLK8k4SnxPoSG7jT
QKiETErlUtg1zYi64xh6iSmey9vu5VHZoIaiYPBloqGw4msp8wmgAfYWDCl3ByDo
kvHARiLx+226jwTMg5ZmyY/hc3WjuoTh0ihr/ij+yWos/rPeco2p0yoS4re3CBFA
zEKJ7C9tM5qpkEWAO0n7x3zvecVLCb28m6V96RIbsuSlMYsy0EuX1ZgA9MB73vKZ
2/YlwaCSF4aTNaHDCncid7EiBhR276l7q3Wg35ie1Xo5yN7OyOo6JLBSeHvxxr14
fpqbtIiXsR0DEDldvmdd0EFfGqDdKmYBTLiVTzUQ9m5/Xq8PT+2N6U2lHURPdPyP
VLwhfe6OpN3cBdSCS06WkK1wUHpr4TAHADtXpdpzIng3NYPzQPTwxulK0fl7RrIJ
TsTAfERhCDT0Q/1Mr3HIocH1w75ju/kRz3e4pg3oVHHBIjYzQP6Sa6kjEO0dCFmq
7wlZ7VL1Ql9JIvLHErjGDdq3ezWS9KMyu2mgsECYEJ4mjlzsccvdx/2xKgCMgdm/
uKcBRhZoepwW3jAH8uJ9wJP4DT34p6iM4Lu1GqipuMdaHQw4OEaVcyDkPPZ7j/TB
XFwxnJAsjexygdlXLctSk6IN8bUX0FHma4COlf8biyCeDIj8IDYOdH8qiLdNIbdh
sumn7xtK55noH8Dx8BT6zaxRS48XZ0PU8og8JFKvtLEpPukiSuQ/CdnM6bvpoJXe
B3lVROHlwLKTD2lgegcfbf7DxPYmE8ABYj87TP3VHYGCUZbRbaHtyIKDIpE5h45H
mD1lBBQ3vfr/7y7HF7f6gWBD/M9BQ5kZEdHckJYFrRSlqOdH/fizrXHBvij9metz
mulmQ9ajdVx9Hl+xriew2CSi5EpgSn6mrGoZMk2+vegG5Ww2knKtSCny+AnBu2oU
SNvBuWuDkXcIZBUrPNRvjbk4lD60dj6W4e3iS10KJMVfUdFe2AWyvbITKQyn2Ppt
vPGRGftvrsal7PkuJZauc5ugqSkD2WcpdGtEXP/CScyzWjnKnQfHTSc099MofHox
zFp6SDwV0DgsjrH1013h9MOvcdaPENdCAvNzleJ7nOt8qXI8RVv2TqfxcfV0Dewd
Obngwvw8lpS0oBzFRgXS7mGU0VT48/uGzNZHsJqks1GIbgVJ16iE6wqtWYIr6liJ
DB3Xy1I1AyeTgwwZXZu/eSN9nc6eutI75i6J8m5bMhCBlg+DSHN+mzYFHICYe79J
Kbvd/Hdlo81R9fMFFtAGfT8Da0QFsBzy/i/Ml2H1aRlu28zyC7KU+tvsVWkcEGks
IWt63G4wolmjT9BOn5iJT9UOUAxgFcSBaaImTj7AHKYb5bXwxegLArecEJkSVPUQ
jeZJVYxlYArwh2CvMhdKWLVp0YgP4AmthsjLjD/zp01634MevwZNgKKMV/XHXKwn
6Lt7VxJFEpaG6M5KnM/8klFoD8zSisA1Ccj8NKLureeD4GgI2dNxFq6tRqKo/l7k
ByAY3slncslCT2ci4NfjpABIPhahEWf9l6OT9xnSMYJUOV+JZ1VdzgE7CK1UwZud
TAG5/kamMaqtJx2Jy8DK+lKtoEyDwxbD9EtpTvkTHqSq6ZHrdDb9BvnaurlY80se
PZXrbuHN75KjVR4o+UL6x+F9PlXDB+zMe+RONBpeq7kysBjaji1tBrY9QYmN0Zg0
6yOuedKOtUK7Bkeu5qI8qKHOgJFVt5N1ixd3E/l0FYiShvcZCl73COK9igrvVmVz
KjnsZ7vibED+9uNvQWgEkhESyoxsdUF9a5tamU/EcXvq2h9z09NAnbU+Xhz8DkfO
HVUCNTSvx21jSx5d/6OwkBwWbWS/7yrqHo2K+jXNishIsyy1TeLHnsyiVbQvI404
/808rRLITfQZ1hkFj3ASn2+NtNKk7hLnVoMHreosD7gGAce5febd2O1XhRjaRSO6
6UhGy8elQ6xB3u3wi7t2ZiUS7bB6rHp6ckLCuSwmqv12w7AdJaIf/sraT4XCiqbH
PEyISSRqImCDXoVnB2Wvq1R3wxI3PbZ81J7xZDnYV7r+un0PhGEAxKx/CBuOFvVn
RaTCRLX9c6GjXcTLYW88nLl0GGWGTpQDLnsJkZr0QP5e+UyW69vhcv3DoQ2ADzfs
o4DdA63CmxsnemP1yYJC38Qz75KHPYrbIREaGrLJyKqTGQ+E3E5sMWSC7v7mEJ7B
6BLsL0Q1wxwmeHNkp9D2KdGRwPVScoM0O+2fU9J9uSprcP3p3Z7/lT4hr1ztEwJp
XZj3uLLNfzHnFew2hIWfDfO7tmITYVrNGRTTiHjmd3IJX4kpyBTsjdxvlMJMnQ0G
4dHr1xHBkjfZp+V4iDCDB76J2umBo95if8h7nCb7tqgJAltnNSc/U5Og8XsApA2Y
Rdxtkx3H7AhZUaHfqU403QFrtMEMoVMu84OSXC7c131TMAM6SxlWwv1eZpDgPH8p
1eUDEJucc/uSVXnHT9nwk2mjpS+yta2wLRWUp5VVWpn+B27D2zDeiSsnzmigaZ3a
rp1lJR0rbya0Hf9xjFGJfBgzIE7Hn8RpJwGwIVqV65Kidcvorzo3FUWdOtd8IACo
wBoonnkcPxWy9ki6EnXnq8L9eJg11Nucu+U0Ufy6xNvFFxt0qkzCe1IaGMZzx0Ae
vGhSJp+ELyPJ4Kq2L2h4J125xKWOd8r83t/9IJov5WDvepwY6aaVcU2BvwNbvW8Q
XymJVfJ2MamLZaBtaIA+QqSXP8tw4GkrkrnG2rN8aXqJR2i046owYnfq7LnM3AsY
xKxyVrJiufSJOPQ2lYuak8msrb30gtVP7e2m/7EUwF8AIPeqdvtelMnmrDAAjRFf
dhiEkUtVNTXHC77MAKv6+34XlUYoMg3p6qpAojIqN/uIqIUuKBQCgodDhhR/1RLq
rQr52bIpow0q4ludUukWQzpRF04im+xcFwu3MVJNWYqonJzV+RBlL0Rgl+VX9n8f
5H3SJCPFJyqVlcSoZz+S8bTAoY65FcPdEGOK0E76zRKNINVt1jYmiu8aOV972BQt
busLO1NqDENnWyczGTNFBgNF1271HhoKaED/7SX5mNXQHI12AjC+kL61ORMBrMNc
+X0RIHOzjSdSVghYZcQhUgLNmiytw9zXnBWUaZcWaxNmUPF1fiwyfXWCKTMCibvC
HWTMQw6KgP274fRSuGPd5poIWvWxSQkGYOpiY0mhovp+r3cKswiuSB4QOlUzZNef
gXjkr8SbM6RiOexF/RDHE+q1E4FKIyfPZEYV7cUorJUjy4/DmOhE9RrOudstcV/Y
o6QsGhrwklis2t46PSW7+9RV8PFmu25K1ZwGrTMuzeuWp7NwDNYQBlYudAUFOxXE
GNsh082EWAOQO8BZhMhwzZoNPI0R8jZnX06+sHMaR9kMvSE4mSszijBabPuiRnvM
kb7wYSlmfKqFb6iwUKLCwxBUqIgsxw6e0R5H+tr1t7mvhqRSmWXCqplPNJUIeaNA
l1Ys3jkB85ubjK5dd9h7flRZdUZNmb/NyE2po3T8Ciw1ocT+kMdo/cSjCZHd76Ie
EMuFmpTEJbg2IMRjPzwWH0kw5o744PV3VxH1sSF6gcNARNTj/tdWyG0FQH1boPbz
nEp+AR7LFACUKmTh4BB+P13e8XoGN7xGZSThx+YhoD/RXlYdls9GIh3pJ1BaOt7P
gsuFskR8d9cUMMj8OJbKqg73eDc/lK+wzc1bW9bw4CuKRGqhOuS6H9WWWl0E5HLQ
37cU0QDUDCmbrsYCp1qYajyTN0Z8x33Yc/x8wZldk2Q5f9fyqZ0cL7QpPNypqTIj
oJhLkNidRl1tMDp/8V+72+IlfhjGaBOOLUYSTq11MMf4RuMHCRqIZb+fMLgCxuah
bkIuv0zMMDZjUEtclBJ8QvPdW8cAFPJr8cqq1H8KtE/8LR4IWthY8/DimhD1RSMl
ks4t6GYAG0aWz5twk/OxwJ+zdwdeHvC1K7DZQt1OI/HRe6WxQIEfRcx+ioK+nXsu
usB0oifOaTqx+iBXjviu3TpC9up0izE3c4xG+DwyhpPwlljlPQZ5RJF1ahwqv49I
tvy9Mc+nOffnaB6kPsKYHBoMxvPZ5q2b5pmb3yLVncMmakUT+hZQG/N1r800uKUP
M2F1J/KLX+lQBvThns55CQXH2r34rlSYNz97HtD4MbC4RS5HBNYJv2T4ReDongtW
OYHBuBE9B8fLskwVOSvd1R/Exq5tH5+umTVCLbMNivBJOQi0Rj9qm8zCegvPVURp
72/5rblLwJAMCWmtbxeJ//HOe8LagQ/yJ2tBveCdbl7GjgH2N/ohHFcBHWZ91CUm
etd1r+yC8KqWqJVyM1BU3QRRKHv6oXwk5WJjCWP/HGXIH/ggIAXrJg+MYia/bKFC
7W0tExmYNwJefhZ1FHhQhtcnFpy5fnvMwm4aNm2HVYybP2wScdiHkvJ9KgWfD+w3
GpONdkAy2486mspaN6qzGGPh9zB73L4ApytqaGz3avdqeQ5iCYZS5lSG2YJc7sBx
6eQxckFP16lkvbj1VWsFLSrc+37ohETVe7iqwMmRJkPfFRRsmn+XWwE/gn+rCv6U
5YATttkbuxHQmhR2TphYkG47x2MJFF3iQiL4KZL8k3w8XU0+9PFqnyHf0SW1MBHQ
c0xHYtowSCdel72E+irDasEoT5WMuSgE/Y7mPEYODvz/Og9z+quFN/AQoXxQ3ngb
6HQEsqznhpu6ojM8YNDIxBYmGlDVXnbkTIM3nHqJZvrIsDQ5zyIkYpV2inlB8Gpb
Y7VEV7U/qQrrpDuDSkC5foIPP3YbEBR2FiWMX869A6bcFiGqZ7pjNlXsph/E7Z4t
CW2+RdIW5p7rajuelzai9YV170ywprFHKMjJaZHa2hczqTqrpY1tdmJMj0rColvG
smEQA/i+Q9zEW+c56sKgmHmYTRc7ydXiiYSyN+itKN7C7bdSlNRBWPsLisEoKusV
B1PrNdpHWQXGw2oYJFs9u/HCL7ekdZtNXZQxz57oN2VtzFb1ZA3hPVvb3BsxMJsa
Ec7vU87lzlK+R0mT7ddKas7nYm2wM1X4fxjn4PNowdnpScuV6AjXghtbuU1EKYls
gRYAj/Q2YCPnJVVbeLJ7jbGyWXyl48MZ3HnMoYcqR7PI8okG+z21exMVhFxSXGb/
ayf7Axku+KliEHjmW0EHOaa7k9oW+L6sHz2bSAlGv45kr3T+tR9W7p9FCD8GWJJM
h29tEOTe74tPCl8TqjBJqLYdofFgHaneKyvA2mZfBXPv6pXwRjF/XGYMVJCgpxkJ
gWDVxaMvo4ikK6ORtJC1bVajp1h74mgjdk2IBepzxQHX7tFUXityu5CYq1pT/khV
P0yUd1whIBZxXpkGjzcWy68b1pL8A0DJmF6EeCGtzScchBhZ9bQGmRd24PDnYFy/
eJCGiolAAqA/q0kFtczsFzpGgNS3sRlfYIpF3t9gzS+lnSU9lOfo9wyAAsemM07j
ZemWT1vvuNhSSGmYTBDZvOCqVYlRhDugf07OH0YS4yD8iUHn1BCifZuxdglRKhXl
oRTWZZNLBI7cSABDo5rrvlKEXf9ANz4pbGyhFFNPcDGC7nKD/CHALvYXmpnkCk5b
RhnNAM21lLgwLbbEQbSZgHqX+3ewyuaRgGDsnlbGRdu48wdkxKFQF14S8VzHTn9b
Z2PT3wQo8ecDjPQqMVwwikfIgSC591NRlsdvGXzTXBMlFarBWebh9pJSkT8fcUmv
E8OnLB/OiWVwLMO0r4W+/hMOsumzfh+dPmc3m7wbKyXrrS02xaqc1W+6rYckTrGL
3jay9M21qgQa2roncF6sesJ0x9BO/Kk90yFTAqjVNHucNJUWc4kFNOrBGNCNB3I8
1iPuQ016koWrSL2+lRhNm/NF7yiR39A/sLkTaZ//JWsOcc4QWgp0RWa3Qs/WxQeC
NyCIMNn2/LGt1tGV75VfC1fQ/Af8+W+0iaPkt3/rVh4t5DFPDYPsQ4Rgr4S3/uFO
lgWDiBViW1QLEByAtqlLcyMTSFjvUIGFGF7RcQhEvL2eP5tXOVVnOrMQa9B4bnET
3P1kcIKV2ITsa003ExKauLpp7qFW2DXvurhGzVYYPrGPq2hNl2s7kHSemSmiGar6
GkcOkjwNl144238lus9J6QQTBSEXISfOQGTp3kL61r8uIKng5AhjV1hyhXtXu3aY
DrBIdtCAUCrd+09MmYBJPp20tQ/DR1SOotThrGfYpYW/+PTjbtNOhuEPSySe3kii
B8RDduCYcTDCgt9aTmNSeyDV6qeEm25FHLJLm23QbyStYuc82UWn3euXLIgWH+ON
C9DccMe09g2+drtPwGn3GklKvTX6egMw7vGgPsZu4TNuS3Rla8yO4nZQM0lXrZ4L
+MrKlz/xx/icIIDG3oOoe5+IsreWCxvaYhWotatK4oiGAzZgvGhM6rYgIGEGWHQZ
vNe01Poo+u04J7y2P2Th/ILfEpF0GnT//Q/fRnBzm9lIwMCYPALSmNpCdNfVSskR
OnATM0nPOiTHdkPtolynymuLQtjTnfSjbXPZsNP+c5QxRSvgv4dzK3/omtA0XVUd
Klw7gc1tzVSjU/csXwZOhBsuD36GaDPRO+sTAbpNL1mjO4jnVABNF8WPYU/N7HFa
PjUKo/SPvVfbiSnqn7NQMYqyh7S7HM8d9S6mnSIDB5EvtMTrLJwdEHcilPNPPXXg
d8Me3QPWeGykN4u6DQHseso6LTdSPiaU6gNLbIaYBWTzEP07oynt57Tng9yNvtON
/c+DCgBpph62BMixVqI5Lbi4LRnyMC7yNUASCIlhM8ZsozVMeGsWaq6aWFk2D1tN
g0Oey4zqvHFxEXqMp+R/60+pMP8GQlRkaKZx7qcB0MBU/Dsg7DrXFtR8o/EZxWk+
R43Lpag+zEBmyy7Yl+3ktEPjTu1+1beZjlqUFLgk/8jf0/2lu1C+ofFaW+dhn7Fy
kBOPwmpp+mAU5g0dOhkTLArMCgia5iFKJQIfC2FxR6v9rTkdQ3UUWxqFKXpiloYQ
eVeCHP64nVPjgEq8jzUioMGjnGexQNOFUsthpPZpPzd4HA8/UDIQhKhlxyyHDevO
nUUxjluQQxZf8WEvzsTpyX3upwpfNdkUdISBpZ7rsUM/cr8qeMSGIt5Vru7wfM0m
fdbzvD7XKHx4UQaOFl4LC1PUCW3W0jNGJEpgbD3XzHwnrsp73VmsR2EkpijwmdOM
izYcBwvhcp7sqo33diAXzxwdamT9ljHzstVj9roIwQr7PYu8+SID1QJttNT1xLz1
FakgcJtF05NYU1MjTAkjctYvCPlSsIfyjO51u4AFvHFcFeJkJmG/CXht9sdKy619
xNX5fh3dtRJiMrDFJMnUj0Id7SSjpKLArXUH32OYQ67UMqxK9tiHo8kK+/HvBOMY
H+xgF6dH9j1hioYHR6N/kaSt9sxYyqjhS3Ek11vzmQZayEn02ynqfTKlzoi3Ujtd
TwPYgth7E/gb8R9t9Uo4QlkhTrYY6IXeRXPcvlRIP8EeE07SDcxQqiDZM2kXn9SR
CHuHEZ8r1bcC0QvKRO81k4jT3tJJ+HTeeWyGfrlX9dOllcT2kMPu+l2fB4p79OmR
Vhyljv4UPJAx6A/gf+RNyMtf/1jpl0vjMicB7VaWuyZUvqRKSWRpHR6p66ZlFl/j
PNYf2AdncLxWdU2bpk8CUhHHbkS5rVvdGNLsoggPXf/m+9WsXQl2kly3039D5PcM
rp7OYWpaGv/xErxeP3P3yuh4fbVhtJMb0SmgylxX31qSnCvrRbzv1WpxigyJ02GF
uyDtg5L8J2PACFiajie+T406iJO/hKMRc8mLDvByYzEjqzSicHgqBtBpSkZ+2Hw/
loPXDE6gdW284I1Htp168LBZHMUkycx5czXCF/k+QabpsRkyS8jYO27+KUgitGHK
Iq9/g+NZ/BZpl7wquwmetniTH8s5KjuqagKhBqIGCizQiGegkThD/CYtZTrCLMJG
tFFrWKzEAX3/6aESPMsHRWqmO3Z8oBFpEezWkWg0ICrKz5Tmqup8nwo+ba1yLjYi
Vd32vtpZUnJWA72wvnCVwoI6PsZ/NWQTeoUYAwdPf8fco7MW/NcPeA5iJGRO+ElM
zzTOytpckDoX9pFjvjK2MqSvPvFt6cQmaf6B+JaG0oy7LDFpxlPl9aGgkKB2lBgu
gZPNPlFtndL4dBqMDHMAcWzEgzknVVZOR6Ck/VoN7G4TjXuLCTBh8mBSB1VpmvW3
hVh/eOsdbwjbLAg5zx1dyOiF37aCTImEHQ89lv32JeQ+YqC3dF5JC9GaXqG4v+3J
Jc4jQPcoxRolxd5XbtVr13UVAqB13D4aCXbhwEx1GvxyL6sEvWR1bl9p3p9oMaZT
wN1YgKSraHwAVVaIEF++cFdT6q3Eum1sZw7MjEi/+EWB0cA1l/ASRffzg+yavRuh
ePw5Qlqb5xKoNAVDyeQcS0eZejtVx5A2gvFdgZrsNGhGsvHiVxj/R7AlgmmCFNTE
XM5kwotwA4azyzfGfa+8BFjUeJFpa3zyzReBqPQNvuNfLGL6C+8xEOh5HDQNgrrM
VAMnVvRo8tutKRRu2pOfh6+Zd7pQkBC5rS3Jv1jQQ+4mZJ8WtD3A2ry2vRzNdoZV
gnHtETFmp02pErxu4CyOPwbQNDVZAmkN453f/fTMV5MIhkB0MN9oyd38m5FePs0/
H0hmmYZyiVApgnZVrWSUOS55WDqmDlDZZuo4WUhf5Ic/tFi9p8hf0bJhcN6wyVux
vB3IAEEa0U0ZIG7/TOIamytf7AAmLHtu/Ipfh1sTC8JHpgCedmq9HhFLo1XiuKul
4KejjvRl6urH55FspA642WRNzx4i3lZX8zLesK+qme+w6iQAzF+VI3QnhwK+nEZ1
TUJ6JKifrhHX2GYYsCbxUDofhQ5LFn2mGNReNP/zFXIsK/SqkbKhSLxp+o/iynop
tk02sc7IXpoawJqoPUFjTbkl4wwtDzXH8uwjjTAJHfE/1cP6TPN8uq81p5Rb4i9k
AkEBTDHorJRdUMX083FtHP9vTpXiPeW0zXRKFn5ovV19l8mHeoGeI0nwNYx43W53
JY8q6PUzWxzuTJQrn4drT6Pq5SQnzdKjF0fJIGRmu2K330lOaHEW27uvfi5GiEgn
cHSnI0R6n50R9vmpxC1hVMZfe9f4CJtuE2D9twVp+tKISrYTadZNNufMlq42W1dd
1skgZc6BMbgXVy/psGwdPxiZ9lPRxxGTMJ3SVok9EnnGGtr36mpecYtSmgvTngWT
xnWYif5fT0p7W0UBl2klefBlKpVt/AMWqBrlmqmV+FmSY4cvyYfrZtHZy9vTVI2k
qzW2yD2sLzP2m3WKhXoo5erauik1mA3ByFRD3Qhktxgw6hZwGVdHFgYU3a3yy2tN
s7V/3GW0cdYO0/SP7lYo2eFw5qKeqx5t0Z/eZj6rqDFsFW+VCnXMP31sgbF61Scc
ff5Pu0isZ5swS2ZwY41SqBDSLa5FL5XiG5MNVd0lJ+f61W5v4ZJsqPgv4v2/Uxe+
QybXlIPPnu3qbPgfFI5rniyg57wREsh5aPMZHmwhi+r4fGBDdiEUbLGxY6PMn8VF
OlA8oI4ZDHn+FwsXJVQUaGSjwKUCjisGqLMTu1w1qXRL2ymltLbRhN6+vLiwcvZK
+OzoLiJGkn8W47kdOhrunFskmVTurSPSayoc1oEPQ5f6R06949oFYSRguDQkKNS4
gP4zw3STP6bjGfByqEeyzY5k8msjFNXwef8E/ls3p2rb/K31qRNZSNNWHWZwe/I8
xgLR4p0x2LJgFuj7o+RVM4Qp3jSRiZ81rP2foIH2dpNX+Metd7PXrfQwzpU7A+Mo
QPIzi+4DMpk3JzuQ3b75ikVb8EhVp9FFuosc43nsYZw/n6qcrm2PlkS9JTHepHLh
iS3YJTNu+sns4L0acH7wt/AKraRVhSCbLDFhIZ5nIiYhZWLfXF51seBn+SZtbj81
4iffTgMTS0VfV1eONtzmO2qQ/3ARtbn4ka0peOqxfHwc0BiMKtRhZ0dK6BFJAv95
I0QexJbX5xtZxQbfZUJKrpien/7vi6dbCYlkGIRyY5a9kZkFO4fBJ1yvyerpBLj8
f7btXIR/0IztmtOJW96o9bORlKaHV9ILAAm32DghLTpUQpf6fvF3cpA6cNe4x4+A
JiSkb/ssMWsMOoBM3Nc2DTaG6GhxappBJw6msoj+sPXGb9ihwTd4JCPra1BEW0YX
y4EjH6VRWa2iekfzWnOGeb7nVdK5FruaYDvjjqc3f5IEp0VS6Uv4DhIobeGxyN8i
y2+dO1qXMsBkh+vDKgo7TZGYzcJpozMgJxnAEU1Iak81Q/YjUt1PQD9E5L+5RDLy
YeumkgmNgEWKCG0NyO9Fba0JfPmU7zjvI9je0aOv8ji+rjVTbh/uylTxWiSzz+YO
P0MoTFVzGwOb/m667p8DvL8i3wm9OmvaPYb/+QD53hrxDqyW25fbSDSkJmDZeunA
YAE8g+28Bks2th03gsFkr5abjVbWm/bVW00CybtjaOtIo+Nnsb2Ij5qyPMRKR3fH
Ntb5TKxFPJ4iLT5Gec9ZZLMUz8cbdWQ/utcOGOoxBXNnF3ghhuCr3JKmAeqo+Q44
iifVbKqBU7oQP8GqYr8CcDGf4a7FPTf8wBqTEVU8riLfNnxkC/IAvX1bnGwjBfdE
wLqslMQW3nQoLS8iwB+e5D/CJlDo2WEGfqFQbIl+MTrkbeDm6DY4eOAtEJceOSZb
Wmt3wEyvOQttijZ7VUMoSaUWVUmhlZdCUX+BmEgvLkLI1/njnDpzgNvwSsNgDO1l
QQLmlb1/Ihdb5iLTCtBq2QRWbbYmPdDXLSH5o80+ZlMaQx7y/w0V3nJFBqsxnnNS
alr29EOM5HLe6HNvZ2AbL6NCL1I5okpBdn512wljya1mPtL2XzOY2DasYHNfVvrd
SFmL1DkDDxnRIq5ov3TcNPchPHLrjscc1E9aRVZZgKYC1+LETU+BKy0UnuF7LWmr
KIAdj5P5KkiZjVytHNLy5Oz7sZQjjg3/CNFcHzSrX346kqRUXd3anAtEEqtFDVRO
huhUFYPQ57RCYsIpQVgIVJ4g7f8wGGxxnpz5K4cndNasJsklqZWytWWEALkYZuYy
cMwHvP3MbgAyLajroeKyqrgCm2964mlrlZUvJ3DCQZ2tQpYAosns2b67KQ7XUKhe
ny3pPbIn7j8BijXFuuhOl/af152TAEevaJs1MKS0i5Y1oAdK4WWjbvdtgEcaQ7tk
dLPJOqfmL6JVViJs6E5vmQeKX7KPgRgxjEDd/OXaEOYGtU2YtKNCFwh+hJlSVP63
6NogCrafb+2ZaKzhuCyWsBTTOxpKCMuT9crRQGcU6glKeu63p6v6MfFio+oEGQSM
2HIeOtJnJWIvGhyrsHqAQWRah9Loeg3jK4d7YqG5ggZllXtHT9GShkEPZpZeIMB6
axnBg3V2jxjxmEdG4M2eZp731FP3a5DKkFh31WmuRE4Hwg3NUNmbUG0Z2skjUG4F
WFvtlX7hUmspX2rTO952cX7FAoOQWW15EIPfE1EUHbpwHQfW8XZgXOhn0JfENwdJ
p2HUSyxci35IxbTKjJLmvW0Df74dBqS3CoBx904j7sSiqc8ep+dZWcMmLpOW6jNJ
v3x5EngAK45rdBoEF3XLELC3LCYtZ+vUCSGPYNYjGwOdDxpw8XElg34QEQm8j+Rn
Qnw/XQ6QHMgx7UkYyFnV1KnJcnTs7sAFjqlyI6Og3hK4iDDBKE32/5V4TIN0MPxk
IXlV0raLe7JsBeFe+s4JApfteFwMP7jggE10CR0uPKX33dOuw6mflQB1LC2P/be8
vXgi06gbb6v/ZBNHsVoSuUS+cKb+ifmAk8AkBYlUeVJqtlrHQH1f+F/Gs5K1KpNz
rGv/WtuDOptpQW1apPnM3Y9gMTPnlrRIx67/25YsHT4xQsXgwYXCifw4w4WvqwxQ
/xaZBA0XF/O6br+wZvawzpEx4zDEaj28KQJtlYiM9J/rE8h1u3qkOhuu6/Pjaq+G
H+UnTWypixox2vKs+etNREcqKckJ6KFEHJgXLa4kM4ekA1u7PuKZL/bvi3hC2/Sr
KD0my7MZTmEjvo61s9V0upCJtGaUypbhv8sgKOLHdcuWtjSPt8QM3CuSUEVg1T0r
5RlF6MT3z3dhbcExLX1B6ak49b7Uvhh8mgtV0wld0tkTsFKvr7xuVPJov9CX+b/t
AC939NgLAR9lvrqd+Mx2kg6ceL0rcf6jTpk3eKzRwYUrc9E8AqMpugQPAVo/Cn/X
pPybaks47qieSTXaIpAtzsA5ih+7ZSFZ/jsTUfmR1ILvydj4LCNqfQ8sjgVxjjUD
HcP1w+wQnKfLDxxJwlTTY97EVwTHd4T0O+2lPe8aTgTcr9gv3JpkTyIWMw1B8XVi
uDLhkT7aQMibQrWJ+02sGTQvL1Q9p9nJDu2QBwzAplxiikcWGJ3IxQqpEDGL9O8c
iWb1+hX3Wdu/bt0PBLNEIZ+ZL0LyjRuW3hROxaW+HEYVNvNnmA/oFk2ujQ7lnTC8
5BVXPnCrCu4kA/tzIikMReDm6kaoLgRYPxRm8NiKxhkbsjHRS89//Jplu8jeJrbY
Rs/W6RhPCV2VCvsoNC8J0rFpTlrAyOeKCpiKF9l2awpkTC4+l/ikJzTTELNVUSVi
4ROzd58+MThjti6sZiNa2dfnEoC1UGIeYAOIOsqbZO8SUabt2l58JpiYWqs4ke1N
tkUuR/22r3/Ojtav4HPyNITBu8VJy3Ua7FauaAoMewzBxLjtTt5xqUHFaWIt3VGH
sUumQ3ZYD4tA+vAOAjXK3gyLhNrc3NQpW7FEDQAwwD2B03LZC9LciP5b5PuKC4c+
ir8rN5ZfelkNxL4e/d9Y0s7rqULutYNAge8Tg6sKh5CIcwawQF8nP8e/TH69jyO1
P3niTY5THYeXUptoQN/npuHZW1Zs43pGo6kkvAF8RAVru7+hmNcu3dE1m+9DhkJ6
ClCgC6ptQo7PnFrllzvEfduwho/TpkbHO0D+T4459ylvEtI7lITtFXhQnIFJ8MkS
04mO8IckSh+hu89dX+byGgvIsPApLz95FKkOMayoMe/LEZC4p0/Rfk3RJRQMs6Ez
SM46d5s1ifaq7ZFWPegy6RyQyijsofnJu3aArIetl6EEEtoYHa+GZWqY2/ag2aOC
ZYGGwAFJ6nrdhsplDosQeZS4CK5KKl9G28U1YIe6zLn/ikd+J7t0R3QOT9ftxmhu
iXlsd8xBXscKPV6buWwplfT79A1rTe+6EvjvG38vuXtdFIe/P0UDfI+MxsGOe0+7
0y99JXCfR/FnKtz/XUJ00M/7M18hU7EaAgCPR8M2umpEXzd1RicZdW6udOjn0B+8
6fC9wMOMsb0y/H7f6l0dsM0w460QyPfncHEIQfhzszIJ/Vpys4DsDL3XfpNb2xnK
DFgKwB/DlDxFZEGJxIP9F1SOyY4hCS+EpmekDQRZ31s3CIGRnldIgMAgfLiv2UnQ
Q+JEe3auHhNr2lLF5u1zrilT+Ivrg54rFl0A8S6IcnqVIyZpOb5VY1t7hyFIxpn0
n6vFYZypkV4zSpYDkZiYrn1+OJwizVJb6FNhZ4IuQMJZ7UZPtXppjDQXjndbRR8p
JpAaly4IJx0yuh7aaW2KpNUf/8GLA/chru9zVRvl/F4MtL0r1E+EtAWDjlZMzf8i
8/0ZhfsMbMDr4JncuBUwjHztjv6o2BSrwbqTegrTCw5G2trNFx1kdVGsg/lU1qzj
HawB5LZBx2RiuCJWi5vRkjGb6OxQAyhg4etm5x6ng7rWmf+24A2oyK3pxYR0nEd6
d23b+E9kTD6pgdJFQ0Hre4tvyvIjiZ15/cnSixdcVE/CZvE5uWF+jQHbsAXybEIX
lEg1IRgZ1nSwyO+Kbm/Iin8Vz5y8uF72MUtFXdwVNOnMNC7DeF1X8kp+VKuz4WXE
GFex59x5CU3qalrkkqvgTEXs5D6EU6mir5UUYoPOkmSgKRTPa5Hf7oXGgPHgLjc3
KEnbSjKPgOEEeFaaL69RZEUhzC85Cg10euWNRb6LM4lbJflXK91RLjTwC4228viC
Pztc00JPW2vFvijQdPNJ5QbOS4iMmfQrWganfXUi/q4pF2S8VFwSCm/mlOviCHIv
3SkD+iB8888tGuJQPLXQp7L3prh8yHw12bTATEwkgsDx+D37Qm0c4cbJ0/lM//80
QdrrmdehRDS070pC4XHaxzm0gQlRHCkpTfO7ojILgYHyjtTWJWaj/m9n1faZLTyM
ldy0smPVi8EUCdRAIoBeiqTQgQztliwfzSxBK5UPq1LkObb3gtiPvxhaaPaMPWcx
bX37i8lEJLcxbqIfDzOb9f3ZYCKiYgLZP9OkJqYlhpYhm1h4l6tNwC7gdTcjss16
fPjaNkDtVzp05g9FhqEUHl5y/MCfLArLbU9v5AUeDedVV/x9sRFWgmsAxcJ5jIsY
EB5ZOnHAj8k5kUJdbEY0dqmWmjJDgFjXM1CsmjycSdOZgKH0TRp/xWdssvjxAHzz
BlTTs3vapar+dp3w3FkAv94S+G0AG5IoL2g+7UXE1yfADs3c/mHpL2AvnyYWHcKN
S8vyRjrF2rCrIaUn3LXkE5vwTuYCR/4JSaDmez303gnquMvEn70xxFtMdE/3YbWU
mK7ePqgW7VweWGii9Pi7hSK1ceHhO66akmznUGfeqeHHbNcM6vSWwKgZN1A+w6T9
AOWBnuavLYJJMOirQ1YVGPm/B5pUwy+63Bd2sEmuCAdVRrZrKPOBqhsCSg7uRvrE
8L27BkcurdrUPOCoYxYnF3e1/tk8tERTKr0ibpXiAbG22eEQKVAAVUj4goguSpku
pd9ZiOA8XQbztnFxgnpjVi7AHfl3Wi5ciV9t07/1uDvGMQCv9uk8bmzvzhMNVGP1
Eqyp5eLFu7tEcVuVj1YcDz3MBV3g4StA+kWC1YhSJeMA2h+CBbyIPtCINA+p9wks
RIVlMDApQxpio8BAt848EctV6hxcUEJcEEJjhpiUJIl/cx0F3L5aFnr5e5K0qqT/
jKdR4m7/0reddotFUWQVIxm40q7FcYGYeD7QUaECXjx+R4SShbLQNsJ1Qe3VjoFX
ZGplsj6iBG2OUxP5PDA7noAZjYbO6vdcn4EcDLX0SFvtUI0Eajd7G7C/31hDRTHp
48CVXSfTpSRlVvaMOgq1kWUgSA39LdrbtxetFIWUfyxvA8Mx7G4+x4o7PTUlb1fV
vbiB1frJwLHeO0GH2u7VgrkwI0D6VbMkAC6reL0oMRxJ9QyokSD+5cllAqA0UGHl
boxWGKON+ifFyAhP+/g9HghsiU/JRevrUQcMxSBA2ITNo6F5gq/OSzlxOmG7nBT5
KvRMcDmwMP4IT59EZfMKrKoJWCIj+mFL2Nq9CdbjxxBKIZ8VsbFVzLOyFALYpP2U
VZqlWmo8A/19/W0vKTVD0JfUJf2xL1BzWCx0xh1OPTH9Bjo9w2SnmktmW38/N4TH
YxSIwwe6PfN4LmZ5KNzhV+nbG9P9y7CNU/3m8lOEjv/MzHJHod5axJnpyruAJZz4
zqhMbyDhcoeKVW8lxhXGjepPGKNc+Oohu+/hirOBvy8Z7y8Xlce5mBGs6iKrGH4F
1aeQZ6IT/7QcbUW7uWFrjmN2UkCK1A6e5gocvQ+lqjjV0eLMczc0vPAvmarK9hs0
pgZXlFIPJfcxi6tC+7mc0RF2ecGBC3Wdw7GoOpihTN/aGfI2TRiwzZBLDEQUSobe
rhL1IBuxsVUqEONgF8CWztxMlJ7CtnE7mC7YlaVQR+h35Ekx3cLL1IK8tu4Gcd8T
+weLvYU/mAV/OAhF+TOE2duxiYTJqm38+hgKGHCtpb/6FhLhiVmEkZE7teRsABTu
ztPzfgoIpYOVM86ofT8pZOyiq/xM0zXOU9aKEGVJkTA9ryUYmDpmQiRbVshKZpte
0yFsa5Bk3JGmGwt+vo50schsMCzybZ9YBE8yCbrZzj7mFIr9YOnTrwmRc2x25aY0
NQbAsxAsZo/wW4PdohZ8xn1gHeKeGBr6o9dj7bRm6+wK0lT9mRoiF3ZZW/8x9EAb
u36qIMc9PJRwVH9Lt+Xi9zgz6q2rbZZO0C1R7rkRVTuTr2Q/G/9P1SCeM/OvTVIE
F+JWbSRx/LCFNLhCgJ9lMGuY0U6DUFpgdIitsq1bMRF6g6XPmNMImwIiYmHEQbVa
dS002eZM2WA8qsJ/fIKpuIlugZpHkGIsORRfO/zdy9H/WoDFgPEKvRsV8TnyCwLd
rEPYqNVathuug0ZpE+r6tTGeY2O1fkWJfghHcYX6g7aPkx72dL7r6q+h1hieLf1B
cJWHZxtXRkwachlFYGKk8LnQyYNGGSVFGPKnoxe6zvKiFnPk3rioLwew9UlK1bWa
lol0coxdr9HQq+yg1CmQTTxp+bdbTzDLSMMdCwtDSDT9Tjhnf42tRm+ChtBnY+IO
lnjeLdFl7gatHGrCDArkyDk7sTUXSfDWXCdH4dKwagRCms/TMT5HAKeOFN1QCBji
pqtkM8c0cpZ7ENcn06qYxXKRt8EgB4+bUhZ1+p43/cZbngsm+ZrtKfy9W/mk05Mh
5A9bRZwn8jD9G5yJzoWq8hzGnzjPkNw+es4hq6ewUIvfns8WRLRhyUUULvZudOJM
RmW1EAy/peIX7ZNzMma01zHOg4KiuIWhcMLICoXKAx+c6PS/913roxO//4wmjIb/
P6/sM433Gr+2avmGxby0s5QiDm0F0LVPyVuFnkQDikYsY1fmUw1fa++M+B9gzBK7
a4ltwFoxOxyVo2duCPJcAF0EHdyfuAGZN+VveI6ST9Dw2lvUFagZFOFdrUV1JvdH
PIff7um/zBMeSaTTQB63LXTPO/2T9M0Ym/LLjRI4+9NiENrRyjaxFRf1QadtQglx
1LOgpZVQfTlD6o1A3MJD/eXeGzl/EnP5fUOoH9TZIU86b0QWtZp/iOKrartdyiTx
wMC1HnSmCbvth//mO7eztwldpZvUFlw0bmP9uFY/CHI09Ka8LZGigRVHZKHFydXj
sn4mQ6QoPTD/Mfo5Ql1TByaki5QH96nxRng2iGDEA+0v6uGBp5zdV5kmzSOXnqQR
2eaReOr5yzymXsx/hkjw6VYeKvZZksn5trjc3RcbY5nWcPdfWDsPwKXtRHcoppV1
fPOA2aKKn4duuaShhL5wq7EU2G/ln8FN8tKBYTsrmGK7zJmOSfOJYVqy10rT9NSX
OXAXJfipWpWAmJLSsnsfVXf95s1F8dQGDTR7NRkRa6TqNmrwebggsgUH1Ibslflx
tDlP35X+L5QjxsRtbQXjnLDdJ4c4O0cIBVTCIZMSnskGPqUWanAZWHeC/dWuwUMC
/V1DdUsRcIKrIw3zXTCAVnrTVNTb/DtrmWbywNTOXWjk92vNjcXPrLngtK0M95Xb
5ZJJ4CwG7r+D4J7bTO+w8p1X7KFisRFud22jthqRr76KvTg72F0RGjUXMW+4W7q1
TYJ04AQRH49UbFOnNvKujd2+RCgDGOFXPUqHF82T7Lz8+9hMeH7gKJTIvJraqiN1
eaaOP1psu/lIQydB23kS4iwD4/4jBHjdpB8iS3bGgCrM0ZCL/cnLyXt9J7HN5NC9
egu4I0Qrn+vYEvl49DqetC39iZBWMtw6Otju2Gmkn8xc2mDoGsEvB7F/jMYUUcw2
gceOgXYd63RaWvd11SX9pHTJhXF1iabrAL2C2kMq8t5bh4U0i5XWaccSBsBQVES3
y6kb1mRVo7JTC7nBX8pDxeZe85j8t7UskCi2hYEVAHHWfN7xei3NxxUUXn1OGtVV
V4VpLtBJy2sLfmCU9kEI/Wvzip+mLPBabSySTV/eUMejhDhS1F6/bjVPHyTe8+fU
s3u74PHAQ3B5FSWcih1dp8rG1/uq9AZKNG38bQdmZcqubSNX9CZqHfaYv6PSivjt
qMzOfuMjCxH7ylox67DsU9jVXwMziWfpvOAJmQOrvfdFPvZrV5tMWBM86MONTJeL
YkOOv123lNPaAWoBmpQJmC/YYbBsMTuS6lL3MmBQYDLJKp/zl5MtDlSPWbTFZPuf
OyrAwpLewlOkr1uHG7z69H/gRZTfgZBHQ289H/efPp4bSyqi3aYwhyT+OJuImVua
fZx9KLFj90JPEZfLKuPFq6Fxp++VqcqZgh779ATv+i5ug3gwG7ZqZw8kvi4mboGF
3N1g1ZUIFnE5pDcJty21NHmLM3uC7mSksjMfdf1y34vNejxXJBGWVUPlTSYVo7qG
V8IfWAi5HMW175ISMRkgdFMEk1xC5HtkDLRNPqjTILmFLDq3/l6t3cf3EtZSES2K
D6V3VJfEK2RloxoJsWdwZI+7OJVgwu4E8Evdm71pxgrQTlCN0hGJG1eF94JPASf2
8ZdlZvlW6mFDFsytCakykgjVXfj5hvmk+vq639dedJoDEW1QQKhLxhVz4B6eWJgB
X9uFMuHoqOV5yDIC+E5Uq7AsYtjmqvOU5Tp5C7RdOkRsJS3OEoUbs5yGmqD5vp75
CKCvYa+liiGzy01UjkI0nM0aQGlPbZvle4om+ZfP7UTd5EcXlfrZi9fKern3bj+d
KAOloCZoRvux3E580Ggi32dqDVv7Svqw1k5DBNVE6Qrt83Tila9n4HkHLtDF6lkr
BZzu1mW7Gc6frPKLA8T5iUDXhY2RcmB8D1MgnxXkK6FD/skD7ORbBPTbVpIbU921
SXrVi4Akj8hgxxwZkcwbZvguRHcWAmICxhQXJGtkUvFGjIr5wg4wHqOlcMoT/daK
cciF9eHZGpxxPzgY7nDOaWtnw2VxtUdymqeL/W4M/5d6nVhwETJF1Gtt9HjY6Igi
rdDaFCt2GnhTzYR4qTGGkyf1uEw9pj04mXcWxVV2bFyPCfGN3X6TAk/pvMkF+xxJ
yq8JW8cIu4VyQ7F26iMEQTemXkkVXyt4GqZFb+PdkRzZkwjYGG/DGfDqTk/AWSQx
pgneqvEbO/u36mO+hj458i/0FYYFCHD4XsWaSHwUJfEru8R6pNgu6l7d+07aJKRh
byOcHwfyf7nmdmO257KjHQcvd8xpRKojOzhi2pTLUp/+zBHLS4HGLTTHYCG7Pofy
5DiZ+4R6/w+ZLSsv9ts6hoGn8xPWhsjpDLTTMYs9e6IyF/EZGORFokyM+UUvD1mN
zzE0aoLKZfkDYJWhdW2RCYhOdSgXSyCQ36qICnv567a8xsjU9CVyoCXiL3qBR+2X
LHeL37LRB18kHvGwASQxJXVwB5FY0tzVXyb7QVtdrM4mwPibmlzzyLWlQviLUOiq
5kPOqq7ImNl0SJZAok1OzUjzvX9W2qBE+tbSK9Y5i4jPfMOU5U/x1LWSkYOk4N4E
mQb4kf8qcYTMiJbSo65aiaqCjDfEb4kaZA6XVmgyMzjdDhoM7MDJtSvedmCv092N
XGcnYGovwhIIlqokxlk5bUnpPDe9wKa0/GLw+GcuQz/ODRQSKSwDTCgpjYoMjrP6
sfa8xnxyoIkkE6w4DgVIl0FwsXYlNxyb2FNfv77CM/xBDX9BSMAKFlTS+cdHjF5w
TsmYywJlo3KpXZFNleV3l8XuWw3reyxFiU54jxafPY9xQBaPsOCF10gEQgxoU11k
IVd4n7IS4uT7nT5nyh/TZNCUrRwKUyzJi8gUAL/nhP6ZQHJQt+UpuMPN5HSb0ShY
hPZIzQC+YjL4HDfoA74aZzWUSNYsM6+0EVcjSgAXbZTTov1sQwCd1EEP2bmz2WqQ
16DKQvslxZB/JNc0GjRSNZez7X5sdP/dqttd7mH/dQGBkKo4NtvJGQJaa/TnaQqH
gg8vr8xsEV8Ovv3wsJLhlQ0A7O0TTmYTPCZCBmdFBm2LvGeZi64Z2I9Yc7NpRwwe
RxFf0VsfZurHCf5qXMjWzU8dPHvsqMNLvDDGlJSqBdWtsd6npAf7Z9DlWkZow2Kj
64hyAEjQpiCmNsPSYzhI3czuIZQKFPDqadfYUz4qt4ggQz47HPAAfCao2hV0Y7nh
6qIFeL6BeA5ACN7wdYttBYZr59cbBPy64/0raXu2q3LJhKVpjJeRfowT02hSM+5Z
YXQ8LsJwtJe4kxVaBST+niaVc1cA1v2+LSNA7MkTtsdtMV2efXLV0Z+ojaYnrOJ3
hUT1pYAvF7I4nLtG/9ksmgg5UpxDrdtcqUR1pmTBSFuUJZIIdZ5ivG1fCpQGdHoH
nMaIa/rdyWUGqRVpDygpWmTpedJCk1X8FNGqwG9vIwu6dqNLMevQSqWZ5DJ5dFS4
3o8q2YFALDYFKnG5nv48dRUPj34jY9CbD6zYKs4l6PLxCrtHc2eaAcyte1ym9VM5
AoC4Hk1lLCImGQE0m/U8xacelLoMOkLP4WXq0oC3igBZCd4cO2aH2w3piUZyzU5v
0qvgM5ey7syuMRkMmbLkE8MIeZ3gCPO/88HcNR3gSW8468FxYw/4JmcvMHoXxI8I
TSFf+QqsOVCtejAtKzu7d7yvTpsXhF4uHDh7i3QVFxByfAvmHGOy+fdFWnQifwu4
VearJVRp3Ce76ACZXdjf1ywOj6BAxxk14m9+Y/Fs6JEA8KtFr0jSYPnLCOAisC1W
5EEyPWb93KbuV02slg40rd2cF4yMlsgcNhdUpbpX1LJHW4AZ7Y639Rl5VjiyYbPZ
CDv9skgkNlGhRLmwdxT1pbWYJrZ+fSqlPZkypCwSNsxPp6jIxKoFxHFuAzBIQVaf
1mseDY+INGacmoU6EsVfUlULTTHbD1OPI5oA88k1452zQPeoizLTxq+eGAgEGW0j
jGu3uWUXYAO0U7Lj8M4MVo/k3VE6ROtS7qQBxU++jnHBM6xLJJ/LaUvrXONIYBlW
M/aWvR9FVVAn1/oDbTdwwZUQoJKln0q80vkCSdinrT1Xww1q/G00VVetQCN/nOMK
1G598xV3oEj+M4BxytBc8kd1+jg2CkViQTDozqmtGZmR4lqO0Cdv2e3OncCiX2mJ
JrXFY9m+Ocw9TfJc/OWT7Vj0h2HK8nnV+Qz9Fu5RPhMij9Et0+49EYswd92hwCN4
KcLKbp5VF8C8+/dW3696enKpjrsmx+UBVzu/7mLzbzBdAH5T/x0qc/3lXuHtwtnw
Cbhl9dSnfzP+nhBXv001F8l6zTeblkBOPTyZUl8eNQLvhTX0LJY6Q9BVkUKeT0G+
OiyHH5WC9J+eAPpMMmPKq4Qe6olr7VnkeZ0bixmyno2BwzrlHsYfo6F06CZZtsSr
nmZ2/nEXxkie20k6d2h7Q/mVcfuvvptz3BlJYFpJNaM4SLXYLPKIpHPRnjI03edd
iM+I0dND1h5vvGFpZxPMJm4xZrNg4N/vSwv8LneYmQM43zz5gWFuQznoZPAkIIeP
X36FUbdS6qWLrdvCMg1Kue9U9LFnz1wKj/Vj/C1HUUwfUvOYXjHvv+h4kub3V5fP
BxeEMPMYmXy5gXGNTMAqfUfu+og/MZk0/5qRI634GfzMC0JIy0v1n4a+Yq102aXT
jh/gfmIgYIIAtpf2Cv0kuW+WC3ZhAydOhmRYWFMZIhXVjVzTwfMP8glWzYXh00+T
H5YJgdjTtHnEcibrt31BM9aMdoVzYoYaphE13dK2TOmF7xamgWdQGBG0tUk9Uznl
e022BdEujpb7JX+LlIXWFfQHrpF1M6mg5HJRnXuK5bOCNYKvRQtu/GOVBwlU1ud5
F6O7tSmfCl+3BbVvo/t5XtrZHsmMb6Um6prcUj6rcF2jwTta1L9moOy6ozak7X9Q
6RSQuAUsQ1S7qk+olZmC5HINHJ26rtFPyNnv6JOp/E84SylOSt4166WHG514MLNf
ApvpCmtLg0JoeVsO9RIx63i2OJPHY6OAT41rOzAMDnA4NbVG+2/GoeswdNIlbg2J
hOqc7Mi1xrn84vmihoovqmUM048HZlKEztfIS6MMCGlXScRx2Fosi8fsgS6mb4Ko
xfKR7OcS0I6UwftBc2gCJWJgvFQzZGaYNXgq4pE218tDc0DSEOqCQm5mzufkD+F1
oWGFJ55k+YrmTMyWxNJkjIjAfWlG/rhJNcShZgJzr+bzA3KWIKviEFpgHeDmDKi+
NFgj7TVslsd6aNAaeA061SjAWA8qcDlVXCOdztrOr8FG4BThizI09NoutZL4f6AW
6QCA4kQ41LEJSrGVV3iBfL47wQi4zPjf1w58gx5iQZZ8Tnols2orKiB7nVh0ux/V
cClCmeySfwIDIglmy+Maucl4c9WH5FXeEeSrKwSGNlmejvPkiSgDSakONT03FfIl
xj50fnz39F16lemIZX+/jRYurCU0ftOr1trplTO+Lw/FPQYXhSNVTJ83gRzDJGDu
MLNzMugcAyYUobi9LJWq+eiHtou3dNTpkG0PC6kocQAo/YAPWX4I1fo+rPNVIywe
BA3+mabi8B3HfzI6M/ua7b42UXOZgrsVFO3E7VlVPx5iv/WpD9ifu+TsOvYOF/RX
ObKFTESH0UBtD4Zq18j3DdWy6/h3L3o77r2Mv0SZIKjPF5Thi3lA/YpB86eqZKKb
oPenPsIP3HyLN3m0ycFUIvAY/Lrf9ObYnCzpRIR2Bm+FOFjBMJ0yi0JocqC8VwF+
piSP0d8i9b+7+XJnA4T6R4cXMmJ9vJK0dVSAoarpb+yPu3qD2Wh7cHVNdrAy6X+h
jNQrb+T1uaUIDU8nf+wbitlicXBozz2woI1COTVtGtJUvkxnYkS5PEsbxIm0l4Id
zA/jesT5JS2CXhXtfmpyvjJuRUTUZU87NIfnVXJOKf7wIp2sboswSeNF5NCs0yzp
VDPzskyifVlIbYuUcyP8LJWE/45PBpqACrFPT7NcYzCegi/ZY+u3d7qEZmfeQvq6
zplaVB7+WUua93zheY+eYlA1N3LW4BDNIZpvtkAnc5+CrqErdIPCZSMlsKwo63FU
K7TtpLzns2TPAtP7TSc4haoVO63fFbk7LZCkenf9JrxD7fIUbf5EsvUqQctuSWSV
1dmtNxL2GPgxMn0oPanKYHz2F+XKAlIXQSpNFwLcFIrWgbLRCbCrHTF1fPQWDolM
jykNCcrui+B09kXDD6saDuGCbpUkhXNc7tj23BhYW9Qth2NuyXs5r5uSUxSouRUv
6ET4eJNgFL2+wZaF8j4R2nmnvgiotGNcNKNPMw1Po60ELRJboftA/vZw+QFUuylP
fY/b7470PCGGOqr0ohsdT6pwM2LB3gKiJ6agKt5L70Yq93TH7YdGEGstFoOttj6z
kr8sKXcLL2FBeWhbgk4rc6rTmTJqvM9ar2ooHp1rjoAiwox5n2FDF5v21wI44rLE
6+XfWnkSbNFwWAdTRwchMa2fBW99xKkn+QDNdBbseLZVvXqTlGlNgO4rhPmGoCI/
44qRmgZWiX50B+Stgg+328FFAxJ+2hdCnhPlK96iqX+LIQgFtvVsVRM5oo6xTWA3
VVymi1MUvCkR1v4I+rlnE+B3vVMVWXzfx9x5ZazBhyU7PeW+xA2w0r/a0DDmaoyX
Knat0iUjcFO5QCEXtJn2DfMbgAyUxEGUy2jD0VqX5Dqn4hGx7NvXTr9heKEDESip
26IqmkYyuJ4YACyK4iZlWBkd7hXT1+2byDTaTk+bATt08UxVQOh5SoEm0pCxM29V
1xijjYkgU9DviFpvxzeFNsTN+ft1BhiMHH7PwvVR/iOv/8tvqZGdJ4n53JQtmH5i
N71blkZ/LYv/ngPo3Pfsyu+gXmOKXa9wI70JvvIvlCDvXHP3a9WtGMuBwb56f3P1
1S0mXjvUdZh0FbQ41y4NhJcXqRAyfDJHKamIU13U9nzQDzHBlPCbCbp/fazJevoi
lW8FAPaTtGhorzjdH3YQrW21dxC8FduYvq2dKesvT65i0zBBuNF2efiCGLlkY4D7
qo/ZknumybDYXiGAkE5iRTYEHFSglDrG7Mj99MHqcS4w4hlC2zpQd6y+0OIqvsG3
dWKSs9r2BonUNGKIBTP4WlsbcqCFIQwV2O+yGp1dmbawSGLxjSNeuNwOeV3+P7+g
O2j5rTVij61by656LXB4yfKGl7SXOseiG8c6yyBjfiRFkaHFNcrf/WR71orYIH51
hS2jYN5/BW6hpd1GmnZlYde8d8quAERbk2KPY3OM5lr30njDarY6Ipj43ajUFPnn
wVJidajSyFqITX2/GsGGKwLvwrrw1pXeVe0c51B9bsa9e5plS35JplAQNOx82spa
f9hOkVydxAqtIYJfFBVm+XaTqLW42XU8fYUtib20izBuQHpoto5K0IyYh4mtFOZD
7FlHl17BoiiwzEtteLY0Kn53SQiTmd6yu3GkYYxYhjqO/czQECA2fMEHNQzSbjck
nAT6RXX2amzMrd+k5aMO/nw8FnLre2zBSk2RJxeqO8frO5oUoXr/fyqe72Nk7SEw
IbsfmbMqhEvbNiXjZZry1bB9Clrvs4SuCE+iiW3d3AsanO12/jvj9+0eFFA1SIO1
mdXxm/9/S82Brti+atwdpxOBgZ6gCBPYKjUW2BXcdFmrIt1T16HIRTAf01XQJy7I
ZbWWZh8zZBREwya/zVi27fxzxAtzmCsnN0T6J03r4oPFTqdMtPP/fAQn7Nhnp8kM
m7d8ChkYxdnep8pKXMLPd6DVCisVsHpmY3PiD842V4pG+P0P8jVKzHpfC4/Rb4aq
UcuWp9I3nhwE2G9G+STjgvuEEHgBDrEoCE2ipql954iZuB+tTJc4arB75jc1DO1u
g1gquzu9rQbA7I2/F2wKVC3YkRBy5SQ31x5eFhmQsR4kiTU7KILcBUbvuj5ifG1x
/40GpLJIf1T06BID7ZJE4gTmm0q6Gd7KvdYp4cu/jdN//peCvEY1fs/Ocp/YgIKq
LN5vhXbguCSHfIDPvBFEtHfOt2lMBxT68cWHmfnZ5EuF53xxlftjVXtQHY8jyMxt
lNUvpl0h+GWFZ+34BEXu7XAd8HEJyTqGxu8slzetRFNjmse6+8HJ6DWpUjMOEWgW
B8mjD3B02BwmZsxcV2hGp8O+dWVtO84DBO4/BZe+6UQUBvTSA7E866rxtNuvrHQE
+1N+f305oLWR91qplJ8ORKIsOBY1yCeZ2rdNuZqmdsZqZMCrli4QN+hTlF8PLQw1
GIGYdoqNfYkR2j06kUhBe3SNRPQajiIlADNjfu7wGRGSWroDkNERrd9l9fXskqJR
w+pH3QgIg2WdwJ0U1pT7gRgNstJNYHsWCd9qIuf5WOV3lspXxm9GpmHlNHb7yDXh
ZhEYxEhAb2Hq4R4ilYUgW/IZmhL/iNI4dRMwMpqlDWjdXGmr9uSyBJnndeISkw7Z
0s7VG8LxuhKL7tIWHHYo0IISYw9qBehJ5uG1Gh0G/dvZytfTkeGxcafXcSvZ/Wge
PBR45YlV7fj8T0faLaakBYOpdhtFyiuRw+U07Zl9Ur0CWAq22rrJvwqdcvTdfkYK
/UwgwhG8GhuNl1PK90oY4wG28qm9rRor3kYdfT1ABSRzz72Y9bnW/fSiayhqdfAk
oCqPdazlV8rroWW495zKRuART3wxLExDN8nl7Vn7QzOhv41U+BfMlQjKwGRkaMUI
u6YzkY9DqPqFnDDSZLpKAeBXkCh8xO2PR/io/WO25ktpU8hrd12lhYOQt3cWH6hI
GO59Cs3yEkXv5OyMrPeMcLx+IhswMTr3wajNeAHltiNo3rOmniosCl/mW4jVDuuB
r2DbG9Mncye4rjBSTDjPYuXdFk9PFxaI8/qsJ9k2nBY8T6iKEP9vj2x4+1hPG3Qs
x9tT00xjFgmvxE1nLihloRsO2FDklJiBFJeFfTlvKvzUkrPzJE5g20JEZoGeY4e7
Uowxg+Q2+xjlPGfztjzYNUdRRrGa7o/fs23KbfdOJioqy/eMKgKWvUyzN6CzteOg
uhJ1ZekFO9+V2P7DARrOUGEhAQF4EaIC/v98zIqQGLlN4B45TtctO20oYmdEYwWZ
50h81vvd3fDun+RvbN6eqgxQDMbETr+guUOympr/MriDitU3tgTFO7qpBIS+sewx
dRn2V9G80irStHlD8aAvnUoPWXA5RmNpwaUW4iY/X9q6Z5M/J8BtLm4N58BpwpzG
rv/7nUzXJLrUDDGsZamlKp+Gissoy17KUOuGuUlqwCzB7MZCC+/j87C9R7XBlsQy
+cjgdcw7qQ0DFtV/it5vAUuF7hQ7ebnGQRjZKU2D+Z89b0ytPAPaC3Uoov5kllrL
tvOQAPCS/lxDNqYVKFIGy+gmdrV1V0U9YzCHwfj49jUnOqchiBAGkQJlSM7ihPHG
FpMBp9UzVVAeE8qlWmy7JG06XxhcbnYyIuwrri9DBSSQJ0UUvDUGoM1QF0ONvLS/
BpJiKZLcVkh460YKhv2H8oMLVAvGbcgffR8xmwe3trA95Ta01Kbh6IeM1mVoUvAg
Fu2/qyH436UTTAgqVV7j5UVBOX1gF3P4grsVvUxHJBglHqobLmH80OAn9bPlRZbH
84pStg211Mlr+gB8G8FUd/9JwT3yYiobgcM+0qs2AlOEbiBbAHNZSrx+Va3RLTaR
NuIAWWrML+z/dGY+IZTkBQV8hPCAJwnCqk2EZudUhPDtoMkOBIWa6Au8x7Y9eQ2w
sjjd5fzLcFxFbXYZx1Q6ztisyUbsIhUBx87CmWmZOUydafC10nDwcaxFz8Ckj5xp
omDH2Z2XCtTM1I6cT2AFvUIRRiv3ax7PkZzPDAAK9lvzYZwTmDOrBW8Z1x61NPaR
Al3jHRbv0U7Y53ZWplpWXSfBZ1AJ6E7o1Zf+/duc9QWLGP5mDev0DlwyZwf3Y8Xo
glt8lgjauS3BaEEAD5r3nLVoeWkMctgQswoH7A1X53ZqZEmMqF2w5CpUKudz38yC
NDgDdn/J7m/gRyJsi8j0kQ5RGpLQqDGo+zs3Ulp4Gtfyeio5D3Ne4l2i89pjw4I6
4EequstuIHy3+Vou9cqcZOLFooqaIiFwM7pl5fbedgl901celB60W5I9Ic4eAKX/
W6s90ToEQORe7WFS+64Pq6An0cb4eRLASPoChbg/36MtHdJ3StXTBt07ilF2czOW
nXLizNiGZJ68pwnx1AGgb4YtTAn7AqCHE+fHXd50qcAIhCCME7MrUF/sEM1XGRJe
uy67cu3AP2qABx226RuNvV2K+ljDhmkI0y33IS2NX3mlf+ne0cVnEALEEAA+QoU9
aDzW/dlpZbVYUTAzUJl/vJbnVMmiukMW9qWBcyy+FX/0PDvNh6g8jL9CZHkySXzb
QxLno1uXJjWuGrFz0mSrwgIvXHHnesqpH4TwBBO4NYG4eKnb9nTAgg/2qm7laMXg
QHpv588pHwRB/4ce7ErL/eTcIZXh6E8oqeJScsku869l0jBhSBbhbOwtl8xLV8pv
wSZoQdTbhZNHGU7jMy09x32JbQfH15vA1ak/W285o2NytodSK+erBVPtgKHl+E6W
Wx0c0NvVxI1u5LDL7Zu47LQEifzCQHVEMi5aP9YwQ7CEf6yZRL7dJi3CfsscETWt
vERZyv/Mz5niKESHIydwq4WwJcKmHu9cjt5NcYfTVcxSNJOYjtbBjAFxBeVc1R1Q
JRiwQinJGrmKGcvFnyLgQJdn6CC8620BGvmzU94Dk5MgAcOmOxNk027lyjVzR9AC
Qk+9yQV3SW5xbDgjwg+ZKqibOnW25AUnGEk8A7NTgjCJJ6VI5n3ul9jd/axr0shs
C+AmrVHR8QjQ58qlZAnvz9FHfJa8KM3GwhTO2lZpcrCweOgX5+vzhCnHbqrPWJnl
U5WEUOTW6EIOMFUXz6zvislla65ZKV3DT24211Yf8ksLVMiovib+jSFFTvnx/beJ
pH1s9mmWH6ipmKatmBHkNLWstvR+NTrrUxaHo8ZGmP9BhhiJX6NwnSWpht+ow0oY
NHS5mBRrIkYArAAPOWxRPT63KLKtgO5dC5YlkbyZGWKFuJtnH/3BBSwakNb0HlEz
JCSn2iM7T3k8hIM6iMfpJk7zXm97mKIfZyyXC9na6qYauAfpTCHgBxW2MdHBZI7Q
kjJuv1rCgcxBVwgnVM8QFuJ9FYcIcmxJEIRprIIZ63TJ4X8fSQxOB3roEBdbPbDF
R1MHyHXaHKCvYVa4720Sw+Of6wogj3Ix081OPhToDTYehjqY3QLpBaK2+o4WRXqV
hERDYCULhscFXgEqhHzvth/JE5PGTmY2XEhoo5lAkSm8OoSuSk4fKlEVVC1Avu6+
HpZrHCZpzbSBg4dKiWIETZHoWzX0ry6Da5T6deDGAx5/NiKYQkKf2HSAU1HdYCUO
QIoQvjGPWt2aXFLrfOsNIK8y24uzpSApVGDQRlHS3PwJECIkLGGN654BmbUx61nI
1wsND0RVSyXnq24+GMtY7sEmpME8Lz0kInFlOgVaRusCMt7/n+5xZVJ62X+bz+OK
YGTDOV49d0Vt2arFnvjpi5c8707InPHupdTdx9ArfKo/lAZIcc4CAB/g1rnvLnPQ
xQB21BbPMzRP7bFAYTl+Cn+xm4AYcv7LvY1w0ModFeEUG3pZU8OA5vYiCaQ6ZXjl
IA97nPgXcMA6nzwHkBlogALwW9Z+wObxosYeFCmgKna2KgBnzwjeO1vpeoYlkfQB
lCAMJTVkvNzt+eun5bANKfWjtdJPJ0BwkO3VQ7WvyuaEMvw9U4sZAmxLMJfpi2Iu
us9fgaAU7HTo6WapfNWmvUHG0HBrjL767Cd7cQJr+OJW3i74wKILCNcVIeRk/19Q
gVjsycxQQhZemxeGtjLFv6JAGR+V4r8pVb6Vdl8FPth4iRxmMIsQJ+SZeHaxuUd1
S4prslgcsdW7HrNvqnXy+Tt2pWNWVQPanKHEWStkveAE+zXq1Q711XBVa6HU4ZEE
Nd/rj+31TKcUcds/YtPvsgR3VFJt2ZEdz5hkvthEbK1IJqXVwihnZMFWNsc9JZKV
uH5aukPuEw1TdWJ/n0U63ShWzOAbc3ft6tPEf3CsAeDO+FK8w9XnD5CEvHJzkntN
5H//vqKVxgpILlSEiKfqR6LcFOlG4s9/tO+YMqMLXRwxyq0x0frFMIzqN319PAMA
BrcCj5H+ldWWW7JvGRmmDuEa8u2Oy2S1D1Quhu61IBymMmqwFQbGTC8ARYoNg81s
gfGGaTMxsIcPmrRsY+C/796kD9vcc2ze4Mcrk727tyPnFTb1BDYQMsmjWIECBmBh
bobfHp8bHo9JHCMar4rNLfY5d5hdEcjA9jzPUYwfKK80FWXB86PXZd2rmyPDKKCm
6EyqlI5P41AXzRdhHvLdYy1fJUyFZW+c/K7P0hoSWkjMkLY/M3yWlBklhZ64cf9W
/eVPzvxCAVAC9LxOIaEGiVfNT4T8FV9MDgGOTNk8oGdvZ2DmggS8f99RfEaHlyK/
498lmKArvW/5ZI752KFQyDvrE/9LUGxDVqtci7xDu+inHwAF/XFDwcMLakqBo8jN
MKEdMOIQUV/BoN2GI1FEtoe2B6VEUvpapZtUxTyulWlsCVUIGSnRZfcF+RrvSYdS
RPy9Yb1k9Jq7gTrGveMQGbJr5DXcZaZ7xY8w3COsd3jma2hylrlTq09YW+ooUM5b
f4E9QzUn6VxrUCnpPK9YvNwQOPMp3lwqcqaoEH4XY5Oxiq1HppyUXndKz0/0I5YZ
c+K2z/q+R7PKtcEQVvGSF3NYbJD4IHPSei1G2UUktsdvvzA0U/Pokg/NxpTMi5II
+IEfFNgrcmZYR7U8LP2LKXhnSM3uzUBOoCcLIsRa3QdLH16V8LDM/r8q+80Ad+S+
KerZioyIROV4Wr8R1njUnND2VsN2Ji+e99YkynH5qyEveGujT/bhXEcCvHk7XF2D
pYmSUDGoJ2zXgW3Zcv2M9pUJCXY50sDiTquK9ATt51TSCOHUSOWd7rh1/mSGFTJ0
rfmBrDGwQ0W1tcYgCJnWyXbG2Q7Rqy5jfedY/O0smbMvKZGZwDn1xcdvfHKnxPIx
vcBpj48AXmngimr0qnTlv9sAUpznkcOYPzqKFmJcM/KsCbR9wSG94JX0EyNGJv5y
7+rHMw3suXPOO4lA+yLFtGRupP/YIlr3QWbwAplCI+P+nAAC2BAuR7I38KxxPYkr
qj4iq7+IeZgpvmIo0qi1liCBLxHF3ccS8FiFwpkc/pIGa9BTZsQyRPgYr0e170om
yCNBJkz7+B7P72vLn8qypNxwDpdodd0tA+Fq0oQvNj3beXAA9TtrsK7eEeVYObPA
cykQ9MI6oBJSdcid8iqoRMnV6ERv1gHQEUDGJzYBiChDr+pP6IF8Ucd2/YsEPH+m
Fr8c/3PpoJ4845GFhxSZMUy8mefYqrPWP0dCk5ut829aU9xcrL21qkpxCvOIl2/9
pnqDcof/kvgog8RSUMwQM8hc5WuOJNHlIXJLxNTJO8NXGwpiMUnrv3CuN5rMOa6y
SIY3mdeBFQ7ZF1jY/MBUQDR9NAgJW6dzOdNxnRXfAKRbkf5hPCukue6ZBYR143rt
1nhxSog6sxFjw5IZ5/EpxsgyMdKydJI2PZRlvkw+/tc+YczDbfTgx7jAKf38hpTm
dgES4mbz4PXH0LbGGlLw+M8ezl1hQzOdxXPKcyPI64iX0sfHFElyyU/oMKngpMOp
D2u9LiLVBQVXdZhZd5dgnScQbpP71y36AM6oyXyeyf4BUH0m95KFmbIlFByhWffI
sLTqW//EF9qPxt6qv3sSmXkmXX2ITNdXRKONCkYS7Ysf1PeIjKf17lvm9FeNUXtm
vH3JGinEFO5bErpeBZ1AW1oNvv5CnnB7FhwlZjfSMblqusDH/79yod/pTPzV8pJj
IxmnKU6m0TkoqO76/U+upQUT3jKRPRH6t7PVmCblILp12BHhwNsCj6VcJXwg9SG6
U06wDEY6bYNd7JIk1EsCVJBmrk+BnlhGl6HveRfsJrbb4hcC0LpifW5FjFZHPP6n
Nwh94IqvJ9Bz+yXudZZBr64WsczEhFHb7bj8zCRoo2VlirGoPWP0mtZo7whEl1LR
5hfv9I6nKXucHv7naas7mhB7QiOXWe5bkGpG7k3v1N2hu2SJ9tJ6UQ+NNXNAZuO3
NuDcOGNObA+kES5kQ9powwezRlKtQySxDrRW4GSk/dkJCXEzZeDQ6c6JiajmdTCF
BRzxx5LbJtGCc1OvjAE2pw46foqliAgPwTsYmiTIVsKSrq/dm5euoB6rE2xLx3oM
7u8ayYgTwj2hafa3QXNzQOPXMzhJ228WznaMtAxmOIq4JIWXQ9wa5dl1bcrRHAc9
OoiFUqMaaKQ4eIPf2YzOfp163dWQV2rOu+WV7tap/S27RTWoNtHSg0uTFUZKo2qf
DGlSbu5vdC5dm6IISO5ZZk6WAq/UkS+MKuotLms8Mw81yR4VeD9n41Hed6CMcO+l
RBvRU7+Xb0t+Fl4QhUsFkWoEu/ii+y/WOKPCO9O/YU1n3ve7U6JxVB86/+1+ODoX
QcS3+LcmWHq+xBNF6NfOdhtU5Au4xUNEsfVtoFg3EBzU0VRYDeBeFFaiURveELUz
Ywkxsju0624beDxfdrVuBr2+CdmchHVZJkq9jnpMKprmP7evXAiOF/VNf2bCy01u
f3hA4qpknZMZ9rGqIC38WSnFOmQs3F4vkz1EO7GEgbtG5Iegb7stGh1EEACSn9IE
l13vXIafM/V3R+Ob2Geer43cRWoIK+5CZSYpqm749XAHkbiIeZeixA/t65xAi2iy
WiBs9nxYtgQ9x4LKwE3Ef1LTOmAqW0aPv7ZDEAJn3OJYz/pr8nAQl0LaFSbIwVto
tjDftjsHbyu8LOsX4ZqqttDcOp/3yv0GH/7wqH+xKdMQkLUupQf6duxFTemj/gwh
MpXRWhJw1OUj2axp1vsF3EdnMY3fFd8CYr7cXmMq8PC+bMpQH+Z855U3fdfOTisg
0fK0oxenC9cEJs2TxKjSVdY9hCpF8Jbk0Y7tKzNwZQShfT2bEsnJS0lSk8oxEaSm
6NfgP5siFGR7CGrJAuIgeBjrQpMRfKdnSi4JP2Bjwn8qk20zauUPEOhEnIesRoLo
TOcV6FPcspvouSniH6FLGNFeReCE5j4Jc/XHdAoM340KCoa90nQcW5MegYhZPkoA
qT7Gx8/XAqNKV4wflT0zQyczfAy6+ie8afWjVGKE2ZI3SDDmHOFKNK7rmSJ80Y9D
PHso/pCaiOq/gwXpqTz+P8moba+HIvH5KX2xPZ3g/6H+OSQZ2VcTahSL4NlEaOWP
E7HI/5P4yGTWp7ET0K4xBFsOkpd9kQJ8yZ+FbUzCXrb2IyJHqHh9iwWfwdn7L0Fc
Scqy5DF0YTJm6xRe43eAhAFYNsLE76fO2LHFBOUJEMDJNMnzSU2riJMt8hlXfJzb
LDxKQPQSayP/lQXkjBeF/6tc1ihuq2ojNZkie6I2czSXAlyHgLmw1fYFenZeGAqk
PoqANbSJfLOLR2aBdLOTyggBSbv6hRsRK77mfa7KaGOPa3Sn1+Kah8KHH3aTJ2a0
SNorfJAG2mHmpmwH+8pxIqC/8aJCTg+2A0aUu/L6X/rrasd2P452Zt+rDJ7rB730
SWoFFRXwuiA0Plqv60xxfPVbV2GA3uptFye6JrkJPTXRAGJRA/d2J8vl/6sDfAiy
ngdkVdUSuDFL3PJNseGAcgz4tzHcapMx59PIVxWQ97PM+OM1ztggDjpshPmnW2/V
30WRlNHVKpfH1BFT6KKuKzoxYqd4QQN9q9MxT4mi77c5LaU92n/EQHHNvhLAfUCA
uAEcJq9dZWfCnpknFCT19BXcXEAPbU/IoxQV1ABgmXxqH4ViWYMSYg+sDr/gKflD
0MWmmovxwqQBjMK+0IyWtCAkdch8+s+IG8uk8fnN7zhENOULr9Xrb5bPPYnuzxat
t4HtEg6MtaMA5Nd1SIidmlrULQa403jwGkehUHtp2S/i/+5/fV/3vQHDi/650QnG
HYlv9C3iIQvrx6gIPQc3afqKefsOgAbpzmKIa/8wJ10jlQxZtSVpXNdulOwzvZew
BsrS0CwvCOI45SDn3PB0y6NhfnDQ6K7T69o+4EnPgtpvZtZ+sOkuLtMdUMGTkSjA
pIYgTJcTGUT7uHIvm+YELt9ItNGHe/j1ib/jeIeZf5ltIOwrT/YLT9PUPBjUXeFb
B7WV2rzxndKXcZCjUFyzhkoBSYqw+n4dkyhYMipFIDqobJ/zsdNsJwHN7bbzBIaa
Hd38cNCJm+KbTZ20ZjQjE5V48H7R+yyTo5pfFq/3ql/HnMfcXd5fVPlMCuLP4pIx
+U8JdcmKKLY3L8Eye1Q/hsbEpnYmQgU8syvY50V5zk78chQCFqeuRMN0LMyUgSnh
4xWmVBsbMapCulMEsGQLNt1CErPMGdEr8whGTAZbUWZAT8XQYWAsGFgDfEweBdif
4TXl1nveY21REkl6ewrUJQkEjukNvvzfkRqlp7w/tmLCp8Wu7mCS9HmC5w8NrkT2
L0bUPegFIFHNcKDD8Tc2eysRA9lYNOtLHgmLpbH+OdhQAtaLcK6s8walRsg0gG9O
pXKxe9Y+BeVRCHP43RsRwcaF4t5iwQ9FxPiUBd55yxV3BYdCBu2rzP+kXbVlFUJO
EGFRK67xbj5bdpNPvT3dYWxV2YC020nvLbBa4h9iUGR/S+pTGf4+McxsqqATxbVk
C/6IjDfe2kTg1EVc8Ke+Tg4nrkclsBSxoaYMxFOi9BVoGA/Ve6I7jGrT8+vzCl29
6bjnUBLOnalyas48ZHDojMyvwBrx5fzJX7zCdzqutpPHq6o0mB92z4rqDtCZRFrw
AGMG+uxdzpX9nU0f29PpINmp+VrpqBZKEoi8v0ImMRVd+CO87F4UrSf3LVQkBg2p
CTyMx5DphJJsvHB3zzjHpgx84w87KD+drfuE68B+BYpj/ZK24QuX2LgweSD52hny
onGXi6MIyeXiIOsUTWyUbUi5v2/vDTukWNPaP/r3dNiBOfNZcOFFv6LvzPkJqM4L
hVY0CUkF+YsloL8Zv5K9zTIeqLEWleYEYBriiq9Xm34dLCf/wBGb+ISnGC9FnqP2
LMZ/adPVf6E4YiRVcbmmcsY0LsHU0rXAK0G2yVLYJMlUFBaN5CaZGZgF3fjA1FLZ
Mgxnpu/vGUboqz0meT1pXJ8TZwdjNhdXy3k2Pa7rmqEEym7Wlwnl/+84DRNPjqC1
O70EErcbwqzhWbAn1vo7t0eyYRSTdAOPNPZ5mtXKqXLsJsDPfwHPyQcRL828hp3J
dNuj9Zv4M1t9EzWdi0OOFbCt+FSFbkV8BVg/Nxyc+lb8pqaKckVpMPDWg0iZ/Mzd
/RAf6zK4WXpXxuOGg6pq2Lt6HfKzV3xW5Ar4YMjuZf8LGbtyzosVod7IBybJBQlp
P/GcEva9gPRTrov4Sv0IHF6v1IKjDm8Y8xFK+M2duL39NkFV5bpDGJp4vHvTWOEH
SOHKrg3q9FZr97YddYeWzz9Nfkc0cbnPRZywCT6mVSvcphwVf1U0ir1Lxxh+GK5U
NS+VrmKRZwuK35lvUkfyEXfQEuRBFL/vzS3ZY1pC25P2+Uy6ZfZgkLtAEFlvxwcF
4QsW5A7AwUy7V6Oq615j5si1OQGDjxV/nXDukAK8Kqvr5UFgGVsJ1Csv2Ma7etOi
9Q0UrBG/Ng49GPx0jFl8zGNSUM9E5BF4/+vadXZHpfgTv23UNOoX6nOxyxYDhN8w
m4Qr/sQ/G2tdl4qtkfG1AeRXgw+uRexAU3NBw+j6tFS03NZLm4qeR1hW3uc3fw2/
kNswKG99inw9RhwbpjM3GKq43QzoP6mOvq9lIZy0E9pb9CK4Sckti8SqKfKISsX4
ilrHB++YbHproVGFI/bqB8VDnDUGnfu6sevCevlTbmtZ+MlmVtF1kZeYFi2zSTkX
/Wt7G1CjverasJguyFFCUTpNOlS4bQ+QFk3+BV6lorDZ2bzAOHz/TwCqfOku9Wj1
1Y7C+x5ZsW6/jTYmeh8DFpbcJ0wVLYKhu4aYaAIDfr9JUxfVL3yBUefNXFkzH2/k
S0O50/57anraU2KgF2zElThy3KkQBk+IwOYbXgJnTs09Vo1IcJ0+zXMZkd0xrfrL
wQzC1wcsoKNrEF9YRJJIO6i238cjvV5xuQ7JajumJencGU5YuYZ48iMje0DXVTlI
+XZ/KGt7i9wQCvTK4mrDiVW3mw215sX2RGqouSdttnAKHuqbsZaz+EH+0zHq6zB2
U0lfXqjs0/AJRe9Lk2+ybQhzneDHVNCItH29YU9CmMTVz/L+qIzlf78wRKY2MQrl
jwEfAXQPOL42Ie0em/G2Ycja7zoDpKikzh44cbvGI9Owucq+WOBKdsFvZWocd9yS
s6Y87gWHR/0GgFMbVKYoMq2J8oZCJerN2AWoaMnAnOzrKJ8fqh/ZrsQQSHTzO/DN
EXa0hR6aJbqeBWcc+cv/bisk6x6N1yAlSr7bg1H3RSeGVZs3aUhf9QFi63O4Dj0A
XieeIC4bEv1L4TWTmbvMdfxf7yGFz063URFcesF5UokEOOcIsC4ACCkOKhiBeHsS
4YCkzhjykIZwEip+/3u4QC3meEDuAfcyzHWCOJg6BTxWUdvIXOq0F7mpM+Ot6ayI
WsIDfv1JU6lUyIJea6obS1bsV4WcXvprTO3TOfOhNwuUoxvyy8KCMcTfLaMR/Ye0
bSwe2HaqmVtxtq7BKPAUWXzvlh5tVdZ//02c2tMr75yfD8D/3lvvYXe9uBNVRPtz
UAxvWnEqg8kt+BRmPfHPyE9I82Jdz5ubEqtmf68D1PtFqbah8ojV4silNNRRtfR/
6B/dMG2c0EBU05N6vSclDAFh8s2F0hLJc+Wtd9wp91B07yn4He47yefaa0rcjvxT
5SGnwKMQeefbkEXLP75BCrv22RtjGsQlFJz/aFcnZmM+L6+RLnT0sZHJpIe2NTPD
D2VwoPAUcdntxXi4xS++hgEF9EyNZzI5oJ7CV5CyR/UpSPcICyL6J5ar0rdf+u/x
lCENnW9AxEiI1NPrvGodLm6oTdduwuTGjLbSoLuERupSq3xuoZ4yUyHcl0bJVvSB
l7/cqJdUBKfpYdkahadRJPEJCFOceXATT94ZFWUv0FfN41NQuxtFsquRvBvqGaBC
TrS6PNa7zTQWMAEcMAsKORwJzfKGLt1vN5ultV0xQVEq3fZGjPKXWTILyiHASA+N
5CqkzXcfgL15rM/4LWaub3GfyLL2DdSMDjhvaDxpRz5RqjhErXBkRF44YDl9tRvX
ZyM94DRyg29gyJ5KoaiLIf2VB//wgA9MSS9TYz+1S5Ec5VzlrI5+vnfQ/7uaxHqj
APKq7Tk15L6fI/dcU6012tIqacXQ13eDaVClHXaR/HtErX1ILuDfmo611hqdJP2z
oV9AlAPjdWXlBAtdCJjEfQ1wZ+BIAruw8mNpOczbIu5Wn7xhmSLYoWbKN+wnEaak
PgRCWce8og2WwGK3CcDjStrEgixP39MV/5JzC5kvNf/jeg3DFv4u9XrP3FMNI0yE
1k/PtPJH7m9Kwh6tg/lut1wtVmqwb+yakBZd49sTtM/HFE6SynoBn3SFwyrrnwxV
Bzj7m4Vx3bVxPWp8oKKxfwz/EP4KBy4F4PUn5Z6U8/zdx3MVMHytC+20UVdLNpzo
n4NW4zT66xudI09jlV7COpggTjDVTl+d9Ydex9VhGaCSQDYEw1nf3FYIPb9kvZZF
d7fBs0WVEeC4U3Ra88fl+S1RHIe/w+/BgQWcYjtZs4ilqbPLfNxmR3SYByzc7NEe
ljDfVQC7YzlLlYwEaGcPVfUbUcWtHUNKqDDC4+jdw7hsXRA3xqVukgWQuqXliX7j
CSy0O01LeoycFV49g2yGWjNSPYjoH3OACPKEXiumRTO05WWAd+EHeE/1R53gBZch
PAem9oE3uJGS3c3NQs9U1gMvFH+zWom7mDULgMgL2ThJsfSOksxZ9+dsGEnGZnrj
YUb0/wCYH0GCS2AJ7dQfKckzM+9Dy9sdeDfizb3m9oLlOg5NrUv4GgGH2mTz8Fku
4cG3Eh1DpBgU2FMLaFf3PZyCMQeObh6U0Pn2iDFPdJiV5Cu9rD7r4+cuDoj4OXt0
tOM3rzw27oQM4A239sVCnNhTXhhW7Gh8ze6vqoKTi63T67BRgV9xyLNcxruEivrc
wMJiQT+ZYuzOs+6ZJuRJODqIku82sKxRDBbslZDorBUyPPNb0dcxDEsIjrDO/HWP
bWxSZi8z376rJlElubS7hykySYo8z0ZCZRjavgdu8vPTnOqhXLfWlLO3oQzETMbA
rukgY5cVJWkY9YTqf1gb+dop45tf8W8Y+N+XKFmygPO88srMXirZT5yA8BCRL1cU
LjMftMx2bwQNio1yCYtgDnjjujPebLg5+fTX+pyQlUetyg/jEioWoAi85BEGu7Q/
YVS+YV8MWnBWKDnHgexxfZo3NDX3WRjiltyFHD7YjlSwGXqg4+nFCyW4kt+k9HRW
hOSf3u7MBdlaMwYSrnE+zmfiYpRpKidNu74YFcrr/oRPcn8qNtWreQrrxpCtvQue
Lt1eEje6jMLjBauoYF43xYg8/PfYSeL3XbCCdHYsmeCGx2v1GPnOTD1H/8B3eiVS
mfuhQ4I21qT3xxowGUVTiKyG9RXMtKy854ekjqz0lQWQ3H9Mz8iePVFNG9wciryp
Ypr4sWGYboLHjtyI81F6SzGClgGez4AR3TioDUyAO2FJUnmlZ6+FtNIZZr0H/UK+
t1AxB4dIRgNLyuC560WVziCP2Xx/Re6ZD1FPc//w2vtGjZ7iNl9EA8p7iFEHhwuU
xG7poEjhurlpQX1ZZ19MSd8LGefDBXdBugp9XJ+2daGysRE9MDHT8kXTzlBwFbNx
rPhpwh3fD4+hQ/ve3dbKUJfAHHw3Qo7/65NsWn3Pjz2k1GQJjDVZ9E8EsuhgpLce
PbtpiGlCOAwa0CnKuNdOThbfOpnGOgJ9ic89A1nUGlBFr8WezHdZ4v9sD3YLuuyz
5VJJKBVEB2UbXJB39FSUIKehYgzCkCjfJCc83bg4FM6XpB0b3JVC2Cfqrp7mmk+z
CdVmBi11wXrBkRHnLlKpW/XI/FirjLXMx+teMRlBktjgDEwUcnQhTtC5VVjBrrje
0XIktiSgCaVxfW2wx7EXl1jDbS1c59iCJFRlDgcj7u1rJrMkBTsIWOuUBb+ma4sO
zxabhN7qpwHj5iSsWJ+2nl1nmfrk02m6vVgNrtSRa7TpLhRZntYD9RvzFQQ19qUn
/XlAdVVstSa8pj9ZSqGh4/PMZjzuMs2Uo5TUrxBPLzIVh5y3W4VYeMgPZYYwcoBx
uIrEWHt8dhNA/+0YNGmnYgxuKunlOsh6d2orNbAlPt8fVXCff7Kh9DtMJOOe6rRS
ChyzwWZBdrxU3OfTYJLoG25CSbCO5fK4y+9KtXWZMqbOs9IZLERJZKaVIKAjQiVM
UUgolbRYrQZljeBgop18/kEQvBuZNRbubuccyGZAxKX8PY6JJTR3x0804VgTtT0F
cLNK38DXqh9NQYI1TwFXESMSwv5xduAukMm/N5Chipi5mRuujpHPcb3wUTcCTu9j
Avrcf4prukLnDAfH0RLHAgZtUmFB10IAOE1Nu9i8I+GVUtDELRP/3oxw4mQwntSE
TEkq48ysinishelm01Gnl3tehfLfYGEb4554uQ9V8YpAv5lUFJbWUTKzvbWky5sS
mllfeG8+LSLqNhRSvcZx6Q6vd7qxdgPIF0S1Y+8fnWSkeRjXYFPYrAHNiILl8JTp
EHdcM3Qb79YzlnsmB5YoaYTCqluKLrXPe2lhNXEz2b2+mmAOU15mbQdtBSitKdX4
6dAvZknkaLQ9hK0J3X5zdOrkNJ0SemK6ryeaGNyXF9UakgfYZZ+jmB8vX6Mg9B7q
2G0s5rB3uBt+0RM78EwgN+Zb2+oLDdmNBw8lIpJQbdKak9ouSQ6Kb/M7sMWp6ok3
RJdmJJtL6FjQVfRgUaBiSzIbv+NRSwe7nfGgdc+aJxHNcphcbrqO5FFID8bsLf36
Yv67YeUHZcJCE0eGgxLpj4zUuRn1kn/DfRT8UGgNzrqwIS9B8Dpzq1jNO0h6iDVX
OwcfPBgdhMJJJwL3r0qlH2oP9PtFngrNNge+nAZ2mTdjiTRnwKaPjnlP3XgXZzaG
+3cwsSRpWi1O+Vt+DNSMJddAindogkktUu8odo+TJ/kpVW/bigLoC9edGTS9yKdX
uQb2UU3cxRSEn+elFwtwUSbY6TkiWeTmLWGoa6GdmAoA1sha+pyiYJm8g8FtldHX
T+c/Gu0f2t9Fi/HIUXhMouBZupNSYdaVb0i6t51TZahBwhdcQDOnO6vi6dyiACc4
CzkWBcG7OYQ7+hFvVsYL9E6jnjOwgQfRCT+Ac/0l8k52EY7W+7Hoxj6NatRr2OZk
DYthd8NOUiooD67TfW/5osNIPowQb65DyPegwFxE3H6hPUI4iE1ck2n+XDmMBkPh
oWbjVUGC/n3d4cXD0OBxlcQ3SGxPT0m6+28GHxNNOUshOIa4gSwLtoy20jddbSjZ
juv7G+hrIvJOOyUVdvCa5+UYKT7Meiwq+oZEmwldu6RHr/HEq/LSLMXD3M0Bu2PC
pTW/Ebi8G5sChMr+Cps1ri1cabh2kbpYpZhC9k86PeKJPqmTyFtYnXcSFl3rylvl
cqJ7a5+4XR06devch9sErmEGd0pavRFi++Tm4C8OjfKCU9ujoI2AxJw2XbvV1OJz
g/p7DFlBkLQtb4b8hPr8S3XVqTzkAwaelXlMDsIeyY24r1sV9wmY05/hEKJ0jqGk
aAVaxPweUmtHLYsYHj7bgEadMRXP/X+Z75aIXvElw1/C50e8lbMiECChqGXFhpma
HEN6J4jwYnZl2qegaPdirJkqBsYNeEsFgaz/HUWTBYFyh/6WILaW2E0XBrK3XEca
x/UXqzr7VCxjsq+9MIq9ddwkUeNi53jGTALEwijAWprHDOhE2fZG9zNOQQe1mVoY
dOBDpJdNt5tHYrXTzNs0UxWUL7S7JnQxwuHZVLxu1fTS9wr0WVeSHf/maA6astHa
FLrj0VYvDsolzMwAXad0DX0jzXEEzr2P3CZeewqtoR0x38pj/TktsGUBCyyYTs0C
scevtAyDciSlTfS6K5kecYsszl/gVIf5LSU6BYrx8OKjn5E1jUuq8YyFNqXHpZI0
vsq25qxYQ3iAms7hQZ2EaPGGFPsQLYX7KWefkVZBFBR6/gIibnqqE9sGUmQdSkjt
YUm9OAAvhjGcTV3nxKF2BuQ89fXzCeFmfydI/peXi4V/WJFO2V+MX051svZQ5bfD
WqsEcf5IUY/fK6+eBN6ldWigVer9gurFAQWL6aZm3K9OayDq6Xgj5vwuakndlxPk
Ud62A8mtIoKInx7N0MjLUe5oUxBqRUln8Hln4TpcqUKQztgrjvK4fZB0LbG0QAze
q6aS1QYBlL4B6dEjLJCJXYJl+RGa5F8bwvGl6jJwh3uAHYRN9qrYzFA6Okd4R7s9
JPOecy4Av7ZuOlsDv5DYrdoaBATYx9gvoNpHA9IGicg4QQeu3YRWpOkLbWJwcBmA
lcxLrU4GIIWjILBUXsj3Of1wyoK6D5KkMA/TpnITVTX0H0TaR1QqvCmvFxU1xk1V
unGlRvxs4xf+lw2VF4cHdVBk9mAK02YrNvqLivwW9MLqtBMG/CbF5nQfxUlIn3J3
uqqbVflytVNcEzp7cGtpwCwgxsRPPlEBXLv2HWcXklClmiJxnQWsrJvsobpfuKSy
O03MqVAaN85wEXIk63sn6iYMvfvCYbuqj5pLSA8VnIimcEqJXMwpUuz9nPFl2PzJ
4wfarEPjHDTcz4ane8gu/ZGXFYEipvebLzlLOcF1+vER1h99KdIgPxUwdpIdWQ6k
35URtNFGITLwGPeDjhsjQri5pr6JSlyISBzHsqmf5B6w/AJVqiJ+KKNMAr/BdtVh
I0GkxHy+7grZ68Aw16O7irEEpJvLeO+/+yF8l9UDobDS1kljwHZQBlR4J4340LjW
GRzq59yiz8vuTfknJql1ZO4Ny7HV1qcLxw6hAf7tC0R157Lxyo1HDXKFbT06bw47
Th6GHZXVGLM+xJv7cLkywXkamwg2ynO2co4zxLpRxfPRKmlE+Ue4HJq5RvTQIE9x
+zDJUEj6sTB7EdfbHLx3Tf29c0X0thUeEuD2/0nofp5JZrT3/7WPkb+CEJG1dZlA
SH/P1MKIk2atcOJkLr34n7fTAPpW/TEaLk5EnwI2kuH9cAJ1CUMr/e2cnt9TzXBx
jgm9ar+zXPojEQ9UsH04XIewd7gqS1e7H4bso94zhSy+BwwkNEONdoqfi40ovvpS
AV/JxZ1CfT/E9yJ8l7CW85WRKY4VfcWE7VZgtDh5PN99DCqw08gxBUGSw+KBrPe3
6HeilF57dPZK5swO0wYa3tcf2f5pF5JpxRHV7vUu8TCtYS84Lcyk00PQiv/ISmBY
MHkQ9UaZDlQqmnbcHUEac25lgXFS+xBcI5bSfiMoA4z6MDj18VIEFqCAe2dO7QFs
1NrRCp07SE1Dc3xulSiu0uhN5W0q1mSM8zOlLHxO1LzZHwyMQx3yvI8+8OTf7MMW
l1raI3nC3RouxSxZBdCUnjXFVLz01BdK0wyK7ImQ4cCKV+1fJ3B57V/qpd7ovUSh
TuBRUdmz7GiX0rIT7sqvSCsjnOvWxwui5UVwMxFWJZwG5ujkXJRegP+Cb2S8tATu
i+eWkMYtQ22HWVOnlHCdorsRl74O5xWVgSBSt4jbgmWrhfJq7QXWsufBmot3yLwC
VKkdBlZAZ5e+tSF3dz52pUPhseYYDgTNgfUqS6fD09uTuMMFwVqqk0zw7dqec5/c
PTQvWh8TwkppjzKk4x3+SgikN3r/qiuUF2hJ6dyFRaIjHHBE77EwcWOclno1G/t/
ascCDT2BVEhFzNVvEYn2/eEyc3YgqGhDWkJ2iN36QqQNJ93edbREnbbWciXBpBw9
Q0oMg6nNCQWbHMEhmR+t8D8AvKEUsGbIAKXgB89rE+JlpT0Z/YJpLZ1Nccke0TKN
If9S0SuhNwmtsaiiaBrs+6yO64nmkAQRMtFzqYjUlBFe+k5gOiBMd25cx00+M45i
5XXeGAaqV06Z1LmWsdTG7s3AgTM3Ufns3lI4n49t5i7W7YMNa/H5nRQUp4PNI9cg
EMs+cOLm4cY3dLxYdKrbZyVzF3aUU/UThuN2ja/Rfb+xi26DcjKUP3Rd3L2N+1XK
PSlg+BkGjcvOTwOztriDj7NviCPojgzgDK8ZJX+2pGsJ5mcjDZ/67iUOnUSXtZtO
UTBqCpsqrNhi51BOSVWG7i+zAXVmpFiKyZX2oP44a1nwLUj4S9DHoPgybTD3yium
m7H2D3jNMBxkXCRfTcco6YfXAyyCic/visx3TOWaMLxGxEJfx5StwQP8dZcQTR4r
sTITaLbBt1FDPwfwzV6OJXowZ4OEmpng2NBAJ+ybDUUgdIsDmVwSLeXNc44iz30j
O6prEhysqf1kwxqQz6gvRUUgpMZXyuwDoAVBsGYmPaxAt+TbJyTSsXE1DQz8JhA4
rE6ZxdrTX0VPmZhBW7qJBVSHNSL6ISxMGTE6rmQF7Cpp1PlLjDvNUKGJijR2s4xU
C6mpSuRcXLRa42b7eZRaNCgSUs1Y+C4RJbg7VC6XDlbbOunCRaZx4iTC37RQUZ/C
UspAA7APXq0Lpk9kEBEq6WPmvuMCgKs8ZaYzRyrfBeia2+Uoc7wlqjlld5KuvhdV
g5e8HzZlKiAFF/BuKBFzSEkYxUBUAaU9ZiV7ph7Rj+4RMLXK8WRwlRJK4P877g53
8D4Jy67Uh6q381UcdxBsxPWbb4KirTrYDlGFgC7FL2mM6EfkfVrQ2opB9VuwN8yS
y2jk/MasZja2I02ox0H1Mq3TQ9vGfBHKsV8JFtyQ+1rFCB4EO9jT/t1PzzJK/1L5
E1e+W8+lUt7vTixIDR0BBlf1mF7xfPkQoTdUWxDrDZgaW6JzfchdSyaGa6Z2oyjc
oqEctsnqhnq+B7nnxwmzuNGz794Dx3UbqAQL1pekhPCYohSIn2W85n75apFyNnca
iK3usd2nq1RR2ULaTRS+tbkUYpwnDssT2xKT2BAfUYmwEB7Va8N80AAwLz6SX2R5
y27oe86H6YtpLv7rJpZ3feI3jqRIpWQhgdb3ybA/74OlQMJaCJTrGMVCQ/y73NdH
ayWam92ICfqWwmnp3gZ6pQO6GyR6J46rrWeOiM5whu5WgXIUUJmRDrgFm0PSAwuv
vxi5XSKqyQoWLLEPNWK4BK9diWwz0Hqdx2xnnvcxkrLUunpPrfWcdp7iB2kLnoms
mcYDNOpba8JyoQMsl2xdnJYVh5nW+zhlF/L6bU2WNsaB12tki3ULN5rD4c/mLRfj
NWbSeBgGHRntyDfqxSwRZAKynzRyn5Cw7jWzN70HoO2/RBslcpyYCWvC60ONXQ7f
X1ZQ/0Q5AmTOn9lIAL3l5Lay0/e9r103EsRV3wS9l9QYFM7taH6/4XzvrYxtvCra
PIODzsjVhBylKWde61UhEK81nUvSxxtwFnr/lSGInvGMHQph6O4PZv8UOMDZL8hF
idQuNoZmNSdjaunqqcIjvEWITfpmvGALEh4pfSOT5DSds5C69QvMvzJDv6oaS9NI
vkdnSSwqdPLI7WZSkoNlhPD7NNlfe62xGA52DpT5SNOQ9ZViYQSKODYVDakn4DPH
hPHYBeLi21Bm9oPGLRK5i+YqICL5N0kqTYtAobl5xhi+HBdPcVegsJxqZQBTL0Nq
zsJ6bsC3QmjuwkIb+TDN6GF1sXhmfDaEwGhYfU0DAw4L53W+ANqSFsTOm1Zq+qJ/
q+832do64UVB2CjGi9fasRQafa0woTWQjBgumgN6C+qobpigN6MP3gBw60tyExq6
RR9UcgUsLOSQhn5D0zq4ZW8SoRrne0YjFdakUPX4X8bG8uH55Ax62fKv+XH39q23
Gd8aVVQRpJEeF3ZsLj50p5ab3f+WDsq8Q4NdRdZaD7Ka8JM9iQ5JbQvVWh48MBqf
AjpJmVxoOqvVnCbJrFqgeguBt3+l2XWPllClFqaiU/lgcoWIBW/s3tmJLe7jQ+l/
fgkRePVrTjitnlW9xX0KleJFHFOr0Yp9Uysw2glHyjCTwXcPpdIvx3GtzouYRvRT
+E+M+zrxpuICUcG4JlOV0Dx4BI1grh3jY38v3qUz8YTatBC6LmgMKU0CscL6Rb6G
s7xcnD3/2KSbSHQjK2fV7FoxisLSu0MKhlYy59kc8KwTem3GsjVUPrEZXeAAKAtO
QCGjkbov99f6uEBXWvtEjUfJLvDzKiM7CEyOfd66qqpbvcZvZHVmGiyR++L4pzyz
niF0lhXNcJ+ZodgU3vfXDHNr1fM7SUSMOY0bxvYaHEUE986NLrqB4cHdC4PnOGSt
3lZLU6riwfXMFxVcwQqZg+dyXoxdhsWuYfW96fy5kKtm086ACbWpKd2hxkfEZ+jM
cwqufJqE1r86tlutLCZ7fxnX9NesGwAjvZyRaE7iDkGTWhjU7E8YBl1lCRXEVnfl
3xdGc8QE8G6G/dvrgTLDEyjpEQcasuXALnU0kyMQnZY2vPb6gcc3MGfcNwprpBzL
9fT/foyonDnpfr0fuDjbNeboVaqSNN9MOhi2M15HRQRJ55myPh+FzZIWlhRvU061
yHRXpasbTnSxd7OqmHTC32GrHt+ZUUx4zd8UWJ6/8HWU5cm22V3GplQGWw9ufDYQ
1ahPOFfjhYBYmOhF9cX12f0YyEDndIoEeZAW20zbjsZzMDR81tsGXfclsHXfNxd8
i/MwgZVd4ek4iTnu+2z9ACvsR1BtKdf4xyc3RU3EsyILoaFDYlQHp5Vd8ho+uSd8
OMFyFLDlTpL7qTP2H313nfLUHovQhH5/pnMR9BZGAqzu75lZIljiSk/r3+vrurmx
E3drUq7FlMiyeaGMIi/5KFM908HFXiFOC5CuP9Wx9Emuq1Y7/nTp7+SiWvW7Qedc
2kqt3lXmQWJ1LwZLp3DtZQFz/yqNQWViwKDFEeNbsXpBbkMtfBc60Uzj/SjFuvsv
yORotRxPSq1eYHEYxbMd033T0qjowdU21jRudIxNgUhWOro378dMjmHbYm2rYZZZ
FXePbMt7OW/bXqU+CBpbSpf6ABUh1v9PVdDZmQmujfnDpNOqFWR5rHfBnQ+v12Eg
trkUKfhVd+lxTbrBeB1Ftqmca5O3xuFHxsF6NuEh6zX2SyGeqCwDJv/wrihgykkZ
mA2R439GNwh/Id1TSpXHF5Z2j/CwO5gDj+FJ0r2Ru5HoXxAkvTu+0ARasKpdlNgn
baaKQ0Xvp3KzWU9vfus2WzIqZNHSKXStTknoyoKKd2y+VGctr2NcRKE8RxgG1cQL
30hH6Z+W/qK0kIZCZkE9ga2ZBwLcFRkppFykY/c7143Uqw1uzvpbPs87jWDkuCyy
O0wB3OBm50iTEHt5tVjNAa3M0+ydXznkfYOps2WqRDHjQD4W5eO+4fxJ2rT8g0IZ
UwWxx2/Lk9KU0sEfiEwpSP+KiqrN292eGYfx9vnjSWoNx02qtX3jXERAlR4NjBDG
LB0lAQ4otdAWC9kvI+hb0omf/5M91mxO1rI2SNCB/WY7rg8YCU1F//YfOlhF4mvS
DWrv2KkrqszQnnYs2BohdP4Pg1iiFU5Z3msd+H/vrwhbEwd6kyve2vba5bB0UGab
zLSgtkOu3WPLQiqq5m7WF1Qo3RrxIcSpIGhqL7cq9R0Usb9jWsvd0lLTaGIFmH+2
0py6IGXYe4xrma8uyWVbmpniPyOK/ygjMJAxU6eyXltIK0vtJp0XP3IkTmSQgi2s
JL4c0gCYO/mudf9oi7DYW2lplATdKeCjhZidJ9ySK0u7NXfzYhZQkjKLUyL+t86Z
NWNj+ggjYIzWrRzlCaP7qkkIXi2IdHKqhuiEbEDJjAI+/1nnz6OFrTnpA//d3hmT
bl040loTDRYfVWf4sFCNDt4t+Dfd0SVrsR3dc+lnH0X3eSSafT/Eibj512yWmTvG
JCN6Lvi8u6vCrh/qsDnwUgHWBMoAKKYk+M001CZj+vX9q0RZ/stKcRD4oI/efTZR
983S267IfVQOFZ22lrx9G+A5Qq2CvbpS4FyWpCVD1qrNDx1AwDIJPzCGglzGIeIk
aLVvqnHIs2pO8K4+5oKZDYsEEkwSQIX46Jkwqva/QETwolAIvT/rcfqBNnWNMiEI
snYpTbgjH8mmDt1cTQfqCHRdjyw7oHFhhFO+ACT+/VQ5kr+z0ddyu8WxAt05sb9H
QOeKFgjKWPTCZLwY6abbH73VCHHQUpt+fXErS8TNMvUwpaVQabBqyo6/pAGbVsOv
8VGqo03/QMtGS1aDrp6nlN/Sw86au7Tprv43GeDMbpSbtI3+banijDRqYyLQd/hj
EYrIeO1meAnHvB0ZqlmPpZFko59MhO0lTmi+uq/NxzEogs6BT3Y23K3CMESRwD5a
ahIcbjJm+I4HzBOPGLTQ1YdFs1WR4FfW8XE158jN/d6N5gPMcbf0muKSB8d4xS+0
Q4SR76QMm7m9oy+4twGHfp++Be/aKY2pRUpMfwGgq1QPCPthE+QQHYWGP5cdeXSE
iXOiulEDPei2+TulwwfWhGS2ewIDQ/5aq2NPBU1Vk1jlEQ/ZMVrk/waPIWrenxNO
BijCZQQFnm8g/XInqVFum89sEYQkU+Kk210HGARvsa9KKyAjUbkW5dLsLW17Tl4X
FAGCwtJEleaEW9mRGAhHQ6suPLaz23rYAiDbY1PqwzAkuB2Yq8MiApfeykMnclno
F+5aXEd8/E017iuXgczTaoZzdWXQjFG5ZSiHmjBnKDh0lvTDKIcOKp/k1A4W4Nyu
kb4KhPwS6Jsq5Oid4EM0jnr0912GtI0sqPSjpwdU1Jaz/VXbUNG3xMq0GuKPBDK9
5g17NDxqCl3F01ugGAlToTiBwvP4/hrvKDQFQRZXPXo2TAOX/z8pY1mSCBWuu1Av
4OBZZXz35LKKZ4zWPSD9jMAnAGCxa4tW2cLumvCdp3qsgiihMD6Tuxo5TD5wrgdc
7cgAPMEnY746kyerlWMJNwmdiH5vd9YBLtV4/eDry63f9ruU947tVAMxvGahQMSE
4HA6dUvYzcGTsdlZ+eI0TcVZXh9N1V5150zYLM6/I+/EAxSAnoC1O+rBxBGwEw3i
gY1VrfpQfyhDIjW06Y5TaEpmdxiJtlbjAd72Eu1jot7NXV89UEcEJrH86ae3Xuvq
W+aVJnaJwRu/gu1YrUG2/WDlUoTLKFHDzyxwW4f9LDhvMdzlzXOzhP6vt/mUIdLc
MVgwCYwvDQlgiq86V/2X/G6W/p6G3/25dC/UHjVb7tjqTs5g8hButeUJPwcQ+bsH
xSzjBfOr4tssM47kLmzUFXKMVDTxz/8G8o7pDva1eGH7cYr+S+0BtxS46X/hTYqf
sprpH+Apc8Jn4jAnYkyfB/q4BbMX/Ti6ExdKwfyJcagQz9cyeKXPoWr8OBQz4SRY
jeVrh+aw2QDIt1p+cprx1IFZ4OF8eNf6zLjvmWEqLs7Corfey/OIS6RmPaltTDn3
BwJec9FFswiPmNA6LD8MyhYpxj4LqjTbgR9uYv4PW3b3ACWmgkDsiAHdvxct1fUa
PT6Pwjmee6Z6PbrbA6Yv9ZcsoJqkUOV/F9n5exSVFDImqxAiNSaOI58cY9mJmgc/
9P4MTB0eF266zjrSVp+V5CSktG3LadKuEPV7JUIevekX8dyYWQYKkVBWfG16kv0q
VeaFKmEFqdwKKvpm/SOXXFtn2hG+j6K9RyYdOomnpYGE8rVowRDMDuEa+Ac/cmK9
FXOBVqVR+K1Q9+YwPoGseGD9FKG0enTvWEN9Qkd2CqmlMdAi1Ma1M3Jl2jB2AbSM
fNfrFASfMrAcWZmE9IyWt7JHu4uj3jSO9bprxadqDfLqvQEE/GCcJJ5AWO1+cC3S
mGm4UXJH7S6s0gBEbx9hjMzy72TQRSbrPEcs1HjJ0wPxuZGaFHKvl0niOOpnet3a
I8WEDd/uWTrW2pj+TlEcyz/p299IYBO4fsjBBRyRJweFrI/HrvYOdYa1rC/wCwCG
cMyVWdHFKlVOG0M0f9Kaamz0x8+Hshx6rVHDXSfYaoMyTGVghKALdJ6b5GzZOlBj
ngUgxoSmk/QQjcDEPiGzmw0DYvDoA+kvcOyS4RQSlIAWH9wU9r6Y7NDMLdLHM6To
WnnMeat9v1xezTGF0BQPxBj59Tj/lwWWQluUbFjc9vyb2vXWoFhbfrLKtG1imtLA
V0cJicxoZ/ZqLdSxAxkYz+7PW084Q7+5ft3WhMULeJ5T82w/qhjCgDzfYHuZhBKa
oyKGYik2L/nj4R2QamIdMofKyJgY2JiUkD3b6ntIm5EzjPGw8ozK6ZTFxm/Vh5A+
AePqHHXDnbwtIifRdU1BCA9KYZRQMEneD+9WUV3TNZ06bZPWs7n92g2VDGZ+DE+j
eJMxce977dAH2BQiBeraVJjAffAcq3wBpVuEwJZ+ncsiymqzMyWLX1yzMvofChP1
iIHKCaSnkC5RQoRdVIJilL9f/v2n0igdUtQfNLJym43nxkWPU5+MYYnpjDcZvtBp
S01qe/eZqFWOp/RUhIStUWR62lyIt0LXrDt6d5SXTe3x5frtHP2v+EAMVjkt4IHq
a35Rh82bkoqs01f0EMTCbdjO3oyyTCR82uKxgd6I84iTGvDdSS5WGundvJCv0dSe
KaUwt8fbVPU7oAcm6YW1vtcgcgXBWv+CItF0+ik4s+qHO3qFVbrmJ3kU7QIuCic/
6gxlXTwNaH6gMc6UJ2CisKDPi4kJz9u+ei3Yej7h0x8q70QN/tDF6shAqg/Y4OYA
eukapK0cMakc0OwKNaSxfLnLALb1yAeOO6I70/J/a7zgOcV9iuvxUZqwhZsthVNf
8AvX3zt5vQM9UE0BuaTBFcsGwCLIKlbwpzi+niENf8kncT1FuNj08fvp80i+VnE4
XgaSqCf06zY5GW7JnKDJf4DN4f7+9RRnJOJB4WXVM3yXmSGwFW5QmHT2wWoDHmKs
03HVle2IYt6f/HsVycyJSe8zJtZI1m6V5W4Hw56q4QlVEIIRQCaptJBOggedqdJs
AaiolQjBRdtGfgEFsnO+Ri/lMWYLKh8ezqug9IyrDt1kH1KytBr2ye7CSqM5Yr15
zKrmzfWc+J7r7C1+SGo0etH7E6ljEqos3UETmrG3Q0OZh0rqPKMIeD14DsQXplhS
iUQYGTZZ4Hgiq+VjynUET1z+Kxgv6Dnv8v/Gn6YfYkEaX7qX/DnAh4QqbRW3fkEO
jJ5PmhI6Gg31DFbUY3rBStOdfGzawlgVKKa5y9HPrO0t5bW38lIjwHGguKMMlMlN
gsGPRrwCgw4PJxfZdExbMq6oaQWegyhWEwMf2g1VOoMROBWAa8mVxa49Axti8FCq
JDU1VHLf7BoWScwMeKXykBpbe/WjL884XVWH7mVjd1+jYPmzldsmkUCeEcUjQDUo
woPPoDzaDVYy4lA8ckTtGdSxLeg9hx2FQSwT+B5GGGXhTo6Y8K1FjxCqnwFwHH8S
OAZdBaD50KObzhAsb+KTwySbQ2fhz4nkxMSHbDVn+fB99oXlTnNfMUSIBJapHFyS
JQbEhevC7FAff3Ox5NzMP6z7EtY34YXbvqmFwc4PqTJS2VWVqhqBckeAa7FbtuL2
ky/PeC0CQ92JtHpNvByrqbFFkdF8SRM6AIJaIklQf5vRmN6lKnYxODU65RVGXmsJ
pDGvAimlT6omFxf+4/qg7uI/gZBQfs7H8GlViQlYWR17aW7u5xlMNtcN3WwnS+iJ
GTeq8qLAxmmjif52GBUxgZ77h1Nt1QJleFrpkprSEoHgXCD0tSxWd9aaY08WjHtv
CMD/v2h/23qJ2AIBkA7bWgwTjeAzNaX7lWM6QvCihAdSCOXx0UwKacM79s1rViC/
d7kDzgpUN0HelJ0xMEowBz+wIgTtgeU6mDLINeTHtYY4Ragn0yML+qJS65Qi+n06
1pOLw6m/VS0GYceuPZvyp2YR4FOEtd/DhALpAgwOI6HNyynvdgS/2LJyavnUQOM7
T4HKXthE1Tr6uocIVo8Pvo6G8nJBQS3u9sG9WwT7QkQYIwzDWdWDBSyQT8IxShr/
MKycENiUbudw0SkqOONA4t5dhXjKoMd+iLo0lE/ywoSLtuVt59AxC+3CnnhLzqmk
1stOE4ZvB1ORQk3tT1bzUB3cIfwwe+wUKH/+GhhgYPkOO3TDUh24I5thIvqJ4dam
1QU18OSRXhiZuPK5UbGgAlnieKPwFYCUQnT6XqM/5wuc2VFPnqmn37EJlzewottf
CbEM8x+Wq98pZ7Hnjefu78mCw8mq65e1oc9wH58y9viRF/1fuSnS00291Po5Y0rF
+z5MhJW09+yPFO17N9qDmSbgfYN3zIA5eeOmmDkom9QKvaR6mk52vsZ9tu48h994
21mKIoXdubxup4HA6yBxmWVRvzOvPFy/Km7Rer08ZzaD9K3w5HbGJYgq/lXoYe5y
pg/WteG/NHiPtnm6zYQ6z8MrSra81GwRvEn76M15J3Gb4ZKHoCg0tCZGI2PeaqUH
fh5nlrXQH/IbnoVnk0DDVhjpXCn4qMed4qLc4OG+IJ7jiMTYnvfUAG8M1xrsXu75
TwPtQ/anYlz9LGwUCzd8qjS673BW5o1Zjf6/tS2mo8VrB6MZ4SSg5uepAZxi3pic
pyrGATA/OnAxqW4zzE+Cg6NmZ88V+GkNrw8MO7p5vc6OHo71W5BkQVzlpBBgruXa
Db+JSpWkSfsJHh3ia1ru/quiJnClNIaptGoosRtoAY36fhSKqq1ZLQTNnsY6G862
IznT6irhCJGezcJS+cCXj6GSzdBgXtHG94n6riTI9NSwwFhM/eFAmmfJOsFUk2fH
gvS9jNJJEyywKMWroR+20bqsk7e6nxTnfSiPuWB/Te5QOS4ZIG/ICYeAdr60TRPf
PbbF+PZ5cPT+wISxtHaYjbW1t5LFstbT9eC3YRJ12c3UiDPxbT8CY3Zk8ynE55D8
lkTj19EAuRekrzaRV6scW40u+kZyfSwuv/rmHohtGB0mdE70DcGfnCcr4a4hfSpi
oWrywCLrjrKV738mwPdvMRpAA/omN9p14qKIv3/YbzksxrQyzw3Dz4axZH567UNU
c5bZCVgsTsObnSahh/a8tUptFSMQeqgMRnxYo7+M3XCQOGQn/MQ5nNQ33TBEQBrm
bdJ5KxlB/fr/5sK10uD4jtsdAurRxHxAZm9eVgWzGI5OoHwd0BLUjOH+X9aKvECI
TiltyTWxhSp9t0bJ4kbhxjolnSEKwK0UtrPehm/lw7OAKXSTNtBCtiKhR53aJw2D
BlIfBgf3sqAztJWP/b6KcqQt+S50oINPs/dxIhKSemz+ECX6i+G+OIpMwlIVxP3a
QcSLM4R9gwCp/uxaAwckzSpaK/4nvItyBSEAcV0fvfd8ByW0Pxit8sh1eW91mg+n
rXBnV1ysG6lA/3N1Ct0M1qzIL0SsWGUh3s9UhEv9UfUbwEJTCLmf01nB84rKoaAm
NdUnWgxrYRr++m4ga4uYp96h4pNE4SfoKCeyYZ2EKHh0UJnn7lwuxDK9CZtHkf9p
k/lyUg/uMrwUkCsoUN383Qjdd+vX3Ljz5djxQQ8IApY2EOhReCJ5y2dnCMn3oMJH
gHFB0NUqtil/8YuWl22N6wQa8/Hg/GSL41Q5nFo2IIMS6M4nbzECIukKYQw2cscT
tiXbNCbCKeUyPntvmGvaaAUItPeDJqvwMMMyqCLO/xvtX9Hf5+9+wWVvwBa3kinY
vY5kOFgPcY9w/r2jF+phJ23pQW1qg5qwjTReRgppgjY20kdj4Ilm7ffYCmqOMjOI
WPwCuemOUKeVbKO25+avJvxR3nSUFZRZyR+LcHMpB61bfmniQXs5zuS/QhpLA7Uu
yaX1HQU9OkSYikP8TGjFdwAGxpILDArAMDEtioK3Xs5+4YQIXMg+4kXAvkIUSYHo
oMS8JIXqET+TkEAC8oBpWHOirR0JnlZQTq8cpR+Cjn0CDdWVpREE4FMXZETTYBlO
v6mq7JpTMyqbYXwxA3Rb+YTc9Inehwudr9sqUCP98zPdLpvkzbmzd59H8rXCtlrt
rHMMUa8d6BJAT4JnyCUUgLwh5SA74lCgV7hxnBMQBENPQQe+sxL4It78b3zTXz7A
QsaxRZC6yWjNYDWyQUBK01TiK0U0JFxnO5H1j0nEtiKV5R1+WTeDd8omaAdwfCw6
SGgAVXh0tVu4gNQ+TtMKQvTyMeNbvJHCbkvlO3koMXEtdB/iMaQVg+hPcfCk2sfp
x41QazEFuCKa2E36xtETGkD+Aaa22MunT/zkONeip/tuz7ShagAqeawuS2qr8rxD
FHWaJqzjdUU1WFi9ytuY7sT1iuObO0U3ETD3lGRzPkBvY6qB8aGhKuI4esqDvjeH
yBO9yHDqJKyebFn0u82ERFlTOyJO3ngi5P+XpMuF7UuDS90SEFiTVOZB/Hq3dXEj
uBE8WN2wypKRoFoP62xOyKfcPI4A9e5JcOEEJT1e+AWLbT5JuxAfvHfTYVFDS4cA
tatcx00Lg7mc1j2lkowFKbW/lZHsd58NbuMhMJfPPBE6G4julWH+0Y/GjkxcEwDT
s+NjWdtOFsqiLbXxYnR0cnmUd+5oJ+tqjdkjSj5acnr7168n19AVCghPoC27fEbr
c3tBiM8wmT0wDjkzWgM7X6QAabxLH6P9mpQqfYe/kMq0S6gBk9LXrhP1tklkAOw/
33PYQ8P+B10rSnoK5Ft8VLZowazq0Yn4fWl0A1Xszp6HH0toPpG+5xMyGbQzgYb1
kLS4eALWBqqta4KXRq5Dn0cC2pHM5B03S841w91vNv/3xt0pj+T89xuvJACCkEQq
BmThdUhoMuLsplJdj8IIqiMSl22r49dc+nOOdABANPi9yAebYFtAW7wvwmmZs9zI
GzOxywvv5ni+Xj4yAycQ/hJSzHv2P0cV4CfEaGMluuypXsnBdIyoaI5mr1rVLe7e
PbBiMmKQCkmvJDeCF32M13P2g2TZ9pdSMlPNsqv/DiS1HUe8aE8kfZ5v3iyDiedp
AWtypJnpZcX3Uu1XuJnrFXMHRj5jSoFpMlMv5jDSrYOwiQYyyvQ7+N3VKViu179M
d4z/TVd8tdjlBzWCSkqqTIoSz2yLo9buVi+OU/aJlOpPEPT/uR8KCWBozC071ROK
TaW77LFqru2LxKsNVYTedIv2IWbyuG17hdwowyREkV6SLpcy+J2Tt1oGng6dUA3+
jvlBZIpR74Ztaih6QqF8SbqLFL/CQtqSFzwrnZqKx8CaFqzdB3wP9mMOtaDdLMvV
q80TCiP568paCxIbJwKikps141+b0JQb0Cqz6gAg5N9UTAkjYrI45tE04i7l9keI
ZdjtYZjc4Qony8UGdhDwbiXJKv8Hk1yGuL5udv50jbV3dji3jiko47NQu20C8G98
ccBCVNFFMrNq7J8tgiY+ZX2YuJp4wPTQ8k3Rxhk8ZkshuoqHsv7yemyu5Pfvp2ik
5Uom6DUMsj4N8gFgHs2NIpXIlGvhYmC+aHkdWaULIWZyUT00a58MIXKPo8qaCcjW
21Y80EdgGnNB+rPpEIqg3MXoFgER9zPlbP8spdIOAMqRrUOdAHPIMMp4Ko7rsPev
j1Fj+QNs9ZLJy26ydHWy9scVUwAmJDwKl0KjWvQqLu0HPIkTd0feQpBzFkGghaD6
nQvyG6fhEEG9N0N0czk9D5zSrfcUapC9tHKtTKYtC17NgOFFLvkubsidFHy4Ov6z
OC7pplprQj9IQ4g61Fd1xaq2niFNeGfWNWP6H2UyLDJJBVEiqlQ7LMC1SYvAUIur
Ud/OyOy3wVmFruK0CYbB+G3xYPJgANaV7m2/zGkEP5oGBdI0LIncM8NU9kyn05dp
9Rlygilex8Kw2qCg4OOP3emXpj/auTRX0cMOuiZv8DnD/SncPQkNF5xM2R3wxnle
x91PPVK9sZseLvsU3dJ+xrkd8mimkbqLIo1TOvdVI1O+6uUGevT4IEjPc+6vWv59
iqccpYFUEUjJnxUgz6zAOwLaYI81/2hqAflvE1OVoeAVEB8Mra/dbBr5wbiU2XEh
rBlg/be5iXD+oweHK0FJve7DgPxrh5ft7T7FTzxDFAxYm1U4F06wmN3nAMxJC3GK
LUTTUfJpybYQ6HSc/HS4vUpFt7MrfFW+uJ/y84Y9h99E+EgE8OswcpIEEAAIOemL
oFp6kYD19nyMaqaoY+s+pVwF3oNCBwM+y1ChNSde2HXQRLTdatbyXLyiA6Dsth60
rHpsY7kMuLxfqTz0xE8kgl+zuEa0RL81VdoPdXofHRLoNfHv/3q7yK7N2ABjWn3o
l4YKAgJgddjd3NdA/IQ080E8nUYJ0WNxiIMwWwCA8Atk7a0pOQ6e+AL223Euq3rV
t4BbAGV9V3jV1EM3j2JEKnRQH3lRv7U8jKH//QAFdoPtBcmcyhG+zy80weUcDxb4
5AWtuD2TF8oEMOAazEUlN7DPW7rHwUYC00nIrANCNkk287adifMWjgVYZyKR1b8V
coSnIBi4cre5pc5A9XhL9w2b1bFArBW1TBVNvpBHwP67rKIUCO8m/xjcljMmcltA
5JnL6sxQyoLrV4eKjIodr2DTOSsC7f6wKRrpfXrd4MibTxlusN2s7Mi0fBPTIsZh
nac56OsFkpCDxtvgFDV6V0wvWZPX1nhPWHu3SnBSPub4cX8Zlwd2nEXNOerp8OaK
PyHxe8vbulcmkVujzmaLoYJoScdLOFhSgfA9G5Ve7UkAEASAvOg3Gr4cda93ckAR
40XpkqoA2v7uiWVfyvrxrqJrvZAxnOCc0maqWh7SIr+V//GN21svTRepYX1OHwNY
New1rRhufbq1VXHNz9pERufXpXCkdtYlFJwR2jHoRUd2qFiWiT+cAsaWfmASifrG
Jp5hkYPheIjABlSw5sCpN3Eii+WpD2vev8+CH717P38jzqMGpasr1CX1kpwsm5bK
Eoc+aZrPTYP/ZI/OMOwH/8TD8Pwcf3DPWQaGyeP1rscl6jzaR7ceGMv/mJawy/rc
sWhOqX17et0RuNz5t0eK8IS8fytPaxQ8qZWHlQhmyAnxMaphbLirHyKen34+rM7c
bOGnV/oYmPCC8cKF0BH1JjP65fB46e4MSMZW/dMOBt8A3GUd6sL0v1ocPh+WchIN
iNpCsmNNe1V6zT+5PaScKfHEDycNvZw4UHDuqBNdJub1l+TG0F+xtp2jWlWQmRrI
QsLFDXn/wQNxfVL6dzDi9wzlRe0p1E/lkixfoEFRSVV/9VLHb3ltqKjdifiz1WG7
1d0EomL25BplkOOK4eWEDxxSvDmk/LSIfnVPmB9Q16niPefQakwBU/kXW+sksy1q
fWTRNidsknAAnb84n2p3VZKoyCg7aSvIReC7rtO0oFXVmkI44t7aInpIpz8OlnyM
r8QT+3SSTLnqKzE7Uq8HogMEtsZunoKS2HydMi7/f+KdzAkMd017CEjJmPUjloCQ
Xr+9AovHC/BUtzDlgK/DvIoEC+qCHFsoq5AtHlmQ3t1qKHbkiPE5Ro1soNvPN+iN
oCzhSLRwl/VpFHtQ5riwpTKPzmaL9lQ0L90INHFEcSMQ+U9GLSJZDVpREdRtIviW
+c0B6cn+fCvgUVolsyM+O9t/4UAp8gyLUHBSMDArYCpnxrXh0Yd81cV3M7HYAmSI
qgQngFL7fZBTKOmcX14Zr0ICkGG42iX8NP2QE31wixhdQDDErdzIXLGZBscRFgyM
FhZjXIG0Q7o2c92Wdws8+LnWNcRJzK98z/AyxsluJ0T8JTGnmTh+NXSIVfZQ1P8A
XS4IQUSICgOkuazvP3iZvM+8OCGT8qCA8JJnOKmkibJnxfh7FSn5MQRI9s48m8GD
W7PyiheZb+v4/Yz5yDrHzWIwgaJoDIEAFSIt9jQuNbdxhLVMyB2x9rNApFFfyYAE
ITV8wj3KApDRB/Yc5KtNcHFSvA8PuzzaHnl3iS61xZlQ88h9vHlTXPwdmEToS3Fa
B6LoeNigP1h8Zfbi25zhMwp4A55L/LPWvk9VxWvheKgP6mjC78HZArSJlabruB6z
1UeyaoPxhkpoU1KKUjFuBVXLDls4Tk8zixUPoO3sF72FlNQu7SsNQFvOETeU8i7o
EArPlKmW5/u3J0InTwxLmT/RRKjmvIERd2iTPX0eYnOEkxljRzIIRVCJG52gUiDh
HD9MNDZalG7EkanguxP3Jz0Vn5++zIttSE2Y7vA1W8/Kh0Y+f2m55Llk7WAeRUqv
D81Yr8NyVRe4q5PZJjc3ohJHfiSB6YjUCCa+8QXup2H4Zz/7S+FlSZAUnpGTG/F1
GtT8U9yWWLvMuLtTBb1AdpF6I+p47kEhcuoIXcLx0BGh3h3sj+CIZ0440euJWdYy
9B8eavPUWRSlZtwilDSpXD7wFZAayH+L/2/0KtCLA+U00891diP3srkBJezZQgQF
qw6TTlzh6RNgkXXQbW5fNUrQ1GNCOFg9wpoEDF/dz8Og8pHd5nFxijT64UNW8Ywh
jyeby9wKTFzH1loVOoAXibsp62+Qx1R0oXvo6blKhmThp84OljYG82Km/rVWN1Xn
46FyeZSXhg2J2G/dyFYrr6o/cFKaRaZfOL9ylptVfrmvGQIBE7YvfOPy9tH+KShL
1S1o0RUN+xlnOcZWvmpkJMSRJxO3EfLon+/pPLEvuOxkfOAdgSOipmBAs9Exn05N
VNIw1excQe/IsywW8H5C77hUNT3kgJNvlHDjjwPjwwbTrPJwkxW88P8mckNneNfN
tJcszbZ2kuhpu6EZAW+lrotrbpXy+TPBJ9PZG48YRsXhHNucAjGChHgefASvFRVO
2u+eC+TRgesqNztSrrGC0BBT4HKl0xarclXsjPsDMWCpvQcZBPMt4BEqa9eN13Jx
Wzz04rYvT7HodfX9JcIhrzLdIRHzfjVDzVmteRa1mgDIGu4UoOpNXEYdQ1xG5LC7
klc/MNNBXPrJ+o2ykxbTomwI0umzSFbrp7GfgzTei30K78R5hOGYZd+4LV9gEc1h
TrxOxejJgMtfG0TrveG82LAbaUW8lapvXquG/cO7SaStu5w0Zt4WIJHgeB/0oa1A
tI9l1v4OHGutdFJzYPSg8T1aSiDnUhu4nrNQT45R2I9r/dsRmqgGjr7D8Co6dqUO
x9h1s7+Kr9dCVdlTqRCMBzJZoz7BypU/yLr1msSflLlZ4+Lq6lZLZqeUm3MgLUkt
MvoHCR8jkpK9GYLt9VFNWltaulEfOPXQKkmqgbz2mH9LrrWc9BQfiZAckOIqaw6R
Qh9gs6HWjLxGArwcYpmUgDaa92hUw2Ae4iIUZ2/7qTvk2PGxW1e4twpm7ez+24HK
PheWBn3DTxQhb1S+artgvfhZrLZkjgq5ZNFPt0VohtgxkipQezC+Sf7dlxhykVXH
7WP3/GSefzN4ffTcgw1s6ZkQk4ZGFD5pdrQlnAryTtnuPQ0G+8T1tqjxFQiGsp9+
Fnf4vY3m5bHJwQ0tMhxKI6hZhrgQYw5q07Ke9VFbi7rTP56dsEOZTzu7k7csER/0
1dLTUHb4n9JZ200NaRhuxhVvrAGsFmzUKEU0Grc7ShZNoLrtr5008x2plmghk06Z
6EOito+MSR+gCffYB61z4br2raJVE+9WEu1YFbT7MYpVG304ujNI3Wk3s+Py+6dn
LQgG52lKBEvhKEsfNCTT8gQM/HlcGoicbYwHNYRSkOZwDp06BN5vMpbFhn6KtYMh
J21nlZsLAQcGuIWSpjlsHRs6mE0feoum0P8/jye/D/J92Cm2ocL1nM4xBje4Mf1H
gYkT4UMVe3FCcmNSbJpY6omzPnru/qm/ExOPGxk2Umvoe1J3NAg5+hEwfNghmQla
k99nYw8uIy+Cygjg3vFESFU62uV1PHnx8UdQnhFyLQYBIB3bSS6BeooOMsS60zzp
/Vth/pNNEHmCdZAHzJQfzDgnzwC/ESDOJ04rKyCFEhRsPUPM7nF0RNfZCrCWd1y2
2mbZgrDeRxlQB/+HlY86EJGfj+bKNdTJM2l+16FHQMhIQr5ZDBwKqpo834urTUYK
QNnG1KMg1gPU3JDpfHzBL29xozOHn6Z/xhQUpPCYgWRVzLyy4Ra/T3zwzcYyamVQ
L2Ns+p2CBSe28CMaBGMMuJQby2mUfFym8SDoE/vOgGzUw3iAH0BjwNamIXwUgs6W
zITyHQV2niBhYNnEmWxMNIWmfRdq5IGcsD9tY55991etmxFcrgFIHr7QWkGb8Kgp
KCqspifGr2Fhp+8+xRSpCAqoxJteuf5P0dfCuw3dzpC6/ZQWogOX94GKZqpj2xk1
Qq24/nKbAfPLjV29oPnXQcpSnBVNvd31GXv+3nB1UKmt9azg9E3ZUSzbUn0B/qde
pJVvgfI4hWt4pQJ48LA6tL+Q+RZggnQOqOQwEGbtItB0hWvND8h39huUSfsCPyT2
1oqgublSBekIuTTqrySx+JkhEw2EY9FjZn/aZsKfGOjCaVIhkjA2GWQjq0q7R9tO
vbUWcaF10OzN9CjzIZrZsDT7ZU2nyS5ngU7xOu2QV7f2qa3Nv6xvaptGZtSLQ02v
mUQCX2A5UqXh6a1CwEOy0TIhW64zeQBB0ECTaiqxfKY0PPOrVdz0SQvM7gFpKGIQ
p9E9eYu1m/dscnpbGTDUWofw7YrCvt9M+ZfR9Q22uzV4U687TXnSi4tD1QV+jvjC
LqdniB1+1wb4OKgtTFPz/aOoaA/Ugt273a7+gQ5GnoZ5mGdILMGIXXRE0XVyUKTv
NuGaa8N0230jJhzQi9I2Ypfkk52/ehOs7K2Kfmd1t+jDgMfHlszABNCvDoMMPHM/
w1HJtP1Uiq/UgddFHj+hb1DqcWmx52ZLLY6owia8IOi1fPk3znmBK8ApJRwPbgRe
ZEW5KlvEHwGgipZhD4PBFkNUr3wpil7mQXZPiBbCYLFuA6uT2t/k+isFJhT2t/cY
/mU1Iflc4atJ+RXHaalqI+geJNDmDjR6buX6KRSXcsYlcQki8Ss3e0iTyyCwA3Fw
hzAJCc8SvotsXDYDACPNOYS1Rqs8Mh866ofAIhpOrGhTC0aUaBILZcXa0tlQZRxK
q08mPsgNcg4kYzVS6UQQteyYw5z76lOwg5NL4Ku/xBAxr25orZsfm5fgN35wjP7j
Lm4tExsI4SovivuoIPTiPRm6JbIIavUTAVMuUZBnHGw5RT/C9jkq/itLwIcD6nt4
T9ImfE3gJo2FxMOmOCrk6spAg8V+ZkPf+Whke4OqQMO51mRpJuN9NEJMz03jeoUh
R1fkPJmyA1Gmi1lqeTKWhAP64zbaLR2/aLaLZ5h0Ktw1oJdsn5VTZFjIT/L4Uj6Q
F9ipmSwiCI41gFWsV09HUSCNNffIbkdv23xLQ97gQWajHboOOWkCUn2BvyiB8r69
1z4PSDuARB8iMMCFVJu+c0ZjaI0JOWO2DXhRIfEYgfb2Pyf0O/ruB0HUsuO0bL/z
5wP7eeFOkc03Fjpnngaw27r5Zr91KqQVCjVxAwNwafVC2TWkA/jE1n9iqaC4TpYp
oCGSjUu+Z/EgLJlGkMAm1SZCuGLfWU9Rwffnn4aNfOoElR9tWbGG3XHVdN5nquuG
/gD90PpaMvdawN5igXI0GyzFTjLTLFFeuOYNZJATi7fU7jUuzLB9+/Knas2cR2QO
n1gNx6StFmm+6zUpaZb3nWIGeUesiG0/4+Wy17jP9NFyd0/MdOAsN5Abb+I1FveX
wU9NOCqVBgrhgTKa152VYaPsOVvgah9RY2C7fS9VcDoRVzuG3SGJkhsFn9BY/n++
wrf/jWT/NbGS51qaJxGjyWerrJ8eKrJ42rE9HPZmdc54qhltQ1Ep++SqMJakf69F
Tgig1RXwIaWzTdnEwp9zDrYES/QNMdtLxCmuAZjneyOJ789BlFomq4YhKTD/uqd2
RgkHisDo4HLTLVUlTbttE0j1fyZvKZk9F4zLF+RWJme8r9kHFz4fovzhUxjOs01K
+CcsIrO1px+cs+FJFKaDJOc/kZJJuJ6TjACugNb3KoeDQhv14XmgVH0F2O+I86jG
6D5yi3dhZx8Q1F+2jhShhfoYz7tDrvhhMcn60lwTdl9QTOcCa+IL/lqpaKs5I/3r
cynEYujv+VvtAbzFUzJ0W+f3ja9hIhyCL7ZYRSTb7to3IxsiZ3CkcN3Hq94MYcv8
zMOvXmrstzVA8SF1Tm6jpthl6ZHqXoE8YhFdQg+ktRxlry9KL/PJ+008k+W7CFYD
L37re+npuGwoY6zzsCuwH1B1a0MOVhIKxld+nLd9Eiq+uUD4o11amsYvxU38qdVC
qE0MMv0tGfF+rOebBI+8fu+Sl2L69pSy5R6Jgw4n9q5S7gfHYCzYWkB5fYRS+06P
4Qv5tylmEk2ynzdPEp9CulxdJh9Cx+NFJIfaufX9dcIYw4KXBxiaVO/ht2YdOCJE
syP9wH+WaZgukJfxtnQKVRJ0EC+aHxM6vdRlw5ESeIwcnxB3xPcObgxFSDpN7tDX
zzCAmnTdLtqbfB8ZSWpWtnFtMHG5MqsEIcLwO7fDCeP2LyU+cJFKah8o6giYNHxp
BqoM5BRj4H8NylX5oSEX2M6u8fyeUo+ZqjGEB7P1iC9s5f14bWiiEawEYJPhS5Ml
oGwh3cGPRsSzcVLaM6gu9aUvNSUttZ8JH5Fj0dFmw0LBJTCpS+2prh016qDPMJ68
shVf87B7eSAD3DlEvnFqNGEl4n1/J0MH70fEfpyQu0p5ZVfkqpc+iei4biJ9aZhC
LpWEh1nqvLpwuZ47ZAjGfu/lX02TzWeehePwZr6HOtQFhGfsOWJLKZAIFkO7ILLd
u0C//E3WbHU2vIfkywtFsqtInSCbqR+RT2aplhpyMbo2u7y3aY7qNCwfUAquL0ME
UHhUTXaE648302UeA3UiHzB9FaExw3W8QmVilEv414odDr2Qf3oT7EUaZXZ8UdQg
4cW7RU6aAsrHfj+TNAJ1ABuiWx2HNcHzZq3BZkRwlZE/XdxxE0xYmcqVGnDuaqWS
5CCF5M7uZZQ4GfefwD411zGJL+bCcZ+4RnSeCI1xp/AI12BtpklnijsiUBl9EFpR
T0nq8RBQHG5I2R/BRbSYUQJUxdPJXfZ44zpO8gfsHly4UA8eC1VZPRswVgOqEcwA
5tCetvoFAzMt8wvrm6Onx1PSX7CEFRaSb1yOR1w4NYFcxSX9fvplAYhHWvKYblCZ
JbPmZHLJf0rB1l27Unw4m5ublAOU/kuaLaKJZvxP3h7J91TI3rb5FSjL0FG5tM5N
rcOtiNyGjms8WMQ24JI0Tq5Fcy7bxAbOUFhKli4bMOVO0oCXUKLaJfbWcQ1SFRpM
dRjsp1KN2Juy96CIJOp5vecUQdN0FnRZ/8qODBQspRp1CH3s/iK7uJSm+NGEDvVO
fSxUV2kxxdGz005XSKnSxUWI4dlmme3CUJrkGqLsYZQrJ46zbDn/GEhi+aZBGyua
7jbv4c6TYNRC1ViCPiN2Y7as51fOU57kV4GZl9CD1fJlEKTmX4zG4RwCfE1//f4Q
V6ilt4SZOTuLHVq0MHdBs3VUPbJTGtJvb4/qqJ7NTLd9nNR6/O47ZNaoBxp/9cv9
tab+wGlZUlRex+K0Y2cXCXihkdKkDRLtnxI0dZA/Bcdl42VJu+BAApfNYLi14hg0
CF7+c39kLUXKi3+CqWjFZrA/AfbF83yX+wXY+4Gc458uPrg9zYKCLNtpnwECcES7
6IwJ+Gxkav8OlXgfThxt4gMU3gPTXBw2dREzPvn/5fpvtSmyEKMz0RGZa1XpcGKP
wS2Nk6Nfo3nqsykqGjwDTVEsqabZUNhRcdmal8+9biQqMlTfnroYQEdBSqBHd+Pn
yn1KF2L7u1KFvwdfdoKc10q4pMg23/nSfBgg02NGGRqJJ7IraiO7gZkB3D4LvBI+
dpCN6FgeCSE47T3UQc0Hf3ACkBzGllOILm/ADrrj7J+zeKE2GT+xA/128IsnWL1e
zu/xDhGhvcpb74HAiFCa4XTtqdvltFcNxbIqAmJHkb0P/aoYRvJ9owqVosQg/tAy
rhgjJeaBBSmjRUAFgKhDo18IH60K0efFSG08tstRp50m465eqo+qpcQ6DC8dq+9r
aF+QgMSK0/TaU6E88EihQjLgQqnYiO1knO+mZQibGiCgMPM87wTQZJ0dmU8+qfaf
+WC6d4hs4mUYGR+WRgo8aqBsbSixcwu0QfSG6ENBgqPlhs028JbPm7SlzqSJnmWa
6pQoxllj79czlZaBxjAf5kVWEVdHee1CXUxmeBc0jjzp1R3BkJ2kWu0oISO3szl1
jwDOrB8W2xRQeQrq3jhuacAGoQbiaLUVL03tJc+M6pTw+052sd7Vxqp0/sr1mHT+
mh19f3kD2jlqSQ5Jv4zPWyrR7mS155j7TVqI0DpwAE5t2tHB/IuoyXBzWF8zD576
kRL/fvcaFgTWO23NCzy2O0/pRejaqQvP/yA8wTAVBvUQTnHuoxDohL1eyyrrOX8P
z519MwGF1PJFRxRUcmVOELRgCPiF09xzCv81Kb5BrCjOqjIXQUHi7ls4QEzWO7jv
0QTj346kFw2uAv7FVNumbKiDSGdV19IFDQE0spRvXCImR3iJX7fs3yy0whCTe6cx
ToSg86spZJbW2pUVtS7rGCV0HMrHU3j6IoTZ2gfZOFBPGGwJR54Ed2pDqTqtywtE
SrzVISir+0F+tNgSQSkYODSS5z4C47eKcIBakY4xu3b0AqBEhNbBPVHfjRhbT+mE
COav9hQH+bNbIJyqx0z/CFCHVToB7h2Rwno3sjrtSoShwGC0SnS+T6kA/HRnsZou
8mHzsEbwudTsw/DPr9/OvIFQ+5tDBKa3wBMtuSz7hLzRzJu6dG9lXy3V7vWP6RgA
29ZEhB3ekdrS/DCP9b8ZY83rhKY3Stg2PPdRfIY8lYUWyeZxEwuvmdYpKWySWQKp
rOFPlvMk/Rl/Xs2ugHbolperI1PQGP3oq4F+gPIpQ5FY3hW16VMwJ3lacchl24k2
ARYKDVW2/aADpYLJZP8UxRjYvB9oOG5Oyfni3QHD4AYy1wkbTOFsIst72kk1ICle
KOsKeN9/l50jqjw2BHW3r1AX+sadIKEUGTn4cZrPAiR5OEf02scpeeIRKJubRDkg
W3UwiwAanyFeZr3MZvOlAMgH3Oa2gBp4EvBNbcXQWushqafbPhS9zEaxzqu3uxuN
LJ6GKE52sMekQE5Kyv67vXFRiPN2DExY6Q2+k1msumw4+k1rfnCloS2FSVpa4hJg
GKE3j+MHH8iPenFuYXrpWN3pyCo3TxrW+ExF7jAkAwlJ7xgHelKBZJk3X1hEr3fP
K98YBGGXDPIEaa4NxUqfPkOhSyQ18vcrY43XSQxtNj7QIJ6aiwoDM2AABWpS4D/u
GZPI1HEWxVIhMIXrubjwEkdE99YMS1pvWXpn8zvcXD8U5y84lC6b/fgW3p4ZUKYL
aSZ6z832a2x/7oog6VtbqBmB5TJYZCYpEXAlPMi0VDlgcj3WXyjiKKmijOAlMXSQ
gNYwYEX34YSgTHy6yeC/2Nu3k70DGlRizYQBzCqKCchH36Ff+YgyIkZBbfvP+14c
JINirBejQsiaO3u6rWYJF6vz3yyg/V/deHnYhbr8Y9TB4HUW+KTYq9xxmaYgN6Wo
Qdk3Gl6IbQGh2omAMb1CGyY/xRkTw3ROx0DT6rKqFvok7vt0+tgTsefP5becy/cv
r9lF0v7pNZ8EOvVeLQL15a1Faf+FEUY0aHkcbkJnyOw7Pw0dRllnKHQP6+OXxP26
zpvwt67MXkBD+gTtB0+S3cJdiFXAriENYMQPxPsxxu0ba8bbYONpsma41h8W+hJa
2I9/gEV9Iq0Jgf02YNVc5MnnKQipV+dVac7m7dKZO9YN/hbgA8QCc06yzioVQtqB
acM4cWmLlzUrm9u+E6vYthbRpKMB4ZLHKrpp2MM2ZgaeIUoPLinhOOuOlIPgSIUh
rRr8AWWHkmz4UNwLKV7oR0ppYncGgQo0aeQjOmn7qm2Yw57aIb2fYhlxd9qieKl1
G3Jt+fDLgJV0i7Gpqmi8uXjnK5DyHqrukPD/Eo83YhqZLmq1jivmhT1nLu4XGG/Q
FDuQq7So8AnDkvmhYx3zypXkxpQ4eiDT/Ucah1/BIJ6EV8FmpUowE1GhiJVO/W67
ypMsaCXef4tiCHAjBT39mbi0tlG6nQWF4MxAsXNRdD6lopQkkf8IRgEGE1guS8hz
KSXuGRO+2AnkcEctBNkwEYXt/3XJT5tDP8pK9+5TQ+aUlQjGejs/q++hxbPTU2x9
DT+Vr+9/Ibk0LSJptCwQinkk+mEgKqi6D8b5AMoNyF54VhcHu1vIcSx8cK7HVVNX
lNJpAWaUM4XgZFsfvEJAYMYMxE5nU4sjFJ9DS3DTLfLVWPzUdUrsIxCkCis7Tr16
WHslEW0cvMpxPfrlvyzoudGdfrBsZZ7Wb2DIR6ufRI24UzZx9yBct/Pa5STJ/NbJ
xDQuoDnneeNx97KNSjKils+FPin9sU8dysluV7GeyxQp8dFFulw6jqR52BKILkpp
Wxs9QhGx0elbr3ix7mHXp4WZfD+xyFuutN9faVK39sJJC0OVOvfqpHPOAOw+j3nq
nNca24syoUkWzh4rySytiK91IBcOmeFspa2G0yOgOgphTaVnA/pwYPz26sGIRz4D
mcbd1rRxlfj8l6nreciz1rBwzwrnIDz0zUo4XboylctK3qnizg/fM6wzKsKeWxmn
x75feQUf8n7Ui60gRhsbv9HtvB7EePf4TmOSZ3yowweBmOrwak3phA1pGw7zzVBN
PNSKPJOG19Arw30u1rnyj32yic/45NZwdvJ48ajE5/8kf3TkEhnkUZSk6FjJ4p0O
kVx+8F6Ip9C5OMHAslBUc4HHjeLoHdr1CpCnTN0bvvHi/UaLQuePgZzi0IXDq1SX
T6cWcBOdYobSIHw9b54Sfn0gdz9lwW3inFere7BmuYk5Am0LiYo9YMFP7UNytBQO
3OAH0FCuTsa2bL0wAWQ7ARs5Pafb4TiQDmgBRev4VK8TjiiWi1ZJnzffDoEGXFo7
Y+joQFgvXdc6j5Lsz/wWccAeK9f58PZw2mcLTbQ2YwEOUo0OfhYnNTsZxFr2ZEda
YZ7o4XlxQp8OiPlZEEBAKw6g8mFAqX1cgPJELNOK3U5xvEh4O0x9u+cT3L4dbwiV
vZJSc8JXux7Sczwc5ATvceoOtmvgpUbGMxtdAx+PSe2bN1vlezvz+ejvVaZsfdqY
sm3V40kuM5w+EY0/iuMAIBmNL+JLEXoDtW6aArnx1JCpcKrZ3LPauG+fxxruT7Vz
Y4IRT96FPqFzNL5sZmN0WuFrEys0hllmj2dx0QWW6Vjwy3Clh00iTwlXLkwEMWBR
gDxhG5bex7vZDhzm+FbXU+Ha6LGNaJMHIA82rFeqqptdHOeDXQ927tS2voiY0Fd0
7R/5WVgO/nWKy9Pq1x4pt7VAn5nueg1jMjyFxsd1cK7UKmCWy281rOiKMPt42ndz
EffJuzLJRejdGiTD432Oj6WS9bgmvL/NZVQXThHLNquB2c1RiwsCV/WlaB0eaE3h
n2Vrk1Ekdj5nikfS4IV/86vdix71a1nvB7oebPbvddEw/2iGwjZsSwjUP2oAdm7w
GXaAGEAQdsrx8DVdH19K8Qn7YTypTdtro0kQv6RnDrL1OvcHfR8WJw5RNS4GF5tM
BZowz9bcHg0GwymwAeRDk+FX1YyJVZJhS04vCeA4I7WgT2NlZXvFRiK5yE1DXhXM
ojBrYKQs/XA1iXMIvnL6xZ+467phhc+C6VvoFKaQ0YUHmJr60ttdEEeSw1gvYPg0
epYrLR/yQCzB27XlZRcS1w5iNXgGARFlolE/OrLbldbag/5tTV2Mn3cFnburSXhH
rR4m/7gKQXlHQzvlhdfqFD7ckrxkPER6HCEfDmNMMLBtNfjEiJSFY85Qq5Ni2UMZ
tRzbhVR2VDAlm3OHW6UYMrxAs7A04DyRJFlEH/1Ru18RvqBNDtMTUCQi8BO4jyUS
E1F9A1KGAE+9Jqp2N2FgEoc0OA8MT/AcafB7OMB0ktdyelmK8P+00E7sEvaiUJcr
I6jI2JP4sSkrb+30P9bF14Ta/VqVPBXHm/TjY5IVN3drEMbwuUv/RaYOW9OitiCr
f5FBFj2WS9wetFtldPy6WT4jWC6djJ1QqM/4XhPln2C4qk7CVP11LI9LU9snXfpC
qecO+AhN7DbgZXA1TQcWsFaB3PfOaLWjvElSqnQE6VtxVrrmLEQzhsTa5Iajp+re
e1EahCKy57UMTaUqGsJHxtiHbWb5Qy7rVdyJ/kxW1GqOKH++B5OUL6VPPRsYvzQD
KGRrfHAllEWST1irBL6UPqyT4U8iVOCYp3RPvCyLnujYgB1NqbJESutAgFYceaPo
QaaXJJ9La+BvTFBL71LdBRieCJu2AQsroo2AMFEcOAf+JMn7Brya8UdLklOCyE5m
sQ35OkCr9vvoB20MJoLnyjJT4W54eusVxkzGcbEXOveoJsD+Y9yUj5IYk6MxFpdk
+c/Ikrskc4pWzxSdlnUGnBmPxdjYHBSUlj5e4sKg6heWrzgbFNOxbt8DYBf5jgAB
aGvx/yl4PZeOmkPhh0Vq91DjPUUf83impFHhwU/+lw4YKKjckAmv0REuDY2QGbtO
1UIo9tHEPgE8pfBLXRQAKGLcmcKBGx6pflfDCtRUUf0Q+PRiJHp6717piVMHm3f5
P9soNM/CepIBn5HaWq3VW6iWXw9Pklms6QiNGJ1q/hdJpcqxIezRFsNO02WzI7Jg
i0w/TX+EyGD+WXukqQ8Jbol80DxXrOe9tmbasMKNleTEmiAEtBufvUPWQA3zCBA4
qqc83tD2VPcKZ5H69RXgFCxmzrLSCK0xj9ogNk4r6UXOu5ZDzYN2KHUKKcbdDn4+
cR9XRHGKSWmpO1WNhl8MFlXn5jY66m1lqR3pAcPittsiTJ5kN3tZD8SdnZZn3Em2
E1+fmIPSsKdv4yBn5WBroFY80TX6/rXP4z2gnXef94vSvy+7hLB5Bky1Gi7349++
2fM8/SRizXZoHdW1QchmLiN+K20RFpHlSH4kPK9ugVPljaCxqU2qA/1g7CqVnEjZ
czmN0e7fdzTanysslM9l3+fPEz9aLRtgRv4BUFqyNaTc21wxEsOHAVDLJnZCUFvI
6H7iyUzXRhf2jvwd+AyYGxPA17dZcrSZdLmXWejYCSVbxp+OBLQxyhugrJB7+6zC
dwDgfbd8XbvL89v4EtXd7J7qhGf9AmhHL7STp5ThRJaJoxJ1u9nzt2waOIXYxIwc
YC1+D+pjswdjfeKv2soUgGqIjSFPBBQmK2MvoUUm7Gu02HMQiD0lhlPR5ZRuwkdt
kozD5nAP8osG3zYO+jMVmGrXzGmwN4KBRyypUenOv5PBIpNuqu/meJET2NLTj7qV
cV3nJ0fxt8Qa1ppXFxicZgtTqLhazqCFD+A1WXPq9tXYz407mK8jPewFfJBE4o55
upG8+iB0DrigC/xWb2bOIhQhh61tNesOXeMKQy3MMSSZxeGKPeMnNmnuqWi4q3zZ
c+zVgXtMryw9AFUjQ+a+s0Ce5w6Ic64rIjIyx/MqsPlIPc1PAI/oKMtKC8n4brbz
8hUNFWWUw0o22ZXs6005NHx1nsgVUmQpVYB6G6udWdIYNMC/MFJDxJL1zACyvgyp
+9yHgO+p2VT3y7HiMLs6x5+c22ALJ6LMrRh99xfpTmtP75nT1IXav/b5my2bQ8Ov
k9iDqLRQTwW3cKVcac8/uk8cLNIa3Pld4QGB1G/7ZG1o89ZGYqmgIbj7FMEBhRcH
ivhWckeZwUaGSh7si9p4w3salgpIC7vwLXoEFENuR2SAgwqA45A1sCBeTKNe4wPj
jeQgpGm2aT0fQAqqwteuqSAQo0lkbQRp8MT7TkNZcrZsZY1UFvPx93nNdp18d4ki
JG9AZTdlaJ8rEkmkf8qGUNb+PFCsZD6sXpkU+b/yGLrdw8R1SAfhqp5AQ/9HO9eX
dICZQ/nYUK74i6QV/noVLcujpALaPKHg4m7SroT25mDlF9G+w2jxqLla3ox6Zz7L
PYmelW27kVGR7GxjAl23t/0Fq7Yb6IgmdNG13+cGzY3tdiCVNza+s/kGYmZ8N4FA
hnMdefXXcQuZZe3rU1qxha+N/Xe9tDubaJ4vFR3zR2x1Yjq7hJ9Jfg4PHOM0VMPi
Eh4qzGaH3ggUiovMTEGyfXg1sEr2QY6umrUgvUlpLQVQsP2S0ogjNa9VA8mPYYZA
ctJ/gXB/yEyPf96dS9RjedvsF0qX0vNDmtmbAhW4+Hd5Ip3QxarqPCN1ICEheVgY
qk5iH0NL5rX6+WUmQwyoKKQf8w8cc0qEIYgBfTMyRSeuiLT2OxfgYxpQHuvQjf0w
JKBvo3BLn3WJ152jmzypiaLrPcRfPCpMDPuWCYuUSgB52hPKR5VMnQwfitwY5baQ
YWj49xWQPeM5aCSEv4df7MCkaLbck7pAPmRZ8nLYbiUkCfkU6fGALPAcGd5MixtJ
0HTuNqGb/b5VFxVmDZhbMa/0AVRbzQdkjp140VXmUAjnDD0zbRujk4+fDBg9Suer
9Ps1BjxAceoNqmaWdXTQhakppn6zJmUuImodIur5TeINEd1pOqXqzOw6lpj2C4Tt
dHA3bDxwJpL7EvlW4KLL8ATIJQAnXdBUqa2jWXaTfPUp4v3Ja8ev3OqcgSiwO0sH
TLxSWwbkfW9ZCeTII8epUuW8aZAc+IzWItCvgVO2HSESmupfjz+4PrsX/qbUbrcu
E9jqgh57HtGXidsjLcL70XeeijIMBfMSV4qpp6YcOr08JxvG31A/18onXAltgbah
IJeqxi/TwbI0oAoKT4uyYXnDaB7GAKNy7MBuZhhFYyYYZkWZuSv38LB7FjTf9twh
e7MrzARp3UKif6LpBrAEtjkbdrU/wy9BM7Ox5JR0mExDgNrD/O2ET0gSuIdt2Rjo
sWavLd5bIQSMfylzWC1gyw/zr8RqxebIcZK8WPnetAR8wb13FnEt8lbiIj6hvCjH
OJ7z2aHUZQJJs9ypQ13Ff7i6koJdx77FhdlwuTs5ghvqRzMkS1bUSmoKQ7/31N/f
3oKk4izTICSjPhCFB1SUAg5ZLx39oh0CeLw4u79rS38CwHCdLk+U7RupX9wcOR5N
wM0jhUrc47mEz952tZXnfu3Z8N22r4Q7W5g3sPj0l0A54Tgz/vkKQRzgs3nK/Dw+
lIFUpRhFfcnB8Sjlhm8JGtHYockbZpK8bytJqoco+l+oJ6NQQx8ElX2eVuApeZQI
eTW4B+DEcmVrLmyqs01qD1PctjsJ9qFuk6JBY8BSegevGdaW7jF/wl0tOfvQmELV
HLN5XubXuYBKKZgY9X2txPNfPfkv8fXzqfG7ZsdqQBInuFFcx2gjKRoheiYEITHN
2EghkJzWBrL0KpgSB1YUycF9wZ2/unBWRMxKv1OqymRXg2Q4ISD1aZa8Ppd8JKew
iqzVSkxNqoH9a3VVhUnUTliB8GHk2H+dc+7By+yiUAhUlrwkI34Ek4DSXi/omvJX
o8kht8iJDl6Vh3uuoJ+ZPP+gU8+aJOv0ZuzfDaECDBtrA0YG53QvBKVWlzIoUYLz
sS70SE6TUhwd+3fjgxVc6K2k7iBHsKdy53jbJaWtu1evDfpmix3+Zpv6hQBHFcZd
VKkJks7g6rfU7WDR8yMUBXllQFLyg1KM64ya521ezl7ElVPmECEBNg48p10SiALh
54ZMMuPYVYbAEBoY/DmxpMahpGg7xDtELUdqXKMh+4i9q78iFE6fc6bhM/EHhI6d
AAdnYPHs8ByTMb3f7GC05ny8+hgzCrYybQ8DRZAo/Oig4fOEoXaFFFSyxxEoD2YS
CKg96u0a/cTU8YpeqUeeKkxXYg8n+tKbo7Hg2pVUQUPBTmkPUc2b3wqAaLS+07cd
53kykzVlo3xPUO7HyoLsnFDmhlsTdouh4F/ZGPJtDdPBN88vMeiPYMMeZ6aOYl7G
NuNB7hDvRd7UeRIxR7IldkADTk+kZiY9lR7h+Mt4IZTTuASFKn9qO7jM0xwJQBNU
c6Vg4YmOBUpp67afpkNgbovPTPDORkvfR4HjrirY+4cdfUTul7wTutClxWvJpyim
hKli0ZpaU0kSbjf+le0EAHCvrrq4/Vc5XYUdGG2bqnN6anr96TgQMXVZBUsditKE
cMeNkBl+4UthI/xrut+V8V8Do7YiZ6ZZdbpWnN6n/bAIJumuSfir3FZuQDcjM6qk
+l5NKdCbDOimD5yCgktMuO+QKwLDE8pZ+8QPFnFYfrEJg+ulJMAePCGTHnK3NMPR
76eJvqOAuZP7SBLqDJwVoVNu4YaC61MTMwEypI4NOpwylvpymPHm3koMGAE4hgRr
LQECBtJJ4LyDYMtDu+cSk4zKAOVhbjr57hZMEk+1TOEH0oSvdCDmAKUPzCBYBoGS
d5DTgGaLfr2BNxG03ezoRgYeC0RJOtA/F42blkWANON7n77NMkZmO8PbubeasUSc
OAtHldnRxyc6WlN0Ti+YmibtpibZVWSfdZ0ne+bY34cA8CyF2YXDSKX5x0Xa44tA
WnlqxO7B8M/J2bpkTlL//ObWAfkYVWSd6/2+/VPdX5DCrTKKA9PnKBIVzuveZxd4
6Hb4yXEMk+ftiZ3rGwSr2QFXD1k1qZBVALedm/wspqnfW4M4R5ng1BdngQyYIlcE
L/9fVMI9QIUDYICokKgOTDHgB7cfFAjE+x5JoK0GZPSR5aQ9SgsTj6MaBN1cVTc7
6QSDEuoSbkbEM6d9QVoUz+7/1EyfNcBKNYb1GZAPYj54N33BSK8x41sogflWa1ET
ncw/4p/zPmpbkXUBNh6XpDXTxze0dkikjMmRKx0BuwxkrxvQPthzhVneJwbPHqko
NDEtQH9xfMkQenGa+S3n1vzbPzzHROIOQNJ/YW42pMSWXVWXg9FNsG4/7Dhp0ByL
QnnrB4AcJ25HBvDJCpegOOqEMhsDfIuzLe02RP4NGYfFzyQPIcnVh5ojRT53vweR
Gowlxq8wjUtfNHS3KkZ+EHenlhkuCXeXldZvLTr332gq4K7nCvRz7jiAve3cN1L7
0drB7T7W86dLji4F35fDrCVoAod8bscaDbyPxJsSjkGKzs1XBHyhkVHufJ+44ngO
CjKGXlSOzg4cETeHC8gi0kqRdSmG1GHVuSNt1s56kvO9X4NJGYvN/VMk5C09h69k
9/ls1TLltP/Ed+GxQsK1iClynJ73tKDFOd9SnwSCJqGAhsKFvOh/3SoOrC+yWS0+
IDdwKOsO2ayE9znJ76NheJUHsLRKymOGKbaRF03WjVe3dqb2eg1CZkDYZaXIBUSN
ftbpQj4pm6bNIlRq9VDN+QT+6vl7GKXRqJ9Eswo3tyTlT6lKIQJqwtfiiVk0tgtx
j0SihwlqW1VPsosyK9iFku7yMgyey4zBqMww5xXCYljJ+6HQNm8TL8m+k8n9DRq+
DfZe9OO4dI/rO8CXzXiv9L6xbIWUH6fZlnHyY/PaZXSflmLsSpjznB/VR4bOPF5e
vyMOt+/wjXG34SeXSvJQBR4Md6dOZDwZ/1GcgWeb2J1WjHemlOP1k46RHVL8a7JM
OauSEWa+oHB2en0iCxD9DnPF5GD4Xqx/iD4NpeeXHEI8fEPzsSJCnoB9AlyhBnHj
ofPA735DEf20dnl2S2FsV9LdNaLohB/GnfSsw0FiMdUovbjfGFYpsoZ12AHY8Vhe
WnzortEtmwNL03oyb9EcqT0XfxCIfhwYRk63T9q1pWz8MPnQOU1XvHtpEj/ClKEG
e7BdiemlV1Uv117k4zdiUtlu0dhNkQA36qJeaVVXls2QKxb3KjxgOJw5zQMoim9I
oQolc+pH6vN+hWto/gluFfSvfU532x07rPZflehU+tO2FxKXfgZKmSm0YZfArHLV
P0NnLSNeZFpA3OKLuXufEV4p+0zhVPfGf4rpuHXhnxp3SFtU22eFAp8SUR8xGN2x
pf+vr4dYRJms4iFTMYx8eELHWaFcE+QXu+6LZoqkjkcTh+UEeNSl0sP5fel+kTN8
5HRnDAk9aGF+uVa8Rydjs7qDu7ubxYx9Nj3EAHH+UlM3ciWKtpUfL8FwD8RDMHU7
/vrhrGj5/1IjR3kaDtXajz55hfOG/avKxajw5FgcdAZyghB8zebOLBzL601nReYp
DSNlpac9JJHs4WBZHkDbocNml4a/Kok6UVQuARINuQbosyxbPex/LkY6LieLWyUw
JjazIejCpOF64zewan4E9kIxzlIX9cd8tEWGZbp7PCRSiq+VZRz/AkdI9UoTWHN4
Aw5xggt/VA8VJFO6L2ZSoOWIWysrAqagORtB/z1UHReb7EViUY3xN+vvyTk9EM7L
zI2cweWVmfg4DGrluXtHincmJ/YVZaH9RboQ08DhOk2//ML3CiLk9LqUyPG1UkoO
Cwiut8qYLK289kaJ2nFRpC+n+a1E8gHl0/S0KvIoHqvmnNEkR7a+MmvVHL8Eg8Or
PWSC96+5n01IokCeEhtsPLrSPbXnfoUzE+sntoS6zXo3rA0FihuJdiksYe+YV6y4
EIyPGeGQJgGEYCChH5Ne6Nz5/homUr3DuPbWX2ApDS7babTgwUzfDjpBi3afYb81
9ay3C38q3apC/Qj9cnJNA3LUFCofLpD2ZXZ25GzsCPCK0Iz89WT9T5eKXuc/Ty1f
yfDP5v8yDYF3/PjkteOeagDg4ibY3kkaRuz8TBSUDqNfK9z+DbNGfwSk8SstWBdl
wlAHCp0xwkBaRMr8TtnvtZQVXYdVOLvOm8XG+OuH8MZDfFOmt2eofNn2R3N4qi0s
pa/cddGJkNPPH8K048gnsr9IUmlE753MJ8V29ve0YdCI+c2Miv7VrdUsacBcM9of
QNgDbh1IohnE2A9lhnOnX7XWEJKX7r10AXSXG84Mj23uFhNzV9OSQ+SdwTOlnRGO
qO7MgSzW/rmIe9VxKIZBPhogXS9+Xv8KbukKYe1WZVbdoqZg3ywLEbajr1+SV8pF
l2fR1emIPIjKe2KZEZjcPPNesEIRWGGnsexy7+l/ELosuDMOipm81OLrOxaW9CJf
Q1DnVElA6091qIs7En+yqCR1Mj+TwGKL0QJLQ8/nQUpC+xZDBT17CkP8P3doBP3d
JnE2776z1ymf7cnNK+9sUs7Nn92Ldg9JZJxr5mUJRGUdbxn+yqyC6ahVYHhmiss4
FE4Q/1QStw+nOzt43K9677kO3mp3Of3X9htd6WV8O7NVLuE/qVVJ1QFm51lmrh1g
5P4RbEB+D254b8KEzVbvvhEtNIzDCW6RPiuEotDzve7FZW9Ye580ttx9p3GwXQF1
mh/v6Qckd+2wPMafo+GLI1x/0zljEmrOySV05TzsuM208mpxvJ5Dbe4p34UOFV+H
uRGqVUWtweNtJmBEHorK+K14PESxMlTqG7CmLAqZkTTJXu5c5PYSU4YHVqcRXKsf
R7OcPZBmo8bLcYxuPhSjPkPDIc3CN5gnVVNv4YoC3EnPrkkSwsONBSNZHdp8llCY
KdqErKXpSyQ8IXxuF8bgEM62EppOftdTu6gTz1nNC95bHEpwx4ujcrYjD4ksbMB8
2KZcPfMFYYscwAsmaWBCRlzCI01EeJg6xYPvQpKCXESH8VY0zvgHOESBcpFSdl6M
DiXtF4WK/wfFeC6N+dvruKEijh/1zujI9PmjdZq1WVWrWCZeeHxpPVOgjMO5AiSn
ha5OEmf/NRAAEB6bKEJnVFhBKT+h3cliJCyTKZ9HUhmFQKDctFXq7OWQpTCNeQKl
xUrIWvpuYALAu1Nihcdqf09lWPKjfMB5mhTjwwfNa/1mHIYfdjgRUDmdsWsTdZiV
92z8UIjhfPjNGlhEzD2del94FNlP5HFQ1czZbw8AjEC+HT+BVyDF+HRa7R9B9UUp
/Tf3yut2GWQRoIQJTxxPaVmPG1DmaWYMZe/OREQ5BrdZdSp2GO30gnjZwGu4w3AL
7XRvHnq8PsEeHQwUJEAI4EbLkWhdO8ByKQ6vSOg89KxxJem6zMyKsvbI46Lo0Pmh
AzQQnbOovjyfyZlkX00P2yVkno+jekIXewNimYabhQTZbquwuZGn/u9L29AsD4zH
7dYYy1aQpHlvW7w9BDv0qSBI3QWVMyLmkmc857goKrHDWOkVbg8Y0B1T/D6eF8a5
tCuVEcZo1vCFCRek+1vOPx0pK9MsHlgp6BaDv9Tk/nklu8Zcqr1cobYlULR6y+kQ
CQV1JCBS2qayEeg0qabEJGBzXxLtyJWo+3xqhMs8sc56F26MZWeqvWVe4WLXekAz
PJGi4y0KfVaQ/gidxULmgKgQmkDplcsnfS6iGodo9fnzNHyxayQvOm15Ye42Rswk
GfugNCPq99zJuLwUOY0ckX/YrCqx1tZCZSTJN2ti8fBT2e3cwUxdq4TEJSxLBJao
t5Emj0E1s8tqIEbZ3ODGBlBp0jVHmyXsXeWuEV2SAOQ/IdgTTgefy2n3HPxI1mCH
eunmmZRZtLrLEJvIHq1btP5RamkY/N8MCTN4RhUbIurlzrkxy2UHGJED2t+Tbl8k
y7+Qp4Ig00CTZU4VIHKlJ4Dwf1H0Qcsxn0FieOp5y4+eWQnp/w3DaI0eN6YjMxqu
wkYsHF+p8vMHskUU/KzhsAimk13wCfdlq/j5tY4kAx//UBgSO5o4ajRoVWkufd5t
NTx3+8bFayE47If4YACMsEjIOXS/ajYpnvaiOK/VBxpCkW72qJnl0uwIicxWF5Md
YhSwqMV0yZMSUzjWpC0NWDNPERC4nYAGly91LWdPyNEf/4/KdQq+9CH+HxxMACXM
8QuWXNZ7XyNE1fHSMbbzmONmGbzUArGuDJSVVPacx9DirDb207oRzlJClJq9rqqF
rxoSZOY5CgofEoHMSkNeIbxSqPOI7I+Ayw84G9Yp/4OdCt8tZcQf4P3nNgm+oS+H
XQJ0vuUfAuod3jB086l0LqDDImmPMFRwbDxhs9jYiVvsGC89u8pbwe33hCpaUrsf
RXAm5xIuuzqANLdzA2N2EikRABb0uv1C35Sym2H1WIVbLsvA1hmxTaIEaZB/fBG9
fzIUmHLb3XQ0bAai2Lr928JKJC3gZR550wpUorTlEIbpfgIdlswpBWRPuBDCB5p6
DbwG3ftLIztWqgz3MNpG3zKvOneOn+pcW3BrUz2j8PiI3vgfDFyfT98XGGUS6jT1
PINuoiiNRrT0+xa87NrdWuJ825etRnDCDVq9ob8F2fRbErkCOa69RZaNKUtlTCHp
un7G3fT1WMfJM9OqnxNKt3q4p1NNK3Un6v5GoN1tJHrOLqdBy/u29g37zRLovtP6
EAdBTcptJqJi1diL1en1BJptZA7k59DT69dnXJ56AYJBrwJqX7rz96hqCSg95a4Z
d9zEncx+jT+lrfhY6CVmHFoVkCxKmXRGFZQyhwRjT2g/+7RJFBgvSYvJkMEit5Om
sq2uYodJlohzr9EwI1HcAadx7a7pflDYXERs6iHwM/cO9KR/nLkbdrrbtfYCVQoY
F/eDk5x5bceqVYZ8h0bYa/VJKGy6lXY1RNDnnFBVPBAA48c1oZWNqbcKIWnl7eyW
ZAfkEK568IKH8SBsTfGjlwUTquT5eWSlMScrqHZbMW+sgiBQu0MVfUG0TerdLOdA
UitssxqRnguP7P5TSBoGu4or+qYR+JJxAKQpIRnmdcFqfsGMpcf40iCFZ2o3ylZy
USs2iVHKoUL5FKRZZ035eEuetZXEmGthd4hHa5bWD3l29182ywG6FFUMJuSZys4B
EtlmAGViRiiJHTKr1HNqea9I4t9AD4mkrA3MvaM+gTfIBmL5uZYaDw1WBEc4D40x
aay8qZ8MA6Bdp99iizQsaXnKm7hWU8WFOjsvctgXHAXtuo/D0TI23QEnffvYKXgO
IfzTGQsb3njAgSE2+oFbfbOBwXX+ry17SZmCFCnc8CQnE3TbHozAw4J81f2v4TGx
bKR0zWeDMTil7eJsxAf4jnRTWnN0L+rl7NH3O9CpnJgz75u9YyM3wO9lThS+W2Zt
qWj9GYKpumwuW49nAQGMvkXNXQYAHVqsKo/FA1B691TVSgVjj7f055v7ZvKiCswo
rWoxA2UQmUWQTqNETkOwk1bSNjd712Vz74kfTDC0lQlFoPVEDFi0OBMQ9mrV7aW5
jv7c3VJ0v1rvtEzLmh8xvKD2+cAxPaLGjbmTRDaBqBW2Rb11Lu69+NmJbOcQgztU
fl8wM9zfvP+IfYdvWtnJYYZyZTCWSOFM8pwzGX9NZIWPdn+WCTm0KOakGzhpNzKi
MVDzAYRr32HsMreTtVLZ/YqbHjDMVQErwd/mGESdl0f11f7KZ/BzTbiHcsTAbVsc
3f7GFZOpnzIbINONLPGNEqLDZ9x1QHmBe3l5wHqUZRGlWkp2/v1TBZTQYCkT0Jg5
bwg8BpvqFJFC7K0/KP+rT3lnPQBjsSDh0kjGtp9u6GAqy0DU6pwtgGzUnHN6R9Qo
PdGQMJWdjfbWKNADJAmroc+OIW6Ndcri9g6g4q/OF5f1WPcD9IMZKQHxgC1EpACw
PwfhuwWqHAAkYwyzyDLxqP2kmO+1/zu3wGck8jQEuIRpugOyz1bcYBS+aDPCHbSY
p+qdq9Ui3XTBTWKvClvLAQXPuHXT1xdkCo1wfx7rMu+UK3kapIsPM7KERXFNzord
4iI1FekjP93+OBIgIX4ef4e1567DOjw21dD3HMNl5SltPqJVnQGKzXOZtBG464m+
R9jg3j0XSdf2y2j8TYn9YM/XAM+ROgkypA526ITQPCFMeAshP02J6GpTfGEZ3gHL
8VFx3gpLZSI2CgJB14XFOjOOlOwhJ6VXTq7omBG+MfAUcZcknsJF2OqQF68/o/Cy
7eVthxltz3Zf8cHQgZ6uzOCelHkk9SKtAn18lpnw1Cb/TsFeFZejas7x7/WI76vM
VaJEAX5JgQ/lL63hHyGdjcwKAiISxN4rCIELnj0rO2B3HtMeGqSNVUyjMZ19f/Cj
daYjheDIWHa4j7zixTBniB64PrkAZU7/4nWohY5j8ekdBDjWhks5fB+xQWOeE6i1
Q/1t/FirVQ+WwpvipOt6AisVtKHdX8FszSqfB5NocX4XRf3IRiCT0vezhSKaOCaF
nGxZxFcNbPp8pUP7GLPZvoQHj2vpESPi50FwBcTGej7myRAon8Q0sMAuUjMcL5a6
cpt4uY4aBgSAhCKy9tHy4rsexel7nQsulAyfIas46Yv18XXYNM2lzGi9myaoKVEb
DgSu8hXzbpxhig90azsjWwyJOK6dbhUI51IL8icfOA+CwsSqvU+BI21aYTNAYFcs
DgW6GsN6XBzeTCKWkdIcZ6atD6/IwlyqEGFIGYhP3efLffIsiDLpLuTntlKo8TTr
RJaDiHKBirs1rpFuTOorOva+7IC5PEkee8CBKmNSKLaWT4D5584hGyWnLlnMxIJF
ClAa7goAwo1fLj6ByGJPFwFYz2UCDfs4H3oYrs1bzOeFZG8y9k869UX7gbj6PEIp
kz6HxdOLMBYmn+N7atLxGGisUGux8gK1QBqy/Oi6ew20ffBC3RjsJD0x8d1J9UiZ
wUmO/5m5Q4j3OrO0AjlKpGf2J6B7mBrtis2p7eoIdcXPeEHk1n0O3yMFOgxbIYzr
bwfGwI8pB4hAfUaXf74ePelM7JD7nHM2udBHIgh4w/Ta5kqVt+UdD5rPpq+FPaxc
u68MSz7FNfRPdDB8pQ4FtOceCZvI2cvjXhnIRqy6mTLwM0KymHO6QfaXLCI3uIT7
SqkQwEnvdCp4Tl0pdPrd42QTbE7W6E+ZDzPbMd52hPq340ZbomlCGXJ8pdrKK9c4
V/8nwn0BychX/riBdi7g25mOxzz24KeYIxPlyQkDksB5Vbt7yGr4/9FawjmU9kMv
HoLWGSbsu2UfcxWoe89j/hzA8ZuU3jPQCYtVZWGgHJ0cuw46XTr5dvPgd3V9l1/D
0SmbBj1IVNEEg7UN0/vyayrGOM5zqbWO2XGkGv0VMivTcqDQlcDbEEWl6dQuoEJP
fEb1wRXBP2H5xVgsCjofhQyAecAvurIeP6j2g1Eay/3Uwbj9LHo+Z+Xj0xn66lmS
YQM+72dBII3QGALZbA+127EgjGUUW3LmkKRvuQsIJFEa1Q5hmU6wBUqnjzXSmKiE
6hUmi8qX4vVNTxe2BlwMlZvgBWGCrd8UgZOBJIWiB0asOQ7x7BmfDbh+NTZHS64u
vZIfiD6r3sYAXleAu8K5J1tKki3sCP6g32X4ceV1aBO55BKAnT5mK+7VvAaArjtO
6K4CH1P526d7O+jSNx8TifXaFZZM8T7Kujjlkon3CKR8k5V6zVQXIbJmgBXA4Kdc
J4qaCMqoDsRl6MojTdIcwiM3wJo0EAMHaAkeUKlAnVe36FUMCjsNYplnUI1reGRb
8yBjNrKSHgO+IIdY1qG5L1LpHnEwH1G5GNGTvbMz+EPChDn+QgkHNWe6RHbnBWC9
Hhk2y1DAEOla63Tj6N/G1VfZNyWLEonn8n9vZ3roPnKb6wBV64GEFaO0ll/fDkUO
9iusiM1N8qij6fw0nfQgckocfBUo/AEQWYIwTPxeHJwvRgCqn0HzMMKuUyKzlN/L
i3JBRW+1iUI2SsekQ2UcotVm7X/u9rzekHQCjHMXjQaIz/UOj+pkKFPzmAge5d95
2WHs9tX8ZikngtrxM8oUOfR/AkIopd1fx4QlzGQ2JX3xIwd7NIRfZ+tgsgrgE5kd
7XOC+vLqiZGSO5f16x/otZ6Zbkv9Siv0B3ybqV6hSfmDJdTh+JfrWm6d3kXyfVxD
Y9kWe3Vf4WZ1bG6H0Wp6921d+z6SxREM4d0YvMoPAGV9XAO9Cua67pxbrjaNCUO0
9MMdBC7N+VWIn+dRW5I9Wp+LuG9wrDs+L6VRnRy5Iv7SXj3odL9W44jIHMPBM6F5
KPCj3CrkXzAHHRcJR5BWtJbdrP0pfuEgzOa1hDUkRFlNYArDcrqf8uJAYJn1A7Aj
L57nSmf4NxvxmAW77vYVPYLKc7qK1cs0bd8YLGa4EkGnIe/UEineOl1YOGgUN/qN
/m5T5JwP/EWEh+VKoSzBchpyeyZApPwvne2vmvtNfXXfFpO8Yj/pgA1nuVK3WzPC
M7t6sIoAhYPnDNUcX0w/vY2ca9w6e8YKtL8BsoVDbzuSRZbSjTH3IGOspb2zKsQK
Umnou9AmWE+5L9Y8OVWCF1nkwpHOhK+4ZMTa6TqfW1MfJ9Rpp+AlAGDKyzy3o6Pj
MZBdHI3brMMakABHhfnC+PO3kI6VeeVjn1DnhCkFNaWUUZ1+5HNwQHbZ+N1jwEAT
Nb1X3Gp277XLMigcQ0KoL58OZbnbiC6rds073RwUl/CrgjUCu13IOeUKKh3u/rrZ
zhCm9MaHvesGy46Er0bk+QHSCi4xO8KdVs3s+BdoVq4fFuJlrwx2MQsjJTtj8l4s
ourC/8A7CHC5jdetdREcxVOD5RDvWSQLgYCLEXL9AcMD4LhQglWTVRznHAQdbqC/
ZFcZnEk6qzFcvSAKC412DAsS3JuFuFAqkGjmewy9Q1K0iN3Kg3NQVaIf+xkdv1UG
C1GGfcpo2Ip+haJyotCDbKFit6x5LITl/TDTZU6lRgM2dtFdx63B5zO0iIHL3Onm
NJZey6sMG8xw+biNB/N62QPKP1X1R0GWucYkypNH+VQa5Nv07M9vE8b3a/44A7OT
Ov+Ld17xz9Z49JLMizP8efNbtdZRFzEgJMmnVdaRVDrdJlNj+JdSV5+ZRBQzrnLF
PxgrxmHc8m6mibyRwx2PGD03We5FkLUB2mTZaxi4i7SousaLqUCRyXtAfcBp05TV
XtaOIZNQYkwy501JZ+3HiJ0hbXc+0gLrHrqZcm9icWfusz/9iYFqGfR2UeZtBzIT
h+qeUdRFKwHvj+UgcZx4Uu7OMnLkMQtl6GlZTM8Zqw6PeMsvD2zmBHO5taK8+kwG
6YhLXqyJ/xuFQTckKnwfeCTonyFtUwAxe40EHgVP3lxJMGCYvz6Mnih2gsr34wbm
Ef3L8HAohmEW+URoNLYvy6FvfJX7awaZnco2Wa7q6Ww6AK5DHkx/1V8wuIx0PMU/
YSnmnROLFJLSKshld5XRMvRPQypUyfnKu5iiM0+TJ9TzuH47RBSvb7dIoZoKknK9
tBZ3ufCt6kbSyP+uvVO2L6n7zkkJB46IdgGyF5mcPdYTQUQ8+vyjrtHoMvCqbk5q
fE2jnzvVYCxpPas2os1SpBlFDDr/Q/gveGJ+W+/W7YaLJRWmI6mx/Gx/GO6aXY8y
zOOXl2zHO3GNsyjIXCw1q34bAQjdq1cSL/DVqghayfFYoTVKLJi9/weKQGmDYZv6
j7ifiI/kYtdT8eCs4PK62BRXBaNjgVXaDd6+XDzc97/HcFsrurgfZXZzDlN3Oec/
yTD76FPnuMocn3ji3MgArie6ZjNQAIn5VDpI8cPr/dGsyZ762kK7i+jslLRZRGRO
5wJ35G3HBhQFPcAmSF8s0ysRmF9yI/9JxhAwJJaKSgsdQQOjblInEAGKbj69El4J
a12+BWk0NxU+0mwcVxCGmXvnJd6UG7AvGI2lBVFxjlhFf8aEWtiuvzPSoQUC9RJv
hRs8TnUBGk1D3/bKhIA6eU6IY/DcCDIWRu1um2TUCcZZ2mgKIf7fqPq4k32p3Gc+
tNOXVXS+yGHuS42l3eGEY8UHZsOv8cY76QpAvHccDn6pJHmsyi43Xyn+0JzMCEXi
5A7fHEx+d2EPP1TCXr/Ssj6QNU0Vt3KBVqrtrMhCOt+OHt6ZTYEpnoiljz22iIut
W3tOv9kPRkqZwRty9sRwILzdRyUOC3qAW+1Ne6FbHHOOiBh5KBGJEXApPdaXteGA
Aleg4T/UAqCeJimtuYNRj95XpQ29cefe0iQ+ptky7W2zWeeNw7DGRpKB3Xe9vTrU
xH/8Pcw9HRgxk/VhMoMsxuNi9CubTpqZx4vRDLcEKx1Fz6gI/6Ydh9jaVMfwbXch
5oDC1oREE0Ss0r5q0A3CvXwAWsMIp+4Eppq0WpjNfLanPMrc/1KZD1CoLZlFWUAE
uKitjdYrad30wPpOJktmBdYoSPB6zh+oMnGy34W595OEqHvqAseupxJFeh1F0FAI
NE+VqruxQjUiQK4rqpvqEMvjzCotg+BLfHi7phs3IzlnRXILAMoVuiFGmz08w9Fx
hrvr0Kmp6R5zqDzIhAX+d2xNT53XqzV10WpUN+Ua1N+emucUwocwYVyZg1riGBAK
1wasrptjo/BAp6CpeDsZ+JuhXLn4VEZ/D0o5pS+LKdvjSc11ZA6WkUlyQCq3mh3T
ZHj3hZbp64ympJNg1zvk5O6VgtbtwKAwYfd8unZXDSgCf9bmKdEEYYNHP48Ox+6R
DRnJIz4XBDvY2jeGplo8+R0d3QTpP7dna0VjZyzH033A+trTdq3pA05XbxxuZgEY
dngcYbhOYAylK5nXi/pkoSBncK76B6ET24O9358rCB5UNsNf76eqKfmesub0iY95
fOwo6vRIFRj2BODPZab/i+UzbIaMqeJWt/SySemqRNgYlbEyIS6J6z2yDYGxpQOP
hOxKS0ZbmXtKOAxEZ6mS9guptFUYb5G4muI3gOAu6qXGJyhRTf0sFjVpZ7XFGmjP
8SoAyoC1JtUwjDfIN7xa/UprRQYZXEZJAREy2K4sJfqFojC1xyCZE/7DYb3h1mu7
9m5XIPSgDRYCbrZrUTs9/GhrtYd4NxJa8/Pe6EPpXmUmRkIOLcXO98/KjWsAa0NS
moXjp6tPEOqX6BJ+RETwlwXoKgIKSl6MCTehPTnC2LWeAOmYtd7PafE15OccF8Nl
wrG1mBVOsEudMIJmevhFjw6rWu1LDtKTvS2EfGUs0r3r+LiAytkdn9KnS91w7rIZ
mfIVnuzgX6z1N3KQQdhFweY6pgh+PWMwFzWwiOzXXuOgHqv7BLd/Vja5LO9+SD8i
B1nCx3+IvZ5iT7dNnm3QNeoiV7tV6AUmGjO/MbDzVU2/GgBMFrJzpVdf6aKYXHtZ
fWqByUKA3XdFN65stA/DjBt9s8Guib28W6rpSw+3E6sgiIfno3GS5ziVeOas+/c0
hCiSIsOH36616U+sLYlYVonZxBs58LpmisjXa0RpfE8B12JQRO87fQOdkvciAtDb
Nnc0Wvdbn3CJ7w7ocGmQC8Imvl4ZJd8/ipJl0r0sBn/Mq357NSxPeuNieNcndZ4L
B5GFJ4BlywTspi47jr5PMsg4zk1VOluDv3ZOtDKZZnp34WqGat9JNPPAU2XTI2vp
43kyVRGtGWr7g8Nbj5VTblVEWZKKGuOAljz1r9CZDpJ+XY1sKwtAsZHmY2OECysl
VqNn0hA4HWGFNqSLJD9Mq/ffLp5eggaLq/kQXKDz8K4NK1yfEh5gz0A3F57ySqej
gjR4/nGYddVXSO7hIj2oK4ZyvNAMeM4A9yLfKnCJJs+2kbRX2D7UoRa2aPw59iIx
K7vsA5kmbQ7YmM4vd8ixvGirnuC/1PF8taAWzuwDn5k/4Rj7nPbMOug3zovIvVo/
dPDexHdsThyl3IUU3GIYcgqsSYo2XCZ/bPEHOsp3saovjW/F+lP0Its6LXymuo3l
m38HBH+u6ev9LXmpjVQGzF73HVbBWbAfhzSZ8q3K3WtRD/2tVjjOVsxUhRVRu13e
z4ZSVlrz3quTDpkcxVrvoLFnDvi1EvPDFgm5BkAkKcJ82ACVLh/yeJXpSO2dMbQD
1X4mooazZq6ScFNvCvdJu9w8ZMRw1akML+52uNFnAPsuNAGMM+NseMPqMsI7t8dV
DOIskF1iGQGhMwsr+6C3FlwJE6d+iZpsgvZt3XfGOqAFs54v5SjxaGUXk5LLJ8Zv
4ylZg07yl1Gkj+dZAr1rHpLiLj/xpssPUeCUwmp/GESk+arJN/vg7B4plyHjJIeM
BI9rMJnbY4v8IvEBDiZRlp4ccRBRPXjKac6PIyA5nZzWcUtN18aT/4Z2kZkbvMA/
zUcl8PexAdO3ITiPPQ5eaSIlJ+5xTemHTlmbA8agUTbMzf8vJLm35qvp94NEsXln
OkUBn0Z49nhFHuY8FF5KB4HLcG+aWPLQ1J6wz4EoRPpTN6A4AoIibsxYiFJfl4xa
MyfXvA8JSS8gQu0O/lEWB7ypC+lNO4ZxQAl7sOt/kxVLqsqJgpclvGmxNBNQkpoq
FJ2HjFUzafk5VJM/ZnypdkIfYPFyleV2xnCzAipRRqp9Rp1wIHFWJjnQARplw/tq
Bcn6BzCG+3zRu0+bGbLmqW08i/k0sgjn5yC4W1xaBgEXYnsDt12bNwZgIvrd8fUX
p8G6cPFTcJwFiiJCR3Jz+vxUpuqfXDsSv+S1HAt+vWfh7VmZWOMNHgtvI9fbd9VY
2KNMZUSFCz7kUmF/VKNCTD8Z44l5ii2fC4y+XN55xAJTdVwyIi8jdoIgrzC7jcek
GqC+XAwLyptbI1WArXgMvfFj9lHrIffv53j34aM7QzxjOh1+1k/+y6u6OUzzrhMx
5AFALyE6Qxaxu2n4ikEflCkB00jHnz+J2NJtMef1Fe2KLz3m0Trj4matpunsOCHz
DPLbfUqeLAwwZSByNdRVv79vgeKKJ1wDnI+eSH4CLGatGbgNnIvHRRTiCxFo4sPy
FRvu6g26S10D4lwRtGyIkwWf1Fv9Bj3u2pZ/YRBwETFBz6hTJprd8+FVSzn8Dawl
2tqq2qNqgqrnMGvVAQKW3fJwVGky7uaWvkkUeZFsCh0hyefiZRRNst1fMNxexCDU
pe4Ycdk01gWUGPDpi3RMCgobXyc8X/K1oV3+F0w3Y+MYuHz829LlLo7LWAPB8nK3
DdGrUcvRFHsFNjjl8USYHHNphBIkW8K/M1n6ptUEat9Xx43pMMh1mCMcBsRQyzzU
exsAfBmakZJ8OfbgZUEhu604PPwRKX0LtjOyvtnVxCoRw0z9AqP9i1e+1d951lyF
pbP80QJN2ytt0U/SKIoL+6FBJrO4rDkugSVONcxBTbmFVWD+Z5ikFRTZjdccfts0
APmWG0IkbmSdgNVfMgScxFuOxToVJLnK9CY+6AIz6sKfyYCANsZXf9xqEkQ0pLtU
vv/8kW3nx4mxE2OBkRLb7rSU38hCo0NxxZjZdVfSVgA4vQd5r7zhRkVliAV8vKRl
FAKdKXGAwHYYL+RnuRwfWws8JDnnJuwFzOMQL14xsS3AXeDdCQlEtI52EwxYL4Qw
3TGQDknpMpW2BHO4UTRwqJGnKposfmmq+Ne5L51ElKZvS5gpLfD89NbazjbA6pBK
lKaDBAtJk9S/Gw04vFknOpCFiN3/Qg0kGfkonodWhiyWg+iQiF6W0nyfLp4FEwUD
/XbzoPLIG3MhhiVfqieaT38tckFJKmA17p7YCaumgBgXYsVp9JlgBpMnLDjU4ca4
kd/01EgV2b41jROld9xzMughBEVQfmz8LI+pfxBpCjCPgi8rDWbhcdB/RQhOMkuB
9jjYV7fUsOmX/tOVH/tVn5ObEkN76fUgFt3Kx6sh34UBitwYDd1scrfgdS5GPutw
HjOYFqQG1nEHuhbwKgNKVfBUYzfce7rGL4dneb8oretOkUz//f7cfPdUtEbQKNgk
CQBhOySDoczntKVmgmGIBxcB9US+BOE5O3kHXDJl5j3YUIzsQs9ttxnY91Hs42Qo
j0EDmvjhgM201GMiYqwKVVhvxik/0dotZHVQ2BmjVQb1Ht1hnjqhdzGx8JcLTAtw
vT53sP1XMhangn0KyQYFXIlu7MEiHodh9PIhNFXXaNpRcMR5kdIi6CWHKsiPnLJE
5+FhOKwwDeRDpz0r8vo6wvNEI0ROCjvKnl4JabElI/lvFNhcTK3cu0isc0twnapU
SisHU34v8g3l4DS52y/eXRaqGX9FMfIG3pGdoRrmYd7qvl4iVMOwZrPM3E9V7VgG
dggjpdwEMZVm6QXDQ1KBwncDIQIouZIrsNXXeeWITZquPcqBP016dr3Ktis2OAal
DCzH0WsJ4Gebjwu3HSIk41A9SZjzarXzLoUZ2abYDNrpJR7VNd4UG42D5V1Vc4+r
SvF5kegPI9tSG5gH7WAmNSMSOqlIGObob0uqAOmX9QFA9lKylNE/bfu3nKHstClm
QU9ew6mYAN/55AAysx2LCArl/AEBZWlv3uEMHLIxST5FYMN5B1MvDD/bjyLS3HFd
IC7MZjb7eF0cwEP3m2EBsXunTKpFbMLV5M6Y/Xh65006oAFbrRtVjCWGzAoAMQB4
gGsHOci8a+VZA1DDs9tD3eHkB6VJP08Wzlpn3EilQRYEhMQXl7ssF3h8CmZV+P11
/BpJUymiMpcKUcLrbgyCh6R5XLwZV6g+vo6Qn11WjA5QN4u6h2SiuX5r0U6FMMHJ
Wbne3QHh/gX2+fbU7q8TL11f9qVPb99j94O2ret3BrxcJeiJ27mKxzDv42NrqvqB
iM5VwrF8QzEIMvvD8qXmHnSumsNok7+VAxAINYiHzvjA6uTH7YrQM4+olKtn27Dr
gR5wJLikvUzXhRjCDuFJqgKaWOr/0doyuhfdIX8/HO4sPjD9FiyIMAviJCdLF2C+
tvmkgsmPuqM6dnSGuzOZLI6c2I+PioWYnM3edZDz69g+l0tNx411eYMdZBKKD6am
7czrrnnmBXnUYZA0XkNNSNUIP+U7Aca29BF1m6RlSGbodBTZxSEIIyFHXQc2MXUn
SlzIa/BqfSEHI5nH50Fe+NJAH4QKMKfsEyjfPgRl9PJmix47yFE50bUxixCRlRs2
87BSNTGafUG5cP2qRosQv7PAXrZaiUj8usKEQz8uHEp2yoWTet0X4D2OLx/x1696
mPBMSB7HtuDd/bnwcMtnQGG3sfTTW+ABAIuZwduqkQDlNHibJ1UrDmL9mrH4CkUy
nOwTZJXcfFp5SUcUKWYCtRB25csIIsBcgnOw9KOonBkfFbne2DElTArFEz9G2o5H
4ls4qUkj+xFIrVX4e/ZD92S/7yMQ36qo78X5V0pT2UB6xDgfg+h7JIA3Zfr5BNSE
guaQy8pSO+DqOvyC9/X23UdtFHS8CPTPkNlkvTJ/FARrQAvoGmeW0hW2yKE+jer7
/8X+n5N9SsbATVhpfX0tfslXsjEXb8Lvmc8hOnFLnu12aR08VR0YSzxk7akyzOLo
8xI6WgmaywpLfc1A9iDwpZWK5NuvlwHhnGEcwkVu/ikzejkdkOGd6VxDzFhfT0/g
SXHcvHZs3Hm0XxFlKTt05Ub5CrSl6DWMaRMOxRJ6ujFQ607sgOjYHOzsB497wInF
mX4zicGadVKS6UoANnPdhoQFhC14j1P9Y71UGeVADSZFgh4bv0yQGDTNbN63PGbg
pya0fzq2FhYMVI/cbWDpbQfhYIE/y2N5ujnN9ToBFU6CoDsHa/FyhZaUmxCn34RV
ijQ+VcGdQT6YR14BmQrWmcYYOqd7gb/BEspc8VPhCfn5Rug9qek2xVL3N9Gb5cj3
vaaDGA5/YEa7p7g5Naa1g1+G/tRxN/8KKC2CfLS5ugZLfCPUVbkYzUKkvWs5DJJL
af6mrZRj4+WBZMM5hlm2ETYRdATFZYsoSxKha8Jy8KVb3OXtDxrrOT+Ss92oP2c2
Vl8W3MCqcJVhwljscJp0NgOC75ohMnVdfujIH2WozOYkbzAwhCxGjaHP26NiksGu
d/PMKOIVkgWO4SEDGMsa9UFAYktRHWQZBppC76xGGPKWEu6M7phlxRodzNu4IJEP
ru+YC6Ck0jH/kuG0ifOA/T0FCjjamhxTPu7+h1j863QVZ2CAa8ig9di2lQuPxgcS
FJCwAXGiqlOQHLiwaUxNapq+fXqMBZiGEvMGwAajNK4ykYWhs955dXUicHEMZenE
3qecdzhESv26S07nbPaQ0YtDQ+8v8uXSYU6MDc/GSvah5rfGaphjX3E30fRmppji
9P7naj4JuFo5ZC4LXkGx78zBcfTjHs2e9KH3Jl7xrF/g7WHHnr8BneciGTJx3xB6
zekubFVuR+olaSKU/IEcIachWfLdEchTGCs0Rz1GX2flLK/p9jroqWHUnM47/VJ9
7UsamA7JPxMlJXFB6qIA2W9zFx5vPA0vnPcsVPc0DI92vpZxczvQS38BY7QB8TRf
3QHh9Dk7In5kYtceC1LfMi4/UyNM5L3uM7Pyr1h5NfEn3htwaa/qdEAOjLGASHsu
dCNOAREg/L3v784sDqicFQCWxsjmJhRbyochu8XKwRFzaxlV81QUeOg91F/UkjWA
aAbA9j54CeiM6cvM/O0KQpAI/j0iqQ2VKtjaGWktGUb8QbKjezsslyVdb76cYkWf
FLqZFOp4eI5p1+YthKRBk9I5wOGLZvxzBq/m9O00i9lXuBTbcHm4ZnUg+ZZdeRZr
+D9zdkTjZpM/FnVOj5AifU/AO4oty5Lui95Jjj/dJ/ln9Nf7PLDhPJwZQjrpXLR+
gcSuM95IqoSULji5HlnS6vDCQP9gAf3qsf+sYFr/58bcK3pS7Vv+smO4k1PtfXFi
94twCr71w+qX0tCAO7cDNNNWXqmljXJoddJ48oFGtV3xjY0GhM76cZ04cDPyiZEA
KLPdQDb2cmeILFVvUSs9ZLqAxH8Nx5pDISH9REIAigOcEyeZjTzj+mmnBSURhPGl
INEZTiVBjstROUqg9HtZlpB3reQ0KuGYacHm0idsAnRx14J5s2vga56i+Kl+q8+L
wrDUF4iZL6RZU5I843GD8BvA4teZ61K+hLO6slK9D4XICDP7ERy8vsvRbb2YH7RL
EGZAxwydxKi4qh2A5iHEwN88NbAvSglkc4DiFYRqmO9UpHR+y0MFwkzDwcR5Fgaz
f16VAPbyUt7IMusq6YFi6TYHubhO9L9Mn+YyvwYsa88GQo/3SDhBr45WSLr4ciyN
2S9vQiMkjQBpWUuaHxDG+OzRK0Lrk2TPlaomeah+pd1iyG2sgZSKwaAY6RDuUCo+
/9drNX8CfsONERGtX8DrqEERiU7oGMnucUnLwdYnisrcIiSDOuucynid9CXDOmuS
U+yLrgRvcXb0y/NuqFnJE9LP6KP80hmiIh6VNnDAs4QoyNjxwAretRqDa/DohZdx
tZbjNwklYopHMHmleQ9LnhnaYlWNDo95Ucr4GN2kepuxAiGVJQmdK+yEXJ5HJBid
JZ3N3AgCYuAziqSxxTcj1PlTT1c3DEdzEUjMjAVC4eaSfTpD078ztTvc8LHwY/IM
ToIN/bBzN/7gMjlRQd3aOiuQvVK3ABhrWRvCUpJaJ8mJwcMl3S+xd1w3nF+sei0c
p6ZlCB5MQJu21o+cpM8vNOsvfxrKmvd6yDX2O7SIte+FUaYHpVH8l2uBGoFCKJz4
WZcT5IDKtbaj2bM6+egr86UJ3YXtDRXeZdzbog0kFqu1T66JcTNC6YUd7if8dmWq
mcRFDLsyc5JgiuDNJjWgpUehTBstqG2XDAuui9UShLt2lbwo7r6snMWoNjQYTEN7
qnuoHTYV+ERjFoprcwDhb1XKhk3UMiBbM0S/J8d5ZkBuFPj46EvABodEX8rEdixv
UsXC9IjHajsU24T1k16+rRIPItfyspk8Vk3ffGksmVt99tTH7EEh76VowafojmAP
ErIXOHX4pRaEnAREsyPbnhXQH8hG2hdUXjY1UmhTyBm3K5I9emOgm4UazVMH4oqj
cSUgm4p5hjtqRjHexCkFyE1hk5AWSs6h20ecogN+glXooIGlgh7yIVuk0b40scuN
/7tCYx/d01LOxCeuVM4ZptoNrqGAYYzUPO85637RPTsmu2xUsyK5NOEUre+hoTkJ
pfVUvWLl8FdBvorZMmSEsfht21ArDZL59gmIFSLhHVhnBVd2nrbBhFSqS12Teyrr
lyFtHN4obLHvZEzgHC39uCIEYfSH7AUiZ70ZrTn+G/3CScuuYMGTayF6hipF+uyd
K1XnZj71/uTBWwzM4WQzi8Yq3Z1dsKfYAIHoQU/30WRyhtAoaSHR3uSO4LMMiaWp
OPNDA+U9hj7AuaK4FnaiXMjXQAE0T0OVtn/uGnrbL8wrsQ7qS/ynhwVoEd4y5h0w
rY2lZSbtHG2jWZfd92FTpt4rw8FOPPczkG7L9HW8z3hEepaTm9QM/4CbbFBfEWoR
fwo/G5kNEKyk8w/lH4J6cX+e7MT18auqMbF76VgES+YU+eczbJpL6j7rFgpATOzv
H5bIEtsBpBfoaGkx5YTT4ZJzuWYZxaOqF1gxWMHg41RjK8lO/TX+3yYPktJ9Fzia
qCkjmBXIcBqYH6ICUBhfbr+By8LDp4zmPNo3ONRLppGE/6mBLzcUEndtuluqb8Ib
Ta7LCPnYb4dZx/k4tfpXEoanxHZImeTTvkCGnVO8Cr9CtHanCL1COes+smHiD9aZ
kAKUF05ptie3XGlO2NxTe19+JeZUN0FS4RmPg18yl1zmVvlWFyOPKBJ7UNKS/K+u
iI33g9vAwrjtdO5EULWTIvaJRmWVCwaDzfyVFFCBFezAklUjkmR0YZ7jIbNsVaBJ
fU0lO00DRJWZIVRGt1Cf+C7xG7sV65uPXuyycPFtdZEgy3lEr/mBtViWmYzB1gsY
KvkzHF9Ow5Ekk5YzT7mdiJYCfhhtXrbnJ+RI+aM6yyJ0ROpMSt4FjS9HPtbHTTwH
dZFixQX4dJcsQxZysk2TOTrjFmc/JMttdwQMWKBAZ747pR7fRZ1Ab0fA6hk7l4bq
+aUvmABevDAiByPL8eJzV9llj1gEZys+29GmwwyKx9f62OY28FDXYzC7v4qgPJfM
6mRRNgKD66X8BjQG0N1KReog72QI8fLAgzgXCaDIaTGueK7M+cWRIiHGsLrLjOBs
1WxnX1oUPkFOtUFDl2+LenhS8zCUnWGzBPNZmcNUaEI7RwpM2A/O8+LzZZRfXGS/
YWJArEnuElvDXL6kZJPQaFrFaghRwwDucs8uAib1/It3cYvgLrbzJvAYjtRbrOPU
SrDCFS0QLScC91umjqzVydDGTpJl3o70TNjV0zNsPst1PtnHCxDm+P2PR1//DjRH
K5gPdQJ2YsJBTYt/BXuomq29uCTnU1sbzbcAbD4tieBtby0kzlVYNW2mf5rqV2GC
wWzLFA7f/JHlXrdh28Kc9yCK2bjmo1B13lR9IFj1dnXnKwPRMxyEFVTcoTjOSsN7
QImmzFioLlH8oKstKENFmaJl4gNQhyARkTFDwbhZ9EV0QtlXF68h/pORnwuOOKrR
FipCMXaISt6YoxxIVcfMICGOUZXmgNAQpnpFQkpZ4CyZaKL5+6tng4i2fzROB5e5
5B7LvnqsvLwPVgsxD4poNIJvGyOURFXd1ommiVDldICSMy/z48NY1cA6sa0YpURt
yTsEJbKwdKqMxcs8V1L40Sva2jrJX53ZoLbB54VHSJ+h3up1wT1g9rLtLoFxoDHk
6X8g7khvZ2t6JLfYlo2TysaA37bnB/79Nf6DNDKh8dmoOXVpIH/qvcgbPuXjfnuI
DgfY1WpVyo1kUZ8CHVeEWOEJB5JjrETAM4oPkuA8vj7AeuhOhg8EdqwyLt8C52zo
LHOzecS7chjrlsKoKKGmET4NzJtKFu9Dbl4ZnWc/+ipgxe6D0i8ewxL+MqzoosGl
P7rvCrZEJgja8XnjZupZGnkcoLwUBunA5bWFsgzeigd4DaJpWl2TQl5pVTe9FTA2
Z0d8Tuvpe7f93BKLJQY0qfhuo2wfNI8EjZXXpAxr3E0UpXCrPilyxNX3AlkQ1snv
o4+zDcnIYPKRfuygvCDlTpfqjwc5vjL3U5qNV5f8kJiRvO6i/JX9w9LXA3KLca6Q
bsHVMTbhaWWr+Abw62GBgO/tKR4fBdvJhzNuUv+N82Vwiyu4LW124rgrMtuX7959
jWXOlozxmviuWXeg6wiaBfwGmW0zLhFp5Hqy1T/qBR2MMmOsYc/Qt1C7azMXO4rD
Ngl1hhQr11NAPGAJG1m9ApaGr+x/OIQA2ENadxX/uxXvC86En8+naVmmY9iCVZbB
yI6WWiQ39WXKdFKxs41bsAKevJJaV4ANYT+EV6K/XjpduKBArvblsmiRmLEXeMHh
I7zYTPVPmDWQwTFtLTtTTWYl1XlroncjSPD+9SAZRIgaHdbsA8uzWXR1mRcoIqvC
8ao1f0ABooWoWemIUBHjvVozb7ROIPQkpVAu7Xj6SrssvpVUIGpSxtpmG0fsJgqp
A4yUDs/z5WUIgRWdGURfprFuYcP/BBuHmuQ5Ad8fxOUxGHxL4UtoZBalHl14h8Eq
EV/q1MhMEADvYu1uQMkij7hq0t0QY08e0J/+dt7LhvrJpzOC1wvlOPvRiAD12zNR
cwna33ZjE65sMLolilAEisUwEQvlPjKBUhrBqoM+y4JTFQ2KydiIDulLYFplgy+5
3YH27y72buKpbMFEblPQYY5/Oyf+C3HDSgQEzWFSdNiLkJxh5FEAU0OV4Z4q79wV
jBbBL2iI02gK+65g2CTbucNYJ/kf+Qq4Ccxu3gg1xa095YaZbuS9DdmVL3FpIFaX
eVUMKce6EjzbzKWsD3CDb+EwWD2oCtE0OBjo0t2PDT+aZbrJNN0Nw2OaeB5PBrYg
a9OkGJ9hHJhVyAE/w2J/SCbQ/kHoYhZRtcFwH0vgjBdVfAwy3X5xk3J1TtEP0qvE
RYcW2WL1rRC8gsqVyyLaHJ/ZdO8WfNh/eMYO5Yg2l5bTkxgGtmbWBYuIMcCw22Sa
AHiBp3hkQ6BvCpVQMODselk2UzKjnhEIuA8o2ApyvgEN5H1DIEBWuRF2CqYgBlB/
nVyuEf3j+kse6rFiQD6H0rjU5yHubyouScrKAiFp1v0pbH/YQ+Aj5V1k5tispiko
KoouGILvkvW/4ajLukQ5wCnjTnNZqIqRC4iMNW/aL7gNNWMqrHZB081Nf5T1umWE
RJVrs9Gg0c+Qv6iJBYJtTGevMawcYDDiObN8yDxDtdQSxUl6ABmVqE3lVxReR8bG
d9mpfowM01qZKHP7o7c/pKokTCoeCgeVXLWUmaOkemiKHpxbk/oQkf+QDpcVj5+R
YbGi09MY9gmdE0USqTPrVc1Shon4HvwRTwRq9KuGjMMq8I2zG4gxqjiLIaOOwwzY
JsZXlpNmaRmklLVZpU0tRe5gB4n4EpFNj8EcOiJ96TNZ12lLZTJHlRigJuPrUBgp
PHzzHxQos+9Pw/rY3vgLBawzNQE3oMPS64paD6+p+EdRiJCNZ0Mt3V08Dm2Oki5p
RUwYgv1Ghs9hKAD6wEX+VOUzL+iOVCPSp/l6eqhMWI7UT6aeM7tToDS0ci9mJkcs
sB9iZXIBqn48NVXZbQnd1tEv3jXPTXN0dwi1c8bOM3yKkYfXQ+QNWJoXUTCE701D
XcM0zBCyiNwe43Kv/rR5ZU0X7rRYOjS4j4sWPRoYxMJ3eDAp+oytHGu8Zm156x2O
HvX8vBI7WOb0k/x4dSDyjkHGoRDdrTRuRE+/k+CXY+laIxszWkj/qbeSF9LzQD3V
dB6903eo9pImArXDny5LCffzwE6w9mBV2GL8TYjXBObrvrDi/5MAdPaaiidJAJSr
NGOCP7SDdaFkzpXtcJWwKrzRHjlXdvqrk0p+wSL6lmQg9bE+nEjYGG3YtUpJ7gQ/
O2Q4mt4K45Hqm0NzcA0/dUQxm8qPo5jmuG5lL8Bym7xQ/YNVrNGYHftk6el8ZvoI
f/zKS9fGOgplabvM1CmYPEecGz5xpqCaCCy6mtUAWumpoNBXMk9JNMzNvDL0hXTo
QY1nG8j+pbEGI3SwTgAr9OOw7L6s6y1VeTBB4VUZKogKgYD6DiIHMF0lCre5Q8Wl
egFxyNWN/fK08+M5L15qXfjTLy2nqo7bxl8YjSYKk3Ysruk1ervOtDf+LAr3dNsr
kGl5YR+6p+YE2htOkcU1Krl0jwx2xX8E79kTRMdF63qZBzll56m2DloSXVfwgnF/
7Q8kh/Vi+CpDOkQICp26d8RDUzQLjbs+HKo7Ws0+kKu7ZKoqfyVX47t1YloJIm56
sZvNXVcdagxioPQSKjXcpziqbZKGmytaNR4PUBlmJyo91rukJxmtB+yEnsycw3cH
seFN8LzmgOHE8FZRRxD4UlFX2wJQxc8PddJRzOJVjw3o4S8IxjYf5CkXnqGF4/Tw
LTUaX+lJXSr/taSXAPxQUtzwvHVWnY+3KE9epomPLQPR0b19M6QRRMFbu2oAp6E4
RKDrZ1FWJqMNreDOaTbvCcmt3RVhXcZuL0Zz9L/qVTJNWMgxCHnGtWBg61F/+5El
u3b4zRT65/9D8I2vK/0xwwC6xUP3mZudjai3laNvyEyYekjGKil+gTdTJhdtg27A
zabVSUnMCvn46yjZLMqtRBg+xhDmo8ri9AdjNbFG4JI4dXvd2mJkMcLkHWoCyIiN
20r5ndSVF70I9UbE7ImhM8Bp1k6iWYh2OMWqRLYaqriHdMwyrJBkFWJTz7GNmh/a
FWYig65LMR0YrCr2h1wnCSwZEOiB59ggD7tpxNbKwwTWmztWCsZc2FbtG+G/5+uU
qQehCyP3fHy7BhgSNDpZ1aeGRlV6PU392KAHmBRzAcXOB8CURrchtUEXtf4VTRGj
1NrLu1ZhT+jCpLvMMQ3dWaFoZoA18Y/X1M+PpTKCfZXFz/TSAMjegx6TTGSzEc4h
NsZdpGU62DRI+4oKL/mv3rNtPbyQq/72ja7BROsJPgOObGDlUbT1cbRqOcAUkqjS
zdF+d4Ucgc+dr9hJLxCR9lXRiySL6IuIqyjE/+dFRBKQ37SYDHYBrsyqO8nwebhS
D7LNGxeHtjFC5kV/qR2pA5yl7WZsbqBL814phXcOQTpXaYLBblNwGsJNHAXdvsQP
N0wXUeJfKtwS0mWWI43321wxRoaB7L18x7ZhQQpBkceLyLLVjR2PFO7RcVlq7wJo
FnZOC1MIPNlc+g5wTU68Z9d825HFORuwye4CrEejKPNqrnJUw5iMKLf7pOclG738
yiKNfqXw8DC8OY1ssfpcXemKwhBXQY3RkgFykqdaQ4zzl5DrCmo1flbqZ+3VMHKl
Zd5Y/R9SHcsAzQvsThDikKXZbAnJ6h4hwDWgsm0v1pOmgAzjmUY4imLjO4Sr7dBw
kzTNC68dHAmeGe19/z8KmArFAxC/cgS4IPpCnKtHU0KTGfvB5PdIc2xRpoJytx3i
RFWAoP+eKxuw8W0kf5J/4c5phe+eW5FKBmF4hmTuEbS+BiCj0l5h4MH9rDPnI6JN
UH9LAgrr7WN2cOTJQc1aa3WpdbQb5v3Oi3tO2nluUSt/M9EccGYaSjJ6v2h5yY1I
Uelnt5mWE9Y/iNlQbcDZQCmUb1U8WZTwD1McczkK2PGYORvjln/bSpOA5ZkBk25B
BC+lIAfNdgAfZe4UlIS2B2ebpckgsFmCJ2aJc6yul+ci3Ogl8NaJDt0VsUZrjIS9
D2I+yCB+nAYIPtTxhW5guZkIj9b/Jz4b6bo5z9VzAQp2L7C1FD9KnStLl2XQBsV3
gsq5zJyaQLXX/XP5ciQ3JWqTMAR5mkK7QwuvPizw3Ek6bPF0IHblU3Zv9m5V2Sbx
AJ6snSuWTH8szn4Lo8dcIoxbXvMRZWCeWeQMUOhIY8NoIiszZMk5M+mW9vSyatVN
hsXPt4t4YvsYkoL+OvQfw8cYvV0h/fFAH4B+plvHVk14hZ6B963vI+9+6OBbPNi+
y6kOm8E/VvhZYfQGjPCPbTp1OfVJLlf5qFZIRYYKPEtjz2WFjRotd0EqZP8NumLT
SNFA9fyenJUcn1iif1OYqWQWNlmSNRRzYsHlDx+tGj69/PvcYP2oS6PNcoyxe96Y
XiXGfv4efvWs7DPxL/uM4MlLsYaJplFfDghDDwKS1hXratKnPIr0puWTzQdhT6ah
Jh1ABoIJzBl1Wy7CwpB2pamPj1AsAqaFD/q+oO/n+0euCrT0Y+SzHISeX68wR/no
2o+IVNNLKTszAa2jBjC/+KE+4n/INPkBQSwR52IXlFNckHrFZT1fGjWhDoONDrfz
9mLtEbL7IsgS7ye9rL8TClEQtWYRLxPgkl0tvl7hw6+Pqev2ouxxutQF4ZuFyjsE
+Agn7AILZCPD89R8J+QfjXlmT/NahKGKvefboGo1cuTXWGHXYODCVv+qcsTx0fi0
P5m+UKWa4cYTQ8NEAI/JqK54VCPWpdQ4BPgWki/U2DRRQtVuEn6n4/PZRjlkuaF3
6DONU3HhkXRhQBfK2Csmzmqoyvf95LiXpHOeea7pXTIOgGvFfXkDCKtv4rVPE0Y2
LhBKW+1LvytsqE0qWGe2fXKsWF+tAfh0eFiC3DBviOwurp9546D+MB7R2vohUpYP
t2nNkHx/6+Of1aHO/bXk7zrtaNhwGaXtUvVje5EEap2OlPsGvTRNN2n5stFjxLO5
Ja+/BwUVRkoorPuzmqSigneyDLYX9Y/Ten/0PGoFrzFd4biHz24pSs9fmE3JGyAR
/dhw8xZ2ZWFHpcRkQn7rCHgi50b7KYz3Zf3Uyryt1eh7Gi6F7pFC6rJFtoaX9eGR
Z7JYEykYsK8G31il3XFgSBbS1JH4nqQn41mEC4OOYiosLoa8lZUS2fVk4f8cX12s
sIXMZzSvNJYnzQb0LMAG0ntMGtvkNl21LixXnHCq6XXiBEFizmp4lD+blMB8dv3t
iQLGpiq87EF2FDOOfh1m0mRi33tMVI3wXEOHksSPNJh2Eq2scj5MIQ0X4/hSQaF+
huzsD9rY58Rx1KNwXcRKIui/hakdqy6+ch1tF3FK/+SMnygv2TlgFcwUaKgcKNiQ
Zq9HQYrqlj4RG/1LRYVfHPMH5IvgotIAEynAdjuTGpOf6Kg45608qJqhbmg5pFyg
Kv43PRCbGkWeJQ2GutQTGWuMhj9e8w7J0LhVQv9wsAAxChuvfta9riU2FL0nXeoV
xacT7EUBL/oaXs3XJIvnkB9famqhC5H8aKDNlerzgoDn98r7vAWkPoBn2/SoChXS
u1MG/+01y/JDvZCa0ikXR3UJUnLXI0my/cZf7s4p6Vm2f4AN9Wc1HDFJnuqXM+gJ
d0eFQDqFDb/YuZMkw8V0ZhG6Yt7lL8VOWnVhLZSnjD8sWAW0mPqcgsgvf4j5RlAd
ZzcCjURY/NA3rTzG07/Jgx1nT6GkEgO2PiljEzGdLDXvfdS8KLYGTjJzRCcAFiMS
+7UPMVp9W+cPG8s8IE61B1Xk2bT04Ll5iA6JjidU0iIvdIa1RLgniTEnBC2qHsUw
f9l1KadGKISDPs73ScVoA5bKalrD8dTMm8FSBy35JPW9o5H6la5O4RoGkUHTYJM7
hUXMxzNl+m+HLlvvLJYgEdc3V0vSs0VexzaRJZDNLJxQsUwoV1Yy1A15Vtg255xh
CJlv9TuLJaOGWAxRuG6whemkPWnR3TYuQd1P9LiwSYF1tVETZzENNFjielnO6h5D
NM/8yhFXCx0mXVS+4BmnyJbPeuC95BeOqdbK/DSDvaEvpnZfaMk5L4Xsuf4ZaPLd
unQizJPYSTiGEeI1qOPpTW2yuAZoWxLXRnSwysKnfJjLkSQGaT1hiq40Lv6jyd5D
k9pESZwNxEflyD24vKDaWnHmFwMe1v3NF4D7SFnxZZ/ALNCKy7hQqlhYkXUUwFiJ
hDG0jC1PcnzL4x1FWH/UoeDjORp39y+LGuYNjn4fbtI5RXN09tiMQzRUybtnhRYG
K9btVMoM5kXp2zPfrnGwvick24+CHNBP3bB4gjIY0tMfo57zd3Ps6t86D3aynTGK
H3RXAlWiyxZxuhwEx5E7+F0JGGJARB3tBynW8OpGLl3Rgahm1+Co/bTKOTgaHhEP
xK1Cp0fklPlBoSoTU+kMEdUmNmZDI91svzI+puRnstE3ZbShJEWjTXs54+T3LXfE
IeXJk8arez3wFzqv79VFya84TrNnJ9bGiEw6MVmgfMpDzIxWWFGr2dQsyxIYZQc1
bVjYguIh+Ld+rQMbM568jlCFi0suYnxnWynCSnW1+9dQYNQmGy1VnfMny8Uj/a8I
TzbOroATKKA0n7ey0fTX/m+byvkI+4FbZdiMjMU8ABCwidXTNrS/eZZJymNzAswU
kBytA2te9hksSJLTEm84ZlA550tmEhG/PmCt+Sqz141vlLIOb5NiIrdfX1bBGnL4
f7VLESLj+MBVUW2TZdJU263vp05WKeMZ/5hzT7BQUQymWbVgQr8qw48UH8MAwf+W
kvvxtYWc0MGKBAzbZg77oLjIy8LZ8NskUpFPN2S2cVqnl5X42ASMfHhfek61tLAx
SKKzp7of4WeVRErmGa2vGsf8z4qgauYvI2zAHj3PCr0rwh/8RR/Yskd+108LWlFl
7vRF6U9zTDFbQ6ygwbybOKd24+dCTfj9sH1gZRn4ZgDzBI7qozWpN1Qn/PKrEfPX
B2rFpe8zoIRX1p8zU23xyqg6unh6jJWcp9p4gK/sNdVR936ouXHG7RzmotvDKr4A
RxsMmleFRIG1yJRAiEUcPCIs8lOHif9zJhSCOBcQlzjsaooh/4QLWw12HTXqYxKA
YaLB67onHee/iI+wGVmGqjAQiS77LpdjzW2vCaZDCm4T9cWHEj0BjKN3MYMJnvnB
n7ssqAgXThT5RD0PSpdRADw9CwTPBW9+6wON0olT99EAhDeKjWuXU8Q8ytRWyPum
Af/UpzsxEli24eHf0rU6nmEwvn3jCsbt2aqTTSfRfawfc63er7+7eFy+3lYGq3Cj
UNPpgARkV2MEXEzdG581PPIyXCLL2Y/6tbZfw9g+eixVWnka7VT4F+zCf0/2aV5x
0qAtvRd36yJuHGuYs9gEedDe7DPh6cZuoWS5UI4Nm9aJnFIwCTCj2Vdup842rZ0R
CCvza6Jx3pBJ62t9gdhV/40GyTu/tdjIhUPm2eKpeZAEji6nydMddQc42ebj0aLi
l9s2IZGrQ+R+YjZPAF1dSVnT2aLuVnsWbItitQXs+Di9221YzUUs15t0+DSHJ75X
Xffm5bfQ9ZQp940JAlH2uC0BXxlu9EH78AuAvIVFvGeBTlzw6+tXlVTmkmXKy9J9
toLl0pGm1Hk4MgW24/S7MyVCcm83ZbLXelhURqHwzSxO/maJYAkXtDKsFaNxiHoJ
ys0oGGG4JwxBPNIOv39c9epzPBOxK7j75NjYo8bBCdW1ilbPOpXgfwr1UsMC4rJC
XHYeGDF4O58nnAumy9TM9xuvFyofohFGCzwWtTDfOe5gMw+B1um2ahZdRl3TvN0Q
zfjcnQe8g6DCCMRE3ePpqK82p0yml6XUed/UYlfiRFXS6hujjaYtRGBveER/O5Xt
m0GShk8uVEDvAfF/2+ENG35IYuCt++L1Pnbl2aeTO4WQhohGBZkRuc7OPQCXcdgX
vpzXOx4bPN/qv5yxcccEpnRB64EQuAw1jYtIYGhoFlxSCfFxfzMIwCPYsJ1Y596p
EHiDkf+W/K4wmQ7Yt/96Wfo/X4mVnomB3BA4MSIc/JeRzst7OuiLVy/GJOumTlJC
yYkxrNPktHy6S+FMDjPSGb1dDn4rG4tX9MD9Yzq2howfMsVSjUOOe8J3YTJhj/ru
I8aHsnj5U8yUCjV/53hx+HaZZaigv0HLVFd/ItRtkrZrIsuM7ddH3+vWeKrLUyZw
ftEjs3H054Geo6uEqv7/B1s8Em/MzRxEe/gSc9UGmhZqdqod+Mecn18g834NzUGk
+xU7go+M2ptmCDAX4lWuWsmR0Hcgc/M134cRVtwNYkTogWA/V0wsHBMPYAKfDvfD
VIAVQN4GTDX3YalrQJCwfvDhfFU/PwOLuoZipiUjn2D9JystApBh5hZoaxB493YU
VywpsONhESwvzp0FCFKSyjnEuxacvzJ7d5AeRE+UmnQ0jGKSXEB7FTNo7jcE9ldX
cRrqIA160AdnqObBQ6aWe+vDKBSRCM3HmBuM3SbhXpIyUH5Q2fjSkvdQsNLpwyf8
bVzyO3Rrur+nLEqqhX3BgLqwGEEvEuRYsDfEVxKpmNi/nSYZ1V+kMjJT2uL3pfrp
nftOI4kpPwsNFGA+6Z0JG4m84W//RNFo51m6WByk6Xg2vLMR9Ja8bk5N1buLqRmd
tN2nVLw+NIVVYPmROKN68SLrNGTj4v0J9pmXkJRE0XgFSfcRIpZQ9GzNwNEyl2xv
g6oavZaT0w+rif6EG6hbx3q9+lpB25aJy97liOeKK1pNR2W3uYADZVcdoYU9j8OQ
AhJYKD72maiQCUqeLVlCebrTanwDbTM8bV5oLGf4WNDd9ZVTkyZWT6z83we2fUcz
DSd2k/tAOw+/o8Ly+zAHFCAbI1b/TgzcTo+SFcHWxjqxtR0MvMo2cqWMu1YHcycO
cIbfLZHPCP59Ov8s4QcDl8CPjkt0rvCrc3B8rdIK9Xh42xk65uHLrsjhBOwoPTFL
nzicixrbQCQFTjLj9dT+sqZkvvOMVirrn3c2N+JYQacgo35IEhA0t3Z277FVU7Om
sHVJL5Gud9aCY8HipKIrUi6kSAwQ24JsklUspTGDyM5nOyLLXqs7L8ePGGvoYfyr
l4XUh4Gb+7FPbzRHeOf4UuDfhiXEoccwS1XTIZX5xCQ4xvMWv/HF9/LQ9nV4fDnn
BIS39xtWusiswOe6s/5v6vfxXFf/FqQskReXmRcndY32DYlcAUoMXJAD7UJhzgEW
9ACT80YjUD9YSte0LH1K9Y0vONrJva09A+xXcOppT+t4riZXqASpMkcgaCFKNO7Q
txXeYWgNTD6TlFVzCc8rfVesJlNQxmg+sXnmLNXWQOKLlXhwCX0OCS3Nw0puABtz
uZarmVnujM2hhlUfra1ud/dk+W36XTiulkU5wkuhHbIPyiQVDl80axbXsVc6hDTd
9NP/F7JP/2rdJLnsSZKt2znHuTy3tOdv/VBu8gCIv2zPcXVDnipskf3OkSmnT27S
vglDchNQY/xedn6l6WNsIw5b2J2KPp8p554oFPNMU32UH8qyojNK6T/ZP+Onxw98
U+by8Ytqi5gvQDfW1KYF8eiBqla6OTvI0ZMGbKNV2CXpV4jbX1B+KF2DG0Zt6NJQ
pZ1rSkLpugCXUHn8eTe75byWbwQfnJgkXLPB3X8Cms2nj/UwAqne4+0s4vS2T7Ty
+0YNmhbLtftbU7QDtDDH9BVGrSuVzVeXyfUkgkXy2tQmMWfNRm+4Dm6mkVciZfEB
jQS8flfcbfUCXBZWxhmfTwE3p6efth+QWX67A1kM6RVPa5yP4HgIM7u7y7H+4T0N
ypgKLpZR78dD+5pVzL5ISmMe37WYEM4bIOSCe3aVsMd7gMnmLK/P6yhI3nL6jhds
W4PLX7jBmF0DiyX91T3KS0JvuoMQ0V1t/q71T/0FTCuwHRop0vw5l5r5Ne9NTc7A
4OFKcuafDgr8r/IPOD6J1uMpvlEUjGHB3yNdqaCc859wiY//dgXEq/+QizdjcELJ
v4Q1NDzwd+hEZLZMgNRANpIYxrN5LnlzWEuV3QwiXZ/9Rr3+h5h5JVNIbBp5yeZn
HHP0H+Ex4sTQFkeynWQDtlIwSGR+a3Vm+W9q0muwXBcqgjqnsSSc3vyPoMPvEibK
gHBhg5s8cjXZazdTstjLab0Xuduhe63GrDqItgvZAc2gBcXCc612OAgtPfOCSGTr
P6I5ZHYX9ZFLKCvK3j/K31sY6wk5J2UeRZcyDZWFb2gZ1MCniRizdcTL6ZN03Gr+
WsolSNQo4b1DTZZ2n8S3NRXLA+EfVckyMtEbuHRhZsrGh5pUrBtJbyUD5K0m61ca
tJz5Tuo/s7tSrjqrWK5wrOlBzU84ClVZ+kYKdbURPeNZkhYo7SPBseO1ihiDGjyR
Mp9wiuI6fq+/Y+acL449YG7tmtHCw+lQXazAbKc1jjTj1AVXlt0hCh3b7EtNlbU3
/YAW2Tjw1zU4yD5ZwQszos2fmKwF3ziXLlf2t6NvX2MNLrYjyfOIDN9eGNLYe0ev
ZW3ZIcGksUxSG5DjU4DPCgf/Yw6uQtd3AZjaEo+H36mXnKcCvkCLUNfVPdldz4n0
RmZAGKX3BFsDxstpivvJNAixOykZ64r0gQnJ0xvnWFnwos/0bWqoeHPS+oc9hkhS
D7trysam15nWMyCCfam4QWEibF40lbeqg5wnG20gdaoZ2eRK11TnFIQ2ab4tpdOu
tpfkn5ufrSi8sFjjPOx7RywOmMEzLvmZIYZ66j6jCWIfcQjEp+Mv9fmQTGYxpzGx
VWQZvDtLJqHK0xem0dqE6Oz43P51tpDdNDuzzQirQS5TE15RAytdDVTO1lmIpD9D
LwaZmtksAf4O6vMI1dCSuU4vBteQd8DzaevuVH9ONcn56R3ALoXPJSeIIZG2U9FF
KGGswfw84H8QjHWJknwMQbi43VFRtiLfvSfjxikTolc1k9sE5CJdFptxRdDdUAgJ
xfhLSXfPZZOxVjkrgAyOchzYNnXhQpLExWT9LEvN6abtK4anIluIHEYX6NQP3x31
xYeIOD3QdjGEiUMHNfb7wHa+AMYlVmSMYLbfP1NuuUPhmp3fq+Gc5l87IRD8kDWw
7RGZ4tzrtzG5OujJKA2Zjt/lmexDW5K5hUTnjUCwpQVertyCRlvLO0CN45kH+WwV
+y9MpPnQTku9uwAEmHDvdTV+0YCo1xeaR0Ii5NkYc4gXhjDb9YuJqEOv6y4VvUVg
/Ahcml1VMsfpuDON/HZG6P3G7CifLOytrdbh+oK2AMz1BDGXc4jqRPwluPFOVmDd
ASbTxaqZhPvoD1SnGT6FpemkbaeH5InpDNsdCX77xV3tWftF1JksRPzzCTqOUn6s
zk/Z7Zw4UON6wz774XD3KMveQuZBTSoePkxoO8EgiilmSoX3T25m4D//zAwUw6xQ
o37N7hXVg6tcx+8jqsZ7riBFdRMu2p9arBMn+TWzau+S6pYEDUimBzBsDtUgWv46
beE9U3+LQ/HzWigaPkA9WlPg3KpW/1VQFaUSVc/3KtPTQywPx4KUL3ZMVzPOm5jw
GeV+tQQwxJ2GT4/x/xUajT2gr0oO2z+bzs2lvzQqWZCiBuKfM1JQt4zcllhyeNE3
/X2kjWJoaERnVxcJVg+LUjOObmOrs3yi0j9YjFgkK9Nn/sbVoSkUUv56rRrNf6M2
jhcgGVw/Z9bhHRZDEA9zrbTGB6y8PWM4q5+D2x9LoIUu9TRB7+OxZLA1sWniuGHr
v/IN0mByhzMSn/uIJ54x7zKxGUuwcd4o5/gU/F6XXKD7/r6ld0a2JxmuwWmSqUCv
7GOeFOL1o9JRNGXv9d69xalD2/5TTDUIMdfkGInkl76IojFpK1MUTrhb57OLDvTc
6p17Jz2EuEHjKNsIb3DM74mAOKyXg7fSYvL7T5+JwZNesV46URbyiWhor4WsZKpT
vRG3dDr7nb6eygxiXnk5u4OxdMNgXTa9JpBKgtYTCtDXRY9/LrkoaGVRRnpjLP6T
oYVk6gXXCN4j/ieUtZhQyUxxiqgp4L/0d3NtyHIS5e3ZlaRhSgzGvyqR01zi/s0O
SzIHiiDmO/EpsJl7jdYrkufnzqPfCmRWocuSQQO9DHkkjmR17OX2I/SZUy2e4Izw
aqFg8qqBSUi54dAVQ3lm+CRHG8yqZGBsfeMGAQMmBNGhBb0iH8o5BXMAYe8nXMnc
AQJj8hPaySByUcDkDVjvEmACLUp4Lx2VchoOtAVKmWib5rJRHvw8ygqU/kaHsntK
83LfQAlhj7TD8V2sLCobKsgmft4sD27kMiuQWTblgDhPHd4Qyd7i6K7Y62nJ6l5W
/S9S3D5yBwTLED30Zp3IagCKitwvcr7fOhATjAXi6kD/TRTWUQV5aJBW8uI2T6w5
36mDjCDD6g2/3xC18IHORIqb758Q/Wschitinx+STpFT78OmsVYoxLJlhkCNQeSh
8/81w2aJS0ZDuFyTu84kFyKG5O/JIdIyNLhiWRCMTi6SMsnlwu/0mLQOYZ+Z4F/s
BA8sYeRC3eFTwYkmoP7TceBFtZKUMaEG9cm10lkpgzPwQ943pCymEwaCxBcIVEee
gr+X7wo4UyFMPjQAX/UUY6lvHxfXeZAC2t4KXkwBxTzzU39db4XkPpFfBgeG4PYb
mlUbRlRkl6usywvFFyBOkN+hOmJEuHZsFi5MpVnrHisqbKPBFr0jdHwmmmJhPqPi
YU1SdTBoSIyEJZ3krnS0ZN5redGcFGWezvOhNxqGm2uTq3I8+t4a6xZLe3SXuc9G
vz0Dzbr+KBLa1/IKiNwXHsl6aqIxGUsS4KvfrMgimTFzG0HBlciQVPbYyK2zEmMr
Y27XxNg8G+cu75QJQJ3nq2mdIKO/CF7dYgNInhxwx/tC/aPJ6/7tn82Xt8l1lDco
/dWCw8G54Q4WTzP2vgA6uE1M9evnvjtV4YB1t0+ns4v2iPaMORx7lVLLGczOs60F
LMh70x5k5JcP/1gP5mxCZ+O7XONR7yg6CZ//+TPmdG4jTUza0iR0/HQET2g/maj3
hKpHSdcRqC1kcec6FQo+CE3Rx1ECJW4PDlei13YEzsmQoMViH7m5PPljFStEUc0e
9fhehzdniF7KQjuNepNBfNRB8f7wnJ1ze2evvhZpHylZ+X3jrILm4py/45jjlnnV
9Uytbm64/faO9dyoQRQsb2Y5pyEB/hsV2yb7mMvRmLG74cHG0vGDtqr0n+n772cR
DCz7G6qCfAodzWwN26qdGcbs/rV0nt2Rh4tQypLEKkJ99FhvJXHxpK/PZSGJln+T
EbvMGBEjcSeB0zbi+X5lQLE0D0AXaJMWnrIEeN3QIKEq/G/T2NND2qvbf3qr0Lhh
zRrVr8iRc0D6AE3kNqtJKVZNAfj7V6bgqCcfCS+STU1Js+VF900eO4sQNc1fUftz
PjrQTE2PCpk/s7qUilOHKz6CwmE8hjxRYxtVIjn1WjVQxvgXlKrrK2QnXdAW9VKS
unO2WIkc0a5m1FV9vJZWjUYP4E9Ma3NdNsarnPws+DcCm/9DjXeadQ8ZjYwRdTEk
ybb5BBIXVXxQ8LqbmqbL3K1gsrS95VcNndwfvu77qS3/tL3gYOyoyM7Z3x259NB7
xNtQ+gOn0cpbopr7TX2gO7OxviYKqJjHRJULhpJHNoBq8Bd1Ht34UjR3S4Up4w4d
5It/k/wgz8cY8T7XsSZEt9GvVq/mFN04fIFaBnwMIndJ4Wt87YIGDopTrjEeHIV3
ez5vtvn/9owQtI+egBxH6+O7Rr3XnyJaxGICV+cnCrveA5IEotD5Xm56p+HNyxim
h1jwj1NHNiqhPXRnsJ+XONaztox9/a/93dRkkTVx6DOAdK6kPuo/wNbOMhzrUkc+
i1WZZRYtDLegJEL/SbkCK1aCVsnDMj6ZNEumgRaKKbxd8SC1KqFo9Ch93DJ8TSux
RPH9RCZEw4rAAy4Y6wVRym+5vnQBoq4KxPo/LMxlQQ9H4IX5aOUiN73HZ6REYj3F
1xUGpkjUdEbOyz2Lwmy7av5YQ89o8jmx+dGBE4MLqoOMVQmO0Yw6ooW7osSofPG/
E0suZWH1K2rvlzLh3XN0x+4O7RTajySORsp46i9jf5ku1G0NO369+CE1IiCyzZI4
UcrxT8stD2ujRNUzSAuK/jxkKWQcdXraZb0MVMjHde3fhXsNQVn+6oEmHSRtYgQb
iDqpPYiDFIbQp7OTjp2XYgDIe/Gv/XOFfJKMRpLGuEkk60mBv5HjVhAeeXQu5/AE
B+n7C6yN+W42sC39Pq7W04WDTo4RaKAE3wAG+2dAaCgZa5KarUDE+Z0uVJlhoxgI
fFRN8uN1R4AlKFzZozTSR4mUfc83W60Ef54B9ttUcyvKWSIOW3jLR+P2ZUAe1tKl
m7sQ2TD1R2yY7SDz70E3CIAjtbUFsOz3Qqsz9n6SHE9HuFEl5swcRDmn2TYejl5V
Z6tdva6d8mXu0yFA+93Of/4XxEMGEQDe+rtJLxHc/Uk0o9U8EEVY947Zm2Lfv2ei
6ky3VVaBdE+arwBvT3NBSmEsXKppMiOLfTtMvL9vc7rb3yHK9ONxWjFZ/0Foummw
TOFr7cAz0L6iffxUJgR30tGtoiHPaKGIvRg/GumwnDl6YhajcwJIpz7j9tRWiFkK
9Df5ZPxixFfKKmrky3JBHjN58HCXavogGO45FszrkGFOJ5ATzkRMqwO6HPNUDKds
/Qihf3FPJ0Xs7VXY7vjHteNx5jWOkdIwW2LCi/9mzykcIppz4j7R9sIkPLXxtf/i
VqTJ7Aoncd89HTnHUsNgNLJTHlYecXvyVF4+RrTMAI/PAeYiYMUcj/3g7y5QBlnW
auKybzWfF2vKHB04Nr33eyGQW0JtuwN4OILdCtl4uObwkxy7VrQfxJ1qVm85SuuR
JWkfK/E5F5oHMWKxN8XpA0tOUE262m2JHdnzEv3GFESUC8DMlGqzFryf4rYx+cf8
GtH1SPUp/T4iocC8SbXDk5KqwpUkS8H1Y1zhhY0Y8k+zLy1arvumVV5c9XoFKqw/
t2l/FtDAZIJbwKiJ4yi8j3Tyu7PwTU/iniXVBl739Fgbia1CBqOfRwUJ3oe/mvOK
k8Opq2aGDbaAWdnLfyVgar5cycvjfRNc9ZrODJVJi6PttA3jo3L6W95B0IwYjbsm
3sZTQpsgtIrRwKmr1SOwz1SfZ6cNz0eQhR+HC4gvFLRJ8x8YH+D4bWzMSPU7/Keu
/xqCjhXXGPN2s9g5HjrUixP5I1A7ZLmL83TpFIUBYTmvbTnNvwfNPi4uhb5ft3OO
W/vkm1sJcRkOd+sDgQfdpzZSMN4JiQRjqueup3OxGaC6QaLMKe+ONyzHx45K1mym
FZPcTbYQcQvcEMfcT7pJ9ksA2PitGkvWVsEWw85ckHM0DjIROjkl+zi0JCFXhpyk
1nawrPd6+AxDAR2qakMgssJwaw0UZWqcK/TdcA1ZwymP4OKgzgcZkH+B/Oz9myjm
7b6P50v9jXwgPXnbtg5YEwBrcc3MI702T3kG0DV4v3D/yn5ozPkD533LzLWYFPyk
XyqUba5FpHbR3O7Qi7jAOK7Ra4UfnHAo7Z7BRxHdFFund1JZ1WDGjWXoXucvCTlT
B1RQkLVHvC0G0g157WC6CrSrEWvsj4GbxFFWt5SI4lSbgnLlqpE5mHpXJMKCLToH
ePjzMGeXr6nn7+vMV9/nwe9rQxyBmg46XY6tGaS9PaTeqoJkLcYnASCzsBBF6bFR
lS5qxqZaIM9xO9Rsv5fopTRqgN9pdPJw6S5f1s6KswNnFtG31+0dYpb1qv/a8I9X
fQEpKVa5m3KBdhpK8dB8dWEjrzLu118Y1o3rErQpVttej8jU96qc0yjJLNecpw6M
s/U8Lo1FGLGnrf+NmAlSX6wFJLtBzY2XlDDZzmMFPis/tZCFBHZaTa+V8CpkRxe2
Qkm5tZupjmik+3KSwtKogb+ypUuAuZsBPJ1dtXFp/nSje/Ly+TcJLIUr4nrDoGgg
4c1q+eN1r4BIhcAFiakRQPm66j96ns9FxWuVgEGTCGPChgWxNBmne1+YK0DVpD3M
mF+QFjPCmlvxpU2mL4Rps5TK//nGk2dniHXaIJ7Edtxx65xrgwi+en+f0d6gIVCv
AlKyp96ORYa/4/auy9K61bFx6tTdcor714Q82PZxniXxv8yotlOy+xdSLQO4aW4/
KAkrMNwcY+shm6IkWiamge+GP/8swXLK0TfF+Y/sYZQRTXV2r3GLGPhHaFo66Rzs
3uChLJxVZ8sew38axe2J05eWjMqwldjgeDsSvhk14WP1dEPrLZvWRgXnY/QT7XWs
xz0PWKUrfvm1PfxY6EAHWOBpWzgZwRIlNJyrvWD6acKtoEltPoxHBHJgmupFydMj
yfv2Sp8XjrhYCmT6BFip9zBj64QjkleezJ3riERL34o5UlMsWlWCduEfr1PW5rH/
PcLssQzlBCTeG2z9H92fW+7S4zHiBzbU9WWqM3KyCYY2Fk58BYFJpEbJgw4TusMt
Hk5JlqqGl1W9CE9U2MRkY3SJL5J7dUtS0JBxkhQEZkk4yKJ0w/cKyVB0x66Y6O1g
cU1shM30pJYZUjPhtWZtgENrLntzffiYtOO3w5oibHP0v8vfL5H04EVvGizh8qFv
jn4x5At0/lqs+1vh8ldAGmvCu6G6zk5DSOZxx5W4aUbO39rULpICly8ROv8akOt/
4uIKcKFuumYuGbRcD/CZD5ABgFT/hMDeJLyVTzPUhaMB4DPRegrA+COr1MW6u0EP
EQK2xu9XUe3gtPmPp0kxLTG2nw+cLPA4NKz+KaeeERn4Mvb/MncrBJmxLt24xDZg
wPCGFiKN+hlXG9Cj+4EF8KLmBZsj65/jusdz6tl4A18ExsrOpK6VlkMRwMKSv3PQ
7TzyP+aLp9gPyl07CWqbFFx+oevc6mc4BJr3evBsJknFrYf8VSHJqXopi+78L9DN
aVgrKTXREYFtxa9OCbUfFOENX9N51n+9K2HNrMIjZLdYdNd16JvZ0qo7KaaePkDf
XVobCoFoRT6wPjN7L0GAWJQapDObRBWALJhNG0izB5WlKep8bIr9eRDpt2PNr1PB
V3VRDIjRqzIEQ/MnI0Kh3eL9J46il1dMH0Gl8US3GSfaMNV5uZS+Psaw5WZyqzjA
IJTgEe6r5PJN7015kWwOJz1g0V3Q3CSFr171NMqXaY5/ZgDuMfCV1XX/dXfBBkIr
ffX1XYPd5DySJejZNILdsTfuV7MpPEBTEOPmqdVJaJvBO6FnqsDmgzOzzEDe6nfg
+9kVlHmWj/9U9zYweizPCvLxEMKym1rIKDBfPRZKGgEyIPVkYTGt4tus0fMwJBCu
NFXHNITjY/aL5KpFfHNMAwmPN8sNgSJGZM5AZCK9jXntAvGk8Exzxe7KOrAbVSka
P5jO2EpxBcLSbebNzkCIKFWZfUJy4IJ815ixlw1BxVzsHFObXMB3zQptzq8CyKuB
wGgei9HZUaK0Sxc3RgcPb2vF65y20h8lU/ymu1vWuiFAueyQ7P2FuMUcUx5IUyDo
G+WtTQ41DrAEOqPIV5eDwq+3bDtV2kE908XG8KuxFiHVgEURXALw2Q0L+7IKHU+t
t26NDcdPQ1mxiQzJQNRjNfnpwKIXDDyCVdL1070GT5+MS9sWE21xnt3oKy/1H05l
K228ctumwt6Pdo3QAVml8FA4PlMFYT1Dfy/nZt6FHs41PwF+4weSyJ2BnjaPrXn5
TFev3jNxg7NlwXKkGQFalWSa5qR1MjiFHIQZ6MCSd1zY+G970AxNobbdKXOaRkLV
eDM11pMPc2jrmtHtRA0hntzKgW0JIL1eODSlm+Ai6uvqJu62ZHkpGQ8NBlSXzwif
DaeSL7NmoUpcS32/VYgFX5lTMMu52lVNCpVj92i7dLyCYBRMyONIfgRXvKspJThd
zzZ198IYVnvPH1lirnVtfxoyg+lS/fc96CdxsmxKCq/w25uFE23QpyQexAQB3+O0
GCHtvNxtesUF7S8+vSwCC8+eq2lRhbq8OGOItvRSZa1nYuYE9nAUXk9P7uuueS13
80zGYlmFEnu/fniflT7j772ERlkGILeYpnD9zz0HHWKIlD+SipcMleGmb30EU4+e
sC+wvOaTTnKeZstWnHBLPacgXAosv5EvFl11Rr3k/oS5ynM3XFgVgFeZkO8uZ/a9
SzD5n5GX2G31+IX51xG3gUFZbbamxZ+tOAjeqRgytA0JxF9gcCIjfAufvFsVo83E
bVIQe4uN6KvExES5aXZN2kz0xJ0KQJe0CAMF8fyqvyqZ5TXjpyWy6TKx2wvVkvb9
mNiZikaoJCqDuQnanYUwZ5DUSWJrEW1m7Jtm+OqdYdaXuH4jRflHRmSkK4w3VvNs
VsH9AczN75MqXjjxLgcpbR7cAvckHaSJrDAnt0aswRmSC6EnQ4pLZ6jnaBsbOgN7
ipTs4O0BEdu73Euf5kbkL0ScjlAP+6CaBcQ3qdNLu9hsDwHz0Q7i+HQXy4t0/OOy
9t3x6Cpk3odGotjUxZYqVC/QtK6nnkSjPg0pI+fi2OblEvPTmU0zjj/eh65cz1PV
QHu5v2jz+JwEqppS+QG80KqHqX/mzvwqa9ZaI5qWEejMYjyE5KxzDSowYJ5igvZf
ISfe44dRbcknpwzZxEweBrDXhpzDvsB/iYeKIHRiSCCY0ybEmtUCeYogifGqnG7T
1pKTJ7EyljDI2H4Y3tJ4liD0SQ7voGNiPApPYhWy0z/6b6cjM3xhVp/y+WVUZsdW
asEJlI2Et1baGUc+C0axmxXTkvnotsypWvIVEGfTPe7jaUfFpLW60KIDcTulZhs9
pmiyK2UhW9T23dMlCPLVdz6E7ykwXk2ELF8IQfDVozKUrKGNavFEOPULIDVDpR+l
JPg0LemZX7hfRT3J3BAyVWU9IoHPfoaKQKZJD5QllV15y757K/Lh3tcNIaYx7Fx7
R0/ocfoIMqa9hMGX3vNWD0F3c6uvjNiCCaAfc4AcgRrhlJj3IcqmpuHq4liLXbiS
0j62qdDFOMyYUeYd6SjqPnCVnkhvqVI/zaAGPhmuL1h2duE710l4x8dXffVv6Oe/
uNbTyYp2ah9KpG+GR6qdqYTQOjNPGi0m74qwbeljvkYBmE0+zwz/hojLUU+j40Z7
bIc7KRelpeatTwHf25Pb8D8MetGDXY19U6HTjiqSLHtiumy1heIROScG11AOKW9/
OFo1L/RO91qyX8/86I9lmWYUTVHp3X/Wbf/BIIKsjfY1f6hVF/FVb9Y0PNzlftt+
UA72FzObchL0kX0ikB70CjhjDi1yHravOe89N/Dji0lDFLbxJlXywdS16PmFjzGC
b93CO3IDsr8swv2JNt/e85CsSpQ7xz/l5cDH9IsCu/HPxXnudtY0G6zKUgKuBIAh
NVXtPFMH3pqh8yzhsFzrHgMIS26A0RiLXuEFiOccEKDmSWx0gvvjhytzkvcRc6ce
wqO+FeTMdPr70978tmc15qhofa4mIzumjZace2/p9MQ12B9XveYh+/H8jtdiMor2
iS+kEUV4jc6TxreSmYpCItRZNWnJynlz1s0jXg+xD/7BdK72GHT1bR4buOnTL6vR
ONweBWVh7nNK4DxRvpoWdGGxlnSAEBrZC7Lvhssj7k2L4ueTTFuhLynwlqDByaIb
SvPv6izivAQ4ZhAuIzUqD9GSsMutmBARaJwBJQJPnnF3h85WhHCqOpb6lL+s0vz1
DurfTPZwZ7PqknUtfuba+YrIgqdGJvPjmlJuoJCyB8cF+nzvhsQR6hjl6SjWYCrG
SSrKff4XRNortRARrm+j0Kfsti7lxv9ttvX2XMCXfEOjje9HK++X8Lh46Sr7cnUC
zp2yyOZ/SVdt0R38yWuQYmk6k5LBb11LkMhk3QYBWX34iQ4qmpO0MDk3t8B3dmv/
qObbm2zLHx6AUkpJIuBmZLri6heDiGyhr4/49DCcxRYJc68uHN/pdu1gEnK3Gs6R
MGSyzwFtGzF5LB8g2hk6EGUU4y/3NSBDMTaVGO5fh/c1U4eLt1HJCUi5fGkCKot/
lCd0sMXpIjj38WE4zYFWoNE6RN/phaHjGxThMRibITjAyP39mNAyDCvoxjL7Q+g7
jpRB7RKwZh1eMCYm3R86X1jlFRnBDcDRZqdHcu/Li89A+y6do4FXIo/bIfqrh4ts
QpVXD0//fhK2C8n+87GUckU8791dQLZ9993cSFidgKTrj14UBipeeFi0gEpWtszC
lWsJa69u7ckPvn1QXm4fsuct6qxrChRp/GvdOqMZ4wg6AiqDV5iA8MPN8v+WjZYB
fkaum2f3tGTa/sQhQDpWqNBHowtNURMJgReqkYT5i3gFooP/bIx+F8htL/GMO4Wc
bwhRhBaZUoDo4UiuuJkzctkeW6Adh9JiA56ZNX3JOa/eBmbTRkvblh5qG/uQPQtJ
BdT1IVCGI3HgCmx66ABpzD0+0wcFGYwY9mMMcBAjTDbEYiYTN1z3rmm7wbUafH9J
WemSioxeUTWMIUQ5SWw1T9CT4eKJHbDBdXD2lRqx1Ob8Pxf7sMrkWzr271Lc8JXL
Qy2ToY64GaDlNzY8rUssvSTF9NMaCkc6KZxuOyTx7EvikKhgQE3Y4yJF4zAYcWUg
3hOF9fqXFbfshx6y3LV4jP41y9IP1BnRRRUw0St0dIvDGNZWwE9y/KRK5TWDCrAO
ddBe46upKpT3TYzaGm9aJOj1TZiAWxu6OO7QOzxeFgB+xyM9QbbNjfhYDEIKNgKd
Xflpx1mDNQKeOeD4lLmOaxoQqAbpzHF9XWa11EW6gMoirnrTlxaOZMGQGyjTOKQ6
4B81yZ4hiM5eV4GVaUWSp/WbasN0oEZR2Y6i0yab680NniXMipQu6aTJ3JC+Plq4
QFng5+LtvIY/tSzATf4Jp9APg9gyusi7LTL4inkP9KlAmwoXJtBOQjkbtpbWTUy7
toURjHi/zUhaU3q1u0F8UetqpdGKgt/7hgPZUufPItuSBlzYVEe+bKI7Xk1slnoE
oYSSMJ0vfQMIcmijwQ6k9plmQRMxVwYMxOCy9oz9iijQkNzCij4u2vREQgSnBmu+
gfbdviMnyXhbNK0K5vSU3Ez4pC/c7wis6kUIVWfjtzDTsMpkY/7e+4IhBgLLCYuN
RDcsm96LZlPXpGqUsHTiM1xZIAhdtP9bqDMZrrQ4fsdek1/1T10U4zAbChvcdoyB
f7wYiQu3wHAku0tKZIe1vJH48/qrq6QbWELJ8GONAUu/d23LmYFcXU1XeBajq1qm
a8CKgIWrOHG4iUSWQc4TNPFNXP8v2lPSyyR94oKClT/yO6gq4nq9GNWJMyHCGXz0
Xcx5PK9x02uMdzBYG4bD3Wl+0+v9tC6MxCrHTD2FdFtzMHq82CIuaOeNtAdKyojy
Gqo3Nl4+JpuR81jp2QkAZ5Easw7E7OjwFpxOlJYoqC82iCiXYi7S6+Zaq6o4M0mt
vUSktMloiI1+Ema+3TekWJXxdhF0hep28W9LeKhBQX2Eh/R8G/o8hLn0MXkO9rQc
ml0kejjNPbRlxVAo9agpt1eP39umSuyX4ZLvIKrA7FlyGt+xyhe2WBYsLCArHDiO
gxVcDyUB49vggnq0jEFcITW8ZBBep5W/PJ7zEm40lvUEA3wJoSbDoQYD3D9HDWMh
YZbACMhjnCqPRAS2veKiXrpsQh6ZnWTO/CKvNqzNzog1vL66U+N8QvT3J4uPoOQU
r1IgVRN1cEEklY5JBMOfPybur725+5mwx6Y07Nz4+pG5qK0HQk7ikh8qCAkBXn2a
2fsQcAiqPGBQZZOwFe/t2f/pfbjwQodLifaYTeU/Cw7hixBcDv4EJ3OC4t1nzqPK
5CWYSy8/VoZirG0L1vIkPO5alE9M+crFwIdN8tDxW01Uy7NIUvpJwPTqJPSw43Z7
dDnzTOIrcZK3UQXL2YVhl08LL/EQTOpNLU5Ye6s7zd7QOdam5yW9Hghgu52CEj9r
SS/5Lotqx3jKS2hwNvwuzTNJ4b6sh0m/OAub12n+bu+ftA+FEk7lLWEimXfrvw0Q
AiKLul0CfNz2owEaXxmXkllOH4Rl4zUxV+JJiPXV43vAQm4gjKeuHz0gAMgzx/FY
5zxKTvmk0sJTkENrmHE6K3eXrycsSNBtasUJHP1reiRZ79sYknLdtcw1kyjIFcsc
gZyglRaBpka4iu5rDh9EqV2vxAaUc3i329xdg2byghiKBlGTnfVHBhXUueBcCpb3
yWLg2znt5GUSmYcvjrgWeym3k+cwZy5FJ5DIbEjGkLC0qyBHsmqDXeyEL59YOno3
rZ/3f4hbUCgPITpbY1o801aBtBGAKEQIMnpF+P27GAKE2cc/lGRh1SAMWoMW/UvH
zg1I4UCM6XAJAE/qqiJ+GgJY7KUkkB+6xoQyNBRtw54NpR1C4JkGRh9gUkjeamVF
+5YG041pscKZeDedNAfJmq5uJlt6EtqYbAVihEAGTouZ9/vJvDiOSRy5tNZUWHQ2
6coho1O41R/pEmFcfYuKpG5ZRijvX8EQRn/4iTSTFKj89wbtJBHAcVYb2TvoeqX1
5VKW9C4b1Yw8Aq812yC8zaWbMsCBJ/JLyJ7Yi1AjTUqWLLhNNGVXX0alQqEWwr7q
/uR1B+WjdWczqqZvqpb8H5jtb9o1gQ32JQV0kMNtrPu+dYdVONhBovJS4LkIakqs
FNTECzBOSVfQoS8LXMlKSvdP/8ZSRnNdvR69NzCrhXpc54WJBw6YljjS34pWELt/
UQiaRYQFxmWUl5T4TInRZly9DT3TGdNGY6XTbGC/gLUm87/cYoYiW3mSqKbCgW0x
Pta2ihfnDe16qwXKeaWde2/BHV8NfqiNyZXPR0AqDtk3bmXd/TzE+7Ku47M9CKvF
PnEcbyw/uynSpJwzkM/sPm/S/LwJxwu8kOAj5SxtG3ighaF2CXbSvoxe8tmZ5fXW
lyL1fWMTcELfnLOxKeajvDbUU72xymzSex6tilQ+mCeEOHM7FOjQ7x1McPgUhNUw
xJGTvXACLJRjJLwouCDA9bEx2ExnqkaL/3tPKWqGjSybzmazLEYuEj7OcyKarDRu
gJdbvVFatHeUW6T171uZqt/37naKqkAxnBMWQAwAIseBGdihCn1osrFV65jVtMJQ
OvsqJkKPCo5SBRqZNQdDCxr+K56C+cPrS1sw9dV6V7ho1NMuS03cvl4MbtTukNDz
kvUsgHLeC8qyIRMyPgdYTAIKPbBwMps/p4/gFCz335zuqMKCLWpxtqEQeglJIlxp
Z+56i/mAnVs5oD7h3faiFvA+5G8klVUrL+70g0aHAiXFN7jO2HJiQweuDzp9AU1Z
OHnbFmwKCgHL/hYHjqH/5hcxqbpATIYWpNQ5/+GLoxtf7YpJBJrb2QICfZN8+iTe
1jA3aoQCWBTd6sj9SKaMbzGcLM8T8w2ElP79nCI/YwCr3N7tUDP8jk5KrGS1TS3o
S/nmZyJmqUza1Or4jf6Iv8CaUYCO/LKbaAUvC/SwYCdi4ppOR+Aj3eIl7S37j3lx
z2CtsOLSRqYA0P/2agRo1qvMqSI6Bbryp3kXeC92pKkAu/qZKSK5B7rKyOOwyrx/
tdlskBpFA8RB80TB0PgZSiGL7XGOvu5XBfoRS9d9C5F+KRxQpq93UFVDAAiSY5+c
O0GTSaewj25KtmFk9NwbwroYY4zRzeBW2Br280irQfu8RLzFST8bi3eh+cH2zbIG
w5z5cFV/Z2uM8ZsUCKYoc0EvaMpAw/H6JC+xw7cSooND5YAupnvseS3GkRsuN3uw
IvbZ4AUTGM6q9m0iRVdr1wxg7MNoBIvufjqVhi9M3HW2/6cKCNcjidJnN+uy8CCq
Z63k5BZXcpDCFoFhn5H4Bq5SqoUvE8aoY5yDht7rq8NsYnRAC08Be5Fnt1KPM+du
AvQkpdd/SngT6kfPoiQFDSffUtHxcdmwOVmE66J1vBvHrkua6R5igVSLE7WQzxjd
zaL6hLBQbcEZFaaKSFEyTimKY+uDqQGSCKUkLj36o5nPj0mrH7N7uFWwi9yhWfaR
o4vN3AtttfGbWSmWIn/MvPAr3/cSJjsvrEpmLs2m8t7GAC6NVI9i9bD//PEt1qEO
X3eN6h0ZFaw3mzNt3SRmGo8srW98lE9Nc8J3Q8VCvv830US/hQ/6Mq4YYTZAPr3d
DIJAQUr0/UO4bfpHsPYr3AQai8XzInnjh4LNJQsGMrp+pEdoW5x2QZ+fd9VKlibF
Mxhu+yluLNkye1sFAN+uA+XyCMWj9VDtqRYTDo/zxgFpKYQmSJ2S4ml6FZ0Woogn
vrTSsQp2g3ej8/lpO/J9IoH453wyWotXxkLttME61M0hzit74oP4VF0JKr7hyBbx
nS6TVnE6NxASNEv31MpLtlvKmvT8VI06HqNbvCSwKWyMeSZlRr55OEJA48ARASC9
hyg7BrudKb1JNsLkOV6kXzVWeM4Ufyo57AI/+0RPFcjC/+/fITTYo3i1alIkQlvR
S9Md/NEgwicVI9nrqfuTGog3CR+URmRLZzovTthDnsm6OXCt0ufSgNJLxa16Ce36
watwre2P2ggAR2afU8WBhlEbGG7Ykidt2DkIo7ydIpe6VeMBYhEACKzIicaR2JOJ
yaq2I1BCYi06auoXAGpSxcjsq97uTd8Mwh/xebTeMKx8Dj8Bnebi0b2XEY/Ztilq
mZULIH/hCSi54yRHyVDnwbxnlF2iammlgVhKh1Ff/bVvLzyjqDMNhTaHWSEzEvMC
vYbu6XaWeINCZJv7RsN+Lx6RuhbwZC/cIxf6lI9a3D+yLWnkGx+uDVrlkPRzLgDI
yRH/Nj9spyl2MmmXiVfBF5lv8v+oKXlABSUZ4d760jbsZAXyaLITF6D5CGVqeWz9
xmoOgZDxVfGcuOPHBPsLgc13VRGbX3CGjZbCihIWEWfQEMajh/YaN6+AfHiy0Ipf
5kJyi0jyCFYzF2eh3wyEySYhb/zmZkFBd96Iqiqus0zIZ2e8uYGhGsVk/QbuXMJW
fdzActJrC/nJh5gHaDD1ikE2a27zzb5Mz8dUp+YQFWLn7Ra8IVAY/UYJttYh5yZu
MqPH04hUnV5Tzk19C7dMXnGS8WYPwe26VzF8sRPkoWVUcA3pu9WzDC/ZK8ULI0bo
Vaz8sQRD/24VgzkaaBq0+e2A3d3TZyHTadqC6GG80cBHiEEOxuvL8nJqhf2CpwwT
oYOh+Xr7QyRIL2/AdCh7GYkL6uTNlKHS/RMTCkDETquZpm8MeFnh8SaR6YfuerZs
xJ87NTjDB+Ugtuv/QXMfS1/Cwyaf+Gb5gJZFWNm4l7/laqr/8ot7KbmiOmLfsykj
tEMU8BN+zzEDv78XdnsuMz2lv3XnjD19nIH5eLDaAO1T9hKbFb/MpYluyvucK7VP
QCRArobq0GwxyD1IcRm3EwuqrJ0eRdT89nmsz9fswhAPoK8pvVSorCWK/aDu42DW
g+JKnqUh5wunK7tsvxV/opVfRhTYVQL2FCjLlrwz8PU+YN0dib+AQ8Q7piGybDgH
8NBa8l7A+qfXMOkDFU4aSscRAhh/8zqvBBHVWcR0w3WENltVEvF/tFVwdxawO8EL
GvJwItwM/3L5xbUUlf6xSn+y49ZL4kwg0ia/FfiRS6NmOaiQRcs5EV+G+nGdIevM
7G/bc/O4bWpX7rtRYWxe4dQ1CprNjMMJwxHb/nETskLppGDKfK10mR1oWDUxDG7L
eaTNoQmUXIIry6h4Tzv3+R3K/fbVS9CNTAvzCf2bO9XOyrbWVr+bytfMI1EXizf4
K1ub9LUZrvc+nqD3WgEWKy2e3rIwsfZZFd6bP8orppOMBSUs48HRw45M7TXjoScE
j1XLnEgB0/rkh1SmetRmhFhwijTUkLBL9pN5f6X3/E7xLVCNh5MdaNIAaQvTsWvo
ELhyeirnMJkUi9SwrhC/hxrzsUjmbw+IatL1n8rG3B4uEo+YAv77/w4TxozLTyl6
REFYNBtMM5wGwhwcoPXY5Gyd/CreCPbxjZtPGTg8ddgLu62O8vWx47mOkim8Tkld
WDVcNLV9BECH8DfXlrhvX5qIdPatCkyhBZVOHhUR9JJSP2/exAfUfeNqid5dPXNS
MrreBTnbI1TYrkmSS5xeYXJOKydrVDrbWg/EyCLrp/UO+oBjt1KWRlSGOHYERuzj
9BaJ5dpPFLPJz1mrbhrN9Vnt4Yt/VtMwTSno+VUV2QjJCHjVMqNpHt9C0uRvNhlc
DgDRabQW9ZqrrXutOJRUKgVoel/gQSoYfy1qSup7BJ/DCQuOdtZuPazity+0rDyX
uhcyJjIhcuxz2QUeFRGC0x3GOpUFrpJiEf1JtnGWomnErL2Rno7KbZfsAt5JMfuH
YB2FrymYZDArfXahmqUJ9ZTffHXqh7q7c1aQ8UKpLdqzjqxJj9ocaJcF61bPqaVJ
JwIciCW7yyBlCydUCXr9oyG+cfggvY28M8h2zNkB+Nj/UgZzdXMd2mK12kLwrjN6
LS8UraWJ+nrKGi4nqCPky4oi36164idF2dHjjQnBXkoanRXF0KJRDeSAuzhx8L5l
yBC44/EKWrCB0B+aB9VWK3vgUF9s+nInOdd5h47QhCNlTiT595mBQMy/BXvMNbmA
6B+keyD9zICEBJoLemjamJ6Bnet77TtdAuPfCe5TQbNuwNm9t6DnhSB1lI7wSf4Q
yNgJmGUaXktj/qqieyrEHq7dZ6JwfE69P+8Xqy8CQsvsX/Kc+BT80eGgkHAWozMt
/P/3ZOcQwPbRsO3uRkC7CYuqAVNFyKMG7G26cvkHyyGLpi7yLVMc3Djtyx645BH1
DXFZzyM2ZvGKc3jZiGjrATmajiFezHebtwarnS/BmywrItuvA96stHQz0TaO498F
IjULoep/ZpqCQM8W0wLhqhTy3KGyRmxyzkne0ty5jmaY6eOzRnxDrGmp1sokdZsQ
TVtYyFpLUF0jaE0WFO+9m4bpl2r/wHtos0V9DzGv77nmelyd6QEqChAxPjjxYQI9
A5UCOQcJO/QBk6lI1uHgmBqqABQb/VE6RWelPwXcOwgqko5aUmNdYTlNy6OWNjfL
iuaHcNC58D1b/UzNDZDYOnuYNTk/JprgqC4MMKA2In5zSnsF3cPyxUXP5mYTdUQr
iAjOaVAiuOALEJyE5xuOr1v3iijeZ7vKWl3C8xwVuxku343lLnQPqq5zR5Ae1+pM
Tysz8b4tyR3kUketlYshNEY6F+af6klUJS+ULa6ZHeT1S57kT066ktFm9Ah9sQFD
6jN4PwgLM5YZCuOMR+sNTvmSu7qVJ3oP7s3KYVo0swdPVG1Z+Xt5SQ8J0i83XQRA
atMYeYEPbt2JOqFrPY7IQzhTilOv+iPkMtXjEVuHYKgVCk+qZdxANAbKj76j4DwG
nuhaeVm09PBhlbkXCClf0JGkinhlRTplnPd9FWFZe226m0sDPeLHQB46i2UsEEHZ
D0crSAR4DZHa58wrlrTMQBV7416foKHxQv6uCOFxEYZdItvlEums54TfGdBZdhsI
4HjJTUSsVxUDeinakfy5S27tDhO8HVp+VbRixXVIcHvk4aRYJtPC+4Hty9iLlKxt
JIxSUk6TjHtroumYHYBluv+gETfwQ0kV3Sl2Rm6+D64UzZ/m+zSzXTkT4QuFDikJ
iF+JHECzqAj+pDiBvsld4y5+aHLR1RCQzHsoEAX5+pIiwTgzZoBATZ4sLV+4u+oI
8Q1NfJW3RIcnnt9AcUU0soACHMQGCqVLJIuWEy0WgTRlS36bCAI2NW43aLDy9DDi
EY7t4snlk9DqQqZKnIVDuupr7lGAzQ/b5yD4Qfo7qyOXhGBz9/r7xrcfFJcXvCf4
H9+4eZ/BxeNNzuNZtUPCTbOzfMqvTK1swnxro0t4ul2pF/rUR6k6bcXUfsJ2SfXk
VSO/ho4ikvawvjbku8gpgmXq8MGgjZz4TWmJNpa/j04fXRU0oH3LwWVodemgfaA6
MWU8RVppCOX25KHmy1VzdKuNGcaH+FUnmq2c5FNRFpzneiExNVcMPQqpoAYsTWdf
9mkFOQVEwRl65x+6VUYgOmdYG0ZcCj+i3LtrBvLzmkDKFFMLYdynbzDSHB8IPwc3
QUBggpJB5Z7ONQA1J9BRos5xAUdpdMLHXmXq12g4sLzdEpXKZWaGelUhpVfdcygc
aXKaY8emPFaqiW15MohMxG1r+hykXBloe3wAu9d/pWI5WyLtfe5c94i8X8+M+Mv9
l5OPxhWATuSF9W/TtK8szBE5i48QdQD+gNjJ8Js+INJmo0HUmcHp5dTyOFcCzCKC
/9V3vkY8Om1oe7viWfUubpHNGzmWv/gfzuqjZgbAj3rrYkFR7gv18woOHUc5wNA7
7tGOF0wD0wwKOKWhrI3Xxo1Man9Y2pfBpQx1PVH9JqwYE9/TuNsZw/5Sq1DoL7Uv
ixIuijeQsBK1bhJUtLRmscikNSjQDRMdLZ50JdkNd5fexUkyPcUmEML037oroz8U
BKEF8xvPt7rzreY3+eQRJsohFVFosmKKZRu7KR41sLySWLqCTqlbgoCPgDhwIGFz
T666hH+nXLts5Dj0SZlQkJhhqsoM+wlK2pxn5/SfVQduwEf+wolWD95He92ZCY+f
cEIotDgdguIRd2BMMOnhCC4WAfFG2lSd9hVpyDNfuoetsy4kx82pKXHwbyx9IAsH
2h2OsA/PD5GRXQLF0+2DXNTtMF0dQQ+0YNTsfbjycoDSpueoyrbEi0Kny2ZHauJk
7Nodrq7iqajrc0Mh/GHUD44UeqKgVJ5aMHbF1qARXEgfTUhbCr6cZMLKskwvURXJ
jTgpE2uaYToAyhyEovxyeJiCFRp1Jt27Eg3c5rf5NRvFuvWVr22a1BWfb0ryiTKE
yV5XXk9NnOOSl+U7JG6eVtRWv/WwpY8nPXD6JM1InoWriGXzv7zM1N/im3JkM9nd
cHTvXMhH7b96zO8w+aTmdPeQRx8zrlC3rWwcwg07rnRoG7RuaNqpzmcIluCF4Si1
RdpEraBB+CFrHZlktdNo4RfDAeGzczyvesLUC0+a8iNerT2LVrCJfkBmIJTz4a44
z9UfZABpA0VXDujm3/9csquL/cbfq3pApcskk57kFJtK9eZzgB+OayfFhJ6rW4wZ
U+5dxJhMesOvmhdPUlsrRKYJPxWqCBMMw2gWxAsmGWTLM4tUhBc3XHsiypqkR3Xa
oaNVAuUIZiz5pqg89ytSejrNLl188s4OvLH3wxyPQtDZGPBNWA4WvuTypgPgnFJM
GdB1Im52MQIuP6HUQ0wY2zVQKnxlXIfaiDOOgPjSKnfSrR6i3V6y8yQpiVIkYZXw
zzdFuXQmvsmNnMx1omkAD34Qpn+nUe7hNEzOzRmiJqTNd/jNke+1YxJnesYrtCCF
kjbUyjpHFBcm8U0mr8TepFmiYFIqkFaSt5Rd1MHvtS5SYpIpf3UU71fGLjFMxm4l
IN+KpZZI/Fmz/Zsq/1yJZ5bqSnycLTeMmx3jK6eS/6GwqHDjR9YwQ4jyH3gxzIgp
shUpJFbqlDhq6Cu7hCSdjYkibRj98e4bCXm7z3eQNl1xFKKxQlOiWY8ezLlen/CB
X/gIzhGoe9jfVpIRKV1pMmbslzGq4JolSW2+3A5WzT9mFhwRNOzFmYNxjpIj+P1R
CxE/lRMiLQBmDPzB9bXrwGgKHbpPUjnONGItVl3dkGLSQ+xL5JERFx/Pzv9bAnag
4WEpxjH5KwXvKtdkyIHS88OvGSgyERYsciVtAdlJ2NGjB19bMfdiFl+wrUeTWA+4
UIcvuWcpbSJ8/6hAjTX3Uf7GgiFxnwZKGAsRPeHNzrcH6NHTyCF1JKoPx1z3sHoH
2Jne3CgD2jbj5UO8FcDDS2w0fDqua8hq+wiyq13NGlvNCVMMyAfJOvKZHpS+r+eb
fmO9MLzuZarBGvp8o1xIgq1HOb5YeURfUDXVaTFoo32AAHCeXBvCYM59I6/zQmvp
jiDTuXpVUkWL7QvCRUU8ScZjqvgE5Ays1aeXEsb2+4CIX+gwbEnixxUbSsi2BEmq
8neQOlnW2fibRGoSt2bzc/1ONJNhKt3juPBxOk3WZ+sjAauc24xfEr+Z7+AkJfQt
JaVV4/JOTk8KrE8etVTzVsjCIsxqk+EnlA21lU9NYgHwdLjXwPyJyHjr2twe+kF4
Nb6QFFX5PD68hH3aYsoTPjM57ZfucW8qRmszZs7nKlv6gjxtnu3h0yzamdp9jW8H
ILS3YF3acbabGxtQlLNZoU9XsEy4Be21Tgbl+nrY0vaO+MiEiRm9hcooBp3hhlWs
GqCrHPFIWhHBdIxnHq5XFDmebWma/Mf9UVW3WCBw3ecYW+LGJbTNJaHltc2o814w
UQOAxBzCzrhaJX9I3sA4BW0WSVANUa4IrT9Rph23rgbZYyP0oXnYHKOjGmYKfCyV
CV3pBr1V6xHtAYIg58HNVszVQuq1TgJg1wrWCXIf8f78q2RPm6Ta3XIh+SuR324T
3mRNa5YSoP8gK1NI1dwIbwX+3BhEUduRfNZeNdDRyYbR35ekWlQgVawqDkq2P0Ue
RvJ/hmfcpSDJ0PTn94+6vR2NCJYdZt3uR1A0IZw7B7NVUqb9AO3bPeEfZG+ZUNvu
DZkw7OBm++/7no/a8T9nLxu+OoLI0//tAmTTC511esEKQYYNtiMaCHIeNQIk3xp9
8hc8tMWDKfdkksXc/zcb4IuQaG08KpzXDOL830PKf+9xjF7mrx6H/1cIXPmpS2+6
1fRxKgwTkzFXFTI/xp9vBQ6MrdW2D3nXI0SmO1isLWVL10HA/9L/9RKqzljNQZbn
ebi9ZfDo+t0Ni5fbX77ky3//SWQaKKb/8pFP+NglrStdqxXwBT7rBquAWQtGyRGj
bAKwipPJ8XTsdx1ZXOfpeXObCX/62Ogn5PGc/P9JZMcd40zwpX+DcFlC4Q9aYkZ/
3QFu70H/cx2t6se0QXJIB+5CuRApjH5RF+wwCJB9+g/S2BHe1SKMATkitybJe8B1
/+WGTIBXN2HAZ0zXSThmc1LCze3sCEPTZmBgnn3U/Kntn7HXo1ptirxEZyrSl60l
2L5WmZvCDtQ/JK1EojG0kwU/FH/EgV2RTYT5q09wq49RZD9q3/fJDqVBWb87vTU6
kMymlpffz5hOaRSroBm192cS15V50Ht/RxVJYPRyfvVS3oAbOqB3q8BTtYa4h7Af
UgbUxxMD9kMqBmALb8jyvHKUwBL02yR/VaJfpYK448QF0FVgPnV/Xnn0fOpAwwv0
z/4XYwKTT5P39SSpA2ayiRXuyKKfikoie3g7a2PcELHlNy6orLSfc3e0dQfx33V1
lbgjEZdOzx4L62HEqxr99nIpR0274Ahas6V4Uf1CjMXVOZ3IfIU+OO5JUzIBEeeu
BEn0azNJgzQNz+zFxMs+Ahufb6ZtNtrmHgwf70s9O1+tsjvvyvmboZRChZj8/bpH
kt7PclQtG6i6mDGUQvjgsD3rv5PYqvwOFw9D1f4I5uX8K+/TyYwW/OWQdo3Iz07U
b7hQO2IkfZTfWYn5G1JvRtWkXiRfzHpqwYBCfzyqcE3z8M4xDFY74PRfTrNQvHXd
/O9z4zjfi2Kje8l7JE+lXaG+YEI4FXxl27OBPAkKdyiJhkJJKzvLV1Akb1HSfEc/
TJxZisoI1n7Ksmi3EkA/V5HPblbuXmfSFF5iOQlY1DU8a+QCrGy5Z+f2v9WGdbRk
B2x8xABswB5W3z4t6JGCYP8HEdJoxv8rRLd0ktnwjtROPCkYQDbIgTz3zFz/CSKQ
D8yIP0mFvG2Rwj9RtFxoWsZse5I2+3c2zUXlj+7jqE3WGHt1YTHn3ypfa0VOgLdy
jzU0Bq+AELyfCHTFT25kb97D0sn9PS7nOkUGTIGeDub3xR2ThL8NvGZ1Cahhv/YY
eSTNxiLX/6Y7CZKkHH9CPpgTyR3wu8NH9tNl+sFmp353rPkM3bmgX0oO5nkiO4hX
nBgVbF9Az6KvCjImyHa2mKQrxEszS1kWfs6XeROXsrpqRZDWXmz+CLWoP2JOMu/3
okESyI5+L7w4KXSV/rGY407Sg7NkSC9GGi9Ve1LfGSpowTev0Pprg5k3d9tZRLXg
OURMNPtohc7Oq2ufX0KDTAYcISlWRmur1naivnFk/Qyc8ZbzCcy3OzydYOl2tpnX
Hg4NajHa8HqpqAUKv+PeqQpNEVYcfXrdMy2bvpSDY7DkVoCaZHajt+Vtg92XBEx3
dZyJ6CC0YfnQxVwocWnEHcCw/2nVxujc3PP/XYTONi/ChrlZJSH2XzOo1DohMoS3
hwuMka+uTj4O1bV6Lfbq/ts9Hq1suiq/MgP5AMCJHkpxiDwwiT70AJZ/gK/pdCTS
wgLw+6Cu9/MXzLfdVmbaGCCtxisS2uUf2EDk7r2DmyoqJTvFhXn4gBnEZF4cbIwA
ZwkLUCGP3no/AVEKMApR1Pl5/zy6BSQfbA9g88SmmJGEmeTSQ9Rx8ckJEC0d24kL
nhYABFWPlyr1KtGymmrA3p6BCHrgjpk1/+ls12kJdN4Vw0+yZHVfNXDJXjBPSAiq
RehBuzy5pJzh65FR6nyGVLx4/tk168phdJxl4ugkA03RjJFTOocVNyby1/BeWaMo
A7Nl8LFx971cP05zw0Zao1wPxH1peF+CWJ803zZSm54K2zIl+wqFn0k6MqsY9/WJ
L0F0tCZksWBRCGA5N6fvXadV7fQ+Tc5PTLOfTWPj0u1vyybVnP5LG765foJVctax
PNWF+UzeZspRrR2OJ7rqpEJDctjeYFycVb+S/WNXvAU9U6ZIQek0iSWuAiqi8D9z
yPMGK9gaMzCXRj832hqul3RCFo+V48TGeJIZpz6UYdiiEHTuBINtFEjyiegttElp
xqhKkYx+E4tq4iuW4iki6XGrr5GR21RTDRdl7rVxooxRijQ8sfG1uVCECrjN3Ey5
vC3Hdxz9MjDiJc1W6DrGjUClH+zyOgcPWvwo+3ilQ+eyJnCVKOO3gfZbsmgE9r1o
vzE1I3E1pIK9ejt6tewvDzMmdjJH5tPWueLw4WMgJRQvEN9Ykq8WhU1PQZ08aOkW
/PuqLd9Wiqk4RzloWlvD0enCP0wQ7tCP1YQFV/gMsQb+R4qjDUVIVwmeIpsu1gF0
y+cvkKJ75hoj/VT//OX1VJqFWZhIRTabx0F2oDMojk2tHkt180/jx9pMwsaSOOTE
dQ0dq15PsjejpsaJoj3dUUIadkdU0WlF5Xr53RgCXyu6bIKL70AXNkyjO1V/20I9
DpDGxbqAzvRsaUvx1YwnwC+8V9icfauJBcsor+vAo0Q/EhjyVmTyNGAAXQy063oc
uBB761EEaNyVbdChFjAPIOHCeyLOhetD7nTm9y1n9Z/gLVFSDm/xo8SfrSXfv1i3
7yRHAWsbKOrMIGDKfMItbgbYT3QToN/jj4Aysp3vzmRyt2uqrwpCh1NEhZK08jD7
70nIPbGKmziu8SY1EszEA3Q/qu/4Qq0U94D5D1GI/dq31WIqCT45DzKMZxfGxCFS
xlc8KUWNwVj3mA5pCDXDEBvLuBsfANbHM5BW0TbMWRkxLv9DuypSazQ+m73ciQZj
IylZvTW79KV3yC4l2ag4EDoVn34n8qE1r9OshmUjJT8RhkYx0TD29HUNZPw/hr0X
dTtDUHCi2Cpo3eJPQUILh9z81pamSyWt6+bV1pRImAEC6IxTzjpmW7rh4JRFrUAP
p8Zm5CLs9NnmtbnxR2wA2ChZ1z+pvibX0x10k0nssNWHQR/0yXaZ+nc/PvxZJwND
ireEnRz2zlvv4LQyDcErsM5VDmgxt00pLrN4qyR4XumfIw1DHJLmfWCK+LgcGPCA
uI4Xh+TQy0zydfVvOnN3n7ZoqG3nKPhS/sWGJLaJRr8KazEh0XhFY9Ep9j1bGOVT
0PAQSaF5QDdrmBXc311OkNWIUlAb3Z9sGpS/m4XsIC7yi8/g3SWlBjxW1cFkOdw5
rydg2AAVutCiFCjw9XHOZru/Snxz0yHcV5W0w+PSqjDtTne4jmgv41I/ihityL88
C1cA1rl4xxylX+kQuRmicg83ZlaFYaOUTPLLGZDkg4pv1aYtntKYpfiZLzGQtAmW
adFdN110kUkr1YROiewVBD21Kbw9r2GxfNu0pxxhsEvM2CADCoUdFxI/QXjAeccm
6/Fnc/isv2x3uooCzdqBPp4z1eXfVeq1AMO9JBb5fugEiXf5ocm50H4jBxBpWcvf
18bGGV1C5qwmfXhHgmeXzupN6zMJZwPt2EtMfV+JtO1i0xBeBYxt+a12uQGHWg8W
h1KYfaNhWY2xJzBnRd0bmnBvYAAA7FwJGAnvF7CQHrtGozO5sD7D4fpt0l3T8Lai
fhSXnR5gVDhphugfJB5CrCoaGlRAd4ACyUI6Z3U7SLgBafk4oQCNllaDiX7KwsXQ
th8RrAeEpkAhAvmX4WBIY+gKBgDhVgmhxTl2SIM6YoI4heDfYEE7ivN5kzYYNdxT
feyCOpQr7xDk4edGP0Ty8v4WlMsB2GwI9Py1jrvWR7blJBVyoFoYZCqeNQ0e3Bt4
rAG1IQvJwMOrC6RoGdoUGhHYjiykFMfpxv9jZdxqNVKKAVamEhWtLu7m72L7UeAE
FTTxZUvOE44NXXrZBfoagms6jxwGIikZmZvID2CuBl6Afse4poSNqprZooi4uD2o
ATlZOuEEQftFJBO00bEz9shVAmEZXlcWqQihOx2KdyDU+Ce4Wrvh5gaCpcgQt1Mi
BYuBA/pXfb0Gs4uBy/+KRHPYRTuSePSfEapqwAQhnmoOxtjdIEzwiSoDaTuAeLT8
9fQBoOA1qTlIwaVtoy6TZ0Z7WPtgW+jgljJxfPfo3Ep2VLMeAcYd1jKQ0uAWvmUy
egdzi8OEUhgI2wcpkK1gg0Bq2LYQBqtIlMOIkqJsGAl/PjSKfI+5HQOwKZONXS2V
SNgBchGZJ7+/iEQbZWsrWtVbymxSYkTXcUar59tdr2Hnpl0JiZKTy1IIgo4w9Vrv
Ch/k13M9g7Gwr+Q/fJ7PT7YBb6lx6Ho39ps4FQPYhlARRDQP5f9xysUZh+rHTTpN
pGLiC9PypgaxG0EmS38W8UEkQhKLJ9qPrfSkM8u5kWDmxJjt/kZv9BHdle+rb8SS
4Kl/NsppLwGVAxgnL4+nLAhxvHQY+Y70rpt8xq+hQq0vuLevOS6JIVRfMd7iyp7g
bZbY9PnKddWRjbtUfIvQf0iBjXBsi822Zk6LAUkqScbKAjm2jeUHsERX/SwHsqOe
Vx05UOVw5QXzkGsy6bSB4hRrh0aATeE6SlJ9Ah0ux7x45XaoiwCQ+l1Kamowuj5X
7ErCBKcCSTH748VOJfha7tH8y+ANqPVsLfDVnhxb/4u4aSE/DdvYCKegDbzgRls2
+HSiwKxEaAqfwMzzDuQ1dUob1k0MpCsRUhYBcGOsfH6cN/dDThSdo+OyMOFNKb7l
ZGd/gyKJLWMn+GWuBCT+0D0AhtO2iAEyfYhE+KV48SAhYVyv8a48mtX+q+eTkprD
1Rn+1eKAESAXF6yVvEuqLFicuz+pY6i4dL5wu5iHDd1bT1snvzO4fNNXR4tE8DgK
MaQpgMsUKaghcbTdiRsX+17W+n1we3SR6ZUGmUWf7z3qPea/sBntbLf90D7o/SGn
1LoSys619Ux3Iy6kGG2Yp/UBwoY7G+3QmJYY3JopQcSuySfiKB6DRVe+gMXTvgEA
RiPBhKgHJyPeu20xLLl7/ygEmh2f7nE7qPAFVUS+DE+2s/kWX39BWXIdcD2s4NWC
oVwfJU51F1TNZ7nxdy7GTVTg8ACtGvBBDEWdO/QQXzsVqE3pqyLmbHf+Gule6d/a
AdQlYZdbWJcF/UHuDxvLCPjWSPEmb3UW9xBV/YTASzJqlhmCGE4Yyj5cxI5G8IWh
4+ihGFSJ5JNzWXXuZRQtl0s+9s+zWgQme9MSoYy43hYZZsPgmcgIaPy3PbDc2TIK
ISqaoOieBzaqH76zNkAxe9MePZiObA8GzRhTmfqCp6neySBnM4nXDBtvjvyNnjxH
LqogHbxfdSkWzr6bMgPZgtB1KV48b28K5maVuJya4nz/n63kUaNZ/7qKgk9i1KNk
21rkqb+3Ab3mRHIxaLW0uXkcBsV+XGeafmJipIKjOrIegdP3Zzn7RSlKR0CApe2J
Oe081IdUvjv/eg8IM7urqpAbxE1aoRtmxlsoE3YoOOQ1FvDVR7dcop3lwLMKiozv
D97owir9K10hHnCD1sjfZqkq8qxtNTc3dTMq4HjWjC1U3G4HIWVV1tAFLtt1DBZm
M/i/lJGf0EHlCYpZeFh5DpyOEZ6EKrtmMT2m2uRIihvBUrLO0Np3oVDPsQXB8s+P
+OsNmMOmyIWoWYpU/AW5M1syftArDMNnUnPotIm3yltTC8F6zOxPOcRCSfxaG5h1
7VY5sRs3qMiNuRK5ec0ibpz7ArDp7IldXygj2MuEGTgoXk2KfE2ucH03ht98RnAl
4IHFcKlGpyUlTcwYfy2UbIioXR50H1uI6734L6js6iApNOkW7LVGYgaIYGG0h3Qd
yGq9b6FKqgKMVDqAymUuK+Ymks/tyumL8pZmqdydZn6HFcD3pRxyz6uQLZLBejgT
mWVa9jNNS/3UABZ8kr+QPMaXhoSStLxSHH6GEmlDOL0nynmJlYz/36VsmfbSui3o
Y21q6rpKR6MpACMRa7K8SQQv3umdf5MxuGljmhqwaZYIyf31qe1duzMXGbWuT62Q
B3HYNfbQpzZMA+QN3c2Dbd2mRHICKgkIF3gj4//rtPU+OPQmRQN9IDx26wmeKedV
Dn/+YUHVtERR1Rqe4V5G4UMrFUiVvqfjsLB4YiGy57WUQ4Bjvnwsv7s1unQQuqwl
aql7ZsrtNnFoaTc8w0BtFzdh/LeBsUc+a2uzlhXX76B7JfOnjsKihpNjeAzeAgPW
TErCxhpkx7SRUD4Uyn04+E5Fw+dyEabIZHc/9BpZpf5nH0nbv52awp+2qN67SV69
M2AH/ig81IB8uuIzF+bCJsIMzQeaAkDQs/3g/MrDnJpJmD2JFDBLm/kVRf2J649m
WRGOY2qn6cKdWpKP7nqCNzJn+lxleBBX1cqXEvltHOBW4iUXuFxUkJyyZAXoGNXh
x+PnBcXSEdhpG5dmy1bvEdn8OU9AaL57HaYkcZMyXi3t7SHx31Ho+SVZMtI3KbG6
9ZeWn/Zhus/GKxQu1oOb3CEGIg5nVrXSH393QVy0Kb4roctcFlDtX6AGozA5JRSS
QtCAD7HazYYPCgGuEnE0RgBsfg0dtEggtX4seXJvOIQcRog9+TgUkL12CL1/eYy2
YfZrtUwpHxGwFG6mB2FV1lAZoRoYSl34b3KljucHLkqlflAccMYwYa/EzqB2odwQ
SeNhiQ5PxwLfsYZFizRkr+Aj56P4O/JUWWtJE+RS6IGhoSffozrcZiKhc0qbXu/R
bSQNB3xl9NwKM7YR1c7FvogZNNLn2ucDuoT3/IUS0+9rcm++9v2medVcPP6rU42S
Jb+lnvYu4YRV7HYD+DOyyPpQT6roN54BKeXc5UQSSNg//ypho+i7Z+d0h3V7gjn4
1o/0ha6RbHiQQWH0oz4Ad3wXK/e/oLUO6eC8tCLEUmRBobRx7t6Oq+x9P9KnTra1
qJxrFLEhJR0WR8ooDgihxE4HrDdEx2qs8KAVE16tyyRFu3gfFj+X8ZWdE6B6b8K2
oIxf2hKB1x13VZVoMrcWA/kUKhAqssWkC305yliANMnFugSpw3Nsv246kxKmX3CW
HCoqJWbMNjJ6vmV112P+5/H6PV+W1V035lBd4lcflgylseN13sDLt/IsRKrAouWP
Hd/G42+6HHX5qLTdsHc13geXbBLHRK1SuAPCSbwbMqX7RQeTDT5IGlbsbVMSXJLA
XPnQj0K8HumDMKV9Uijg1xWFhLbwg53WMuFCrCX0T5TRQiYM5rCMYdRMtmBdk3AD
FlnCVBP43Inhs7/JZ0DA9lbtkN3jbcbQxSf4+v4tNgd1QV0QDUvSJgq6hvEDRxQJ
Kwox3OgpByMLsDOOUFhk+vn5Qwi7dw1b9mGocdiJxmxzZSv1J5/LDbCMTgjqcPoF
i63EZILzZdRWjt9+/88x0i4IYl0XSyiUWS/t88+yoJFvWbV9L6THp35GR7IGSKQi
RwP3phv6neKbx3URpe4iKccKyOXUQkKth5LyEujqSb8tKOvEZnnJb8+mmGWsAwHq
IvIyKwZOGf35OM8rrbyPSMqCrH98rKJCmcKv+EFxFH36KQhD2MI85FwGyfhtCO9t
aKn6aullsvpJfINSULRt7RcDHl0WrMjoL9rM57Rqmw6yxOfRNUNQmDnTY57uGMaM
EuCJq5Z4JSGxqY1SGxhTqvek7iLfL/GlLjZpFAF5LoZ8vkVWXR0o9EeBLLDuVC8p
YPI3RzWNLuHLgrCU/g1fWSYU/KQP9aIkAHcrt7wDnjrlRJvFE5J9Z2jwiaBaZ7ca
aLCTc5Qi85ug61Zfy/fhalyDYyv6kqvgjlcjFx40mVieasfP8yVJtun3YfelzWnz
N+L0AMxEnFXyHKubc3qQxCKj6XFbtXRkkZu7nc+39cRbu5sbU1FgEWlskAT8tE96
029oxJEJ0qSP2+FTVmGdY8ldNTyY6wLgXIVhDPY3co7qkubTrFLk6R16v+D1Ecob
9ehWWi1cm3kRtuWWuT+6tr4yfTrOTaW9XZtC06nf3wYpMwZdHsLU6N6cKAdDT0aT
p3bQsd+EEzJlLIrPziErkStKmWms9cKbB9QS0RROd7zMo1CIcvurwS09Fma5KMoW
hOKQrM8+MBfJFxwllZkq27xtQngYsdEohPmOzncXzfBlshvhkBdFvsp9YeU+Rq7d
dsezoeWNUQ+SwGFQ1+lQDzOdQTCs4OqvxxfUSz1owm4UjqFBWB0SjRTfne8UTtMK
VkeKGoIePtat1Jt5w4QVH2KRc+HG/7cYe6XFMjRY6MYYNT/kpmQSbVxOAIasUDi+
PUJe3VEza5mGWjqkOUdmCAUREqGnlm0nZLU8JPakuItzZpHFBcG0wJ0qdiu9s98j
7p4UpGpGG0hZ1NYW1oBZleAGB0FfChk0Xa5AGnsA5JOLJOVbHp9YCH87URzCETUO
MrXxYYBzjrWwZDX77scCkrHtxC5/AWi80tkDzf1NPu2IGufe0/khQhiusyu2A2Q2
lCeDQcqFU7NmxOc/GsXRQkVni/oIo3L/bzYUkAc25PexPmP61wA/psaq2VGzKaDV
2VmrRmgce4AGpwTW9UBBPMwarrAtCcKk/Ymt9tJ2bBNvMm01P7LLKK585VJoIs15
hzIK8O4sxhVXKmnjxiuf4v6CvRf7gbF2kMk+sOk/8HFJUeOljbvgpxVyc1NifMjO
+Jx113T4hYmgPnSn9fgU8ks/Q4Pl++J/5bXOwT6EMu/ywehToTVXAiv2+L0iE/6H
ghTyJiqlK61lHC+lyNBln+hcYQvSY7nJib3wOVEEwnAcwZuIISApzUlwc4Zsf3/E
LqpfsguSfcetXRa223wXh78Pa7qk1dmByEW7c7+A6tRzWp9DVxat0kuA+FV1WEZp
MHdqtUFfU7+18H4UPLQwU7hh18/9HAqahoudHl4rW5v4uBjBlZwkptouJMzWHMJd
v6V5nFVR9vRbjRb57sh8ev7+bjut4k9eRnhqOA5JdgNtPsPuk6ZLzOVV2FZ8b51S
0qknn8VuLwh+qVM8KKGgN+JF6A4ENO+KDM2GqHgiYAruR22L53DbDntU63kb1luQ
w2iW+blMSNXqtOs7SVoPu1cqoyYQy8JPymrYIA+QXkCAmFqte1Qt+4jSE6jNQrA3
luypE6CovNK5sPpt0qNkkcgeObsX6keXkvskX66hbbM70ivL1JzhF8kzXJNSxFa+
HeHBVEovbEm0pvGjZOdULrP+HfdFOLFJCVilkBEjFURTdy37spErKTi283DOpQhZ
iQGBKYyRcdZ7tnrQu+eOwLSD+d/qJzgV37gSKmaa5vzrcPr04ZiniLvcL7l3HeI7
jmVcgCKGY0+uIm1FU80fe5RDs4Cu+mxe2pVIUE1i8b9Kc3dok1CCg1+D8hKTXx8/
GFZqs0NbpK2OlgGJfS77PwEiTdc+MGzwiYDz2AnJiBbPKY5zUu8Q6nWiStdo7UkR
ZEH7zht8chi+++gjRIct1YIjXUVy32IfVj+P7Kkcp4IGPbWscUtNIk8rn2kdUOp8
0VnlroVo7KcJ9iUk+mKETGxqIMELZrrFNjcmTn44jlL09N4gq5pOHNboNO2BjIJf
pFGoAALoYvAcJjejIv4c5XWe4PSngjAhocZoY9nOe3AitW6dWP6oZM8Su6rDTObZ
1/MDfHWPVTf0AwbMCA9kpF5+K5lAwo9h+1+9sdQgZcK7KYeI6EMn7L6iE5HEwug2
QhqwYvE+Egh+oAB//C3DAOWd/nqkw8UG0VETPxahMD6K2oA00heFtCZxzUh1hcsT
Sw6P7qOAh542AsNqHBWXeQySFIoEKu4L6NgTkMB+M0VPoIUfW+iqfbv5A9d0Wu0G
+rHvxv3kQWoKxP11kJk3mOV7KXPdnecAR8WemQNf+cqnR6zRXuWxrVZ03w0S6/r2
nZ3y50FZa+LSv+Ipoi3iVvPaxHGVd7f+GH5KJPn/mXqbxwnn4cRUUSJtm/5V1umW
eXEtYVFWb9WK+olPQ0IBrhwY9xhfO4X9i369HZf1f7+kAFkp2BibSDwlnl4WZFAo
lAsWv+1krCwkOvcq0wySqGsyfKo0D8IfwWx41q6CFAse0Es+H62QCYWCsm8dWK+z
kKK3Tmo3FsMm8ibEP3CWosXI8/bYhAs+1MYH/yBRRhx0yyM0qjMKkvFght+MromS
ighlHKH7XLuhbT/sS3AjUio8EtOBxDnRY9FeCZsGav0gulMUfPoEqJXx/Z4wgfWM
ny0lythnIx3D6sz2n1Av//GIsO562vBGzy+SirzgQA1s2GrBMwyOWiWfP+t54ly9
07Ih4E4pAMN3SV58ZWyEvi2l/rNCxQhVZIT/KK8YzaT0240U9aJLkH1XLNlMjSKJ
iCllPhtr7nJxld574H8kp89ifJ7bdMe2LUfNfF93KuMGRKctFn/N3q9t4iM0FqHE
iO/Xu27+mJYEvRnh8JJCnLtLbibGcnD+jhdA43FwMgqLUCZ4X3GRDbsgkFxLfC8n
VPtvCh8Sx+gh3C+dmgPME7ETyTao2x9mnTI+F+oEbInAEbyEkWUeAlxfwY5263r+
nU3fc0npje8b1hslhOPAWpPDhD3IPS3puV7e0qMw9kSoWBLmxZv/jkShjPmJ0QBM
qqi9XhNVqelP/flvqZTQMagSC5J0ASxSXmetbTyPZ7UQMU/YwSEdYa1jzidO8JC7
eIb4ehIkx0P1QXpsoGk+PM65wUxorxJjflcC+r7W9hc69nzivid7nhH02G3RGvvQ
x47hmFNNggaJ6ii97d/nQEOSW6IGRKaq/YrcGg6JBZg6g9wO8eBGONLjA7TUQbV1
rRZxdlWBkOxZ+grHwzwNJ2gdaJdlNJRvNq85Wko7aU4LVekjRonA77svol/5SWUD
ISzIrJG8o1/FJkF2KDaMY3yzjqiJsxLfH79yXjjR6ln0wLzaAZ98Mx9sBON2hJE+
uXGX8dNMyLhslDgvBCnszUV2HagCwO1W5zGi9oiLnd60lf1fO0QD6I4h6uc6JyV8
QQuw6jXQ6mqc6kD9uNmom0AMsYeBtF1Knyea9RPjyR5eOk5JGMM7T4YKtkqGT1fA
52ULhM7XRfeZcVLDcXONCb2srp03gP6xrAS0UZUl6TbeVM22Xx77Bs1pucCRyRWf
w/mTXDE1UbZk40JGBOAADq0LBizwC21XZQvGnvdVgefvKjidih8/T+gUUiNZpjaq
amkeJlP63Xyh/7V6cu2e8M8rs6mcsvTslZK4iv4aw1IdrrLTdobBgILWbDCl1yNw
bPQ5VhFci384V4T7niG6Zt2J28gLCzTitCPzrby+QeOrEvPwNkvEBJdMVNgfy6Rs
28I/o8z91wf5C5NIeyuKdKstJc1EELrl4UTOOAhD5mlXkenOJaztCnWHiwE0NpvP
IGY6fF0hA1ZJ8I731838rci0q+NTBWR50B/IGniNNtkkfiBC2irBz4pHsWa4OQtn
kcFDPnhLWUI6ygwTUx9JMD8lEkj/AK84yVOP22zkAq4rEnBO4pJ/Ncppr4BIiYRJ
HUIBbpKpt5UDJDNyzvY/On6X8cxJBpYSzJM+CDmKJPIU9I9ku64pB1nnLtniCaw1
AbvmE+z8B63uLbvUlH1c6WryomlUuG8CAaCBuYG+O9lTt3USaYkBnbsLN0mkQTlc
8oXbiNsIE3XhX/E61xjEKbmC2UQ3p/mSWNf2JdFkfe+msxhE+Q+MwM4Pol6/px5g
PAUY+rT7Wd4W8qhyo9n2soiBdo4PPRdq9Kf/0ooK67hMvxw2I9YHHl0l5k3z0m3x
ZPLMs3EPQ4+ho/KXfgnhlJlBa6aL/JNUOjVw4WVM4GWjd5EtRk8yA4YjBqsfChTv
DvWbuZbNX8HHtE7VVTZ2+bGqbuxSQsPcix6zb1AMK5dV3hygoMZYhZeLEOZeG8Oh
gBetpO4mfl2L/5Rltwwb5Cnavti4UPhPDtkyaCidcLNAKTogJb8YRltJDFmzo8ly
AyJhqrb+GhXkX6kQCNTTUDlpjWc4773xn2aNWVIbdR0xfsEgKmuo75hPJTGt2a0p
P574KIuZo4rnD2c53aol2QxxfWSm9SBpQ0qgcybNpmN9HqTQ0Jva1A4XqFT7T9gL
gXNz6ze+bymjAukt+CNMIfWDQT7dsaoMqpFtI+s9EpdWRmIg8ViXokaMvqT7pEHs
LO1gAcAoPadKauTQQXsfAKb4odu1g8GLX/7u6zekM+GPStLIywYnvvyGwsTA1FGe
gq3dVJVuIy6RFJ+X8iO8uHQxVoJTNyd+p+AyhQlSVIw0Ng9us4ivLcNvHHW+XQ92
fVBXkpGDhTMl7t4wi9I9ZIJfKXxSRlgT8RBxgHJPmeo88FXcSH0NGXTCf0vJPI7v
LhinRraToe/YVWl0dLLd4ddEjIvWcyUzSZ8hFIid+wRux2fQLD+PIQ4v3Rf2gtD4
rBPrxI9vgTsVXFOBoYAEwTUHkkkpsZf/cnaMGJLlx8eH2qTKGUo9N/4Ox0BIbR45
Elt5Kgm7N1GqwvsEBJwxAFVav1NVXlv6RDjzRatjwGLW7NyOju1lhChy3SrgOEZC
yasYXxvRxGQtCZ0MMTLLXY7ChzyHnGM76MyTiV8FEoe16EmDwo+mVJG6DrB0btWv
rmwCLW1nkGebnJvTVHwlt/eUiuYx0vMCf7tAXMgQ+gKx5+F5Yh7352mcHiWTc+S9
+qhG7yHFCLdXjr7Kq7S1Jiruct5ja67FK7vw3KHep93kB4mKbb5w+fIabaVYuHGY
iEmZhN+56VqVhvnyK6iSrYP0Yv3S3anR+WYKoUF4GPf7dLvM6i5PCaCASf0E+EUH
K3URCdWPllnGG7+RoxAr7Qmk7rzcZ1O0e3n+hGliopJ+6W6XXWOINKgGgkBZz9vz
LQQbGM9c2rRctneo38EPkflV+mlrlIZe8yo01tlJ4mbCb18f6VN3B3KHmPxSy9wY
SsI8ct/zRnLAa/bovUlKQG31qUc+XYVPtQebhvzxC0/cOPQliVw3gHFBDasLLMxP
BZicfNq6gQ1lgUQ4PxWGbtEt+Tg0T6Uu9SxrGyMWePdPszkr8oNSRcBrHxIFEXme
hcJ5kOIv24Sm128A2607/2bvmyj+9Ay7VTG9HesvDMtw5cDdWRPCkkRAL/x+2glX
ZNHlZkp07GAmKeoRF3KybdGNJKjzlbkes/FgL2GTRXQzY4XQHsEnNx4rlPAHLKQx
gnyemmBCXEsbhw06sySFOkD61SCrF5RjssP56PXa0infVowD9bDDi0I2PJpIgpbI
UpmsXaqbGt3zwNRioUCqqG0RvGdP9H59Y46n5UG6BoG1I5mwdn8oq4Bl5nzGymki
YAKnnHtTJreTpLmd7EApijIILc+7qX4f5tA1EvOK5lIN9Y7fvN7nC3Y1KPcZWSKm
MarrMAvk2qZqn/FjOk/KcZFihE4BC1tft5L+Kt/VUcYFpRrDfso7u8mLnPNVq9nP
/xG9Viv46a4qiV84ayAlYuXtkd6oCeoHh8aTUuSqI79M+i6AeRcK4RZLxcKkucau
BCsgzV2M3mSWt+zl+5KUB2jEqkQz671FjK0i/KJJD+x/fpIYcIGyQ8JlhasALx+S
qIBLXp6iSt+uNlJKZjC8cOMV57ubUoPd3av47HI+MA9HDb6ZDXb2ZvuwnUQ96uzq
4f35hHtm3hhSWT93L2u27w1j+bQ5Bg3FlYKyVIEolLusUJuW3Yn6o1Jwzr94OnZQ
Qsm+Fkr6PzHV00CvDCl1yPdUh3OaeQ5f2RHFnwiY3V9sLc2fsfawqqHdkrb3OGXy
KHxgkNLj5otju9CYqRoWgM6QJ7ebTafzCD+XDSsUbeeI1HCqS9cUkHNcOEUNX2Tw
E84PFUse7/S19HhYwQfpmbhDNTIDa1BB0lba2fmWKVFcb+247/XZPZ8L3xyyD3hb
yY4jEwFUwAS0WpC6sP4cfWJPF7DyTvl3UA/Ufm91DsopcmDt6+MqiQvOySGZfRQZ
MvwgoEH7Ge3myK2XIIhIc0JYgEj6lFL+QknKVUs1GCdbvmIOSXB05BTpZKLJmZn7
tF6RUb/FLgaHc5ID2eJA45D27hjUYgJU5+UPkU9XVY+ORSJsGYHHGRGp7JUeHMWy
TJkmXEpo1tOoXYo96yE6qDTwbKJ61m0d2Zf1ccUbxKp24/JAAn6KJKL4ZTnWOR25
7uHzYZBylvdqXAYfXGFWpJbbSSSt+4EgYWb7PuXo5EXc03nD9uOdJV3fPs0qZoFu
fJ9HTwalmVCXyG6VkQgqDL19zw/1LbKAVG3vx/RVo0V+gGbtVKZla94S6h4anfef
FjKNXEnvUF5ZXgVWu0+SxSBl3IJWx7fX1+93D/1oZ6k/RitElfqBGmBKogR7+ttV
9A4d/Ayh4Cn689Spmrh5PQkKiKdoE3OgEkzLGsKtqlI4ALPSSgOvMPYHLUBv96m8
sOJOj8J1OljwCn8Bxf93StpTEBfX+8HO4pjDyRpGtYTqGM1TIAvONw0KB7t1iHIy
1aJqCF5BV5maImYr7eMmmzx5ZtTRcGiwsJm19XdRIzcQxTq+CeE/jRaj+ep2DaEW
iioaaTFHp3YZOKZErnCxXObR+6TAmPC+HMQK50ywwYBAl8JsoLQqRKB1Kd4M5lLg
Pa4NX9eHxIYv9jeMGR2Zb1fAeuZI7euQ7YxVN0706B8NRlBOV8n8bJ19KGJkoNvx
EpUYroYUSdGGFagT9SluF/34clXtPvifvBz3ZDFk1OONusd4Jjq6fIM4BZEj3Bbk
d5VJPcwQ+8wBFRDTWHlVb9Np/Li/FUol0hdlCsUYdpb+Vm3OhGHC0cXOuVxowqVK
WKA3/PICs4DidrtPAF1Q+edRbx6HOnT3BjNzvEH8xUSibvD9FTTaDYXVo3Eia7l+
k1E5fXakuTxDuCajljxqfONWVM0ULMasYurXQqHSuf2MS8yTQ0XfC3OpHec0Y7pA
y2HXKU8hS8xZUL6UnYoTxjnr7EJg8KyCO8UxC1oIrbH9YUDDpY+t9qfYmvz16SMA
txpSRMIv++hNXltAYj+zoXSfdFKcwo2sUyot+zJixjyduSTSMsrgvl/OfIJgva/s
NVlocR/zpbrQkHPPgl3m5WdTVMLL05+PjBpHKTeP/VNOQq2KzkSSl4+a1OyPDVn3
pdQ4HTrjqyw5ITmfV4tXWC8yaRZ00Msxhs4/X6tdQFcIMZoO/22Ovef2MOGIhpr+
mUFjpib4p9KvrEEUhCMGZRLZ1qfOQ/1FrirdsZeT/M3J2LMSyhszeA5+IB0TIaEr
ig8N1Rzg6BtRnMn7RaXVL7Pa4VAd5jSVkOkcG4rRpHt66vtF+EMXCJ84Vitidid3
VdjbE1bUpVelnBCACx11ta1Q9t0CpjoocnC5akW2DyC3ZHRPZl4lLe11Fsq2rXTb
KyLgrDZZizUamKXprI11VBQWA1P+VcP3DeupySIFvETmAGfyf01gL6o9AzQoksGW
Ju4ldGjWmGUf9ILfSkJzmk5/UAHJfHvz0k1/giJeFh8c68DWQySWlHPNOCJCx2ur
FtUc2dbXWE8+VIKJ01Gm28P/qbsk7vgJL+/t+eem6YxFDbC/G/WNLR54x+keFQsH
B2knOYXdH1HrBKM7SC39+G9YA+mhdTTwGoczOpLDWgcnl7h2H88C0///g4R6FDky
Hra7Kre8dV6sXIvO9jZ9RdDWpjl6DxQvK5Yo6KPLJmu/rMZpDJtuVeVNkUzqo0p/
p3SPBP44jIEeUa8Z7YrL8O4R5JwIR6MekHQ6a8czJ2eBQ8PbAGwmf9aK1cb6tVIG
qKMHLziTbAdBgshJJjaEylDirh+8UHyWGbApCcurJqIcrbvyIUyMAoQEYjduCa0f
25tJkQA4X6cqmCVt0cKMhdRn4z/9qBgD5/eGSsyG5Pi6l0xrEsRcZSIz6OG96BSU
JBsk7LAnGVKmzV0ZchcbC0lFMBAE4iM0ooGqLiNw+gkaDJLC5728kVCiHEXyX0E3
ViGv/LP87bA83cOlwzdT8gD1D3mUBuD33Cb9V173ChHd7W2b37wYdPNbDWUJhTJf
Lbsb4AExPa9jFAC0DZJ9ngNiWtF2Nt056OKxPlWQ3HYLTt0tMQ90In1iNRGYk0J/
CjbcFwmrFprWvFJ6fAai7GixWA7DWsrYBdD3xm2pRtmL8UNSG2+VhzMVyTM+iVvc
K1w7XLne3iCAI8V8ngsXDK2FlDl785MbVDG8Ww834BZikHvMhfxK9CcMtyXKN1wr
ml+3sH4WhEK2KkKPLFnU4yqLBiUi26lBtXoAyxaWRI3Kz93LLyze0Bhuc+oq5B8W
Uds5/QvVvVh/IXaB9B6dO27BqR2nSFpHWQfMxkqQgV51GXmdie+v+uCucH0V3CCa
cPnfxHbLaINPbH43i9PcWqTeX7kezaNZmR5/9aeUB0hwVjcm7dsyPjdWafd6W5S4
Q7bIOHLCLSBR0unhJCxWSH/8xqVsL5XnSTH/ty13ZsF5cu3tVQlcyfZsgBW2w+SH
GLYzNqJbaWjD2cetrWVSkIHseYiQFpUMKB9LZ4biC2DF+b7fwmVo+WVCSMc98Nx8
x8owlgn8ZO5Fxy0mXsAG0q6aW1fO1s1VsbOXsqgnTlNna4aXoXt1jBKfmDVnXXZK
u8ZSd2sVXLazoPJQePFCxXcJk3httqOFvp03ka0wcg4IABuqfID/m23ENV3C8nHD
jMNewdPnEMSH3prHMVWUjlfOOYEwBV9HUjkMa3BI7JlaUteOILHE5EFLQERiVVJd
xTHkImsMJ3cQTHNpA0yBoiUmVGAoYT0pQkTtQWf/iujxRrW1Q2LOcH+nac87Qhah
Fo3ACJtJzDmg7r93YZ2Mf6GlyfsdaFqRmH6bxk0ruXG4v26cii9ao/CYcwqh5YxE
rgyOavG4WVHf7MakH3D1TzDnC06r71RF2r4rwpbs+TGu02IjF9LL6Kpvib3RLmlS
7AnT6Hgsp4zucMbLSSjzy57Z1EsCTnPFxF5JD19eUAulMw4ZfNCFtGVaJfR6qCPD
M2R/ec2iwgzHDv2KRDqTHfpVKTRm09Q8rhD9hut+j5C1DeOjuho9X01ZTA/NvFsx
0KVCsRaKL+SmalgvkCLdAeUQAAeqzKSFdRDswwcwNuAoxbekilbAe8oL8SSI0tuK
SgqWmBTqcuVyJj6hQukdHqaZ6/uEXggyHndUQ82f9vrizvjR6SyIHGD1NFsBvWAM
XKaCh2hAoEL7LN8sL7IiY9Uw6WyYZ7z2yT9t/OLZk+t/UYtkzfVjR9hVmu4eM1DO
Kbuq6jc51zza831xfXOb6p7gcVPfNz+duPr9i5WW3fmdbzFSuXdO51xq4vvn543J
oJzxfQ0MJ2OpnPQkmKgdqasUkuQhQvdEF7mjM1PdQLSgvDtBIqP3alOc8kWBlmo9
CuVBg+O5qI9zP5em8Rc3/CFUai2mUZgf6TIaKWj/ijQRo8Fflngs6u8OgqnwNJGy
6T0x5SdKKG/ODkyELq/eQoukrv1baiPz1/4kb+mHWH1db2I2g2Kw8EVvi6cY7FpE
4S+z3iVqSXbUGEAFkQM5IEdro+0gUuEHe6r8ATAj7IZle3/gbcYgQgGpiZUH2m+X
towTdev1nkPORTWdhgzRZuHnIotv555WAJpdd/zI5FvJ4lnWeO0Da5BuZWZHJFXm
LxN3nkriOAp2g7SzxptIDrIQjh+LU2b7pL3vdWPKCE7+1Et4hKTaVIe95/Iwtnvh
4p4bVBlLRJhwG2i0G/3RBVA4tvSzr5bdlKO8wJhycXljwH93NX2sFThrkmduzMew
zjCIvNCuJhLnJ7HjZNZNV0nU99jgk97bjw3cRR2kKwQITxWShNhNTt+VptvtWIlI
iB9wNYFn8liWUX6UU2Xf4GZkA49944rvLiOf9RysHBU2STEgCZW1OEBFJwo+g913
T+G3q7LrMORe5cxawKOedVC2QqqP8t7EsoG3/dp2Hv86L/ieM7BiFnmfDfBAJ1rA
Vw5+xEilhUSNvTTCDumK1fhUNNA03H8IkWsF1XpTb4+t9gcxaP+pEf5PIDFSkLFm
EuhOBLAXx6jADuP/woCNNhj+cF5Fgwv87Gc4FtCZpet6iMgz4kzi/JSh/69DUEsu
9zk4C6s+eFTV9lVdkPDxkbmMGjzE39wFYwbmxTuNFh5NjhVYaNIzHzHBtAdkjIHy
KA74BZHQX4RfwU5gAdNu71icy8LIYVl2AxIk4R2ao+60jxnq2zvzpaJ+xJmgWAQ9
BnT0loGAz6aCtHWg8QW/SRwe4/eNF90sXpvQrCAGw+PyKEhXuLCnnezeSZ44SXtn
JX0wcSVMGmqDQ/4FWIAUOLsJelXQVl1cxBwQoaZ0/8Off4HjlJlHJwgrn/DE9dmR
25xMPrfsdbxXc3rnXxm0z6ni0+Hfa1HnxFsMQ9AwslsZLgYkkvJBsw83IhlzCQDT
nNBuunhynENChAMW/47cVLoAA52f7sLnOs5Y1EYDAlqXvInzOT0sUB4ob1hLGiQ1
UAlL/K1b87VunWjQFmOge6b3nYmxxyflTs9p0C4vhnPJRFWXnmSyDbcV/OqDGaWp
v+HzrMScTmGWBqzPVk3KNWeUztKEx1HB9nH0ntS4sGjgRvn4PotJE6d0mi+oJ6v0
s+WKa79R7dOf4DSX67kFh3Atj1J18gVmEqMtG+c7Bwy8kB+FvU7DjL3yV5c8kqo8
hNsURzhsR2w3qyWHsd5NJ048aDUmuaomCAyyFsYxhvJRY+Y0nx9jJTH77y6piGWX
gfjhXaE+FzoLtsoo0/QMomtaciJtAJWGrDKSOfAOHV81ivUuAqQx+tisKfsFhh7e
B5Zl6Kua07PhUcUSUA/CZVA8zmSP7Y4nsqZU2pyQV1Y/pdl4D2M80iOf3qKSyGgl
dZ9t7WlsyQgtx8OG1AhN1K1Sriu56qrET34oAFAFNlasgdzD8KiWK3ykSX6yqbmC
ej6s9fRXf9J08MntcVFzfv2GUEaLC7mKoRG8GiusfJp04Dvb0gZdecQ5Oo6wGqAq
siXSVMTWjYJnyCf9INJalgtMTrJTlv+fER3Bh+2AlyKBh5lJs2VZsp/49NvagWAY
MijIV90jGHqfbAEYLISf02eUHcKSoUxkNFLAqz3HzPfQ6eKCP4K4cuDHzyfsUuEU
etgYsfj32fwdZHUm39bj9ZOz12vOL8BKihn/8hZOncXqo+AgAWBO40wkUZDLNsfx
dm+NJn4WLpngxxR8rC7VjLmCvCk0mHS2EvuN0ZHYjvouPpLjBukQ+feR6lRD9GH8
3veRoQ1g0kDl9cYCryTLj88H2c5G+D3cCItKB5c/q7hvzqcez+LeFGiFQqZw7zwF
t3r4D0i+12AiYVvvV8woE6o/54ARQ2FdOilDN4TTH0tQ2jEQRgJvOQd/pTUllXuw
t72wWI9tCGnSeDLtVXD6myyLy7FfVnZKevSweUV6DU3VDpRm5Bahnt5pFbYDUjtN
6tWaws9yI3iqwgTcniEDbEyPL0u64d4kiHFYnh51q/PI3LCOpbGglqYzAwtHZMXc
mLmG3IF1KOEmQ9W/ir6lxRwKAEjJvJoNE7l+uZWhBABx3MBKLaBp57xP3br8hWm3
RqDff2G7B05VpX7Rs8Ka+y/fSQcxZvLPgvj3dCPd1c3d4YU/5Tlp14xTGq5chRLG
KIPE58GRULu6itPKUJoLDbPx08eHvP3NRD+L5+9T2m6AQu+JJlBJ9D40+mgetWmU
83AFgFCD23f/7NawoI/Y/JJL6mSq3XsJN19ShkMmUW0LTrCGxezYJvL0vKe1uEW5
61PoK9edN6yIbtjYHZhIrGi7pRNCIGwIa+shPomGDfdeDL0x+Sat5UESX0tNZCQQ
PKohWxGJWBIghA5lS35ApSciFB3lwug58P7HQZH0DduLw1Bh7rk1k7a595ksJQYi
Rim1WuK0VzWUlSJpOrsQq+wd3WxjGxfYcTX2XYvowtDFxeCISrJW8ouNKW19lSS8
aKsWGRZV1bwmATkM4FmdFD5sIggGQxmnD5v9n5elSuA54n1JhZSfY2b08dWp1FZl
T2DE1YSCJFoyCv6wjXhw/ZOnCJ2lkroaEASLGBqYvRpYcFMbeLiQU42u5jevI8cX
nZ5BAtvYsH/lUz+07Dwz4Z9NOzEX72YCVWq+4qODNBwF+3O7yj8bofiIBmeLN8Ye
D1plK0gEufrl+eBGGIl5mfWpMkT3xexB2TNDIekEdbSBfIxRU77dL6P7Lvw5Ai7b
M1ddM1PxSQKxBmvP36w9/DKcBht6go5GJfiKNFUr8VHC7FPhAMsOpECrGqkOhHUD
xTdn17f/2EmSbkaDHS6zqKW2g+eR6p51eF8SoRf2KqzZ+JQjCO+e13IICmVEq7gR
0skz+QQ1ZudELel3wN5gWso3bImkFTzj43OfX0aBCLTsTCCY0arD2cfb5lSHUzwK
ybFZX2U/83nf+BhR3A3HiX+oCovvplpb8pcE0Ssc7FxLRqEu80VaWprYEMCbFmZa
9qNHD+dmPyXdlq98fKmcIqf+RJYy0IrQ9jY0Faz82vRE/qFHEu0oPK6l+emkNFvE
DNeukWJJlf+8mkmL7q1jdLPr0Vl28enu2AlqfvTt9PoPMk1A+6eLYKVNWiepGxvI
lbNVzfMbZpJjBeR3tUgsCavWW9oeZjE1KNiqa40dQUPgd8pFCqNaB3DDJOG5tbXh
1OB/frjypqSpWoETr2mmTrGtLCTAo5t3QDq361eU49oDDKcH4hhZSEkOaBqPg2tC
kTrnRP4b+ZaJKjQZsW6MKKbiFFq7yU7djMwIUBzbEvnEIEUCytpBfYUh+IP3j8cn
BkTv7B/84wNAGW0pXBlRP5xb8sKQ+PTS9AvGZwpTePiaWvKDD348YsHdnPgrmHZG
5XxVlLukjEujwuPIaUoifUNA0CfOGkydiAMk2O3i8rjpZZ55pLPTP6g63iNqEHu0
5q75PidnE+2FpwQ/lHcfruE+w95Ko3X4Gl3XHztDV/+8j8ZbJoVtsgnyibbT8g8W
38q/iDC7vVoaCVJ1P05D8KsO6KHUbXKjtmi12kWd6M2BAITMYdkwTZjJtihMc0WS
KXs+DeKiHn2I3VHdTzdxzLsLILUkdSapNCuZWK2Ie4g+ybgYde3EQBUs22945Dmy
JJfbg6DebfMZ5pyMOckCuh4lSGBRm+UTohIp1tIAVfXGa/8ZoWFIUWmtSG6d+O92
INDMak6LwxaSNLIhYWxgbcZzq+UAwWfw4xGUEJM+2YzYrM5eGc6fPg4Q6rG4ZRhW
zrfzSvs5VKNdjM4k7ZWW/am8ipF/cw3MVO4ANHgjBf2QmqPHIIIxg4DCuI1IWZCo
acl7H5xTyd2RmBuxHMVBxz5GndRIfHAIEtyz6OQCRyWEuf5Su1dElxTmt85Smcs5
zRgxy564JtslfyJQkX/9I1JM0qlhkdQpvLngXeH/JN/Mprw6TEJv1JdbRm1A/Imm
nj9FuVp3U2qidDB0+vHLRSL3Fl2uUYrMGaEpmxYUq916T49ZYODtS/mQiyBauiLb
jswDyxuZnTw41TEF75VcYi80rsRUO7t9rLH5/DQYrJs+DD+/ZaH5he2OUV8fNwF7
A/hcx+ONWgm37QJHVKxpL+T9Ngp9WbUNRT750nIqyDHUbt1LD8qqsPmTjXIIOmm2
CsqHB1WwnfbRAhkL9RODQo5VPekAlh5YNJSpZKnR2jTzZkp6R4pJP/508O1nEApw
ZdZS9Nak4lXXxoQ1l8YIl+akhUwTcAJ9HneYl7CsxFKm4x+yL4Uj1+dnit1GyUBd
Aw4xfVmebEinKveQylt6bzec5X9+LrIPaU1cb4aRaRDcOgz+bZttaO37R0nOncy1
RbRWEexwldMBdSA17GOAi8GfIyOsPbjcVOI3RrOjahfpFaOrvh/NBdImYOTrXOEr
nPBMB5t8M5fLzl1n86OL4PC0NhDwvbyD/5bmxeBVRjQX3+k+ptvZBsHmvA4VtFNh
VX9VEctvk1AhYEcL2SJYCTL3yQ3uZT7dL2dY+0r5k77KJFv8XW4mbrQZmhrL7sMq
5b7y0AuRop66LKE952/mNcezB3wy/sVZrhzqCYAeuE90hOdNam3+tlMNknD7qJcq
HzgkH7+v+j38SOdv6R+Xyp9+7ddfhlPzVj5wau8KZwOWnHJMrZW9ugyl9JbL2F63
ZmP99EU0h8Xliq2EQdMdFpdyzqpDY2ustJCQVMzQx9V2EaHNuCKjlAP0TxvJQ9eR
c0gP/k8BEqR73uKZHHhzH8fvpjZOxXkpITXAE80PoJWLJy8DwZ3jrn+ZrqxzISD7
HNwkh28AbfQReVJesFbvdCT1Nwh0mVS+IdJMvNx81m4HaB9VU1eOqfSfBAJk8gqO
cO8zAxrulJtdcduNTDaCOf5NE7+VG6OvAbUeYXJYfzVKPNRPi4dVbkqgPW4NMYt8
SScdScsP9qpEgTizsHirgfihEe5+ak3M09MXHMtAjyV/qKE0MAhUUS36qh7/kCNP
iAXMZm8qb0rVuulp9o2VhhKqvp3a3k+md4rDBRoKLxk2xfz6UlA+3uFoN4EIhFlE
tvwPj1CnNwMuiXA0mLufaHUvmcqaVtOz3zmHt1EOsv0WtsG4OxFU2D9HTePQmSph
JVyteCe3BojTO7/OZPrwQEn7wK8qKTpW3KSIul33MfldX3glVaEfMpDBFaPwmohd
0Dunb4+lVWuM7boeJSrQPqxRJQOTyqnv9OHCJfyCu9YNqsONEJXDDWWEJs3IH8QA
Qb5RLP4uFQED6Q8X2egcMaVK2qWhpS6Q6BUKM3N7rJxM6swN5QNSvyzdqxuZmIp1
z8fjx6Xop9lLs2ya4Y82ePfNJcbaY0molfHTXeuBKqRLA8iiJIEGl59v4QhOVgtr
+AehxbIEco/lsFlWw6JkgnsuqBaRVNzHIPHiss4BNpsP2GSnuPEgd0tVrfN8HILW
K9laQScx3w69O3jn1uMGK84bVeEPMXnyq8Rj7dcQeJYw5lZK6vhFZmWZPmdfi4M7
Uw+uCY9ylXSo4SG1tzCR88CW3eXCG9qIoGEskIARJkgBHaAVKUDVzRDbP1dnpY0o
NO6Zlucleixm9ZaNcLQAps1cRU8o8UalubiCZ45FJUAfWxsjWglrYXd4RJSBw1V/
DS7bgv92tsQrE+vhiRtRo8/v9hptGuoqct37VoT4kidcYPZJ1mT6S9atyAGbPHZI
QuhEGxPy9xZjEYvaM7ynmE61FCrE294+9fUzD/Ludm704gi7uinDFMPj2weSvF3S
Z6arCKGwbBxY0tjskP3Z3wLtI5Ihfj+Ovwz1MVnXpXYADonfnQin/CQSVYfEVfi2
nLNZrlSiCeb4KADdA+BtBXKHDXcOrVG9Fo7Tx4GuraGQcBCEjrHLO/ESAiZSCtBf
5QXFb6C9Sazm35DZA4imb8xf4fJ4+XwVrFeqB084hIqYiKpM/mTKeaciGA59V5z5
wM9qMzm7gmIqjvJZWeUIZiWVzqzMGud2IXLzXXlAdehR+x1Ercqt+JYnsKGQ7gvh
qklfPXM9DFNF77kAzNtKiRc0DYiUOFvDrqy4leSFGhpWRmW79vR+0ASlRbmGCAX9
qA1IXKvIz9t49k8yBJxgZd6fZw+gZNFee2IAuWahmjT8qg/Q5B+UuoOSNLy2/A9T
5G8Pyw5SF5vHtsEW9tL66LAAhrSq9KwqFrb1gyqaBDhSzgVmkZsoj0kNfP2Upz65
kGIUMgHLyDRfNQfSu7hMXnL+cTbnLt7mEjdf8Sg1ts1xnN6Lp+6As2OfoYu2n6sm
YOphaXAAUqkVxFylWaM5BJwRvjwOjjxokGfW/3qWM+W9j7stEre6o00PWg7AfZ8q
Pbam/HymtJ9zBxG4PULDazvEPiS8xRW4Ug6y9XPDAv0pnKebHwbFrUqxdCKp/BqH
/+wFg2ZdigSyqs+dP1+ieGVGZlQOjgc1Ih263eGK/39nbDGvNQ/FI5zLa4Gt4xVV
t1h5ImaxuND2mZf3AaZ+xoGSgwcjm02IA26jC5Z6qTV8Nrrf7sG4gREAkb+XW8h7
kmgOUic9HCw5ywpVAB9tZ1wU7j/8XRcv48XiFXWQMHaR7MXN2cE+vxk5EXYm0sQb
pUiZTo2P79iK3AfeRvsFJT/UjpkRIetMe+PnxWRSoTCcEsER6hpK4n0fIXaOmY7E
ByyMqU4fY5xGi28tawfOpCBc2Ky+2+mZFdHrrNk3Y2gfQSHlIzVbtfOgn7+9x8L6
duCVVKol/2RrGjfxrsO36Rwyd9bZ0xK5vgOcmCTKxFy7u4qm/i+GW+bsO1RT4di9
xXjFiSycC9M+L+rIX+9Y5QnsaKqMy5+HoKcp5Dg1Ap6hULuXt2+0pdC3eQCM6/Zw
UDVPWYQjy7Pk6lZmGPdNao29owmFMsswaWcxT1x8IQu8whoRboliZrfPuuekZr8J
QM3+Zpd87AhuY3gGSwBy62Y9bkldgfDhCLZH2ofA4aPvKOr3hgJeWikPRZiS9dCs
IoAptmlb7lGV24Fj6eNzffwunZ+MMF4SEPIx03V03fK5xltNywE/oJcWkRM5AuEa
NUt2cyGZvTJUeswlGdRYOke/+1bpNN7fSZNtlz/L0oQiiDo6QxayYGLJhGw8Ysqw
+qcOV7Rx763oIOypsJIvx/gOaKLGe37STnWmFnYtfPfMmZJJ+Iz0sPjFuET/XUkL
IUe7sjCavcouxEZlTgexCCfC5IUxipWW5mKGMqc/4o75QcCRqwX9n5E6ZCWEDe+w
lXYXFyJaJkcmhjYHm84mluclGu7Ra2D934PpvJkcJslOcz9shU6rLsAovWXUE3Dv
UpYFaCd4f2SPsHGFwk7Row3UHsryBMfI/1ZR7O0b6Bywk7psJajKspBtiORqqBNS
HxPgiO3EBpxG//iRk/qh/f1edQYfgpqNwUQOhb1vnxxn8HD85jjyIIfzaO8OimC/
ovmcWlQ2n24mHz0b1SpDtQQIEeF5YTkpyGHWYeY0DyjBLre/PzEcMKHWuVPPveMi
2X6F8vekei1ChfHUMo6O9rIMgQUzZQ0hWjFsa3u2+IscpsAEjysBapVrkwuNL5cq
4gNfAXqXSwRdbwn0RAI/0gpr/5kBtl/U029HNgWDvrlGysDRewhgHQgCWQC4ay6Y
cj19BmCvhGHtiWdQNKh5fxsNQ7Y8IIz0F/iu3O5TPY9sXFhCfmTJLaB9b30lGpkb
a1XxdZeDd+J67mFcGtYuWsi2CbzXD8cewIvmxzhcwnj/NJYr59HNCQ/b3WLKpn4d
3VpH6u/+QOAcbLKez+/tdG9cKYIxyge1PYdDB+/ZmezGgi8mxPBb6n+42gDFRgHf
kHoUNBUSczxX2Eyz/hssegCBlgufFKdyVDNf8PfNhqHKgMMnhSQkiNM5y4l67cRl
P+OJGu7EBBfIBft061XjszocdwPEsvfHP9BI6tPmSEzHPRka8Eh7Goqj7zxP6Um0
qFilqcJNlns7yYR4tg2jEGLFwv9tYX1jjdHMMhyUq92rx4rC4dHgITqGH6J5qXAx
KCWITk46Ty4uniE6gDGX8Qqx8FjNHSdZfd7y2AILHvrBTia/QaoGsNr8xzz47Y6O
gtbbpKqrgOACSybMytS6Xy1xP0jqoeeuvJnuFBpEeuutLz+yFyXbOoO2Sf9ftafu
DdciDHom6trSvm2BDAdBgF0UU0QIWfP2/UEiZkZ4eihTmW2QG+NLYfjR82mYgupQ
RKSLX1WZJsdEU2f1ZsUcktUcbh8eGNqkd7B+e72wW/a1t68yFdMqNwezYwhZg8bb
b7wtbl546R+rSdcOAV+8gLW0TYvSqUuqacdJELRijPtNes1hpmOnhzfgKNjDz4SE
+W7mPvGR2g0J0k90P7uONK9rAUg5YsSfG/9WrTv2o8qqs4d6m6BMaQGTgoW47I+i
kF65TJ0g8EEodIGR+s2vRBSENMq1L0qtMf30yuZ7DtDcd5Pf6Snf/Bf5kTI/fpZp
W+HX9TK7gBFy9yLHT4sUK+WKUCjmPI6Pp9C8RPiR4UgDE4K9aLyDuIdJG9z6QzhD
h7VAwI0cXBj7ILuKSfwNAyRpsi9Gtx08aNpfePO+ioUXsSS0XFb/uYN7lGCfxy/F
y2hcpXTTYMnztZkQ+vreUUGWOVpHpHOBDbpUMMRLA0ENkvhU0c/xt6hoFO2faTod
yenDvpj6Prf6+r4Sh63b4CtY1dSpfhO4Jb09NqZC8jX/UcTozF2N1M7QdBhQ9qC5
A7jAtiLMz3kH5jhx+xlOydb6/n+RJ+3Qf0V28xmyTfmuaFDS8voF5IvE2Vr108em
0ZuLS3PRc49FikAEl+MgrRGEMxcCx7G8yKfnMxthtEGB5qdVdoLFZ7s4xYU9nNeo
s5P9fHPezZaNGJ6ZKQ4jiyS4kylrXmOfNxEm0Epog7cg/9qLI4WIiWfjkwsm+GpV
6TjbTXOMihh7NdTgzNdaVwj7NboUCmbRyKyaFJ0GsqBVwtntC+F98fMj4XdHqaHt
6ldtbGGJt/XGCXUDhY7V8FqUS3Ms0Nz7g9nXYhjjWwDJHe9alonO/OFzHuLHFKY6
iXCbgGo/V6xobXrpwcANb7Cz6/7AycNLf/W9N2qqDxdLlju9boRXtbbw7NQIUKbf
DYaXAop1wt2M25Fe5OgIZby9aL8XOo3wn3SPWQCgzz9Lfmp/Dz9Pnr9UWr3PQc4U
XEnvBFwerL+FjtoRBVm51LDBrBoOhozgtO9Oa8531tFAMqdaaXDC2TF5vX/eg4sd
r/smWZ+fkdCt0kiS0FnmL+MKMsmF/8MMsSjXeIC3d77i4HCqKneXK+xEmc2faTW/
sf2AQIn24xb8/14urjFp/v4s3/mCERG5rLrMsRvQ6FJJi6t50IE0IqRjsBRx2cup
HGb3c7CLJay45k3iUWRxJrOeNF05u767F0+CLvtDzXxtO/QTWCwenujRh7wMWWKN
FRy7pLrYAMRaDJUAWlWupQopg3R5DV9b6486eOHp3zY6esJJmk6D2sjQ8WAwN0A5
OR1c0bO5JWn6gMg7ujAKqa3R0+FIsZG0E5UZhnBLKntmA+8ZrwJB5iPEVldo76ly
2DP9F+GwnBCvD/HpGlKcl7zbC+nYIakiGCA7R46v5nZqKubP8DYSyD+qDo3YS6wE
J5UdSuGZR9Djxt7HZBE2jqPpSO0kKmfJHGyB5Ok0UkmkIYt2lMVlq9YjDXsKUbgW
5K9NsB1QJMk27P/OgxKgP0dzz9v8uH92yxzy6sCq5S9ylwlC7msvZLtB175Pt7BV
XalDC7xmCC8jGoNxHGnz9QLGpFJiQtQqWnHnuFrE4D5g7fkR0X05/OITulQ4O9Ii
Vh0Bls08/kgnz8Y2FCZZTh65Q4kS4T43iJYrE19iPLvPatLbI/htKuaujUn0YTim
0iYhZ1jsi5KItVqGO3EzVI8dEFGcr5V1eqaZN9HtIQuTGUiq9LjvBNQSQrms3M4k
CWf1gGlT4wmN2rRIy53e88Xsdo437XwTV7OHi8rgHZerITN9LFhsDbugCgLyKtHc
YDrFluZNC0ki/aCMnDM/IyHzG7DiEDChbP+6kncM+vZihTwa/X9mUbn509DE2SOB
QSPJc07glLTfkFpzoXxIcVEvWcnVbOhymHsEhQ8tIYll9mPeQDCl+j0iRS0qt8nl
ZQberi+/Gv/GvGO/Be1ftLGqo2B76z/yGJNSgM+I6y9vNrLzbBmbYCUR9aBB48uT
E573vadM17jEj2SlZ65O/xeA4suf+OTehu3LlM59DfcGY/M9FrVm9TH8G1cKWRpF
GSLmovHyuHZP/zJSeKZwgC+QdDN9iNPuLdX5HqD7H6ot15mnLqHKSm+hkLuHJ/ka
4Dbm3OAV1ii7UhuaZBK7n5qmlc8g2GDdKuL1Cm9ha4ZqaQh1cb/ZpN69LyFhYI+S
q6XUgB+UA76tofmk6Q9vbVJHTdg4bH5hqXyE70AQ6VeDuqZk95VhqmzuLguF28lo
MQ0wOqc1bNFTpFkRuFJWGdWXBFhow8w1Busn5SYNySmE55UCWR1S+x+SoumSn5vP
AcJFu+ELVhMBiz2D0gPTs+IxCSdRVdE8JoeE4IZDq4d5XaQ/Dx/E1AuHIjYTbCT9
J3+7lnMjXMYkbaS9hjO/A9K3hkNzSLLYzF2fSv/+V8/B3U1BF58KzbMSfQ1EHtTb
HY4WmOnzJOx0InGOZkoWGgYBqLPUrYdT9apWDW0qQSxAlDM4lhmqkFj8zyB4zNRP
cXfn6VvPMpDamtbw97ZuWIzZBTsW7c3hmsqsdemoA94dc+odU7Ai0IPfCANoNeHI
mvnHO3/VUZMTL/6zBGqE5oHP+pkrmEHOsJOhv9RaXdwgKGzvk0kAbThlr+Q3caGJ
N/D7HHjHb5PGj12e5n2qACp9UnNiaNkmM6avUXMVNjsza2HYbgJm88IhduPD4i0W
YOEwfuoNQa2AJo3yXcfbfmr203OoZdhyYP8b+Sul1c5i0F+dtQeDoPR3f0n3N8yq
jKv9oHDqVae96i43luDPS6kCGNDY65HmHm5CJVGg42Ap31waXeqeKpOmXNaVWmhv
BfIdmJgBCtMmxaTD/p8RsynCRl119IIcW7q5SsKdykxWT3bJ7dXy3S9f/4HPSoNY
lLOqJ9+s6B9XcCdcSBqj5FAfY4H1e2T/YkbCWtsIii9JesCxEm0WbqGj36DbBdZU
iZgIF/D4Gjj3lKG6D5c4fG1JAsk+SH1Y4n2ijC1ub7wO3eiWQgd4pRx0EimNz96n
P04nkZuBjemrKZXottluRzI6NmIFmIxY7nvCxBdrnc27OM7vaZ7wLQQiwbuL99XB
ABzgCbsQv121yP1ctOqbAoSwL/tclqrtiGrxuI9P1Ppi+Hfh2oX6zoHHpP9aTHoX
c/oZvanzZdz790MyV1WN6coslKF6I2VzKPdYkUaUR2HM5XygX04Du6PNt7VzKCTe
H4kOYKWbB/pUZpcFHtE+5K1zsz00Ji7zL+VIAxT4HIyexrsXL58wdAKA2gwUjXL3
HDyhUxHQtZpeLWWAgCSDRHsu+0HZUAJjRFkL8sbFLaQqWBTpzT3D01Jq+N+iVCl+
KtKRQ1Hobpjd0e7sov4wJu115Gl2ZHQ/URwYqYjWC0CxMfb5Zw8qCqOrBPsMgCfU
FTiD1xrUBvG6rd+/AZXcuFmF77KiDvfy/5QQHnHU1JCIRQOSm2zoIhX69TLykos+
muT7ip+kWFF53pJaG4ez91Fhe5kwWRyz314PHz4jtcInYmI+PT2Zg86DMK5p95vA
YK0zmsArfTpmTZDdqfj8+dISZB5PzS5exeFEcR0MO7CHFlD+Hpw238tFjRekH6aC
IINO8NhMJ8SRQtwI4FzFuay1rh+QQ/LzmsAW0o6Z+by8H2l8zc9GMlddM+yyaeTr
SfumbixbItu0crPw2YD/2rM+TbUm/F5vN7bzlTs/xx7eSMPba8HbPBwXvE78W1S7
cakzTRWqNcfC0CUQyYHgwMWHc5ESzYKvfdCREQSe3VbKEO3/h+tioOSh47ZzDToU
csDpr1SROKSfFEqgGQRQsMWIBfBwTfD/fdwrkpzA+Rw7GGRpVLU+64Zx1nrHS+VX
iPyja804C8ZO+Wj3gCvmOpEsRAar1t/adPbUXlfyik2RApXyuVK1sx0Uj4DIhmKJ
bzn7WHwEXLUATmjmzbiJ+DIokRggU6kGJTPXtfDhcTyRDMtkKuDi1W/gNclMFePX
69uK3OdFwBgUvQEmFnWkcFLpjmJIUCZSuFzrmXQz2qlihtc04Hg/48v6bv3uIQgd
8miFSyYFtTCnzOdnOHahnNTZ67Etzmtg5b1+2ra+w4NP//2YXb+JWqKKuemp6juV
G7xmImF9dEQ9gIRHxuids8Wf6UYYBORWfL3eg0QtMgblo3WHp9//mMkn7tbksu+u
OhbtNoXgQ4tauBaDzdz+VbN7kgMS/1/IGNvdZFx8NKRixCSk2wBLW6xIR/EFT2ba
nhlrVvML6xVahfmqMK8zE7xUOCFDlFuE96i3laQ+oxcyVHvMkpt5Z+R/UYFSFAlA
4dRGoWNRQ6GLl5Npv2K4enVWaQnpceUE/Ksmw32E0r5d4GrHqcUwMihz7ZY+qY4J
qY3JzkdBJ0S1KqLbKATEyw06c3AAvW5efPDwwhhJORk7pr/i9nqu5nijscg32sp+
zaC4zs07Sc8OIoidlSucHlQZGPHt5n/TSpqWQ9uRssb2IEPJXOFMzAW9CEmrfKLV
WIClY38DNRJJoboclRX2NFo9dgypQ5Cxy8F7sF6vqipqAiqq4h1SQJ6Vyp11ODfE
wtMRTVIz7T0QSa58KwslNg2mx2zopoEcfrKwRhIeMBtD9ji1wvmQfEegTAtwQewn
l+Hf4dyt/ikJ1THQ6HuicSR0951OyaOlpmfUU9W3BRoAQzXqMcFrlqGJIl01rzz/
0xm77wnL0Ju5W3P42a5UKAiXBCJNKSKINXVDHMTgltVkwyUpGyXSBwC+XxzigC8P
pFW6MIJkNz8ORvXgLRH0qeNqNAXKz/wN60NxNZZSwzu5SS8cswMkufIjRCEy6euo
/EJdgIzcta27UQJWD9xol5xXzDRMw8zsl7QQMBXo83eisgLbV6q/yz6QE6eBcQxf
JLReJmR83JOOiH7ys3f3I1W0+SnZoPoLPWWbXj8YGmMj67V8buM+mjrkceSteu9I
YiupLgZ0x5nAm64akQcN3SdYQcjLOC/PwJ0qu0C80x/4lVGtsgKhgeVqeqFDrqJv
jGkL/Wy/3kcNX2xUIljcAi/re9KohUyGKmmIEHuFYCyM3mBxjcRxWcacOcjO6zek
etTQhsxnMgSNyitqjMkZcAuYl9b1X5V3C3e2BUpM0MEcTfRW/36x2YEqoO8ZmIrD
t9bmVRBc5z2z8/X7QcDZXUJOSPJ2aAw+74Y4WbGdPyE7pAxrd6EkOZMFIjY5yw+C
K4joh+N5891Qkelwo7G4pAaQUEy5ke+lopZoEEZFaOILMTYtLgiZp9QgDM9X8Zyq
smIqT69SW4LzBFuuRRJjBJsb8266eKaP0yfKdqPHwt/M4glLKb6kJCP8Kp7PcJX3
tVeXVGifkSHFiz72/t6IPVbLqbRBOUrptFnpp061wG+PKbLQYjBq/FMssAG7Oc64
nZkMyYq7nn7Y8BEB+u00ACo0mC5ML6/iz6PJ7OtfS569EFVeLJnVCPdTeI0RpqgN
3vlETiIccTkrVkOblWIezdOb9nBB56FNt+Z5w/dgiTg49wA7epMMpCy8WHL4P4Ir
1uhNKQpRA/IdCmGrVh/ruvb1Ue0cqOp6gJoB/yppnRaafhwvBfOpblYOxrdAqlmz
YgRN1VHQIrxP1WRTvRQ2pyEbBZHcVMyAopLJi094ZQHLhdgaPFapM8qczrtzZaEf
nPfNOmLcl1u7Z784GylUfRAFgLDwDscyfpB/Sty/Ib1Egqj5w3WKmXhcWuSa0uYH
cvzOZmHeuHw2TndvX/UfrP4ofBHxcBW8ueaJ3dFDbK7CKCXk7JVpsOeM1jtMvbpY
/rbCUmkgwWxF5qsCpsiNnHMkFslRu63HNCyse9hPYNECulVN0frWP0UaXnl0GFE8
rYXj0XkVInq9hFO0McF4dMBFYcVmgdHgwQkEyvnA6POt2mEU0KERBd/nFlYgNX4q
HyuW1x1CGXfmVO5AFfRGULt/W6QEyQ1haIlvdm1z3/DK5FsXvc2CbLAyzouqP6Qa
aa8IVwkNZJb9p7LbJ8SG+TFmLQhamQeUBF1QZN8u7kpthbaDSs3QOcuFZUTtY3kA
VIU656suoIILbCf7z8IJSxCAeS93paOpHn+1TV4LD3WCyUqYB+KwQDdoWHNV+sNM
KPAAJ4SkS5EU7thSED4/dzp+/PH+m3zTCYEYrUSaGsJ1Wu1JkVricH83pus4VLy2
g+vpQ8uxAFzVlA/zH6n7xWSo9q0wyw0QIFbWpcnbX7CcS0a7Efw/hxAVPPZ8uR6l
ZzbOU1gPzAq9yyCwT8LvQ4s6y9iATyzevcFTKR9yZkfdtFhoE+7PrULkHNrJ6C9N
QzIgUqq+oaxhjz7GERvzooMuqj/LZ0AkE5v/vcwPcE1kdBM/Mqa8O9IP72+LssFt
A4EMbvEZbAy9NIO6HhorJjoXDWMfHsqG6BpX78pEMgjw0hlvzF8Vi+uxUKZoLFy+
U8GrZ+UoGq9BlPCA5hLMReALVDklMahsiSQBj4/d734rLTjYAXkqljDZev3neU/J
Hz+lnW1sZJveAN1+5ntU2+TVPfD20+2vWHrCty8oB8Gy1FbwSF+IKaRkbbDjQ/6P
CASB0wZWsDZ23g5MQskzwLbk2wLRhtCXKSy0NO6IqgN5PjCkA3EbbZT38mEm0OxQ
hM7vw/XlkKMna7KHghDrnYzlHI2B6XfcKG0E6XJAfXUMiPA1NvibVAAFtHSMT+3X
jFoqLuBXLdAKPGoGwBwiadoPIQ6kzu8jEFoNQ6Dj1RSUi5WAWrcCvZbxNderR6HT
Dgt4zr/iWZM6tOtJo6jHC9lg6iu+2cmlLf3l41foXSmbTNmvvQ+JT1koQRHDpKNx
DipZo2fw24ZqXq1rdutYTc0mJJ0JyDKs8pAdNB0yVHuOlleZwdU655e7YYIjx1ct
aMz0dAjVVm4NZAjlNTooz4NWUsYe8yRb37hDA2Dw1jfxnH7kd9JFVSRtK6em9opu
K5G0I+wr2xSkjtg1A6dGodBpoME9IkyhOUYSlLTxokNoo27AD+94Sdu5ITn53o8V
op5pqPfjE5GG4uuKXUGDxH7rza+pwATU+5fD653Qo2Z6JhP9I2jmLFVkY/P0mgTy
f1G9anhASZ8l9BK7seYYuDoDFI/tzjxM2XRCV/zwAxF1pfIzcN8MiODvwLtKehgV
jDjR5cSg9jTffFCmpbuxdcdLFPLRbhpMrDSMkI1pgqZSdRHmFespBs3t5uORkOHX
X4iCcF2zBW58QvzX+5JdWeAfhYcVzeEWfby6IYhE/GiE4v/yHrse9yOTTpgwGaGS
oHDIPtM43qRw1f476NYHLMq6Jorjy1HHPPjoeFm+M632Lci/Uy/4pTxA9iFkbUsc
0Wjsd2RsoTl0be+kkJhtZBN5qWegeH1Iwp64mTR1OlG+ZqKcDL/PPqQtUM+giIA/
zur20ejHAjPx3rtFe1noR3OggnlTIHVRZQ2fV5XbwAviPpHGuUTyDKXgaZ7rrnTB
YRDyR/x/Z3Rzz8jSyc1kcpU6Bz/kU+CJKkWRdcZ4DtvMlpDYmIN5ySM1zBBmI6Oo
vANrl8SoW50dUzPmMhf/LSFJnsIH/uI9YtmUXTJdQiUBcCFXZoNI2ET2/qNmyWkz
4/XKE1ZhEo4+6RtM9KgRcId3FjfmEs2B+BW4v9E6lpMAtq3ogVElSMpWQHEwYoM2
ylgPHXpMvBz5LNz1e+jaLoyzFdvTam2EJRD7hD3OPAH4EYgars1MwnWli6NG48xz
MijCfDr9QUehcqH/8edbs4Ex2DDg4+iJIKrZdipJP5AdimIZTjDxMwUC/uss2hrg
VHLC6//nbIkIBME1Jn+hdz7Gnmo3CnRQaYPlM3My/NFlyQ9EwfpSb10Hbdr2CIIq
EDEyjgda49+0afXrpS+e/2yT/fe2xC+tujPFLP6bgjj+rqxyg8WjGw5RUHSJoxSc
SqDqvq7eNRow6PRapR1xOuSXeniXT3ec7kb9GP54aON3OYiZDzHpLQPvz38xvRAk
7aPcxfZouV1sLvBPR9J0cvgGAgeUqI8ANXCynkaLDGHuDdAzsol3UBl690EXoaEZ
MCxTuT2cameMUopBvo1ySxcN3uUmKAMUkQuXdbQxbX8HFyfi1pnTbrl6p2ChR1xA
+1rYX7oJgeiTuW7Tjp+p9OhLPTrfAJ/6ysqXvdqLLEyNVEyNJj4tz/So9gNEmtBZ
uTrxpLz0j4MnGdCHSAc89ZVjGp4uibBCW8/Y0z3GCq9PYMP82TgqXWeykaPD2hqw
LecVi/IC7JTgzUWbD/O3fy6GpugpkCnL7hzUbRwCwLVkgSjLFUwq7f42ewCDhEDC
vfdbQxJyT5xQ8YR4UaNLXUQ8gjZSw7+bK4JTDp5PO0RDr8Orkty7Q+YxVekkpg/c
xxZdxs6Yua9AIzTlGc3Vx+wQJfwlkRV8QAZIR+XgmMPH4ABsuiLdRLBa7IFK+7Da
6fmTOs71Txhe4aEIxMinKr5O4G9AtQkhARj7FBygqR90fJkb3RKcfzzcbZK5OWhw
9smq+r0/5u5sobly3rAbK1dwXZJu7mUYnJ/+K8y3i21cKa/4UQG8t+Dmb2LjXLc8
tgQCIwray/wGboqFGJe8+V3VHweFiluUeFkq3VX7iBM0FCq3ex0HnUJbKUkFjXko
tmixdFvtsdotkWE60CL2nqWIFicmwu3BLhHOBt/v+8vOnofXU5tb3GRmmlvd5zA7
bTsf6iX962R1nIvvc+DjrhdVsgSKjgXDLtezdGYa0ZjY1F/vtuSDIotorNV7mMTt
NCjFHcGhKOdkIbvSml2aqmWydd5MbFF+GTs9fZEhIu9MnUkvbaVGgXaS/3EQ7Uku
UFAM08gaarErxPyX+p1clGg4D+j/qqGexkYbeXc4p2qENPUp3Fn8RPBJLGs8N7R+
pjl3K7iVnfQ+T9QtmRT20B5eFyE9MVbD89iWtc8NsvV50/gHR5ehFYx9rLi1iunl
tIP8J1Hfb7u3MYsEbh/+o3+ywKAL4zgMTfvKjBtU7h5lHsPD4bWWDcpq3c6nmLJ/
1TpbMR0ldeY7gkkTL5zu6KPR8TfzSS96uVCg2O9YLFLvzWxNP66HLwcQCUywKDye
grarlQLCv1vnZU5mTDcEtHc6fJGWS9NXG/BAfqCfwvCWEtZuIPNCNpMcRVCSDwqp
iOwkvCnRJiXyT+8I+3Iff9hQQwBS1F+8ke7yLoZmfIoW2rLnQgJU4pd//pMJLTsS
S8zsDGLpB/nPMIzUqnDsCrTIxxrNpM074RHD/mrdj61lfh0aOSBYX1lXAGO6B5k9
8WLmYYjx4FKJDEnY3+EMtjmFxRJ/7QitAVKbR6/lV54NtF95c9Xzr8xt5I8U0Hy/
NtZ9XwAl7uEW3UZAFIVhRcsDzzLlMAlk6sxCTqcBya6idrI14Ay8fDTC6qnNssRm
31oHBcwq8w5t8spwMuNOrI0TANhiQWvQt2w8ChQ5bLnkrrO7JWNbg1kavw/yNIG0
eumie4ljNm/6H2qCyC3zQpAKfHHEUmDa1lkKacNJ9b/EoQbJRKDDr+JcQuguUcSz
zZy5f71WQAH4jkRwRAwhDW5+HYEqW+F1U4yvPuGqHIbeIiN5vMGctLpH+1nyIjAu
svOvvAmM/HZzK3trBWeFZNLXyWg6IhAdp+Kkb4TDs6ogaMJnTfjSKbZRgCAwmgsh
lIzcy1vJAFOH6N3ewOsGNG/RiolnaVY+PzNIU7NmVBBgrd0MsgxaEJ/qZYTmTsuR
1uUcH9hk9zzlJ7SENx9oMaGGdiZi5QuTkdOJ/KnyZtI1Gtsg9vso9xvWsGnR5ymO
O0iSuLoHcXcmf9HimAvyjaStCun89taeX/vZGgQkv/8e0ChSHk+zfxb8rUVXB224
RiLeCfBtmtBu1RpoylaUvzhsS1vNBx/HqE7yiCz4x2NCR/cybjaHDCxUn69CaAk+
9xiSp85ar0Qv/34sWRO8tTC4eP9gp1JIHl1Fty5yH6NCdDUOngrzqp1MhL0hlrNr
z7dHUR8CNfJLgIsFVxkLoqNVVEl7+I/f7xyXNDdSjwcPWK1j0EzEMOehtstLuhNX
VYzCgShGtiMM5fVeSTFyZmL/XWTle80JCAem8aseYD/TS5g3e19DTdmFO4gj5Bo9
G4bMiamZzVAdGz95OusE9F5sOgj3T2rKRzAD1rM3SG7ue2rfquyk7QdUVQaZXKQT
A8r8NucjBf5xpku/eIYovuEk891MMhzmETxvy4IX5npFcZvCD4nBlmrvw0ZGqOf7
cDjagWV5PCmYhuH8sjvq4H1nL+Rndgi/nOJ99ly6W4Z7R5cQ1xiZXdS2uc5jxdjF
4kbmf1OjqDlbBpldgdE5nj7zOWhrLntv/gBLcGn38CWpm2q9PjP6kq+4QigvT1/x
gZlD/P7qpW3v7hgBwvkPWTdVBlDJXwGfLb4U9bWj8IITWfFyiWD2KnlZf3ULv+tV
FnJ4R3Slrk//phHSvVr1LvlSd9oOOsHjQhPBNkRumjzl8ybQw2rfT85/rJ5Hz4IJ
d7rm5HShpVhHy424pvcS3I5Kty9BoBOjOLW0MzkdJevbjGQHnx+L1+eO3F6OE9VS
t8i5zG4Ee7wSczy1WkEsXYyAu4wCV4gPtZi2orxUfW6WtiHSwXMn/9Nq2YFxPosO
G/flR53pfKu8DdJNyzSXf5F+ixsuJpnDEK3BCsV+txrXqwSMvU4CACARrFnkpGFP
JqzrXF2+r0GJ6ae48Sf1cpotG4/cpavZevi9If1H9YOrdYOa+gznV88ygOK2kl/B
hiFl3vZm8A31RNCaNCeumxtK3pBMAY8tSBnfMvZLQkaIFDsoDxtZ9Vh4QYxc9YNH
0PJRM7T1G6MVN1t4Zh6Z4sX5EgT+u8bYu2Y9F1i10ZyRTqTKYqYB3wezs+31vg8X
ajMX4AOyDIPV9c6O5EEKGbHA6QL+C52H8npSat1wsOoS2PzZ7MGaeCue5bsOnW3Y
syG547+fxtd77yGZo1WEcuw//l6qzGiQRgo7KSEcb7/DZCbH0wc0LOhPilJcp8tH
qoPfu3Q6z4aV6at1gwQXNDWfZlYkHER66kNpUQgGOUCglig6hACOpJum/G3+gF6T
ogvdAwU6fY3jyHIkpiQyDykswUan014CSPeC9QntYc3ZN26hpRjU3/E4UMbvEl6w
fnweV9cSpdLw53pR8ocuOfQxcP+yBwq5lTVj2RfezAaKHSmqUbMgueM8G9FSn9vs
M1d4NevUlf7YIjNafXSRCh8D9rRfXExB54ey7I7tVCiif6Jx852Z95IjQJP/S/y6
VzoJBXmysBrJQGXp9NTANGeW1V6PZSwq/tAVvaZVZv7jKPKOa9pa8FW36qzM6FOZ
1j2CPQj2aOZl0Vu0vmyG2j4ugkyl3+UtYlF18VhCO21OTLqojM5GRI7ig8+mowBG
v8VKCZBDSzCicoZ7MJ1+s05hUUh+xqdS/hlk4UxURpDJSP+0car9vjU3hdBe9phN
kMqW3hFhP8Qa2PUG8gOH2/El1lIUZsdsUlELxAXIqufYycqrTCiv2zqJuLZmUt6u
BzQ1jBmxiV1m4xcwD/Bie0fQlHdkFvKx1VLvXGPqiVytmMUUZICAV1kCmm7PXlbH
4+men/CgLy2d1LTYuWeXdvAEu3+oBFKN54kx/jCPNOXIEpxtnfD6V8x6Tvp68HZ0
NQoypm7Zb+RAjy+4EpM5zIzG2YmQvz957bA7pfMmky3gm0Pi5IW/JSRl+s9/scqh
XMuyjNX6rSahpatRmJgjfeK0RVKs55qvNhV5YY7zQT4uzOxstS6AMYSG44j2Qmzr
ZKqg8sNXjpPDXTycLgobtDIK/IeRlWCj4I8GFl7iUwsVU+f0y6mZFpJn3Pthdbe0
BP430zEoX1jc7AW5+oa9BrMpxijwauBkn0sjS/VCPXKNX7hDIV37yToz2h+7LMPk
1DRED8xTA4WG1Zf+lQ1AdmJgopUW/0CpQhGscK+LxRCz2M7WghBABboSGiitJH5L
Ie/ch3lglDpkZQeSXeA4Eufh6Dyj9dHUhu73Bj343JvwhpV/UBt7LXj5224zY3r4
YtCvJqpAV/40zdkciCgBZYY19M252DpQ7YJ49fxnBv66fmDAGRwReqW1OK+ywbgT
d8SGLbCM9KCX5LtSL+ukbaSReYusFdqlhnXYgWDtop94NC6HaxALJzOwhrgMPLbW
R+4UzJLoe+P6FCiipOZe01SQpArU7Crb84G6CRqtnOpYn3poFlwS0FGT+66RJeT1
7RZVJnpmx45s26C0Nph9BFAfFf3RUPUO9bWIALgS87gJYVRGikz2NgSSaiOD33He
HbGo7YSn2qltUh00DolSUHcizi8uQoqCq0jTOvs2nHKb5ohYgewXKhAq/1ocm/6E
k2Wq3Z2mZHHsyzuAghnjK5/WWDq5xfjRtQMOazLE3uKBP6vhP6dnpJN505PQ9lcW
tiqcIzQz8i1QxLEn13CY9wnFcSlcvSK4CcMUaaUMAz6Va91oc5tOMXpqZ0zsLvtC
uEk3q4BHZCeBKHDTh+TFT+rJWk78kGRjTBm9J5qo6YmmjP/kEkTop2R0a5F60oou
+ek+js2UCQq2KblYb+XZa7PssJ0kLCY+qC4rZroi5uWPPIblUc7gWOtgAZPBY4QC
8VGQhTZ+uMkOpcqBAj9+4GiIl5FgKuk3F3rm6MAYcfebSOMshntY7lyJbzlOjQex
Is6DT+CHwg8chvucfTpF4kimU3WwsajsGqVb+EE1Pg+4PPlsL7ur4w8q+K7T7vS7
GQEwckAGPks4rKznkAYFv95/+uUHnCRRShYJkewpjbC5EPO4XbOM+dht7xd64yY6
kNpw5lN8NfUR2rpNKRXY404Ffe1CKOiWOyVaZhGz/fkZjtVtXP/rbvGFM6ucykRg
fYz3qR4FHBkyOuaIStPeYI55VbjIsomJ5vx1zG1oV2HQO8mV8a6Hx7vRZ+MD0qCl
4ribBY6E9z5+0KIaxPyH4vK3crLwIg4wOYJEL4nsoE9cuTP0W/UYkmP2mc0zRLCk
3fhD/pkajynBp7xy/4JGEcK3IPKzkAMQn4/qHXpThuBhqX1dR2pZuiEDv7/Etiti
bd4AeNtcA/3+eeA04yJzUZlxTBj60xmjWztji5iJ4OuhL0gm0pd5mym/wCWqfdln
PC4g/6FxMQ0IXVbLEXmuSDuoiL2pFiFqdHJGBLR0dXSjHgsWEGwtS+FZWkQ/ZWt8
YZb1InQ8k57adxfPGkhZM7sdZNEqDh2Q/7RvXR0Q212SNXlkUCCKySsNu1jxppA+
WwAXzRKXWwzpSv8AnkpxgTCg+AT48qNLbHEqI8uxAtgydmlJhoxUa/UXumcFDkN5
aA8Z/8fMPbFhfZ3DJQLm+lZ3PCs7VmZ3YcobdqbqZLTPZ/BJa2on4CHmsMoeIB6f
elchml1uFf7PhRJ9YIBYSsM5q+VywwnxXHiwfdAH1l7ZUzBTL/CiX6y0XC4wxBHl
ITPz/LckFHHYbAbnqN4euNqC7E5uLiawqvRmRUpq5prpYa9uXGK8v3qsiTfRwVbX
5OB6g8wUOjBnRChfgb8umhzK/c6jZ9+Gwr/JVQt/CzO27YD64Jg35gKyP7PrLzi2
FQT6ZTfsQ3ckCw16Ks7+Ey7aW+u1VgNNRrp36y1yqvKIWgyo/cpMqnXk5/dyEOs7
7EQsEG3QDyBPut5QEQlvEFyfCsIWYUszwjzUGFG4dYw611XbRzRsqJroKj/yp8n0
o/e9qjhaM3w5prd/FM2LPaUQaWiQD9M9ISOXDLP1++jY8xcA/idoMeETZB+XjIkn
5zsJfxp7UU6wdLNGMQi/7O6U+TeADNgylUaKEHqynAsZ32P4k64cO3CVVpZ3+cKc
j6JJogGdZpfT/GpCUCwO1dnFOqQnbYRp4n0fHT5RDQ2R4vRy/n8YX6LQ7fqqoGP+
MGPVy5cK3sfhOT9yksl8KQ+jhXgrnSDLceJcUnaJ4cX6L6ZmXqXcrp+w7pT5O1cN
hOJtr+vkkaI1k5ZXG1L2NaK97dhAO0XBuuNNEzengQAHllrsT6uRjqNcbVMtUWT5
UuzJt3zhk4658A7Rx/v8WemLa+H0NeozR1ho8VA9T3e2bTUR/1zvhCupDyIYoZIM
NjRAtNrXfoZMoUoHLgjqfG/rK2WMgSH3U1VQJ95ruidci/FbCEjCmsqbzWtBCwJF
3pt+LHgFB8F7kAryevZhArovuoStLrXvwO4JX+xO+Yn5OfHGUDAfs0ZBVl3ud0+K
H4T8MRF22GnFA/x0xMlEAysYQjGCNz+kVUn6If1gA11S4sDq7G63ztuB9Jym7rzr
WvlL/ZlCAKbnspvr55711M2MPlwvFutpWwmlPgdzXzQ6EbNbzpioar0axHHszR+5
O35pKSTB/T7v3Adhv3myQkxOW8PDqzP/FUOzgKzZXbc6P0p6ZeiC14XxTpgXKAeu
8F1m3reQHrbQXzKVnLsDEWuhumccwGpSyRzReXUWGB05e/vFh+RyKVpKBbb5W5rg
B5m8C+d5rPlp9kI4Rp59x86N5WiuAxCknQ2WvUKD+nj8D3FGlius+JkIOX4o4nSg
GeIqnMZfjHFu7hw42FLyB593yH2B2JBr7xpwnkAG0G1UlkXYUah0aITlTgNdUnGh
SP+jPmqOmRvJ2e8TllW+Xus6zJl+yrUDVvxIO4zKH6DEwVuMQ+5ULsE7/pxDDMO3
sYVgD/SP2a0Jv8e2QwLmRTT9Vlvvg7Hs5wvmknK0RHwUdl7qjMV/TR7RRqEFvQXO
ilcGKWEpuI78ovObat4aLbXft6lHMISkRLlU6/lSKXhqn3nndR7KN29rW/493X9e
bQosfOYmmPgFheanl2agkj1zZ7IHk+8KgmbaFiHQA9qZiXmkI5zTIM4f4yUYF0+x
sweD5Wfz+GVQLDgUaOaBhrUDt5c4OJEDFH9qxV4Fnf+uiTpBg4+DNF6v8J9sR1Cx
/aPUgwg16yANEn7oMrgFEfwPhVHkWtuHV8OtcLp+CC6oMcbCTglL1Cuc6K9nZ0SL
cBKiMxR5hfq9SZKoWsJFuH4h+4LtupFqmnqhwJx2soj6Vrca+ag9kPuLNefViD+x
THGS10ZxtewotOFCLOn3ZWZj8euO9/UOvK6YGP/EOlntHMihsASnyPWv2q6EJ8Un
fOuQPT5GdszzmJAF9YT/D3Y79DzgDH6mwrnfJZd4QqoZukymP5NM4LnSqaDTfJyo
Bv/rrCTpiVNY6BgabAfdTKdWymt/Q2HF5HNvpFcJs7EGK7hXW5rtPfZSXWhfwNr/
0Hka+EdyT5W+SxPf+BE4NqUSs+O2lSOp/BL38SPByqayXbF4NEDsFhqEY1MEJ1lP
yMQ6JqTLaj7Fw4VeJDmV5gwpW2bDbl90lh6eieJ0VBZQ9c1hsbWcmN425/Gyvj0b
QfuvsW3HFiEOm+4Q//P11uwN/I6slAt7P1o++/8cshvC61+3RuDIEDEKVbZX7Qgp
/G26eCUAyiUueolxsdFxglLZLGyQ9Uc2PUjCNjPwHp1Do7sB4SNE1hUF4M3njOzc
3KcnSTbTrZoL4ov/o467fNzvKGynbRHMPZGuRXXelaxbJFFy9BTwxiMsOeC4/5l4
ZHE1KWFUifLWbJoEMH7P57gkrYdceakwiLIWHGY3nGIfwQCeyTMPCyo7EhCG/jHI
l4KUTVGFi2tbyXd7EAoPg3t7IduCyHIm5EQYd4dp4oYlPuArWuf3VgT8CtXCKxB0
3sA6TUKw67dSd2a6TKEqGvrnVDH7YCZ7ZcTaO0AhImbF/xojL3jmg9HkfRevpJhl
l8/5n/Z6BZ/LDTnRdJvey7MB/dfxpWMKmCPan6fLwayKAZ9sAOMOc8yVdyB+pP6z
r/8xvg0UcQgXEbG86Y4cAfEnBCj4YYlQepa8CBUrwPMGckdIOJq3LZzcbTijIFSL
n1ASzV7MEOvhE+q9QFVTK5gI7URlMsgd1Y/2nQ8Vvvl4r/DeRdx+pTpobsZ/biYb
6ORANutgB+9gbFe4dpyHivhDe+yQ0vcbkEKS4IEz19jN3oY87aBhckdxLAQZWeSU
BzkRx8ucWWwxs5/1XNaraH6ZjX0n5BUv7efEtx0U24BxcLuqKh9YUAcEGtovpw1R
EuZHCkEi0Na8DCQhgEV1k3KplLS0eCPoRoAxK0zWlMfiWkTYsiYr8EjY/J0B6Rhc
LK5xU5KzSe941wSEQfCc4WSZraSfzndJCf5j644DjHF35FpGzRwVxhiRxIkGxAHh
jLrpv/bkbolJ2m2eFkCyQd8DJeb0BqkB1c3uAcCXQzvI+/B7zOSalvqIZWx8LNcv
ILDpBWbS54zS582irNjCV3M7ndFedUFYucxgy9MLyA1/nbIyW8r9P7g0wW3D87w5
UUA7HCEaOu5JEMk49B/g/64EQorZltuB7gquirE+QYKXTv/KZrQPW2t2+Uzmhg2Z
I2jeRz5yMFwE6dt220XAKBodcvhpAOfhXnYt+gTcCMSLrglvyNbv172eXAEkiE57
E+Hjs9Nybx+Wt0wA2pLxJTDUF/Xcn/Fg7Y641gpOhv++cBKZ5gWv/gdPGqKzlIFF
DYNS1fMgb6Olx9qAHu8COO/PtM9dN3e4kGWtrTQTLrMT6rxvZLPf3D3LkDZBQZ2C
iO1KYhXF+sWPvdqLMuHviMIZBtCiK/sVICuo9dQJuFNdna1jwQ3MRTfDQasBcPZg
89cP+fFK53AbbaYuWOJdq/t5z82Suvcxi5oc8VlQRs2CtGcuzLoJmfe2c61Gh/pI
kXB340+GWfBmMwscTgtafVZt8ReoDTTh7IgF3mylqHpkYcSgHDwlXd6pmTkSRzrn
yKyzi6tAmSLPJyLZm/BB2f0j2NzIvK0jMFiJmBNx0afOvhnrfZhPqzih0FAYartH
tGTwIs2sBtE8NxsgCVheqRQeFbOIlYmYkKXfYLh6ahc550GioHZ2s8PFphGA/dBs
TD2+3/PnLgPczbRIDDcOU7SQYuWWSh2lTYJjcykwCCm8qhPRBc3XqhZSzt0ICsiU
VzsVRLxG1C6XsqjGsewXmKFvBYKw6QE2rpSd3/42AQXShjDbqplcv7zvbBoPsw7A
CxcQG+9fOkCGinNg4mhsURhZQrjZeCroM+VJUzz9p6gOTGPHF2fo7YWNxScwZjLt
xewK0gwJb4UzGzeT8yVwJ3jLjIg9w3W7j3zoxQLVLT+2CRgdPbbesrl4glFW/Pk9
6AN7gx9btlQE2b8R88KHFrEnnTwnVTl/mq551Gxv/1yFp38KPZsRJiSfWA/HCcFL
2J3edQvaq1rvZJOOGx/dFU/iYsZ6HJ8O8uytSuLtC/NEI+LTuj/NKAGxzFc6A6b7
LKlw88iG/pwcxQ8eXw2dJq1VETV4CE1msraUNE0NoNFqCNhdFL50TxWxGRDwY7tO
IIu2/7U1+tVUGmvIk9nxulEco+5rgSw6J0xTQxszPkKfOG2rt2il+ZRiO/U2bVV1
ELDt4Xg+wCtcT/A3Tcm+w9dMWhyuGaIOnQxRQNm80LkT1x9lqbM0Z2EzNoSNg5qG
rnmc2QnG27ze8LaZzImdY7Axi5mJmC5v1VFYCiVOmT0C4m+TF3NrGdHW390fSeFz
0gLTweXSYSPiDCsRnmA3dFjAJmZNKQbNF4bdAxnfA6DiFZuwjQVm6Ivfkv+Syy8W
yY52y0XIWMnfhlFlLg4RwIGCteCt90/rDPfg5LSuLkU+sszEXIGd5uG9zEMsiKy3
L/C+NJn2tsFdPiyMXSv643MT0Hu3fzM47AvERNGuNPaSWBjhd+MswM8iVgAxbpZm
9/sBULb1+gIqpVNfO4gqJHXA2S5GlnBct5GKRhhv17iobUxKcSYVPNpYgw82AN7e
VVEhVVfWJ4Fy5YluV6VAXzVlWnFZlMmg/+XNw/61f2FN1BbzdWzBPv2rC9OY20dc
mv2v14xAirsNNkcvk+QXXgsduvh0aAU89lwFuSO4o9qgBiAS0AtG1F56bK9GgLFA
+crohLv2Vo+BWXxsJxsiWMsHY8yaCYb21/LWd2hj+udT2qogg6bBgTCghLnT/YSp
WM4+I8CZsQFg8hrcqJRoeuHaPsE9anWs1SQ0RJ8nNQz4+6Py1n3GpTrjRdoGhG6Q
njLKusGyPJlHfyRiemaDq4lcOeelyEtXIbAf30lMll9jYMAeWB0aY4KH1DxFf0yO
a/7QnoJh4tIlxhXyL7DBYxOc8kjmjRtGDtGofByFCk7jrtOFbElKhmewP92Rn4vZ
naPdHekssQHz3mgctK/mBHBiKXw9OwPQpTWUXMfpc5jtKHCKCy7JIIfwBQQ4BIRl
dx82cn+f0PZv1fy8bxwWoFwwlALI2z8ju2LSeFQt3xaa72IVFNLBMYO6EJd5GDMR
Z2U4DybFz/0oHPMjEecdTmBoUqOcfdHyZLq4h9u7jBgnRnQ3RT0K0KCXNjDgylVy
HTNxXpvWOH04IbV7WRpxOueosHJkKWtgZUGVToKFkUYoyjTrxVi5TwDHyuskVsc/
v6bXjFqw9StxKe9hvNc8QfHq7RjBHYj7E5Bnr5hERloLmSKZ2nYZl6VJMGGuGuFE
DeTJf+/OQebAdeGUMpzfEddDTXD5lpt1BcPyHdgada+11mEzJK6fzyzWGbGhvxen
T8vn05g6l/FgIlHQrCL4y0z4BJnTx3JUOzuvbhBZTurK/8JSAsQ57sOc9f1TYJeo
nVLMmTWNkyuuqrMvqz5e2EECCVQ6dzfj5pCyy7lw9IqZJ7wD1BtMqmQJJel1kijW
w0YPK3VjK2sDPFFXS5w1eB9IacX6aoef/R5OC/O4/j0kTSbccunfzwZ9N5tXozRf
GSU9GAfNjwi07ZtmNRggYa8YUF4E+NsMUyO5Nrv3MBXz4NGC+LKV+iq7u/A7p5oi
pqr2aAFlEuVevXA2T1Gq2z276EpwARq7i6OhPDq3/uk2ApVAg4YhNjQnOXfW8slN
7TkBiad9os578+00xs7bMf5FLclzExjL1kYMDlluH+uerVFW8FvE8Cmv85HEx+2J
bWzN8x1kt6rje4dbrc/bCZ4GXaJAh+rRiHL2bYheD/eTDXtkgcudwivZ1NPPsmOY
PdIp3Dw3PVNbEEP5lwMSxlx/qEvmwk512WtfU/FrqOwWjRIyf+r/VODt8gTRtWnI
XP4NJmPFyO0+TmjKtJ5xL1+YwBlxMWola7OnJtKWqQQtZOCpszMFPppnNIpvToIV
1InDX2Kg0M2dGO89e7gNDlKlQWOYjyow2FcoTNM7mg/gSaBII6epyuAYAHL50Kkr
VNXEhe3u110NKpd4t3qAujNHCWtMMa+yIYufbzsxvB+ZPREi73jAtFPPjgTtM+la
prQ0s10/5vsI8iQXcPtahHoQaLlmTOQ2jwC9KyLm0aeELhNo/sU7ZCu2yhyJyXk6
tL9R9wBfEJpuT8xlQXnU2gnEpA8DxNn+tcX2BDq5JZooFs+m8YT58SfeiR643Ptw
fF4I8O466NggnWTCkAA5JskdytmMbWOufufRcDW1m/8ds3jUIMUmu86hG1m3pVzh
RrgsRz2npt8kjDN2Y7eXtxLVx4eRSahnyKt1BwedwM/bRtckNi0P4ff9KCwfYUBl
MPfnBbBXd7/xmx2/ZQg3kRS/DQaD0K7PiPguoFgEwvE7pNT0Z5LO1HbUNlvsSFbS
5YLx23hVHJiyY8ffv9gj7ObUbW9L2Zu7/r4YUV05siOeyMZGXnLFYMMmyaBhL67M
3jRPSEbn4liKWhP/cjlgCjuXslU4Za7c9OrA8lXANKq+SRwEiwDm8I6AfkbthIiO
oOg6cvH9Er/lS/oong8awcVPhCBMtOx1McinYHDFVK0bidaNVn2YN6UZQTSyd6MV
meNwUwP5ElzbX48+KYIZmOWmForrVXp3E/2l/Px+RPoZy7yosTrkp3PaWuQsL7Np
l9BMryUNVXfKNtw1WxpI5EAvKQ9Cr0SquvEgZMBdaFykdNrcsuTamAmO/agpu75r
HXRMR/aMPdbikMuj482vsrmawLyrErZmBnqiWeUJIjl4kP2iY5vlisFjUxpQoV0c
JntofO7thOGdwDTjf5wowUIf1UWQy/a/hbsrXzri1TD/ZHAQMUK+ObAMJpaGR2jA
GTNEOTv7uYeDs30bM3+tqdCSAD5w7jc94NNXtVmOQjlUAyOZwAv+oV1FV/Zu1LXv
/2cc4K/YzRwECKTnF+p0YBsOp98ZvfCfoYpzYk0YW4zJQ2+1Tbml6u8T6S4v0a20
O79NPmpkQf6vVL91oMx4MYVTcYlQkYiEsEX1YvJ0aSKn/WI+c+F6vlf7UgZcRgdY
kYSou9i9RJCJ23roEmEUFsy47C2dHqFa0xEtUDO0O40P2RTADu6s+gZpYbO9LBqe
3BvfrPcEnc63MoO7r6h8w0IP/I2SgnihGgjaNdRG1WkiC098Vj0qcV/ssAbLyHBR
FvnQkqqTh6exd41WHDLL8G/BeEOlOpzZBXBqkVCIzSq/4d/yQshZEh3R99zLNR6C
u7sQjmhrvDhjsaCyhrnpObcSipbs/1nCA9LZaYY0GVOIRvbrmLTwpoUErabS7BZH
x+YeYb+3aS2hE0XZar68r7aCgqRVoZOdO9RE6WCWFCwR811E5i2QsNt0QjYwOrsT
nOIS7NO+2vLZXbLIGbtZeWbirLI+bHiuNtohnNtCdNmTqFbP2Sljj8365cVZMUZ7
HHLcHv60KalsmwVP/x6IOAOcD/t5+zlrBEfevKn413nq/l4ho4DE8kaHUI4QA43V
jBkvkgQFdxeUKr83MbJYHVw7+3dyP9FunyHejBX/oT0XtqU+jQWOCA0v9KYn0EDn
I0KAADgv14RSkUUTqFNw/To4AcFTZCBMGi4zz/fVI3cUDmYFAB1va6XkVSKuSW2N
ANwqb/fsKrj53s+f2TbRSz6/ahAI5NaPc110NYZOnoayGd6jhWg2cCMgK6GX/SbA
KZ2AJlFHk/qG1GjMt5OjVyDp1CFgzpd1Jc5d3ZuSy2AoDFdrOf0xE5ATsLJqiZMD
EMnO2z8iPP5S73JU/iGsFGMhLiZSi0g4ztPjI7Izq1WME4fJx7NgmbRRf9QXQYVg
37m6Jlh0fIJyP/IZnQc7N9EhUi6hJkYj8zkBw+UKRY/x+/EP3BZJFxyEOIjNbElM
G/bJZvGG6AAK4sDs/lmy2p+eVWCoFYEfIMxzZJn+BPhnyqs+rtrxelNVsYfK3XAC
jVnO25CNSAt7g5ls93KuZPTG6ZdoluLMY8NtO+Mc4IcEXj6RXHc7VxaGeHN49ML/
KpXabJh8vJsTSUWNWNZmSu3tjTxM8mh/i3GMnKIh+h2xZq0010AZctjA8GqLcP2o
WzVki/BQ09Zt1KUe8PMHMCeQNEHBgbRJOsaZ/EFAeSXARKXVnntn8jFdPULO87rs
YfFsyoY7bts2P0RWxg4zegSaEw/qYlP3vXbq9qAzgzXo4J0jZHGuJdGmhj302cjD
l6xxFyPTwAtAdJ9JJr8JsM636vU0xoOey7Aa6g5rGsmHpXxtNLLeA7BM4+J9uHRK
HHNN+DczN6QQjO1zL/l1cQ3M+w5DLP1gQAsFH8Tvl8IBDBlWuSRqGbqvm3JgN/Y8
R/BF7D0J+dxp5dHNNf1qcmOFXYWK6MuNUMG55dzp64VRO0HnNHtguedpdsgmJMcp
rfyLWewdDxrwC/LV/B3kpBEAm8xQ0eQBt29E2omBW6w0sC2HRkM6jAzNM7kihxPm
IkiAmPEEh157LFJHlO8xzqlfo7kbv+g5LMUPLTFdWM+aSQQjh4efTnkpox+p+9ur
Dwag89TpsqBokKg3mQWVhfuP0tqFS6ohU33BitH95R3N/7srQ59aiEfkHbMVd77E
f/HyJDvsp+b/SYW4NWB6dznvfrRZgfhOMpSwqGzMhCFy66GGjGFCfUb2mBJTxCM1
Ose5vx3EY14wKA57f1dvzWdN00A7foG51Q4B3IYo2K90BpulOV4HWufq5BjSNhG5
aGvIm4KxreHo5PHquVcsP1/OeLdJ0XyXbWw3rMChQLRoJUqyStxosaNbACDI14Em
jc4FgoSwR7Ks4wtgnDintiKG2CDwQsoIBiWih/pCRvP8OOYbLs4JlnrPt5KCU/Kj
WJRcem6xLBB96X3t16bNMf3PKMna7z/ZVl1UaUkKAa5FjEjZPZuX/XuJO+STw3nq
WKbDurqnEZ9edx0iDFCxPxUs6PB+5q5m9Q2JhvLIowESSFaAKm0onhs6JCT7SWU9
3T3OUg5QyD8uJC1VpAJRfajXEM8D3+4oJHc0EXf2x2vNwM2Xkc4AfYqFdfIe69cG
eWhumElwT9bqktmjuS9lS4Rlt/W9x+vxWph4/SvRXHzyS9X4J7i7/ZcnDI4BI334
QuHEonEEDgWiWVw+nx4Y2AoY7ULQbWPWnw0oGy3Cba/Aj7qwIS9CwjtUpTD0Zhoe
7IJIo87NhFkSFLolSGEx1CZfh10iIfHyOz/+343zkE7gg108sBW0JzWC+l9btr+C
IeIiYGj+lNWvwIvztJJRqiZdFjhp0WimnPclC2OtremgOCP/xr6e8MmZuWmmphTk
DZpZENxtq7lgsRkO3XrCsx2LykxWcevc5UDTLTImTXFrzLq+Jk9KZz9XryjD/4lv
kMqcVoJ+110D3nc86KWK4cei+u1fX7OVlB+TpWqA7tatGwLQ2OONn0xj6BoVT+gB
tnCRf2FztD7gM8xzPsB2gFEzvQ8h4HNVWn4fZxaZOcDiLqKjpuxFwbz3BTqBovFH
5L9X7uwlWMid802RH1cKMN4oUAJ5gYqwWp3ME6/If+QjTC2sK3yf5gnS6Rpx2/zD
DLyqog7j838ujR8CUemPr3UrBg0SSkiGN8teEckyVrpBljGXCnPqAQq9+wl0RAOK
orKwobOY/n19yIQLw32ylnOuxI+04Lr3zz76y/aAo0d+clP1c+O9NSRPtvxMPxy7
m3+Rnl+kyc/A7fpxY43FAuKrkuaOXkNLdeGc0Ojzbksqc0FLmkXQMT/Jy5CIhhlh
lbwnbIJQ9alqWMSkGJEfsEyzeo1by94IWvWdfJuZ8pUvdw05HiZxX3BKwE8evNmh
j/WuiGYL9y7nki7+iSQTeZVnD5nA4xOSoT3fQ7fKRk3AKvdkwMCQzLyfB9K9Ek1F
yb6PEfw47n8zIciGGt5eg+rHG/Zd07bG7kNoDqKNDnU7RIaR4AK1092dZpZ3bbBP
bY1nvXoAcIxkTwljnXE/KeVXC/1YpxrwMqXaS8Fp185SU0g+K8V40ZFGPq4NuXOi
ybfUE3pf0NaISXKqMWR+mIodelccBPFDL57bUfX0UDVfE5ml4GO8yQo3tmJTVLtE
ss9MCcHjS38WoC4LJH6wRzcQQadkBiW6D1nrAqZYOaVZ5MrCxGKk/KceKO12Cwl3
eLDEKByNbn/D9InJx45ye//4yahnkogH4VY5YMtApghYOKNfnLyj3DvJKugrkxxS
EmYj+qnZEWWbDYxFAAWZakfjt727exyc1t9bLO69XSwbjNvzTa1Qi7ep/uwY9y43
YmFihNvxsiHRSlfrxqm26cSIlpB8mnPOZERnoYZzFqVd2RKausHfUxo4BdXSkXYb
pY1ycYpBb+Y8n7bS765JThb7kLXmieMBU07llwQ5Rj9IQi1TqBNAm4aPetL+eKks
xCYUPCdMHF3FXDtr2peMshDN7zm2JeL+4U8w8hUMTdSjEfbDr31s4QisruE0tE/a
ZZw9JBPQKvPKtulzSDp7nWJkDeatakfcHhZF9oNzvWOzVGNM6TfeWxLMItA0P0El
QkuBiE1aa35ruBouGHQepxyEdAYdQpCTR43ndEoBzqVQxZh4VGGTXo5RlNWQximz
fI1wuVvSAXXJLR/gB1fkqjAIeENEk+06XNpmcieChUtlGkS9W3ZAXZ1yDzjj/eI+
W33pncZGAX+h9m4AIBT7/n90c3pJvutXrb2+6OypdnUJX1Z7Z55d6d9jktNzXRFO
87uyfhynQpTS8vh/ZDGm77qWkCbwocA5Jdhhqj/GsDEdfA1s08zKrNCU+jtseVZA
wUf28x0fyNOz8jMFLcwbdIGIvqXmP1QUdwdDAGhEqMMDG5wC0RxtTB2zbi/q+3MY
/NTUID/U9dwA8oqvI3jfl7jldI+sZJc0tyhUrtcEbCNc2yTx+ZwxaDlgJK64jyao
XcJ3g0oZlkz5BYvImJ0GU6OEEDe5XRIbVrrqwaR+sO2EUrxQ+5VYr2mZ5sgmF8VQ
de4rpB6I7rdjIAHdOMvI7uuOnFopS9gHfD71w6cYgmVzzsVxD19nz0tgD9fgXP8Z
ox7xPLpOHtn6nDqjah+De+/bD/DqI1idat9uHEVOJGx1qph5OisCSVpd7H/N7zEC
9DW3P/NnCM1v7WIt8sp/w81vwSo9Ov6L1fpVWba91w4cE3XGjakufqlsbi0EnDoe
O/1bc2AnRsCde8YN7NixYdLhSMOJGvqo7tVknZnc7akFljRA07h3oU5p4krswHv+
Zt/dvrkKgrG1C5upOZDmvFe6CX07ZKxjf7AQc+WUCdjoVSNH4xpfBNYNe+sP/Gam
BigojpCOl/GfTrRg9ez7Iq6+G6Ku5/liUe0ds5UQ2908XK4eQAIE0ZGemk9hzAzb
CFUgWXhXLtiskfuQo3DdSsLxCoR5uy/rYtDIL347i+4dGyjcONgOk27BLeja+Rtq
gE/zvJxXcVgyV6fvEAAGGTMTlJShHvlgCr0xVOedDLC5o88u2xWw1mElcNtwklKp
9weJnRdtnZh10qyduOP3AZoKpPyq8mGaFugKq6rdgEhfqRR/d1mLAbI8kZGIBvNl
LCswyryMDDPGu7H1CG2kAa8eA06LOHSfHJLnlHFVa3TIGGdRlbWwKEm8ZF6X80Di
EHZP2UTQDDHMNwgelmsIuTTo1azA2nAHe/CWjlmsynYWRW/oe46oTtDTgLdOfOhh
L5FyyW9+krqwMTUB68hC9HWTZxFANOIkxJxjkusuFuusXMfIe+qROOsOtxWf6vOZ
RQ2Jbbc5cEUte6ShM311XRlSHlkNJGZQ4VNEnSsqc0c98GEhKdEBrWHMMv2Bkst7
Uk0Lbe4wK3GTPtVBDlZYaUn2KJo7C+hxqEhFt5Mm+6f17ORgO+zbFINko/dd8XL7
p2FzEeH5hJoiAoa2LvLPioG8JHBp20w7IReljrJghz5nTr9BoxyjheXCuKu8Bl86
V5b+Cs+gilsDmg0+XrWsSIlsR3DqR7HIpJAWKL4jyS+Vw7H7FdQa0RKBeuWYfgbK
XzUv3GGCHCDhrzkJHUo6aUenjM0JSwxid/NLyDmzKSIgSgepYGsciuv+Mgsq/Sp+
fefjBLn/rGUv0TG+0Xf1QAA9D8aMi8HNNFQZpyRgILqjDqX/VeCiaQ5t5L7lhMgI
o9aWqQyeb8/P1YL5XAjtM8tRylUaf0c/w2nCMcLweEStOxPbpCP2TB+zlTPMbxJ8
Ep8zA78maaxD86KVngKirgdIDn8RRG0b8gSIYlKh4d21VJPcZzPcP6SpomMVQJgp
DZ+tYyTRCuhu9G9JSxsLpige/Otp8WX5ieH6aQ7wgNa5OWD4DmqwEu/333ZzwNLO
QlWqltGkevr4PAtVvnpVN6L1Fxfegns3vZFX/HXUmAWU6lP0bQna0e2aS2wJnlzM
SOA79spkNYNAq0yUa/9HysYzz+G7HYDjG62eUUPii2eOPMY9z3Hw7BLGuLvq1fb6
+QjoXT8bniRcjwuXgVBagkTSXPdHCxFHw2BrPIJ573FxngPvlDmQ9CFw+4l/IxOi
q/Lvuw9QMENOiPKfFjGMzOLzCOKM83gKU5v9aIO5BRe3W1MS5eCHgs2fZ4+twFrz
W1MZDSvegfsY+ABcu0c/BVu2rB3/sla2oXTzuvHr53tU9dlXrmwcIArHusgVJpX5
SZI8OR0XfNgQjFyA1MHZoVWAgwiVg5V/YPnW+N3jw5bml/9/c1P320FixQKvZY7K
hSu5q2qH7mNlPssipdK/aLtdOQtSo4VhtCBXcYwirbYMcp1T6PAb106VGtu7G/zl
YAhm+kF5R0dPDQWSQNGU0lyVCrA9thlMQ5FnOTpqutQIMSRIumHtJKWREmLXhC8g
6m4W5WDbKgkdqvVOM/yjETTd5ITjMXsTqGsCIX3xKhWykF1O3JwC4lKxY1Bv7iVi
WRsm5rj892eRvd5LeUiC3FT5L6ImWQu/+/U+7l+yYTaAopVHZmqm6YKFc7EH7Xle
HGc4FL/saMyMiZDdNeygNDDJgNL5Y4vvnUhgpgNiRnYFzg6XTRtCW83zTBtrGJXv
7bWXoiqKs+CkCzzH4FlVaVhXXikg/UoeASzbjScK78uQAdofZIkp/eqxOVJw9jRn
ILsWEAb5VjO2S1HmN8qRnefSJctb3ln5A+eHs/Eo6BMeWyoiRR3gzVwRmIcy/s/J
hvT1N7g8PxOLYRNmJhrSxm5HUhfYuJJATK3hMp1cOtbC9c8w+/rwRSihWcmBBwFW
j0RgVNGdCmsszuPv0w8BvgsInjg1bv3+r2VFXZjne0JxoH0zPCwKEHnlGjwctGlh
JUd0mY/39w5csKTPILYLaqSCg6jTvAIlAkTg1U9fXbGAjQt/RuxNuQQcc9Xzkw4d
ZnYiKNfx/eH23pwtxhDAlhyHi+q+mUtnoe4rc9kXAeWLymFxFn2gX5p7OV696QTU
VdnIQXEfHUezJ3ENnEd0w5skrKMcrwGJy4l7jyBtkeZhYtBga4qr0/qHnF/rlFzu
FBdYB+4gMnFou32pq2ABYR6SUrEXvKjqbKGEu7ITvV6jeawTepN0Z1ZtWgBT5CD6
ywfST5m8/LEIblpfNHCbejTf2AUXHaWUakwI0S+PF+ZwvTfH7zop1PGZ1qSXvOXH
ljRi5AlDJEF2iPLTjcy3vv6YJoV5qk4zOVkca/V+ACxbRICWULmhe0GhIU48jJIe
PJQHh57AEqkDg71ALMz0Y8SjGi5fklp5gBYo/Vydmmci3PVqD7aczkc/aRXQnLJT
VOMNDM9dBoNZJXqFGIVubWZ0MWDW0rFGCogKU26npfflGrknKI9hiXX4CYKh2aif
9sQw51fpI2i10gxSZKilkObLbCH8tbrVS6gi7ObJ8wS7Fd/q9gO4MFCHhcqUNO73
PBQuF26dT4zM+xjd0KJlIqyjmNIawU0nYVhdsaw/FL0rChScCmIvB6EiN6bihTWF
98ryCLmUmGjegc7hA6eqZUW6ml46FXjxbnqUbMFrwaGY9zFIdMsgl4ZmvseywWwt
Nz3pbxSwuAOFN9xRraa6/24LkLj4BYAoMhK8kvL78/szdPDnPsBqHc9xzs7PJZku
8A/vXSA11R3SKkwu7mjI71AdSsc0iU5VSwUK+veYTppVVOJwKr+232ixovNqIlGb
0mQhR5RFG5Nd5H+qTuXgJr2PZjY/fA7ujoDzX7hs3QfwCUzoKgs1N8BgUuEXIxDV
BbjGUA9Wat7XK78OaeE95H2q4vzg1gAmju13dHWRK01o0+2qSbAzmE/ahprfa6Vz
gF1uk6IbQG8kawJwUmPMAVBjTbbkpgtd7+IyN1i00u4sqR1CMPFymJtH9Qk8uRBm
PCPFdBU5kqtIo4lPQj0aaFW+vP5g4TdW2oMR2g8mcOPUx3C/4495PGBwpyAjLsSM
+6VpkzDUEXE8ad9RGQXD7wcD0OGJL6tKQNyLH2dTbCpcMmfoa2wCL7lyF86Upluv
yENyRiWcCgumTUOSo32SwFpopjIkJZzjVy8lCQFqsMO0f3HcB2QcE8wCEkDk8Ee1
5VqSo21aImuoj+4EuiUYq7b/GXrMWPFcgfQQFiLzlhzltq9AJFAIMQMZV8GToxTL
4EL0mgjCJYN11DKiJWXqlZCCCAmSd8DFHvF9hNMAjll9vHdgvhTHDtloj0mKs1Ht
45NL1knc/hi2lLOWWfCUp8CRKBKLDRhmWC5KJLmQR1prDov+2AMa0ODI9mbwxq+h
xErd93B+4UcTR0uYoVr37kmZY6M+s4ahK5296QJlp8DpyrrfryRJCVm9UThaqVBU
zouxbPdib7DGvWmZMBgq85/nIuQF8W4d9DOSc776wmDIHq0gNdksGCzZpNykD6xw
yoB1ChonptezuTUjnFcvvoIWvCwS+zbPqhPGqQKf7jmAjKUFF4heuUiN9q2Pp2pF
839VzbokeoiYeBXP8iukITXC2yc1UNjpa/0VJ5mxHpP2n2z5n27HIs9AqWwXMEnN
7D0BoBMC8rJ05v4FnB0GGhFn+ReavacTHMnG+2VKpcbcnhLBJcP6C/YLHJ/L7dqr
tkodGA7q085L5zTnHbormX6aPjkn01OVYp5wlYWK3nHNdNbh76A7MZyNIrkf2Wpa
0g/YtWbYnZd4bahvlAikMoZ4xuHCBtAtlPoLCfpSA62Dk5adrEroMnoPzz+PQxAw
k12jtYbJJa93gahNJhMiaU+e/HAIBkRStNgGhT/Le3gHkr2DPoj07IC+ovcHkmMA
1CNaaKbvau/9eSPK8f2t9AzrW4ljMCdV/kEuCB/4/7goVDMj4IpflkZLBnDKkUqK
BSUjy0aCAd4e2duYsZyJ5McK94Wvu8U1eBLhAv71bxXL5rVFqlKCnvwWDWJvDiO5
vdHSlrNYdyEt2p8S5OCm+NbVyrjGiXlntlzINaoyC1wfHhIvFltfK4EuDhvejMPu
vg3Sl6O/ZpJmpaXIxv7V6uNP94V30pYwn346OucmkvChXAufnevMnlumHi9VdV1S
+63jLgAm2cQq8Vk35AoEH3y5KY5IZyO/pFaYjgO3F1/TEBF4V1Xco6PztFB7wkrr
fKVcB09HVDUb6vR7rPV7I8G8Hhdr6/pbjDBNNi836vVE6VDhvR0vEB9eDE7DeiAR
Mg21obMeKDgU81Dvh03LugBKCKJiwOEXMQLkY2YQ8TBieR2j91xd2XMr4dedS8ZJ
GMncm+X1nz2UYmtMtAeNUfQFKswIEdl8nLtpEfEXCSsK7kaCpWpIAg+mlRZR877n
IMXf5+IQHR3ccAvL0hCSRYPUh2AiSyqmKz3Pi/bt3R+I0MLKr8RsPQwL/cmOq+Es
2u+fQtHfX8QtuA1PqkzWxlwP0XCxjiJYkDzsU4c4gCXGXX0s7MSK+AaiZ6duuVJN
UdK0eG7+1HenNF+GrDuMGKC5lDIk8dg64UcEukcvLFZb+5X2clL5coDijfrp2vP6
SrsmuMkGSxpYUq5w2NnKDf/49fcgt/GqxuI74og8hFIxcLl64AldYOiYibEJwyYa
jyCGwWWvWacueF99ghtu5AtuxKLXm5p/cJKpapAtQhAMgiRWaj+XKZghKBFBnIv9
5+wlVX3qtZM3bS/zxG9mwk983leFI3d3LsE5m2ZD4bH5YqS5PCUHFNX89lIU90WF
FipGW6TFgnn9Zew3YHDmOI4xw3mJZEWikIF0pBpgJHwAulj8FZKK9apD0UIEf6qX
+N1L/uv0BJVIcgy8LUuVSD/48EqK8smg7NucjytMA3UmPok815WK0HumDsN+94vw
KcoAsKGOmisa9JxS37iCHBbvnglFNwDwHOuBAbjIeYNwGSWchpYShleXQSOGzW7h
sz8kMgxkxErhxY85SttyvKz+/8aphrKiwhWdUIvW8uUv0tA+LJeJIplhXS76YTnT
l10Lv2o7+k9OF1HwAy/swl0RHZRqnb3R6zAWx/U99ywK8coPMzPWTJ5TEAv+YinA
kqlTdAtKD2m5xZjtXgqDY7zlrDLOlqYjfTHtWfSuQDQG/koRZzn3u8/jLdFjpnNp
oCUOvELbueDcrMeUq2lsB1+Px4P/fBKkpwRFNNtNyoHbXCVfFpgfCFC/o6R6JFB5
e8m7+mpdvMULTkd9/yQsUwgVNpUtlf5WrhrCEX5OA4/SaXy50qtnMytBWNDOeTx5
etCxSGJFviR5veTV4cqwAvzxeSCuPzC9iC97ZaBahaM0VuF0P4agYJG2ZCPNE6hu
+mID6uuUGbO0h+HKhubRGE1qfbpoRSJrj171fZtv8AdwiAwE/026/8pJjcaZT8KB
huK62tVQ03uQ225n+zIj9b4X6qsjlRSvvS8gVr5P8b9BcgN534/c/ni6zt7EHId6
A/OHj/F3rtsjHxGhDd4xRhBpwbQWI1xBwY0qEcBgpa+gbKorMK8COLRdnBBjCRI4
zHFrLXku+52m5C1/pcZncT8Laq4yYzPGnVp3RktfoSgPGUVkFyDCK6ekD78QT4/J
/88323pHOAOsxerEHaH/MPcdbl08LOcjfKtXhiV/aklYroM9OGT4w4iDW6N3xXb+
pCpgLQgkR+sbX29sAOsXjQYgknlCh/g3D/8ag8bJLKHzHqXr9H1Zaf3YvmhdJODf
FG1T3SauntxlVdJUNTu5sXWLftmH4SfDSBI49mt3GRIFJK/ZAIE/LXtEutNV5vJm
O1ZXKBL1o35cGsubi3xBi+6kpxC99EwEjaGq+WjuYaw1AP6gq2iDrg3lnG4yUmF5
niQ9LfNlv7MML1uz1nCxpRVe8ckfkO5fkDvyVS8Mu/xUsAS7L0FHZX8lrR9TXxWH
MX/itLVgtZzvYdbsd9LKE14NIjHal4T/dCjILyH0DSt+/jtEpezoCfPqGPgjvNYT
ArpZsfHTFr0BnBdplEVTDtc3F3T4/Ze28oYubvwMMn9Ci6Ye0+O9Sz7lvQ85ZeZr
zXu3RD1qXbYXVgaAmk/acBZ+Y5souCYt6Ik5Wfhnw7O5FOc9Jgn6J/cKQ6JZ0ihG
PfLy7QYnZZtmf9CVttFA6xSLUK3x5eIDPPlxFi7UUVMcrC4+9OV/i4SdMJkdU3L5
WsTxHH1YdRJXFHCoAifXQ+SSr+Usr4doNIqDmovVemzbSU1toMwuurjq4E8PRig7
YupRb6L0KeDhwMhdruQ1jD9V6iVa3OxVgPTr+UF2+KYCKBoDuLVdP3tt8bTYmI2h
SVnKFEERd9j2oDWUn53nmaX5kOzb0ikHFbERsPFDTBJ5Q1qa0LnHnhir0BRXQafl
xSoFTRVidDI2Bx9e5DfZVrsj/oLixlQdLbn669efqi9GU8WdAVS5ueIjxPlFzYCS
Kt8oFmMNpQh1+F6dfzXu9xvBladt4vBZVB2hvasCKczlXcbzpN9wDqBOUVSyTNsD
MlUDeMDoZ/OrPhcPO0ROAE+UkRRR4OXs91nuMbQckHIlWMIqXwn68N409M51brKT
3ldHcbpVSOsm6Q441GaSy+52w7z9gkSiOsEI2q2fzqU782Dw8pNMQ9uxRJ1r5l4w
LBUuczLw4LzgMKsSPK3orfp8IZWoU1got+02hHzpbfySkHqlR9bIYfThAUmW9u7w
SfeOu/ldAoiCdN+fcsVPvoLc6o8eaGClLg+awHDKt8Jp/3/WpqTlDfgRamFaFHMI
2yZlzPv4PdtLfphRU/A2O7AmQi015QpzHF3BfQNmfUv4gm0w6Bc3leuKwmMpKnFo
jupoUUwxg8HuQzpEOm79kuL0cYK1O2Jr4GwPwwZfG7LmSdbL+9EtbD90GXlcbPM+
S8Y1U6M3+u+sLLPCa/D1aaRqUaoRccBOIaWkY8zZc8TfafwKaAd2UFGcF9h6KVf6
eSatN8k1uz0k/xBw6wbwIZqMX+6uR/J742rjuQF/fwCFS3f8Gr3R7OKJrBnTeI8j
xEIM3AyQaDVazm4ieC72P/mYfX381mHYSQdOiXrlh3A9bUQGM+xc7ysLjfM3tYi5
WJsTjvkHfj8r7zl/Tu4G17OmhGWF/F98+I1QitwaXN8w22UDK5rJqLtk388ouTub
YbE+/qJM91p6ESiim+8nFlJXvqi/yAXBb0bRS/c6+bP1N9juMBylUJXhplwWtCwJ
iZrusn6eS/caLZh6EJXoJghiFBQO1OOKeI+PurBe/MK/kBHd92qteU7RaJaRIC6x
oPVcV2+suOVurpps2rkPgZRibnZgY/qEou8lYxjnh3lCf4LH9unGJismfz/4ucDs
RCjxFqVvSYS5TA20l+tUUewrC5J7l5r93nFskmmYthEBNT0WHNw6A37il843j4DH
1L0WAqHATejY0cykUtz5xMd249JM+dldmErQGI/+ITAxlrnWlhkjiyvf5P2IvJZ9
JFj9sEW0a6R66PzsKAdYwWtEuzcQktup7FtT7evK2aao+QBxrN+HFOMoSAhcmFpA
yL2ZwYXZryB28bazkcLa1EsvN4uy6RZ95ecZjJjXUyJljkYJw4mG0ootdiHqWDOp
5fRPdPExU8y8VVZOULly9sEbLfstrXHasrLW4fmLNlrMAA7SmgtIs+WU+t1q0pEU
GqWbMRPawrBc58kzui2djtMrVwkUKj9D2iVscB/28l1Ju8PzySC4BXlx+8GrUql9
fD+Rqp4wGzdsebU9t7f2oJQILYxCAxmAb0fbhsRc6kSxMSiJzeAwbyZPqwxlmio3
f5+QUrHWcLh0NrX0b6AhfhItMCJYRG9pCNVhN1RMcaFdPm8CF/zUlskLPGdkSd2n
zjuKnP9ZocFZRpqsgrooAutpFCXLJpyda0ykmhaSDDCuHVqogfzhYww+5HbZ37ex
DrnnD6jJUneNK4sgxOLs8rNgScFJeZsLuSB1zqKXVeaOTfekGtmCHoB67NMuXgOh
8WLVC2HaZOtB8larno1dh8N9Y5TAMKOyC60RQjGAriMHMs8tK6qw6k2hsVPoQ1E8
wWdtArEZRRIzU9H/vGinC1MUNX/EpAZ5kjxeC4avdWiGP+6hfv9j+Ezksu84tswf
rm1kEo8KGQOerQU8i7ankie4D5TQPhRJ+/VxXJ6xNCseUXEayTbeMC1iyK7jmOTm
YB6Tn1uRGmAUtbApkzXYHW4GYsxtFdAa9YyJHzPS+Ghk4nC4iCHt8CCpKitGE56h
kKF/lKPJg+1I5W4rhkbCrCa2RnsVbk00XEUuPQk95QfRJxe3s8V/QYvzXrhPAZYm
5QTULjtHZKJva4omjiNoIQH6ZEyYTEX1LzsahA+a6+Q02lXbCIrMXXoqwYaznljJ
nqC7EPhRuJ5xV4SwB9GnxyTGf44MVqCV24ddNCN2THZSxXdDLW2s9l+AH6UjcOT+
i1f375fEP7x3RfvMRY+GcwQmpxKg25ILjWWfsKC6XHUEGvEBNsm9075klvOo6RKo
NMfcJcBEAsfVmaDjAWXHYcITeCu4YN3JrArROxjUQ60DEcNpeirJAEwYM83N74Ej
Es362ye7ahZuKEHWhBHVEcDaTT5/msXSpFn7s8RcpD84tPwoGcSNnvVFoCOVkEGe
N80gmd4/dNc2EfGqyRbmHdEcBo9HsVbpN3QAkA1y0TTVc5TEz+2WxbIy6Ff3mWnM
ppTwVquS1E9hD/YFO+31Rb4Oxi5eVcgjCpytmi4Bk/u+g3p2Sg0vh87WLsuhcIAo
j4zyS4t4rW7oWNcV920eGTTHyjWPxaMI1X25DzN5g/5iX3w3W7g8mJtOvCp3hVFl
Bc532qNNRGGO7J8Yl2YpSZCIhsbWLiZUvSmC41rNayMr6MCHSWcsbQIzJtPAtwzb
gxLcyJA3fTB2WDZsSJE16gLhs7fHEqMqWo5qKUZ374mZfcWHQ8DSBswuUOjMxgqz
2iqF56qKWL71Trywx0273idjg71U4Ilxme3T3zcP4TEnj58g8Qx2v8WFCpUIjcnL
yLvxQ904MjhdCWTTFA1D0wGMjcv4rWWbbRPNpDEO5+tyhVHdWS7+HycpBE1r2Ktz
jjOD5ZiiTYIUIrGF4U8eS7AK/QAspRzvELomEd3ZXpgGVhai92rl7cfCWNZbQcWJ
tGdBih865dGOFHAYLyJ+hGJn//h+HlPq5U49t+GggAKYzsjQktmE9UWFRI2cLgIO
aFNQ3AZxkYjluu4BAMADINCdWYBZnsIyqmsuDoJSr4eh6+JaXY0K3j6XMYUksOTd
DY5j1ip0GkbhDqKJXAYGwCwGq6UqGd8j0pCXxqX0x0O0TwS344NE75gckm1zFIDi
Ha0wbPsBcV/fOJ3CronN/JYfr0NxD0mNXty21vL51eUoprBVpB83QvzbPdMwPkY/
WQj6+mNUI5yQN/FbLLJN2a8S//090ZjvTtxV543ld0TNLg8aMLQ+zXyaTQpmW2cQ
QOQqR69kMgw46VIKpGVlCqalBWcjBj1RPiEiqygkH7KZZkfwDSjKzDDllv6p7nFs
UbNYAKaFu0S3nKn4iHu13yVYqqgCw4i3n0MXWZt8s/uNAQ6d/VryY8LLXUBxo1t4
8X5ymgqgbo4IR1sMPitw5xmlNfRcExpfScZkkpyOEMWOVK33z6aQacv3B4wWV6AH
i2T8u1uIBZlyiPI5lx1M9ZOjpJO7nIoSPzDlk2mF5z2MEyU14KL+/yBp6mr8DRM6
2DIteAP+9zki0RZCz9iIqplRxs/ECwIQQC7pnGsmf1fFAd4qIeXuUBtzlJWAlr8V
LA4oj843b/lUw1lAufnwoVc+mInYtg8LZ6uwVAg4/WBc6ciAGPFIU+AW19y/78UC
FC215EkQ79cm5NaMqIldw9f5TJbyV4f5hPrQ5ozh/ovryXmfaeEocno63f8GlNsA
vS54zdq9ZYuqsS9UtHlGf5z+0iTidmvkXNQ5ffGXHJAymE3Pa94CFC1tPO1f8LOF
dKW6Qh+PwYnPvXiXYlmVDIEZlg07mDEcEyyo/Prmkbc5Y1MdGB951d6swaWMlBFj
mO2mBNMOvwpD0CyKX3zl+7O4JaHeW+In0RoR9S7a4CX4PXvY8oyJn0jQK6o+In1d
kEK56RDvvh5v2SUfWNkMX1TRBLFkfGbo5HY4jCl/7x2pm43TBSzt8o6msFZsPS4f
ee789sd+SmqJnjlw/lp4eF8W5pMb6WstFq7S6Q6I/4kTPQm+FlU5jTdsWof6xpBp
aUA2jJAKPJQiJwxnwlbMsZixSXYnOW1ibKZQmardOolqACA185coSJQM2txuebcb
riFr9Dv5OtOTPkusG9WYTgtFyYMlxsgiThnD4lQPeDQFb11d4kn3r6RH588Z2kKK
jeeDv1p30xh8nTbCUJgXMDHEFe7VUkOVs0ag5z2pSMd0GFIMPkfa11duGH87NBs5
vgPnaCA7/voXVoMXgN59Xg5SI9i/77AKofoCD1I7Yo03GJUn8qOQQxPGdLQPWtEa
M0popuzH0dKrajmErj0xFpaICh0eWEXjcDqjGcldcmDhsIZyUdhNQNbCYiMqu9du
RFXO82yO7S+oVwimFL5AVwu4ncO6Yl4DUhxDogndVTXPgEiJJLl6+ECS3jKcgLIe
VRDmN1flr7Eq/hxl7QgYokdz4fiKG4zR9H+u7+g35nDzGvfDdCjBUcpji9lsr+fw
JD8w4+3dX+hft64YQIpoKrYW6Enowci2DLMLBukJJ/yFdrmK8uZbhEUTSNmhxSpv
yzILsBhy4hnOsvAgaG5yklBRzHh+/iF1o+EzbP+RzHnCfZmaM03kHMWVqaHjcFqt
HYbFg1QcLd57VnTyNaP3P4BE/UxXIjxvjw8iREKY0mEKfhoCrC3tx0pMw5zQ7ZB0
iY1ksJEXx8wxh4Ez9rRuTpO73lGnezz4GuNAgu+YnAnYzr2p+uNXRcu1Qloml70e
R/f4dBqIY3N9tk/xu0u4kgJXdc2FZgW2unvVUoV/6V8K62BWjXdVCiFrA1LLA65r
ts4YQf3o8sS8qwz35EX21yYqkFBgYuiEGv/2rIAgwKgUBSgvBa/6z0qucF8gqxAo
XRPXsyR9nNRI7Moa/QKqJ0afG8c8K0egXWJ/QOEoIffpKu4Aeb62nv8TyOz0SkPC
nzPp1tV2Ma9cNKOn8nwXfXZ/nUsNnfkX80VZVbnigBV+LdlyS1fGFev2GgC6WLlX
Q+6/DzhTbj1i4VB//Hx0BAz7biL0aZKDir/Gdmg9xudRbb4zmVpfEmkuI0Z07Pj2
F7jLVklgnts5fWr1Mb+3xVcUNISzUrOXJEBAmRvCxiufwAjXpKIPK5YfIM7zJ3Nx
4BH+tGf9hdsPSWX/3m90qyQ8Cv83/D7b5JSZKJavgT/O79fxQzit9DX/hQsQLTIb
8GiLYyzNI9fy/U0Lc0PObAM2eHT0Ma2KMk96Eq5GJ9S4z6E8fr2/4EQBxMNEmK6s
VqEctRvmY2x/ZH2onBSDAkMFUBrN6M+OQoCi45q173dECAKmmJ3JC8jMakAsEFXB
g95fe5mnt+bb8PTwIegKPxqiINSzePvbVKCfnqsdEBIiMo1WSRgI3CFLSBAHPeXn
JxbjVQUz/5OV+gBoDgPYmSgCY6k6jiLMIQV8S3kB2oWOgtNRTyMsHM9NI2Z7T4ia
0xUGodVX31mdIi8h7RBURd8U2MVpEQWCrOr2FQC9mfwmVa+E5+GbXpyU6V0XwN10
yWnxBgynHmjWOJKxBOkHvXMvEzzkxluT4cBrw1fa6Ig6IidRyqUASjTOTOEuop2Q
6hgNvHLaXiz0ycsHE6fFutf2ihCS49Y9uLsAJbQ3hD5rqFiEY+rVGpqCXQ8gyoZv
096CsYjslxaNzwM1G8ZLeZzwuWrh+LztJbcYb/USzxsdC0w0OraNH2tmGlRAt4TK
mB1WvPaOyV59fSC8hM37KHDVFcsI83CjOgVbwhKQGeWhbITjtTa4cemiSTEA06iW
U316dS+xaM/dOwr47i8TVi6nuyHhlzSHoAWGTXKvw6pXy09PTAIfiqWZKVdC19zI
JQLEZ0lPaUlbURceWRW/4SyCIAsElZ3TRMTNeHtRMOhwPzZiKAXPQ2zZsUI6dXo7
C38etQVfQk7NTsqbQcEErSOXzQJsbQcw7zSdRoVLJS4uvUvfi4ov5T+tneSVgIK2
wO/rxODJOEk2Mi1DsBqwDz1IcBQ8ibE5ZBP8rCS7+WaCSNYcwxG1289noj4sWHJY
RCvOTN4q506uoI7IoTnVYW6dTPR1DoVOgk/+NlRXpLbcpsDJLCYRzTEZYlGPzIfD
p+Tg7IZkkZX4RIIVtcRZg94mnmacAszdxpvB7DFLjoNjCMmDEwippauKGfgRwB6a
yCv1147MF+bh+RReJ++fQtzgB6k0HvK2usZzAXSWAsmetKYCMpR7IFE/d7ZYq2v4
5w33/9oJkaZ5qI3MHUCgUSo5soKx2Fr0hIwFakDL+GDnO5nFauMZD89vOl1Kb+Bg
m0DC/vmF3gKCGhTKQNoq0hlYMM7MWwuF6sh/rHeIwQAAMWsei0k8GF/6dVm6f1FL
igomrO7sZMO5H8rTpxLcnKdG6MbG22ric/aqtvb22j162sFlUfI95gYxzbD0J5IJ
AoRKs0W3IRYkBUPpHlapuP9E5LPcjoxMU1yQ0MDwX8mQWokpOUYqQMFp4H9CBe1J
Xs/uV7adHLYRaX2zim95JKXRZxLjjAeTtOvNqeM5+ZX45NgDJyZb9PDO0BS+Y+qD
RS+VX6TmAGSri6tDglBv+slpLed/Fpf9v5WBp0q1T2+2P1zRKG0Rqp1y9WGm2plm
7+xTmsXf6g2Tthf1b89wANCRDKHSyOuIGA4+Nc6AhZ7oASCOKGqPYzvtyuXgo2M+
ANqA5Hdau6IbakQLeGDYlk1l20CpYFYjLgMV7RZvZadYCGv17dFYFKah3KGr4k6c
Wy1p++UXvQu1GTulw8XLLd++WzuPjp2rGjR3MAXcAFC0gDPQGeBSMWAyPLYo+nGs
GToPwHg5sctxfrK6sk1r3VuOwUDkQoUdGm7HaFmnf1M2YRB/5vGGqwRaWySopD3D
KVE/xmDePUjXiGn+O7xCkUQeR8Woa3zwcGcDNKqBvNQh7uSzsbH2I22DeOigD54X
GylE6wCCUv58XLgwth079RPE4sqxoVOEmHi4x9zHqzJVqPEfzyEEJ7QRNjxItE1m
GJG+9mzugYvzmPgmc0R2ekFYaW7kLC2B7+q6MtMmux6IOUIIBzX3MbMUP97ZhORI
EgTm+4EO2ZJTqGjqBgy5gJSvwgzuR4GIMCiBGMGd+l2D5mIAFSmnQprQ1BwTT5vv
v6q9vOTIrSa9WYLkjbcs8HzBFGZUvjoAAZTD2C7xJ6hI0WBpw0uMKq7aaW0O1gHL
jIdBjHy1QOYBiH0uTf7IsGYZQKerDzn69IcNbPCaZ60KvCwcB7hjubAd/dtSkADA
G623MuSlwTa4Tsg4gxF0TvOE2MtNBiF27siwr/qAALA1n8zwCxtkAqJtNF8QHHUr
IFfoqxI7sk7c2Z6bRGeYBZo0SCRWRmJFcfW21UVvOtillJ69SlgFaI1Lxzms1SK3
oNRySU3fV/dyj3wleaIEiUeuura9xTgIRdPsgwzfSZQrjSVyOXfvIHk4ndVXtgb/
hKkMX1QQY18Gq7bINKt2o4xVacvokO5XBTUxwGBBHBI8xsIcOX3utfoGZX4E+C8u
GXLZt3NEnjlgaQSAM+5teFnMpOR2rKEegyGSNHlrlAsz7cjRvPQdr1RgaX7hxfEL
6uiaD+/178MLSPuHYThpUyZ4QjLWMASjCEDKj+CvDEsb1tqoHgXfMt9AD+pLWso+
paBfXe9ZY8QHm3miAeMXoR77PXtk3o9Jb7gWQodRNjTxSN38Dr8wyvcaBD4XsfdP
Jl2zcPjY/RCre/7nFqEey/rhfbtm4PFCO4x02HRLCwNSEdq1+//hnYOYtQPcudFr
bP2JlGiF3w4Z0QO2j8/gYvjsTbdyF4dc4FxwOuMbLewrhiYW2nCeP8drOwHdJMJs
4u96T7tbNpGyj8jCSm1XhW4Ls7BLueIOrApgbw1sDkWV+A6JxLqIEk1cEG1nDaDS
3XFUl6LSwbl3tLSsKlVkD+cbx8BcJzQ6jB8VThr1up87HM+vVJ1myLB1O4o6OBRU
uVLUuX7dQBfhOnSfnDCxzG/4YBDqRj6aOZY0MavYpuz+YIXg94QDwlDka2IQo2Zc
5fziAva3sYKxTk30ENp4SUTighN1o9w6B3RFgJhzTzmBbiJZLzMVNi9pjnN8Wm9w
Q2cmbSlQLu62MeFkqTZrmDdoYxFTLS2FKBnETUN1Q98JJQYOs9qVVmLH9wJom8Ln
y14t2/vfJ1wnua62D+AtmJi/IoYLXn+F0Y2EFRjLdJG6SiW+v+dmUZ0HF7DgWSas
F/uR/1WDAAyDuIrIAM70LueEDvUfY3QxXmmeEz5AHtlnOHuoMNTAxqATE0Hp/CFe
bIXKIm7qmlg4ad0VLxx7Y1iIKhcqsYLNJKU+UdwSgFkk3fO+7xB1x3yl8Zm7OwVb
qpxgR9XqMwE1tTeDBAPyvFBPSJ7d0XT6VtAtk3/zSVuOiNqz36X5t65NnmZbk3DV
z1KrtSTHa8soO+/Q34pwdCCHsG5M3DTxo4awIo26wPhbZ/pnfp02o8NoK84JH6G2
UpFBo2Dk3UVCnCKe8fhFvac5BwlLWbmZ8YJMAZ/6xTIhZk5m4IdV17CNtj6BSWo3
UEztwphkE7ctxwXkN5u12kXBp7cKvbjNxUp+PrT9k91qg1pMi4Vz3oyp6dLJf5RS
MSWLIgclltRoE4A/+kAQJVU3NSA5HtTWkkOeR+Tsrc6MXma4NC3UodHR0akBxXYl
SqFDJrwNfIyIgSWZRdYchkg6jM3n6n+YTIdPR+mUVumnNFHrrw9lw8r2B7jhVxxi
XEv7iWSrcpILJKfZiHX1c4QT+nQuQkIHDLBOo8eZEY/BgC2GFbSJ09NJsTwEEzRh
XiOMq6XY6GfrWyLI4+2eDDy8fzGo3FsFQVuWtRGyPCPGIR1+gpdpimRkyhSwBI1u
UN3+X0hUK+pXDvaKeYM5+Rv4lAzN8OA36KwvkAK1Inc+VrNpZIUiR6rSxvBlY2kd
voXzsSjgIKIURhUaz05WMZxHOme+ry3wxAVrSqVORFVSMOW9zEHKyePdNRD0Lduc
IqmrEyMpHrcFeZbZZxEZA1ogCi1As1MIgYI3Op0cwT7NSlcUJAsGFiLSSo4JRP9/
szYxt5hiBSMf4j8/cPgnzvce0U9YQchIyZGcH9XZBPbckmcBTy0Q423GcqB4WyPF
mIMBGbtUxpZx80/NQZ6eCIQfWsc8iq0OXi6Bue/lTVuZRNlW9zGNZbv3wMOHwc2m
WrJqoeGYrkLI+DWdt0w+Pkj5P4v8Vrpr7EA7qz/FMRYF1ZW8Fjo0tYVLPHmFJi+d
IU2SnIa+3LNVMYljnYF9F+hQhQIsY9IePhl8qyesUQtYQiYEcbzftde7NpRt3V2O
K9o//HZ0jC4u1e5dgFxb1lh8zorba0FDd3P1ZZR/ScPZGA7OglKftccbX0i/qGmC
yamYCTXvftrzcC7w7IdJPnpy6KkTp8DvIHo7ah8s2DZNAEJOQjimaOvmKh5QIais
O+ddZ4WRCciTjNgks6t9iaMVjCGMs7bwpyvo9mVznssFPjPROiG8yhShDMVMo1vK
mBvYZJ3HH7tsigm8ywXYMXg35zkWW9VEtEcm1rkhY9cK66ILM9hLx/6Vd7sjKBFT
vbmfmMgQxCAfglgZ2r8e4DEilg3jSmLchqBkd5cf19X7fxXFcxfIzprAQCrm65kY
8mdMt12diORBbmhBVdy8pOmpRvaYC4VU3hpY29Veege6DvNMNN5kqg46LJj9oubc
GaxfBXr2U9/plkzzfwEtA687GdlWXy2Rh0Ul4Qdsc0EwmeLyjIELBcmp33GlfWhc
ho/MP4ek6ZZUokfbWfboebcYQNFGOqoui5UArvDAO5IST1UJ+1vwmYAlex+eiZtC
d7NqWT2JyNzcHbfQn54RCloGI9Yaf0x72oSb5YRyosMlT0qvh+4IzO5j55nHzN5q
ALQ0wENUvw4h8wOTmsLjdTPdvk4crsJTvXbH4B7lwsUl+Weh0WJmxayeMVw5pTQj
5DQPL6QMVQGRQQ5JebjJqJUVB3YsIRWHzskSj+yLIbiJt3jLnxz1UOACsVLpf8gw
bRU59jjIGy4F7IeO3EtBI6vTGa/tnCq/SsCFf3djnitvdap25W1edNW0CqR5fhqm
W6abDCZepyzohkt0GMMpPTij0fyvru0BBN1PV81RkFWkeSCyssSGRqjEuLrNE763
pV4HJgu323mv21WuW5NEE634XYiVIEuLay8SdcmYxj0/1paR3IUlPpNBi7F7WFw1
Lz+/WQYWTWOvcCLAxdPayAIvyTkNgSnUbdMBkGmUo7Fd04UkZuZhtcauNz5fckMF
ouauP+UXt+T69GZ3bUXAcL5mN7G4MmTfkjXYeY8fTmyZS5u1SvNsvnzy8AveCm8X
1POx1p0g2tOTT+rW6fYVIXRsqdrM9e2KwtHbubvHIZpiT9yJfgoe6pNrIXlrHBRP
Vp2RV2sTmCGeaoQqPWOqKq9vo7+lfZf2LkC8ZZcGcHMpQ/jDL8MmzHDvpbk0RsX5
A3Kb6vpGvfElhpAW3dNnfLoTdn7JDaWw9aMfpyXa/ZHC8FK4QJ4yV41i88xYtNaw
V6awgjJtocr3JjWm2enXOa7GTfyQ0tSGs7rHpH59MVG6o8BagH8eiT/61ggHdJRX
cMe573l4WOJy9HIq3j9QJmcfmmggYzOfLZbdxyru6cF7bD7bfuyUcOj1o2Ci0K0l
fWp9twErzBwTcAz7EmV5VoralyhvveXb+SwYC2awUsqJJ05WIQWUuzaQrpKYFfl1
cUfP+LDU/ZFpRq+xecDDTZaQjXlCSLICQIsJhVGwQ9/CYqxr3oMkyFclyofa29yC
eTkaawL52ZZo6SDO9AM0pKXCvvYlbbZ0jVtVKMFIE4lJiLkX/sVEyiPgEqlh64UA
CEI0sZp2wxqufJh0ze5pkb2ga5CkvVkOIkS+rOidDXImE4+fBr6vaGoxwjYVrVOc
UCxrcC/E2t39kQk9agCZsY4vXbdO++T74JfkogazswJinPrkxFV6vROHD1D/Hlvw
/YECiXQ4R9bMT0iFkeT4ILfoBUG32i/smLZgo0VC3eawx8XjiaGU2WFbqvmNJz2x
424lo79M7Hksszstc7XI8nixpmjsKt03g/uQ1w6tdcchl7g7zzNpPxdwmBkhDOMe
Mcc6jxzVuEC6brqNnn6O7vszdwua2Obfqkz8vr1rnko/sDHY6JbJNjOCzGQjm0vx
TX5Cw8RRak2WcQIjXj3cWxx2eAZrXe09tKAAFiRcpCCuA3+YRWfRnY3QdSsyz6aQ
Y+81Qz+xonBHhPYOpAd10jSgHd3jtrZrb3Da0kav2igcubzQ9IZf7ApEX2tb8IkH
HptuE31OG2Sn3J9YV+RTUYI1ZpUpCgZohJM8voHNKvfqFvo87tcenuzPcBku9Csu
euSUsw6bx3Acx+A9729dPOc9P9jvQcuvDHy875IweT2p055nBUplewc9r6knCVLG
YkUoaEPnBnfDyTe8axv6NdBy9E9pCIgCR1FXZSg9YVZL4cW2Ouhb/xt2+R03RUm/
N9FUKbcAfwX7pBEe5iJ4aXKT6Fol8WG1AaLzA9y0vxyGdTsOLpkDPoU448lEmYWD
w5hPDFDew73a2bY/ScX35m0gr3inH1TKuuf6Ar/8aDKRx9maVu6WTEEBqdm+gJKi
QzzXQ5ZjZSuCCd9/OFkHNyCdES4p97AhPrrdSwSs326RgTGEQDum8EMOs0V7JBR0
XvCatE9X/Gmc44b0WmnDE3Ezasqvrl+I2WUFaMedzH60i/3aW+axUxiydk4g2x9J
vHLvfaHlhrF2kHH6to9TnHBeS7YgoB7dU57sRuD8osZCVHX+f0/KEQh9VQdhgSa0
a4mekt0J325IxQV34Coa9Opc9YO7P4Cm0KYgrs5S0Rv+inZsxBxJBW71xVQkk1Ud
XJX2fkZqg4ml8RsHsbo1vCPFRsie5zBPGsdDmOJ6PQEQ/Aypsh2oI5gWTgqDl3xX
mrDNrvVFWugswBoRhbJs9F9CerTlKQxTSRmQx9s+W7SMZCgqolZP7wkWiRoWd4Hq
gPUP6EU2kqQxejVe/Qw/xWy6BKxJ3NcJ/FiJLDjIEHX+E70pviCX6ITROZWvEoIN
Bs5DQNhucUelKkMabcfa476Bl/ePnFFEIZ+HEiOy2PmOP93yw2lDK0SDj/F6Np6g
ULsnUw66wiCPBeNq8tdv7sfDsWcuEvAlYPJizwG/LuMrR4bGLvyiiJ+DFjFQPDV8
qZOk6pF6OpwjwpwTZCefZZnARYdTmkW6uTaXg4n7IUzBQIA1zOmee97dDJ+Qa6vI
hZJbddQj938gOBWgY4i2Cx0k+44J2sJoa1ZuRAhuV7zuxQGDLLznNKYipaZugQo1
/enuiw32UfjdJo6T220n6FbHJ1aZsvabovl6X8Qzi1HOisxQ7U1jgxYthpOrHN0f
oWN/EhO4CZKUfDtyhRbiK7EySaqMX3IRDiIgJZpcWrxpXxfNiZ4oa2VSxJpRQpDx
2OGqjNys5GIvjf7LhvbigSJsAErJ/zQw9+Ec9izmEECi05qIhL5am9BKc+gUKyZ2
p56946UgYRoaJWDQDSqO2xQQoCuyFB/SGucNZArT5VVwPZaTg2cHfRTBMrhInEu9
U/zYDcPo6nVs3bp2OCJrBuyEQR5U3bkcxh8NOQXyQNUAz6TSS/FSi538btEA8T37
QDqcAOmHvvf0xWc4XxkCosvdrQsB+pGaItEKSw2vOUnrVYyjzzQFW8O0wNzXeEsI
wLWQTfzGcJfU5ipHxVosh8y7QDK5g2390AO/QXXTuoQqz2BoJtnTbpgL3Nd+wI8W
Cy07tzaTT18Wduze1RgIl0yp3Zh1TTVGKcpAHqS+410gXLIEh9rG7GAGLNz71mxG
tKujLSWsVM8pa+su7ercs5ufwsBykNkhNWy6N8lzgeyKKMG7sg5creDyWmb5d4zJ
W1d3hC094HZEG/9rkM+k5INUMkjkFlXdlGvJj/ZNw1f6fg3eMKFGBaH0hFTfYy7H
OC7yVh6s0bksmlzn2pBlG2Ml5ajyVJA7Fx7WrP8OuxaeTM1iFtv+41pX2wDsfRX+
Um/atnoryjL3k+8crAQlTpzSCIzxI5v39bZiarmiWAOin951q/KuRSHgORikkqTe
rX3YNoXRqfPeyWQ1bK57IbiTwzHFAC7QnpvKeEl3etS12KpV/OuWKyejRw5JPGdX
tULb3c3ki7gfK/sglPeSUgJLnkh8QktDTishKpTafHVww3V5ltly46VUO1aQMceT
ovlRRHhDdmHENI6KaPndtDwvA3xpTH+YPumIzFkf633ZWKMfqCruqEhH7qve2xEk
N+aO/8yAW+vuKCCNZQ7tuWKyWfBB2ZRYxfpKIdLlF9d6/3mLeuLp3sD6vZHi6FSf
F2KUpSA9gDN0JaJTmg7C2f276rZ0CK4oI5Db1OUvkiTUMWS7kyaamZK2e7xkRWz7
bhS//eQ7eli1rRvPaLm+W3TJcdNl3Z4o6bcB1TYfE18cBulbqrfcQyiIljKWBnps
Wq9aqSDUjW0BRsdtFVFOQwR+I7nrNYkJnwPI5Iv/da07RySGus0u7lZOLSDAFFdI
UksFxR4O9rmFQVHGwjOxIU2vjSEQOSMFY+XgFregPZmyRZF7b050QakjWzZR0OkO
xe3zdKU+h/8Dlg2f4tQCv9j2at8GIr0aZ5V6LS3NNihIKPzndpQNmx75XkokuPk3
fe427fhRtUlaRxhCyYm6P67cISut/YAeQinAM7w8ns2X4vcRQabbWc0KoK7IXzvW
QyoF4EJPUOGfETMjJX+c3eszbxwh49wMr+iMm8o/p6ZCfbcLAZAwUiNnmUjZi27J
I8CXUAVdV4rmJhDwWgIl1p3hq/ug3iid1pZZhHRLUfNp60VMF6ejLRO/TyVYct99
JaOhi7nmnDsX20B2oC2G+eYFAmUT99M0zvyZBafwW2Zu/E7Zj51KXjPV9PXZR8CK
33mrQQWsI4MNPo8jaSySJ5s3hD/LItWlTBGVZ1jig+W/rjiBTHbrbzOWNT9j8jTH
2GhRmEkFsY1zHKtmgXMUR4JisBE4x5v3hPGVc/SnplPrpU1JTC26sIcSATG6dNmY
2tl9UngjYPlxVYyQWwJBNDnt1LpVHYc3C5fWeGOHhL2CQwD0T4O4h22nR1oSCBL1
tU5JT8qTBQ77syfj9JoDPzEF+fyWCu4v3N/7zMZydLGErJdEg0a13fz3PUHWGkGY
TkVu/lII3QW8UfmLKgPU1tSJTOusCezEhvSJEn78K3VC5gylLqEYi2eM1dcY4TSQ
7qAhqvS+pCzZ2PJu+Hnzh1DOgjpazzJbPCDElO2SlyOEVOlhHuzChEYa7mEpX9un
oXfM1kIRwqin9ltYYDi/ksGTOkD6yfDbH8su5iZkJpjfRGDdyisMeaConj8JFK/t
dGIS+n7WUkVetKcAtWy4j0llk7/NMDNfNQY/O8556I5UP3RBvexmxHrhX+9HANsJ
rmAH1JBYgORy+LPj1CnwQqlgmPFhLV6wgOw2sthGUyIg6Hcs29vkbsPFCbD5mQHk
amDyPHpcBwRlIYonvFoAN1NLwGg7pBr6i8wZMssprfCHw5Domt2EPSWspReSc+it
5oJiZRSwX8klLO4OsRnqblBsA+haiw9jcx0NzjIYNGnQMiFcvKpBP/zC9fLSpngX
2ZDfDHA9uXTR8VHgXxBeaSThPbrFcNNhXp3kHMZ8SXBCA3NRpXiy371dE08DetED
2fO08daI6YhwUQqf2TcH0aTaKUKE0duaSXLi5VpxwzKXvH6lzoD2Y9NZWQtA2gYV
Fiq6omV7vc0K+4BaBJq12TiXSaj8ET13JFsAL54I1sQjhJejB5yKlr55/HaAAzp+
hrxfowYBoFO1M9ANkjOClBh+6E2i+yMs6OiyEw216AbpI28yV8IeOecEdHKXBNUf
saem5yPK7qZpOriiuLvwAZ7/OTNRVtP5G2hmf9IUDuSlPhI0sEp5E5xg2Bm5hshr
EWiw7kDCQAybpUh6eLhOiMQRWJv8OsPjvzjar6In2fF9PJlupaylCHskG812tIB6
zr0uSnK20N11cs+2epOU13f6nY5F79g7WaDYcKwPPYrJ4+9rSWAet250Hx2p4Sal
SNYnxtog+sxKVuAKbDM4eZhGdM0R6PSffTfFu0SXrV+urmYuGp0pLVX0R23LyXXZ
BJ50B4yMXhvhjSQantlKkgcAvnCJjf8s9uhjH4a/oRuu6kJKCU+aMEFkk2Y6WvhR
N39ozjspjGokbvxTtx08TuiOELN3d81GdvkNe0XHYbrwRIkKtFiS0ajHXi3kDlel
jmq2XKfG9zYYWyi7EIRcYCjmpKsmWmFZ0it+rikemqcA1mTzQs/dp+0ef2I0bUj7
0XyJo0fvqCqB0CXzYIdX/F7eTaJICCS7p8S4DiXbzgCmSdJ2q2b0jZWOu2c4taJG
oDqsI4R2xRfUyDdygdzccfmXiT1BkdQtq4pLaMZplIZQYaESaE5NeNAnoG1hzYQC
Qmz9BC8OA15g0jJREfIDtL21RNbXnb0EhgPuB2bL4/p52EgNJNUV0djs6BPaqobb
Qzzj/41CcdI3NIJmwnrQEteT2ieTaP4427p5A4nWAkDKo9amFsL6H7FdOUR5cX7d
NGdUlgvBebT2P8BWAT9872a0X18ZVqji3jbR/pC3966ivdB3bAz1fVtsieq2R1bP
LejJEv0iWdtU4Kyb7IItZv3gZawBbH09Pb4n3cGw41gW5JdEzI8UugMXquuuMVR/
V0N3eMDpYJrbKmOzK+Q4V3qeGoIFFNxAG8dcy4EP4ivjUMLdZ3lJ4M35d2/QDQq6
YTV4JcCwy06NlhWYv0eU5T5IBmeczRDK8+vnvGjv6Z+jW2pMxiQf/7NfyvE4MyNB
nL4HK0DMfpisvMmnskp4xyIEH2BGpRmqaWBLhFg0xK8sJOhNBftdbrlp5j5l2SKu
YGooisibkk/EyULBITeKRhX+25pcPOh8RcwVPiX0B4sHdlBqZErZPWRr+sMIbfbg
sNLsLBLse+RJWPdnqvJNLdG4Ztn4BHrL0+fSk8TlFBI7NH3p/iAhDvvAU5r6VMZ6
4AfbvWvrdvxvQK6BRMADq+RewqXYMlv0chaaK+M2ye0NejQeUPuzTyLnj37gsaiR
+4JWrRXPh7St4b/M5uqz/HEIvBXgjvWp0H8NMp5Gt2THfq+qzhbSbyuBe9mBtufW
HW6NDG+FwSTG/azSA25rS2GYvmOpS2zLMMbbA6warTSQVm41MY4Wj6Ih79DeftLb
0p2uETMY6jsJQyNkzNHt37hmRlHZGoD6d62u7GHjY57VezCiruJxapOkZ40qj51j
SNmm/8zFTz+BULZhSh6sllbuoNMDYPXCzHnI7Dv4ufnwx+ysOETZQMSzZzPI+ILA
sJmrE3896dXpdAxhhj7AE48QJaiuF2SXi6QHkt6aZbdHeMsTasF+PIhWOnCYcFAO
7BLtErPq3vO5HLr0nA4astXzEKomTo4c0Ppt6G0SVnJeV9/hRsUh0nV+g8vQi1Pe
O9DG0TUsDPHm1v4pYQ4PJBq3s6aamqSVs8JP/wr9znJBn1HjUpyX6uLQnGHJ3e8D
pTVqjq/DtSpZE0xIVCW39+AJONG8cLcZdD2cPrBbkrgPadcyyRbk/QCVXz176s5F
5tME2zhZRnWQo7mTkiJsUFGqErykb4GRqdAgLIdCLM5fHqewQ+UeC4YQlMfrtfzV
SQrSr8Jzl6TscqKmm7gwZWOsyq4RAKvjhiwH4TMD8qtmA3sWXXaa8vCvYxuRlKiC
t/PsK6BcpxxIEMXtHB7X0NdyMcjDte5y+r/IOIHAm7ujwZ1QpbLUKlD7Dh90YY55
o92l2EHQi+DFFc0SSxB7VK+rZ9Ixhi4aymWj8QyHuzMxtje/AqHhqPNBKtqD7cTV
Q3hu7V+byN189qldIvzh9rVQfD9oEhD5OJmlPIN/xWgXj+M06FkwrjJ7dnqNkSDy
drQlZODPhDID9fVtRHLsztn9vvSMwGTDhAQdIcDM8Mutijv/uzm6b2uUBDgGqkXd
XxzDRVIiYFUU+9dk87MVwg41azPhGupP6zHteHSgCSd9bcjmRI0BO+zoet5Fq7Vh
aklEefA96R+iaY76Ry3FqvFTB80SKeMZJaisHPHh6qXqr9smEtd/EaP7llpwhgei
UJjCwqCcbSa8RzcaeJ/IWrxrn8v2mjBeLoND5BPlKZo9gz8BPH2gF4MF50qoRtaK
IKRPbMdpKborcMvNwoGfOioQCduMLYJKmox7ChPNSEc30o+YxlkSQpkYmfTR79Hk
ZL5BOYRg+uk/d7tmtb31vUKoKE/oploRwdz8V+iqLRBddK2Qh6ku00iAzfW1uBWI
bUMb2vX6cRoWYh4y7JUjWxpEkCWPeqqzin0Rz9dGamq1NnKHpdKobBr+EV2l52pI
tOP+dVHBJXMJ+C/kwQlAZm6zm/b5jl2rHoEKM66WQd1pkWlm84GozcvSwyBcDy1+
4W6PAHNKsYeMyxqYkkwcgjcdqkiydcVdA76GbCkh6pRFmF87omOYwLjjt2pJHSnw
XE7NtPaXloeifW2ER/u+WhfA0U/ibwWiezLo/6lpS8BNKO3ciLVSeuQGAKJTv52H
vVn/djXhU3AptTc2G4+SJBkcC+ZmHlaRgSVVLQekeiBb/6TU9fVmnw7pGCqtKfNJ
Frzygb+N/akFLw8rdy5xFOmdeN59b2FcskespT60wSNl9J7b/bEqEwwsOimR/PA5
agi0OMbJJph6MkfMuJOgOJONUZbC3fwWIPRdLq7PLo0XIQUvtXS1uA28NqmqcrzI
8ER3WFkgBiCmExPll1WGjNYJGGNbFuvHuhkYVxMmOCPCYbFZR7zwav/qYFbc4lm4
MR7VFdBbU3smZe0VPs22gv+11YcEj5/DEUYrdFm7htNeH/DIRtTdhkhG2ttNJzQi
RSC6uH1gC2h1xmYjeugklC/FvJPWRcOcK7lOeLphKTDzH0vRp31T7t+0ZutI+1Si
/qjUnbKRO1qqi70+zgTmodj9WktCbVsSxXSTaeUEHnrNmGWfSakGT30KY/ANi8Id
XWL0SYa6BGiSYJVfR/6kRmp2fRXF1DRlNFOwI1WSQyO+vNmQPp0GPiTf2i1Q1LYp
GKfS8CnzlvgabiqoFHOAKFy4BsEiCv6EaQ97c43WEF+G5T9S30i1+4bnYPdO0GYW
y2mDMRl2iqPQkZ/s+RBGS86qBbsR4NfgjqPwF4sBWasPf5cCk+MhvTaaJyWu1ood
1sRJ0BY3Xm5VNi4+ZD7DIA5MwqHa30cIWDbP0V0WhIHG2U7+x/ZukMbsM+rnU0NX
3PK9puOV+MMtkIV4qJMaCIBhtX/ChKSieBrEwK5at0xGcBRMUTDxp+iLZvOUjDoi
1QK5VRnFigjPzXuFsGEnn3Ut57m7AYxE/VQmS9WJRrGVWUEO7tteyX03vdjnFNLs
VNLB8zcCLY2B7cmLKjC+DvcuE526qvnEnZ2S1UWZ2c1vqqOfxpXR8yr9avYAKYVA
tJyZIiJApmnfbzRatgSQI/g7x+N0uTH9nJaX/gtG+XBcXZR8RQxVrYCxeDNLwvQV
+prAULWCbmhkf2VDVKxobMH64uDnJxD6UJ9roTun0qdRqfE2E/1qn5N7Mp1ue4wk
Xk0jH2Ix0J6nRLYhmjqALwWKF7UTPOOcZRAfDch9y+tsz6LsMRKRvww55FV6MZ5Y
tvqlGiqhFq9MxChM0cpRdNJcz19Ol7NfaZyspdBY7fPWQFRUt+r5+U/MZGcqCC6q
xeEx1xDqskzKh+76D7i8E6PZJU7MpFUdvkSm5Iy88HEvL3XYqhlW7xA5V/udI5Ua
SgiUP4EoqYW5rQ1heuNjTbHUlEk6UgMQH5zhxN2bpvtjuuaNznE4VGCYVcZcnDN/
2caSmoVa6AmSMQztU5b2rtF0q/jPkBWS3M1lNie5MOI1Uqh/ltrEMhGtA6sE66t/
gmY0GDxx5tvYKQt1syeeELboi48t9LmDiLQZEXjV7Gie5dQypo8iCodJqaYclRmu
bEXoOai8L01w/EZKrkQoOHj0GAv0YWrkY9AHGJHMr/v5vgnchIB1l9Nr5JK76Dr0
BdDZ0YIYCPXJTOzvA0SFRHNJyrVkp99KmauntYRo65iMumcRbZSytNxyrUcEXHhe
oBdMHHjpy/AOX24wZLJJxahUuv36CxqLaQ56r/urG+YuHneFZY/46TC6pmvhwmyS
WWhZsqNSGXOzcFLbe+T2LyL6qgThLRd6R/vn6AWecxAtD7JcH6GzkMy/mNNOc2CN
66jABdEGG1H1Jv4e8FMFfvwogyMPsvOSqDS/mV5wNd7vUxM4I/7ffTPgoJVLiUdW
Epq2fZimBG6gDY2Hx8Xknn6jxAtpFGsnPcJMfEOolqPXnesqzcRTSjua/oMEQ5YP
mAs2sp2i/PYY3oDWPq8w/GrQ4NQUIwgMwnXfsTrq/HjS+8zqdXeAsp+2FZJ87zuh
cua6rNAbgrKDjfUORQ5p5J7zGasWpvOmsU8Au/38MY5Tb2wV7OA0CBRRsL27hb6U
t/qA/Jh65tYNSFJMo11KAsE5Nnz8rt1QybVqyJj8ZHPyZeiK/m9ZqmxGv4CCoP2L
MvcOmme4f5DJ1VymcL3hvI5z4k4G+zUOtSIqloI2rPL1fQYTb4gthzc02X39YXff
FwvlVE79iOu/5FSzn1cQ7EJFKS36CgQr0Kmg1Tvx7dzPGSbjOCums9e6+4b2GQAt
YOeiLiB8VKiAqIvHCBIQ13ywxKfJjv1uaonRj+qcJfkvhQXyM3Mhj/GVz8Ji023+
ruWkUDRiMEvBLIhXBwZQ8kqEs4myzcIsIpG8XgYt8Qlw/PZExhEYXd4Lv2J/6AaK
JMG1DWrUlllV9pOdEck40GWJmS4FKFSSWSZ0P7rWwAZENVgiFpEOy1Agd9INmzC/
QCPMHhICJY8uiNeq9ueezxBgOVLBx84tm2JYvHVTFgwzG+8DUhpwEqcd8hSaeIYc
SpFZkDAUvNryuNRg5OX7O/+X6zBeStbhF9SGrweGmUBgnNJ7NVRedYbJKTkm4QjB
9XWF7EtZuJBphroMGGkRmyKf6KgYK3VQFNsKLffiPq1x/pbqw8R2h3vJOz1c+BA8
a+n/OuLfrnp+ezD/RVBBA2l5kdtJgtJGuoe2kdZiChEm/JdB/3ibnitM/GiJRdxZ
6Dz2itGStxk5hojG4aklUcDV3qoesFW7k3FKGVeLc0p1DPRJyB8XUxYjLQVNpW51
FakD9nOOcUv4+8KlkqVRUkaypzTkJPMb3xyCkHoI1IKKeWYV9xXgZLVZ1mvHXhI3
SW+y7R4VYkgMfiFH4Vb3klUY03Ke6+RJQV91Ow/6VewzHZCjZIB9FRS1ZXAj0T0o
oLuKfSQPNuXZbkzirvBtvVQtvGPAtjB3MP7ZRiHrJsQtBNYMu0ga20zgyYvylfCw
DKlFidslEOfp4qa+3kgiWkYs5UtPmYp87H64sVGgziSbVhq8GT1tx4+XGuLfFO7y
whoMucUQh5+FYmsEIjd7zJ4K7k12pkIb9F7IwhfEYoYrLf6lH9ng2Ean2VDZcEnZ
RtGkGduir3+urIp0CDOFdLaRAVwFqqAiZUUdGhIKtBSuFGtemRH09FUolYvKL+p6
Zt/6Gn1GIFjoyI8IrH92K8v8iuWrp5qkSzULWi/kpXTgS4D/xHs6UCAd+NRA0NZP
OJi20rIgBv+YuSquPhHky6+v2X+APP3XY+auIdZmMaYARSHxH0Y0LJRVCOPmMbwc
ATh+RmEpxs4mhXomnPh3VneiJQKj09Nf7BfWNAw3txIfZAvrvr6Mmn6NMwFoLaeb
O/1dQsPM9Bm2h5VoFLC+eNzuA7g5gikHnpi+amiBDvBLo++3eGKh64yOX/FTi+gO
FivycOkNH8cA9ZoQaq2MRKgxzUBN1W7IevLzlBRn2f7BBaw/Otkdko20p/aoMA+o
T9ARGpxAVbYL8HKLqU+aVzXybgvofTN6gU/KMie1r7t3XLaZ7pxbaDyrbAuLPcej
+0EvEsFrmyfHGoj1eLrBbc7XxSA8LGynSL0rOPbf86hD6dxHiNGje1QcaS8ylBqv
X++dwjJW4qqHhgj/F8kP7x0kL3TlJwes9er7ifVn/IVyXxjkxU6dDcv+2nezX/oi
LNt8UOE8/QHo/fm6kCWZn2Rr9OOH+GTVxe01DEbJpGa3vUuRnzUSLT0/U0R/jigb
jSkRiOt4ShiNpTPSkyaBPU91Z2qZ0u0AgJPgd9g1dmAoi8VOZraS3WtTRMIss15W
aI4HUNnFQd4XAwix1qDwrRNM7INiryEMxqZX0Duis6nvTsqkXMp/HDslKb35jCV7
tPKeuB1Ar49THJMoiUSQtx2922Wurps9XOWorlD55UrTaUOJP75XyGTDbyLbgizD
32kf8CgBrb38+y9FDyZI5WuYmljK3r9QcKN+mKc6Icnc7D9RR7N+xdwPlIXHcPUn
TLkTxrX/jThrRA8Ne3KoASWyCymoEQz/fgU6MtWDKGtFyDYoXhuK+tqWCJXgveOB
h/pOuEX12hk9JG8cFEdy86RClhUbnJtxawKDu9UkegDePwpWRItQVdBvHuaxbUOE
qUQSw7fv/7HCESrqwSQK6430pmT9iDbBPVvNnRCbzqSbX10EObc87/ja6HMvOIvV
qmt+5bSjn3M5cPPipSveb2mBywccv1hM0PsDAb6+sGWIE96Tc2i9PsCWFFZNK0RW
pNaMpXNPgo78ULRP1oj/V1AUz3WhFB3AqSapBe9ggKHXx+5OAreTs9Fdgsq01Epa
kcHAabSyzbnCKCjUWyUfwNQhgKfN+Avysjj17fOQXyqz2b214FryST6qYpmxAnrV
fV7DtseWp81NIeo3gM7+ikVkKk74Xg/tiOkGaTgsAo39mK+3rN//2NDpjBeaXVnk
VPNTIZow4MuBW3ImJGJ8zwKiq0JcgL++LnPi4daOV6vVV8EItWp2TKJIdswVTCPJ
5bGzNFVmc709QB+eI/rmNp4ngswy3ezr3eS4a3VLIeu3pLelQihUropLrO2X9IXd
8rBYke8HFmEqP+LYbi7LdJCscWpMqZCMHNJlsUQpxkFAk6TuAxx8imofVdukHZg4
vQ1AMtDjUpO7u5NPPLEtDYbELgA3sHERg8/2wcjzJ5b2Lwo5bhAJbusD/Is4qG6P
7xp28HSXzyuRHtkpnMFQWmUFiObXHvEqJgmG+PeD6XlSry56DeUkuhht1S6PxDMg
pmrT8TKwX1Ufx+9KvIUA64nyapoh6Z7nNULhRVIpEpbGFBRmUiumCcTy4UKZ45QR
5cpNZfZn6achrKxSaLFR8qHUv6gXMuaVv+3Qt0LYmP9Kt6mR41BYK3xUlhbCdGc5
KqIHF53fu8flzZYlhPzj4XRLjr3cREWYHuDZCxH7e3tAiTkNJQAPmVXQTqUaETAI
QTHHul43ufKjCv8U83YF6VQ5j4LKPutv3vl1D8g3lRSjgV3aq92UyvxAS92ecxy8
j6os+87R24Y9VSjLju5gadgrWxZynDCDI/nBXwrt/5pWrarvRJNspYXnMIMtaiHq
nc5vf+vd1roF2sPkZfaCWs1wjRIc11Gpm3LbJCEG2YEsGdC6QOB6+nh08jICOzMt
lH3jtvTHnVk9dqS2GNeCPm5gICMKm9vZEL+Ks2wxC0h5qgH34KfXfNpgbNOLPkJq
E0u9a6Elli0JO3DhmW0c4Q9rhNk0aDSEB4EkeXqmFTQhzP5Ex4EzbXAkZXnbWArH
00R6/T1GrnsKTZETJCAFecWqELFManBczMfGHLZO6p56+wlYTP/lCTZftbo6Iy1c
qrZ6Mzv3zA4mob4Pr8p5wipo++jpgl2bn4qwq4EMq6V2EaOKdqzYLUR6/4M8jYy7
di1nGOo4pJ+yKX2WIQyUcYJZDQ2TMlWvvulWoUQ3KnBwBuMygPfFkTC78Mp2Tx/Y
6MnNWy/MAZG4AbIdPXS6+MAirrA7sdVJqremgJnD8CeFMdN5wx9jSnwj094jPnbX
l7BLZahoVOhTHQCrdgGgiYBtuFEfLYwpWSQIWeVw+RjSnQn3mxMcQP4G+L91gZC3
qGcqLuPYYmxMKtz+UTSTnKihOZhg8WbArlAEpMDrNq/zOJjeErGbZuT1GirREewP
14PiQfyYJcachFpwUkOOZYGNw9QnGXBFTvxTd6vEWYctKbWDfZDORnY0uhjSpkim
5EjagiA4Watb1py5bgWBXvjyUq9tx+UqaarB+RcSV+el8ZPRjjbN3/qTyfl9fv8i
pUnAwzP9VpFQJyNsOxTafODKd5oScE0BlfwHb5ERR/Qn4oT/oY97U8i6zTM8XrXg
cRly/gUepEX5HHUm9A9/gV3SIsQN3RLPyQsXsib9mzvwYLH4jVnMYHqtf1I0SeI0
+7Rt23fGfTnZyAf0AbO9qYlsjjynCCsboLX/mBl5j5GMjM9nrbKiLjNsCXqrIyEY
2WBi0rdtMjZ+irUU0lRXm8gy550OnIQ7AlNhxzGZl5V2dB+yh5gd/49CrjP1Tnbn
TTTunPNjEwJ910yBLfM3bqJmtYriglF0cujLICWgOndajM584MS2wFHrovUJHQaU
pjDn6SCnI8E/OhUf5W8eDsPQl3UdbLtKuBOkSkFloS2/xxk7QZW0XDqC/wkVZXj/
DvGtTj7AZdlWxW5izn0g1dABe9tfiR3+2qGPRkzD5LWpRFbDemTnaegfpuTSkgM3
i7I2Ei5W+DdbSz3sfrUa+moXTISHyg2uVCGhOOueLlH9/p165HU20cdLs/fO+bSV
WY0xIkJXlz+w/lIYbAaKRUlwSpYPxoANlGG7nGGT7e6xuA8oHsKg1TtY/9UKEv9x
IV5FOLe2D+yUiFSsmAyZPeqputfqL31JnkZfFy/qVaYk+2MHGY/mz3PHYa5lDmpo
cIFAZh05u+psrzpvAMOsUb3ddkNPwbI6T5wRcP4KT2IElv6W+IUjD2EDqIc7tyj2
wgtFg6mDhNLk0eUth3kN9E5xWLBl5GSf4n/TijOB3uhJ3MN5aaZxeowkn10JgJSr
qZ5k1M5ASi4SUyDbeusIjd1hfC3ZzSKKlVy8qv1Cb4ZW3CJQCZxgApSPQM8sB7dT
7O3/tjBKGjUI8xOlbIdkxQNOL5wHnA1gXmUBTozfJ7NarEJsgRnQVBCs17C6NGqd
IwsrWzFck1L9orlvaVVjHFA+39sntZv7YfrA3qWS865vmrVxVBZeCJRSEUp62MwF
Dwq7sSGGAPCTGCa1WxDCp3+3OaPO2X9yP4ye8Rx7uQX0OTXkI3coV4tGcAKMalTa
O8+VUSjuooMZsmRK9k2D1inFxyUWlv6AokQk65oDkt7PgRAADuEFezL5TA3VBCUD
gHcyHbzUTMHds1Vn3NDjr6eJUymd2jqztnZUdoALjEKLyiEA2+ZSdtNfCFpnWEGh
lSJFmjAqx5Qlluw5LQLGPd94McQUMB/HEXM4aBFst83PFmU72Mw4Y26u0lRbT9WF
cX/5NBRRy9QQA25BFcvrA04h3FoJJsLkvAGJtVZQDcgIgaSByXYzTdnqjQCi9pI7
dnzGL5HrDV8ejyDSRRqBi9S+jWsE8MOOTFFr7l/i8g6GOXdHxFxHiapSx6MxQquY
PIspCR0dYBaiCR21TNTvlvVR2iepPrXLBNIrHYxT3EfPRkfTQNjg9RpSApoSBX6h
kA28zPWYx0OQJhi6Bj8W96AVO9SsJXn4zm5ulzqJOgN8Q6ECJ8sFw1VjSibVQ5o2
5IU62TRtGkRN/xSNEmJnTIbcw2fOV8J341D+HA5VpWjfK7gvG9viTgWffZZ4+gQN
kpnliSTRBCmeRDfSH/5u9GQkPF8NtX2GEmegCUt75x3tbiY+96A7Zij2HTVCdRAI
hdZxB0RomcNW51pM9ULL//imTDJYoAJoMoiLscqwoamP/EnkMuz6PjHggp5lS2I5
lvmWjHKj7FShuzIzx2z9etQF98VLakdUB3RNaXkPDfiHbo+Poqd+lA/UX3JGUswx
H7LCrW///YFN/0J0W5IjfDh9OnS6U+Klu7eVQCJ8mPIwGJQzv2KuvA9+7KBgGw31
HhcKCAIanzxb/ZiLtr4/EImR/mNQeWe6GTWkMXtJf5zB2BSLXS6sWwZTTnTFcXUZ
R79uDQmDxWV2VD+oKRK15mZ59fkb9sHIeYTLoW+KYHrQnsjlWbZfNqBI6LK5y230
kG3rVbCe6MEXK0k56Wvxdj5OfUo/nj3orbxAJ55j14pZBWNAPr1tw2MD869aC1ig
7RjtBb8KpnmNjL+3+3B+iZHDqiVlAWUGFNPqmCT7ca+EnTaFGbaP6dWL+EuhLWAw
G2rNYskdcC8vCBI2p4TOeYNeX/1TgIxdUF9yj4YqDWt7/DzyXD81R4UvR5nu9WbM
ClWSndQnG8ahh2OkRxPHmz9x17epIz2ObLR3ierieTOaUNTbZpGhO18rhkGb3As7
tWhPgTVInVobBl/TCLLOQnRyJqedIRDPmELnxyCo9JlnNSO6OSW2uvqO8DaiXhSG
fmxGGt8jP5lwvxW6f3i07xw8z4p03S5wX8tPkAA9FWSRn0Sbfd8IonRTV+zft80t
4+mMP6uQQ1l0sWeOEYAWKeGzlAREo8wlBT6dCK1LMj5YKhC8ddl0BaTtXu/oZkyx
bbIdpdb4ft/Iu3YQmG2wXqoei1NFJSW0S6aokfFUDJUMK5siE0LjF7GBH3c4MVfq
mSkzr63b1Q96ktpuc8+BIMbifDE9ZrD/ts71BlntB/o7dFgquCL/FSSk5lwpdtzy
oiImbGBgDLCs01mgg3807ZtfAdqAQNlHioD7Gy4Lh5LlNGBwIjQM9TzzLXi8oVCs
gS8gnV7rd09dw/7zKc6xI0BnRjXWlAO6xBUCDVUh2EsFbwFU//NTAXNOhvGEnh8B
xRG+xp6wdF79zrSKwwLpVBlQeTQkXUha7Bp6SXiOA8Z5Arr4eR0xXAMBYYQZ2iZ+
cSHd4OLAi8bA6OzNh5RteZxJQ+GJ1YYzHLyaecFxkLQyQEfzravifzNqrCIt1Vxs
qGTs0UBlQHxcGj6q0C8m8HHrKdyJ7mYL4H+ShhqB+p1AxxWCr8mFobyXT66175Ip
k3T5rOa77jfKsQOpEaaHOmlyQwJ78NlSMyvnMlnMU2Ihzmix6vOe3voUuotmH5tV
t789ac+7Vm/p39vec23pTo6CPmsRMxwfEnnq26+h0xXLEpIN6KNRGpzEYwUu4IJt
8aLDjWUcgkU8twActNoQG1J/vx6C60MrJn8aEvtFyXozQpRIU++Yx/UbzM+1XJsG
1SLL7/Q6DujmduKgq3DA0CPKGtSF9Rz/vnC+zae5KoHl9VrhuvYmlaGFbRPk5nmg
RMVPUaI5bCbLml1hcF3A1hR2JoB6sCdTTqzsRF0L8CrHFCu/sGQJ5ElSPvUb6Uja
E8qpjI/xZDLHqZlYEXbj6hoXiVtdxva5PYIzA70vlGZuKeBMQAB807iJUmn5rUPp
JoYKoeJaDVg8a4bwfMcIR26d/yFfHE+28aDr34JsGKdV1FkhWunBxPlOF9AWyUuJ
A9IHgRczjvcLNpypbBe7SHxws/Xup8sQy2I4TKXo1iC/bpHt/J/lpzPjn31znCE0
mhcKBIjaSifMxUXQtQ5McUT+NZW6uULz6cDDwNVrKmOH/vc62NFB/cJDjOwCW6bc
QwVGsY+skCCRwOySWo09NOI5IYFMYEHFELvCJVCFaw2mThREuRAOrsbMSKGOKb17
c/l7I+dMQLbRb/zt7Tg/A8+qFZOtTI8idy/1DAZEUvkN2oX1WJZpC1eUXMBwmv+o
llzggaHYh3Vh2bNaXuRKsRKdHKYgw5nbs/poGxOL2sJv+U0YnGiIADf/BF91LZYv
1Wj74OFrSnT5gOk/BskpeZ1+JahucYLr0bA9cpA/HAOKYUIlYRMBPPTLcfV6fzBs
yybPbZ3i0BtrMquv8k4MFscjC5yX0MN5tHw7G/8e/kdChr/K5SObk9FbPllZHEOn
VJyjkUyhBczHKScAFfIupKHbYw89r9q287eLIR95EntZsTqisEuDEdyh3lOeQRxJ
1wp+hq+ONxgA6bT6UKZmNBk3QdTpwzS6gE7oRO22Cq/85PaTIiUZ0gPHnbJTlOyp
2cYyldNKHWpRnnvfF7tAX7eqV1n6TWYrdb0oP1nhyMihR2PcETQ24rywdEI4ulhi
A2PFjPTkaNZpcJyONLgZpRUjPyKPIeVPr8vNy5mUHtFOd1WFlkAfNjvH5Fv9OSWV
CWntCcla2pEsEkvKVMDb3MvfbIjLx7KxbRW0kojeDYBCuxxUBEHJ9BF2F5n/9KSa
jKAoU04/Isrhufik3zmQSj0/OClMIv6IB9SjZhY+nf1qpg7AJ1dtD5mt3F8/AalZ
FUynf1rpfoJ9HO/DzNX12ZSDTNgKbmjmPRrMK/OqpEVqcQTvvo8Y57yL98SWpelB
Db+icjUkaH2jlfRrJWCBK1FQY588vSqSylhCDriWMyHJD0/t+uzztkhmkqOZb8if
gBMU5MlB3Q4RHnBS8r5pkJenu5Z7B4KQcdGkCFBXyLpiVKVmzmEYvI2hQr8nzYkO
flsQmpy1hErfjYXe40EKMoXo9sYAKYG1OQuFvWWbWSpfIxAnN9NPfj//7Er7ljRH
BTaZV06MYHALUpZ7iYrgGdggn36u2GLr/7J9iCZFM/W4VE9qHluv4X2X5qZnseLR
2RcbFQZ9SpB2+aVurpHvzgzzE4xoRVXwj1BDL+nPJao9h0K1uKgYZBzFmF/CdG0x
bqGKHWMOKmSuvEgpUOydOH+Z/eWIZcbKhtvO3St6Lgpd7sB6wqbsF67woKSMcRhA
vA63j5cpK0q3ePS7oz8ip0uMAyyEOBGLhmSVGPYfIQ/tOd57C9xcQKPnAZLKs0KI
6Rk9uxjHhle3uxJ1TkadCLJoy+gxDc63HVyZmf50yu/n+u7XFctxUbAKJsJKKBlF
RDkuBikbXgO6Dnh7ZircO3q3hxMEFURG5q0WamrlhJSwwHgx7GdzOvQQR6kIv36q
Kn1avOPGeOIUYHQCyEBE4Ld2hyq4keDzZoFpA2skppQJKGKzZo19+ZtiIh5GedDG
y48Ir7nyiZlQdh2Oj80ehmhrpfiGzSpooyD/NngYt76bg6Pmin8iMBlCJFlnIJB8
2hCTltgrhOmzh9W0w/c3EVogtRhYONPySres/UkI63LFcObcey6NjyYN2gwvLM7i
VtMZ5jVi8Z+fwyOCzNcJuMB70Lr5Ij6Dhfkl+gCIxAcj54jb6hqfzmuHqPrzjHoy
vBHYKMtJl9jE/3hdzCLfYJQXG5e/kWxWcLutBZJlik/uZItuHpfCnO0e42YU/lFE
+FL8lNGyc7HNZoHStdouzKU+9BlJ43erKl40zr9dd06DiphRNQbmGj1kmNwSABEo
w7qdK366bBq8YWHk0RUN2qb6O+SBxXRLnFFhDACPkqBylSYEy3FBRpnoT+J56tnI
MxJ27zub998Q0OKh/8bFdXPLxeUaN3w2gvX9wH/PtfzDtLcFq07Ga/GEBuDKOwsa
Qj+YV8iBmX/fSw4AweiVOn09+v4g/btK+zh4iO68Ly26kp2T9Gd1aL21+PFs/yJE
+QWYwBltZQogj3V0QRVHS83YQQ+kAAnmNidGff3KaoraXW/cKntL+YeijjLEChUQ
gh0c/JhJMO/qV+vIUbAcOYNCoMOwJgAUxbOV7LK2Aw8UyA4W2pA7nXDll3Bg7zfZ
KuXI02WEQtzWbnGNJ/LzPnJX0Z/LBIVUCQpruKbGqdUlWMBki8UylNfPzoIYA6iM
p54qyKBvF3tCo49AYWOcs4gzE6Hu3VKVOZzCwI1y8CA71bOMeDHWD6lwufslkXRb
95Q+Y8DaDbsNWvps3+QDW/PhuLfcm1VVGf4/VEj6scMmmOOqUx7NH1HbPmahFibi
h1Mf6tCuKeK+kmkLF68OXm9js2IxRfTwecxYnFtYTLkz78Ewxt9cxasCTIIJosux
24rane1BkgP6hadMW3dw2Oz2uSiDEfBtS/y4Qg2ZCJXbTgz1qU5V14rnYux3AnCG
naAUuUcxDHRCcurHiD7YQqRI+9npQoFbzD1F5DK/UN0T9R0iL7c+P4cTiBOtNAKs
hsHRmcF8YwwLBYvxd4GZex7CAWdrv0IcVslm+kU2ErBnBStU6fHUlgHQ39mG7Qdb
xiakFmixRpt5KgrRLvIEZMDUc+5uRnHNgqI4zgKPgjwqFR11zEHAgrqfM06dzPg3
s0lsUZFbu8adZI1TTHNeD7lAfuQUr5k+njS+ivXfo985KQXmkmQMWXucvcs+kEoE
l6/OHxZ94a1jjEolHSvg/rUgRwxBIIcMffnZd0Jhpkt7KL4Hl+MU2qtCTxwNPiRd
oMVVbfO04nbx8vS2EpW/WNJj2ssfK7g/H+VxeC0tFXGvyIo/FOy810JUChbgE7tb
uHoBC/vzOf8buU4eEaYb0nK/3OGFuVn/vCBrnaV3Qb9lbcyucS6SqmkXh8dBT9dJ
Eg6GTMdZIeKWCmFR9Ja4kLNfzd7VxBj3Hdc5ONZwd1wdWjfzXQtiUcZdpR4bXFV2
g57Tm3V9vN3Z2xnHFXRMuKnmdcTbJEIShS+f5xONQMsaFnQsk6yftYHH1PJMe0Rh
87o02B5HC/CJqNMbXpz3mpbxaRw8XWABSf4rpif+vQ/uuYbv9hpBQtm/f85BDfz+
Vkl7dOtJmfl3NCw99sU+FnyPC4c7Evc31VzMlOZgud6JjGkfW7AVCs0lGqSJJb4t
Xf8EHYi6UO6SugPnugTGPG2HYghcW4FLOP36bGvJo8Knf6porTOFhGOUmQxX/MQq
wVa9zH2Tk1lmnPQI+Lesay6gTpd5l/Gxer/UAnmckyqxFyGqYABnYI8W1X7ndVS5
Y78fb/Fl49QPibLfEgGzHkRocDnDvrNaR+UJllCudehe726gNh8Kkk4pKROVLjX/
VUVBGiPmMJe0GkagNb8anD2TjSpORlR/IyRyekT03alHlcl2hpRv9/mRnmhqhZ9J
+jNaJMVUJTJi8/M7z3zKiwACI+eATGfuQUd3HjHEFhUjuslhcC3yMy+t7xGu6lWf
J01IDxSM6YOl3AhDeryfkjnmSAiMq0rQsPYT6Lf+4Es86diQk8Kgiy4RgEG1mTGR
qxZWoScWRV7eTOQZ6dOY4S1SkAyStLVKjkvuC2zvCaPt+QHCH1f+o/RW2FfeQZly
GMS0DZQ0SQO5KhKzZSsXwTOj4/XnbUsX5GquXzbwyeImU1DNQ5w4V52syFyuSV3e
P/szt9yRh3esk7DA7X6S98lXUN8bpDzmERSN/Y5CGc1UNcU/0J++M+boUW715GR+
c1UZOuyGGgHt+UpFArIIAJHkuJHSZD8x7/tKDbKNJTn4KdgGL9F5BlH54hev7TqI
6XYm+eL4xh4sCnvoTUwwBkYiv21F11mpMuPB6tvWT8ZxW4U9oMftc2UnLKDSa12H
Kt8aSSGH0nIvbchqnh5nLye46yAAxLLIGCULWTVMIHD90Bev/YxwjA8FK6cHU8y/
ujW0wADzF0NnqBOdvhkY4L0xhRRRaRjYQLAghJkrWJyEa1WjppdhZCUPjqT4Rhtp
zdHT3BREx71gnP4hnqV8HEttEZZ8Ja1wAV3bhuSjDMKwU/HIJBgRykyELhSq3p9n
9XXbBcBD4ruwc448qQBlqgdBmmOGpxh7vSLsy/zWoyraatMTzuZUQa1okMCf9FeX
kFJSYuWLM2pBaV8FOrvpSwgnHgkgk2N1vAJhQapAYN4p3vwcIN3FA4tTVP6Oh0KZ
ji7dEq7KpsSF3GpEn5PAAHTQ0y2dppgn7p1XL8aTeNTpfzLarxpTWYrFMfIH3fBb
fwVUAEXmto4bj3vf8D3IBJBPXoqZp1oYB/uFfJLvYCz568WLebLO9IHNvKO1i89/
+XiV0g+g24gkkxeuvpIZLflDgK7vJJY+8EHm/vyv+Tv9n5q7C3qNuWj7tn0rat/d
AmkbJNMW75J8UX8F7W5vox3kczzI6LcMKVOnf2HH+iHshx3gHbLphZncyRAn6CL6
uOwnHgkz0T2GRZ6QGjGtx2MrYZhFHvlri6t6xSDPhv2521dC+8gnrYAwYN0zLt7a
oSJC5vdGuMQPl9CrmgALqazPR8Fdzh+JnGPrAMWDf0aB72beado02ejjHSM2NMc1
iF1Q9nPX7hgnA2UNci0+moitfMfN0yc4bJAmgo7psjlN8WzC73sC0ghVRh7o5OyH
XtjWLwxRdE2m49hKLNTBZcdw0DrxCLGsA6nNYMeafPss0bViNGS7aryPsS3MWRZ3
Oi4t25eHM0LW5tk5/hYIai1sYFjk4EC/gbxbAhPR5he/tfVO7ddcqu2qeq3XTk1k
4wFCYNOdRDCJgyLFNPyk9GRJPjmG2PaOJ58UMqhuepU9uVp/JFIWuMettvKzBMjG
PITvzcuGSwQPrEX82mf/LGl1Yj9e7EnSyWwQ3ekT3UMMQyuZkKNqFesewOoRb0pC
f0/KHS2SwHksiwyPLYj3D1dTEmvSJkMf+2MUjtvLmHDjIOuLy7J5iDCOOGahgVHT
XapnQIlqj18n8JI3jbsQnF621uH/JZHok+cZQKdvYieGGKylfNXED8f1IUwr9sse
96S+fGQk+ZfPHC9oFu3YUC4HnTrRm52qYScLOuKemNbkU6DnayObaZI1zQwbQccr
xrVzo1TR0e4mUAzPPByKvGN+A7fiXs5TJjc6fGxSpZIHVKQLS9eTDXvPGqfYrbLA
RBB1pXfPSWRKJyEOuCsvpEfjb5winNQsGVGu8+xXuQv8bPhvffoCjtewx26lTO0z
Sg2cWtY3kZPQWEd4PgGB5Wloyt4ENcd1C+IXithJ9OQbyWkYDU6NjbxY5p3bbByx
sSYJag/2knUxccPgn+zTaFw54dValsxRpW8ucFnOt/VlU3HkCIW7Ae/Seeo9mq8J
f/VgT+wnDxD83dn7If/Y3ZMtGIQAGeBYIXyNYwHLn4E/ib4niarOFgU0mtZ42Wd8
nzuh8OLLAioFZxNNHydxJTSNDzY7VyZiuujlVq/jP3jpDfHh59XCsihBRNDjTfIZ
6buMpMDPLO4GBueS3Hp8glAo4kq5Ajwto2EJAcGL4P7dH32cn2PShUIYrMwTUpgN
Bxw2KMQl5IwIZHeCNvS2uxnsGtDWUcdtDBRmQIzw33nGBgXpjSzqGybwdp6wT/lt
PfyFpeYJ+i5tZMN2k3kSSCdlUJbHSJQy+yQVCyKQW5zh0NQEy1+VaAGd2AEzxKUb
uADQS37jxUyqWqyvgkjUwpHM9KnRRHr96k7f1Z8wSMUvCjaMEyk84dN1Etps1Z6Z
yJBlbfQ3L0Z0fG3oweuOIiDvIy6DfKerVzeI8cxqojd9kJ6hk9Wm6TKr40MiXJVt
pcmr3JQdAWpWeensRmtYAhWUF7xP+Ckgwa9XD4GIDu1E85yjkrFzO9510jKOYIO9
2w+TbPucgKTM3N3MY9isE5ZpTZWKkxcG2GaPOz4iIEjqzfv6EEFCM8FJCd+xN0ly
7153KCkpCBLlYiQyUO4tpxJZ+pZISLt9Q0FiYczWlNz2ZCwxGcW10lBHJb3+cw1j
iEdsbLLe4a16Q5UPbFbH+t7smhsVHP7GO/ApP4hvMberZVPaE+KtitChOVSSE6Qe
VKfD39fjueb8nDtCl7ILEfOdN2FE/CK7vXBgtncV24RTiIfmCmLBzEooC8G28d3E
kakclN5DN9MdYo39Eb8vgr4FvETfPz2SHxqcsV9NzGBmjoXUEVxhm6xmt5IKOOZs
ya16chDoLW/4UvVUlUOhnVy+NvjH9PeLWti7u5IMgBVsa6weCFPH2nuz0xdwabJQ
nu+YV8g8dfmWCmyWk5KCNsF+uD6PzIvWzZme+pdEg2aKOmstriqtIkv/WPjuPlIS
BRymDdbvEk48ui2N07HhJVFFasrwEsESeADWPRF9LrpiSRVlVGWynavWBcCdEu2V
IXhVetnZDC0F1iQf35/ZNjIq2WbTEFMuFp7aqpoEYDixrLzFPwkv2wnUvb007y8v
CV+pl8SVOVXjkdUUDu6mXL8UFxhv6r2eQSBfptxjCJBvhgMQBT96IRO0mmmV120D
E1Q+uRpUPTQ0KYsC5HsPhz06TIUA22UgEgoTE3PUrJGPzouXzg3PJ2lzPJ8BF48D
1AvdNPfXiDeg/xeQyyIIWwWY2orT18jFshCm9mdaAEcpr7LCQjkzyA6R5oeucI8K
aKoHGcCHYvyJG5WOBtt+E0QzRqgTyY7KmBBwIlBF+tbHgCo8ahUqG1B0AhvzQ98k
NjJkPqyTQj/xUFF49VMDF6L14svPJIdmy8PAZUEm/fPzipsuQljWPdZk4KXkpN/K
GcY1SEqkdEppyZnEqlKs+gMdyERnh+40Ywk0tjjr3WtBUZ5NA5IQXQRkodSgZhaj
qRApG2sWo4rauw38aCOBfa1n0vI/qYpcpMAKwJGntufsEkbC1VqqNSPMeCpn4wO1
K28CneJ136xT++aLZVOtqqr8xEct6YUqgIifYVv8EGsx6ZDIZgDYbns4zGUJp55J
+foDvzrZyXmAfvoGRaYxDCenQG9q3MobJVoSoYGjUdQbgA5gEOcVQ70nRhNEu0nb
q/wc6v2xvWefOF6zwZMGJJ39F0oCkmP8G1WMetSzt30/0R48XPCrAV/nZaoYp6ti
nIKSFw/hWN416Yik+1M/Ng03jzXLz7bbtZLT8P/N492R1mighwuh+xdHYcxLiuq3
6QilUFfBvdszWt7czroNx6tq6TI6u5lzkV72IMmeQySKK40xWGA0BbHWqjiXJIyl
4hYrpCOeDCozp7oCNeya7Pe+vune/WhstKsUHkZtP7vN6Q7elA5lMpcvjnRWHjvd
Nf4PHpUobZJ4UFL/Hkm3r/pk53LdRUxPzzWDZqGhzM5VLddZoYnRY32TKToyd2fI
xEHXDCr5HhoiiL6KTOc+pr4QU6xcwE+Tw2cD+jg7DfdeUwwKERdWQZao+3YkdJ97
fBRjawFywD4v1t596Pj7rEL+dbJLexG4eRRcwnU3dXK/koAA3TKMfugUBSqRS+AU
MUGNXFebWDdshF04q97qX4dvimVF3PfRvWjo3H5GGbpj+PVhyw6TwnOePkCGNqGu
A5NRATc/W7nsG5m+RdGU2hpMn1LcbHHFcVq7Av1pMNbiZXwjMWV16YMxmLl4Y+oK
BKb1wxgMUEwMnu8jlzZILlbqmeeC87D2PLkY7iAtxl0/VjDA1VHr0j8FPJVcDDna
uymozntq9DvKWs8cO1BXLdC02I2MU946EWVyfw0fNBpQZoNac14ln2pp/4XmXmD7
p4H3mJzLoOXTXslJ0F3wuc80MCBibXhA7GpfBD2m+z7VuVABw0zUIz5BZaK5F9UZ
A201azMIbs5gSuFJjvFtVzhkqaAOQc4sw4s61/cXwJyIjfGsvSfTqfWteH07II+4
3J68cy2LcmP6cspqBGGnhzg0qoRcJNuP4W3488v5LsM0xxqHRmK+Pxg4JEqwTErV
60lJovAUSJNbk410cvPBnvt8lkq36GGfHc0arsdd/FmhrrhLd8I+BP+U02wxoUez
CeD8AW/padUT/T3WTVQoXaBskI3lCxoaykicHQ8jabqyxg5J//+SRIzFORqXdYlU
6iKFMCIiYNCkIuJzR0VhPARcY9FrlwPR9sLauDTTbqoE+eiwyaGKu7p9wC5lkyd4
gPss8pCLWeJkj+jTkcS/h/bDXj9O2/BQLya6bVsHdJimsMZdpYULGBPYmihf8rIv
s7NVYsXCIh2E6aav3IO5RxPOXLw6L53NZsXiqRuHp0RKuKGFGuf8DGgz59EwELxR
/QXS24U3zj1xNTPAnAcB99/nUjrdfUQWeIZYRepZMUC+hnXXQU3lzpPOntZzE2Gp
Z9kn55AQpxpHBrrUa1eJB5m9ivUgf99wctjdAAzRZIf9gYkLrE/6mVyIfNyV7P3K
HwI0WRA7goZKsjBr7mmhSno4GvXk7K4RmvEsyKo65BO1bEDkDR4ZDEcqUCAAtrRN
eqfX9qOrChewySPrJC5Ra/iB5WylE6psHHVoffNNqWrflArlYxDYdST4tT8o/b+p
G8wuf5RhYppx5fCNEytGb3h4e4DeXt3b6cPhrHgt8Wkl4VwcY1K1O/AvvrS02o/l
EsB+sJBuiQSoVE1V/qmyjRv9bC9ps6GMgmjwlEI8843qEFkCBaa/k6Y2jWLWMAw7
ajK9/wE2xECI2esTCe8vwOvKsZNBvdvdeOpPCkTJDcOkp4cf0PrJZO8pfJG0cIu6
oz0K7DcIALEblCkaw4gX5FQ1cErCIH6c1/0NRh3pwRTGQSVL2N0JOj+CmQWviDQU
5PMefybAZbmz3itwEWpEGl1364TxdByC8ei8A2/LuSa5xU2x9u+zdIUfxPk6tuG/
dZXgTPTMGPxTRe/wd09Mi0XFsfbvsPcI7+cbrjvGlB07gWt6BzmFtDkmqWY2aLvw
XNgbleaYjGaPsw+FpRjemjH1i2AaRldVlZ5R3RkG6X9cWNPl1UkTzT4XXD3zqgCe
a6ISbsHI1qIKpjacC2iwUPRq9tCfNAQtMysOdKIeXukmMRHh1qvTOihyEYKkt/Md
OZC08sGiz3B5YEKl9s/L6nGBV2nW9acrfyOoitSt3WUPLauD1FZaeSyTHhIx1Uy5
AhiWx1aaQbrENyDIyMFg3zNS1aBuIlFjJFUCQ7Ak+geKCszhHkb7X0BoWKcji0uT
bl0vUpugggaWRyvVpmBrcKfDr3c+FTnt3hTNLLo+g5JnnUQAif6Vo01IKdkhp4JN
RUpYvFB0ZsQEigCUIZyRhaAPKrxclGUv/qGW7cbq+KxA8dJhGu0TmZvgvs9wF66y
tY+hL1g2ntjLemJb+TRtXLL/+LlM5luUoUXownHTCf3IO2NEp/XhCiK1zcbc3UQj
IpBWjLRZ3nL9zBzJjW0IbPAcawr+hCbGpP1UQzV8no5B5CGQ4gB0+s+fZohfUKKo
o9krOOVDhfKthXkM3RrOuyoU34SCsuIKb8VWN+SqmeRmRZImz7YQBrVSgU45q3Aa
/ziJa9s5hOoA6NJQLvTPWqUD/6PNLLEEoLuPjE8/25vu2ohV3MAMxPXD9q4WqxLc
eVB3w8Y2HhfP05ipA4wTup0eNhsrF6JkVRK5J/nap1wSR3MFQkUuSgsBcaVnBKZX
EYqEdPUTiq9exIaX6OvfXIzJteR2ylr+tQ3fTdIYeBBBfFVXsNEoinqcWVKOGJ2r
r9an2V3hXX8BoZ3Y71DWq7XTsENx/9nqTDfz+SsLFe4GQVMJMshKxMzBvngTTdjE
0jGTp3HOJxYCkzRQm3op186SrfcWfpxsAWliJj/xV9b3SM0esokfCMuums79SiBS
jylWLa4APEEl5dD4lIpdP3lQwPpv/HvCFbdFnkOgs0eHQKOoH/WTG1Y6hZ6/tLyQ
31oWBrtx+TRJWI9enYOGSBuHAYGx4FixZLVguXoID59KWfrqDtjW7YozJHEFQpsM
Rdxyb5STc1t35Qf04ZYZRBHhWwhmAvjW4kV6OVWfOmsjVgQGj+bzl6QWAev+chMg
q/vbjpnwII8uBYnRiF9i5Opxe1HC/6iyVAjysg/tTbwr0dA6DbuQcSDb/aD+8/Fn
BZRRs1+MbK26uXSM7HIKU+NbhrSSvtGeBpZ/3uQOBJLvaiQpdMq8svl05EycC2Lb
zaL3X9Zr+jg2ydPtctRAzS0KlLnL/zZOR4+rrzoIPsKYpZdf59helNlaJN+s94zK
jpSQPanMiXLtV6MItqNvtHQEGo6Nyy0V597z/sfLHt/Y+RHca2nyub02NF+oDkjq
cAjtgYLwDC89+p7HQaB+2oU9PMl8yXN1qu1hjBqeWsz5IaZ5Pb6F092/Q3tA0DTL
G3v+ZtguTsgC1ijiM0JZ9NtBQb6UQfuiaJOEzuROrfMDU+a8rI/a4txEUnC05fDc
4G5iA5EjiSoSFLyIyGHbFoZeoH45ab0Yd6/kRH4d8sl6ju+oliEoJQtUoNvVrcT8
HonUVQHD6SsbLtAKVkZKckdgJaF8vwKB6uSkA7A9MFH7G6WR3gajdWQ8ZNNMcWcc
vkHnm5p+P+JlkDcoaqBqCGEZ+X//vo0XF83kog/AI1D6pxaPTtKN/Jdsg0jFZ+BI
88CuMGzZOVMD/6FraIja+x5kOsrsqB2xzXjru7vBxmxs6Nf/CliRrtYCK0WR4Hu7
bW3CRxyCd+ZMlf1sbEYfqXh+qdPqLp9Ti9nAhZxiiDlsPLV0syjHQrb2q2es8c/P
N0Q+S3GaXvnAa/N0scD0OLEz0DoLxbaXAtfXbqZ0+KJ3WGLkcfi66vbfCs3oOlGj
DOP5Fr9XJAqKc0Jj5g/pZQ9AVo2NCv9F2YfQdXU0QIq0uzBSBTsAjAP7doU1LJ5J
KBciwl/ILNoNSX8eoa+VkqiC3l56P0uSG7QY8b1UBocNs5iEn7sIIEUKLMtX0Uva
Km0KyHvk5oXcSoMczs8UhAqLPPpfWdWi6CJdKlWmhFr5MnVN6uHtIx4UahPwDKhL
z2HXiEpB+M6Iih2smOcCtRdTg0oL8wfV9QehFgduWoCFsYaMtcMyQDFXEduTBrME
Y8+S4yQp7rHvC8U8RVFbWFY6MK5lYPP+iEQpDi4f/8K0ZTpmu2Bd0U3MS2YM0SVC
lxcGWSDq1JMpC6cWGgn14AzQ95sOgO7IhhHjrUHa3eAw22z+Omm0Silu+p0HGhep
BUj+7oSxgvsnHGKZqby3mdYL3ufcdptdYJrhwWVbREgpt49WTzUssslaVKpYhgt3
V1N1O+M0IY3QiyVuv4/AAJt4vhVUh80ZLwFrXBKfWNF9QzYEtF1nhxn51/rK1rw0
gtg3CMKtvUEv9QJVqJn+U49OVoU1IkopmR2to3hBG8Pxpfru8gtV11vkvpSj17OD
ks6l7rBkZ85gRxc8SAzxOwnn6o1+T8ATyfYHOzQVVst/3MKsYGuhEkRzBmQUnEyq
UBCHlT4wnjpLvOz7NMzVNWQycDpRfd1oL5HoKhydktX1PjxntJ4/0gfREAmNAaGD
FlJvyyhfQeXGS7pKyyZZ4Bhmy+Ir0qt5I4hI9CBBVRPQKd3VoAvJTGUEUmaBmDG9
6+gi/Q8OgHCyDjE/Sk6MTRyS8wztPFr7T1IgkwcbjREa9yeQaxPEGo8a+T1EVlVc
5ZX951O33lkvRc51M9vGX0cKgJy3Vg0yv8uIbSqx936H8CP/PpB3QV1QLOxhqTUS
6T2nDB8E3bsYm6TVoKfwsVDoUuVqg0eLlhfKp8QHm07gkGsGA81aXzunThIFr4Aj
K3heonH1AUqnVqpjwgoL8LrFOfgHTFLYjGEj+wVtiAUq5qE7MArngRnoxHqRL3RT
GEC6QtjqVpebs91NY3ghOHDSqt3dAQfdS7UiLCE3MlWwS2XU6jax/DZLqlOvUhux
oYPWh2Akbl1fw0lQKRU9F8sYPetp3KwTmvyGnYVX7UpI3d6OiEg4FFQQBTfkWpPq
iFDQ5cU9fxY0eMppdf96wNCAME5Gpz6Tda3VrjSd/6udLB9VmoNs7F9dBkLQWyw5
6ndbW5m2//u0fZ9Vu0ceYAyPMY43QYTsRM/QjNy9fGy5W1Q1CznDQzx7xPk/HSwJ
ptmNJPfGt3cjbo+ZnKO1FJsMP3BkkLJQ0kbu2+EPYgf4dB/excXJWLWCT+DEB+9K
4JpQOGZI19PtjgT6ELlF+Mg5h9d3HVpKfHuEonHNGLc0Y8ydOHPd1HKp5BS8iEBz
vTWS2To5Bh75tzdDofDr88EkRWY8KeO8pbXKTODwRTmJbDkTzB5AgFQs8IlaUj7H
rRn5U64zHTu/VcjMUNTXHYkpwJ1JO1iXZ1UuJgaygEaXfNdw/IgDUnSjA+wHCZTq
ZFxHZc6g6vFz0fYE5ff7cMF7yPteroCjfBF8vYI6fZInwqAhVwelT+1JUTlt40a4
o9n7ccN7fsoRNiwmc38skMimUIVSgEenCEHTubEhu+sVHK9W8HD0XqgH9E/X1uOI
wlRMbhw8IvPxTKxTwO8BaNZkujPOHnJa5ePXmJPDl1ERW0S3oqgLr0852zwMtGQP
dwp36Rw6CifQCypxxrfAxmiCXQnzJI4PvLmaaSvRaktxqwMHuCiQzkh5yhaFFgv0
wqFn30xBiXV2qt926xWNrEy6TgW4diiJMDc5oErJ8t2sz7H8VVSDmSG+lx3emU4G
/CVuhVHEjnaKaXcoejTkH+juoSU3Txl/J8+k3Ag1/NLu0sn47NTT2gbZ13IdMHkV
Ay9X1rqQuQal9ayAUUhoqL40RsJJcqJhI0XjIWT4kySrWR99lBhHkDkoYIUtiP4l
vNpdXDsmn7TbX9M/8hcQRZ7rXktTJeiv83/Y/GF2s3ZqnugRLCP9jSOfkXa7NjYe
P5m+etKiwiC/74GNvA1/O3Mw5U9ciL3CpAazWjNPfhXMULMxjzdGPlqknYYDSTDp
iJfytAb4y3x+0sPtbD1SIPNSMtlt6uB+XmsG5LFOFoe1AcsHj7BNiU5ebafjPLo7
jVwRRUOBrgaiG+mZxPmjzTnbf2264EjYStnQjbdzFRlvA3AKqdaIzZfowIn2i8J4
oxtyBv/Op1kEOS0hffOOjI7BNdkQv8ScW9cPulDCkuiqeqv1Q8khf5kZ7XjZEgVS
wG5HEGGuPJ2On7JY3RNP3LBoImM+VWn83eqepKPkxuOvz01Xb9xjSR/R7PPvUYfl
8zKTYYTHtexTebG7TXzo+vcMj4qO/iUdw3P/GssTqLIu+2FDqF1s4af0IJoj2G12
RYXw7XiZBHRR/6iTJwBeM3kN5ttABalvanq+gvc6wnpPgY1yO9cJ24ZGCxyRkt/p
VADJDFkmKIwQP9xBsUIs0zmxisRiqVXxLFnR9ZC31CxczFyzCfTqO0eFQyGuK5U4
NB28M76LhGT6CEyas6n7zaOshroFaY29aFKTr4k3ixbo3drxzqhp4W00lg2kFi84
gEE7VNSrhslq4EVAD8c/JawyONtwIFvPvL+kxor37wlNxx/hkorPlz/dOpYom40i
DOQ8SUYWEprUJUIcSjP2qCJlteK0+oOz+IFgfk6k7VTwvly2xNAyj6BGngRHT4O7
1UGyXjeC/OzclyDY3jxjuN0VdHcvC7sKwklgmsFbBEy4ZxZyF1RzwCzuW1QnU0ur
2y0+MsTupmbQlukgW2jLe/JnB5DG6JGuV8iuk+BVTqNtz6f8nRkPdE+b8v/BJTfs
F9qz3SrrJL+JFB2XrE8RPjIVUBb+rYNFG+yHfjaKXUxNiVZ2+zaMB4cnhjHQDj9Y
jzesyiUd3zvqq4UIW1CX4sdbcpG3hlE99fbFvauR82yzM58bYlIPf8OuSFwh6W4B
rtFAI+A8AyurvHRW77QfTVtc2ceHmMQMdInFOK6nsxMqNKpFyncLd06F7/1WB8yw
MBy2PIdG6UJ7ySlN28gofC+1sUqYfDiG2jGPUWSmTiDbP4fAW+8YX9Q2y4Ju4UuC
pFZioEnfaWky4FI9RmJ/MCFZnA6G9L3W752n7kVc2CE7u4TXlfLv3A+O3Mq09Y7w
eP+QeYoEi6CjQb0+NyD3tkyUGCziXqoo4AX1DLA/hqBIe8qFlBCNde5J4YURMTqV
G/gKcPmzo+KBG7X+7Lnhib46vFuDUxx07vAopaZ1eITwAiZqUoVpG18Hbx6kO5in
2OSG/dDVaUnwDYssRnStkItMyzVzxZBib9S4YO64of9sZcSadkjPTd1QdQCQmijn
jBDYK9j+f+zER39EphERmrumQ1zumJMuXnj7UWfwDjAyLgA06y/MfLx5vjonUW1P
eFveO6i2a8Ii8xecl6AL/90wRIrRHMRBl3/6jzkqWofcyJgSd1TP35joKu8sfKvy
nsewYgYt8+jZ3MEfkbkSKwLaVnMZxJAs1VLKjhArQ7e6/4NF9aljsb19kEKOQqVj
esYAw0iOfmDj/K3UZBz3zZpXgDymvGyrKenjeosML/blLYb1i6rocMAk373KdJ1h
6y5XacQJU/KYt6N3zdqvDjyCBW9abKZdEiPJisvKdHtQjhDnEm+tJ0soObjd8hpN
QUP5NqnTSyIN895cDuBZwpGKhMlQbJnZNU2p4mIvRqbxqKHTRiGDMmeNdUKZVdyu
zltxDyuJipe8xI+IFLU4JCkL9cWPwzYGT7paps5KUWAvr3q/S4W7lBK39BPOjv45
yNA/XKMuu6YhzjaA9AksCUlITLRKCc7/Td0bffUCpcX0uEmzyhil2LYS1x0DLUGm
Y5KnynPVw2rGeRoAghMHtteZkg0K5/0rf3yiUY8ASGH5Rs6hGYhbS+vHCH8713D/
x5WyVlzyV1o2Bi9opfioC/XAvt34opFRgJN8WN6W6V5wCtIB9XMC8ATidh6nXxuB
CvABXYOvy6/3yIUY85NxMOyGHDtjDihqF4ZuhvGqJdG774ijtGZNW1xxlE7l2Uly
8edfA1j1IJso+h/x1O0EW/CST/P6VT/zHyQWzegkfikOG3Yd8wrHLLjonvVBa86u
etsY7um5xgIyi0X2Wj8HlTa95n9I9wngDi+X5d1SH73CnbuiJ4d1iUgfy6F7qPAG
MipihWq3Lt1PPBkb3b0cjsOIZ825o/EkDrjxCdJhZG3Mv8jbHwBJSofcZPlsrDy8
dFTScj2qHrMDVSpZnzlxAwVEA1oEvUrUGn+2fTv/v0flfqEQQD9al1chFe1rBaxj
AQTs08jAEdStL5yi1ySjRY8HrIpl4Z3mLdpJbafjXklXAefBfwBi/4JrvP93lwJv
hjzlRkQuFpVNIh+RzYIs+FrxVBVMy4rjDBYoqSbGiRy57KVeVD2ShWu9i9wUcM4y
NZwMvhE2JL6JZlFOgctOLP86gdGSl5pzadDsao2dAiAftoCvFVPigNbIC4R81La7
F/Gia7h6HwNNpVUJm7oFjZ8bH0wLBV3DtLg2ZDAXgNlb2e529Xo6ZxSZM55fUMjE
4EF6t8wlwZQCVXTtA0cat5YHFYoNRI8/qMadQi7YVEfNCVTCXyUByUz9tnAQirSs
tb43T3K+BjePwJCqeXbT5yifsnqWj0UYkOY3UqpPM0WVirp+Jfnn+R3ZkP/yItYO
I3k7pdxS0f0/4JHI4GBBi5Rf2LkgjkjHt3/q1L3lVRrpCq1tE3q3hbAkrj6vFnpP
EdPg2lSnj992SOyYkw5thM2XM2lVzcroOLqNvNCMW98Xe7j/Im3lnFI92F94nxtF
1XqARgmuMMAKz3iBR+wjf395MR6R08s8/H4fNMeJynR48NzaUww8KofZm2dXHQfV
yPGnZX+0N1O+uFCGVW3HA8dHHvqW5vdr4bTdCkyqZjnvYOSTmOffsPZU/7r/huY+
DRniMeGC4qcKFPaexggZSm4dD1sylmwH6yek/0zoMEHi7FyZ7d8Ql2WXGShx5r72
OqoF7r5vCq6KLjnGUJg9FapsJUeVugFYWtCrfIFzsuaf3dg8fLSBnCz0W0n5S+OS
2GINy5cGnUpMjL7V+nrHtLq9ZfV83KRN/ISzALwpUwq6W+e6dZd2dw4fBGWey31W
EBzrvuAOhmaLOSE5gvYjhQxZU2YwPD5tIa7x5+InTD8FcnP2iPNZroMLggoDwFQo
gIZqkECGzLgehCIS5C3yv3OlohIVQC0uaBirUjVKXOg0DeTV2dKFpbXYL6SqJJCd
xTt7Myq+7Bxe+6c713ItrGiQRGX3xxoAHGp9NoJoecZ6ud2vGcQ6GHFHiqDCBem7
YpMH8DPXbXzj/cR+r4WUU+2DsGDfCu/hTn2+GcjvJE6dHQCC256MB+jCXGsi2PNX
yYIJAGECkoHe3rW82KotQ6afekl/m+Zw5lZuxuwrrIsEzs7gJT1Cj3VEs7DvktoD
YSv+TgsByAvZDIzzhuA7vIMdP+nB2nurUBK6B4A2bH6d5RF2MlwuJR4aefBd2Ad5
EhvpQWIfPyGcRi/BHD4FM1kJuCXE5wbmeeTl/dGvO6sM23O7CO9GC/rV1OuUZwj4
XkqvX/YfSveF5+Z+23MjfNY9Eu0RGZSnwVF8QheRQCnEyBflkjJQOpzm4ivU7qFh
oTHoRiTp+PFIERKCwC0Bqy0Tn4qoAdLUrlF4Yx3rWAcFJT+/oGAH4ync8sEdrGvT
qzy3S2u1lwv1Yovynr6W7a09boWoBlVS3d1+URTde6PSEUX1zJ9hDq3UIAqRkuqg
e2R6KeMF9yQvMmpb5RtXPwx/jeHtPGUulFtRvcgjDuTeH4iQNZGx1YQAwaLPVv/z
ioUp0ie6G3iC/mqJRCLspOJj6RLi5CpaC4CYNDSFoz987G584FVuSFL2Abbwq+7z
Hd5pm/iDAtSVf8RgADemf1fmGZq9gG+j1qTLMoS4QQ/+04mAi++lR+Do+0YYIWNx
1puDWv2fplkP7ouc+CcV/ukSopwG4UQwdzdZTVrJHSNEnNgrxY9ZkwG1xtIzBXNM
Ac4Ry7zDf/XB4FuBQD1jjQvJJ5qM4yxXxpTi/PaE4wMNoQLNnQn111828soMb7nf
TmW7TvXm0QtxW/CXBd9znPIytgyD+T4vPpykCKol2GA+CzNQDOkG1cHnMUd+F0kd
jVn9C76xD5c1I4nC85n64vWbf/WoDeIPDMO2b/h2NSJnbJfZa3+JfIu6Xe5IA+ai
8i0YOUlPpmF+KBYL55gZlLlR2lS1lYv/RxM/dNdLsFHA9nW6uK8a7RxvXughy8gZ
K6wwwDtDH9gxmk9B7GWfoJNgv0pa1eL8rhL1XoAEFXwZ31yz1dV2P8iNnsfOFRaQ
kg1p8MjKlOHcp12WCMDHpepNNNLurs9+sk5mW/UhBy0v2SnhKI4VaiFjKFsdaZG7
4o5Fka43NRlJBxTMnh71U82HL5GToBKYZ7p1UaIVM6TZlEsWTiZurEFkovT2dTd2
r2wh0VxyVtyxeub7jSpAHQONQC9QDc6C3S4x3V+H+7PiWny79SHLI2CP1kK+24RL
/3tjqo8FghBDGxHCe75Vq1iHkq3ABj0qQenJ0TLGMNTVaZtEywLr7bYNZbGfGzXL
98Om1oYOX65Akt8/U5EUtDp3VMSIimcUkV2/hbGqydnv4GZB7tCTldZ6BxAPs40f
GQ6W6I8INGAb5n7liVNpO4BJIzmWG266WBJ0BRpDsXKno6NzmESV2XxeP1pxElFJ
++f3C2U8cZAD8QAPUCP2X8/fKuORE8Qg1fQ5wntmDyL4J1AmOvs2CMY0efe/fiEX
lmcJFYbJUe7Uj3L2Tm32RGAj6KczHxSPazQRrJVY4RlQzHgBfxCMhXo1VSNohYuS
JLHBS60clJQsM+sstMcWkYnDm5Ookp/s1Nopo6DmKiUYBHSWbG1gxRi7wPbYZf3/
tsSRfsNTsCyY10pfBiPIWOqM1C8IPkScTL3B0SquSgPjfzKmjKX3aXFC0pBIxTJa
3u83gbdCbis5/grqQ74vwLDNYzRqgGAJgLSa7qrU96UH+/3Mr7cm78Q/KiiKts4N
0jYbsJd/tPA++Mk4q0B/w/7nV/S1E1yGEfGjdQIqCXbkSPySm4yuPgxV/CbBVQUd
20s/cks20MGPzHzWDWO0eJ/KO/BLzEvPpAnn3Xr5OdHrhgZ6GwwaOe6BO1PrQWk5
L+UgT50A2tlW9KuhyzaG0/SvDJ6gD+XR2IFkA6yaAFXgrcPTZHmBSh3u6adHLxTy
BdpT77L3DoVcsNFPgLxVMbP5V5XXHb8r/G22AwHRwnJf7Enb6Onws8VY1f8T/dCF
26G80l5FF5UMgLkYO+OxZKyAXuGDyEQkk4NYAx9BJlz7hW0bE9e/7XTrv2YusoND
VtHFVDr6QdIvuNaZKYFU5+0kxeoOdsSkO7cZx2IvuFssAcYrDHuBldrDRr1tDTfv
1ZRHbPB61sKL5y082xzLYiz5H8o4rUjbMM8Fp3zMKok/qgC9FoOv0uqklD5gZpf9
FEP8obGaiAQLEenPMQKFTZ5NA4Wndq0YZRJ5NyFLGzf7R6KtZ1C1d+9GvibTH0EQ
HcsUS3PMQAeLM9EXvgc3AFRCy8wlLEQj6DjVLqRoWgNHTdkRdMF/g1tjnyirBpbT
oeSxORqFlJJbSHJmEm4bTnWSE4rz227QUCKIVE2P4Xh5+iOelNFl/DAPvNjhUV0T
uqxN2lnSs25fI2VOU7n/g3b1TZZVFnjybJCe1NdwyhL+wt/bqk82GVETHsA28IBY
zWFoyDeAIb6mLCal3T/FEFF3MnZcJq/J6qFT2f96jXoBIuazhsFG/WMliVRNCpuo
VTcxphHH5xKjCxEZ6x6vnYLDhhxEhzLWeO2dta/OksoyTBc6VaWSziw8khbu/Wg6
rHWcHgPT1y+nJXPaKaVpsKuCz5GxANvL7B17nXcrYd9spwvrDeXJeHbKJhLVUU9x
400GAChWfEhkvV1gOxIbstKTxsIvGbfvR+H/WIyWnV63LfTAWWcEvy9j1C6KGMBL
TADCTKAe2LPgnSOeOND+luLolYe7E6vhxncf1mS9gjrV/6i8s3MMhUUcmr03cyvN
LRq8Y3HGBbcjCm4qMNUUAHFu3WWbg4Dg46rK/U+XAw+8JVejTHAdXzhUpTH7fubG
NA33G2I0l4iE1cWSCNz5R4CvQvXYAFHN6PVvw5aGFAMR3/omL1B54vP5yeMgeBf5
oB0pF8uQoNlJvOVbPxg9nOjGOwVil05qYxT/+Lr/2ZcXvdfMjhMWAWPm0ZuC5vu8
bGQFaNElc1llTk90iBk/Fb/0x7y67xHy/cnBVAnk7T+KbxOvuijbLAyUY+O2SDVT
b7v1XMzHj3iJQ3gRtSQpzCFzkzYfyUGaBMxkkfdJ92VtENxNpTm7jri/fV2V5+kW
NLpJZl/jnAUhP6vDb7hHDUsCCIJnrKCkIXF7k2InKSiwk0mCdCPs6ONTG97IHnVK
y8mX3or9UwKtAtEcsUj62Ylcu8SvoCWgyArWwlvurR9feAFFmllRIGRp6Pb6KI3L
DV74FxnDG4vMyqq95Yh1pA6SgjQ2PAw1SaKVAnBCgogfzRkO8ssosmqCBYNdSBA9
PTXWuhnRo5gfoc6mVnP13Kt9XPYEB+MNR1CswemRH2yDAu5blJTODhWWhnKdX8RH
4/4mg6+eZ45wF0zhSyUDfGExqfyTcFwDGsRW9PVFPTWsX/DuDOXEPTZsWEU0F7Mk
4rlJiff+h7yPgN/zRsRO9DZntmjlQDrM396Tn9tRknjwRsSBx4jIvgb8Y/TdV8cd
mkgHBWquXTUoveBRi3ZkG1N3rA5cYaupnEVShHuvByBlyICF5koVQQIMwdqsIRpP
w3BxF2KsIep3YkD0LzAGK3ROS+4Tw4CeiITMI7yZA9iBpSXmA3TKoE2gVyeVduPS
gRAEnqWzTbry5LBvWCIzfWvvx6OpulNs9JfmT5v4HX+8QTZJo1yK4GDcaiNWYVyh
VcV28cgtm2U76354UAD4FKhSf5jjbjMtXEEWROn1ZbESAiLH2PQVWX9VuW7ZBh2e
itbVOEMXMfbfGCybwS9WFz8xz2ylx4gkn7ytJyr5MX9d1tUdshJb4VMUiiD3tKbM
mshz25H6aUDdzOf37zfTGQh86T99C7lXOh2Ng1oGQFWDUfxNiJeyhuHu4szn/sBN
202nrDw7v5zqqcaPznJB3hXHeGFJSVWYz50Mrh2ZgWit4nhxswrDuuWaj2izKk6d
NWy8B0PtKhI07v/yDaprIQwyGasdPGspuCX3VNA1dHlkenxnHN/ra13nJ1mwyoJO
xdrbYYIO9HysqrLXUgiaIL69IDYi4Z+dorTL7DYF1zB05z5ORlzm3P5nuiapfX1E
SIWumMkMwo6fk7PolbrNHsVpAOmmEmJ1NkkvFwq8HgvkqF+eHW58BHDXlzp8QrT5
89kyAXEIznOxujHh5zIJaJBOeTwsrghHQxh9UbM1e5e3UquFH1q4fbEnOqpLtow9
APPMChgDjzXkTsapgiSw3fLtfMx6Agquehuh/o7Nv4/cyjEvF9BWFk5Ww/aM0JMY
FQz2jaofC7brgTvj6L+CbXRRcnmYGwPWF9zvcGvybaELpQ+Zq+PFtiq5ncWcjaoF
VOUY9ceKV97jhSHGM2hAw8hgxOHkpmdpyaLI3CAi89ZR2SkLNdI7NJZrT+a+A2dm
KBUCdnl5ayc3LGkSxVYjoDqyvsRiX7f/1GofnmckRqbqvhwF0pW3Edcou1eLR7MP
9dAlRFdv41mu6zGMy3DVgXPih8GA9Ebv+z3v2nBk4CkJb9+a9GfoiGa7u8mzk5Ps
BTw/KaljIRX1sMu/BdwnTBTHQpu/2mrB3qEUyRKTUbXSX/LKeLnVSOFrMU2bjYfT
I7M479i50EtUzR42y0KnOm8a8QTggeQXHbKAs6/MiADuc84bMOv8nnflqD7AWDCw
pynP90tMotPvcKzIqPh/tP/qxajmRNG94H4FOdrKAewmVrExDu0upi1DRtCzdfWh
egSpffxBDfFVSd9IKkLhZ6qFrnuqDwFnn+eGwE4jHU1QVWHUv4sS8SM73EmtGYpL
MFzeA9tXoOh2olPpCEWL2Sejqb/uUychKG8U2mceOa4QPdsT2WGnqs/QvMblPlh4
jaT4/95VzYCAwwdJ8NMWP85fVAd0hHWwPctet9za/WH8tvPY+IMgdaWHlYjJN84G
p2PHKGrM/VXXrm1JDDShob8erJAdhUIuBXDT7g+iEufOaIWMwdYnAi6VNiQYzjvV
9GLxvoqB7FgBG+qbcVEnx+F+slmFCmfyXiBa30nqJ7nNENLjT8ZNg3+ueLPdLn6A
k6qW0qBCQW+ISWZcbXY3+vHDQ4XTmCfmBC1zGSDmb1sCt7TXAkT3zcdohjVKwacT
ynuFfCWZ3yJNKdIt0FdzUc7/Lggalzxf+M8U8qNpfv/GbQB4VRSUuNlq2NT8YZ2V
KaRC6K0EEtLHy7DgLcz92hozio9589mM6rlITY5lT+QZ3M0seCs9CEFomHczWm+b
PHAP5WFrl86u6x9jy5Jeh992SPVZfx/H3RZ//ujMeE7n4KMkM7qpdHhjso57yoT+
ZKh6lBzXWmlC9lk7Jd54geRfAbpFLCODYK/BgPhbq977xpbP3cTVjVRfEs07Xyiy
iL1qGKzOgzlB/1bMAlUWFMzV/yCs4WNczHhX8YwZXsf6fldhBS0om9WZ6NirzxLx
0cXfyYC+ANnCzL//3SSXYzqaM00QZt0UHOsWG5h8VmaSWPjViPI8YNpgTZ9aTZ4Q
8VrB9/eOBdK8Szzuw78T+2wDGaanHJo5YA7QVAbUiyDdYSNBQq3YC7H+T2V0VJZm
CTcB7aigZJaVYpIYj1F6TMXe1xxZnFZpGwdtoneStUB5RhpF23o4iznQD0nYsIeS
8X6tj3yOU3Zp9J3UN+kGnYTE48PRUrrMv4lfwalGjksQCjrVtvHyBi+olqQxpFtn
u0TOa4ZUR0azRFghP1N2YXXFZFEyZrUMeftSCDRekq6qrPuFKR6pMWMfJFq0qQmY
1nqjiMKgWACoAyr0UtFNhqPoZ6PefYINbGmKleZpAaFwBNREemaKRdZjb5rZhZsx
dzuRXOK6n4Anv0Y+dloOrlOE1j46b5SE8E++I8CSewJVm9OEPhAkekH6FYsTYN5B
GjYNSMcrpxSR/GpAgf9cs1w6NTKGN+VAmK5G8IIdiPWt3dvh18o/4qIjTYlOblIR
x8fsNzvvZ6Y9EXz25ewR8bDOuMiwhQ/JlRxnwmfo5tkX1RjZuMecbjzx6YvVD5hO
5P7nUVF7jQsKEWSHYxxR6Soolq8vFOrGO9UX81MmAfIjDxKOmTqt64bFTyyGX5Kg
PTZEAEy0Jf+faZ7Ouuqxz2onfQ5P/JQ4MSEebYnnBlPir3RE1gEsvUjjzAJm7aLk
Jtg+x9/UetJyItreAGLDtrbqG0DnAaLWNIEoF/YRtzV+EVmuxR/oLet0gtjSz20n
P8Qq5IRfJRFHBoPbM+zUf4MZJXWBqsLqOZU1qYGuO+WgsWZ9jiEVlIWiTvqrxlyf
hmd4lgacO2Jq0dLceQnz/TPDhwausv285CTEMHVZJmmq0VQWc8PzPV9yolpwgb4A
tW9YKD6epSnCUKRIOU0ZNahf4uluh4datlprtg4+xCbuwBHhVHHaUYvJpBanEncR
9r573BH0HURTkLhBB2GHbeYZ9Tm1w8PpT4SrAVtHeU0S3iqlokyOemBlzQNHNIRs
sUgKUjy2qKkWK2x8VuvTJusLsaozGy95YhtjYabaSB5txr3sbdtXW/hv7yy2xCST
LxQ3dOtkExytiEwVWtjR9xCwM6pqemKZ0h+LCsmCQCGwo59fn3RDiJgn1MujogPi
jnOwPBW10TIr6+7ItCONYiFsWf8QeNW5rLfhkfRJxL+kE5GuPfk2sJdg/K9UlgLE
pd6nfm+rjLIqRlLOrMzL5JZhb5KqSUje6YCDI2QpJbCKaFh94bGF5CjhJoAzwYb9
o58FtSz1P4S5OKhmli4em/DrCuSs6iUrOr4yfW6z5CF/XCDi+ugs4MrELLqqkKiC
x4aooRzYrVGFdUT4k09UhnSFzdO6mwM2cJrxJJQhqw8KKHvFUXXqUF2zDKv8Oswr
JrJ5636QFfd856PiHOK/8MKwWPr010hpj32vqZy05j3fZvi3AjRhj+FOSdqqrRky
cmr9MOpbDXn93iHRh6NplfP4Q/o5BkIRIkvaZ/yTUniaFRnmCL+Gb47jmI4CJgnb
wtWnhYtjBSDBrTyTlQH5BLas5TiBJBW25b8njSsFVVeVuD+CJ3mXT8HjW+wmmc1Y
acWutodj/9a7F0NOE8f+xLP0knDaTYfuUMGSIf40p79KAAg3tRx5Tyk+WEamKtyi
tVTQomV7F/LdkJkG4bn04cv19/5lOZSxhkNp0ft3OgiJLghFE69nj96IoXAJmUKV
MosEM5MU+qcy+jVOnLN39WfZZCOt9Cb062JhN15wr7+jj7iQSXph92lnorzxZl30
SfCCWcGd/YvQ/uAGPwHQ0FQe4b8C2LtOlmBhej+inZG5o1YtDPPRBjo9milW3S96
qVhChvB+CiuLAUprU66f/qvZ4mQCT9rjxoo2JQABAac4fOW9RKL0CLarN2debi4Z
TnpcEd13m4h5142TF5PZ685x3F2lZi++FhluOMz8RrsXyw2p96bhf8h3LFf5w/+I
cxMrfbiKdxaLeL/oVK+GJAgZCcDoHqc1ndN/jrsdBMZrswWnYSPUG9A/8Jd2QZmO
6lFwDMmrfOiYRfPIsPWIXOYhjf3PzL9shvORNR6HJtfJTKISNKf2DwcFJAi9biyz
rkywKHE1QOvMK5cIFWAzoGdfGiMhip8gdJdpKyA3M822FcTFXCfISj+lLxdqhEkx
zVq3nGnf0G+qAgyuCxZRLuhXPNIxgkehkd6VlzLAG6jBku59aKKk7P0MQMbnPNLZ
ao4ExWy9quKRziMP0Jloolq3DyDX7WBtmavn1WZ0QlEBrx8GY1lNima1T7njBN3S
RUUzMkFdmz+9TxysSKdqADMFmxtyfK9ZYdjnLxwWyu+mYeqNgMQMTILHBEW44Zp3
wPsoTjV3LGHCoUj5SuDoVd2pwUiNN6O0COmJ1Z5ldwi+/H98lVr7e8bA8qkY+s1+
2BGoWzE6pc0RelMhuIQPADmoES49QOJTBF1Nk/AwSPY9aFDJDtWN2OqySNNTU5TW
eqMLJYtbuDQw1IWRogQXDjMvYEfKi8XX5ySXXt5fD0nYLStI+5zcM7tzE0qwwTNY
L8f/d0WBREm8C7ugFgHc8iOXAIisQk5Ve8FrDchPfJww+ZuACTBgKfgKqZcvCgSo
cpJqaq/rpdVlzTrwiATllLLTtjaeWwYG2bLtcjc9Lj4pgunp64fYuZfgJDoEUKjk
LsSQoEjQZCXU6plS2nykfDwVV1UOhTRjAZTwo6mzCwv9gIeqqEOhREqvN4iU7/dS
NSsm/Cr+3eRdPqCzeNdpB5qJtgu05qfELS/kzXqmKPJAgDiE0qZRegayJvntQKRr
pPDxDbV4koEaL16w0DTinxw/Ur406lj+e8nEb4yiIca0pJHlp9T7JGJ3uu5pefTS
/Bs4MM5uNXHD2TjuzZfcHMIUSoSuj/ihAVz6YoWhyEurnEWDMRQ2p4ycT2NU0Nel
48+UIOg0UHvzM9bTUbef2hyCuWsgp79sealr6/Nzk339MMQi+oP7BZKJRqyC0QjV
Do8yCK7S353lZd8NNbEt7yYHSxPA9cyHopkvvkLRi9HvW2Jb6FER1M7WxQuAlWe/
El3C3oFDvj2rCqmoq1qQwLWL049aNFBtayglZ1ZRdKxcBRjNL5dzTFHPgKaR6kR4
2juO1mp/e4xEB5IycpOst8i6v54Fspy9VIwTMTao9oMGfWj1Gqw0soXR2K7as6lL
rmarOVBJP5hA354rwh54n6tXX79PiAUvOUmHQvpX/mcNOodi/v2HkUxjHIVUDPbF
Y9XbwobUbrnebqKcEjhBn3CzYysw78c5nmBgBkuDeGag26JLdBYf+AhgNgqxwyNB
BW79yi9kOj91PQXohjvHExNPSdNFKmdNoN2FC6a+spZ5l9OJ4odkuNbqrOP5W36j
vEFSBJzb22D7JreySobNmZ5EjCWV/I2hhOBbRh/cQv+WPNWtSOIO3YjmvnteOCyo
WVzoNoZgvtylBFokbGsdT5TQ1P/RsY1uP3UkDF9e9Pc9lUIeQNRbMfUl/lsyut1k
Xd/VPbwuXTo/Bm/Kh77Dl36Vk6y4m3ACYGF48w89aJZika6536OHlyN+M9o02Kf+
EXvlYJc/FC51Dp6or4i7iD72ComB8VirNrG9RFa5SXVY4KB6ARl2NVazmqQgd/8a
Kps1+cUSSqhLBbcKgLvHrK3CUDJadtQaEEepcRgx7NBe3vKaMliILqyg4gz4gI/3
wsIcMIpZGSHHLa5ZtHtP/yoxLXQUamydc20J5ZsrZBZU4tvQ+nmxc+6HDaMBshUC
fQ4EIOLIIyRQDt3FND9C8m5ROcc5sUhVDJnRY4WwMja8pRCu8jkAOwhWtpUUEa+K
A9xxIEXhOxpJhNTsZ07iSjw3rKy9wrWORz3RAks9KPwdzhq7VL0GGQHcCrlPlCis
3DFnF6zEpfBRcGXfF3/+qtrYjrDLFu6WOLqFpCaljAkPkrTOc5giw29VeBk/2Rua
BojLQfp4+1qljezw94ttu36Rp16HvrtRF/F8iG54vg7RH9p3xVz9fmtjnyrVSyTj
egI1VhU3ITjdtnaTZD4csX5J3X9Ye+ibS8vnampxPlwhYUs42XRwzsp3shYrCXlp
ZhIXegc9S0Vf92gyrpT7kSWTc620BIS8bYrxGb82FobUYOsq9qUzqQSMsEorG6Dv
gGTx+2EjZ4Yy4Txy4Qt0ffz57HZaR8I2z6GKauBKoE+T3+fVNbuokofVzVamZ5Oc
7tk9AQXSboiNsS7LnIK8Q5PZocnSnJblc4I9n+nN/DavfJSdESZfoiX2xsKejz2R
Qot1OeUf+qnlAIYchjYrHAhXMxq+8rDv6hLGMV5f10LJIY+z5vFKYGQbuU1nv/8V
o5Xrtt4qBpG++6ytM+dmEuAuBnF+X+/4NR/76K/w6WGPol1woTfVgpIXaL3rE1ir
8vuJThaZpPv2kMKpLN7mUqFqTnY9DJUzjX0xrNFpVnZPS+ywN1ClWXIGvhEnnf/q
hTT7YhNOZ3rS7jXoCjRggJwWf7Ih6CeuiCRfaqnuqwKITY9kQtVNQ2QpjEK+3lqi
uaJ8WFjLgqqke3jh+2WcitUStTMUJOQK8dJtlfmeh3lGCh2pChx44YyM91hBhF2Z
/orChbol71tnW4f3WVW3k0R+I9ZHePAFnHR0qCzQounoZXOxZSUomrlNa6x/k21l
kYjDj+EQqtGRcVpvc0ozMh1EmOYqx5G45oxlLz+E9YILtZDDSzyvcE62rnFKvb6P
cXS0NbEvZ6bwtVFqA83NUOEHVIXougHJKtaG8rfmPkXF7e8b4gEXlnRcxlQ/XD5K
ry/pVhOy1hijeJxgo5QeLZBE9XRl+lQFjOefEe/5eAfIO/0KG8Pvq4x/gGea8CwS
J6hEcV4on445kstujIyuRtbqVq6ANdeMnTSgS0TG4d+y3QsVF4HCOG6Qv7QdSnpA
/Gi914lkAgCzSBX7kWmNTv3eXsIMfEcweTKXMZ+sN4Wh07h5fnMDskLOaFZ3fsK9
MA68X+oeDr0GaHImBX3+GrS4afvLD5AvaBHy6+mdEoQm32BOkMamN4F2esPCgrgi
aDdRZhOrFIrmg603dIsrwgN9rUQ7dIn3uo1MxaaNRjnQjRX/nzWjhUWlmiXjJYfX
Sbfe7y60f1aG6jCgRwunKIQpLlIj5xY8pUv36tYHFRnpiWPX6hEJah3iwg7HXGxj
9QmZf98GeUGO3N7rykZBOGH/MkRNW37qJxJw9Xh5D94OPGqNhLGamHv6FfVtx5V5
R6ccZdVgAuoyYuK3QZqjAIZExCpZ51Np1Ss4Uri0+4a4jiJAlBYSQjiF1zFDaQdL
9Y5i46UiKS9bdAs6qxgfWSmdIcFiniQEho2VQGOE8nkOfYrZTWAkcpBvHi7TCBm+
A63WQCmJG6aGbgIZXxkwGnt3SkThuM7/nP28cSTWh3/ywuiaHXPg0LCJuz/VFoea
llTU8RgqAKWM5Tvn5IROh3L/TFnz29lKbR6qK5W/vCM0HyXVP59lm54ajVYRXZRZ
5xpWAYxrJyEzCRqG1CriLU4AZ1do+DCVCtrpACx7ITXjfplu4+HcSJyesynWWCgD
XbR0BpjbEvpJoPINv/WgHYsALBXswmUwd7+IE7HQKPuNTTh2a/Y5O0qeALNGC6mF
5rU9gRSiLiW3d3iv1QZAYuHrysG/rMdee199sqSeYZJxy8FoBGOkXOuhEZffd0pc
Vfqbn02MUinsGtum519sulYZgNKOMMkYLhb/qu0oa6tP+I+Km/NtvM+2ycTCVlcc
ti1BcIqqj1jGP5vlTuEfFiR7I/j+0V5XsYM5abRSxlnFFkefoaKLYP5ew8ev/CHm
SLZPa3H9l178jR3KcoIjV7G4bMHdig5GoICKZOZFynanzgl+jFkwhVGPHZJR7rcr
YkhJ6UQhTsnKQoDnXRcGJt12cMEt+6r/cjLx2WSWjR5TTfi+9ldtP1jxyU+YViI2
h4puwGjLrv63uqVaBm9yna657762OMfEyswkmEo2RdeclcRGLmbMx6zBNiJxTvxd
kbbMJhnch7xABw/Bp/J/HreZzM4WUMiaiEaQtl7xHPRq6LNsZuhN4fJEwL5vyGPI
0QS+0zbkunEi46jjAX9UA4LdlTVwUp09/tfUwm2/y9xPzQRqbJP3AvlVs+kIwGUx
TRW6hVscxCvBqqAd2Nglhdd2KxDOPb65BC1+SATCjiI6x542cqqdDvEfqHs3RHt6
JB3pyJuBk0diqgnZM3j6ZUCSfLWrrcXi3h6OZnspUorGewVR2hhbW1De9FQcInVB
RsfL1yr/wBj+3HugSaOTdjcuWk92RqUKTfS0Mj+6anHMt+wHFLnArLlHPJFSJGsv
KjDpW1matnui+m5FHzPaVybdnUEhFmuFyKIF1cq11anFglCloBv+i1XSTlb503FN
3lLk5kZ2B0t+7GIciQs4oqbsFOHll8agzaVrhVe1zQgZW0c+6DHt1rBt/NVOmkpk
LQja6MrvoZoKRZkrxqvj0PxHxZORJp3f28fP3j1aNbdDkPaXqnKAbgKPFM2OGyyL
d1/GsWyVf/rwjhN7Z9O9ldJFeFPaEeK/ri22yGn0WbBC/SK0dXCzONjtmLoPpFzI
HjJV7CwHIzQnAxiKmQhCS1ILfXCm1F/ScGKv07hw48OTAoyVbRtGK5Vub3JrZ9h4
lWYpR7dYj1Q+mhaGkBSQAYu3bt6i9NlZta4ePh1qaQGCtDvrIBGUZrOhGmxw2qjS
L7eQO83VeB0xdev5Kc2PF5nB+vXazGF1+aCQN8BRHIgX9Y9aoCFqqvY2dQBSf3RX
yTMwqZCoHLoeQrbAItC7PQRP3u08eAZnBqCsCCOWJDutm6mK2qtvC4oyGH00nmDv
iRqB1vcEXizwBpENPGnnIvIZMYcATiy7cFuFN+SVM/mbyR8rWsvcz1OPdsqFnKaE
MZjZ9OLIVFhBh8ULAW1D+CmCVAJJxSHFoYqcq6NdX7nXd+zWvfkOyXU/lbyMkPXu
WyYUOEol8HfBrsgGppiR0BDISjF59pGuC5hq2C1iQaanwkYTT/5FcxdD/FLOSY+7
SBLeKrLhRqVzLmCw9PwAcDnSgthXXsitg8fUL779WwTwsyCnc8p9qrGwjIQOMXUM
nkWnJSC6ShL/bLh+IlCI6IrybZAvMW8AGFAYQ6uBrOHEPoi0NzIO8b7Zc4F6TM6V
MfknzxJzY7O3iz3Ke3rC3jMr7e/m9qOImNrA2UJNjcgylicU9ycwUGF3MePp8eJv
FEHICZjxibIzAfondf4KtpNwmO38JH0tR69fG7bpHnKwyP7aNQej9z7JgSK05y/t
5rvMABcPsmcYFCaurhaiLqD4YiFeDzZF08o8bMVG1Ech7Ju89X7u7sRJd6LgddQJ
LS4nJUgjPVxBDX7eFQyr5JrqlETJpQZZfQF8zdtKcOSpdkk2jW6CNoEYZgvOuEpZ
XZAq6sfb/oaZfLJX9y/bP9ZT3wjiIpuyeP3VbXcbS0weFGH6uevu2D6rda4WbE12
+64OGB7LutuMZ8Q2zv3TMm2XclCj++tdap2xF4YfEY6TybOmXQzRHE0VxkF99cOv
zjTHK8v9gD+IdlmDf1HBvEZ3KlRIwP9jA6k3Pu+ClQ2DDaevA2tqvKSefbMZCzMk
rEvtZb1rUio+t0Y1sTZtw/h4eNqnSz1PbeBVqmGif5XVAfTLBSB+eXfUv5Rair8U
YjxE0Sn3awbXEgVi1c+oolNeQYTjA3EeXFRnLOFF0kYFVoqjjg+UiV7DFEdg6fYP
lY24HkYWxIxkZYfe9tEqiKtF4E0RnNvky1bBUW7yznNpzfnNOFbiBWyLp+j3SNSi
niM3xJAfvEwjHroOKUVgwsDSpgkq2xpnJ6Qoc/oNdgK3cbkxSXkmq9Z8YKSY7gyr
V4a7rhcz/eI47RsfqZgG6OW9nymuCOpZWy6brl9iybYPxqhYkvTuymvyvWIG514w
Jm9igOj1L4c2+XuitseDlZhVjSFF8MkvQKO0cUx7d58PeYNDqGh4CYzXobazkuxm
KfVUa7VCEf0jCffkghsJ8D7/Tzd2xzWhjJrMiOG+3Yyn+mhnHvpiIfvVuLTyNMkG
rhB5vPQB/rbUO558nLA8MxZBtjx/EXsCVzedh+5JKdRoIRdWOCUa1H4zKEioQZgU
yZUjOPAvcaZeriqvEkTAkKhizs0JsoENrLTdFU+6x9LYz8abW6FZXA2UZG3iAofi
rKbQ3zCYBVZCE6jahHAF/a+G282CeFj/qJE5XjMxhV6q+eCag+PiJjr3aK5cHAHK
2VfLsxm3dyXMc8E2Yzo1hNKO7hhvTzBMPIMKPcCVhUhXs4rFnftlLkHJfm8jJ48/
wORr6+Mu1WfWhE5pcQ/u+wq4NOEOgCqJDVJdb6o73SPYxe3njYoaiBRuoqXc/D2e
fS5kLKxXsiukEbM6hgS0Sc4YX/jOnwFGy5me7v725ebSeDINir/s5g3a4ib30fRU
rD8ttAqiuFBunUkz5AwWaxku6B+IdlSU90F1z1RC5kg5ng/mRSW7OPzlbUave+L1
RBtLUhKQY/kUKCWYEG4tQIAbvHZoKrFJztHI1Dn9htELxPtDNPX7UYmWUaA9KibD
z29lKiL1ZUhViH3e7SrLNgnJAuFEqPLt6Ks2RYp0aDPPY9jbhHs9i4xGo2lXifgj
mzAMEOr/AE5vuyv4gihf8BnTfnovb89drtDuYUGFihLz8FvhJNaijsaHJYz9B2iZ
zKiCO80uAu3g0yAS3KDb5ftfu0F0Jz273KUcgvD8kZt9jYmxqW7cpHhb/QZPRvCv
wfEpMqUEF3U7uO4OVQ+wWXW6MgOvDNquq2NtcAk1mc7BexqfXYT4MuBfv7DSiy4V
sYs9qsGAkLogACHiEKj1y/cdxnXKUyagteBgNMybOyILIUvG67yjZQmFz7dCIz+R
/2pz+lbHPrPjBwqvi50jLO8UfVk9xe+KtOurbhrEhQeDNmM/h3YJzNi7/YB/sGwh
crVvLRese7H6Ct0YcpgrbuJ2VP1hWngIH3Y+UNDCqVlsGgptKyvqNY6odcgAL83Y
Et18stTCvfwxAk1Jj+ydsOxNPDdvElgsRM5r/CqFtOifyUw1CCWg7IcM468Fdivo
7F4NftLtnYDLOWeBejgRVfAn9w+uGyVRBNjOSNMUT0uKObG+Xv6IPOgZMgSJqkzx
gElh82BVR7zEdyNZ3HbLXsH+rqmp+Q/d9xVxDpP/a16rw2h+rNJqbSuvDdBU0l7J
4+8tbpntODmH/8wxQEJbK9PndO6cqG+bXMF+ke0EcmYLhRlwGgmGS1/odHuWRDyv
wKre4zj9RM1eFXfkmSNJaYZSnmx4NmUm8xxl9oScI5CFwax2yYeBvm/ak4hwXubh
niFRVQIxDtfgKCge0i40DSYpxoSzEhkwAAaX4eQa0cYsydUOjIBiUg7V0tVzq/s3
459FPqcWdz2IxgzdXOhah7pUQ/xpFatt7WDI1GYYz9tN9FcpkrtS0xjl2/Ik0Ov/
2mZyKeaEtnRJIoYcDsD59aGary2mbKP2TDGCiKL40d4BagcE3Yx08fCqCPH17eTi
U2W6h3cx8uY7dHIxnoE48OiHqbaLCclAy2VCW1CZQmtGUjH9niEwv3B98ztipaG4
Tgu34fGMLkJqyBEECTEyy8e7wCuQWmKfsOAK42x6fibe97vB6fmDGEBFxCD0vxuQ
Kj8z11KUUPYvBAHIoPiWYSWVtecxLzw7/GO2m9ZJAtBo75FZgmR68oegbbYH4CCD
hIVbRsEourSd3p3Q5dP0McrN18CEza67VEBBs3h/O4aX9rQM0BThc6f2Bd42/pVP
k49m88to3ybbd6LRw4M8V9RLpJu5vuUrHzOd6PppNYhvd4xswMcSxCyc+oNvbuh5
AanP8NLeQYLKa49OrVHzGhBKThhtYQyD829vLuCGxO/tbRIttr6kkuqPgVuJdskz
Yz4FYjdL0FdpNHS6p6bR3ntBOJxFGtCAnD+jEtpxthz6xowOy3qviwT0CNIBMpvZ
Ox+E/iSkU8urAwtuR8FaxXj1w6CH9A3xRkB2ce0In8K2drjw8FvtkAN3ykZrqFxf
NcFMO21R2AVoSHdXkVfeNXtWmJKkTX8UWVmifKyg6D56p1sWMKUYso35AGvv9nds
nbdIOZcrygLCcJVSEvLpiSoHUt2sCWvXtZe8z1dBemuJQdoqgBXIJXnqode2zbjy
yQIMA4pgma2F+qxlDNLllYKqpHi96tLkfbnLKt3slIQni0tb6ftgOh3jfUBzl9NJ
od3upqByK09UoEoNLJYasRqJl9E3vcmdW+151BAnnCC0pKSq0y665FuE0TA4xm4S
I2k7FiKVslBXD3rSklejGLrH5jWFD5Te9V1jrxrVY/5fwRO4FNa4FbaUcxkDZ66E
4QYT2o9DgxotGDFClG7RXbYj4XohohOqdt+xioW/PHPrTLH2WDeRMliaymA2COuF
JEEGzjyor2Axhb0G3J9PXFPzaT1gQJ/dkqwBQRDAW8TTh7IJ/kl1APqwXgBOgFqT
KJTdD5SWrePF1Bb+37UvjM0gQzRFMnc7MKmYuBHH6Xh5RTaayjvlRDbu2ftmoxJF
LfM/1EEAtvLVwa7RuxNcd7n1O83JCGirjq/DilqL+yi+Mpm/0rh+7si64pWsRPqO
bEbrF6xtOoYTa8B09rlpvfv1yUvVgR7ZvvHrKDLD6yX58BA1EJPRmJA9+M8E8nuF
QSGLZWs5LQeD8TIQym9lefrFJ/+34qSl7AefbuJsOfM4u73l5/BKOrQj7l+5ntHB
nys9evbpUlplJNtM783/MipB4D67jWAJBFMxAkyIY689gQiVTuLgKwdiCTVeR7L8
gWWPXK0CbMKij3fe4yFX3ZS+7QTXO4zA6yr7sHavfaxuGnj4QdrnKvDClJEBaImQ
wBylg1h3RM7PDW7TYr0iJixVJmTvebHMWQy/Cz1xQdsTugJDosE/ouCEsOEmOZ7S
KmeK0ADLTHEn4szMdqtud4RmUg1k6y9t2vhYPJlrKwo3yLUX+vkWARLmtPtnBZ1S
NZ5ztftI8gxeYmhIGFUa6IOYKmf+q7/9pN2rud422CxXYYpwO/SQfL/gKdgTpiPY
PzVwScYNI7tN8YeBrB4hOy+jtnkVNJgJkAeDC3L3yLUCcdrbAZMxyTxrJiS7/WfT
1K51vTGV7VHoUifrx+6rQNJT/8YDuiFkQDrMEd5HkgOtjn7nazuYIIIR4ydwF4ZR
HQB2VU7aFd75GFPuaigMoiquxLjVYWGQnuRhTCphPO2SDr8PaaMngzfCxb0sqYii
lwS8gMC3k+TJ+IuNKOodpqJNj+VU7l94XiWg/VjwUA7uymfFGyikBbazACjT7hrc
FntgmWuNW+eofUMWC+CfAt6l90vQ+Kb65MzaJxnMGajc+By/BuPOcHHhj4Zk/l+R
1wUU+BzsYA5n3Oor1BGCzGK2mTUU8yliRR6V9NsaQKfVQVoG1nY5P7E5AFqsG01V
R7XUwsfWIPeQzel9n0CTuCwymFVHlEJhiaLG7ZZ63eO1iu5iuJyzqPpAIaWSKPLS
qJPhybDIPuOJMPuOiqoiWEMUi7HAPQDQdQAvnFoIYXl4sueuRCrQUh8GHoxY+etF
MlsdEKGK+1FddNZX/TsnEOS0oDH4N1M4Z+AlzcUPznMdd5ddUomQb41p7/PnpIkd
xYsE8c+twQnWSLWzCCjayrA5VI/kUaWAp8TTxTHNYGjWcLaJAh7ARCgzK9DdytlX
n+oG7mrmjXZ8/krHqMq6MHE4nEsevyxituQOnyO69T+qE9UKgr5+hn3ohPggmHmU
fZZMIjmUNyLug05ZlmairgkQcAWBJ4nDvqVuqof77BhXSZBx02o7usuep5fzMDZo
Nz7wB3zLgzY0QYDtnvf3LoLEzJZ8AInA2qh4X3n+W8luT8F6Vls3g12UAFkJ3Kx/
xVI2bPCSkDyS+CnJcpYI0IVvboClE4fbkyyVM8PTReIHPxnRTbxMCR1eSBmY9zOI
iL0dhc09AjWRU+gMR0HowT2T/Ssp22I4BjcdfZVnERX5pc/5GNB0eYrVvqw5oTQX
DsHLCL0yAZhAJOfXWY7EPZmT4p1BTdXf3G5b8mEUbXyCA8TnZRMtSD1MfZVHzIJ1
ueHh/ye7ON5T2sqA7vJQchqLassO2RoydltxRoSZRvSIMkqmABZpQ2zocg4KCX+b
5nWUTmIl5Y7VeES+03ECQHDp54HtrgrZE+UpdYZCWeBjpDiaiOZ9YY9ehHFk0jyT
eGHDWhinWkLnKXfRccV8/GDmOe+WqKKhekwkfkwLplCa482V9NMG3Jr8iTuXRfV9
xNYjlHMc4jbmKDbJiDXnD6laqWEDSaZMR//NcZgpz3a5AjAAG8nClZr+3SKMYyoA
rxzFjiaj2mrkbZXwlfSJK2na83eWncu+IHld9VmO4cLoB46Hs3wewuGvHNtQ2VlR
0nfNFwTFmyKo7TyyhdV4TYfYHHLx6jF2bwuya5XyAGQ88Slc88hLnBdHTqe15XHN
/Y11k6kJ5DEJvP550HulTHZIeKMYKnYWctzxKSgCm1dVmh4hhDxlEqWzKaO3sEiN
dfwJo0DsdU4ibsqmM2uT1S+QTaPoxKf75ezX+0p6GCN4H6XX8PceXZfeUrpvPvk9
XujEsJTgdAfcKjTvY1Q+AT9TMbClt9G5gQ7GMuEkMew6lIBf+pinISnQBIpXMOMd
Yn/ZK49jzHOliCJfTYgN3lWsuGYJaOuqV8aT7ebn3UJoLJAOv2QVm2oBHNyEtQgU
pSBRajMABM/JnVlA+8UvPnJwbqn1h6VherFNgTrd+bGlKZc4ie/VOcWfRc4y8po3
IqFwxxqq8KAB5ZkFWDhKy7LZ7E4eYtDDSQF08q0clIQQHFN97muhYuZWnvqFll6l
H7tGanLbdcuFi5nvWHuoM9CpVK1R5szRjzzmse4wXrFg7YTqf7/jaXsGmAIwFA4W
sV0bC4cjKBRATTJGeFmmO8HPfsw6t9M/eCiIBJgmkje5s6k/3ZFscF7j22ZZjEHk
v7R8HCPW3zXhKT/aFxH70L/se4cJVvWSZNxt6g8GJiz3LEakgKtnuomoaiG4tEKo
wLLmffGeZsLFMF5LZFU6ystcAtno0ml8RUoB6an8g0dhJQ8ebKxC/CE1XsJ7VOpH
HS6cfoM7z30WthJcDo2EjMVTk5FVsUxgE/UNm/gluRhHZOXg243Y5U587NYwkwji
9OmluvzrmRqg5IIJhh+6OFWTTKgOEZnfj/hBoxDhesFhxfHsZoTrHVY2ILtZHaBz
LeaB4sCtvZYl/8lL1KaMirE+cDwG6z7w7zuDNkHkJXpfy0fFTUvi0CiXMTHmF5h5
VVwSJcj7bhb6xwbuE5VPSqv1M7rCeuwFGi18cD8Jn/nUEmi8mVcMdrRGAUFqFYZv
Mg7yhOJNHlXeoPhsJdc1LmwEEbpobXLKP1EuEmY1R4g/aXMSDFsIMuI30POZkLMD
KLqFxDJAfVbLkfiMzRY8kHcsOu9u5/AmIXZRRF6Xbpnyab018qlVyfVpcOmmSwCU
Wlag4jiSjki9wRXFWS4HZaRvIP9Hj5kwRcyfyWYGhnuvqr+4GU3ng79qSYOL2k+c
XwJhj1vQ5oYSez//bxvVQ74GScJaeCZ3Z6q1zlc2WAbpbqtSl9d7Fo0LRgqjDeXv
cY0lJBLOaziN7yM/7/M7ym5vxiGAl/8fZFKFPjvnM9AgpItaQ+JZAREq4EDRFRD7
htNmCKPl+Cd5Wf8/jPepnI84cEGRA2JhAItfwbaIA8gw2P4k+xRUcORqslAbDe10
HJ4pAn4INlUu6wsBt4vOXfcP0PxfdA8wQ8CQ9ewaO3BoKdwLyPt6ihXqwtGCNjWD
vGHDtt7cB4lUo700aaX2vGc04iJyhZnLRkwm0gQ1Ul1uvOYtB6qxHffSdxeQV14w
uIQhQx8mWm6lTTm873vYFaQSay2+XDd4zQQ5yXdOxs+RfGaIkaC1urccnL8d/JW+
b9USAkt+wcyigmcQBl/rLtIiLhMww3+V6D7FXV8iNBQom7nfKdVYNpmV6igaJzfb
e88U9Kd0hM5ETpKyCICF+c+YPi5rUt0PSwYzAoU6CIJCiaDfguAZjWfomdfUtdNN
QWHUyPw/Jtz/VUEux039uWMOARqjGWmuIEh45KmHWROVjd9cNx7Nu8G45UEnmxIc
IT+phWD10wXHUXQmrcvOMSRos2r/mumNwSLjA+yL0piuo136189OkEKceaN+8wZR
WABKgd4jnDZMNSd8oSCzhTdsrog47XeLKxMfLvrvvfT2vPsW2gyAOwxryurQQMVp
200TfKC2wDsP3v8cv21wSntJFUWRBIYj1TafqyBbdMyRck9pBZruCl483bPg04Wh
9IZ2TTYI3mS8hvW0sC5m8c1W7vsqzPkUvsmGECCr0W4/1icO5R9YDD1iyspNOx0v
TU7Qb6W2tSdyXnNgCyD8P0jO5BEnZgYZtTRPINrJRkBGgNt+a4vOrms8/Bs2Oopw
wCefVEF3812Lf7cO5g32Vmf0MumYWkzIYbXO08FhMnR/jnLUsveM1YwxK/gz0Y4z
g6LOnP2WP7jAA57lKPQKSC8XH+sI7GF/4V57G9mWfP+q1YX+P85tR47cFevtzh1A
uqlMkgU9QtauvgjGCQPa0lUKk1PDvB5g3gsXkahlvXtSRyqOCTVBTi0tOZ6EJckR
3HXtnf0UPvuhePKXKFp2GDERBGscm1EaS328yJE+m6phwfXkBHLU3h9qGut8qq9G
zrGA9EiUmIl8vig8vrn7qEIG9BRqmrwqkghxe3M3cgOEU6LWizko5qbqJF66OgS3
iljnO+urrrAaDT/S+HolxyT8MtF/7w/AGjQ4eqEyGkcUvALuesPlRH4ihgSRBEgU
YTGebBPBqxz6NxRRUZMP1WLLnc+6jpl64emeHHXAYuGOouBXESsgVlE2zjWKt+RI
aHzCT8/iUY5wQtaTJhA0LL1mYbLmOqvEHiMK7+3pEg0cckfL0d8ElPjWZKhOOGSe
pWSoE+fzIn4Xk7M2KtLubJu/6+aDYJn694v8ntlpMJehD552GuxsiIdTEMKgeGCx
PQNYfPGUWH7BJw+4SOLzlQv/A/fkvorTUg9Pbtpq+CvVhGBZGxGpB81SzTVuZ6o6
XIoXhX7vh+PR4Y54YUAUzLROK8Z+n/u8yKaZpDcoR4mGVXBqitJ2LE8BfuI8S6VI
aecq3K6vC1i+riA/SmiiEpL+IfCmALsINFmZ9FLYPuFOWR/UNltz+A5d+EIHWz1r
3yB2U4sa5cKlgmNkZQKdlG5Foj1g+AQGVojzJuNh6rroawSu4/UB74mLCRrtsVG1
8CmqU33WaYPnkPj90YSk1RonLfM5zJ92iRj60ozJQVbkIUQZmyJyB5gkyRjs9Pl4
aTBjH5Tyi9OBeSvAl2FKHr9/m3HBKxH+fFcYs7gnmt9KXCWACV9rQ/9Xud6znwGt
86YgGnRgIOUvfZu6hUZskqoZulMu8guxT/itXllF61Ow5BLG7lnxOwd4uvVNXy6S
hOu3mmn2iLqINu4kdRdwWtIoaQwjAszneLb5gTiGYMMPLNmIf9oU8fpJCnND6wvH
hvtiXtk0GALiRQFTK/NE0BYYi2PTMFtmjZE80qp0gQ5Zp+n8R3zFosoy3V5ah99R
kHnBCfyf4e2wp6rZxhqGW//u6WxhQVWCkLboJG4o5Q/Wf4a3dmtptsh3yKgzhNXY
ZohGOP9lCnjUZkNMvsGBXWboZQtSqLSopzRhi2TdTVj7rJu1Csg4HRK3R/WRBCxf
Tz73+BwvE+3NQLz/9luPJZyi0hL3Z9V2j8TVFpG/e/0mUvJnwhCs9YRvYbDhdN3F
90JCmiQWO9bVAzDKKs5PpQBwq3HDCKT+Td4VfSQy5ek9GukfVUHN7Wu5MKOXI5xK
bItqVzX/AABOp+mhqp7HVnDx1JImUlZzn4MJEws9IUq8d7gczE0z8BXBPli+JR4D
utTOx7DIXWrh4q96PiF5VlQ+Jc9KIcE1PGkmtYjQ65BzGUTbh3pAL1EHYv7Bd/oO
Pw4NbrFB0w9+P6ib8eDDMSutXkrhsOt/HidoAZH0wm/w+mDlAHoIVDaCTio3SdMF
KyPPggZ2iz6mjmzQJ2YYuDaw0etFDyKJwrodzcWvxNfH6IZ8g2B287co2edpb2+M
WuMKEcGUr/DEq9+d2oZnCUzKqVdm4w/JaOUxw2iXruiud38Ho/jq+kZYPh6vgoib
ROxoqQrwmWx2iVqSESTHDMy2weH1rKtqUdEjLevnNNQWLnNT8PfXbo1Tzkx6VklQ
C5SrNLiPa23yJWRSID0cXj0xFYvmi4aB0A4Jc/1eNxNGo6iVR6nlxBn2g1HyL09u
zbA5HSHX33Iq/0n+5Ljq5L6fE5dhpDSHU2rbtHXFVJ/QDjXAu+Pjl8dsnwj34Q2T
Eh/E6UEj6E0FNaNrTwUHl4yQjFFTMswG9mqlx3XtkIXYiNvOT5x5XvrTe/JPABV0
uWsm3ZSeE/kJdg6kP6S/48KtEsyDJ2gu1PJ/XiAkAqgA+bCt0mqM6gVZhVI/1rut
OnwiPtT6EllDib//UKM093y2/4G3kkWCdo8h00B8Cei3XPkYLiFmdRHgQJaD4PMx
2nG2IvPKpUMCBv0ebzmA8Uc4vxmfai/FcygTwA/y1nPhpBe7ruKizhbHPZu+FTRV
eAAD0HizE/HeZjdaIGAyFcSGp9TFRF5KIqaMKcOH+OyVu+QrBC4bEA2/avqZVb7f
jPiG0FBUeqUgOTSJM7pxvRDJQEHULXtXI0hDU/dvp99FnXPX0zRJrA0PXLdtSVAw
UWkBZpXsByKT145UDaITgudnrMXSuJ9bfrX5PSM6tl/je9bQjOIb14Bh75tgyqBr
YVU542BRld2G1CpW6iPYkqdY/q4BHY8yZQNdSio+9AGhawFWr4Ne/CE9kMiirM5j
CX5clUs2gdb2wnHuXX3Yy9NUh0J2YEjn30OkKp5S5bszsRJdoqa/A7Qa0lMHvuMD
BtMriDjFcu14Sf6VBoGc+b6RXSX+cNoypxlfw5TaxMtc0hQHBf1NbdVtkUL41vwY
SBmUZ8F8VBU7UOF/zxY+2QU/tXx+Wk5QWywCXl05uaaSTElj9VZOW1qNGZ2DmKMw
Ddl+7f8uRQO4hBz0fUmJ4t8hbd+e3/HI1X+C9bNN/IYGU+2ZV9UfLM+ZVTAI8RYJ
E3JzJMwbq3qG9y7f/IljPa99vckIEdAcvvWcR4B1Ks6ABvkxrD9pbFUQ1pziMKl4
5at5fo+mtll9OAIw54VRxFOfu9fD49ymOowQ5e386IfBjvMVNmoHIkQcZz77bbng
MG9ZbvFEYPzm24NmAs2QMBxLX0dSMUEJEq/czNTf8jbC+CaD0/hjuibvubq5vMNG
SbEcJP2xeAVavzR1T6jN3OWG+lOt2GBaPbprrwHNT6OyPW+Wayr6+aYLfu9Fgqk1
tSiGGuD2n61DaKmS87TMq5sgyM55o+rw/BxYFg2cyZFeMMTOBr7tRqZBIphAN9L3
lXrYhEakyjqvpOFpWpG2qqTplfeNtSowA7hhfTQAPxOov3R5KzVBalAIgsbLlXae
bHq2zSEsLeNtXMHqyo+tumNfozRG8DgzQzaxjKeqpjFc36IvksOnMKEH+mVHQLEd
uE8YUMV+ePNJ7mtObmP6HF4JXiZeqb9SK0HQTGC0Vy6iaKNrkhzlEtopKEh4FsPx
YhEKbsgG4IRKOstzLn4seS/vPa0XmHAqOfz9pj98lhSWZ7GN8RV95bds4QZcZ2kJ
MqYQk5IIyAyMapwxuSi+zV2vebuH1dhpplKsgIhrLawjXLj66ze2pKlvl0ONmTK5
pjaxQmcS/1GT+PlQhKLhUgtyhXM6hxCRQFGYzKlUhXJOvx4twjMm6T2EAxSz1/IW
VQ72HQ0+2Jr9H3q75n47HAKFIyKw/tjBmafKU32QSCUnIG5bhdFlh2QLV2ot4NYW
h2UT8l8zZVEHpV/VXIjumlQ45uuofZ3ANlEJjUqiArkFYjWGCJFZ52Lqyrr4gBhc
KVrdP0kTDIjQ9rg8HQr8+r+Ym8lKun5rbvPs92++nsyHuPBNGqDCVIYGIXxG3KNF
kAK/IrQK/Re23BxiYSn/a7UgOQpAuTmczLb652+tnbKyTpmO14acmfiUbrVM5baM
pgkt+hiH+aNq6f/4NvMTbrVbx/4Zbr2LuHuavVGHcEcAAtaF4Uv6SCfqtqYjOBJr
TFohp7Wol1x1FIZAb6QVn44erPGCXfUeflCNsy+m4DSz7gpQZgpw47k44hiFss73
bT11HS4W6Knysk1kCL1Dghuc+2dN0DYqfAdkQhI6fWHVlvsYZ23+dxL8/GF1+tmO
bBq9e/TPQtinfurFIjuJLYDEgGlfoC1/2159mCbuh9ey0VSnoyFKm+oLctvvVZz5
YKZXo8Wg6LxHvgt11PcWwcK1w3NfmSPcbe4OYSbyvdqjHUPyJXPnhHEJ83hGoBb7
cHVMAjaAhEFAgmFE1n4CTpTMpX/z7ULRmmf+ioHcCtsLnpZBZOH1DfDaydF/aF3R
gdIMy7tCFb59LVfiIieskd/CItqpoGFZuAnwEnuf2qjR+XTLCBelFPIL3DG2YLSG
qLsx4FspS5nryve0QvCDTCF3PM2sVzX30nETcFd4sEoxoxQIrefwu0OL+oDp0jTj
VgNZAwQSbGZKbHfnXXc037oqDqVOcC2IhhdF5iCieQP6bnEFS19CX7E72Jc86eWn
PWfRZoXVXukGlOcRIUMK32j46GB4l1VESuS7aVns0+3HTnvR5Uxo6nUfCKxWdB3J
TDFUyNbMKEsRsvRX6YN/DFfHKfDOadlNH+rkSoTrDBJEzXlX2iq14x/Ub7sKWs+8
LBUASjPZaKTrwQIGJyyH7Lhbg1+g+OyCM/wnbv9/EOEaAHagXhiU/8wYFjox1ZdM
0kqJxQOJs2qfMQLPw4IZ3ZNPU2JETIAoAqjMZ/FqQRHZcRFZXz9NlF15ncVLhnxy
wEqPQMHXxtqNnNd1eFjGVBn3CjJ67a0rJSmdlIaSLMqcxv9x+HqedZfewaeIQmF3
rXCafBWnaDEujRyPsRHQ5RbiYxzUjZSk1hClVDo+vovLmmGUTka+vDF0w1Tlfsel
+wEbi6Jdu6P9DCTQMY+7FEe6RE8QHsOL3Gd920kx6fQ/C88ag+mNKFffoAnkyZEs
lVzI1aUEKZXff1blUBO3KJt5WWlf3aObStAU2JWF3MJX5aJXleRYDgBHU01Rea6r
OU3xMedfdktGOmh80ch5UWgmdm9UbIrKif+8VCOEiNzhdE+w5B1f9jzbr7bRVwx8
SE8BEs3bsjGf2ddIy7HmPO/COXVNAT03cDRHYA1ERrB3i7fS94L46qRuF6C/CxyU
XqT/VwHdGWCWy4snOyhi47zjrzDw0qre+daCIxJgFDwq6JEfCsTwRmskF0XJX0SZ
GO6EbmQIo8qQiDts/7+Dm7H3W2CgbGgLVuo8SuXAt1iaP7wQ7480tHi7m02JnCRm
onGLz/cde+71lAJDz6oZYcyf6vmktxotwkMTYtM7HR9TTVObJ+dvOjGr09eFjLwf
Uq6s7miL9u4Vv5SUs1v/Xhz+H3d0a/dOBfQRuPh26t9j6z4kGDT5Tc4wbch31tfM
H1rqyW9pbeJlnRc0tQmTORHBYcNEGft9e4TMVw8SribGtkw+Lv1YaGe2Uxnvzl8F
x89cKrLZbzxSKtSKPqVv/1RC9W3Ynf3Ic28zq9Qc7Y8cvBKUhdHyI/oewGT+BiUk
e23FZcOHlMtRo5WdHvhP5vO/rjd5s905pPmG2/Ky3iY85CAcLpXjyco5yboxFtoO
OzAPH96CPJaAl5RwCmdkPHJymMpQeBMaiXCQe6kUFoAFEuwCE8JjZbKHkCz7HCao
9DqyUcCOiYXVV6TvQBh6pUIS3teM7HxfgU5JHRAiADTbWm5BDzY/8H1p06SgFcoN
aB+3dRBOw/peYub9eviHd6ilk50I9s9zlpuKP57Cvpc+6x7yFzBjd438bSA18VFn
ymmV6SDTJkMzVuVrIYWiGH4vB70WRPIeQfC9EUEpyKbdBPiIcB4Ah1PDWp6dqFlD
x/JGvgsAjlPbO57jXxi2+0ArkNJc3U9aZE3HbyW69++lKBa5QnCMy4wvuynJcM3+
4Oz1CmA7k06SkDGBAAwQkrDml6lxxSfYJQaO3/Uk0y+ko1W895F8iM1kFMH0apnG
H8EprAB30x4oNwB1hQtGIvVutdyxqqGLXcsZLdRzQUjoZbZJ4F51ENGIs8EKL7u/
qrhlljywfCr8uAjU6n9K7xX7GDhpf3VlkM+xnP6FEPUgDFpFAkMHleYhQjW2NTZp
letr1TC7p70wZ1fyL5LRD+8V+tYBevNs3EYihTU9EKNwhzZZABDHiTZvLcKd6fE+
/mtcbZbReyDMYjfJbZ2cvTjWxGIo8b2trwOpSNmfDAftXiPzFc6r7qGbm727zavA
WZscO2Muc3MUeWMCQV4hK89+TYpZgInY7qcJAl/DdArgRwRtBcygPdWBc70TJFl9
xgobEM4F1xGRhJtdAn9IfxjGY/NSljV42sa0DaGWxpCcCJbr8iX91kmCKf2LSPrM
zZBkOf/3hgzLJ9cuJOJT5tmwkSMEJWkWQE/4SwT3+ueWtTgRa8j5vGRXcVkniwYu
2A97+UpuDqxjEZOc+HUTm0XNuTw5y8emxCJ5PCYNnDPKaIv1ylTn6yAoa/KtRhLo
NUeWM8BW2DBqJRz+SBuubvDytN3lGRSRgrrLS+SNBHKy5zWeUy9JS43qG/NG5e+M
0XILXtyMQFjKUXWzCHUfvs1tWK9Pw/kn6Wpznk61B844Za0GU1MncLL2/HglkwfF
URDbxgATwCA9YtSdZj5gA9JEYiqNH0xumlqxfnajLU/Rh3QjtiaGUyNoMU5n08wJ
EnncYMIsBJpHs6QltMXunjsPJNAOX1KhGQSClnx0mAOCQ5Yaj2zObrKOt8FpLlc8
eKex3rZXG7mdz9Qq4MFJgG3xzbdzR74s6/fnv5ttxwdJw4DK7UcNNgwx0fHV7FoV
92TpszLN3ycVz5U1IrrENEDlXp+uAHxOcVgasxehg36u0mTX0iHrnbe80zMay85f
eFxPzSLKg/aZybMWPxhpVZT12h74+oppy+YtdfZFL1ejMSHzkoWjD9PsckZxGJ2h
IsllX2qoUGTvoHOrsd9qaBkq9ckoqTGTFqCmMgqFgAWkvCt/Qx7aRwRKCQCXugX0
UWcfKIDM3YSVCHJq6eHObnfAwBgDNL0VUMf867BBf+tqEVcLFg+2ll24Z5UhIcVN
SRZAjAYcaehQJx5Ekd7bHlYsu4/tPRwTx9d+1MLgFDbaFS827CfJ1kg7YrdBXRVo
n2cy+0UHVwpXsSgc1a2A5H0tzh0dFZ3ArmLtNDjxDmy5s8xTldALJhil762ku7te
VFw4SBYWTchuKEszLaOFqx3yv3DJzs9dWEPUMdvQW/FpgDyyZv2YXhUN9dcvkvmT
LdSuNJDmbahlEEQvgEioXCI6ROOS+QrIACxEkqnfOjOIsM/4JTN2OMlM5og+hfTQ
5zySNMHVnHnWroBM3MgMsSBlBcaGK7sE6qxBcI9mBFeDtcUc8FbrgThtsoBc+DQG
4Geus/eNMusZZLILucwsUMIlvUyxigAv9pqsf7jHa0WbaWqd2CnORrSjLtti9hje
Q/LzUseUIVa+zQA5HewOUSs79c+dGwis9q8xmqOp6zVcoAT+C4D8BblBSsoDfZcm
7LQ7mbWPLsFVAVr84GLLI6lQzUq+6J9njeGy49nwG2jy9oYS/Z/Uc1XWp+aRzgnX
qXekepIIROBbbDyCzUBgbpWFoml33JtFtMS0tvqDR21ylPvsMeypMYe676vHAZwC
4wfRtW5Yo4qUJrVFGYLatzmVLHHR4zyAJqcbd9Xte9iTf8xCUa7DzsrXIJ6JgafK
xpKzEW1NA1qVhpno76haHTb8a0xq8SN2Ux6Iy1dz/JumeRdxQFeUuLh5ttgH4GZc
wb8aZ4ByTp6OU40Z1FBvyNVK1T1eBDv8fkgj8QWgO9yuOrrqjRBq6TiMXD93RftZ
C5q9bZSEZrKHCbVnXyfnNufCp8Qi2RmeaozSIWmreHW2igfsTIbPh8CW7rVr2CHI
IhlBBpfbfk9XqZ/jEz5qiHX5sCOwyh8FtYiGcxqXJrdKzXvRNaO4vVUMQ/WLSmqt
GR/eh7n74Tc7Hqm5r+/XwJjNp+ASyS5kk2ngnZdTIA/wJEZkaXToeYhZ5nq/uwTO
w6OXY6N6lYRe6xPLyQZa4aIcj2gwaiGJy27Me18njTDM71e1ndJGEy+ykS+3NgGj
IKsurhxkD0hL7hs86y+nRCMWSv7ET6PgZgz42gGx+9OxvNy6pIJSfYtiUPZPtozu
Huoez0G0Vnq/YMst8MegdlQB4p02wnhqmRLZ9JMF3+e2WaEXKopDGn4bWdcOgxJg
Y+fgpSo1fR3D2PL4ktm2mIHdX6VLCYFsMsB5p+Cz6h7StM8Lg3jgtU7ex+uZ4ltu
YJICi1rc0HB1OMkTaL3uq5LwM7jbYiwQwA+RJKf49cScVOGVFTm01VwaeSDgC5nz
bXr3QOxi2vsQYBt4E2VVM6vuqGbaul1JEpOk1CPDw2+UXxfAVV8s3vcHvRL0cB05
T0Sqj7iHC+BV68FiqENK57nGb58tTxWO5R39Cfhli30eBJdg+pinpopUO7FG8p3M
LMZCmKBR5dk2SmDJcfmF4JfFjhMDTRTVunDutXBASvbWBSSb7WbWks+IdmeeF8oc
mrrEC/Aq5T12/LvxYcDn3fWYKgTHwVmg2Pi2gBF5UL/75AV2A2vePouc56nzWR4x
AIZW7MfN4Cffiu4u01w4oVxq6vNf2JX3cR9KZBN1Kv71KZ0NQy8+9Xl5vyUD9XGT
r4AaX8mh3edzEa9QMzHp10IIGA/n++V56NlDPgoL9KZDkwUzQK5VFtX84FXTWQ+m
3cA3KmmY8x8iYeg8XRZh4OmkQY78p4SSWFkqwBivBGeMe83L0XNxgOeUwIw8AdZI
bXyD6FvjGaqlRUU9BPiWzA0Wlvo+Cfk2FUsAmNkauIGKqgg3HZwiUS+PbTA6AjZ5
PYMes8WRcvcGfS1f5eFmVbU+tdYMHM4Wfvi9e9d+DyScOMUURJe6PGsndwQTws4X
0aRNoIcOaFLB6jyp2w1ZcHcos4F30IqJRhJtaZAqOSemrtFneRbOuEzvgtk6UHGl
lVUxVu00wfD4Mfem7y4DvuBviula2qZisME8WPL+j3JbMHlDhPQb138xKwST4E/K
bhwpnnZnYVov+v9c9N1WChTukEi2mi9OVUO714+Ijtc95CHgnmhNPM7MbgM3s4AQ
DU+xBExcU1xvs4a/KcMsikhWQpK5Tr60+qKH3KUp0gx4udY+Y6NeSyh+aPXDmOkN
19834V7zFZy0LoPvStp+pNhTkdjEZ4KZ2Vw3ciFcAnfAlfjgaYV5jS5IhiaazGZp
xaP7iUF153URH10wh8/7SPeG0/7swqewJ1XUuGc+3HswMSkjeL14z+96QKi3J1VC
pg9agluGTYzVioo24W9sHFAfSQDbz0QcheOSzzsIhRPYWrfL9uyP/SStpI/6yCks
wS72OI51G7Yj5QE8qi9TBrof13XZvX8lM1g/vW3Fjals72b3oTq0kizrbmvB3Fyu
QZWCjkDJyh3IW2kv15Fpr9BV4PGaN/QouSz6DUxEG9RZykHNg03cQ6F9Vda2RXnm
Wddc2ErtVsIOYXSTyBEQ311LUpUg1eziLC2PULbGNzp9n2Hw119C2LnbqixO1h7I
KrqTmu8Xv64t1KxvGThl5LlQmWI/EE5WuUkaRms9ftXR7t9MdMM16Oc25uwPD4vw
3TxKE8SQmPA3Wo3a7O3S7UZXZSslQxanuZTjRUxJSMT23Lc6bxXk18n6UdXdWs2I
FZb4puJeOIOpywFy1IsmbNKFfvHoz0yos8x5EmFght2iceSxCbE7/Trtr6tuZWAe
6M06BSnI0O+6eY6quSGIE36cXUh1nWCUy8ZCjYPE7oXBrL9H3eCi1S9x+sCEtfGf
qSDy+CVZSNMUdyfFe/DnanCn1XlvXdmHWpcGOVSxGzutX3BjMJpUYVyyC5hAFx2N
xcXoGC2NLTjEGSy8KrqpXWft1C+CBDSH+k85Z8jJxK+I7OlneGdY4K5UE8XvlM7c
cIemGq+9Nsmt/3hl6/OteCl97/VzSlLP/FasXP5bW6w89ny6fZ8A9LhILqdctdbJ
2h4DcDeUHhyHEr5uZ9DXpyx+eKfC3j4ZSnS13RN92s8hDQuU2kwApgce6mz9Ed7W
PPhaFh/FvOxqmiEd1t7rmD78suBWdJrZbD5euf8ZA0gDH2hUnXH5OxdM10xNeFcq
Jwnr16fRGq9qQBwF36zgCGLoYexPmgNuOg+fcbJSwZLteoZrBoPmuckOTLAeoo1f
du7qDi7d2WWMdPYIioLRnafZXRBX86NaPhehs0UqRTgg7gnkz3ILab+nIRqtg/SU
f9zfCecN/5p5PTu+jpT+vd0VwTjm2YvcXbya8wF+u77uETY2Yn0UMIgyNxb4PgAM
jFnX4p9wyFWCBmIYbnmyZu97luglnZNj2WlQFmZVSTO/BQDVa2NmIZOvWxVl37ue
HyTT+LEGTXIxchBOl7VtsUhc/CPN6138oJHZ9Y2Jbil5Zpo1ZLkjc4sSJBemuYjU
kcnSN+Snh5yctOgHNuhGHENgqRKX711/dTxx2IFmKBqvTLpiUUGkyPMm+3qgeNeb
aPXDI81rWwI4wKF62Q3jCpcpzrRPmpVSNVg0pBiW34UZ4BSj1W+U1Ot9nWLHDkU0
bk1P8jhYXCvUCnKkAl3FDHU9/E6/Ce+rtPVuzQTXQ75UTia+9O1t75cwCQHTAbWI
9cjzRfYM4nKmmaM2ck3f5Zw22h75lGHqp2kGJ9wCG7C9LyE9jR4k7DL7KMOLk2pf
PMTI5BlcAAYRYm4JsJRNd077WVkzNBQ+GaI2px3FynHCZsoblJLPhYCBTyjrWre4
M7msEbQYcRH91WOSS4983TrkT60g/hfj9iewSNDhexNmFu3nzCl1k/p1eFfDkcEZ
KjDqNie6/TkEuzecEzO2cG2Q94LXvFjn6xgovgfAXziWtDkLns9yG1eT9CbSNcmj
94qo6WZAznF0reBluIuUVZj9DImjL3is7du6zEKChR44fMN/9W5WOML0jyQUxAjp
hbHJ8JqDOldiX+bZE/pya8ZXKY8DVCzQZca+uz4uiitHONsvLZWeEUUbj55MknuW
g4Z/4Si7myhoTbtJTUZOVmHxOOU2yaMIcjnYbxinvRGsHQrBx8ioILPAzcLamG4S
mwJRaTqE2s4AMcgtS7W+4hA0laKcH4DPP2KNkTXcFi2Kk6hRW7W/FYaQ0tv/tzaE
h50DGT5J3jN8jyd8ueiOmi0Nr9aBfuRSJYAWC+pQYfxGgdEXku+INDUDEAFLtwra
FkdD7dDMoRNfTQNVKqRRgPf+QB/4emloeBXoyG63EoVIV6Kgt8C9qVC550RQz2df
apqBHulFM73rqwg5uhlWa66R9DQj9SXBUtnBYRH8LZy7ktsAGRe0HWQQ1Eh8RCM5
4ciGRW1UyNM/P2DJ9BAlBqBPCDmpiY9+Bbd2HhWV24pPeLXSOrvgk62E3K4UASTs
cWmVOCGRV120yRkHJ45BFpOFx91pEqm3QapT59RgUi875dbo2svZgiBmRzUqND0V
hdRuaxiMUNjuxwTTROYf/QnbBgYAsJn5vO1h4sxbWswG1LJfCAT7yg7rl9RqLDOY
QLOCbzakmGgUZ05PMXp16qih/bkMuH/dlPRru2SkdC7YKOp7UR4OT5rgIDob5JCW
b1eIPBcZ7/MsOV/JM/HIu0Fav1KxPwsVgCzE2M4TRXIfs/+AjBMvNG6MlJBM9Fqg
bSUzRwbOK8iGCO5c/rw8Il58r1mJWDkoVLaEsKoVYiBo7JGNNddom63dymf2MoSN
z8rmnEJ5E0LVSwI1oZrBsMSWiFJgZMbsZ/SYYD2U+bmOCyDrrdOM2hgQeARiHQ2k
mGgXuEIK5V3eUIpuOb5hy5ZZJ+5D7GDXqANVHIE3XpbT2QTbq0t17K4/HMpgsCoq
5AUbAvtvm85gbE8fUwaMykfAVTGU8umAGaeCZzvELllZuuXuDdUd0Ti8s5AJovph
sbJgC3Nd1zx3yz8i94/uIKwyBif3sj/hIpQycKACksH2HX2Q51Cjdzura9x7lSgQ
oj9FUtSo8BHpsEK4YcTPTO3EnY3cSgW+T7prD0ccG0r54AwlHaCjY5qiEhA9j0Xo
o/fTaYfS0IWRu3zYi6Ffhi+PhwD6f4uvupoUh+O816iD6q49F1OXk7LhtiLXMYMv
/WnFlDNDCEJp/p6S84oqSo1+VvZASL+dFyEQdSjMzMfIzoL9N0VS5Jvj6vll3zZY
yCnloywjR48JTo4OScDbFyJbE39uR4pXKMJthHRxeiIsULjgTA5B9kdWP2RbW4Gy
bKFDvpEgGgr68EbnlOSbV+4VofZ4ppH3KgN3/nJ2RUZzT3jVuDJvVUl5dmqH/2K6
XQsG1qJk9+pB+H1zWDxxyVnXMr3/OPuweFw2J05bY+fyqPEq6wj4SDjr6TF7btbK
PDlelnujtnvtM83vMSa4aNa0e2ETGE021JT0/4Q3tafugTfWnzS+y1sWUaY1Lkz4
r6l2e1Hr2wqkPLryI2j4RBC1snffWk8zlnXmV3hHHMM67aWQ/y4ybKs18E9zNA/m
yv4Hoe8NetiJGaOVmq66eYgwpehdhdIVSEamMwoU+j8UYuPaeWcOXTVcUuqF/6Du
QtN4VF5LweIodnseeIHl7g7SrUmYNS13/jhziCmch9C3PXsDPqf0ONbGtOZpS9r5
T4mJZ76Fq1vAKEFlqSnD7XRgZRKjLxY31lReC6fMU1FdU3WmvCnVXsgBxOd/cScp
F3ovneUMTSLGZRPcn/TadBZGbrWmL2kWOuQ++XF+khxomP4jneGdk352khXfUtk3
9YAR8iKp5aT1QcTPqBJrG8rBjQg24q3lgqzghKSx9NisZ+OzmM9Zb+YFCoE6VCBQ
oV/ZNw+37qbfQNe3POJiquA7S5xQgbcj/rdMnKee8YRtqWipiZqFxRW783AvDojH
5fhQIW1pJqZxluERb7iyUi0q4unT+/ouZ23oAx7psQ8Zrb3EO85jBC7gUOGwMLzA
sSAjSwqv9MU5ewKEuPlmI82ZvdP9/ICG6b9WCy4lwGGKiTJ+Rb+rH36Tw3mT00cm
3Ac7cHgYE0m00yZqY1ioMMmhtYOEv7Of7jbBhnMO6K3jqswdQ3dZIggjey8cl9Ol
6CkXmdJkbviCjc+nc8Mk2q00loTnE84njFsYCIwTJmn+Jowsu77MspR+QcNWr0k7
qBks/cjpMNVQFNC8aGa5zMefOk+tNUv+z3smqt7F+9DA9/nJmVkPlb3RL82AkIn+
7qXBLVVwtqb9WF7/s/QvBM4iadkTUbliEPmSJh7CBxFW7up4xVuTxtNKkJhooXQ/
wbe5KKe+RAeD35ennZpR5zh4s06t/ItcygWcLZh4YdLdCs48q2I4LcliNHe3nEV9
QrrTHRV8iJzpzcCN3Qlmos9kc9sj9lASIRbv2bkJkgXgXXlY6+d2Ee3MhSGfki5n
40DVBbCtMm9OjBYmYSG2pEq8xxtyY0vF18PIKTaqsdZtQuh6WEEPXS7PgMKPk12y
/61MJlPn8PGphpXwyJop049AnYO4e+Sz0BA3BI9KW3pxyF4Ks79EWQ/Xr28a6p4B
U3o7sJvuZfsQJfzLHryE0YC9TNLwJuXEOeuGGVJt8gANezPvF7NU9b2F7/fLSQjZ
E9QQRV81UfNxa3RDQvHoZXPHh7cwUDK241u9h/D6kksQnSjFErwLom6VH3nt+GfD
Z1SseukrD/ZohUBvMdfhmFHfOlnOris7ufWW/JWWSlfchjy9fiCtt652SIjH948E
3lQPT3o5lm5ZYh+MjhkOA3cKYx3XYWwKX2jr9CZQLMcHOPOfW401DuK2eKcyX6iN
CoJurLslQy/8nEUHp6nC0cjCft0w01fgkfRFIgf9yTfNd6yXpLxhbWaGCNnZcHY0
MA3rxBaj6uAN/VAmCulxnotoqhyiK9s7ePrsVxK8tcsw83aFh0acQ8fT7INwDpY7
QsN2VwaKKv0Z15mnBQ4fgPhr146ktLtC1R1ROMD/ZGxu0JaptlBsnlVFLsHQqeBt
WfVANPyN9uNA5ViGuYd/ss7NZdF1/3n8qcpuW6RCmKeh/Pb0X6vJiw20pATNWM2I
r6Wtf6nISZNGtkoHRfVopWhX1NK5UCSj9EDYjTI2A2SG6VyvV+eMfNwXITQN7K7L
MUIYptCqgLZTwRGv1gzUxOek+jyt1Ptm7bhlOwC7kOlm7r+JvW8KjttoNNQEICLc
Us9ru5eQPeXwMVhTtGu13x3n+Y7HQYYO+ex2lrCugJDI82gd1SjZNbKWsRvay6WR
iz2IaiSizOVJPp1yaa9VgssulvXG8Hwjdo18IkizFyt1zfUdmQb9iR4ZwhrbPRQx
u9n5Lrht0zH/BIE23UaFRFB5yBdBsTkqwiZ19ymFOVuSxmGgOBaCB9mjtfyEXOC8
mYhv0P/FN3+RRPC7AvpQPhhSjC8cquV7T49UQ6qkNbl3UvwBhjJPnxyJayQMC35n
OsGgbJMx7svWWh6H05FAmQUmY5G9U//whdgg3tBSMA/TzPF+DDrYeUoXbPjVkjIS
vm1mJu3cbipRUPbHOFsdA3sW6niIfNJncj/6WFOBgOtnBIDbqDFGrehPThEjpwBs
1lR3uiZnYtVmtka8C+C4OVMQFuK71JPyaxbO932ROIilJAMX9+jukThedrYOuEDD
aGJIk5U3DWc/6mOpnPaAzZCxclnnlbtFhyrJwmde3rh3D8swGU7u/oQfoIF4b8At
KNLprnUu6FTF3V/1llzqohvkOnT0NxSd51KNcnDVQ7eFSEr+n0BWWZFDVDnpBsLC
jKPb0MbV1plQFIhu+cuiFcgaSQBwejm2rCeWu3P+8EmSxqxlOx1ouVSEK+XUHSHF
/3BfJrjnxEaNxGgQiem+MR4BZKVyi0pOnDaDtfDRi0jnSYVu/cqyvwgehXIsS7+V
TK6/dAq8ORcqzO7WAKE7wuBrOXDljki1tO/Kqn7gjxe4EMNIOBxZErMo2/2xv21H
NrEZRaIur+q4D7qz+vgmSM7LmJeiNFoVQSPbv9oE7Eg3rZ+6kNH18vK0Hl1CX87a
u0pb81ctQx8tzzCP1LUhTKSrGAnMw5MXH7SC2RlZUx81MU30NUrGbxEld8RCR+gp
FJgkdiQpDnB4HwPh2Xdw3Jv8Vf7A0YW6IUQu5ATet7UkG+DIc1LKvDZC0h1vctD1
+z/ibDsfmiOKniUNi526+BoQiqjIgJ0Z/Ae5o6DJfAygAMnig/iRr8IAu04Ox4MZ
LuuZri49W4RcmxGd3mGS/r+10I3UgYq53lrxt00EmOpbyGfl4nChyrY2jg9GDWDx
7OSY7OHycKcsfA45uy3XeNXzNn4Inm8YXZ+W61PnZzS75YkOZQA0D/liciksmIJy
/tKZFTJgXWVtpkqY40f9JiwEAftA1PXOgXx5X+mUiBi24oR9QCTn0HAMnL/1Eja5
C72xfuXPGpGgujQAq7gwKqlZRLjRZgU5sFL27dR0MlZZDOFJQrQD4JIlxanEf8Vq
csLhCfvcKkUekwG3iqdYOjFO8cowbgvFXZeEqX6A0j1Bpc2AUZTKmF5jdy0dN2EZ
MAhkGrLFX6UDFXbukD4dqHQNHF1OKpg5VHDLUx5sTuxNSBkbyKK2brt2LmfA8X6B
eBwU4R3uvwmntQC+o3LY2XQKfgATSuirBLMI2YEcCJXybLT2zgWA40hka0stpcYH
a3SKVxl4smoL9rKun/gL9NuZVNiy9xXXYQ4fz8fC48KN7ODLRZ0ILcla5JzR/PW8
s0tBgePzBpbRyDT+7SjHjAzoUTigigELmEV3nNkUem6gKfgTXeA0w1ZlnAJgwj8B
lvBQdi+Za/LIhmFenogfb+4Oc7JgWS4GyWfXAuDE8mQMYft0pCqpu0sr1EVSzmJP
6vkvjOcXDPvKKpBjzpQvpQcBAvZ75MXta+YLO54P5nL+KpYlZJqy5nbfFEtapA79
IGMMPqIjgv7CBr0jtw3Q1QtCZSfcpKh9ocxO2GV8mCbIk/7SoviYtTbDybs8RsT8
T/pQoPQeStF7f1RuBL7VZ4Y87XdgLQvnJ0ayIO6BlBUGQmAw3zTJzCi7ycjIH9as
o51VKKWlN6L08MKQi7RigKCpwm14k3pZ0rMIQFJUh8A0J2jGXx6WR8fQnl2u/cMW
/Eo+XMTlVXI/7aZ0uiHhbQKA24d6dCvidMfXodbxmOiCnp4/YgugPD/MVqkOrTzG
5dl1e1x3MIZGUnVEzGZ9bIPWVWz3Oij2VGZsYqnwRxMku1VqhthU+byzsvIOH9PZ
QRIi76Auig1Exv3oQbWDoIIsHKgupLsnV3BAB8WXspf1BrlfJxcdKAHIjLucAJBv
H9+VY4C5N4W2eLhOeosErfi4k37LXaB1xe/3j4FHQwP+otUuLPxqJMqaYNYreC3A
/IZnOVYRSc2+y1Y9c1GS0jYGRvD/Q8utSclFX7Pex6RaCylfMU34MBK7PdBtZCfg
TK4V3QVjVjA/TbvvVO4OParwp/xEvBO9KJEPoKxYqldlXh5ajma8PeK3QRcgJJdY
+0aHDTXXsj9Ze7yGmuiWgK+r4ZUY44eAd2w1Hxiif796VzQk17cAocYdeAtGp9nd
8SMvBWGmioDrIbMwuDsUK0Ovv9KTLV3HlVIEOOjTnC6saO7Hd2kxuX8jZfZ2c8Mj
q1DYBqO8DLFrMRnRGxNA8U4ckiGaxZuI0DJ0kEQGWbO0V+BlkBbLiBo9lBzuxip/
V1FA+5ed5uI7zGK0P/R62IccvtDtyoKL42VT6dmvvCgiZCsSFrGTvg4ts7SK9vdp
PINtavc5XxBVa/mup3VvHjv6eYcwiApVbZJTg25GyC3RYPM+62iOOGDF6zBA1cKL
csnwL74/tlkKgESkZokiJ0F+e/gjj4+PhIXfQmaElKkmsAsHk7jK8vMOyyeoXurK
VKW4bnBukegbvVA6MOeo1Xdw1nB6tGV8oza6qV2OYYBCwDeVFFzJNnysYPhlwtpQ
9X2MO5OgJrfEnPND2k6NavXrp/nT0lLKRuvCcSMr+RXxIH9Ltcf0m1/N8RJRbLz2
IDm91DkhD3ElogGPT7DbdJSgQYD/hmDYHJoBbrOQosJ9XZOFk8yX7S2tT/OOGo+g
yfiTdqflKYf//HagR27EKOtxS8tbBJkuBNAOBxqk0te8IzGjidc1Dap4IQv+yrDt
suYM8YPHZX8P1gQWMAVouEodwkxCxBMm4eBc1fRFDZp1qequDqhdcN8/wcyoD1BS
Zotmv/Lxr56JsNleu6ZHBrwaJea0Foa1sYvO7ar4J5oHpje/N+u8nr+Eg+sxpgTC
PvlNyimxpS7j1Gg8dynRRkrcXyBSSxfBZo3Qhj3xh1JkDF0lVp0xRNNK9cNnUTas
h8WIcHOG0MEHv/PtZPi48D28eDlkDbufy27WRkLQ871C3EMilOcYwkqVXXF5seRB
SoZ0xmQOZzX5Suw2WMP0YQuhorxHrh5XAOJ+dPLxZL3S8fk1vPw5mS1DDPJ2dC1T
qSrd1rzjublF4xge6zDjfqQ2Gcn3lC8NDnviOXu6MTNinpabpxbvAiz4+E/LBVmI
G19SzDhtis+j3sQRjjpyntFu0Ijw9sFnmDHng9pLD4NtJyaNl/cKRbNlEKnzd54u
nZqw9GXXB9yQkjTbbWsddCbDTip5Co3dr+bYkiOKjoNxe/alqqljTp6kNV+k5Xwi
4P2UREqztxq5VAOwXZlwoO12kEDLGNxlcHNS/D3C5DPxmCX0twbtoJkDlNGg9Nr/
xuLUdGA00g5qEPMGJgMg+xCOQSuZxk6Hjy9ioD6ZA9J5M3ohJ9MErCTHD3b6XiQG
JrpVMksYmc9RPKqvonA1y3hbNilXb4c9iLQ6znYBTpDST06eN97B2SACppLizcxx
EkA/vcJYKb2zS5c4swRptEpgcIfezdMYbjn0RjTr0ziDv3t7VV8C4PeObx52eaXe
8di16FOgZaHwTbl/9wMVylmmzXkdajGKHH8YdaLw/oygZRymYX2C8dlnaP4EiPt5
MNfluy9UxwuDQYizAQ8sN39qrIXPmvPuLIcBaB/uCtZLjMa67cEi6U+ah8QUvBDW
eKsKcjsWLY7Eu2uszTl4tBe0OcbGtm+VAC+qoOiR7uojCHGAz1FKmmDfoSxnKXy1
H6DC5UX6MCf8E4e0tPQGbR8NxT0YzmIdSqEZoDPZS6JhDjBzctBRdD9P8LaAQKF2
y53gVjrq2dlRzG78VXC8TsdAM7w9t6MPa3RtQKYrG+RAKKVma7toALdLWivlVBfj
6UDSeShylgZGk3DSOhBAiSswsstq318nbaimfmVxfcH57z1XAKQ4W5gvsL2kwOYR
OCQaaW4HVrvb3a7D1W2UgpimOrry5mTPtAxjFRH1OV+3jCtseA8vcwhlGkUd72yD
GF+RqWJXeTOYXT5k46HzTrsHzPdsQPGhzADDgVbsZHa630UWMskdeFCDlPThenxv
iJ50NxTODTUQAMtX8sfR9Dbd7oEuf50DIl3c1Clqaox9AoXgQEDbKWIOkp7xHeVf
YLsMphpSXjE1+ND5RzgeAVUtbZgBypyf5usbjkNVdj4IjlZxXhqNi71lQjxAJUB3
1gTOIrzq4wKEGXaNyejsyIXpxtk/pBMS6U3uAypVR3h+ECEPkDakH0B72rObvESQ
W+BwxC2Mj9flrikcF+JgJ2ED4v1CXB8qf04sBiQia7dii0h66iOYpK7Tpw0EF4RJ
jW2F9akGaooS05xOx6GffPmvG2z7/ho+hq9Iw6TBTVDv24N1T7ChZuc+aJ4Wcssv
CLUE68ngfYTUh8tfVeeeCd4Na+FsJ6+UcF+HdVbDePYL/E1Z4LA6xW7qLz6Su8kS
eT/9nCkcKHANueObDcSqqxGzP15W29cin5wBvnz41yAmTgh14Z9OHuVwGvgdsmfg
/ucM7kKJJpEzU+KTF5yBuMb2Je/mpDG8nHKph/c61qqIgGADJCo0pupaChgqm3rN
QtU3DeuvxzFjVvSYLaMjdkCJvt3DtkCSkbFPp0PJ2UFmGu/E9RpcEZtCzffx3w+f
JWRp1CsjdaY3v3dPs7Pz+aRTNkOUp2tVr31CwpMYYHHKZhyGio2I79BsjbsWxsZQ
yVP8AAPIPmvvReo5HfmErGfvweHvgytBVRge4mBGME2KsCKYzBRJu3s/hAd6DfqM
1FqNhd+Zn9UGRAUOSnn/seJkQj0t839apNeZn/tYFenmrPAi8Zd6nxT6p+9ux6DN
Q7REgxc7YilFfghMWdd90l+K3FaVp6Ixgb6ggEYnpL18CKeuoH6qemmPINO6kPmq
tetDUr+1jz3CIdsivnriW7Y4NFp5R/DixcjkcJGieMmPu/0HbUHOX95ai5gqQ+Ug
98vjW8VxPDw4c5kKf/qWCR5f0dGO1d0BLwmI0qpsvatZzmlhZJQ3xEqKwrDUheUe
pY6T5d3OyyvmEibGrqWvk7LFRQ5vNiMMvkk8pWOZQ2vu+3hg+O6XOsFL+4hG2Aw/
t6x5K03CYCKjDz4h8Q0xdQzVwhyEv6i8R/31hOfk2/yJ4XVESB67b4Zq5z7AHgy0
7RkxL9Xbb+PVccK7/fmlKCSIZNLUCFwXBtaG43fVfkN4xY4DfarveXGMV6u65lf9
14H0yfbk07QtWIm22jqe7eDrAHbpJGQ/3+SgflJbjqI3mILsBaYwWJzqK4+3Qs6S
oDKMwO5pcdBeBfJvYQp5/FW5VajkmBAQwC0CtRWnNEUNPjA5zGkQKJ6Bn8Gp/bAa
VP4V4dpwvDtPgw4GveKqZXlaOCzwX8M2rqLHQjkgvOP/IUiED4gRsOewWipmp5dl
LfEfRoTIV9slTuye5OqOEpY04Dkd34EYvHLTcdOgatJN5N8VCgxG2E6zYfqDQQfa
CJEkT+0gChqhIAMI29icoGQeCa1R4oQYYnWkjUUa37HWhLn7qzsa9hq9P399o2QI
iBu0iYyh0Y/HpH7CMsIwaCwHrQms9cbRL1CGDG7L8qxh8IUqeeKrT+LOKciTs8QE
c8xrfftB7d/vDoP6yiaMdu6VL16m+472BcXtSXmREXAROt23IpTWLDYjQbc4HuQN
0F1znde2xWgEBtUL3e80CgJFzXr5IMh40uGNDSOwrXrmkm1wrjAvK/5nuaAA+I6d
RDeSg7Yx69TaZ2/vgsRpBo9xCkfGrWWzkeM0VHpMcp6XL23ehH8uWD8HFwsXQdX8
+dQFpsmLgH/cBVgesSbS+NreTO3ELAtCkN8X2u9cue+V6hTSGr/zjqtzIouclErS
u2Nh0thpTN634BfF1DxViDZk1Khdas6nbB/DbHu94R/rvS3cRc2mJUagwJ/0+YiA
1ZXxUt82jsSo55B1WGG10qHXP0xSiUWU0BWvW1IZTtGwmm/Po2aGjhSEfN6KvPhi
JRn8o5GdMx+BvXBbo8mDHyz38HSGDVc1o5Rw3Ua7Xt8fLJseSS6vdepPbL9/IbzK
yFUpV9UMbs+GBoLueT3I0nAKqc6K/KdGVB/y8HscCY3MmRW6R42ayNFEXXQO2lsI
KeVdx1SMvtJAx8J4yjTsyp2HmvJ3BiUkU+6MsxNV3eEj70FG8CAYJr3Rbu2JJO/o
S7HyZdDbqvPNZX3zKdn9mZO+9uBlsidGK0UiUXbMw8tfaVw7RZkdsvR3BT3cxWfF
sfVPaSrtAPQGsgOzXpopI6n08QUTyPZaf8j5V9cBjtCWGswTwU7YKADnyFV2YZBD
xJazypYI/d3LOIKASAtcHemrqM7mXGL1Jznz9JmLZrsEnNVnCJlyabUXqwZa8idU
UzRoLPTbYZt146NE7ERbuIyXVJhOpxd+FXWKqXTdx3oyt/hwnNHztKEb1BwYRAc1
Ny7fWj9opyBDbDh+8PlwcD4ZHviLJxffLVn9cP3UNejf9f5yXl21cjs3WAxCNdKU
TmXCWHPEngIUceslQnm5GNAVS0fLR0XLNF3fiAucPBqjXPsZDelwJ/8+YpjXSi+K
TDHsQzwnuQRJz4ktMiwjmufJwmyInmDxr4fYjCwdHyHLeym6HFGcMIDT3XfE7Cr5
PVWQDRtntnyf9Ma0hV4zm2dLa40+pHSxBIx2U3MOhB2Z63TA68xT4KkZBZXvlkEB
r9qplnprWsYD5rDdPQpZiDukWpSFLZngFiOVKJqFo4ln5+qfpxX8l2zVlAg4B2qL
/lKwB/T61MtP2Tj6MKt85ySama+/ei+NNvVC18t2+pC2o3HPr2j6DYtwGaXGPQz/
2tCxBxonsq2m1XkNfAiXweWWODWvS6mqlSJd5wnWPZxmgnN8+Lg7gHddJUmaRiyT
Nzq7e6GbEMrbAzAiQsyvs4sk6lgdNKjzQEi8261uyUbjD0CIRVKtG6nEYqfh+Ajz
Yb8v+FXl8FXoFFb0O20/vvMUrjXj32BE4WXmSSItatIVuMq6DpfuOYwwv8mZUFO+
vAaONLLvDd4xLEjzCpBqFPhC10fWEx64fwtDIM5PLR9CwZck5R7MzetMrnksBH5o
0IiYpNSSPn6LDJXkQV4rAISwjvZtzivcmG+Ts67dLoW4HRYo4fuwTP3zLZbgFPHv
NnRwHmB+3xsP88JYoape3zcL0nvsWG+HuXMDGzpcpKasLsAsV6g/xmlw8pCJpF9X
kWH456P5xhK87AufcPpsV58N6R8cgCtlMIztLlKN3oqG6S/TQIezPNyWQqW4qrWY
Gb0EDlS6oFYzzlAwZvhM7YbA2adTfRV97SZXPLNj0DFp4d0s3oErY4FQc+7YBCD4
PKmqPnKVJxFNXOVeCBuWN/XiQN2wfMqg5r26O0b37SgFlU3lOPhKjHdFWldoF2qj
6is7qpbxN0Az/PmTM43CgbykBiA8GXKQJGrXu8WlF+w0wr3hXLCJYB7Y7SMT4nJo
PPwCqriv/ru4EEGDr4NqabHMZxXtUZR6gRDIEWmMETnTzAAY0TEIRGfI7o+wpP1+
AS62s9OmowuhDHMTQjPtjnXF6t5s9kvKHNSM6/ZfrWX2sVd1/VokOakHDg53CwmP
vhoP+D7du4S35vQp/iRdqLikj4J2JFVVfvnIIXUh1fJTo77arqVx3aUgq0a3Lejj
mJn8fNvnuek0I1ngxCL4K6yNbfIV2lZjKOdoMNTjax5qMAzZeYaYze+L8xX4t1LQ
K8dMFUCNemd+9YQ5u3qxTq6sObltAxhiDPmgnxeLUoBX8mxviMChSAWOppBOtKqD
b5DcYLOyzVmaFvJfL3nrhmxpTVN7Q5ZRZhtHAWyIrWrrKFvmPh0IG5xtk9aLaRiV
E9f8B3aLh1kr0b3Q1camnQrIZMWEih1MyV9gY4eDSRotrCSeWU917MiW66q0LGSA
3yTpuWxHL/vlV414bi6mbg16ObZXewnlN9yfr6GUB3rPDp19Pbj/1y8Pzm9Dmh71
eRNS5aycc4QEwEMwbBcvHbjf1EP1+78P7t6PqmXYgwfl/ApBbFmF6UqFWHknUlEL
NwcB9h+33n4NqaHNFXBs4uBilSHqhzoP+EqPQkkbVSmlh+zJd86+ar4lbOn7BaTQ
DIPuQtujgg/XAnh4MHG20d37GwlozFGs42VWk/O6PxJERFtynj5zPq+u9Fc51C8m
sA6UuphD+782Qd8kKWIaNWf4qHxw3mAtHbY2PYjqKufo1FKi24XVHqpjm2NBH+9t
myCBNtoWHIWQV9XZN/sjtPx3O5axKl2GvC7hrviIO/Lftu9z+P/2MgIp0k13ro9n
3wAfDP0Uf5TxvzV5CO0POGlUEaZP+GzN4O1oAkjrabYLfh+sP0nn3/fnUHLuVD4Y
23FJhNZnORI3A3sHZ/CioRu1zFuHePLzGtV2JWa9aJhbHEBP78GnU+y9nsv/u//B
QnBoDucHKW2tm746CB5Zz2/Kie8Ez9ZejVl66+LuQ8vAMaZUAXT6AYgltxreJoRm
MurtkO4uN21lpiPkoPoxDST65KZk14sQWKYTDOUr1ZEcU06HZxMxMTS9Xr8Lf+/O
HYral21diGmmBiFDFhj68fn6BgP0Gge/p/To6gZMeacLGwvLFVyMKW+eBVxh0HGd
/BJ+QOuhvlsyMHcOka28f5dCzhANbPLKYl3+alnLSGzFSJMbkNw/cIWRkAX8fJvI
uVfqKn3NHX2jkEJfhtoIhSvhu9l/Aw+UbO2HoZY1cd78HItTQWpzY0XRQaQBfgMg
LQGhhBazU7I2tPnhH7uXg9LM0DpN6i7hzwLoJs6BrK7kL3F9lGpYoXMXQlWxXdsn
B7Pa3Wjv/AAHQNLWOPNbEmjOHdiyNDP83MP54qiUlezWEB40Pn7CDpzgHKHUET7w
Zd5GOJbfsLBOIuXkOg+KDfTfjLkPQ8tzCznrjkq0Z3FqNMll8fGjxfHtAd7EFuSi
ljJuMZab1IIUGwHc16E/fZinFhcv0iHyZ0nt3DC+/wl8n7XUkXm9Y3qKCXXHHyK5
tWRxZqZWMkSYrHLeuWXJ2KBhzYntFj/r4dyLArVTICLmAFvlrgYymNLJtI59tFJQ
pw9OGOmyJBC9xdWWG+85tOJWVe2f31tc2Mrli2as1sofzF9RpzBP/BJ3ICiKMXe3
bOc53pL/tQi0Qjr/rMCs55FzJ9Rp4sEAi9aloYRz7610G0fHjuR2lwR5n62oXoXT
PqoQ8/eoU9rwl3xAS7WDr0AX42sPHf20wW8XIsiKaf64amCQ4wZurweE2zEDbeIC
EROlE7XffnG+4C8ZjGNVakDCn99di8gegre0YJOTvZQ7t92kKJWbAJkaN0bRZCcb
BeqPbFsBTcALmBRTRuai7r4X0eCCm0oPtDBUwJ+IL/awfXp2c45Sb+PB7V1YVhG+
cn7RfbrxKaTZ5m+PF3VUH7dJxsYM3MuAQYGzLC7ZjVHDx7sc5qlkC9MxKxKab50C
6bKBb4oRUNypt7Mo0BFr2cIftJinglMBijYg2N0BeLiwLBCrzbrOB/8bWrs0GcsN
MOtB40RVpryIoOrnRddQI2drwhQDL3idYddKI53vugMH6/qUDdz9ovXKsR+6IcpF
2jq5r0OuVFHGge2+aAeud6GP1loKObSKoUrcL7HYmxoMqQNh0xcmGFKzb8lTabaL
jZOrpIWhqqotFgC8MBwemjwTzEChjgF4Hdx9oeM6pwt8Le8pNpqEKCY24o7XAuT4
WuPam8ijQNNS4yppVT3HINiKAYmJ5JskUPDq7VTZU7CNECUdp/uDN0bN/f64XqXf
mvxulhMA4zEC2/NxBwN/7pjWJM7rYbd5000EAWr0+2Ef8WCncteSp3COpccMFwq+
+OwuSW35gVZZF+FRR4ZSnz0gK+tCO5q4vQ24vsJjAFZkjUW3W8AYl8pbf1nhIp2c
GKTq32x8Si8OkZs3pcI0SvO5zd0lJcgAPqDk9HhAK7iV7TY7B2Wi3Lg3+2vryoxl
k9YibAZbl9SkGbK0adpoT0LEZaqIIN69Ke7FQOgaPUnR8LPlL7hrMr/kvopMAK9d
3pjRa0kVafBOSIhpyyom1HOEO20CNff4qCGJlKvSkmedKATJAXPBMGVlyGM3CV8X
d/rNZK8UBjvlCLlFrKuSE5x3oV0xqU4aJSxaTOQ0oSwduv/MA7E+F01bsbsAgWgf
n8IaQGv/6tKZEtA7f3uqmuGsg+0ne8YTKqXBl9wrWkccI2sqZDB7cAfwV/u2oHLJ
RCvAkyVBB0RJp4DCk9jd9YuLXmSWz9arNL8ts/ZvKt8FY8lYh5zCHY0zbtVG+y2s
otU7gSkBhBTRJULjue+HVlPRM9WVNy0rXJIJJTQ5kDvGB2y+MlH325xDXBNgc2+7
qNZgCV/GmqEzOEsigGd76OzrQxCZPmHS2gvB5QeEKk7uZYGl+cD+ubQUNfKAv1qB
NvMLSXdZgY3o8JXGQu1oG0EuqvNrm2j425Z3C/9EpagsPqdbO4wWc/AfXJyCiEqJ
N/GgnVpcFwX3as4uG4H/UvJ8l8fjyWlJTQzqBop49ldYFOGnApHwMzxIGQel53rr
hE2Vzdrx6PYJ1rxJ3aNCUlyjPdDSEMCdjlkT4tSfHvm9gc5a6wSxY2oHPdKrs6R8
yqNm6geLMFEM27HcL5C6nfZsgivFkGwhQXfYRmk1Mt+BWWsB7o8BbHGlJRidJlfr
4vEBvP6ZYGPvkZa27fVDFSfiltgBGk80/OH7ANiX/1D9F/I7cCUtonjU1dNRWNnK
Ox5V84eZRXkBVykjvPjR9AYdPRS3X1d+QxgIlEfE9R2QhC6ZRNZku/Vjmr0xHK3V
NMnWv0vRiYGLsnMOTQfYZ0h+XY98x5vteH4t0MdSJh8jpQ3RQ/NuuUyyJ7zX7fef
WIeG/6v2IU1pKiy1TZHHx1om9aqjjUfenEi33uZ7FU+sPan+V/FkGTItStFtqEKK
aVznWdZ+BQqbbINUz+3fjjqhGGmFtmjSk8FwPmbXH5O4VNtmzLgkYZcdaOLubZVm
pVsCjQcH5bjIUIE4s6hH732zTpaM5ZRpGeEC9HYDzDPjhG5gq8kA5kftVZJLaNzt
mpfrPtIOlRWkdQ7fFX3gw317knml8B9ELh8rsVqdixwtc8selgKsR92Ef1d3vyXt
BMZJlcSHZjJIfGuzIgowNMWn1x9YFiq2Pum2sMIXmsOFhKcQqt2hLUKxiK635ErJ
jJcX6eSHTMSJ+ADU/2GyK2JiUw483kR6zcxYGZ3x3+SsA/trzJyV2uy+C1Mtwc72
IKP2yiQN8THafzwpD1xQaDgr9czHhOYK9A0b3CJldY0gpMHqbuEJlRODdhans1uO
6hX3oApFzR6D7GWPkHCC8HF4jBhriuOL8ebiqdm13aEYkzg7ReelIiKmDl62lmwT
t3ALZY9AoZJBOucez7B3nJ1v1Y/A5NY4Nd3ChfIG+9YZLp7RW+vF4/AVLarjtFnm
J96ikluHgZ5fd1/OCE131EtTRVXJAO/dsGviNFJsxRvVO7hbq/75tfUpRofYOCl8
LeZ7x/nepVh24UmEzfa9ghJYH1qYUZaTjdIlOp+lVdf+hQKtfm7MiOnOYhFsNFRX
v5wdzyk1HI8NF3iHeu0vJqmnF2w5j7DPy6bEdRhp5WY/JQMe0rHP7jfsiEktF5aO
tr13Tm+alWIvi7TV3P9x4z7fU1wLevqN2Zk7eWSB7UvJSypDNWqFo43Lj4OwJReK
Z1iENZgP2mIu5Z3fi6R6MDG6E8OWHkSgJbTm00cnbBWrfqiKLwDrZXiyPHjZEQyD
5Vti0ayrGphNQQ/opVEslm+TzNleVlMRwYy9Tit3FSNJZHM3XRu7/rIVyz8XGYwc
3m77bQecCuOBV3pUrz/VDSLYJtH3v6u3IfY/hVBEBrVM0jFWvaCGHJOOS8GnFHsl
NIe/7JURB6RBC+c0iYSUNjbiKz6ly1m1DN0OMrAJCkoCd7LPdc435oDKSdroFuiy
UVRoBqX0A22s81wYBZ4di4qT5jZhT7Vx++3h4VVPLJm8yTInRrlrC9kZw03MexUV
dBr4xqXH2cQv4MPl4D+bBQsr6AyHxspM0k5FBTlIIIBZjcK4l4c0i1V2/j8fB709
igie/80VcNmxUDeBbHJW8wNdrKUTC/jYwuKfhkotmSNrJ+PnLEhnVfMu6GzgTQio
yKfiQfMMEcpGgU/aVAbIOGOSZP7RZp7LxjA0W5J7XWNeNuOULqXGtH67KhAHpOcJ
6cBcORSM7z0YPMfBeMEnlBND0cs3u0pQteEgPK+k1tuA5L6CI9md9//G72/IFDtZ
6p0axZdOyRPtQLgETmp7xB+C9RDkSLFM1NBgrCnMb8/nHsX6bCa8Jz9MKuHHUpFL
+/dQIWSBAhsJiQ0rikdyTsNomU6j+LQ9eD5V3Jb3ICANEsT1rVTiwW8f8H5Q7+Y+
L9Zjm6mNmL94uYiS37zMg8oMCHgnRlKFSMQfycOr1DPFys2UNPjKOxzAJCunWCrT
GkRAEGuW/0TcRuDJTiaiECCRg7c1OZrHd9ZvEV9XXpHTBbN4FM8CJFzrKxqDfU0V
BDhVUCuVFhuTkI2abMt1vXIaqxyPW2IS4QJS+6gZ+eVSCvKj6voRSTvjZoMqzPvo
yUn/bseys4EEqYJ+hnvDdpVquuEwAy32rIg9rZg9lv1sx/SlzS9FTWxRw78rtgPj
jT5phfJDtmpB1FT1TcqULcBTgtk3FeRwvExzNwz7MR3c83U6i76dNLYhv3P0BKjB
0+rCU8S+n2F/Lwbz6zgLOPYP8T//Ia1E20nLKj3dLMyf/D2DzNICitxHP+T0oF/e
/ZgwJtOtht36pVhgq4tpIv5yy+F8W+UTORY1qUXlJSgtGVKr82zrdh94IaCD+Wwe
FbzNGTBcN5cz6DY6jACB9zgLCFuZo2vHYTejgepqrCrH61qlbvFJSdCL3y1KFGRh
w/BHWYWpGzexP+TfaJVGnaxtG+evzVJI/8e4bxXmK6cIwSRaFEdgJz9Kxn7gOJd9
i1KovHL93HXcZD1Veao5cjX96bAq36STVKuNCMpXCOm30lgbsYn3lxFEp/RvMNq1
ISetAMCskuD80ZLNbefkTMAtGcFbXVvnXGjsXYU54iHUPejh4G0C77pm8rgbFKJR
jwbn37a1RV5ZsrenMA0s7AcXb5FiQM+ddjkCTAuH3B7VVSGN9pYhAYyI9eeG15dh
eN0uLfXRChb2aBO2XJQFNi73HLxqHFTwbrDr1tkZccQzg95XZQnOzU+8VTPLLFKg
H001I6JBUFtD1sbyVUW0gUaFpzsK962wuifa/R/V9+2e/M2Nrlexv4GLMbOlivcT
77wOIHaaNblfW1iTFCs3voytQUHd8UrxNnAQNzjYJtbv9rAOOuKXg1NilJt4ZZzk
igMOmM4wTJ0skNrgGOutxSgnEMxhV+N0G5jKifIAY2f6KDT+4JcLjhZHpeA2usX/
kKocN9nQYZfp+TBqOuYBIDfd6qk79e/1STVj8T5NzuRZif6LpB+qhChrVdoogqqN
gnBw6ciNKnPD5oEM96U/Oea3UIsepS3TTny0RVx+OlI8+FQB2gRoEt9X84ntyIvi
QquzJDtOYHaFF1/R9/5t2IinOBA7LVNqolUMJ3WfVeY4LUevY5dL3IattTnMfjJ7
nlr6wFRiRTBA0UscuQmSjayG0qn73cgIBtnE9GT0BFYqZiDtxHr3LJaimz5GDdcr
vvPZJIkl89nw6Ym8Q3cNSb9Iyd0WbShQLQYz9uc69I6ePoM9ncCkNmw5jbFfI/Lv
AjEXB/6kn6GqAVg2J67oryD5Tq9ypV5JZVZLn51FwpRxJAbxCJPR7z0U6iW63a2h
xjf6cg7z1nXrAbFDFdah9MPII5VpHst6/IlIkmVYWJg215xIO3PF3czRnIlDE/j9
QfKX4tIoavNlXMYIfPni0BOEWgY+Q/ScyOJrOcjoGbNQkJxk8LVQalz7WzEcsWfY
+Lc1+s3NfVY0oCHVBUzqjCvFYYUmuEp4ZjQCVnH9V4YftYdHYlYVzFT6kd+sVwKU
HtlVshzf6YsR9Rq5t9Si3qd4Sz2giXM313/XwpwtwP5YQ6mIiDh7GtkxKL2xQ4q/
3t1XLm+d9IKT9Xm9AeXxvfWm/xgveJLWXntXwp9QPN/+eqQhX2hddbIcN9E69AfR
Ps161cruteTTptLlbeJFUlTPqDNWXB/5m0aESA0fqkzKyk5MsFeVJpIQXi5YFXkg
cVAUKjQmw6veW4gOAc5rsJGTzbacmWheiPAGXPg3z9vgeY4DUr9jxbEIX/iKH4Rf
jmA9+5/Eg3LnABQFOEN389z9MNXCtayQHrYCETjxKUoBzEMTQNDhvYleLtkPUN1d
xuP0x/SNFibUGCOl8DQHYqtgZAHR39bQAq6UhHRSycYge2jYJnYzupGYwgSWNXlo
aAztmwEMwOUfm9sUoHqlfgAo4jBtHvYkEEB+wskznNzO5lR0oGQTQaBBRXpc9HPs
R+bKtJc1zktQbzRuWN7EwOEktDuZTsq2cm2lO8Nppu89gBNDCr5gUeT9w4vVswGm
cakgaan/QpXoJRqHgzO3pJL2M5+rkvw1pq1ng32Z9xg+itG3DbNjnrH1/Q79zbEO
spCUqe12b048eEe74Kw3+BEjkKlLN24/oGS8zJPWGi/q6GS2M4uZ/K5Q8qtuxBWz
39Rz2/f4tp3rbzPuCrLSaBoQdpK2h6/mu4t0XZMl8u5ERAwVPjX4pgS0UA3ItxIH
TsImg6Nv/GH2hIY04Fw26RHtGli1bSMa7g1r+EX2Id6Oe/6XAy9oT6TR6VMmxMG4
kfVg1m8WNCaxKP57XhkZ6zN2KFdTVs9/mg/anlpzvyKq2miGYdv/MuGu/juUiuzW
+W+dr4JBz3A9w0LjdCFgjfdjKfb/PPh0tVPiILbFzZ7woBe/PszbH/BCquOlURsm
AcDbAg+oWxAb44Vyt547n2rHxrB6LCc7svmfRlrOPPrEU9e9PNX+hmZsRpYfF5LX
wtxoN2FcH/qhrNPlngAE99n+uuIs2DNRg72BXQOYstJOGwruNILk38UIw2G04UKt
7m7Dm/BBcWKjuHhLOWJRUg6koQC0s463uwpTQVmHJ3Pr0JzSmc4a2AIAjiVqrwS4
wFjVE5q+is7sbieHPkT46o8oD5ngRo0eP4OILfhvcQa8nZKbMLasp6QhieQp4QoM
KOUXVpt/iZ2xQTL/DjHjD/fRpCMmZXQ6QmmYlPg1IQoshNOadHtFuSn+1DRNfK1u
2z0Kpa76PsZY93idwoNA9fZBGd8zvOVjh9lbQ+eOdagjWBOG88eVFyNAdqSlstlB
E01LXWm7ily9fuc/HXznC4GZUEZOWb3763iWr9/jSv9noWNcWQzfzyDqWxXLOsjf
WtTJ8pg/rL+ykl+btoaMh7SQMy+GV+yhN5Dt2vUqzzjFd12ME7pj0qLjdyiz73qX
dVBTMlVD6rH0S4FOhhEGiJhygg1R8j0/qNM3dnoE4kwIirRi8TG5YQm932jdo0/O
Pt1p6bbzWu0Ec30rmFxWri2BD4e8BB7bfDsymB/gBIQdzVor/LvC+IG3GIVf8dso
a2BnkqxOyvU3OOln0rwvcplMtrX811r+nTFPvjt9loUCJEOI7MlIgUQa9lxXL3wg
URnqOFxhM2PdtWJvV44QaSYKyXjyYzwQKEQ9rYeo+k5pgl9FAwDvurVq+2aJHwW4
Qv5n8rr879ZnNKe77jjBRRUwuFRXdBJP2AsLKuZqJZJfJcas5fxHDwMgH3zHcR9J
4zqfwSpO2KESIpLy70mhjrgDww01TT47A8m5YqENW1VNVT9udY7Fw60gMOe8wQIp
CyNYy+cagYCcxp6CTr+p1RU+rlcYuiaEXdvEkLpYNwXXclHL9cGmZk9DuGNSUDgD
PctoV3rM9tTBE2hk8x1/1g3wqEap3YcInrk4WC1XlS0dq6ZW9NwaXE4qj4fl7jr+
GJqgmyJkpFdXXiWJ0F07yLVTe9mt1rWnzrF7Napws7xq9SZKrgU1hjWHfhfOEw0Y
WutzQCz5S/xiCt0ml/ZAeEXUM0W80bSfCH5cAb3ETficVtiK4FFUdg5LrEFVDSke
B7qT7QR+/ZPambKR43AHrlI5ffQhL7mdnjuNdleuWn6PEUn/kFLZBGHPM8CEEFhQ
oH5lAi7YmTN4OaEpFQ271WsI7Hq663sOOoR7hNOC6C1b9iQMLy1v4biAGC5ByZh1
efeg/clfT/5th2ThZiFH8vD65SglO3rQM/KitcQqb1nbxxsr7WuWC4J9rlnHtiaW
deIeslEzci9A2ksXG3or/HZLIyXZsjHA5fC3gQsuZAsNerM1h3PyKF0Yj88xd4U0
UdQ1Yt8KgyjSvqcD0xLXvNzrRMqOJeV+JuJU+7YIY8ZA+DpSwsBKcoW7v4KMt2KK
GaakbqpkWQ+5i5bi4rCwjC8w9FlzeCTsnUPBFLCqCjKb4PIEOmyRb2GuJ2/5J9W6
1LA68ktwo1ScSmtr1IM83nt6rPRIBGfSSHQhfEaNxsC3RLEtloFrSbyitREjh8Tl
LwahBWQcyS78xoQM+sM6ooGxVpJzfTmkoRwivrTKyLY3M+EKNGyVGqC8HAFcmvKN
L/C+KKoNtKiKB4ors4feP3kUkiD9Qr7TreH6VO/dSU6UNoI00utC/CR0eNR+TvNa
KDRoOnYyqCDhIjO8q/8HREnsUZPzsT1ihSn1cCHJUJw7FrOQ0Qxl1Qw8Q4NS/N5V
2W8wu8kyQZbHsD3eCk0Rws1ZxwsqRxhoTNvld9iu2a/ehupc403DMl2kyCcsn6A6
FGcSg13qL+VlzCD4PlsFxEz1FdhFh8GyDQqAPS9rwbkylKZpGgKmD+ke4b74Jz0k
vh3tL6HdgmwVjW7GzFRjWXlalaLlzUrzvY5gA7eLf+XOL0HTw7HR9YAnaPnvs4I6
KtOCAl/NXTAyNLDRErYV7paELfIhnN8kVl1wxvuvhfgPTxWCpjVZ8vWamOg6PDJE
bDQvd0y7YFfj5+11HLdU7NzObPdffUKwpexwxoPjY3+YD9fGjvdMiofrRpxtNykA
IrNSDP8IPHqa0LQPius8sgvaNkYw2g13V2Eboaxa6e+sDwOyX7cr9fjyWY9zk4hW
3YyJhNhyHUAKvOnrff9zDlaDR2M7XTRYmwin6qNNxZYxMfm5eXxz7V+1Pr8e8KO7
fg2UpO6NGqo8YjTgYblLrut/Ym+pwk2Ol+F4Tx61uZQgcNIx+Vbgv0o9LsV/jJO1
s0h9DcyJGSCWYRQahRnfmoqfcKv+5S91cuJZcnoDYgrC66/BHojY4JRRMIi/y9My
gScdq9AkpJwUPX6gF9URItDDod5I4FetwEvTt4IGbaggsFW6+zEZfC66GQtIVSEj
/F/zgBCTvKypSQCWyN0IsKXhzzRu8ABRcyZ1aze6DFchJ0/tEjdQg01NXlpdg4ev
w13Hr9aRbS/vwoFy+NnC60a7Vnab81Cz0VtnyL2zSXpYTSF5TJSAnciEDNWtJGo+
lMnAJIGW4+BKB+sQ0uzufnfkkSrgWHqCtrWvI0QgsCI21FYFBaci9Kkn5CwYLHKN
/GCf2Pmolq736adD1w+twBKS+g82EdNPc2995f7WAiHW1juKzOLLdOPuxg4N9ROk
rS0yMYfVzCChzWYG0bqdiU4XQTw60nzzB2Gi4YkcSLrk/DAfvwg02EleTkP4vqKq
ZN7ve/3YqS9kULSdaXR0iZerDqIcb6X66dHHVLnTtj7dqzihP4VwJHD7NPECwYks
z2TCprrTTgS//rwt7y5lHYps+XP43B1dqg7TJ36UiStvik+ywoG1NOv2kwa0CbjO
M5EuhW5KqVmLX7XA8rlg2Y4CPdBJABpSYq6t/qkdo7N/MVdqIfGn5JU94NPODntn
hHyzCVQ6SJyrjnMEv5a+APppuktZA26e+m6kCSKW8ezIEhoF8ehCyIPuySWBOXH/
kGaULOWWMzlX4RcJCKqFdx9Mw9g6MA87YT8DXb8uSj8aaZlUgT6PVnMa2zDK7lOH
PjJfBAOkh77+l6kDxAt8BmfDxjyY+S7C7buL6EmhOnBF6Ve4sTzkzxmuuMFq0SxM
UC+WAUJsMHDJuTVxk+wPWOodOU5lZSpTwzp47DJF5fHbbk+lSC3dEmmisz1q8xpq
b/RwBUbkEkrzGrvUb8sIvWQVMJMRodEawLSc/ntmfHwPhxl3Btxog4ao3HKqD9d1
2eR0vBAlXBfktI5MTLsgII2+n2OgjgE4k+WyAcU3Q+VYmUgXyFuQt3w4Q8RTIc1c
Cj96+jC+VWHZ5keoFpPaDYzfPuQQIk/4dMEWwvoEkunHnfYIe2BlHvuEAFtCSOYQ
UbVjAwHVA/E/Vvf0Ku71/cR6wMQjtDLKqs4FETgxeVzajav/7vCJGl6ldyc4sIFN
lTyUiiV9vAJxNt1rjxnLsuiCKHM8442L1Cymk5MO5FcM8dgUycCKWMvjiDSrig2a
I4xYivEfitdxYMRaIol12gMrMnJkOmP1Yl5gS9JnNxbn12vGpoyM0jME3j45iMtt
wduWR8+KkaZXBRhpTQLaO+fhUhQwPNV+6ZFGe1ZFimL1b23FrePMs64qM2uy6/9o
n8gVtu/Zd8sKJaJjWOxj3E3j435pr5gSE0OHbo1cfWpMtbFuetNinACDktIri47Q
/lhdFrBHIVUXxzZdPU5rKwG3jN4w8tQdOXkmD++8LHt59m2BnfHzDPbpi6ZLjyTR
QFZm152sZNx9EEC8c2TbdzC50Dogi0TW+z5NpceEQdIs0/QuwyBlzIgEZsSAek4X
hVNcnsxrnllGKaVhi33wLvF5COaCs/Ff31ionHPUGjeuQOaArAdPDQEJ0S5lwfg+
xCgLFPK7Ox9kjTjLfK9S0qYiZzSq8Zw6q1CZp0JDkDAIjbiMxoE3IfzBXXP2CDUx
s4zLMDiAxO8QFrz/jA4jEXda5zbMZ2C4vBW6G4ZrJc/kzH/ML7OELm04GGCKIlFY
GW//zjL8frx40/rFbWPf4CLh2TJF1wVcUd2LozRf7oWNEeP+SOhh1YzLi3oe6YtT
jOicNpNvih01qbkSWkQQLLKBeJ8yvcDWawkse1rcvD3xrwtTPfNHPTPcTPvjUeO6
k5tkkXBe3Z0mf/1SG02yr6+8VZKCtGLiNuq32SfgJAc3BhAPtqcu+7fIwZL0Aivt
OikrR5HKfTe5vdbz2S3tDbFpbg2KUfN5+wXw0muBhDD9qrlsDb4vmYTNvS1hw0Sa
y9S8BREJS2Z+KrPSrA4qASS7F3Ke+fjtHajs/XG3Er9vdCN0WwdYI5PizjpVd1VW
QNxCktSwxIxhGL31hMDgCpKN3J0NcfaPJTs+V+RyqVUY91m2WW87WzYBGZmmvPw3
UPQrmtXnZMQqqolhNSKzPWUzjaCoiTuLXgnf3NTwJor3trf+yfw6Kyd1XycUPKtc
g+0BC9SQv07SH0Kle5kczL482fh9xSl7SqPlnN735yxi7jVPWw553oflfdPKNRv9
1fKfCrMQlW0y4SPz9JK0UtIPmevLXJAOKSLItOR37eBmn6pr7bNM9ESTpwZlk93a
j1Kf+GGrf6RF1mPeWwjvLsouWdZYIw1q3MT0JbcoPzhwk5qCo9hx8TRTU8+tx5qf
1Nr3bj4k8Cq67OXFcN/6VY15VSmbCz1E/9YgctaqcFbeOkd0CC4MNlD2DO8angJf
ENYW8RBHoVP3M8vbTHSbvw0mzASIJZZ63+MgOy08X7f/T7eLlhOczesfOZPbzTIF
5TphBl+G3uj//7KIxeufvmmSOm2zrBYUOHzVP5BcwO6R8iSHHEmpiZf3+W37iobW
saadokuSeriyJdQnScGC+0+CGFsAu6+9nHAFgkYeTx5gM/DOGWJSEzSZt/0Icpdt
NjmFJyOOjJCJ3exCJVY0d3WwCQZ3zelkl15tp1J+7o9cf0GScX5c51jX6Mr8BT48
c15IwshNyJhyB/MIkt0MNsXv8Gywnfs/tHA2tDcDcbVPRO/1mjzzZ+kzZ9Ae9K3I
U4RBd8kCHBFp5wa/6yDoAlZspdDhWV9dZNzszwECia2RZTlFPJeh3lRMun06NRUc
7QFEyVJm9mqXxkfWcz/i3dDaZLJTxugfjlGTAKskagaJR1t3sROVciOJLeeAJ6uK
CX3Tt4FUvld5AXnYbqanUnSG+yv+wcPzlOHxMkjyHGtHF+clFk1NQYJeP0ztUxg1
e14mV0OKqTIBELtiGMd2qnijh2pwqXQSXDydd5d8qjPzxp4kSlRoSiKCG8xJXTae
GYn7bGMJnavHiR71XHnT7g2+Uyr0d8HbEKW0cVxeY3EZ2IyLY7UutTQAe7GXng2w
JsTz7HjYGcMqjVVV3H2o+MSFzYaRWRtmRLtmhFN7vqrOFXW2a7r1g9jM/B56xUIX
SOhwnAjpe/O2qMJyvS/iUQFycQfsfpJyCOIwh3yN/Wn2mmLN+L37oho+7q3+y5al
4YBVOvrMnIOIkgK0MPFq57K135M5ZfIshV5mCccEJdun6t2TtyyUgvYqqBaLsxj6
V84SvRBEhxBXHzMVWZ+i7VyXHgZjm0jUO7kp+hPoxq3AfRxbGgTDjqH30qlngQz6
ZDwT8oozVnk7aF+yjJNCq+HXQUiYl/ONrEdF59ZoR3UHpJ8FFKdlZtLzI7OhUOQ5
zoN+s+KiU1vjECYo6lrhYE0JXCsMk3v25PrXzR6M7/8g5PlrxZ0rKocpAY1bCcWQ
4J6EruFh/d4SrMyjEZKPF0FDySSVHJbvZAvMjNvRnWwwhrJweXcsRIKC0xVFcD8Y
YAmS3W/1aM/llKJdvuST9F42T/kYKk+0MNMOKKd73i+gfMw++8zxWij9UQR+G5Sb
Lb7E/Yq+PTOf4XQ5pRFMdMs27UE2d4ugftYVfRqSJe7VZf6bzaU74vnuUB7xIXOr
TEIt6lDtnbjv9QOL/T/0QUdeancd1N8zN1FOdFu+tznGn9JEmaJASDaQtc+ECVCl
26lWCAGtcqAOvD+lPN92JJuQjgVvF5nF3i11SJsCtYvI4NDkzK120qlsFW7Ypqfq
IYQOEd1N3672ZGEdFwAhaU16vugzv8yv2EGv+KjTCfIuOhJIjPguo/bhlJr+98XB
LnjACTmsl7s0MEZsOwmM+P+5nLS8vOxzEIzaNF22IMwMg7qsffNfFTPYekSdpcZF
dInCP2F5Jtd18CMYYcze/678fvp1b5VZUkZnPMdIEp/V4TE2ECCQzFb42DhCkBS4
/dUOOF+i71+C7xWjaJ2Ztbr09gtTHadJQKNSm0fKN0gHCGBrq3bU9RUxXp+HAH5f
m5sHlF80+n72DG5V65uaDebsgXH28B/3LB0dOZER0FDoaDw+9L48/8pR0PAp15vb
8mWfIlspVveuXvLAdKELiewypA5CWbVUx+15wGfX9ejOPT1T2QSDeDIFHoxJUXGw
z4k5pTsvmX9rquBpxXbCV41wMmjSU9FpVy8l/v1c7ldFfk1wpG33E+5K/scF/TMl
r9osphSl9Fa2oleUko0quzeGz3ra1UNEdYRxoVuXzs1x9IzP1Y8lM2+LzBqW7FFl
2xf97OtBXu5th4cQd/CrVX07k4ZuVNz+URPsOfAldFcMhWwHKMA+pUJh5jCxvRrh
+58EwVwRHJYGBw/UxtmYh7nK6PSvle7cmmbG0U0xNgbyrAi1fjnV3Q0XdeZ4+jUP
VcHIeLRXapzK8RMMtEfYGDdCx6mXbzToY0zvTOGEPGgMIfCoYiuf4XkYsBgQtDla
E1KjbdAzepmMLoWnXy5zYHd9Oo59pP1dWEPTOkfC9yZALJrJ3F3jDZlvaliizWLE
0ABuBkLuScbgEn2c9zEubiIu2ClU58wTohVIg42TFjgityfBPSrFoCO2muwGnV0T
Ys92DuZKjm2CGT5voESKjWIpE+d9pfSqXNAxsMgb5OgBSBd3AZ+Iysvt/462wca4
eV/4DSkBlnXvEF3hHVWB1O8xbl3z3ivYPBPRzuwLHAD07D7Fwuujy7lX/nPtQgmt
wySsB+6mV1PzzTimEI2ieHmFwOGJqOYGbE5DqCtGgzhGf2XeZdA1gALfZrnUwEvW
nvePlAHVkbAPFdcy+gcGOAn5O9qUZfvuHS5cgNQUrbu/63H4L1r66ymx19TR45JE
P74Qeif8rqQJGTFUIRmuAvIKWoroBiHQrcPcZhuWvYOkvFDSTjy/QfokSXoIwVsv
6qHBaGIa5eF7QmfRmmYczFEli1KOIHbvAsnXVt+TIH9FXZM/4znCQmNmqNrgiPvM
/gcI9GDdGlQfkV3IKdn5UFffAKLxw7uVOBG+synT6WvVYNm4SZBv8lA15/q1UwO3
epKzJSoUO7EYChdIBuv4sNGRr4ofakCmjPZ54oj1TFXTq1zHh/hsSitjkHfmVL8L
yo6Ubb6mO6l6962t2L6UFyG4LB5R3Te25GFvIYAw2LZs6/NWyFDRoBRTaHNdR7V6
pXeLQzVGWcKs7h7wpQcBWBUZKotk0tBRhTvtikR6vYSyzFeip+uEBQL0LnP5wSlH
d+lCXIpoG75h4sc7aEJaxeKD0JxB+Xa5BAohMHo4/Tx5maFrGtKddXvaq2ydrxHi
jZVp96MrOlk3U5xu+u3ZKmTc5sThjtMsJB6tSWOPx7L5GVMQe6VQVmW89Fhqe5J9
pgh0W2LTJWUgAueLFU7Q3SoEuzpdxNSck36Exd4vsXPkSeIUqxdhdIQ3j6cwNxLx
x69lKMzy1WaoC4f9ln8cKW7jdpx51K6aWjKGHpUCeJ3jZ+ChU1iE0yuVr6zVbOsn
pyfWTCHXieO6ssrDtt6vrfunrMybCKaNkNt3ISHBcSnT6LydD5pgl3IclVlx0DfN
i8O+Ba1y0tnrUdjghwfrMWW31LIOu2oRA6t7p932Ax6MaFmzMfP8nHwiooXlf8eN
C8Iq9SR9EIOkmTugCZwnn4qneHVskG0mzWJklofDUYKvo1IcQtsXf8CTLjCxsh67
c+M3ni+/9EVhhUgs+ikR1a1SoLIJNu5REXI93LDkCTMZa7bHX2S+K5MUD536sVdr
VCasJP2k2yoF3zjOkHPh8bI8BU8XDOou0Bn5L4DMUCATixb9yec91WxCujpPkn8e
9Yo0aQ36b7Yo9LiWQE7xc0Y8b/7eh0pU2l8QYfvsQ1WineB9BYprzRNu1sTEV8JK
ihplF8F5LIssCh4m0JZPkyu21o3BbTeM/L9oQrYy63zB/Wp1KHcZJhYOcUfbsig1
lRLZWGlqJFlnLw1KT/Az/kCD71FdGCNjM2q7A1D2r4AWU7bZCv8NTAhDz4HZnnIG
oYE1EIeNl9gx/RyAhqiysk+G9Cn01b678k6gYQVQq2SEN3EwLKMLmzNkQfu5iwIH
tjHG3Ow/JKMfZZ3Zb//ZuvSSE/JTqFTk9bYrbe4eQiDFmcii1JGroAhoSc/AK4fz
F3XOpPCJy5Q2W9Pb1/Wj4JcbyK4IL83ZSGjctfpTqQ4idM9tp2fDDWlAsqEcCCDP
u95/xRqV6gkjYl5OusV/Z7DqDv9hPjYJFFCR19+EViSv9SxrHv6QeiXEfhGn/+Dg
Gfl1KfyVvXfYu/AFojPXHRG7qxzERNb8jaMPuam2PJtUjsPAZhzMsNwAM+BhrBrN
PEcvuMOFbFE/Qzsi0FfSUsesppHiK9rA9nnYJJCR+cPFUB9b563Cx1HA2yv7tsVD
gu3vJqE099suPdcbOgBHQnWFKXe+g8/SJ9BuVGLnZa19HyGyi9u7PXP5hrA+uusm
Aopz/OV6d3s/7kbH077WHn8PciOJYnZ8sS48oxYfxh7vgPDFkIK1XC+wOEgGMrjN
5dhDOwLMy1HoMR9iSLdOjk6fIb5J0MIq7gs3THujh8h0PVLZYNASzCNf4ZR0Llec
raDCsMOE5ICUjFDqwymoHPegba5kaKALWoLHl1HoAbrf3oOxveiG3yY0czEUBn3e
XyOGa9Gott6ju7T32GRS7g4PYmec/Y+xplUK/vvqxuF2KMAccaI6QH+j0B9/NVWL
WcN67fnG4Bev5MtYt8FBES51dmIT3lVKTtTrf8yf63VLfZ08JR5caKPDFXLiqFws
gKyhTjNFJtFTptjrEkItSXTl1CWUdcHovPRUYTy4CE894VABUDbmebFv2Dvqa8pz
18K75LLTsVsyroE9VgpCjZVJGcMVeyX1CsFznOTh5pObVeoTy68CipN8s/y/dxMZ
mpNbnKvwGtdASy2IJu9UwG92g/zZhXZyXmXOAMHGm6CHNKk9UHYuo5ArkUKLJssX
TOl8E0GqVEEPfJixUeFQC8gquFLCppPvoDvMlee7MPBBoEUpmYiYIFXneclk4vt+
2WhU/FcZl6y0h1a3bha5YQlU736tpBsEfnAQoz55eZgP8jxbKGjj/KtqM/yYWDEq
qqJ5rKqQy5clG8xNXEW1nt5FD5ZziKBmd4cgMOjjGpoW4ikndYvNdAAhM8kU7Yx4
Sn1LVWi3uzI/AzaNfanFBVEB29WG66QEI0T33tghqPfS0deGXW/I1JHKXpZ8b61+
OyyJIlwa0hdhadwPDrGobyohx9EgzoOTxZmuPbXbIBCWCdj3zSVqAu9RVi9qXIXi
h1h5ohK9vzK4QgW1bbID3uOBMLgIeH1pshIUU7KXmkdv04ZKOy+t6gj0IbgOxr5f
ByCJFKDCRlCX6OBu53E69MmRnpfOT7T7gePxToEQjKZXkcuHVtiFOa85mvpc5iRQ
dnLN1w7FDr6cIod6SQ00ijKrzHezCAuTeUY1cllUrjXIeADufL3fHwa0L9ij5bw7
FWel4RhpGR1e66owsCXIlLse93O70RoSE1m2IYPaDKyZ9+eKcoBPSr0mPqoRx9eP
qfW0xBx8+UneT/fvOOhLxLJE/zAJ4FTT6qPcWpmI0LqCuy7OkElV2lE4BqeVKNMK
IUAh2tSpzQxqhDhZPO7yPUBiF6aOa6A2nGzeQ7jIrBY18NaATlWu9Sb/zBJK+Q4T
2uyAt+muG1nlu/3hO1K118faON1y9fL+F7k/XvmvMe+IxBSWuUrAEE40qSWCZMER
vn0FCR61mlI66AK8bVDiP84RA7/dkKdLkzrXngKmQN42ErMblztZeugArSNjLWZ1
ow/SJoDPad3I52z8l28QU9zsxrvLiWCg3bK82mhvvAguSpL0G3KvALI53ddluilt
rSFiSgV7gL+NhU/tc1CU4uP9ucR4vabFKFHaxyymIkAK7jyFrZAWe4A4/NJEL/9Q
EgmKdcRG5lim2wUg3itcshC1q8SWztpz08bk1EY0SYxJdxaQwYartP3oDRW9Ii/H
t6l+AU+StR3yG7fK3cPljfzl3MMwMCc4Llu/o0NB0kOayLPB+mtlvj+bTJZScH47
fGytrA0kI8Fnh1L0dJPzjAeLTjN01KP4Y/D1cntnOatdWWV033KxLV1FbbUkfnfI
SkvNX8peBuoG2nLRVlZBzC6ZilDU7+MiQB+nQ1TrLQpSa8f9MjJz1CZXyJcgSm8Y
2htTwP5QbnwTGH3QE9ST4I2flL8/3UhnHDt1bbVQimF679BT8Kb9b0RsCrCihm9t
z/gEd14I1mmwfg13UGeuzBG68rwqVdCmdg6lZnlopksKkp+Pl9IpCp8VhiEx77uo
4LPN40gDICy6k3LE499L0WtnXsVbPAH8bC/wCni9eFL29HK+Haw/8h02ovjNwO1Q
0YeLh53Rtw5mVSNZxoUbqJNMVeGE1h4GDCSjNE8bimTgCBMRHrVjZbdTQI8u+iZ9
BJZq6F+fZlNaRxvGIaaFX6tKxsojnLhr9nTuLLY58XxWAcW5Bt7CAyime/KMbXxz
o3B+2WUGy7rDMuOrDuITeh/jd/iU0nST54kT05XJfsqcHi6acYdtS1PZpG7/XUy6
4M2rVhRinQ6xMaBnsGh1dHELt/n5uaPH9v/3FRBennvfxK7E70l5M1N1BJ6Zu+1O
oSFqRZEH1FvwRt7QvqSnzaNmCwgmJ6l//P+a4AUwkFvikhGnF2x5jkl8i+gqFjtX
Qkc53REapCaMC9bOsyoUT6cUY9eFL2sAJcgaZ5A23tyzu8lkIhkQNPrOjDKJHpbr
iMSzPY5yCLd//eaTI3xyozYk3AqLAwC/XyUK5Ftf6vN00N5bMsVmCtm7nZkUbVAb
z7Kz5+FPsMuP2hDmvYBZg3PJOgphAne3Jlcbb9J5/6HKcHIlUiRWGzuwjD45hJ5d
hCV9CdT6Ry8douSG5XIjzg2sjUeCqzBfocuYNv788Q3nLhJgAoqMSVHW0dcelknt
kJHFT0AY42NTpum+t31KXFJ2EOOhwCDysraEfbP7ZednPVy260BcO+w52qzWnEMK
QhIfgUlsRBgzyFUBJFSg895nQm1IiRCdVdfMB6xvQKaOAPvWqEk7CBn6i8ONbeZY
sp/BvANcJWWgBnezg6IR3jxja8Ud8l/KV0jwjCy7Vs8RvyDuutvSB5k+VXoKasIi
xeikRbAMC1Fkg9BlwrKKQyMhqQAJ9b97Sqt9HacHHz8bc/oEt40Wo8ULltZjkTQC
QlOryyOdp5/K3oAmjD0o66RftutzGpbMKOMQvOGJqvtiZS/2AXI3qayKiQJpQQiU
/gR0C51wsD44md9EG3s0LKdkAXT75A69IYGqr5+QRgk1DgmqhdxOnwnw4aBDiePs
t5MX6GjFMvytpEnMm8pJoB4TigkOSdOXCuVu2ARhMTZcAk+Wp5VjZaE6pjudGxPQ
H1I2wypRtxJLtBG62pb5aH7wll8j03O5Nc+asRwfGbmxmNH1ELy5lfCW7QtXuEEW
diDB7kDiprho4l/tPyt08ugxW4jRcOgGB6EZpo8h4lBsWPLRulWGJwJXyGk2xre5
B671jqwDIeCTrUVUKCzNDOTLjQeIMhbQ13/azF72lBLSp5lVxkhh+5Y2phBhL3SC
nfT6CrJm9HPkV9HBhLsdst5ocIaN/rQfQzH3+ctgnbhBhaXdaxjx6WLgp0bxV8/G
MOqeMbIk6ZowF8Vjl3bewxhLiMXwiLb9Qi5RlSK1hCyzo8Q0ke8a2yjEb9YmF8tc
hlPcsQtSKRDAnZglcqoGrqFFftiKGbOmq5fAMpvlrO34o8jEmORNfUhu+cRO5qf7
2aN+ucH9P1KbY25jP1S/dLNgCcRgVTZEfLMbXSvyvxFaWNuUiPRSFBT5iP/rZi9D
0lwC1Aux3ZtUCahS1EX7lNlwz4h7eepzE+VWSxxupkWeDUvc25/zHqmlHY8J1sfg
y0MQiNgKaJj0IU1SAknir9SxmjM0u07B9jdoiqBYGPONWp2fJgFtXRoWymh8eRMX
dV+C/6RJL46u4y0Ncbn/jMTKQgXaG5dmRXoo5oculIArYcn5GLaSMZ76kRZoOuyZ
YZZ/85jctlfcuyTm7//H/KVCFTpXsDpKDE8nUCbIUaeaDDNeN1nSK5RIsBz3JUlg
FlGIUTOGn6MjiXsq4UOlAD3AHSlBJ0W9CUiaEociu1yH/EiMii1nVNgJV55lY6LK
3CH+EJL8wylunJkKH1YovMHBxp1lxQjbMZ8aMyg3fLJdCQ/ZMjeJkNI/5R8ygs+p
r9lW6G0e8BzVViy3RcZeh0S1clraP7lat06+Akt9wvq6rdDl0OjaTu+aKKKv8Wzb
/iD9aDPmNLDo5uMasDj2qgVisQReMDBPZsW6DbwDRfcH6OXIR4MlMNQHSbFOXMMy
al9vIyRInCzeBHoom4/EJRiPl7lbs3SvfLsjfuT0pWd/fY1PDVkVRnqTFxyiRZVZ
YhBp6BQU1t+MAH+Eu5POqSDmKSlT2OBYirUgLC4B5UvpGWzRtxdtAUeKRYX8RZJk
QbrjrS2tTSko7iD2VESzwVTeJ/DqrT0D4eR74e/xGPF33L0Wfk1f4Xu7CrE2+Ow2
P5OZTVPs8mbpb8MbjVX4TXeUF6QtaZM3Gw4UdfwcFhcWgpOiYhpxzz0r9USYa56j
E6ydSvlpnGpT2BQ3z8/BJVAULydMwFqrThXsN16UUHWZouA1a7JUSduJCOOOOLKd
5J/zm8726HtmugPzSJJC3QemPtDJfBy8aHAfJCJBuI9TvW9ZiaLjI09OlCcK2HZF
ir1Sn8b3Ce5pOP+FWrEmEdjN+mgOfPCGEhL81WgI2f7nusLlHg4TDij7WIDl6T6V
yJCayCm3nkgj3J8Xq68Z4QGpkp6OkOfpkrV5pv+Pt4c8R1QRlWiDzQY5csUMqy0n
T0DVX7Um/IU5DxwCauOl17ORywAUmzDgMyKDmRyRVIjU3F16lQ9ZhmFtDBA83ULb
6y0kGRihvs0Pmpxw5gSxwmrqwsXCut2vaol11Mkz0fnHNScX7qgBNhlE6+zJeozK
alFFOgAGymv/T8QJJyX6tnbVm7Sv2t+tHSpiWKuurmH1pnP7lhbk83Iie4LY7uoi
FnxaOyO81sOYwRJs1CQxX1be/CpVrvz1WhdciLx8i76IljmGK8zyiKfk/f7Zs+4b
zeQf3sD4OK9lV2h1n1/JHOI4cFxsNuXOFhVUEEWSZCpX1jzzPhAWCzUmQfd2EsTv
iDPyN1MjjwKiSaO2LDZu4OVQpEYsOjBT/QCVpFZY4CpotRWKmBna3P8YRGcRzVaZ
5+uDAMB5eH77N/RbtPrlwNyO2GdBUn7E5Ycoq8vgZhT3q35SC9VDvcniGVSSVvma
ftlU5vwQieyzbMyJiH0lUiASlY1EbNc3nAgQLFY/n1fyUvzYNjZpKGxqoznZ+/ib
ZYvoHAiheJE8cDVChYAJ3pftqJXRnZe0v63fgkyt6kRIFpBCfOxiY9IAmsSuxlX4
g1rH/A1HGCrRlsk7n5NVKEHNtM5Ouqy6yVxhLmGLpgFqCnCvM4GUj1gE2fZEX06Z
DPJE2DqrH11dOM9W8kMJ5PgqPChmvovwsZ8B3z6CRQ5s2qkhOv3ZCGqrpAXh9dSf
YTI8Ws7O++hektkKJFPJdxHAicnsDUt1cxPPJ/fzoKTy1VHeSoeaJ0cnD9o+vnc4
zw95velj4YZ/U3ZwpMGAdqMOLCy7vdtd7/GrcjZ0bpo2g88hy+OseIMKr6jJteiA
Uj03J68uzLfn4WvJTWAQs/830ZGhlVx7wko0uGEy3ExUEmLMy83bnQhju/2790oV
hSwbzj+8k2aY+FeSWvOkUUWcnNlsy79flLBJGPvpi9uRPBqKhamDLVBfOFpeSo0s
7Ssem6iUmNVxHGnLN1XZ9f7FxWNd3y1VFEzFawVuC1ErIccAzF2ouEuGhlkjvCwv
+jXIfdQiWJ0bH1k9fI4zvdMFeV91yuAP1jkbIhD/uX+vH043wmiK9hX6EEGBZzJr
aKxYW2lO9BSbx48BVfJsaWoBNGVKJFIXqQEpN0O0kZsmhO9R50yn8tNAV9kVsHJs
UOW5QXAPxWL7O9FGMv58BRoxl3SyeHdKTU20o73YFAruI0OkAe3j61nUfk1aaZ4E
I2YpXLl+jM/r1bbhaRP7w53545i5Tqh9xyXv2ujLeHBzhcO9J4y4CBJgIEWKerGN
nugIc2nZM+T69czk3lP07+vjedAjTCGMZDIh2uSY3nleXyEfzmvKOQqv9wi65DlA
GJHq4zCaq8HMIDhN4b04X9t+al1NutjKCSFVAihrmDJ+wCKIwv1IcMW6mK2ObF/R
fNpbQ/KXW/6qDuccX8xFdBVfH5rsChtat498Hw7CY0aubOISo9DmeJaKsrM7QEPU
jEKb0T0RjeSEJoe3Q1b4MDgF/wAQtRxkXEYy3AaTaqRg2EA9HNdlf7nWkTiLDFSW
NMuN7bqt7Dd9njRXpX5/VA6mv83CCBH/j/v6lK7rXtZJ+y/ao0DtECVq1atqVrP6
5ESJQ0DwYl2uldEXWBLMl40UcP/21bnLE4088vik2D2uZZDas0nxrfmoHeXlyiSu
UdQ99tPgiACAZv42/+9+Msd2sqll3l0IP1vzgMrTcLohnL2VkjvEsDUmwRcV4Yqy
s685qUykXAAMtrMmx5E3UMp7ucbmM9SupDPo6zt0oSMRuspU83zANFFULARes5n9
NzAZUiqfgwMQptTZYUNyuIPMs3XfNkf6RL1WqXtInYjuxCtstDL8qRg838we8+p7
MPPR5AbGA/HS8715Na8I+Y5KzaEdpjvTJPg5ADlfEoPoFlpGrVzN/PTxaKcctvsW
LrrPQcmH15N7fz65E6K95ybi4hTVdhXj+AUgBk0LVGX9ExgdoEASHxLMeipqv/sd
xz5stwiEzC1Omh6RPsc018iNTluYsapevBqCDZwSLtzNhacfT1SQ4UitqTMsFZaf
1zFHZAZ+fByhQodtDE/AbcV6a3BE/kAWFDN6ITgXAahfrm4nYCXyHuOPqzL4B19L
TC1AHcN8eiZwJTWCQVYyouOAYKpRCjcb/oZuXnVPSm9ozNjMo/pJPow495DErCHU
nyjvjs35FHpOsT1BNUkh/GvMqU61sMAFckUjEBsj6eo+LKrYA+4akj0zSzmPlUAK
hhTiYb+VpC/pNK39cwrRu97YIWFVl8e8i51sgYTJQLHD/L5kPL2M3vjXNp4KE6YL
FWEd0LCIAP91dWQcmy9Ftwi6Ko6CYQp+ZcbDoLzbw+L1ibELra5LeMXT01WaJ+YS
zVVBrvFccplgQMrFRvr0yuPF88hw8KmIMPeRPUJXOWqzm3suZoHrZfcNIAG7hBGc
1lXnKmJzK8qnn5Ah3juGoa1Q5vzzK0qNVOEv9tdOKr9WZIAojV04K08QjJVZvhaA
ZyN7D0q3jsbz3BmoNcIoFng7RyH4+o7OjdZc3jYK3fYRq7NAAH4AYh94y6XR+pq/
JhBpEpn1HlckT6zXfN+66KwfBdl/tCcKIRH+g4NqT1KOkpq0i7WeWxbh+cova83G
8qdkywH2FGwaCkFesENJSAvbIg8+w4BQ+/qUTl8mF1bVAcNXP+CQB1epOur4T1XQ
3NSLupticibawrIdob0Tn+ijheedk+utfyB/jBsPqBJR2euL/ejJdufhx98aNBNU
9MsStxz7QDw5bWiztCiJ5D6Fx5RaA4Mq4cW9rCvGukSqgM6BTgzLiuf9ylaQj2qo
zKktt7vLsqWR4LNeqNHk8m9FzVsFEZZdC91PdFAAI8HfCmzomo4ddsDeEiV8FpRy
ZfuTtq7W8J5a3zz50ccwCWO7ygsH453w4DDe8bhO/D3sCYR4vHau2CeE51ElEEFc
FhSyWnWjLp4AHwkilDHa1uBn1gnJC6MhoWaaOMyiYHNJ8Vv17fgPBcejPM5dBQNH
cMSyIZE4a+TdDvLGgHKJE+ZXO3/kOBZ4I0LcsxtVraWxSuiJEBZkzHYecrF0/teF
DDESK2Z7eQ7dmin/YwhE+hiSXXQvFiUTuBzxty5iWHMYCG8JUmoWXypW12m4bU6O
TGiHnR7drV8uAl8fExfBAoDzG9UFvGzpLk0xfRZaFBFSgliPlpZwhhWhedbo7BO/
W/joBslBAcjoxm9aHKANycVDzo9fdviwvjNkDFjuVR/AbkXI+pEJ6ngjxcgvUZS/
/wDUSGRMgXqGpX/xpRWMaUHlHweJVJbDH32rK2Xj0jV/4+/5DR5V8N4XwDmsC3we
4XuMiGxMejOvNmEuWLvFhmfCsIPVq03bk0w+SA7MmjzELX+G6Pqs16OJtuC5Uqar
upKkHASfGH1TZATpunf/ty9o3iflXdMUKhaUh1Y8YtxtGD2aGN6yivpk2EatEi+s
db+et5tHHUCQK3bQUPrNFL+iBxSFT9PovTf16lvtwhNCgTbofg84n984e+0rXNq6
kvZ2CRyXcO9lQsKQphv9FZFQRyl2+VTLLbB/7/kqKS04HfS6Df1EvhOBIChaY0zG
oWGQGIuYuKNqskzRPAkpbrF3OoXpqsTuy3XbGl+Qv9ebjaE6Lm5CZ7bwI0H21al4
BbgKpF/ZvjGgoExrTfx1925VBrHZc347Llhaoqpx7wIV0roJehsPsLsLJY+paYOj
Z6N3+qQeZsEjr7RsrNpZ/+lOYuI1Vo1uF398N2pi3FTXjpVxqj4QPeiD1rW0+QQd
a3toIK5PvjU0khM4SIYutrpjwqEC0nB3lhhfUahrUPFVcO3sSAvAZZ04t+U9WkQD
zVrUfZGKh5LLPfX2Y3x9wEi28XsHoOloLzfagJINlmd5JE6Wdcs4NDutLbo7eyCx
+5K3+Scaenp09HCuHAYCrSC+OkIIIDnlRSgml+wtx4GCAkmA8+Ik3OjSOGt5pWWa
7Z7vAJQM8svQ2q1weBJakc823XYWFObaDBUNXs2gQnDOXfgHPr8NStEwY0JxvtQy
vtfFE2qVnQfEan0677FLC/JuWnPbSOTumowqo4bvcPMN5WcWxqUPuxl0w8M5srTo
VV3RPcrcnrm9matpeVSPMghd4+8P/lrEP1TI8Cnc8tJXuz0Vx+X6MxUN7EyXkksO
TKClffRSd+p3vUk0B6lPpRxY/J17xt/h03zNHqpSVS0Hf8QW+S4Ho/7cM7EK4i4D
vcwdqrDGgqG4rm6grQauvYMrnNR7dH4sY4VhlKSpwKp4Lv3xXRFeaakR8OQp0em/
YxXqjume3R67ncFuuHFE0QXWp6np1Kbh7DPW74Leli26In6GPp2dIs0omjoIeaJW
//o6SGWOXjM2S8UXtzQJoUw1uCNGX5X9dxm8rMe4zRuKWPZ3Kt+52egp8Fyt6dje
MXxRZYQXWQJgOosWDOo4M2g0T26GZpdwSBPm0XWapueELHh6VZcV1BXr8CROjo+I
VQmujTqF1HquY1uY2IPvDAa45Chc7tQyx+C0F/EoOM9LGM8YDj6Fb8TecrVr6fnA
vmZOdmr+oIi7eMZKGL6zy8C+Ou2v721aT85Z+ubc9dkkZWpt0Lwuq7iRc9qyW4ni
OhPbY5Bo/3HpA6kcCFpH/8zCbJvZZrAELOsiMdpMe61DxUnr2OKXG/Wxs4ubixdz
w+FQqM2fCu/p8QMpfQkDLwi9Ai/ph5fFfA4EZYLlfzh3kivbPOLjECFkQ2FQDibl
LYxdQXqUl+ciWwAXj8kAiMabxGnQBTjT9eSSukrKQdz/B56TeA/8QF/W+5mb48NE
kTVZzIsIgKVwuLzV0jfWEka8UCdmLSQLXc/fJVEjntllb2+TyMzDXdj2JYZQbqjn
TXEpIq0hgJAiG+pQDxwFTl1Ddikv33Ef4aSAkLmNu2YYF5Pnp4AAXFcF9kl+oHwm
T0fLucSSyDbKixBpue6DvTTN2hw6It6gRVnQTh2kz9cZ1xpCxkA4E4G2uSUNcUuf
GepBF7EB99w2S6eNRY7BUyv4M7++eGF9Ru1dEBmjtJ/Al6D/mklFEUgBaOSVhqYD
VNpPfuTAA0ucvk+DOkZaPJBE2pC6iUJ5VRjgy1hRqdWOMKEmBCMTSDBbIIZK9o36
SjgpAqCgMwzYcaNgM+sqsoYoYIIlABXDxjHwiHeaCAW3mehZGubxt3NXakBQ0cHJ
wJQ8Ur9sjDi9nvItkNV8bb/DnKPTgAz5EmFMNVd3GXzSJEFrL0t6MaEG1YdDVyk2
WkCSUWx2dIVlgBXIOHcFtE3bsHfVLohaP1oUDwBMbDlVXWPcXgNneRDpJXjK1bS9
g8s33IUna0FQMbVxsxSW3Ey0zbGBzLrK+WrzG/Hqwq7uvUcJJyXrcTY7+lms3QPk
RtrXaMUiLZSC8XJrOlnDDZWiWGfbOlEJMy2XDjL4pd5GYg1p/VFvSiO5o+JjQprC
jduPr/IVEvh+JLHKYQ/gcyTt+60GftzUVxZPcYi0fH7yVuSfj6Qwez/UlpjPIX/4
cBXytT/8Yh/2MyuKvDfSzIconMoKINv3PYKJYIfclRtpSa7viHZpr2AtFKy/eXmg
utkUCB6qAogRsbvwqPrU2dWPMqi6zXuAGg/Drr3CKKNfL8AijBxCHZ1jf4L4cRt6
dJOJew0A1emrZ/KnlD4MbpdyvNBI/LpxpQ6CDqby4fnD8HHUEBA7xag1fXTY2vRR
O3bB4WfdyXAp5MSeAymlQq1HibPSL36EyHwR+VLhqnwRAALX8YEGayOqkRYmVoh4
ag13uMve1JMUCTbZle8VfgHfqvxKandC3DIDeARvtoFEd82KEdLDqatRd+ZKmTHX
whmp6t98HZLKkYbPQBpn33Kw1fCVEooghpuPAel7o64TCl/AlTzfAUZpqqBoKJuG
AU7R93qdTfvy1kS9N6uBSBK6B6Bt6L5PlLRAUoOlXBNjjdCpDXvG59IqCUuQqY/3
ZhC2U+8a9mS2gqSutL8Ljz7rOSrt3Vm8hENb2qla1ndUmn/s3D6pLz86Xsau5nIE
Dpa9NEOttrNfGV8cugsAqXdZ59puXcDUWg4Os2t/JaUDzBvO1fAGHCcdu3oTSPbP
z6gmlHa2kJR7ZsGfFNn7YA+BaLVH3tnRo7PJ1wGIQzNWBi6F0v5jj8Tl+Dc++siz
3VZzeM3du0qQLIZSMdwRZkluIMlrHSukUcqEjZKyQFox1ExHQH9SBjxq8I3i27g2
yjzZALvA/Ilw1iTfdyodOVOkh0jH8Sm/zTG1eWtTEkzO+MPy+VCmMrP+/RpgDfkt
AVpTe75Ar+xIkEPOTRpX+gDHxnLkxr1a3r35JTiIJIYd+8jAnzeYBDvZZKiVLYwN
s0e7ZYVo+BQFKhncpU3h60twXaha+dTdV4zhU375LEJxIHNAvirUrQVTh05R+sWr
q1pvWzJ4rp+VHwAEKcKKlaGe+ofx5vlXyHrPz+lN2d77bKfDMR3Z5+MbZfi7Omch
gsGXmI5+3JXP8s4JrreKBmWwROmNXqoXoR16QapsOuALFHv4uHCrFpBXe0bOcTg6
IWtuOs7fLD56MEDh42UsroLZvkvLe5mYsTlff+e15+gg0h+hRBC9sc9BbEzB1qvG
KbqXDJDY/jZgvr8fqm5oYC/Fpktux0jWJkahgh8mIgzbsZvQYESnbm0LWoHCaylp
DWWHVUiXy2sS89PjHJUMPL3Tx3gYsagOh/n+cjFqKlTNRznWhPiDpzT5JmJCY9hf
ONWtSOxUge83uMSSOFPOWFJlFYgYtOK3jqlZxDayKfhGr5DFnV5HhFYYO0k34C+1
AfbKIB7hiZstXFYyNmtk+s6yV+xmWljbO218DTpjbLJ3IBG2K5weuifEv2Zn3HFv
0x3/T8MjwiZ7U/qLHm+odTPsU3xVmaoIgFpuNbyzm7iTIkW3B43zDnFKgjAjjQEz
IKHDW1778m/37C1mN03Rn8sYAOu3MX5cXdkzSgCJa84jB6tkc3BnTxxkFdvjmrQU
5bLqUO5xZnXQ4lBfjbk35gfRz+nDdOFWazoI6la17XytUTDtuzOg/oNHqD/qQnut
4aetuaMkKs9bQVYfwPC627Z0Yy+8i308uSmj7IsHkaVtartvtUL9/d572vZnPUPv
MO8nm5EbqUfUv6j9Mm0Dbqo7MqQzN/VNk9OKBE27kHStVasTFwXRJxG6R0WBcmun
jSvDcJaSit6QbRJQ6aiFYSnut4OCmzzyvm3/8xzMBNzm9ekS9apj9oDKvSVAEnZb
6+cX+BNkF/i7WLW2j57PlcDdZjkdcilax25ugdeMegHgwowg8Rq3jTEwPB+BjioY
6ddeluOxrgNg+CD9Hq9kFK9wWHlVcB4DIwh2eByVlKqntQeTXDAjMFHoLPXr+nGM
DMMgh+pxLsa0NGVnwz3fhbYet+x0S2Rz6MZg6PbFuJFtff755WU58ei0jakY/s0d
cjalSbr79TMVwuZMzLBZRSTXXEKByoE9VHPYbwcWbIc0Ib+9Z/mQRJOXFNh2PD4x
tVv20YTGZU3CMLUpNlIw6Q8NDzJBLdffXN18odTZWv4VxlaP/zEr4Pr0BYdry8mB
NhSF0b2KJXU4lTcZUzjmchJyX4P2P+tLuE4SvzeJOikXFWcPIvI4OzDx+2LZKOmI
9dPH///FaBb197m7ytXzy31Wg7v4psvYpxvtRDrXU2RmoHQ6jdo0J45ISh0Kxp5f
EPz54oU+vADcdK0LFy7JEJjEzQIcThRZ73GT7Zc4cogLXZb7/hQj/2grMRnhQR3V
QZvRoA+eDIT/8BBB67rCaxPeYrYHxZVaxZRpearxt66ud8L8TSX5PE5vBM9hitX3
clw79V8P6/+icfy23GKKzjFmRE8bZTOKNk+7egmi53CFXR34nwxKNeGUHs4J/dXv
peyuHfqlaZMi14bCXlrKLC/dGK+sRt58LraAq7w0gNk3S2cBnYmoWPjKhsgSahZJ
hb1wcZ1AV8SQbcTJdOd/ZdjPwsImJZXfkLCwF275sIqChX4tZtYePe/L4uRcyn9f
ZR4vQBQ8UFrXfWOfsX1IN4HW7CEe1EkvzANHQMTOSfA8mUbpkvxIaRA74UpBQYBa
tYsW29WeVhwsMRNpeKcNuGVoUqTmmKdIyWf9YPZBfHZhkz+zwDnp6zwMEnF9LZY6
k5ON+W9ZDyHtyAvmuaNHQr5+zAEAOWrxnu90WPrBce8+yIjqnKfhjxi+HgB9sD9q
2HIxtFiwlXKZxt1/IJL9/JE0MGpuCS5/FypAiQOPf40omowPr9LhD1haBzMBtMSt
nHGUbx1fYlJnowQfHYLx9cCh3eRzkiOPTBYtxBKKuq4Z4ulLX3DxWLY6A0gl0p1u
sFiO+ZdeA90SrNwgGNIbcICTW40WD+3TGz5TxvQ/fWeBv6k1KtGuT2SQ7DqL0MJK
Ya0i9CnPlDpdRCPvM/v2+yS30yOwujcysu/7KP9bGKA2VHHisaogGf6PZl5LyySj
TgsJbQ/R5qm3D0nN+qlnKNQRYtkTb3jKAvG0jA+cDKZ8koP0MEI6INfWBABfLmWo
S4vZaY/njYp5Bztxw1IGYixnyTj3CLgFvRr4Vn9mRKmGAKSvPZr6WaQrJKDyMuzB
J3iLXA/lnPF+0xszcjfKrE4Vn6nIK0/9WPxGv/XdCUx9HEdlSwr/FGGzEoyZcrpZ
Xkx7AKlqAsfbbu5ZXPBFsAvWYH5JIAlO7Xh2mMswolFUyrBI2U04zTJi4iL6LiSP
SBljgwNUNriG/S3iWry4P2Cd/68oOzSQ3Z+K15sfAD9nXqJRxF/pzHJpajctCT/S
zMayluH5EbePFJwY2YU87NcyCseGI2fDA/FwBZQ+3oaq+7cJA+JPq+AzOOVNl17N
+zdG/WUoJHbDHQ+SMQcmlNch07WPILhJnnIrjV6Umpor8JB3kF4UvOpJR1V0MHGv
u5szZcNs3Pu+v5RRbis6NmltIlZe83dnNcpiDFPPH7HrV2LskVbej81ScWPvIkO+
frfyFjpJeUSsAMVDOi5lZbUCV1DJ7FexBEpxy01Tg3kdzXpO1QWdTVSnHARbeC9n
J9oCnugcNsJC+K70fMUnet4Bkaae5iIuba70EWJmO5g7/9nPQn8KZ/28lbfrvCfa
3tdfg9teEdcf82uHuIMKSe5ZKy9zxGys1kvWjZAr8gaxLDwZcjsuJvqFlJef4WUU
YjPuW2l9ro7s9ikNCeoSSpqYFH4A4UN11OjOsinByaLw9xj5e0tmYi/Gb0DnqmsY
LrU9jxeTinLYD/4H6Fcii2Ip8XvGEoBWtVfd4F09kzNSNlrAx5hMzYmTLp2KWiHR
DQjFyk4q1FN/gHU7JA64ApKyDuCEcgAdnylm1r96pCxLrCyBbT+lrAjFF+jiAa1m
/sSDNCROF/SmMCWcMqEayeHTD3au9qDUUbje+24Ua5ql1PiBpFjOM5gQ/JeBERjK
dD9IgKt41VpEc5wnoOFPJpiq6o9RQ+dIBrhxnZu48uv2Ur/ioYP25iQH7Hgk9gtB
FPDV1KK58DieHlVSd9nuv5XxfMEyncyy5/Ow2wEnoRPfo9euNh7MI5MO96RnTjd0
g9wEYV+d6wg3g4gybRAFbcx6fSQqejyZLL3A52308U+z0YbmoZ/f8FKrtm1Zb2GZ
yYpprq4Ot5trlwEZmOfQumILFiPtJpEcjvh8a880bBYjnky71T7DvVIj7o10SzkL
s31Er2diixxV1kFN8dnnmpsQZb1E5yRIwGu0TV2RArGCKlh4lHLE5RcUI1uEX4dz
Cc0WzOkVctfIzeuj1fLnzRf5AiwLr9LfHIuWCBIG+r9R/IC5XS0RdOUgF+7MCab9
WatQOQorKVvetA9P4Bvz89XBbGtYHb4aVL/01vaeNBWYp/KEKQ4XB7Eqa/8rbrk5
nWakAsYJDDcZZim7UohpxbSBG7DvAep/A4pE9nOrW/4D3ofCwKqsIb3v6lpamvFS
VuAzUzIgdKJX5829q8R2Nuw4H9JICaT4fqYxh2Ce4hMpPKeD0akRD2ndcQNlHRMM
KDxVcyzqu8P5yGJwOCmzT8lxLZUt/HyqeKK/HysILZAH7VW1iP+zBz2+QD83lSwL
yJx1U8Mu5C8bP/Oq+4+M8TWvvOXH6pOHD5KPvwKRc3fLLsczDyt25cxEbxyucfPI
ULESyIop2gEtPhtAjTV94lRRWpYlxwuSPRaybD/OqSXFBUjMFaIWrgCbUthcMiik
7iedPwrr1Z6rGbHtRCUdmrYDtABgLdA0gkJegsO8VpJZvYfkZHFUA8lJLcXhTLGe
3eIgl5FH/djUfHgF2gEPhBOHniGLoT8aNjtzaR90fd99QTbbtcLVoWY68BJRYKV9
APZRAcAG18mF+k3uGNgpi+LqZbztfnTOhxtLNE90F3fTfwHePWpLT3AtRDtijMZC
44awQLw8XrflY1R0BfIfSQAC6A3rmmjSlvO7MWDL6py9t4VQ3NhTVr80Pc5nXcDd
43NU2DwyIeNzCD/wSRIIuhjYrgExP8P4y3IssiHAbR3JqHFG5a6fl4ddD6z2R25k
LcwzoQiQzIkfTXcFH2O7opaPCV7lg/aewpdWkGY4P34pgLyEqx5/MtwCzJjAYS9Q
XPRCF0pYHvKh76Pnsk4hv2Div5adt6xR0bURtuH8qiQy9H2gsJLdzlTEa0aRmrl0
2ipFtZBVMIGWWLfxQ6B9s8wQnUatkfKWzhXzT1EX4qXyX2xGFPRl3rIXonsStitn
qAa53J20CEdrgpVATW+6QU7YdNVz8MGNg3fKhic8vEasDZx7k9cdUgmCsJBWUdz/
mujKQQpjbEkmNcas5Nvp4JpgNIhhYsVlIhWMowTHitP9O24Pz3BXeQvzAkBsZY1q
eOnnH3EukM1ZeR9b+rbFaZsCZtMtpQ/ludb36sZxehVf6LmuWVLcZJzKNtIco11J
w2iBo0qma2cyJRo/ET0H1nOl9YAcqeort6z9YR2NTvSK9zc2wSZ31gJjy36AKmhp
ZV3abrjWkuC4OE0PlY/GGO8wN90WyjkwK+4Qw0CDR8x7OBNmMitf2ykyUj+yUTm6
w6l+elsgKMoQCqm74Cny514uyaIW8XBKf8ZfcijLllZFjRKw9FVOuEbInwh4AEHS
khRs9JSKRJJvdfvSFsuI937XR8e1h+VHoJ3qZq0ECkVvK9fAQ5CWyfhFpq9XqCYs
92ot5JNOTrnbw3erLzgQW+z6HP9mKTxxnGtoAAN1HXPmBucYQjCwCXaTELlq7eZM
k+EInQZOPS9V5AE/3AMCbEMe00pXRhap37M4lkB+CdaRkZcXb0glfnF9PdUMGKTl
y3oGo/ZpBIIa3Y5cqdq6tIQ+4mTKkBvc1jzedJ762gVTWa5naAF1YsV6a0r3MyeJ
aPAPkZCV3I1aNOX/DLt6Zbr0NoJNH46GQtRVTiYOG4OwRlAOgKdrzoUEfrIIjqZT
d143YOPA5ZgNJo55Egfp5cMBaVuSgK0ZvfgTk/nEBz41gXHhtNEzXUWXtx0UkRM7
gmkQoGERlsQhd/8efL6ayKxNozZSTeLKTvyTY+b+ucR6zG8h7fnMzhIYhKshNtcu
dwhBFfZhKOyq/6y1UhfQAdDu8tpr7QLgX6dimRVCxjMeZBtWBs4MjGt2kLTB2M3I
K5+YKhS89NgpUr6jpXuovjG0zWtcW0HzshSQPBoIUQT2Xuzff8vQXECEY+MHSpUR
IGjsMHQC5gfKSPRijG8f6gODSumkqegnBbRqIhockrAhZ1ghhMRRnurXxQKm2uUy
fJ+I9iFj3eneiT7ZCoKVGw1GPReF5fT00glm3KRuzCeeZvhU82HaZCrZ65B58xfR
mYbackl6O6wPsrFs20dbYq21a7HttSf4mfK/AyIiO9VzW2yOmPOTFZuJ8a8DxpcL
1jn9gZzba4vKNTPAyadMqWxz/zlKnyjuElaHJNznFgXQpmSyQ/2eYyeTNNXASvgL
mlWkBrTBFNUdb48JIoiJQ9y4DIy2Z3X14F3QwUxdHHUVFH0Db9f5NXPj3ji7Ila8
8Lk1cgbp0jHHdkECqSLwgZXTMHleOZswuGprYGZL6wesBPnZUNl3t8aHiTkSdjDQ
Eo2Hec8bl6og/+/+Bp0gfQLScZrJ9KH4HKBtzR3Z0oUfNz93yGtq9l14DFuInKKg
gkUXbD/QwCAaMEwIAr11Jr5Km7oRzYyIGRfAlsDHwFemHeqB6zQQ4V2Ek6z7DzLf
t3cx5akdSl+s81mLsaLxMN9ylBeZbOa1kxcaGFvfBzdnFc7bCMpNWynSLe9LIzfU
BVsy8mRQMR7ZZ0S1a5bY7BgBJiDschNA31JXgDLD60hXwpJ/I1SxZuS1+VVpWkgX
b5TeQB6fPueGgympbNQ/DRn4V0RBtwnBkwyikLwrM9RlqZ/vN+Iy7nw1gU4zs07q
33vvGCJE82ZZncRYDkxK0v0IWu4nYsDO94KSN5vmedrsvcOCREYOg7nBADj8qND1
tfXG1x95rWlGhoj6MNN05CN1Fuu43Jq7MQFsKQ4hhEBzNX5abPiO4hoxNaEy7shr
sLESBnxLAQP9pVrSa+Q38nSDXoepBY5b5cB3pSajhoWkbBdNLmEHDAI1d3h6GBEb
M4ICVlNtvM9B8bU4UkOEx3Lvc+ASRDOaYyVsV4Bk5C9lAUKAqCoI6hK6iQf+Jlqo
oRVd7ohMY3cvXbxAglzZLqFjr0T/u5FCQdCYKYnB5ISAuIX4tCYRQqWeWeNnjlAO
9QmUDETyT+tWXgRyT3lcj0ERQ7A/weMnnfuxjQj7eNM3y69mtSfZ2aSj8jw7CwgV
aoDY1GOs1z0brHprG4LtytUXl51ddk06EZse3yz2dXUM/yUA33l1WoM2nDnRq0A7
LngRHwEfqptWiu7l0qBSzkyalcxbl8tc1DFo+634Bih+WeUlKjOwqfWpGxfqSRPn
N5DLTPnnSbG4y2hDeI1IbyxhoIp9bJQIVH9cwQScN1hiHo0VUZZEPZ6HPyEHdkPX
cwCwh0TJhms3q5/sFQHU2gT9SXmA6g0Rh0elr6I/usc559xiQ3DOJwHjoudSp/ll
7fRFucWvb7s6/qjh7TvdaftG0mKQjmigBVfwUrtp0r87PRyGlR9/x7XKMLvf2l+t
P/C6akt17mWqoitGQQtGOExFNJ+Sk8GK3pacKH5S48hEFeQO6cK/bphutkUpDV8f
wExCJK5isK6h6Y0RS0fhWq78X3ceVJDDLOXweUi5DSx0J/BfL9RkwBKFeyDGVSZA
kZ/gi05mbDvtc/Vyqy3EfehuvLfn+xbQfi4XoN4d52+lJkDqze0fOowqj8evqL0Q
wsUrXjZJSqJ2uTh/DZM4p6MxqBQXt3WQPgCGos0LELFhj6BFRLKFNl9VuGT48wOF
+G2BYZGKuesB6WNOuAU5z4tFGnvHEfCyza3DyFbTmDAW8OrT2Byn7xPSsHOa+XBQ
76x1WioJYP5nh46pMucpBz5cyjce6KVRlRgRuki/3zowG0rcnyJdvmEx3xkKIbn6
BfjU4EqvslXBGpgfz7QA6cICSh5BngACdjo+ezhia9eL9BGigtrTEuPVB0wXG2pp
/jGqNIq1+9F7wWr1ZMBYQ5zMDwSBiytpbVzcDjTkruphAvXWg91ei/OaRR8uyKYI
1/I1iXi9W6UWYkXWrEmJjinqI7qpNVE9BLub9xRgBsFl+Xk86GgO2XFJ1WJ+eYko
gGxOAXJ5iSgE2tiSuFMPmqG7SV0uIbuRDA3+J9HP5NsriQOoD8DzAZdbx8S88jZO
+MkvL/dFeYHBBkYKyn62zz/2ThxS2RINg4EgTJ4NauTEjfVg0tHqsmsFlWfkILCM
NfPb+uDPU2zP/Ff7Lvc6Gt3jpIBLqXF6gNrK6/pOMxakYXYieEPaeP8PK+muCtLt
H2UpOxoRg9RSuDbJ2UcdFqGZRhm0JlzebciMRPENM59/wXeRFQSZuBDvmhc0aQb8
VKlM2SvG8DaOuM/F22PkVmiqUFrqsE++5Ctc7HepzMKr+KHkHFBGpkuDDJ0P1ccy
OtWHAkCJft1agLiuXHuCNC8VNiMyMZXjGlExY53E47I5vvCbEiEVq8DPvUDDfx7q
JI6v4wvLGeOxLMN4lCY7LuYFNqMl3fYEhkPQOa6wjARBXa0A8BJ3zBi+0PoAt/wj
BsuECUcWQ1udKt+pkGksqj+M2QXc/WV20/3axAtjOpt28S5BAF/FK2gtc3bjZnXo
IgzwRb97fE/ua+uHlinjACi8z/IZffc45cpXx54QGgSsks6NXFKu7Y//7lHhNj3U
Fn2OMW/hdu33EvNGBBJpVdHEEJDElZzbCK+Z+2hyhiMIyFSzZ5ryG3PxPUrI8axq
kJggwBXH7bs2sTmB7AY7lGvcTjZZl1aVSzBNdX8cYcIHW3PO8prs55/alvvr8Lbx
UWsiFWDIlHfvcanihrmmCNoaaDWqdxjzoJxGw/z+YvnH1XWdYqmKMBWNftVU/20h
8Hqjj91uvcV90CgLzgEE8qYEKRdoraNjvGTkgXzxW/JaDPXuVu0btpIRlhUWjl27
VUF7Fak/zNjaUkJq8R87i0p1juPiXMsDKrDobt6FcdpjJ7v/PMS8+ShXXwxagFhJ
jk7EqDaY5LiYwl5zgn0Z3JupvJzLDhjgbSqMWhTjiK4MMxuA9BEITwENqdltf0By
nV1pXRtsIRtqe8vd+N00So5a9oLvtguJqhq4Hx4VbC//YdP/qUVppXwfVpFDuJyf
p7XIevu0fRkLSC358pWGP+AtFUOHr/jTcCqi9SPC77KmLvuMKgN04GPObU9dspkI
eX06t6ul/wQg2/GVtSB15eY7fO2OniEDvWI0PumEQoKhhCxti9HoYvQekSyGpnkF
kjMsccza682Ln6BIRiVBlbUKxp0jxwxTn25/tsRTKO6RFCVsouwc/mq8qiTMWM9O
yUCtgdUMj99S7eUQan+56IZ1ae8TzVldulKzSxdnK8OClHTj5L3MTYNQmfMaZBEf
BAF8TcBIaL49YvBOCuchxGMGOVcZC/eaKacstzIxPU5V5150KR22Pw5MFf+IKYeJ
DJXXlMUKVSslpPLwzrYbPjFNYnC71B2vdug5HVsSeWIXDY4oOl8QPLtrZc7wovyO
vwB8RSlZwvIetrZKCDzeVef9PGf/baGlANZO6GNqH39qCll85ZOVxuGAdpSEXrPC
OX0+O4I+LigDsCzv6maFoIVDhfRxCihByrlQrMIdYa7J35S8hmAzcr6kLciib1Pi
L0rrWbynj7WfWCprvUosfGL+w3Bdtge+f+4VHA1Bjbt5OkBoeF6bPupKjR0nDkQ+
mittDENd3OH2yumWla1ZZrVwVCQrN0YeXfZsGlNyGxrobbw6tPfGtxmaA0ddlSvg
/cwNUV5b/G8bSUmQsldnOt2eutYi5/jXPJw4U4BR7Z4c479EoHKY3FOdwNgyYYHK
5a62ZeMX890dsHCMb1lq5efLpDE3HlwIExnq+qOkj8Sc9CWearo1EoeLxLa1+F1M
Krs0hio7KDL0DhelZQ5kktmNmkSyCTN+TXnnQ1ZTnFo8bjp/2oDADoxjC9Su+6QV
6CokcDYRsliy0eIBM2Ej9lp+RhU+FTQ4iCx2MLVQJVPqDqtjgFUz1peLE0yeK6DL
uTZ/iJr976oEQjhhoTjwLoj0vTBefQlNY7cKBmbgPTOVt3C7NwZer4K6T/310GeS
PAJ4xGGHRn3Sn26UB96cIYuIBk3zsjZ3gqeUKpCqTlY71174Nz/+e7NatvGyrh93
x+1JVGYQqaJP70DLXAcJKxh2cBrUqeb3+JyIPzXUzjRS5gvh1reJCErE7FaXf7V2
3FDhqGcw8Zbr9z0tDVWjxX/05Ts+4BZGYCHbBebSrwL8h2HFne1pxD5vMNQTqlCt
VO8Cc/BOgNEJW+KAjOwV+dXkElkl8qPThkX8v/xRTG6Hw+Hk/XkGyi3nyrUnZy5+
Vq8UCvcU2W/zj8vFvwRIJKDq16vsNoOuJXwStO2TQJU34eEpncwS4CxYx4vD78Kd
JCXAWOYPm2yCve+HEK26tEwjp/bKGKanVTmi2bq+MYeIqkS/mzigxbImcjggFSl4
tDHcLQTLob3cK2KoqbWFJABlEG1Uma3s6Qvh5GRptd7b1N2cewq1rcP06ubKl5Q5
OJTO6CYuEoO1SjAt4Q0yIsuWianeMel8TSLJWapHGhiY/S34T9b1ybnYJ4ka8B2R
uE2JYutc5BbfHp/14Wr/DfPS9k03rvzDyrd6jR6S/NOYrzSJ8SwgM5SoDZYeJf4S
h4UH4iWjMWn+l/LoJdJX6ZfUhb5az/kSCkZ3sL5q2ejnTz0XHP8M2ouslgGsZKMq
964/cidST9Xc1HAqQrK+i7q9y8nHOXwptMwIUTLDjFghb8KeDqiSC4Rbh7N9JXkz
tui/7frTLdCdjD60YU3mkrT3tJyoCF4kqKTDYx9WgdBedjkRUQgMvEkdbe0JQeN7
SravqdIN7foVIUO0m9HDRe9Bd1e72srXN7toGkjCUQH7EhaAe227EtW46NMAFbY6
YGjtCSaa/qj2d5Eugm5G3LuqW8oVY1RblOrrwpCg/WAr1b6msSnRKi10amhck6gs
r3qdXW61zS1tnyPLxltNwIEk0PlSYvHQd1P6qUb/Fa5PxTsW5ZkbN0+IP7UW9yTA
fMohnV8SItLMbopF01DgRF6LxvkRi9GtATNdpYlZxKn1nqDXPadmGOU03QgFzPSK
0fAttGibQS4sGHUTPoH888XkJby1TgtTwOZTGLSWqNXoWmCzHxyM9xlWZMdG1+SA
PmrGKHcWotrV/jR46Cbcgmh7OYmvio6KYclot5ptTsq/OAeCwkxOxALgY09jO+jC
05lcxAW+nUTZjw1wc0RA0l/Q3QZUiEYg1jYENChSSYn/oT0WbfBsmT78mL11CQ5m
mxpKhytmbfSuk3btur9YrhRdz4tnkVo+couulXdzx/YnUlmQ8Nybc5ihDxovKKyX
OEDbEF5PZVMp9lQMtg/TiKs+tRD4cj8QltxvH0asno/xoWCk+Cp0d5Oqeik5cOKF
qs4rXa3ZG6CY9A1RiNyEfMkodqB0wpP+EzwyPwLoxl4kzXnG2ZepekHljHq7d+dS
CzDO5FN3nJfyNR5TvsNuMQ725rZ9MWu72D8WOnzvvs+RQXQlnp4+0wfpTt0vazWh
iPoIezgPFwqm0sxOA5z/KR7DF0Fhn6IJ4ytqj7Ylw7Rb32Xuf+IC/ftA0gyw4FQT
UbBjH2yv93ro2C9fVLSyb4rQGKuzzoFXdVRtrlPnTorGamcFFTB98uB7f/8sxU4Z
NlR59TqqRsX95bCAJE7+eu1GTAeUhEtfyzXxF5KVCzClbef6799+eamewQQqXxK7
ALoDSkXqTZQBYjQuUGMpQb1bTHrpGyjLdn4h/BfD6jrBne8gdVMpdV6HsWP4bd0G
5tWEyyupv3q0VUvFMcUDUzSiTVaqFv6kb6kFOqh7SU0IEvWf6ssvyCoxeYohez0V
Xvbsm/sebr1Oh1XELJKc3bAlqvZo2OK4HqECEd8oRA/mNAtCHlVEInxFLlG493Vr
w2cWi8MoIFt6c9Aw7U0s5RfGaSwFH4ZLPY/AVfIuYVeoWnsrLm2oZoqpfWVZrFQy
yZ8lfTj0F9q1uf9GAXKXOcZGEKIhc8OlC5IgILRxJ/e6/U6kjriTcEBX6DJZn/sE
F55WM6oditopFzLBo8QTuoCJtTebNsk4kx85tHEEM1JivtXh1TA92o0IF+gfOVjy
dmeJMATtqP4GExz4escVe02KcdTSvQJ5C3svDSjoIESwtgrUCGlVzU2D5AoULyK4
5Ga17YoI3mXj/mIxd9MTEF1EbehVdyBsvd6R34wxQOmMk0PQqts6hWV2PjoNp1UL
YmKXByShohEPJw+whpKZatetpnXFrSllJOUFPfv+EQ2jkd0vIwaod6AO9JWdxdpS
Wc+7N3JT9vO3a2F/TIAGrMyWjGgf7naTaXY5Aamvi7utLIOuglpgIU+i5rwDplsa
A4pY4a2uAEC/uIIEOWS8wOR9hvm+l/mcCwtHFz9HJqhwFy/Xecv76Ljc5G/nsvB0
ajGm/k1A/dPtsuKlXUbZGJocv+zT9OSF/U6OpvArM6deYe/a1mjWuLgxlGnFUruW
eV8dz/mNGCxp9QNIbYHDrXYbKN1SP1wmXrks2iuAlK9e16shVSmM3HcSdrN0h128
gEvfk1SxqXf0mQTeJkA/NOoHwOTOddPg5BwHxKsCSZhmB+svmHUlFMAZexFTY8ms
4nQ3FrIxiZjreBhKwH9Xp6mftceGManAIZi9GrTtLD0fCp4zW/EMzRy3DuhfetdB
6itrRo9CdxmTaFlv4RokNk4Pe36FNobgyBpD/XYIY5WThDaQ5+K7luZhgzSVUmel
wFAYpOJMztAhblk5imZZvPqNwrbcqOhAwwx3HTutnuS8+IbRqg+yJRGcHrG+pi8r
xwpOnTk/ZtoEIXQD3QlaCjFMulIISWFKoNSx4OQvOvJdlBjdWNozL0H1iAYB0+bN
vECrgWrBUE1ppc8lZiwxu8vo1g+ikSowr+cyOrucVEzHWtlKfyDxkiEbDOewjasm
VAUeFKDVayyBBG3trzO1BuyDjhgTkreSCLVlXp4Av0LEamKygdvidGFxyjOJLAje
aFyKVu6kgkBjKoebyJ3rO1AiSA3jis0XX7uY3SNnKcIXDnTkvkMDnkY5dt9t0vot
3t5NdlURj9ktlSIgTKKHTzF0dDVB9VweF7OyTcn82vv1yrXYyHXKFYRGtIMjISxB
M/50pViy5qWboBK6ry5CQPLJxLiqCD5igKG7y730A5twdti9sDZQ7J7GZY+xwgdG
5BXj2mECTD6Czir8wRFnxZ69o2gIJ9FZlsX7euH+8tMyWBfiytmWex8L3yGtpjIW
Ou5zLPWv+NUOByplFvOQKIyANsiZqlcMDGkDAjLiovFnjb0xQ4C5bhxRF4ETfC3L
D1uy2Wde2KdHSJFhgKS6kVgY1SWIyO2nmLunrnOL4XoguHB63f1tAQonZdb9cQ3P
cymKxCAQnz7xgyVk8NNV6FydwkxggPxGBqWKDlKKpGlnUBZSq3ogRSrSyKDccn2r
TZYIzYsQYEBSwJTdxfM52jpicqYOgFI11HcnH8qZNJtcD4+9QY2YpLmgtIvjuBhv
F5KX6JZREGjsNz6bqUGqk8u3hm72sF5poQfK+tFMBASeYlPxTtMqpzsSO8tYSKMa
ym23VDszLedC1ex/Ffz+6sj8M9nPkxPk5ko6TKRL9ZCByCOOr/S0IMGOlAeqlwYm
1kaVgbfFmmINiBY5k2DoWCLbTfH56D4szM1hiR442HsWMWwIVoARfLTczRAeRdA4
PXws+MRVNGCslcWQQcK3aXSC/zJXflMfc7fhRgwh47pRyUV9QYo2JY/dCs9kxm1q
v+BG1vVOEtma81Duz6oV9aOs2VvdaNi9TeKn0SycbJdaP5+fy0V74mVy3IQKjq34
wKhGLsxacG83RrJ3uZ12iQamXfVPE2NbP1HLj3/tv6hs1Segxu78f+AKXy2mHsTj
R5wtfP6VDtGdH/PFfXqDzmOEpKVL/X+tFLjTx0lu3J7bZjuHeM6DJOr9uASFp+Lz
xoIhJBA5wQR1onRiudJ9BWU4wyWhJ05zvSxJyWrCvJfVPX8KGAIFbCFwZn0gO+nZ
uVkPyxDlDOF0qdcz27pSYv25sUBzL24cGtyfun4bawkaSGyZM3KriV2KwM/bWsmn
nm3MZfaQKMX5IS29/iQz71jR0s8Mzx4Gq10FyFinWT37KtTyRWLE+oQABoTzKn/1
g6Iqw0T4hz2ppTm8Vutz+oIIF95Z/ap1jMGkkvSVL+VqqRAqkXUIUs/6g/KAnJMe
cRy9vuF1TjfpsYbBFznYCCPdsVqFz9E9RfDP3T0IlIkO09dGIOZ3QFqs8tgJpvoL
JlUF9YGOxdHuXauo/exC5X0/WU+6EVRlq5GsI5ERSlWLXYbyk2xgn0txo6X0HR5l
7D6cWYXTSjCj00EX1wmCGiwjf+EnxU5KRZJj7/rSFfHUuJbzTMF3QYVX+V6JwdLh
BKxasTfTJfCro73hj/5Is7grePH4hiWBZSo6JlarKMIgCanbx2tPo+xRyfDRNRfI
xLsc17b4AmNDmNvkCDUsmwJTbP8hN18XKb7V1amSctdRGjLn5UI4oIwAfEZQYb4N
u2B+vK8Pwqy16TJ+zSVFprm+Mb8McXuSyc9HrtqBijValbyNZGMUQu0otlVcIyRm
bDoO+pkjKixp3CGTilfkWcKktbE4BrPVN/VacPaYBlURl+7U1x2TNtCOQvaJA6Zf
n8377OfHexorjQSW2hZLppkEn6HXZS0eLCMupuZHztJgZnuH0xLKMXe2562KFkND
ywtxuU1s2Nygj6fOV4014O+rqgfks1h2Sfi0BSzBsJnsAXugy5p2WUCDas7wsp1n
Yh0uzTGkIickrxqJJrw9HyRSrhcATvqRrBR8u+YStLcutOp8LAMSyGNjXOvdWlgs
5bY4tNhPAKO3FfChW+J47OyeBJFymIl+DuYvH9rtF/iirh0jtGf5dOvlLW5A8lam
LQYhSyPIjNgkp3p/Nv+TFBf8aQY3DtP1BMHFduyafE4vwNxjqzvhaHrjr1U34vTg
UbPsc1zK+PjHihaLn7tNxsUF+w+WAH1c3TvqSwGmhj8cRzUumVZR3YcOp5Og/c0d
DEXi6pBklVwvuhzPLwsERbNeYv7+D3EpdoI752NFlq/RJzfUkAhN7qcjcSurTG2Q
opuBToRPCQ2BSXLfmY4NOjIsumiuHXKbKxgBH5fcCbhd2UMfKiJX5ZRvCerkbJ4q
nW69ws/kgZ/TgeQ4IqyKLOnCuavqp6PBHzuE8rXXkCA3ieFm+WJO+lNuQllkMvTF
ScvlcOv9wonFzqlFlC/PndjGyR1ntOHqP4G4ZC2ideRFsJ2Wo0EC+eLGhRpEZpVd
sfac6KJ5jFWctB3KqRSIek4hFScegJwEoVyCtONfTR4A5gDyFIrej96asYJigrrY
NjBiBrTFHPHrxYEg8IkwN0VvgjiclRQ0QWfgq7XlDXvxF8d0F3W9TB3cPV4i3kpK
OBqdWT02/M6E6+WpepJA/2iK5ybe8333ensvIz3CShuBXJ/dDJJQoe1N3rTEoPT+
vLbgQsqAhylp8FYNTZn7Lu+CB5UWdaEYRCzy69NjEFyu3q6en3fLtr3Q6S+hn4Ie
vURAlIIjZsHqlC/YztfLmh59XVMX624plv0DdA2v+8LoxtrwNx1u1o4/W1B8Rf3J
RODkry6/ApTdUNTcHGO4DCs3rVc1SClbpYLuIcrSKc1IFqXxVgwuLBzsIVhg9Xkf
YI6rjfvP/fg6y7456DNZnC/vml3yczAbhDMfcS/zx3kgCdxsFENqfpppzwNr7otH
KyAj+qpTpl+sCRSdnx/Qx6olBhCvO8coL+HIGtAUga2VkWTtNl5R5dMIOhfoYqBc
hqUt0RVt1GLQmiC9P6bTAVfWWqjk4j6Uab3MfjgqdsnD3E1waTIgEEt75QwgnLRO
DN4YLXBuDO+/E81LxC50Ev24zMZHYbdJh9jno0EgG+hd0458KP6X8EGmw2wUwTTu
j1e0HjtcvoeA78m0+ZrXJtQ+fNDN2LGCeHJADGn+6/KxhOG2DrPTaAKkX9oysF4M
WUlPDNOys+SR1eDhTX30mSjeAcpmZWsCXSZlzC8jJlfkW0g+IcZDZXdpbDaaCzE9
hkM9IXbcnZxBMRc0Uqa+zQv8g9oZ/2AtZK4Oe7Wsiuprp/BEiFQCzS0nRqYpNB2R
kVGKubVtrViEsPiNY9ZMCqW7jZPZOAns6KFR/JuXRm5qtvUaA9INrxOBt5ojbNo6
FrvS+yooHFfmRj+SHvyYJ4dY07rDmtgLpesA1KFCp9LcYKvBWS9D17DoKJS0E8Hm
np6euvah7viHs7kQVoTzpprMWahndO01Z7hg/0cfEplkN7yzYW4Eq03NN1KA6Wst
NHPl0bf/9VbWhe/VDhTCGJ+RG2cwsWc0N5Twg0D9ZgqVkRQdmOOrOFk7EPm6NzCe
vUEppJoolLUlzF+4+25wTvXdmOyUnPvq2clRIHDRKsciejJo4J95T7NIlm0fT9WJ
EWNdhbhSLczitIazGBC9HeCkJNVs80zTxgo2HZXu87AdFHem8KcPcMM5FX+5zhn5
bw9dBgJAqw7mpULOqCpqiX7ENx0OjMZWEr/qblfxRTZj8crGJRNOil8GNgT2fEOB
1J6JQJFuk6QKI9C4SnMfKYuB8vbmNL8UgVWuYulqYENJUl8ArjcNl1SNtCbn+3aZ
cemQZwXfOQAvclJ5pOnQ8FHAxgtoGtDcwbRWc85AxK3ZYBSNr6m1fahsrxiDGX+f
HbqpbR1+FLAsoPijNzqJER1Ly4k2MXUsVtRz+J2CQqsPCmAUyVRr8juAeulJRfHs
mC/Gd7p53ax+y13rznciZo9e5M7JN+JMifaYx6nHzag22ur1TEUOFTS+MAqzSjQG
dMl+iEgu34b/IexSWDaRhgLVl0jlGIOqr7CcrBOb2E4um5FFNqa6kPoJvbaYS6Ds
UMLDlAQxZKql+qyyIGwHmp79XsgtFMGWHvq91QB3LrZMnxp2YoKgHyUShuxuSEgW
PUtsZYQvk9gpX+akKrQ66nnWhZMLnYmz2O+QWp3d+kwYNf650N2lQgpkyjUNojTE
g4QmSR7F+UDn1MrFa108wJUyJeR2Ml3NoU/RSL1YT5CQ+TPPcOtvdVRH7bqJ5Fys
ko6KAbhLcwaTryibPEJFTtEsMQNZqXrJLkIhqzNTpAktkKYRBJwRvjEwpZnobKie
rgF8t+5BuC8NMVGZ7ip73PDL4DgV5iAP3Dfqunlspys3J5egVWH7lOTdt+C8FxGl
tpLGzGdPU2RtRDSP6Oj6rli6hWfvBaF2jiQhm07a9Dx/PX1mN52K/Dy2I8LsrVvN
9y33qqHYecAAaenbavrMIrCY6Dna7Qc29GD8pCvVZZAhTy6ogqbCyWw5a6j78ep4
cYFSBPR39qVk3+Ygw55j9p5wPIC389UmnzJtAoefx/6PFreYp+y1VhAyYJqt+rk7
+L/CAz5lqvvzZekIueL7/mlEWP08sVMhch+Zz0puSHmMzJSBSVGIRVfioKy2MpdF
xwHFgvib32wTLS0fcufLhcWwdDqlLmFjpJIOcmcJYvDOhDe03Rr+n1SCEZsGxGEA
63gmtpGZqQVYYkRi9yZ9052c8KOb4FWSynAd7r7MUpYw8Agk5WhZYEtRF77v+df1
aAPD3wtYYgcUryjaaJ4KO3ys//pqzz1rT3/0TThqJk9yBQXdfebwmjadoy6xGS1R
SybB65JPK3YGNRAc04Y3ijFfTMVztrTozTA0TcpW8b4kyC3cugi6Wuv7trF0rmzk
iIGCGNu2Q7StYhS3gTGdeVXhjK2tKu42buZ1RxQv6M/U6Q82G/u873BHiokXScfo
zZly5bP3BARjhNrQtmEY4NMASxb6bRJ/tyMbOjdAkaGImxRK4mKSHBV0A7qoZSQH
KWfRqSU0S5Pg5rIdlpkPBCOOKe9pJHHAIb+PQR/nEfOBp/DKsbVf5TEEN5emSgvt
45qLbQ5inqWKd8DMsAI8YQY8jipcQb0RJkeMUfcbnaw5C7s8n9O57Cixb8eDgJJq
bnivQD9UcTi/eIU9PnzsxZpS7Ds+oBCX7re2o2k5v/UzzJe/ncuuIBHTDFb5vTx5
8kof15ZQxi4IPjXIL/mzQeu/s5/vvdMN/EkiP6HEqcka5959tz1mgp4O47OVydL3
FyMT0SvhHS8hEEynYxhxYBGnFT5YxDogxAQ6DguaGDPJJ6zD5Tn/vdiVdVI8CJny
Q5uobhBaTZU+8rdwrnu45QixKaGbRXrZ3K4X0H68ewKX80ijBvSJSDZtUg6nVZMH
M9jrbJILg/hGd0HzsbMqgVeGboYXZ18Vv8W0lYiTt5AKogiERN1aWVlrVLGc2/kI
oc1KEx4zJ6n5X3DIZywoXn98pBe8/bbTk6vb9464Ox92rF4BDRsKCmmmk1BqIJgk
RBE0vOE+hMs+didCJERhO05onp8Lxtxgh4wkEcnlNQy3vSyIVfN3pb3A5A7W0jae
qvUjSRV6/xT5GQNf5A/ft7tAf5enU3Q1uQByaPqWnaBdPHwCuB6Qhs/DkFHQzj9W
/YLn/cCRcDiPIc9p04K2zk8OFgAhyfIZ4sLY02dMThV2xYjdUB80qdUTtmE5o4Yy
66aTCwHGK9IOiDSDDTF8bpnft3+HWZuPOxFdin4mxGzLAOBKbAFNb6IKrA2zhKbw
7424LJw/OQDrws8C0DXQNrch9JYBa8xTSqi4O8/oFh13pLYQyDJehzc9IvUGOqRH
LeQHU9ZsyXt7HoCmsuXUL7pmlhvg5CRxHrX9xAljResrctTxaVHEQ0TpTe7zdAFJ
YPGsEgnQfHFiF91Ty4SPKQ4qHXXx+bHCnDVK7eiVgce3GXIRGjila6xFrWSgRLma
UGfM21mrD5RZJAvSRAsgf0gItYkfsaJq1WVhLOtUauuY68cISds3V8i//YtSufVn
Z1s1POo1LCxZgv6c3ZwPcMzJxELiz66pnwX4OUIGAt3bGMXYJElYdsQXZKADmF4S
9AvmiSbhFvQJEcZIYfU9bKfjfYv4pJvfGyR3LUfyjHFIevlHzJdhgLrKMbkgUHdB
nq+DXdYri52eBR4SJ8wHjKiP9bfhXfuGJmqYuph/blpb60pkBG1jjlsMC6Xo/Q8x
7hoTUGhy3sgvC5HWnZDVThD4cQ9vGAS1TVdxgbMCi/9YKCeCDugpwEXHXyipV+Nx
OVxNaAbUv4P7iaCnvNORCCaWneHxQQE/tB09WuDKmk4jFwVqc9IAdP+ZFGrQhcuU
anFYev6JgMYk26yOUusxR4mZPTtHvG8Brr+K1OqNBt+GFLQAoN+jzw+nUpvCcbe3
Sa8gGM6eZrsFM/hESjpdKqeR7K4FGNkaL6caeE8ojR/m7EmslHGC7l0rrjg6YReX
qOmbpYDI76Up05V70OGvJdy7sX8GMOd/D4UwpAQc8jEGPSTAh/gl145wtx0MBywn
APoUaoSm69XHSdpL5dQzky04Mdou+8mRvMYmXqAqtMbHrgTWLGtUfuysn26mLAfN
A87jg5kDfWlblf9FPvMIDmXguJnwGNqCl2KiCb2fiPyiHm6hzJRzAXh/2oB2u65d
p08gvQWNe37WpinMqbEIYUwTcQ9B/iSMZQQYel1MBW2gyf6vM8rqwPtA0S2qJ+JL
WwiF7q6dFvwgDAgv/+pJKXlLTA2U4q8FOZ4wKyDjIOhtxIcwjsl+usxTaTJqqFLW
uquZfP4iNv15L54+PDpFzZdv4QUmdkr+wFPd90wuOtZ43BkmdswX9oD7URe+KOck
66BjH8sSVhuciDiLCMybdBIyhx2hP7FWaulBTCzzwMnOAzeYaPOQUhtWYeterfqZ
WURden9Ln1pdl7IW2GDEKiyLcEgwJk9DNyBPnvD9qBPkDKp2oVwylWygxS5CCF58
yHmjZNSfDy6AKrbnKe/HCiq4c1u5exWO95/WEszCx+lBMyJiKzjMGypooXKeCrXp
/uRio8Gp5f12lYFF2BnKiUE4J4INl2HC0p0AQMaoF31ClwoXWxnc8+YstmK9lfxu
UHNKjvhpy3hHgpv9ZP1OgdSD1jA0Il9Rqzu5U514NlcAUH2mztJMBU0tGLUafRoH
8MhbNr3P73DqPiTmzBnxpYl7jZDvpFM6Zwlfh22y7lI/CrWNoRtCs5Hzs4lZPUDb
6oF5R342/w6CnZIlBT1rsFe54BdUj77zsELVU7V7XfPWo2orfEaDIivGz9GujNXg
qChnceToRj4JqEzGvD42mL2SCaehJRwjNPUeZoRLtrX0aou858F9wtAEAW0jupzW
plAmUiHCuQNatEugG1M/Dxy9n1++6rTySB/fTNyjLOFaZQ0OouAKkx1dF8IJ6A5v
38uFZa+Qop8UbPwXjiUvltuYhKLhP508uzXrdYJ5SdQ4iDWAB6DpV6xfnsnwVwxY
0TSYGwdyfr0OwZkI7ZAh9+uALCWbGDsK9dWWkOukg4QHxlgzp72I6IoBljDVQQe/
jwrdRAxkSQnkpsfXBYMuVBlDy596P9apmvEM4OrdrQ/GNyK6ZqJNaoEtR/sBnOIQ
vcqIeEvZ1lT0YWY4WbW16u7hHMG4svQ4oDHMPYZQ0xpY4BwsSJ2NMGqmiq7Eq2pg
cux45Grl7bYJTGqoy4zl37I5AfHvj7Rb9euuKM3pVNCUcGWK+Pf1JW8cpqRJs86m
zAYVGn3ag8rdfKbcgLX7JN0ORNd3/SeyGfhW+MOHJQD7B0ZySFIA9oK1zg+Ptxep
WcPq5+Zuc5Yv9wV3u2TFdR5rhFGvhzx46p1vkmlWg/TfLKsn2x5tVW7RmIxefk0c
nwYpYTLT/+Wnj8lHv2ul7+LQKvdVIHGazeiocKaMwAyRvpdBUUgx4HxTFQQouItV
VogxIUI30neyM4c3oPIBzHFwHc47guEvzAl6QJspQh6ZpiCkL6wF6NFewg06hYRm
gFJAUAul/PYFZs376zkQ4PL29SJ/0WKvTUpJYLxAPlApynNYofhx/Fn830d7jy5p
3UCXuGqTWzO2mgvttRo8t0TXI2ilYqKi3DotwNO/1IZZfG/+bNGGZeJdnXy6B5RK
DMqnd4zHn9ajrPXcgCVeAB7ybWJeUiAA3mjJhyTEdFaohcmQwzZyooMKQ6Pt+MRf
XZQcVKcXCV1N58Zpgx2JrsTLvQoVjTIkQ6WdXdEOGMWKkAjJm+JbnUmnsWFPeaZr
HLPiwz9xTgDSzP0NZWiuWS/Eq5dXxRyCFvoa/iQfDmbiNFrdZybP7uPKe1cAKi5p
oQwTWuTP3pgmAVrEvv+kVsJK50BBxTGLUTIrGFhT4qgrjaB7/P076nUOO1f4aD9W
iOY0L66k2c9oWHleWiC4LfxeE6JLhq2OXbZTI/HBUwilpdL19vz1QKFU91Ca6zTm
uelhQo8bMzNpHoTE/dW9HAKh7m0h6r0OvosyuwrBjGlkkvW9X42SiUBPnpZ96Vih
SjiJOssdlyDPLEK82Cj1rLFfs1smesMP/nIjm5qvH72xrR97ia/UlPGIHkyKsD7E
+iXmRSzOJrAl92icqOKEgkb8ih5g7v72fhxsbzA3vMBGLSTwuMRW2nZJx4eVpU/o
1gdrowVp0+tLP5jGkaJcNspA2bdPWyYfMrz88uaoYRu/zF3tY67MiK9fYT4XeZE1
rMYwg1TURFdEjfdiHBbsI7/LJjIazJkn3apoiZqqJxLmUoLt07saJYRxQvx1MQdB
eKOGOi07gz900SyjDnSHgqdaMy4gO3ByQt4jnKmmQka/R2NFzrxDMQLBaFpBd3OJ
Rzp83PT0tcPPmMPINpOFSmNH61GJXTSvTNjRVDDPjIBy4CQa3d3w/OAc1+e2aMKf
RilhZfVYFcONiz7ckX3i8V9rgErq2YeaqbyqIakPylXfAObzNO2DeGD0MHMvFWVU
UTmchcESnox+d9DPHQve0m7c75yUOGuX895uK0jKUc4/uZWDIUSm3gsVCN4SwfNp
satuD4APgmL6xJKlw/1EJokLWASComWvPVryyAnIY6A2NwViHHow8ZvLfDuEP3Pz
iUxFzWlTchTU6ZVUTlSFMH5TkFz1l1YmgeLcFZ9x2YaflLdUugkQ7l8PFW49DTC5
SD1nu9xyGggzEAG/UjCC3rEc6mTgfGcy8YmCxkw+MDeIrWb6ybkIHpVWPlNQrc2o
z2LTJ9pIupHeI2tH/weKulGa/SmKm+0qjXvX/mxD4GeUZNzq7VTcmMlPbQD2dCJu
YTFBewIixYvhBsKb+u7NBUxX7sHLi+aSkZcb5ZcVM/jVhzL5GMosP9hdJb3eyd6X
/MwEq39r8beLqwz5DbyWwZVmyYv6Wb1uuiYHMegEbWLDxXk4/xWV+F8wxmXayn99
YtH1+ztZkLHPni4jP0qspkoIPKBDa4M+6I7881DG8XoND/pPIoDGrlzGyEkl7P8+
tgM1Iu4oW3XTaZ9eKWbc4vBfZpVmoSM1xgCu/jjUt21HX1UPeIShOBieX0n3pf+O
WZ06ocSnrFEu1mfzR7toM0Q4ik02071o3SoLigWXfT8AASufutuSNAWDDbEs+zyD
ADSr/ajmA6QujqTq2jzks1COTZFCpOeES0zYWj2GvuYGknCpTfPh8RG80o/D0vRD
qEuogWuQgmQiVt8CD+UvuRK0mCqsj8ib5beKArVw77JpYa47tiwNjZKSE+CyK2io
hocSq7rjH4WN7A9cvxHTBb7823Ct7l2+aXe1Dn0UsynsnAyueXOYseobOFdTpztO
jVXDp34ffZT4QTPCHkgTYlLPjcvcrqzE0K41GKqFLwa0eBJwpCZBKcvFh4LsJZ1C
PVrfX9VenEzMXf338jeT69dYwxn0M3NjkhbPR+EMQDJQEYuoz0ny3+CWVTd5plRB
ubK2HS302PNL2GRuI7DigjbiLyf43LvUU5Rf3hrzUCFgB0L30kVUr7Ob71Y4fkMh
qedQ90F2tbwRFM6OHomrXiDF3FHOWrAz9SKY1oMH4VBXY3GZQODRzlUR4GHO+3qU
tF/6c3LW8O5hP17KX2/aLrsT5SJM5J3f4lbVPRls+nzo7DlHlOTIQ7wO3i+2yaLP
Eo6LenmJ8YDiDpR4/pIFG/mOr1lxInS54sL2m+uVOOfaPBa6Wka/3BLdsJS27+8W
rpx8ABkoiZ0FQ+/pB56drA2CMji439fiB3/C94avDIhUbDOGXoZU5GqPCyuUeCtd
Y7d3BXvyGOWeJQ8+FmrdUK9OiTfvvE0b0XHU+8EftfqvzJo3z/2kldZKegcuklFq
+GZK4uKU1tuj9Wna5Qbgcn95Yx4neCdFaSY1+c63PBJpFXB+WM+VLKrYuLIdw0jo
1kBmlBZdj65ujxVZVA7jQjIIW+ejr0j51J84KRq1khH18ZA4U/m15s9lMwTtHA3y
KowX0O0GkeF6xS42Y96Iv77o8ex2s0XvVKYZE/EGPMzZcZ1khsHNLSGrgS2vOz8l
qyH4kcFZ4v8cwa5FW4K0Fej7jzi+f+J5/ivMiahE0y/7NNrum21w0jI+QKlUTyAq
oPl10iFUUw8QjmVtcCJBJrByiQn5ubynFxdb4D6Bu0nWKh5aN2yVus8ZtK9K0fW1
8MyXHSHDXeq8tB+aKV5p4bn7D7nvHK+AtapmnyF1iXHxPsA86BQ/59Gf+yNnqZB4
uSMNA13Nqzu/FP17ny9ADAezn0GKAiyKi9IykHNyDuo3GDV36Piw3DSJU9XtSO+8
ngsxHHbHWBzssMI7FkvYm1ZzdC/lvIjEaXdZjstDIE2ahrV9q9dtHk79yU3ogzc5
Z4MMdP2IQeuPibFghL512X/VmxC51vWhJOlTvQcDLb2LHqxkM8hBCY1rksM8C6Yt
lDaI42lzlOAp0Qg/KupZMthequUoXwk4inuVqfSs2LBahch2e877aurXep3JoaDI
4/4vscrT87u8QSuzA0ATRJxRtf6goAZLYIw0wwvHKmgkO1DO0qNDZesmGA1xYJaN
JD/vV9MgCOQu5/owO06VHnwHCbEdaxq6PNSqG2k2oJG4jG/9EaxmZMKxyCbPIPIN
exK6OqTaR4/kZXGE2eiUuZGjRS+I7+H713PEhLEcjsbe5ABlvK9fxtsz+PNz6A/W
TPWyFVWcdeCfHJYCnGLmWchKVTOJu/uw64JwgcPA/0Xz5t9Ukgp6j/L++AyqY/jR
E9HyxHjg/5Etl/BWrOEMRVZKuv1OzSK3m45fLapEbc1xjzEreMc6pudjNL3SZJ+L
IUNYeHfMCXYQSuVvVtP0FfV68V7dMyivIsMTn8KrOao2GolvWoeP2dEUyfk37XLl
ZZx99wkafrH3t9X06zxzk0CYFG7NRb6do2WRK5+s42KW2kEzxT1PITGOPUJ+pV9u
z/5ktIpyDPLn0kkJ+1K4g3RLCXD6L8Dt3Vn2+wMVdh1MVyOcYb/cfh1v9DtzbiTw
XYnXkQYyi3t69T/PfdAxnu/PvWUwKnsM2n/CDS/P+/ZTTTzkCM0DIDuhh9WZjv5J
4V6dPeUFI82lEYPB24Bgx+/oVkQUXudgcI3PDOHURojaz573waSsuYsYeLgTmriX
AOtjktB9XFh+nDVS0UebqrYZUvUzr3MkF9gppOgDLH6azGHaO8Lo55F6IXPy9GI7
7tDJmel200eudH01M8aUKLvRG9mh8ze9WcqwVnPH/nJIDdA231XuOvE4/z6GFYu1
juPdkXzQiNOS4VAAbe/Eyr834BH60PduXYTU2BTPFjLggdpY+Q7J/HNYyWcVRlH5
W2gW8J0H4G4FLaLYhsXHCAHJCoOlgalypwOYcJSOT2HG4JWx6RByJjaMdnX1TRmH
pvXoUDLZFZd+LeCbyKWxGuv0/U8kResn4zcldte0Wg0EKagAToIETj2c/n1FjhgS
CKtSuIsq3z/OvQ0uHqs482NJi2ezGORf2+/R7bHAyMroSZdWtguBAZMQenFd84Jq
OAensllsPwWTb56YotdwYg1e9IGRngrgHfAjK2TmRPugtlLCWozmY37GijDh524b
V9kkLfVTgV9XH481dIoVOiJOWe6OSLzXMMI14j9xKGUGoPuPZuWtmH1HtzolVZE5
u5pIi8aqjjorDUVS2n78eY7NSM9tLS4fdWcLZEknwXY91FHE0Ogt+GoUGqmFQbqm
Nn25XBWc3BW3waP6JcA4k1mTYraIgqnW/rj5fFOwA4x6vdMH7kgYf/B15gi5hgIu
eMknLNg631z6XP+OAqDH2dlCJXIwKl6wr6OZCYLVpmSJA0BybxooQXjpEewp4abR
VM0MKf+cChfYWIz2qTeJLYHJebUEvYZOLvk/DbIVx4kwGqnjiBo6wb3v/FRQpcTB
p169IK4TDF1BT7/UmGgtJDYA4tZkC+XL8KZ2YDVGWMdkZ5Tg5djhiungbFzcmR9e
yHV4yLs+RgcAgQoHVzyPzVl7KvRxbmI6rQas0i89dL8uKePqx8SaKYBkAkQYk11c
64/OwG2l9k+8dlVq1JuIrRMnkfPb2Pz1Qdsn24DeLY4SQcubkrKpJiuGOw7PItBK
sWmimCCD2PwoWbOf10Nf//LiBj+b4/aCYnBmHAsWzZR0TLfmqA2I7fzISyg1quhU
7etyTVopPlTEZTS2DveyriCUDjzKzTKhqNw4aTy8CMd9PtPFMTNHU9d14QQFZorF
8zH4OUz6QeJke9Z1FDcMtMCa3fAIvggEgyB7PMT8UGb4uFcJbPpzbqXvYDAQ8Xcb
MdRx5sqEhWivYdAJxSYn92ZFLDHO6JiwuO5l7d0aTNIKCEawIf8eThkapFkAQk1x
RIBQRxjHZRLme4CyyzYMIB3dgx2OnSCk8RB6cS78RWOV5BaqdDgjiooB8xJVbbBo
noClKo0QUNsY0aojTxjlFffVnPFLBj1dQUK7ng37y2KrkQgtp9uTGep3quqencP0
z1RJGGzlWke6kVvM+XNqwEHYO9aVpdQgaZlAHFokB2VHw6aUWC04sVpyNDjBOtVv
EewWWmwW+3ougM0diMz4a7+FHT/5jagtLS/Tmi5EirQyzN+uwv748K5NJoHF0GQd
nJjVH/u6I/l5D1USJZ9E9mNJ0tfry9hG2qXBWvEfhSjmkKkvhw4VHLIIUpTuaOKC
ZGy3FFeVKQLkiE2hW0rVDSpMdf6hHPK94ZoHlCKBHFBcv0JAC+3H3Ll5ekkx6qCo
g77M7RRAl1vqDuruST+QptqBQLAkh/vEXEtu6hO6YlMsf1MaNjUpXbBCgc2LwtU7
4YOJB9W0JC0kY+ewaxR564MNMS1pbjK5CU6aRH04MwTNkZrTAHQZZWIVjEbfdrkY
ZoKvjqI3v7GkpVzf80Shaew2jxtDgekFxJoNKo0i4VrQ6wzpxl1h8rrVVLauypv0
AYABHvEEdGagGF1yfpuOI9CREOmpRCrbYboNxqTOMu5A2CqoyjR3bnvsAVXsaU9R
xJHqgBgOyg/y2YRBxUG0l/ql1hyXGxnD7rJRi7Z281eMeB/K7tBde2L7ybheZc2e
t/tLUTHjvAWk9P4KZPiwFWr9XJWX8dwLRHwTQLz35fc9sdPfBdk2ZjRPL38k99/G
QlABYAyvsNZ+l1hg1MU9RhsV61cFKGO112KWkYkQdXHq1oEi2L9ZCzw0DawuKW9o
zg8Gkp4WlkwYuvKjNNNKOyPLWL57XrqhGU6961Zc5SamYm6xs8lmwYIiBJwv0CvG
rXK94wukfOgSn6bK4U6VJvOVjrXQtm+WpeuvEr6cG1IK+j9E91p+G5eh1oNzZMjt
UXSV3WOPLyk0cafc/rU19gq8/vXDSPTuxHpMjaqPyGf4KXZ0c7x/dcdfdgNhB+D0
YgEcACWmVW0bk0ska6eSfq2JXlsgRaGRQW9GVvSk7wJJ0662SPukW9tvZ3Kng1tL
9M65zmOUcUUYNDJd1qWqsNxmqHZ2XOHfkjgYjqWIRFMJnPvizwd/b1KWa6VNQhbp
GZYcQ4O2/MUIEl5q5iAWUcPcIlektWcARxrpmZQsbvYeJH7II4O3VqfuC/8HN0d5
vHLVYM0VzC2PrCUcD4VF9uh6KBcmjnopaxXTxb5J6Pey4RWQDF+rNBfwYjEM+XSt
cqQXy/BLIm+1rn6TYNPHgvY/ohMAGnEeQE5rYLvALKNxTRaYnpanDskGv5gAPzsk
ppkN1AkWoh/sLCPIRLK0T6BUgtC0NNB5v3iHrK4MRiG7lWD4LKXdTVRXmFNWSLlG
J0FbhWGD8gMDrADOCI5GyYsrdh1St3A5kk4esRecJltBrJ0fsGdEfYQJJjOzBT87
q4Kzmj/eSNEmPs3FPT6Ip6u570PFwUrJXsdfGhLI7j+Wb0mTcxLbFsIbM62e1nDi
tKAuZ8ng8nO6DX/REYjT2Suz9ujfI9qtf0eBImIDV/KPHg9YXfQbtOHGMyCiU5gY
mpbojErgIUKfgoxqwssT1XPJ7bLfA62QIv95sgsPTuZ4GU/uz3fv7nyRTmt7QTNM
qYIqfM4+PSFTpvo1SD7IqUpws7uLJhzHLi0dqHDemKGz5nsScriNYRZqzQbqOPI3
3X2RNUURyzUHY9WrJeG8xKfLP2dnaqRpbZqB1BSL40iYmJ3BzdUuiejzgUW67Mqx
4Fs2oTZPAtgsxmf9+V2p2wSswAhRFk9FxRGU2dq5ZQkqL8f7qRzgfBqMKOb5Gm4x
YmM8TlL74adXxfsNpBZcgg+Zoz/u2ZAur5pTPhczQGzqvZ8ika6rEGDBLQGNFyZ9
1/GKtlg2ifVnSV47elX7NdxfwHBjniINiHm56AxsS7vB2sVA1RK7HoUOQJYF9YOp
968DHaEN6KmMKu7s4+guEdi9EISZbvF7Py7rDplfni30QRLXpCu79HiFEPxoOmca
7MZMEfCS/Z1dOVvhJOPNHvtXXkhGvHlfZQj9PGojcA5cRpf6KN4JXZwcVE1ZGipH
tXeptL7RzTKneVoJmg7aodtKcIdOqd/lzgtKqYAPlkkHwDzbX+byuG7AA4/OO3MU
pinQ84VX/UVWdhBaumph30mIzlhuxoo1JQx4JexMrgKRb/8+DolYdKP3iR/L/Z4N
ogza4oOTIdN/u6wnKrY8uRHP/LzALsisyoE9gf9DCqRQxY0b2zU1oZr9oELbXg2D
VAcvOwW3Y3ok2nrS+Yp9azgLKaRBvMI+7DFtr+bDW/UfQqsVKQmhEkIu29TFvm2x
swyzfgbKng33RiiKiiuGzwo72FMDWWq0IOME2oOMBrbvJdSmvRAgXh0koPL8ceHa
kaBGx9eVgtXd3AoxWtVFQUmYth/6UQmnKA2uYwA8/v2SR5haa7+rqDFM/yU4wuDS
qvp0faxlxTnfJksGOjiQyaiJmux635qa0fIXM4zDCezbk+hNqhFHb743JJWKKadL
iNCqq9GGT12zZ9NIO/wROcbS1jouYcxM1s53Hnj2Nqrfs1ka9fjJvRwNAe88gWtE
axZkjqCF5rFp8AIMAKC44TiwZsqIoWMY7BGQ4jFqCBlSxBDWWfoG0TJdSetERavb
0CQndjZn7WkWIOdwPWeFYZoWTkdIrMofNeTkNOCVip/xcu4JK9I++bJDt2H9lWJ1
j2kqx+ZIRUTOCdvAaF9qQwxAMZFDH4nETMMCW+LqmAw8HSKn53WSyt4B3oT2x9CX
OW1q/kRHhBksJb//pqgRhVFdyLBx5tVNMYAEm8cGFN7YOeaKhFQUgYKf07NGEmDm
cQe5l/tedhb68CWh0Se4jW+lzLNLAAKDPLCipBGQ0vNP4FjZNnxztyGmOU4uPClT
W4u0Lc4qCuCyBj+PAa2OrwYjPL+rXoEU+9eqd/pmE0O/LGfq4YFB0Hvb0mFXqXG0
wZtCfdU8fo5f5mJA2WO4b5pGlabaUyVcQQBAsIq3Y3xjKPD3rXaMajO7F280o6xZ
LffdsEo7a04cPCuWglrv+5PX9cKZAomzFnR9iUIfcNjVytfHDecvYp4wAswD+q38
OrdE1jSYNfK+VstIxlM70n3kUqTR4z0MSmjeni6UH7S+87DI/O/0gUKkgQR2HtYk
W+XWT+GUf5nmzI9HPDi2vuFtVMzjzTOD5eANQz6kNbCAyrI+BL0tdImYM+scbG8I
9pGCP23UGOs9dZd8wliyh1c7Zn/w0zoj3n1jtegUOGgzCpAl0RWBzAU+GMzVi+Om
ukiLAq03miNAi8KULuqWRnlNgT0qWJ6iekPHxV8q2aLwkQBtV4LYdUvZkW5iYyAC
mDg9rZihxYSyGp00OnnKJN2ohwBsdy1qmv/1H1Ku+uZ89l5Ib0s8aAj7lvEo3PNe
jvZNYiqSdNs4PuzT2Q1RsSkIBo2Lgi6Y7wWrdd6bg7Q/K2o75DnPwjTwqaiPP2yW
oj9uD+9TQQ10CMII7hNP1hWWXTk4xIctKmNxtT8jXMhCVnGwMtYYPaMSgxn+pXOR
uRA3WiIq/IDBOdbH3Jb+15cz6h6KtDUv7m2VZae6zom3aASlkQVlupG4231pYUlm
+OWUBxKLGyeR9iMgwSTFU8XworpcjT7PBZBWctvXq1KnhUZFOfIK1FsWpeXVw1q0
PeSV5ZOik3WCgfWX3X1CYQtZ7BnVGbvSY8QQfeP3+LhP6Wg4bJHFfWxJlKIpimpq
AIHpGlFQfCSNhsV2t7fSlfr854z/KlybX64zmEqS/28XswjLRVBbxzUjurS1f/uv
AxVIC1RWUem4m4XlcQs944blXedJKCsX2sEuir6PwzFN3ehIHAwXEx/SaKJmwtvS
s+1lbTXfmynPllWhBL8mzxs6dvtGOC3Z7zK5EyhfwpT1QGe2IbBiJXFuylyGj91R
yXOxIE2PAhIlKjLbrsFUXDcf4BB9h4nZlEnsVAYA6VPbKgpRQfs5nkfDIp2L9BDz
WWkaGbC4Vqjoz1YHZ4Uke7/JyUQqdDzfLMcgr9wt27mdHKR1Hdyu5G+sbY2Y08vC
MLaIUGKrRV8BgN9hN6qfw+U/dbl3z/+P3jn0Hfj9I95uQ3YQDqSS3uslG9BQIQi7
lmLxHzoE4Ju1jJBZVlYdp6ddnIX3K06JqfJjZB7GY3AdRU0NybVQ8Ai1nU7fq/Ug
LurOCUoAcxpxYXF250qy6IbE4s2jlZUoSCEFkRE2kFxqbMb485nMDEz9/nKa0S9/
UisWjpy2wrvuqQVIYzXWn4pAwZATZrXp0cNvHIqIqk4YYGDwptqF1wJnWP/0EmWU
q3dBh2b5AhOuD/o2H1POXsqDi/X2+brflJnaLMvU2lFWLByHKRrsZH2hgPaabO1Y
PpLkFgckSAfff9q+zjKEtFQpEqNmBSl0G47jvx0nPpxN+Ov2IHXsNSZmponlKl9w
vOUPv38ClNBSZhD1LcFjy+E/p8ypfPaHK6tQKPgaWYeW+cBXUCa7xYUcmmI9US6L
9mTbs0gIoQpl25CDaTAh6ViKnB0+U6G+VK+i8qzoO4xzrs6fFlrMaqO2G2AFQeV6
SMPgpaRFZWcqp7vmTgANe4s1NC9gyCFLmnS0zuugUMbb2SeJKDewPmuzo+MAC1+7
O1s3q8VkgGhqdPAUWDt6cWc1/Hl9OERF9e6RDN+yNRX+yObCc09rLlQzDTtxDCzs
QAnUjY5mrGG3arvAefk6dPXITSgglTL5eWTLNQwF8PL0qu5jHhOI2gOcr1Pkfhgs
o+9RvakoM2odr25Q+0qzFgCaRi4PpKQoQ0oyy3A+5gNTKjcyIOvYqAsOHZi03e69
EaTCwjAgqmK2ad5yrQag89SYz3Zzgb6/iKyhbvvK2ZBMqhts+ToRsnyjdzRiCJzZ
h51KLtj4RSqD24PbnZf6zC+nM1UfwgJe0pruuKFJaawzadM7tXO0lLHXUHcIudod
izkeUmk6EG0CK5kcHCT4nXD6gMreT1/FUkwEm3erxsVg5jY4F9tozxVEc5Segj9M
FKn9VuSVJadh8169yVCCWnc3Fqe1ZNkWFMKPX7S/GakGSOr7iW7ypUYdQW2ipOsj
p2o+KvuZcMl6e0aWm+UT81gYUu7ux7B+uEVBfSB8+9FylDx5Zu9RbGVd2gohOQ+k
ULuMUZL6wxtHXOrTqOa3uQHxbUyRTiCZlQ62BfRI4d+hTl/1wGS6sgMxp6w78yaK
WlCV+9XcLi3o9KGYzSa6rq6RYnSDF/tBeI+qGyx8hIVaJB4Bco5XcrYUvDyN/6IY
hWBVxwLofso7vsTjRQhLnww/qcDl8phuhmhbEYkX5f6ttq4WFgawlBKGXVK4MiL9
EHpeQrJhaFwhm6G0TyI6onkh4KOV1V+7PUFUVx7HVQDhxYlhbuqi8eOuxdlipQv2
Xc2PmwF1w9XF14sNFrIbgXNJ3F30wHtnr6ih2HTIoXYBhpjBy0ZlbHVbLGkdU7zm
1Wt4Kj41Dx+lzF9m819JKi2kwmIr1brTkTxpHHCo22qM+37rcpfBQ1+Rp+47YEFd
YH+JfgNXXTbCTBsVA1leBAKER4U7yGSYJZzO6QMn0BbQqmFybJHt8hAKHB2cvx92
NWtHW1+qHHhlOB+nOGpYSo0OpOKQ3dRHc8rQo3KTmdpJtx45zs4wt995ofhhtA8Q
wKXWWouTACma1uumj7VXfwYmjKXQnj3nuUer1wBtsL9EjT21JcpiV70DC3wOYD/y
7z0UD+oTANU7L5IkydDoA0tnBqNx8r3LoFT+m9D6xIoqd3QA46MA930Gs322ryBo
iOgtQHLIbA31jtLutNPNDMWpB1d38LvQhvqHw301AOm2U+mLXfDX6wDblyW0pfpv
vlmzuTKhjKQtQiyevRFK76/9o7tky+xNogRC96odJrBwejNkDz98DekOtLfvViDX
DsJfisXQUuE+uFG7t4f1ILQOzA/Q0VfnrnD6BVooc0pnG679+1axTsq5T/ZF+b3L
AftV8MNHCAuzjl6VztpR7wiK3DGtJENl13IRZxTqUhiMO8lPyyGOfAXoiVpxp31s
lFtQuFWTU+ACwtl6AQq6C5Fzn6oXzObODPpPXdgJKQGFjm4M7FaYn2PI/G1PntUa
/HB/u8/OCKqL89y4etXzu+qjbHbY8NYMLfyM5U9aarZz7/b8MWaStXmwzHEGopMq
dxD6AaYC9JbOuORbGJw27NFLZBgSGbYV6bNSjp/hLDl2sixwB4Q3BbofNa8fyElP
ghV3U08vckO1dFmt3RhTudETEHRVr07Tdx37dTGHDW7zzBrBGGvNSsoxmvbf/1pL
Clf1nds105AgIZRaedI9M5GjrmkeYhhLbb8B1nflvLeWtC9RN0lR53c1N+M9RMj7
8H23NhGU+/Xx14c0q7UNYZfueTJwfjNpWOQsir9prOzw1lXTNI/f6BBTG1ZlZ9DQ
fpt5t4u1ldHKYUnW+ohv880LuzI6pvw+DkXOg2z/p0+eB+dZSA7689j0+5BUn8lD
cgSNiGrU4Ps9nRvz5TWuscw0CE3ejZ0ZEqSVOcmV/dp6XXQGR0iI9lg6ldRyMJKF
7teM86Ap/82Z9YhCvDlBeahcSMCQ8+A1k7lr/nKWn+ne74b/Osx48xpy0mQxwLkN
/AZZTk1sP1LFpI6Es67B5oqq6qXwKzifxVKFIexN21bpuDqkpr7K0zLVW/PZ91bR
mb5MUNFUEYTfheIiOjZGbO/K2VqZPE6PfNJCPLcRa/yLqH6OQaS1oRnH9nECtNDp
Tl6P++lkc5i2tf8/cEsQxv5Q8F5avzZes3VNXDWImC6Z+JUwk4ZoHBFNPobLz+M+
9E1v7Nbs4maxDTvKdWnPR1SwIZVDHhklGCxT29XSF5xK3ymckN/fBqUztBUYNgB/
ZEG1hen7f5CSsWsd+EUw0OzE9w7dM0XKjAkYrsEAVvJKhZQ92TETX00kCCGaglBi
tcEAcidsrwXAd7J1NLwI+19a8xN1GrutWehGBZa+/XcyejUTgXQU+uD4YwXdxDn1
QhPKjzZdj+r0p4+07HnYdqzute3DiAGEfmGTAgr/G2B17GpZSOoMenBGZU0uGk+A
ThYd9tHDaP7je2u2/pap7ccoMDnoxqE4YdJC5b60PSOpUtlzYaBkTFnIPti+3T5Q
4CgtcVp/aMhpt2WTifI5hKwFvovwz1SyeIR2JkzyLqo2XIp+La3Z+n1cWtsTosR2
Y1LaeDlm9kNzF0C4IoKvlAJnizOTgx1N+v4DQ8eFQ4VjcJaHTkkFVTSojU1OSgog
xe+vZej+IJS1/+Fi03no+z1ChtVYX3PHKBG0I2USzR5xi2F0AZGR+6gVvjvufyQw
Ser4/YROK6B3B4uJO3gienLekjFgkehlyC/gy45FiuYeJk0uBpj9garEq6GiMEcH
z2yfhRMLnhYxceKi/55kzwGktD8P0v5GdB+3grF4S4gZ99kg2w0N6g4gU/AqxfSk
9PPxcTODAk1qbC66/ugByt1sarDQscOkAMnBgN7a3zmld86pQOq6t1oOMUWINHGu
r4j89AQsN4v6Vs94LRpR28aOFVypD/Ly1HPXQpFC9QkS/5aMW7tG007oSrhIlfZJ
UQ8ZubgKFgt/zm0DMBQtxFZFtZ5QlfsVg0lWIlzmqZ0QoW+T8x7tap4kk08l9/jx
r9+1SYne/rBaswSPOocUSGQ9X+3folvWNUriIxixD7C/RLz8OIDSblWgCC02T2Yn
kkncfTeVFKJPs8tG6OVst4g6BAYu3kH10+O2guYjJcL/xzavziGsG+ZjvXExIlrX
2k36WSsEXqxUiZa9e8bBt0CheivibVW00opqom1CDFXpmQQ4DKrFBJyuBX1v3Vn7
AqjKWcMC2d54H5fyphJEvI/pPaHI+xKNrG0p7WMTefcVS3pt8DyR97e2Tkjapj4m
7vXkWRNT9O0NfZd43exbzqeGcUz+wwTN0m97sLSGPjo64zk2O/cJIVKyzFZkeODd
eWSUN17CY/s8oT+VRcF1Lernq6A92P+9EoGA2kIblbG65CyGBp0ecQ8rp3AdM0oE
ucMRNiC/AFRHMnd1MDc0tnFNBzzUQuGsOx1EmBNCR3Bz63bo3XpYJGpcq2mN2jrp
aRM+qqRTmZcpCI74tXuzmai2g4WZ2mKEItAVRumLglFzaG31MaPCYPrWZmgu9AIu
86VgNBOQdu5oU1pD+Qk36X+Fhg+LKaWEbWZPqy/SRHZ0MPElKoiSu+aj6/FYfbJD
V2a6hQAm2Knwe/NTY/laLTp/m0xOiogiFj3hyy4Ch8w5tOJ4AJPZCZlws3Te56ZQ
EN6SrE7tWuYTROl+LJ2hh9SZj+ShuOUV8uvR13ZSlu4lLbu2upvv4A8N6leI+kM6
bcCs0OLPw9LepeDwb9CyQmzM95vygH83j1kFTMZmdnTM2ipolChJmJu88Ncd7reP
aYblZp0XG09BbdPhkbASmY3tqijryXnsaeySquqoeNr4TyF//pGjHOEq6jHs9S3j
w/7z3UxjQT3XgThlsioX5+6KMsiUIvK9xQpRJomcaOeJ8vAPHYFsugIUc67+t/gf
MdEBzw9SuvIDkf7SIKR5kDdgMeGNf8TybKtWxEsLc2MHHn8+H8lCP7ERr3MlHGXI
YTC6hkc+UyWaWPE1GknMWFz+OGpYEeCUhP89PXDIir4WcIUbsLosusjVs42hgdgr
8HOFg0kpz2sFfyC7RLlRGTDPlRzsiZa2k842c+Hxfzrnt0TteEAFlJtH3F1r/vbz
BNnKZYcdvbX5yofYwuqIhHYRkymrAc7PPiajCQm6MB325YoZBmDOBREj+6yKvqyJ
48S2CqesPiPwRafY3nI1gJEEbpSMEzp9ZhRTUU5vuWD1L0gVP69uxZEJESMbxrcB
gcTwANhjclBUetq51VCVzAK7yFwHJZdLfepXno3RbvEbo6LLXsG9p3zPDzLmv0Bf
fV+52mJZkn8tAXYqqG3CHP8lg1NFS7aQ5tEE54amdxavHFGBnAD8Fv1FJDD+AIMk
lr+k3BJjs6d8ChV9Dxlan/wD6bAQLPCUBEVf9vmFrbEPC8Km4RoASzc6WHOLY0+m
utNlWafpK53Wi8nY7L7ClhCAOpoP0B97XNKz6u8IazP+4Bw2Y1JmbX8QeCNIFUHr
VlJGQXyhZCybhODnMegYYp2L46stX1hwjJg0XIRtn4VQQ2N8ZUlz3jwlE8rYwp3n
4ortz9I9/xZMHeOOzObliWTIKGKYdruEmL/7ej3AMgglq1xGMYl9HP/gHWRb/3KC
d8PbqBeMyQVE0JMfoGCOADMt8woxoLywRfln4AIzCmhbfFcnGaZfW6xXfMlp7NFZ
/XLZO0bkRSUwccwT3uOAwJz66BRXPf3ZFDHH5oqbWfH3su4AEUmG2QKeB6+SRFHG
0jPTUad/WauKdCt8IQI3CuhvLK4hbrRn9ekP5LHahhFxKMHrec9IMSaddlSl8HEr
M0edevKfdQuSBnIvpKXaveJ5fWSceZlQ4SzO/V03mVvfIpmzjSNMJ3iucoq5so4C
0e7i/VhkCsVVbxeziO3Xhckv0Sggy5pDxO0BmOvSdBa4/nH4O/gDGeaf7zqRxMWv
gImYVLUYV4eqthybKMZyT1CNQhpjzJIuOSIbtaf7y2SR9UY4l6WuTNQoOojFrt2N
114hwi6+pmGUZaBhwfCw06UKvbKqQwIbV4X7hrLPLNDl1JHJ5g+PPqJkr0jq7KTV
HykfCBQyv74q/83TFueLOHfpYBXsQYBgyUHZxrbS5LsJrxzcBuOPF1BO3tqlnjhb
6uwvtZnZ3m9rqyDnsd9oTO0Ckm/S/CQexkNCPDumSnS8pCXuLvojiJ1f1ocraIOm
EEsivgaZn8GLBz9q7wqYXZd2Xg5xTrlzf8eprjY+HG7hLJ5zN1iJGl9LDgwEjL2z
GGMrF+3p8Ndr7LjosAlUkR9pmA7IMcPD74b4FCii5/zYAgq1rroGfP2KIMxsyFhD
qfvHm1Til31HqnPkPj6vUu96+w2kMBhY82oTMFIckDnzzjtAq045Nm3s71ROEFEb
kalr6w8ANWZ2Gma2/09vofE0Q2R+z4hD+SVgzD9qLLyJqqZagF+98vtvpU32X+Zt
b77dcbndPed0XltpzP17RvhhVsNEuh+SzC8qH53LGfBaFnqX81FpNxJIga/BP38K
Os1tWorpYG67yXbYIPm/i6kav5x1f3wFsfUFxY8p15kZC7dwSjF/sSufOLCKkkvz
Cbr51JIKwkZS/p3Bt4pdVLRxvACgqdkNHkyutVoCceCo1BIS1FHskefr5vx2UMBp
uPC9EfxQk/zbduynbZN0RMS38L2+UBhC0Y7vA8Q0GebB1rOZ5nPfVQAk+/8Gg6ry
jsfRTcIcZr3TmsI1dX7yAM/1NjyGyS2xzHSfNJc6AMlKJc95yVBKUbssL+BbPt/9
ctJhXmsLjAk+Y707BNxh0KGq/X2g0OFFTyaHzaIPpql8W37xeZBP14l8Sq4CEfAq
sUovpTGy6Rsix6b0Haaliws5DtK0f6ORW4ZzR9CszIKGFsDrpiTwE7NEZZiIUqVQ
McuEcsPjBJWP3QFxC5DIxur3ZUvDb1MRFbbl31py+Xrh9M6vdsyw2FLIR+uwIsUh
Id/6Iq0PlyO+0NWanupS/itp0FLepBjA8YE+XeYXI326JoKTAiMwVB6Ag9ZtIKlv
mRw7Pp23Wpr2WqPGVw/q/AFWlMmf9A5nubiwmdBY8G0+QS8rL3p5cYQMlPUWiQMe
iQjITyr2D7Dk+wB1O2WqaId4qAbpsRZvnhiOKWuOTaLJgJBU1kucuAGP/QmF/Wa3
/8OykI1TFRRGBHmuEY/ucc5XW/wRD9VoYHpOhwdgEyFEON57LM031U4+kNLnt9Pj
lE/OYjW+SGZ06bsdU18tdLQCN0mKOlrmkZxr+YMp2vo768xzXJWaJYhhrPZuzR4I
/PTFziNYeUNGOUt9ZqCklZ26nYXfbmCgXcArZKCpV0qwlhuVNzyivol8n4OIcKL3
vqz2ehZPUPjOZbSl+Fr1znnocCDamcUah5E2Vyxz/SGvdVjrPWPPUGECr89gVHId
I+vhNd3hBkFrBrOhQAfANic4sjORQcBrxivsKk00nCKFAjUae6ZS8iYJprrFwkH0
Txfz2RYR8d20LSo4cV1vpF3p6PWc8bQNfz3qUWhixCgSo1EtUsaXRak4Wber2lDD
/MDmKfzVWAWPJMDmW/x15TioxfSnF54teVNmOMsJGe7M6DLhGFE0JfGKTqTq9zp1
ch2jrXerrj3gUXmEpiLy+wlA9XALsrYYpo7mt8SxM8PTWwtX0JpM/WVFu3sqXlVX
AXFdXaPDpW8hTTNMzspCISDz7sWidPD835ZNBaliJvLE5WFWMkokadHq9l+DAj3W
Yw+4KiIcmvgWHdCAuzVATSfQc9jCJsLksq3n+L2KXkfjr3AmbhfBF8kTW29V/0Hy
ju5pyfkOBFS9KwKAhnwu4/xvQOKGsCBW5UUPvsoThJvG4/lmG6LvccmS9IDD93lc
JC0kh5fosDteTepO5zl+XuYqYOYC/HMAQfoVXHA782A7rlNDEgT7+wB/XqrKAkBK
TENDgUw/Cj055jNEKb59XiKcANev7CI9s57Uq41P3O1U6fHsPq/NxdPhxspsewpQ
k4XJqlb3ayjmigzddXqRLe/xFd8BhatA9OM1c2AlemrNjWTCWxa+PjJfqdfRCvL7
KVns7BKvdpkis0/uEyfpxeTQ76O26ToS5jW1W8W6pSTTPhb9dW0AMZrrNF3VaF1T
fko/q7SOetmIc35ef4hkuBPBB+Fgh4adUZ9f3TXdue0H1y1qPnEAy16cdJTOeMSX
iRBydrlrdoGzzWYT/NeJF51VzaiUXMG6zLJ5kejGIT9GTqsVhKtY/7Cm49gQkQM8
Ib3wYDVICS3aTsfrxwQ8+6dhN6g+tD7rEiWi8X8AS78OQwDTP32IUyPrVluPoKuq
Rp+HjFNYpt756LgNaUr5Oo2DxSzceAF91VqUd4BQJRtxHP6CR5a6S544PInF80Xo
o+8EqazF4iSQ5hy/dr6Vs6ERDwro9Phy45YHkZhDYxLNsnI62aPcRfsn//Zy7Nbt
RbrB5N8kCYEGofOTFMKJT46TVDALki0uXDp2gaeCgGy+qnKhn3lbDjXmi3yBSHgL
rTuZd47rtf3qCdciiBLDp3WfzVCLzBHd7lWdXjXyx2sSmDYNCcr7r19E5KzRaeqM
NtP9kH+8KZJNfD17+/+zAVJqLiq6JY8mhffAWj/q2da8m2VCc54RntW8Q7LueDPx
FT61AJ8LB98RqRaRuW+S08ehHp1XPmRJDBMnJ3iH69nfv/Vacsr/JXZx7B4qqnug
N0s5X7WPPYYUJ8br2j0uteNBRVf5MgNeMuzfHbg1Qegw7UiKj13HGdsaDueEpeLI
plix0Csqp5FxlUwAxklDV6gvBQzn0Pkm6KKi7JjNhix69LuGybVEnacx5Q8J3qip
WtGO3bDtte7NTCqkiWcW+nOoq5NHx/Rt01+ImzvfS1s4Yd5loK+LcyJZBp5nfhTR
xLEVYvnyX5mWWRqDDi/A2NwgudUPQNCAGTwQpNvtsdfAqd6bg2d6qNOw3Q/Van3C
GiPItci4bLg4peh/wxzHWEHJq3IFvYLi6GifO8UedfsTwCcrg5MldSShuF5E1li4
N6GN2/jo5Q+riDDrELjtviutqlUT4YwPTlYtE8OF2eHsYwrTbipgCUnWPAdwEsqE
/hTwBkw6NjothxwH5S3On/UHTQGuFwIiODvINH9iBgbUrASK/a7t2OSmakqKILXC
jtosXkZDtD/Y4yG7oOuGzWQ4rKAGM3K34aH7jhy5QpwYd5dIieENMkS09Y5blQWW
fBFYEt706xEG+4y73MooNaFL6N8bQVUufuOAaCzGDGG7/AwyCYrucKhHrxws7czZ
F0gB4bb6OwvzbZKI7Kp1WwEgfy6pUGoqfU0xP/lmrVRN64JfTYGQ0efxJPL0ZSJQ
l2ODCRANLUX+8UIk2eEtZ/C7IFDUu1QJQxbwcBR9/ejwDC9dV6PK01VPvBiCi3BE
2jVy94aWGX8ipnjg/lSS0uyKaHOUoGqGhidu2FsQAuCqLFnrFRX1a2oc4JHHR7WX
z6lsKM45Zp/vuWg0eH9Ci5SGEK17kImcqVN2LKVLtVNd10qiZ8oS0oJzsa9vA4o1
IwPy4s9KJd5dQf0k0A/c+RpJcbaLAn3KXyMCLEHmNtbblE5lplCYyl7FY0fNfjbq
meuYKIo91SsUcYiHAVQPhCpBXj7wY/qeKN1J33LcqU+QA435+XKXz2hqXH3uvnac
IB7FQ3/BWxg/3BDbB8XSN1ysYZ3dyzfdgGPeJvQNsTi7qb8IeJLaq3H4EApiwU/r
SDzBYy8TYLvTDUY6Ip82Z4O5fb7IFXiER/2GT+OaUelVKSzR4B2KXtK5yL2JXWw7
K3R4sEIO2xKtgcrfA1SUxxmclKTLm5TpQp4940yBynt8Sn+iOCxoaSnQjD+bsiCx
0BO5AUERdyk/wZmtOEsTGFiNeCZ7zkU9vvs5uP12dClODFF+3FzCsftDO4McNi+Y
E0gkscyp0LuuaCYYruZNRQ7b23PRecgpHZKRO9mVLi5XcbPV6qwQdTeUY7Id0/b/
V36Dx4FlsY6FNQT9gpwkB2ir6JahDq8ht7zAgA59evaUN676rqVACEINA2XjypWq
0NZziTRDilRFNbbAq3WYNILfTCbQAGgRwNepOlwhCNzqvQxmHW75CrMMHVRoPV+n
0t8BGRr3Wl6MYU15d0HhN2NaQWB8XvqXAz4YAUblWBudAfp/yRiE4jxfC6GU6sv2
xnfznHRYTaZGi+VDPmb4Iw3G8ZlavB/qRfLuTmuYE/TTe6nyJSi0Zg0XRROJEDC4
rvECMhbm/h3UMoD7eDkX9auSggvcjqvcsVlGmNv9U+VUTXgJwcBIZo8Y2vS8FVhY
0onCMCMjffxte7EjckIdzBakePVwR82vJghlM3a061IXquWYnGj8BhKtjAIM9v/W
rwq4q/wQedwT7ybrqV8Kj9zcJgJ8/XC57I8eeSuAMUWf5uYs3wrh6Ir94J+AzcOH
+ddaYgqFjQLd1ahWhJK/9DF0q3ttkU6R5skdN53yjvobKAFtxVyp6X4t+T2t6R8m
hAZ5fiS7FFxbwTy7ogLznRSyIWhyLpleu0Cxya03dA8omMVkbDt9z5jorNVCL8jv
pH+lvrDLmkdzwmaGXTEd527pRlY0Y2gRbRWBF3VW8naoHP+MiuV+eEGcF1jj6mYO
o5/W9MSKpsk1m7AndNyvvkEOcExKVCLGLcf+/kGRAXkl//vha4/yG+Nj2+3bxjkA
peiOThHZd/JgygUbvlun+rVzgEFUcG34P9J28CHafWGMYoi0WbpMpb+NAC6keKD1
Yn7PztzRL1++75Dg2b1dE4qUI7th7LYyfBFdV//2/PSVyzTBf98C/NhnCXJDvzJs
aZBH/9HQjtf4d3ENQ8cV9t+h8S5heAgLbonvxiWL5lG7aBN8gakD/XdBNlmYi/EF
WYlP/A24WPLOAZH+ACBzZkKzayHnE1LNiZiH+IYkQpsXxaIRzlpjwO5TpOcK06ij
6CwbnGs8P5UoibdMKSosi8mUHsr6ZoFTOKlWA8hzV0T3TjsNqEbl5Wqavkt5On4H
1+0pc6llE/kDryC1SshC5wEHkpclwgKt+Sfsc1AyfKZhjppB7KvLqLhxXJuxEgbN
U0Qye6yBd++brSRCy+ve9+tZa2OHx9QlO0HAYPRGlpSeRckDfz8HhgxAoKp11ePe
Ax6+Rg1r6WF9KAnmL2FwfMACGVd67jFrQYBIV9VGfcOR/XU7lydqqOosxSzR5+eD
4AjCfV0khbrIz1SeAl56q0VKdDTKtBO9Wx2kCgnvltbavraHB5fLsVOvKTYOXXJH
wBFervCUsSWovs5lXYP0Yx1Hmh+tMtoMiqJtl4RO3zbalaRB9+TE1NEc79z14JV6
eQxUajJ3a+2INW+RXCIwRdPnY1kNx2+/kAY1O5y9GPewBaSDZZ2Djxz/KRtkA8YH
eG2mHDFKH/5InczQ+25cML4hhdPo++mFkOj0tBlye9sTFsmvHBbqy2zjbnMwhJ50
GHFk74GiedgabQu78sw1M46dtKo3zWpzu03hjZDuUmBxy0qEw2xowO0XMcrEmv94
y/R6x7j6xIUJukh4VExKjFflXT3w+deRH4KolbteiQNi0+CHtrzquZQ3m7UexCOA
CSPaMOLjgtmGpM7eCCSR5BkY5GeNUU2UkknGPZNvcRG6jQlmzYe3DuATgbC73HbG
9SvPYQh/bXKHPnWk2cG2o96T5PNjys4qCNojMIEY28vWqkQzjQwFgxzeRTcUQnNG
sVw6hhKikkeK9tko/BeLUIZar659Dt2/0gAtqORowMN7l8MHuhviItWazxzUqwZn
kW7WuM12VwZdgTOGNxD0eIrcQUfL05kSRCUqivSb/rPrKwq+z97FLwexuecCywyg
74nR3XF2X2cK52Eb+Jn4TO2xj6JpoZN2Sp4jKmhcSbIMhbuSGeamL5er0I/KweTf
/WH2nUOPtDaG8ywxw9q2cCcZ8Dlk/z7BQaaBL9oAABA1WjBLQngc3P6wdjsDCFjt
pPbVPcyFtVIMIlIMjsd5xRr2DaKKCqCgbCEfqNX2XBqLC/OFuZNthR4bwgr5P0xH
iK8ajmxAyCmly4vvEoZclnAUGHp2Z8x8KICy1aADk1vdAsoL95R/sgxpba8eYTQm
qWN7lDhk6fOCoZXSab2ansbM6+S/kSCtCZQh9UH60qogUIrd0epJzAU1ULQfjWXI
1fxY+uWBzcrSAPQGE85a4NW/VDLHiYHc+MHel713FVfXAWL4MUHzhHllfpYKWac/
hnOdz4ujEzIW52u/Hu/tVPBu5gpaoxPOdkhC+Ibtg4KPFymMzBMPgQlaB2JCfLkI
kUeUaExU0ieB6OJpfWkuRUByfjx0kLiM94lLETMZm2HpGakEjvdWadfg2T0zC6dT
FlkJ6Cudv4+7sdGB0jVTfLfR6LLeBEGfJAPf49lroswqUJ3n1z/KpfFj9y6GrgsV
m+2N28gZr6WxMugZ93q0u+cLZxb6suR8MuiCiWOPMiNVo8vT9FIjpX7IoslN2Zpx
OVANzCSKeN3yrmcJu101ldFzmTOlocHuuMgEUgFpZfejExPfg9Hn++JMn1Q+1HMb
Ipg43JfD821VcrOMUxoNJtexUvCPGV0QX2g9tLGEItnTURpOEml/kaI6WHqTY+RJ
dpXuL3ZXL6PHJuKakj++XSmPHbfzi1iR64WUsTqHpEiVt1+ZWVRxusGVKgCrf/Yk
7s0fWW1bMkDGmG+mxuOd/xjbtXkgPmHiHGepuRvlMWCLXnrVwje0cIt4RG3It8ku
JHzcf/DM93KbbvVAr55pnd5H+nFSjNoxoowIuLT56w1sCs61DR4NMrzcdY5iuvWM
43LmWRxm+2Q5n9gEcHCSVwWMtZyi351mdhCwL+72UF4+tD35A5cG0hH/PimcofRT
oLmcUX7aclvLoDnVLY1jHvVtYr6eDRZHIrnXAuh9t+BLfdUFHxIV326bho8BNSew
N8UsTZltdlnYLoKISTZUbm6K85jakb8ZzR676TYMcqa9xIXuRDvWTt95Q6P4VnG7
+06GfKBElj1iknr4Gd24bcKGEj9pcEKyJ5IbOiOwGDEYz53d8uD0VSbIXJrzX0bF
RakD3W9vCoHs3eI+MP45/zDxH3lwdB5bcviZ09jukIXsTRxsaRHjT/+BLi3BnVal
2nEK/z8u/wZ4gsc7JfjOjZkhfE9fH5W7XVc+GToHh3lqGqcLv9D+NkfMUFJjQRgN
8Np5mauJ5jjVFJ82H5MjCfoUmf0Sv84i7nba/WOfpGHwlhgNnSSIxyQ1P+HLhjcY
ONsLARgAoPXpI7EzmnAv0SE5t8NiWgqVgDTD4MRXrZGp4HVKK7fylb67aUbVS9m+
4cp5nk0eKYESkgoe5vqybJqZtTjN/iGJ7fzk0dTMnvgXB5OOTrBDr/0+aOuDbS0T
qBNQKFIWnJGWFkG2RHDywlyH803JtMuGMIEfaXHDRcyRoB4M4G+a70wHAPZdLu0p
D1s1sPDDYfvPOKMzIjNZEKEivWXgzLWF1bBLYEbF1Be0wIgq8KEaeQlBn+QABA00
Yoxg/gwyecSWMgaPSCOVYjqIe/GBThmu117m3A7UvGGX37osl1HdPPaJHciL3zr7
kAb8QC8A8MAZwIolEYDq3jX2Zu9WQFL91V8Q9scrPS59J8QqetJxd3+5qiZIGOx1
JidofeqoeqC42YR7r+U5CROQKWAhhKsxYAhjqOjeYbaON6Uq2mTA36VYbDRaGQ5U
rIHtptwnP0KB1u7jmiJjuBLSUQxXy+7sKqAyn+w2TjfWL7Izk/lEc5moMydAfiWq
43YZXhWbkEsaj/x6rZD4FQiIQxGrDBH0TxGVmhDtp5kn/lNt5xW7Fo9gq4Jk1+wI
/+yB1dAKrqT8vw9o2ryG7Gps0tohzh7hl6bOTz++NyqxygrZRyjoTqwTN2aqx91b
vP2WmxrZzc6YgCMYMQLbaEfcn8QzH6NZTLWmNkZhkeEJ1A+KSL/9aYTWlSOIyB+D
v42TukDM23j8VR0jyEfEV3aL43KBfO7pBx9TaoVQJDXrdlE5QU/p/YA4zR7FD9nV
pxAko4Ax7MvGCkwm1NZ3JPRtdiY+jznY8MPeGcWkCLUM4rGNyG5GbKQpullON/e7
ibiBcKNArlaz3D0Kjmq4tsQu9pGxCcTplrwIPZ1ezhUwQQmlqFxixsKiCGGDbmMi
ahMn+71sc0cKOB9ziDaSmLS6RtYSrvuHlm+b4hPyaqj0MZNNRZS2AKAZZwAlLrU5
7Nch0LiRG49GyKJFMx6NisqeGsGNMOdJA1a8CGt1r2Dk+4Os3jGXoIw+26sgVi0m
maenYLSBDscAeW04FXv147WEcvkJnkUGhq+GTEj6El3/jtcDw+CMSd32l2rk3agU
F739ZO0MZlrjyLcIvyJd+HdeW7WWJiK17FbLqc38dn0My5xpnjjzjxoWTAfk1Ioi
PSwTGvGZm61PG3LQg7BYeD26jaRozRh+mSz8lSrYMkHDdHJpWtNVTVpsFRC54v+l
qh8BuN9An/SxXn0xpto2j4HWz04CRAmQRV8oOyG/eT4lrxBP6pPVNV1DNje+VHy3
EPa+L2XdTdKYD4PCjRwX8Z04hKl97hQgZskZ65YmrI3gkno1rwC0QkHrezW0TMAc
EIUN9FF+9MqiBNJbT2EKF/kIFt/atKsapwfi63jQsnocTsi2V8/mtiiomnEYgMcP
CZ7Qpyt+a7N4JJ0omIkPHSemmJ2O/kxMgyT770grBpciFZTthWIPLjA8J8hCWH2W
6TmWtmZA5CrqgNysHAtxKnPXkr7rUovZmpp2bHaBJKya9ul0DjaMTl6vLttyU2V4
OBlcbP6bJ5N/W5wjgZ2ganzM53zalALeiR/6blOWZQUn7T01mxsOErl6g15iM4Uh
QDnGO3rxKJ1hJfWfjHvTZjH/s2Hh5mVsgVlsB4WZEUhBYObmAsNfO+6F6y9k+NTp
GhZYZOC4ZRePl7a28aVNQU5mbKdM972YNjKjzdZXycxp1ZpoEpsrIWjfMFYOq+NI
SDW/ibL/kdZ3rQlpXRec515koreLh1YO18o91LOXZ/4BB8RryIMNEUt9NdNrnib7
dEXXUWPisS14ZqY0nY7//P8+pOjOOi9j2G0QnTkpK5QiMKBn500obuqua2/v1Q5r
SQiAoMKGM5S3w8uajVgJ8A2Oskp/BIhNCvytzLz2tjfNj5657vSMVMhFhZNKvnic
NGTNX1lS6nbb5RxqiqTtWiQYPYifO8d91s6PmxIVuYNMmpKZ5fjrqPK6bVu6LKQb
ttbgKfLWkZ3WMNuhCiAG8k3owPxRhPsOulhrQCRtMyS9yA0hrNgQQ6mFnCY7MuoH
hoWfu05WhoKUMizxR72l+o8l4wenP32gQAPLu1YM5PZR37wSV5r8SaqeuDJBBamq
F+NN5kclqeFUmwb+4z6SrPZeMYsDqVb2HoEcG41c+MGE5bRcCvCHKH4WE5JBtTFQ
o05zpL2IsY/ccsQAQ+94923PI48IGIfif5kmbgq1IhoBuxiv2wGchWSC/YXHkY3D
2PM5VZbWs8FRIf/dyeS3WDhUi/9xwRyIYyFYK66vRQ6VS6DWXX4i/UM8CRErT0oC
OfsOfYui7KpgAz/UWYSaEONxa4HLnRJQ3RrbCB6eMQd3doIXasmT3ipQ76u7f9sm
fJleNrkTnht0QmS25Lv8GsH4/TxiUuEzSjXf+qHz7hiLOCGIKlQ5ZZZZiMccMh0W
ZgAaOv5JzhYH+nU1FzHobcEvbCtZKp7MMjILB9M9JX53KmsCUFlWwES5wiJFRsU/
TPBhVa+pzp0b2yOr5xwQ9viGsxzOBHZT7QvV/4iMs57WN46zDRFRyHCyEIthmzrn
WSUhZWW0sqG05hJpvaZtnUt7gI6Jcd/KtAT4AZK4i63BsSeLlzDVVqU6dkkw+pzk
dYmgRsR6i+WcBAm8lTNHka9FbawnWWh1ectk8a4uxnddhcdMna97rx2hanawO+C/
cWvRFmNoPDZdVlpRcG9Do+0hg5/SweOCeeh2BX3nTnAxM6hmMpomiN5eB1H3ReF/
161VcOag/bgPqstlW9U2WjUC9QLa504ZX23jaxDlullqlbjcELBiP/wODVuGCQ61
icTKcUIqQz9RRKkoJMuKotXRsEm6jSVUUY72Qnzn+Kv2vkzr5vEABW8WCVC9v5oa
UewZN0x/rXe1HggPwbnv4ZXScf3lBFTaFI0fymprg8zMzK/ik2kq2bYqZmep9xSh
mMYKk+9pd3ews0lSQPlH3J3TDzuPFANGzpiUeX/xQXiXFMxAWl2uo0ToHQ6wQ7Cq
t9Y4qbWtzCYujK4bhG676Ypu2uvNITZ6sSY1SP6cutljD30Tcbdl/8nkrkdO+xmu
HZX1AcQinv16ATAp57s26vldh3wKUOmuoLYYLo3KSB7fHt1ZSoNoj1CLKf6tTU9Y
aFj7/GvI0EiLhfrcEYYWP2O0MzQTJXUm59MUg7g7a0WEICKuhWOdVY+fxKD4viiV
SxNcUfIoNAgU/4LErGV6fGViR1CaNymwNTw6LTFExKliR+/6hfWuPO/nVL2ss3eX
FNXsp2EJJyp5E5GClK53puyQ6ZxhsbaVc4ohPHd/HS80g9ADeCrRm4+3p8kLm3e9
sCYaLx60Wn9ds8/GJ2MsuSSK2CbFlJLU1arHk2+XwSE4K/gfclk3JjMntlmVD4eB
FKgugF/Nm3DVqXhHf6CMrgkMmeHw7qHqMsLXvCjRy1pdwSdB6TJKljeHk11HBpHj
jyRb3AmzC1rPZSzNR2lYmBmDJ465bKrR6/1GT+KRjD5tq1htWGPbpDwLQXA58lHt
uO5RBNhltjXXYsdSCH/W9Lty9H4RHvTDTeBQXvtN3bUsuqdVTjZewsyIDcYbjPwX
PJSV/7lA/yPVHq9r5HTidkpQpTU83O7OXFBUtr7TpO4ppEB4eDEAh6iolyhBUZAm
PcgLtm3FTV0FAiWAYjyeK2G8jKFVrbXNkzRHz2HAJp3h8i01XG9adXWVWgLw3621
gl59sJBBIQ+EUhBOcuCSlm80r/zvUWJZWidQp/J+EpBW7wxNL/tUT1heGhWzEnCx
MuhIZa/mngRDy2O/pkqAxRgfHmfvvf9+bmvLKFRkM+T829GUN+pAuc44hSUn/WST
zTp0Rzvlv+2wf24w6pZJ5lzk/0rj4vGl3b2KAbDhehTVXvZzwe+1MjyN1kfIdBzS
S8SAuvJkJaus6PWMOqlEZQIxlYgdQENi/Lm2JKjJwG1yvWhxk12dYaRqRqfZsvfG
4ZyNjx9GRNT5ULR6NwZidh6v3U4C/q+xHDIGt6mnoQph+5EgMHOnvNNuS0uTHI4j
obaVggGX8y9LUDe1PVtWParlGpwxxDTLoGqvPicZ/UHpbYsj2StbcrDuxlsiMCE+
VOpwZ1+z9nvKklN5t9EUhAe8947PLcLTj/kpdT4P/HfKLvTbiEzcMwS35gq2XcxW
PpfCh7HLDQgtgHfoXxM51poDpqcDgD9ZoralQT3359noYbnp4f1d9tc2UdaBum0F
vAK5FNJ2QcR9YLh0WjbKwEL+4oqhb99sF42wnbulCh64ecSbApW62YNR4MvI1d2w
OvT7zAjLcIoFHnl2185EocwNSLEMvxVH2jjKqA31KzZS7vcS4uHHuqrCFIaCTDAd
dgxel1u3vU9hl2PzN/1IEjoNbGs/JUMxIUsnVBuSnXXxOBao8Pm2MLeCvNLrnTGb
TdCex9X+3cuhB76EQY+oeY8lTYykXDmB1vz/dX+XDe3u3qoxPfmJ4g/CFTqrbWld
EVu7gMovYiTGyjsRKA6o9MJSLuc4yRomB45qyZ6RC2tMPiwkma1ExvV1gz3zcep5
4WJVwXCPILnIxQIBnXjMZDpD7NNyvQ5kyQ/ar5yTfGddFr+SE3ltaIrxHt/nWIne
JNb+zZpYus+wwvJvbCSDvIqtE5Ii1rVcHPnP9oBNSZWbv4f+lZ9FYgXHfs3csxGA
40CiJnF5Whnf3vzzePlM0OMzBA/Sr0Yri5I/Eb3yUpM85hndeJfkYeUy+U0lC779
nLIe5pTpXZrDDijCvIJNbDd/T/Q3WfOri3/1v8FbSDZsJCNg54epDYaNBWESNGOe
ZxHRDQ9WbLMSu80h9qMuBXIcFH32GuNkzQ9HFk9kdvo5YDBRQeiyX1SVW2al4eRL
Eg9Z7YTCoqUHUpJNkava5rUdd3GpcR5qUUfbA36NUJjdTySBA/kppEdlcHIOHEp7
t5BgbBI/DVAHIFXYiTuHkG627VDGUjELUp245TFFAS0z2Vw6wNFCVx6sBoZXRIDD
IpPZZgMrhQEdQw7GdnOoP44DCKiL1tExhdzwLOuBdV3dWy20wzU7Wk2ONjMYjjIU
5q4uddo3zLzsCFvuTfQaB/dAPVcJiSXdphQLo2XsQasV3DJjKcs36DK5iDSTC7dR
NR3Ip97K0EWFA6keouE/6ljhEDA8TEAE7VTjmnNBG9GzMzJmh3nfXY/DWtXImXsv
Y+h17GYeWVmUxJ9txfPvl49vJYD8mLWDq8T1wVdInlcy7klVRzuoayr6N6ga8Lkn
6EaYRoCcHS2dO/FTmx288I7JU1uJrkIozJah7xTjFD7dU8jlCa7ZbLzt0P/qKXV7
SM0sKKbDm7kAbbsMyb1EOt5ACfonkGdeT8AhBLHmhCO8+GUuOMWQ1rqA5t9UR5s5
+4gnqPeoh8BigALKuiX9BODrotv/+8UozTiUugkoK78c/fhj9vz/CM6DvKLZfMG1
BxTnpf7WZjU3DE4FahXNjEwlgpFGNlGRJ4ur6OPqeilgA6OeVX82bxe46tzJdg6r
/argPPtqH5JW2zd+ZBjw4DdE9QQSY7vBm/m9uu7VEu47vAX6BH59iDcWSKHURZq8
ppSbPxlkbbXxCxHz4S7X0miZH7sNHsv369iIVr/3y4XDgoKkvcRFZysW2nsdEQKS
dkFZ16QAvGbvUUv1V0UzkWgsrXezpfkhsMsXYK6zx1Zv5q7e0JgM7ll8dANygOS7
aEC2ixRsAp07a2CsixdfruxTeYeot2jHgLDHqOFaLhlOAZLsFUnvUmlU+dXON8P/
ZVrux2mH5+XUdrE76I2IACvPiPU1QIi/cCyfbypSiA66Du2kekvYEb+7V+j0woOJ
vC3tBWH4jslVTAwWqisRyqJfjzromACocaRNBsy9kC7SkcR2hHn/5PzItHmiCysu
YuXFqse5jpuhLZvUCnUuVGfLOPzVCN3sydnCj2szDByuMyLRLv3c5a+teIAA7oZU
D9Pq6htZ7yzqAs3mtKsFWk6i7x0BtVabMKRP5xdR7O6tnJIGfKfxq0a64ojOf/jp
rwasrii71NAyeQ3hAfOPcJUoCKKK7ksPlO+/58GhVQnzB+gAg96wzBNsNpfzLodu
9BmdCckfroFlFVfA58byIl8rsgIiTjZSE7HPrSOa9LWjgWbm7sa1kS/W8ZzeUWqf
pJyhlVvte3MSm38Xscrw2TnGRTZB2rfPWTcQBtn1tuhq0m/mkmLG476n8J+3wo3j
zHsGSv1MNCBBUAZ+vND8mEfdeotmxbmiwWKC5b2UEwXusWBHSW7kUQhnxEGHpgGd
VwSUCyBz+lrjfB+D+lWkSTeInteU1gnQzS2bv+oCZGGWpxRFzmvOyxeNHARR5ALa
tWWqac30mrnOurHJ96Rc7I+RN5kipMDNAtAl7IZjngZE0Jeb8Ti3+S6+Y6PL9wHa
A23/HPwuZ4WoautmFmlMkM4CVzCSfAo4/p5MeERnDmbnsmkCzUDJl/ewpf5x7HAT
xmoNxcsQhC0SxSW//JWlHKj5P/AirUd7TOCj9YD5oLTz4tR78fQojXqVUEflWeJI
GZEI7OQdWFD04yxftzdt/HJWmq+BvegBrjMbXPPVE6j7kUGJH/RFHekA9wOkhAq1
mTXB37rZljWqZTK0WuEl5/oBP7Z8/b5d62DT5rb7QDuPJODw+dtlT+lXmkXdzWhE
1q9lfqUKaPAmIMOuPqgQvCx/SNnZXdL9GBjaSAi7u4sdG9QXKo5bpVBquv/s7fEs
jnruHZJre6eI6p1xlRCCpnvFRIkcPrWJUvPV1ppTstSfqgnfXuN5j7lZ3+gYJ7de
bGOSTVNwkjZWR4EsWTP5VWWbWfR4k5ic/rgXye88g394eatelmiv7AbUJ26DQqKr
2WhxkRaKoYJu9MbheFMcsUOt8F4hql+DP5pwDuAQFmmRkaJiVR7c3zOpXGA8nnaq
wLCGg36KXMy1qv9FDWDyboxWlDOhoXmAxMTbmKe6X8uty1uH2Ii8zFbueLV20VP3
QA7cYVQ0UkdpqbKpEB49CFf5nQhqupOU+jVpLM8WotKHa5yWfThVZgcGqzzvzwmI
FmdArku7jOhfpJVYnbbYVkKbtNTOhsXb28srpmvOwfwAlzrLzFxlamjaPHlJloy4
KAI12jEaAFx4DQYCDw2pzsCQSFk+tbkb20crdz3voriSnb/ZnTvDIgJ+yxTTDs6P
aFAutrDrDF4ysh0zhCTrbzTP0WveXAkZx5kRhjQLdFXTsmLNxZK6ZeaoBdr/nKft
g1NkykMmUjE0Gz/9N0+YLjVsgaG95TnWQtIBf1j1U9VvxRhL0ypC2sPGlt3+Eu9L
Q86C5ASXs7O3NNUWsIrl7sRFJVka2DlCSQ3NqkgujuOn0eK55q+zESVnbpzuI8+v
BUe99qOdAB/RBdOW1FI787O26HeJTXZht3noYKQmFou9O8sXQ/dOxBzfbWBHHeUV
gtLqw9YF0S9HhC0W41Es5n7zaReaUnjU0Yj2ndGEEWu/I+P/tAt1bI2DyviaWAHK
QiSvcf4CfMItAJ8Stn+gE22LZuHws0ncHJrCzARerAtQ/cgGkBlxQKaDzkghji6m
3M7boKEBqozbAjWqmLxm2rqjWfHW8/rM5uHcZiBrW9L5nrUhHcqjqVZAFIqKQTaM
pTd9jt67CooGD3M4p4P1xwaiT04mDBIi7xfWBGvQpbzXCCFtE4bPeoM2ud2S/RSx
eGZDQy55y5Rqabt6mJvB8BN6hpvN3mVKvbrUR9NyjGOVrtWSTYIVmxZcyVGDat7a
ytHBg0D03jYuO0B6EtxcfUJbc49s0bXPzvVqBQwofnCVQQanyxFF+3+clqQuHTft
FfJ+LEzpqEJ8/9PMxCnGRd+qH+/5vBZ6jIKxCHoOSZAXr6fLGT+VpFPz/SpzSugc
yipT5O09rPCXB4vIDWihbj5FanSO9QiO7jkqeMC/VS9ZAPkj+c3rXnNe8x0EOS4V
CfBjAZI+VC5kbnhU1+O8KD+gVHiW53wpCh/5SZeLp1O3Ew/qrUzfNzKSjy5VSIqQ
OPjYRy/y3FOEEA9LcctmcdWRwJS1l87cx336PmYiqOd+GcuP3ZoYUCkYkBszgwde
pGsIbhAGZObz2irwkjU03ZkjUe7I2TI95VOkErdJqanTJpKiVIWKDsdHQlr+IWEH
cXxsczZxTbo4A2FO6yLS06XMfAGttYYtPGpC17B61jXUnwYi3U3RJPa+q86hTgcP
Sn9FcWJhv1PnniF6tf64MGqT3IHH6FisqePfI7+wcaUqjMfqRGj9lZlbHfWPsvGr
hDMXcUtzpwHkpul/7LhkArsLK/z9iynMJwQJP/CWjUtZAzXFCjLMDF9dPZ08RdF8
2t62pyaF0Fo1J+pcQQ48rmWOoMBuDFX2NH+OigznonEhk7edkGRCY0t60WERfCji
UWIe1xEGwe/rJchxrDbBHSPF9KVDhnoWn3gsyL9f8f3LJF5wnzs8Sh5n1gJyR5hZ
49k6r7OUe4hl5deKHBLYHKMm772YWpqZMFXbyIQvJ2OYEwVJ1w8MeAVmrTkBpf8+
TjlJXNgjWlf0XXv3BOCWibLu6w2Ykajo6r62sY3v24QYBKdItRahaqueB9dgW6k5
VB/MXGiJopYSJSpnUMMciUX9VhdlufL2ui6QfmOzG/2eZffOYbrycZFvOuxHUvqC
89Ys8UjjnmoVdn7+0sCKS3dKEPEzN4QOVDOLPj9OSuX0fUEOkLDmT8i6CqwwEyeG
deEdpahzRafngrKLuDPQJxJ7ETjsOR2ZpRxNm+ebqy4WoGr4hxVp6XUIzYzYVs/h
+rcNUivY3/JHol3FZ7nNHuYarf8fFUt0b2lbeLLjbC421ltRyKRZJkdl88pMqBaX
uQNmEOLVRkBmDh+JAbRJDzwt7dHwGbCZsg8/BBGIXETPy7j0eOzFKQ7x6anzNweL
OlfJ1mwcnjcGrXkDwqH/bXTJ4Fyw4n4lGFDMfLPokg6su7zK1PHGQ5R16E26k2ww
//bIhh122q3Djq8yf71wmUTdRp8VfTDUe0t+FPjB4G2SD/24Jdm7kReIqnYL2x6K
20U+ljK011ev1hiby0Gi8e5LtdxKECE1f6kgeSthM/8JsoirlUg7WfoMv/CQpcym
dOQYmSXS79Vy4UrOkq8HO16M/qzzaoYF0Bj/9SYAPmArPcTLIVj4+T1TZrDfBF/D
7JTrLFmpyxZdA8aJYr4P/bpaZhrCDgSb67YdB1DqxCxBYrQSCX5S1ShQhwglh46K
ScoDQVwzobX8cUX1Yg4BhfsGb6TmxKyByqjPHZmR4BK98QroTPWfHVSMo/zo9KAD
c/ZG5YL26DsWneF7qwvA3kNE2A0uAohpZKyKJr7eUtr9iNTPHJijdRQaM7PfrenM
8+48Xg3Q+xDcijKSBoRKlJfiT27L2eAaHru6/1k2PUq12nV3iAC71a4Eg1Ftoe1j
vkmOOeHtUa7Klwdzeuu/amYYvmdDo9aBmiUGcd9mmEiHg1H3Q3vGzbiYYt/dPaGt
wGUyonNenLdYG1pzQr0Oyv6ZpUX8OcIjWmDeyWfrYKFSoxe+I/bfxGu8x0dZYq78
jvqgTZeVUQrS+YXQxKW6fWnwtaLQQUM4yen2I/WZT4Q01iZoHlYPFJ0UvmNuz0uj
rEXfZ5SP/62ooa73Edlj0E/dA+v1SNLN7PIJtWMELhXzNDtO6iFLF7sdzEsb2+T8
sX7/50G87Hys7/C4/zv4sjsVO9w+TrsgpHKkqeXS/2crn4ymOsncay0sVDbrukbv
oGxGz2FpzzKKmp1aU8UMhKNTToUh8GUKzkNO00k1ps8BZwm7Uuio9sikQzIRgmpq
347xE/rslDQC2rWyIIb9P5RFsmxxJNPXSOTxWMoXQm/yVwUF1zMHF+Ak56HtGT9I
6z53dnjYaYVT+1Dm+ZSsJRJGJJnDwmnB+UDjxkMlrja9JZe0WsZy1tApgDLP1/tX
TAgVxA+LbVI6eRNomoNuDcLhTmhxWc/aMSmZuKni954Lt1G2bDaAxy4Fwqj0VR5L
/cDbk5jll5ME17iJBHyOw4FmuxKELeyOLr3cfErRXnQe8F27ahaxMTWru5QUw+GO
/OWsxYJ84SaFaUwiboy9IIB80UzUNa1JSDIq0grjI4madlxkbgwOfHhBYtdzkZMP
JKvHoAms8W6XH9PWWpL2hyusOGm9wKNQRfFCq1/gK/CjGrwfvoUBKZPtY9p6gEWO
suwnwrxui91f+9apy8XjHMVv7/IU3iQ8yLH3DUNsgkLm+hSkTUgozlk8PTLnTPEJ
jNmRZKhufPC4wZEvCHpxxnB10ES3CUJ5qFsoj8LHFH+IYhYZNol6dEV/OsuxWznI
7j3+aqSKPPm/DY82Zfdjck055nXzX526JJIzFchksWPzF2K4AkJ7lxDsiP85PORC
EwePHEIn50u9rwmW64SODckQx7WPVwsanPc4M8ve0F+CyM04/CLBCFAFj2zMtthJ
AUKgtOH/oXQ9Q5sJHJDclKiYY3+8EiDdOliDJQnVe2xamn6HWDcT/KNoROnP4uNM
SYqDpaPTVirJexoBHDXZCZep613PR+LPLdoyNENCYLqTqj2sjyGb3hpFF77MNzhP
d7JRY7GKdOTcsOUUcYTu9/sRzED04JkEBEBZI8Nhe+0m7oxYLFUz3djLRoM29xoq
lcZEh88Xwaujz1ofyxJMH+g0nqrpFX3Dg33yp5F5GAuhYP0VJuCgF/xukRSNN/x5
dhfsrbAVjtTy7s7iuuyDzNQ57loa/zYRZhqPB0QqSS2QkHh80YS/ChPvGc5nxmXu
e3sFLaCO0MpJLWD1Nz/0DPlS1OoTdtMVCD9CYoxSGcZdz6nx6IT6g9bdGC+/Tcgf
QP7C/RiA5j+ReIslc5F+XvaQdYLOpdMBSDIGXyezKOqR+MkJyGTv/gw3HMD+fLDD
nV8QQQooYK4zc5zKiKNR5X69jXc6SuGHee8CdqSZhSBR/rl9fgQo5jlX/8HIaeiQ
k5j/g/d7k54qfvgfB5tNWbd2CTH3lYHaUrcijQoSr/ZhT0JgXBLScNa2f7uqCYJM
F03cpdpl6iFvaHmDvVGusV5kZ+tbsfC4DVbQoYG3iNu7aKl+kf5uJLFhmuNy9OQ9
FvsDAK947QX/c9vr8M+x+b5MVvIAIfVKu2+zcxnP1ahFyWz/aY0MgOjhyxCEVSG1
olAy/DiksqlwVhYN+VtdiA/FQBo/ZLbT9aiTTwqRjylZJrq4pkUfojGG3CjJDHj6
I1YCO87+UKiziqG8cg0lsrgVLJGmsNYM+ERtIYxHVTMk88yFukXJ+t02EgjjCW8Z
jqeyN6W/dddRB/Xf5S9aHXJAJO7iVz6d+UdodNT8Kh3Oc0nBNG1KKuDMjMb9AHeU
wdStJxDPD85f9eYNimZ330szWZbafcAzwoIEglt6ryEwo5+jVS0zJgjnamlLo1cz
H9ZlK4HLF+mVHMbphxMEfS5zWdDuDZSWadbvbJ98pfuewdcLblMwPKIXP2va/heD
OJwOVBDbPy73P314GOtZUKxfYCpXnVlq+xQPXO/6yeNR9vq6tgE2+DafzModaJOo
h2eo0s0GAlxp+VsSjIREVjiFT8Q9lkjnPo1X1PZPuhmjnj6WK3XazxBWjAtn/S9D
H+2qflGWZutPqVIriVzQzLuUUe8ZNJzRdnJCClrXxl8+4/18/c2sSqiZhRt+sg9k
xOO2019PRSpc0Mnc3Z+NNkrmyHO46zsefnrIq+tLMMFRxcsIoo+PHWT+UQ3W/4s8
g4+uGJj4KRxEQQ43iwXmfWvVAXCVeqXywUSZVEx+KP9E14pgBdin75qWVOSzgQTJ
baw42DvqeMYteGbUKM1TXMgtB7QPZLzK0hhWqGa2EFYMDccLQpmJpeUK/t1Ko9o2
1PoyQJiRuus8x+Oaak0A2RwQC8uWZUyOJeU4aMrXsuJL0gKOMb6t33AA9RCHGYpU
I04aC+h+IVCVNkSVtYmGYsuiOkZrLTWMsuN/YrIYcPGG76H+s9dqJaDUEcyERjo1
dQq01qhjKSSUb5QtJE/TkN2hKlryXZQe14RV35ggbNvh7MVBn55DRkfAYlihM1pm
08W/gSuwWkY0saa55czI7nNzm3t4680REzrrwVtIWKf4V171by5eNfhwqBTIKbxL
G9pUUurC7V5766B6u71lkOLRTR9n3xzYlfF/68tMvKl3v1yCTuSqGil0GIJ3daW7
Fm+KVsk31mWCnmjbuyRQK88lG/6D+ahPyUbgvKCEZ4JEE3DTHXOVoyTdXCP/Cfw+
Ci0PwDogl2CMkRWBGUGefwSHv7YQz/OhI+eCCcTfgkiS5gULVaxB+Jym/Ld3leDR
davkG5WbuybTN/q7uo+gk2MLrxJXOQuu01J3SAziv7+I+SRO16UPH1pUneDREgXq
3098dvq1CVYJKKGI9OjztdX1ZP40IevB0xF2ZaVth6pXvp/32y5+j7x/iNPL+1ex
tXoEcxf34RgBYwA0Nup0qmvOSJV5cD6S3dq/SjzGS7EZz5YWtwmzKeZpBxrMEiv/
D/VajO8PT7ePGACKy+lSLduIM1ERaobFrcSfLNOjxfmx/RB2WQPXxIrC++vN51h8
ysOl7HF+EKzkvwgus7KLbIJdx5G78CuNHO6MUJPjkKIPIGkTH+x9BdW43y/VNLGl
cAlze0/x7ox+3eQX0qsK0oBB9So0/jb3yPv9Mo+i4ey8LyXanVHdiXMh6CKK5ek/
wIfqqal14ePpjuQIeNUIDLtLkCbQNY7bi+wXzO5DjRiRMjtJFOhlc2Uz3g12RlgI
PF/O3eSeM4yPCRtLDbj0HxDaZ5q3d2KeC7NhPEVbekA4htpJBgETrzyyN3E7BQa+
IuqQEFcF7wxe5UC0E4jakB1vm8MDE+wLTrbIek/wu7oy9DdmTqOZxj3KnA+ZGS/M
ImYoEt9HJEmewihS0rmhbWlvdDJl0iT7TYRdt7TIxCxkfjIbwRTwIkv9toPBD4/q
K+EsQWGUfUaDlsg3FQCjQalusO81nKqgsgmi17KV6h/fzB/LrttUGWTroRWvcQfQ
dsNN9qO7GyPOgK3HMcBMQdbvtXEqgBxb4iq80fJoKcJWXhbW2bJsxMYO4QWD5hLh
h7MivxsCtNy6dRQ0Zi3eNQl5ski1vTo3oMRXYdIaKDXToAhhfR59AaRJ6XFSlIWD
nWyCo82whd39d741oWm/3o4wkAclcvywJLovDrkIwhdxInHJJo13/HEcPn4dvAVf
+44pPi1YYUeRe2qgOQlqGYArLRzMTuclS/msyxgDe9GQsCaEBnOO68pZm2/zFuzs
r9tiV2HLC8S0kQR/5WvadaUxrpMi/bf6BNy2QLD6spBCKHeIH9T3JANXfvUJvbQL
dWh+x1/VyzfAI+jtfismhWRnlz2QAAkXxi7xvX6xTTOF9FmuxDBXMZq1ntWCMdov
rkDlhKllMbcKZ3TckMmUOMG39qBh0nx6DOTwbyFbT62pWjVvv2zU0syqbNkFR3cl
nKDRHIcG87drA8ni8ieOnTB/p2Pv7bdH2agCxX8zilJjxC2B61pLnD2uJFOBeoiP
wKDs6WaNLPgNQOhwCoi9nFWU/IkVR3UHN5MzgPc4s3yskYoJIkbR9egUHRRebSGM
4CEFOSLcANLoEaZxGBHZXN7QTurWK58jzl4/UnLuWZqGtuiAKPY3VMeSyeoTmuDb
C2Rf5aq+I2+JBTRneYS5VG4xRq6EO11wCVY5bUE40o4VdxTtiRRy0AbkAukIaPrH
59g9ecdtgflc3Dr6XlzW9CusLBHkzDcrmo+jE/IojEkxU9L6UCjg/ymLIz1wl3hd
KHjH1g21fM9RNXWnEhpDsmeSWQHy49cKIrOU0k3j+Eq8y83waO6N/Sj3YVXMsmWv
Vj7jUy9gEyxPy5Dn098yjZIXkY0X+kR4b+nh3BuUkmtGtxN4BKXnSBFQSu1S4ab7
z/lj7D0pVbYHtLrkEKGdewhnSzup6GoVNi/17ty7JG6v9TErUtMZ/2jpEr5flNFF
+DQO2U33+BPJu16UKr5sYrBCKnrpDxGeMU9TSVb3nfZECJCXVPjtNyKGvQuCtUH8
7xU9kn6iBBaJFMPghSBxsFwW9AlySME1upMuICTX9fVKKiv+EH7/vIYXWtmbFDQJ
TcLPZJIvIyP1LSJCAmOSdyVjs/gio/7uQwP7YXyO9FDu2qZeUTDpPzEFWgPlix1M
qyDxUuAjYWTMBoxBoGhGlcbHxFexYEoN07Y4NMbtgjUQPOZgJ2+P/wTWikxN0o8i
GE1Lkwq7Yn2ngh00X7XiewuYQp7UqxjRwyjPvR5B/9JBXlyWWMAmieYK7QfQk2eD
EWApu4Pj4LTGoV/Uwjt0AhdXox88y7P0qrD2X7myZLKwHb3enQAX62nP6HWzopE7
H5I8pSSPBNNcpbRpQmrod5Ol7WPVEkKr7QlnKONsP88lKN6/tThs/Mr3DNuq/ukB
hMQoCTy7awPfjD9eAlUL4ygE2aGjW6BWpHQtDHv5tQ7aEUifWt81zxvA0Y2i7kCm
IL9l66cOaEcbIUqZbV8C6/0yXzDvDJLToZg/UNkPPKMkcaDVoO2Z1REn2N2L/Zg5
H0JqBP/zrT8FytfUUsx5SfG2UeOFmi5tiBpCXJXxanQ49R0xClAZyY0bPbQ3AgAq
IDSR+9ERxRZG2NOYTlXrEO61LRVeLNSs92GxP5Uf7TlsGPbtCnSoWZP1HipJ77o2
cXWWlP5mFEapA/U+uqHhqWvUNUEsbxtT/qyXRcMXs6Ff1/3SvWgQCRq/PB8t6LJj
FephYsV8yRutCkFjr/34k47eIA5CK8IgyfTHIrOspMo5G0RDAdUwDC6ZihjRZO06
QQvwJXXVRaZ4Oi65ph7a5dLdzlqEAEk0Qjmv+SgHlRcXZeTIJkO4hRHN17Efx65W
asU/QI5MYXL0YXOTUOmv5EOknPlzaCc8OHcdmqMREByKy+GJoX5CPucj186GMFk3
0vtiSIxp71j/5df5pMbOfqRHLgLVAaVywRKX9DmZ1nHV5i/TocedeUdEDOdiq1v7
IR2X/ARdH6UQxDhhuXLDhBTNCjj5uZZKt6IpKMbxb7FAj1s5Mq2tFfTPIP6tEu/a
hFuSsDEyhz+YLRnFtZ484aXskpVwybQnAaVWLvqToGt/wUC5q40YgTRqhHDKgwW3
JbFvVvBMEOP29crwPmkob6ad8eTkbpGm3XoVJJVWfDSU47RyIaN0X8GYxTkAWPlP
hLHCGxj1NPgqxHGq6n6E46J3u2bvcZxcQT5osqxE/Q4xWVCb6WNNOSAwH1tOxMqS
ps15k5lqIzuVaB37prMZvqkWKADB/2jr4w/g1iXq/l5aTIQJ8jqAVP6JiDl5YbzE
IoNX2d+XOTm1rtSoC2nPlHP1qO+lgJJGpIXZTHQUKKXoZluhibx/QK6pBBr42pRh
gR7x8wse86HdRzdSDONr1KZ6lQ5c6YHk0hP/EE8PMEzbD3wGpPjXxcaEZ7JXMTIN
9fl0kWAiL6EOe+yOVNorc2/tr+hAwe7T+qRqbHVpaArFs/AhdBPvTu9tzeatdTjq
2k42u+MKusz2pKktuLJg/zR7d4VeZFGfKLeTUqaBfcoESAUFX635KmvJY1G+XGWr
Y7nL9/ut7Fzix9hHMVHndnHsD2LdRaMQmaATeMbACLwts2pidbz8zhhhipbNLst3
ItzfBP8jlWamO76QTPDPbpAnF4OMIxlmSN90mFd3yU+hSp0MrepLEkfO8PlfT2QL
h7hbSkp6j5qFxwnZR9lv7ihvRcTAEOrfED4VXv8ZEHQBCuYKIbkrYjQFBBGZLxro
4q+B3Wcvn/KHmThhDpeWmJOh95qoVQMixIp46ioLmYqdhqUdjw6814WtbLe0x0s7
gcH3WO0v63vM7EZ0yWvXHBr9m4j/5vncIYSYdaR1+4AaBSJRBW4JaN+l+HSyOzQ+
4k4o4RG184292ojATT7H6wj4MAPbVhDehU2Cvx4XFDsZC6yIdEOf2kFXNHmSy9B2
S0J1PQgiCmgiEAN3dh+KRA3P//Nez4p+5MoTlZZA+gQgcR7FNNprRDyRXM+IPilu
yQ2aoYfe35Z3Vpihyd1U0mwKJPFAJPFDLSUUQBAZoFxeGZUwf9+MvnN9GBQ/l3YP
/96Zvok6YVOLx1LGucntu2YkrwVtE7+z8kHx7krh6YwvT7FEYOt/NhP0kmA4AcYN
f4STAcB8XzjCtNrdGuoaT8t84myecx/iipF8BKFPjUX/jsrP9Z6KdvCABI8t6dRQ
Rh8GMtR0eZdpBWCSJ1PQLJyhT80zJ4dS8tFuipWMnh9oo4EhXb02I1re1Bv8Y4t4
A5Lqn9AJUzHc0v+RQNwWe55nf3fHTwXJ0KJxQCUlPzogeQJVCjaEweBKjItPsXMC
39n+6ZDram6+SQT0CABGk10b2IttyK/la52468kzgqsM2CYjee4w7KCWp/mEwNzf
ypw3Y7xfTRy1gTubrJdPUiTNd0xufdjOPbyMz4jgVbKaCcxoyyMt4HpDs7F6xgse
rY67sy4mps243qvp7bfXEVi54QC2jWsl+6J4cNWScR4XUVaKjkr5McaLpdJo0vEb
dmmlqcQTtvH7dHiyRNBMMEbhSkKfnhF2DxJrMIBczyDZyuGYlXTpOJvfMUuRf4CH
qF3GnZPYoVMIkdVDJQU4WDnXxqXkcaA9IzXm/l+zm3fv6H4QvbvbQCp950g0oNH/
CdJfkYtwil+Q37Kqx5LPa4UZj54FTugRfbwIFp1cP2PXh3xPzPe3zOtNU/CHQXIO
kPemlAPdaUYhYJavcKiNNh7ErZsBP+JjndRKLjPklL/U0WUZY9dX3ecIAbLRTW5O
l/rUCgefoVEvFn2+tB/xrhstQqLV/Vjc9CdCBKGQ8W13ZwB2uKX/aXWtwuFiUlxa
O/IjtoahaV3zrX8tQOamCVW78c/3K8oThmsXKDtmUILoOXJU+1opRHm/jF79ax3D
t64wMWARrQOs6W+v027iTD8hl0D0rnJslmHq2Tq7+gMI/zknLGQ+zgUeg0WtrdZl
S33Q0Vy2sYuDL9mg+qU6kmubOK5PvpDDjhs2nBlBAfSDkWSDwbZPWpI/NbmF1xb7
J0cHRtqnC8r7Hc8yL87sfrJ/GUfbo+x8AyThVi6eyRcVcceMpRfHt3oH/AiRuYpI
oP4bqR/4Cx27Zf7JGB72IxnK/8KwbsphCSUcbkPE5h9js2oR/PbU0Icj5C2ajiwh
FLCQqlR+tpVYRgVu81BHF+r4R+55UjsXPLKJ5Wq7UA4Snnr/E0g8e8e2Hf2IwATN
97VHwFzn5eXjIzIwJ5R0NQ3457gm/4wTBexe89y4NqyWRMRI/32SSqXs0KOd9Iul
wKcDgyoT5UddQUak1GMn0EBHBGO/6B0KTqj7gc6YWpfrB4cr3IQK/0EbTQc2iFzg
hFPO78sKraNghAKMxuba7a6cM2svGH8VvURa4MwhpfhzFeOphhEyn3eaba7B6gun
l3if0Lza6irNWU7Hj7RsiPngloq7/BXOyd3oPswC9oXSHUPhxM55l9rK3E5IzRVE
dPeHgiqajESQiy6WoBWJPWmcJr/pjQG0XFDnOND8pm9ODMhI965tBuUan+4T0DZw
3r5153AqsjqkzPLiOnScW40bO/PA26V2vyfBo8wKcXFtHEPEilhYi9F9dgmEpU2O
7KaN1UHuKPUPTZLM7YV0CAVZeK1ZOKA5N5JYd3XylCUxHvUaoN6bU9+sZfGi92+z
tsfwPEL4xwn2C+vgWT5PxgPBRP2yhAY3IXtgYpbgQMKxYvnEYENDSFOdTaG85j8g
2TkWEW2eMzGXkRU6DGkeKSQaFwgeFzVofuaNR6ZbbtdCQuhraR21ndtpoBNWPAFT
/QQHne0nrk/19Sg4xblRdbUT4oqHscyi9gWrEaZ491uNnpeWXbNla2dljkbH5Tqo
9dE6b9cZ0GIALw2jkpivZMt9gxIZGoHkuQn4Rogw+AvbaEDyOEH+ulmImnu6yVNd
8GpWDsP3FIi+IheyFNtcJ8QccvgVaVBpHhWKDWUaueLmXhZ4usAU9ORG0230+gP6
DBuW10be/dd319fbME6TXcfYmf6j0Ec+9h9CizPEeQmcZXBeJ/8MjmWfCGZrDM1o
MwBzrluQKQvqPzJcBXWNgI3nAtAddxKhPp2ae9cknZoTP4AQZf8hTAFI17flkQhZ
6i2MRQsa2Pi5bf9Q0S8njDTMiJ8eTRjhnKw4YqfFLJRwkbOJ+3Mz3TaGASM0+eBw
1MkoLYEkpxMk3JXlTO0c/oKA4Sc01JXLCGCLNT9Jhj9cibov99zEteeQBcnIZBWL
3aa7r0H2qi/yaeSZrVWWaGtHxSlgHsFfuLVZpMTXkhWIsV8b4dMOroOpAP9qjloH
TjPtgMz4cWLYi+gZYqo7YHRZxMB3KXbJQXouFnV1G8r2yWxXzYSf6ODrUu/X69ro
syDsBkhSBuCgK57iRSs1sXQazdhMGK993HAZaiFAhoxNzcAh0/o8jCdxHAHdT0o2
fr5hlW+I+ZkZuVnxpIuv2ogtOY4tivo6KFzJa3Prx6AvkiuLUoB3r80pOPHIKJHc
K4O83y2LjXQd42X4Fr95NEa9zbSmGwDMwr2ALOIeQ9aYZZ0hVnCOxtdPCk4zZhBA
/Y2n70OkFWTtkZmqQpTgfmXkrfP0bReMCsfBaXpODC+yCk4g0ar/Pm/5TUVnMZyl
3rb0j9LcqtMPZwfDMakEJiZmV8T49HHn/b+CxMSf29sc9SzIVkmqJ5SrdPV+WW62
/vUBZjnX8z/Hlgpnn1yoxtIZQIYqRhMv8mXaeeiAhJhA/ndLhVKQHG41h+wPx9VA
tifvhWczcxB9f/s00zOIEvtg76eggi1iGjEzqNJwd6FL5iwtktPDsy09rwOutTrb
ZvvAYEE3LT+4u9+VywMhNYouzmM7F//vubFgUXOw0bBuXas8T1pGX7+HkXePYnDg
1O+IcdEr0ow4BTt57Ak8wG+5c5tql/mPQp4JlgAoqJS6NIgfPJTgMdYilkhqpUOw
2X0RpPEJdIgI4UkGMH8syzVrAJxsJa8D/5JlhwqxX1cVTE6pCFbyjsQA7CEwxuJX
tXIy/5A1y1HaW/rs0DYfRlCrrB9iI1IrO3/SS6LAPdBZbBsY07viZJjBEfOQ7GlD
EH+clnrfoDgj1nv15okBul/suAeggWZPAEelc6uESqwKhNNLngqDOU0SK+OAinmf
yPbDEiY/ejDU3BKv6RxQt2oybc+eBZS7LUJD+jb5/48QTJmQPUBgX6+qSg4Hy2df
UFvEATWQUXd1n0cQNQdT07WoLoesBvKhkGkmBA13oneCnAPGB1RvQVrWqpycefxp
H6tQzSC6F4J6wR5wWUOFg66DINTfCxIJn/OpswlNMaeXQ8D1Z/KQhOrcQraxqoxu
ee5n5dHKfRdLaCZnekNAbtfflnpYed8lT1y0Yc83jrbi6xkWQMCO12BdPCs7cBw+
/vegtBcFa4+ugQq/UMV/aktz667408NZvKXus5biEzMBVh6xCuydRuw7B9uacRJT
8IHNYmlhHTMZwR3OA8Ohyz3G2vEkqIZcXoIA+5L6nYHW73+hB7mLIUmDJOIlnhcA
Jp/OvhawKWmW/w0p88fPOyf+1F8/9H3L5GAQN3XnaUOwP259TO+MgAhrQzwZzf12
f1nIURyhyO01UARAyKrbo/D9vy6atZUkYQOSvkhSKW3r93BcFPjOs6bTdrSdkqEA
o8C31yJg8X4rMYK734MwN91D1D6bk44ZSspdkm9xmGqWuUqhn0Bk3yGbxSjpbTHn
osb+vydxn00r4KC1sg4O8In0nQFWMmmTGlIPhSo5dLOsiMqql0UnAppaE7jkVaRw
pvbURws7QVna4NM3LJkXEKBEX1eXrAszTGw9kFCp/4macAX2w5kBnxQDWCRIbPfy
CHT4+xpXbTv++C1tU1/OMJCfemBNH/VNQZwKj/lOfWFbTwfFss9+MF1OJ/vM6sbu
f1EldyT+mqgzraFF/X1lChQGr2PntOwJ1aY1AIpCayk6r7OKq6HlNuCetnAiTTWk
EO7IE2Qj4foWQ5yWZyDkJKSRehEg5ppY+GE1jnTVZ857bjcRvLINsAyjWXMNgo+w
/t6csLorVFeppQngj9h/OHu38czHs4tOf4mELWJC51YbBaTrdhTaEJE4YxboPDZG
GtdyVxu96SCTAGa2vJJoijFKIOGRRhSwOME0ln4xqr9pZtVanR8A9BIx5bHHBDqS
fhwQ29/n9y2wepXZNeXm/Hd40T7Rzfbhfi6J6lBCf2iTqSRI69puMjHMMU7T7I+K
6152EuUkE2+PO3gkz1yVfNgqQEH2WNvjRTKixjJgBfKAlMfcZpVErQF9g4SkMn5s
kmOK/2/NEwzLgaIlAL+XWMARgMZettH29WiIkS5QVGjSCKFDIcmHUFrmoIkrXPdf
kyKaTbRSo2s9v94SbmfYlYUPCvMN6uXo1GPpOIULOyJysshkuEHONavF9MNcvUMv
dHPRN2w+1IiyYDMOwP0u9koJXAMCtL1A6PVWn90ahP9aImslJYQw7ySLlKRld8h7
QM2REQJ65rO5eG6Cq4mEKgb7GpXN7yR77GCNbf7mPwyj4Pk89dDKTZTYVTzZcD0n
ETsERv5jxyAvE7FNe/ia5V4igV1EMOZPxpdElTDyWXTRHmIwhVVSnrxaHuSYPjmQ
FehDBkQiXaZIgBg3EClV/AvBXYIu4QPla0DaIH5p6WVFgwi1CvK4Oyg7aye1vtLN
XYSWM+84wIFBTu8VZCHFvx6yLr13EssXNno6i4b3eyr0o3g0IC55Rcch4iLwsHl0
IPyHtxPNyvf5w2d+sodgoxplYgv+37sq3sAIQq6gfREZhKgzbbKPMad1P21V8EOr
5pnJoGmQWVT3eON5cj0R0G5l0slvTrWwu+zrnHqJTlkH2Z0JUUkZcILOYy1ISqN+
ZL/BARR6ElrBRxfW6gxcICY1PgbuejNZjC40HvD+ya9aQJ7Dncf8qRd3LA4f8tJK
vE+73BJbT6DtatbE7aCVOsr/w3u+xqHzmwUBn2g+3XZ2+aCfHN/V8P624qoD679K
b0Xon1ktEh7OrdwDKNT/DYWYKzFeRIfFJ+26yqI6oKhVJ4nVwrw10CBFaxqWKlvq
US9vG3hL1+tkkhc8OdCKGLP21y2clL4o3XSc/tJ2ZML7KP68auuge+GZex3lNPBv
6bPHy8jRzQ4Z+UyowQ7lDKsqdvnWsN4aSu7c79yzXpCfPWZC2++peZlge5pAqacj
iQsRII5ZVQWG5sTeSp8AXwC3nk0KAhyTP58T9B22IB7Mk6gTvb5GREjhDzRA7cjw
szU69zXqGr/7Hy4Gpk+qAZ8EJ/HV2GVDDA0wnOioI/GJQsJb1cbhx/lSCaJVDU6H
xTG239GLOvWLZxb9pchA6X4twCFINfQ51oJ8wlEIr+j9lgYkRmnFwveRTBdM6Fz9
311gkbbl5d+HHgN2EVOx+adcKd8B01KdKgsr3JT+/ng50bEcyYzeeTSMZHyaBbRw
MANiLdDK8IOn15xaHXfDyrOqzLjexRpt/R8JyCLi02vGtGxOj3N5vW9gd4gYTMdD
XHBdCuziU2XELgUL9efD0XKq35QK4J7SVvICaRBcj79zoTL0odVF4dTWrrwKuRxd
F5e3OH8Sou2VgcdX1HdxzE1GNamKM15N4FhCYCmwN3iFZnT+JXjoRuG5W/9m0VBw
POHTSjMS7+LOQ0hvvcPFHuJJAg6PRSGNYcLgzxB1ejpZU3AwoPQdZSRXnaoxaXys
E6tnJ8hRk7ERuGqItnNi7x9gocu8Jbm61XC7OKNqKgPeRT6D+DIwfdtrq8QAHNlC
y4FHsStH66jX5PrTOv2nyLRaTAlo1dvaO8N1IOVmVYaAPlZZSejZXk1+vWQriTfz
8DiukN8O7nBf5sG9Y7hJz1Ti9ygZhct+tBsGdnarkAQM9SDaYNNvkjiMppEUR9cl
wdhYslZW8kIUV0xxncvfTRj1g7ZMnA8LJKfgo3MUtRSB71GPtC77y7vdmvUGw+fE
DCkrimx5FTi78TmWLbThgDqhfVgIVpzCefuKuNzAuzMQ5SjKPgfpVlN7nVfNSPpY
dXggYO68br4Uctk/A4XOIubhd/lpjHDeWRZXcUrYaeefUOUd0fTG55RXHJCVVEn7
8ApoJXRhc+rH12h1JZixgwTU2ERWkD5nfbQLjkg51XklsRBqMcCAiELFyIJFoKTZ
zWXKSoLs48naPlvnA90lpcQaewZRoIZsyzY4k0FRlWbNAp8UwvmgBemS0p9tUE0q
QvaHxYzuFSo4yhGOoJ+Q5wvr0cKN8aO80jrvkwSLkHXTEbqGqvzojo0ovk+bAmYA
IkgakJhKljW9CYlaLOMu1vMhUBm0kobVJNa6RuwGAZ6M9YBYY+5mMW40tkgtWm4h
6TNJ0jY+K4c/JWt8pFNG+r7ZLsfQ7AlN0sEH9Fq6C+QiZLWmY7ff/zLNHgB7FW7F
IgPL7OnuAWwEHvsh1oYFiJGxOUUjPlaO5ngIdIcwmOY98qgAXie7Y+GAoajBvUSc
dcCNeg/c31Ses3Cv85wldSBkYVaBtZDOYZym99Vm0vncCW7HrLmKw+9E589InO5o
ywfIp5DyhAsf9na0zffoTmHOSeoF/vMnNz/WQqSV047I8h3oojdWHj7hDBBJc72F
72jNOnPkb31SgYWfWXEmZ8EF0zhqhIIlOAZKJ2ou44iaR6GTCCW4U+uH4pVe3SC7
zGdTNT4HWz9/wmfFhM45QdGJ6v/3tgSCskhSywi7CD6iB18NLIO3hUASe0tlUfKy
I+lr6rX6pOUX7yvLo8MrZDsdCWoJmRtAgSnYZ40UNIuQVxkYIG1vTFDCpiJ2fxeb
f8RcsVMaitpZgSyDdRI514ZWuxSBQWlJPvRTNk7lzmwwi9s7BLMhERS0weKy51gZ
+SPR0YqGDp/2zzqg+X2TTcLIkWu+RI2P/qP3lmr50FivjOBRwxMpe0MXXEQuE6j0
JpgGdmLzBf4LwwEfvbeEJ1AjCyyuKOgIETSXuVIkRqnXyITZHgxYxQ+z9kG9CKM3
s4U6F/2PnHvuYT2zZ0R4FCCH2Rfu/QF7dUh+3QBGVHLRvQ4eujAADp7eRLQ/1kBK
2AoBsUb6MUlou8n3EEPFY9pkDZLxOX43LU+ebKuAYFe7e/EYG7PNWja1IDRgHRh3
bp0+rElN8E7KTNsgYNHx+foOpMISVqqzfDg39P5l4Ec0t/3wj4wWPvbrAGsyTjqT
u/qbWo0O+QM1861xmY2JgNu1ZXa7zhiEstKVxDQfBuCJhhnDZR+sai0LPeHi8Pvb
xow7Ohapo1Qmm+uKPn87d9HlDHtoi3yAk7dO/97wHXBmGMLfm3LzDhDEcPK/EZ1J
lT+2Z8DnXrARbIFVNMhqL9wDc2zfdfWsKJHehkPzoArsFngAxQP28XV7iW7LwDeQ
vO8736EPaRE78J71AICR8HONrge+64tFJhgQNVEqHt53qgScSH+lQYALyC0T9yYB
LBvEEf9K+sRDZwcUtghNH9bBJ3pgkbs6/2F7QOc8pvbd949nmdy5M4OLotot4t9h
GM0UW3Q9wVrW5jSuZOXCLoGf+R2+eJieM1qyFLbY1aanoRedO6xARlvStmQDOGCE
kkN2bWK25pUSS8GLhdDIgaKvipl24AkvaV2YMgn8b6qKlhhKcvZzdXJIa9B2rr5+
tfm3CEklW1oxUe1jKRod5yZMCbX7x7WSXGb0eCU/5kUg0ICBkUhGlEPtrv0C1Fk0
7eFOqdQxJZb4j2Lh/j/oDdBeVXJdEivHwnx0pp0F+ohSXgONrBHNKzcdx1vMLdb/
YqapsOwCZlFJ11E30ABYPwTABMZpKzMtXRcaiukQLzVqRPLjUbmhg1Qf1gV0Pt8L
Di935nB97wv9eEVnNNafTxj0j3Jz0wofpxf81tZ3JClMgGh8REYnZJKbAOnqGMbX
uxpBB46MDB2wtkdh2ifF2F918g3Y8JGvcpu3MAjwp8//rKy5MgHfKctQDxiWObfL
eWcT9ElvOUcEWNKKDnscZXo/yaNKxADPlBIJ+4YdLiZ8edN1HeHIg7Su4A0TjPBG
+ooqNAnRl0Km/uHQdj14NwZXNJ0eOxC1DapxUM9JTVCp/WtdEhxLrfKYI1xkEMI7
pufqnPqs1c5tkbUVywldsoVbnLnlusExhxyrdAiJQQ/D1E029gjCHxp1vdqSfAI5
lp/WoiQHMBVl2E9T4Qr0ePHFu+8Y9ba84za3IGKybQWZhlYhlknnFrdDhuBQNgDW
OYmAIPVXA6ZTWCdgwo8sDfoOhZoOLpWojZHi8j1pSeEClglT+F8ZL+igC+I7IJTP
O/uE26Y10DB3mWIdSd6D0zh76T/iBsDRw/uL1jGIGjfOaSQrqntoaRztpj9H23PP
QXen5IjW1qlOeHFF2Lccgs5/E8IdxvuP5Z781e4FJ04xvbT1TCoBAxpJh1Fbq7v8
EyMf4YIN6f2u2JBlAJkVZFLJiYyEfi8V08xIriAwFw4eIgjuP521+NFOQiwS7SEy
f8HB1sKMonWREzvH5si9zrom0In0wxEvrznw1pELsOMjwcrX+9pUC90dGh9/Q6rA
wKiLMcEuoYm1hR/iftWZFpQN1dCUrslzkZn7TYCePkWAa1JnH76BWvyZ9Kv58R5Z
hsQH0bhLAVGmV5krtxdkPytZPXdbZKUYcrcjly+siBeJTx7DRXyEsgVc1+D5Z6wV
RL9NLgPcXNqElJVi/hwSglIEy+Dy2aRGXw9V+HZ1jbkCdAqwyR3zzzthIFdad7HH
TemprR9bAwqcVEoYdqgtcUFOwWNUpV5sXlje5zPVlTjpiki7vgvTmFEuWi9SG7Oc
iV25lEi3Im1lHWp3MkuMnwDgwEMv8TjhEZa4nlsRbOpa7LkRZoh8tBoNyt0UPm6w
0liyobDVAp0KHL86mZT7UkShrQjK59nj4yjj0DBPSA7WaM7F93Ii7rJBwJzZhgcg
s9whWjh9ifjqUr6YEVp3+Mewag48/YTAuxdF6wFdERyye6N93YRvjaWkLKrIyOPs
vPlU6M/UaoY1a1jWcngH20TKTGdi7jTUJJH9CcsILiW0wFjSXzV+IqSC05dKHk+c
WBF8rnSpTF26q+8LjtSfT39nC8TdlsQ7Yr0tFcCQSK/hvdlnGWOLmYYtJQaDvO44
FQzeQS92WGy4Dwzd1dkcPNoE+r/05uhB57mVTO5lJTqPiOq2EQjyFmStddNJxZtc
7o6R9ij4RtJ9dPfLoswOc+s59Owc1pb9RRdYH7ndisAQVyX+FdqSg96Yrcli4v4L
BLaJqhU3IcVLEYyRBWzocC90WXDYVuzof8yBI09F0DnjpsM2aJaJsp1HLYgwd7M1
ik41VfmMa7VE9upL7bGpPFT3ZLh6sfZQRsK2HGQMfREs5+1ou6DmKpgm1lSuTxyA
FCTDAMqLRx7Rh+tvJKkuvqf5/uYIo+VQ6QpqY+ChJFLK6iVWgWNLs35FaFHG1Ox0
7v+M8fYXZRRqTGPyRehFIXlsDhMJSmHFTtJEKJFkudUqgJJ21Ly3LZjuZPaAkAKl
gImMLufH6dCWiC0b3VNr9UE5O8GmYjrhapjm5878Jb+Df3K/EQOOmTU52xwbd+3d
TjODCRK6RmBxAs85tEPwaNPWgmz71ARXUHtadM8LwKIHmSAV2A2Q9fDBrMnUdexq
0XWdr8hLcMJ7Uj6lEBeJGrMPU5M2VuaNsZtl7PBZVB18aY+t8WpHnh0N4OrqXUeD
WwiglsRkxlzZAgToGbZbhx1kyv7Qo8G78Mw2oq2YYCB2FifqNgjFec5geXJHJA07
FM7JBeUZuEb0C6/BHQpdvI7au12jkTN8dxQ410uk3p7uResSC/dQY1cvACtCI2CT
W0KLQ77BO4TGZ9k755p+ugjr/yyofqVmLGNdCxYSg/K6JhtQQ4CJMHquPgkhmeIw
sLmIwyu0mB0NV3wb0L1M0DsVY0npiflpC+JC266s7IB6GDs0hoXM7/5KPeWjG4Aq
oKOUTe6ZQ4Vi99rir4eP3BRroO2EHoAxAlglglTQYvURzEwTLP2D978HB/XRlfAm
rPfVwe5abKjJ9oXRN58518uMtwplaaEn42C2i+BSIlh7E4W5rftVPMDlEssAW3Tg
pmeCGPy+in57yQG+/j4XYYcLnxvRP2OIPs/nMVXZgiZxrGhzXM1AAAcFoxUgYGEO
KX/ag/VjVgScYEGAVREWKGSjafUcsuFlveYmQUfrbh7Lv3R0fQNl11fZOrg/zaZo
TsaL+Xf6q7/J8GVwFgBmuAQ3j3zc6eCHXAJ/XYk+jn4vuBoGxDz/ys5ERSe//r5o
ScCqVGqcwKOQdVZYdSB/ErtBkkCjEr1v4/IbBeKZqFNTXscXtxp0tt5bN7t0fhRr
fMEBS7RqJ1zCCRquspwbBtru13mrqKChyYE2OSlhBkXEckiVYS/jwxeV67QzQ5w1
ZDPfr4zYgnPMRvewDcNGIGNOfLtNh65c7Q6Grw/2guWnjBfK1kqWNPU3PpDh+LY4
7qo8NutwPMAA58QAGHMtqcWaj2v9hd8wQ73+hITgxuoQ2TMKKumGVDuFg/eOpWxq
t1C26rhrRxqet7Swyl7isqk8HNgGafkmakhQvko+5MRNIfg4A34HtHl4DRd0uT+J
XymTpDCUNab0Tas5Ky9ovS6w+17poFTUJxALtL9u8v/mTkELb2/xrtud4QjOiGQZ
bXHECtXqIQbz1GlLtAvDrix7PrNcymKD6VKi88bPs9WUiRKGRBzrefYYrAx8jnw3
EzyINlhgBzg7n2wmlaUBOXzQXaV55btWnA9q9aj0gRIIMuAyheWQIEBQixYWmChB
i3Jh9H1qJ1SPiqQpx9npeYedQfeLvDa7qIrgqMSZ09j7iYaug9nR1Dn/ndJKaQX3
F+dWTv9XfEwNgd2g8ahWT/WkrPkEOSW7DMhl0M35ODSYjMgMbAqMCNqYMoyshZay
n/s8nulrDdjRm3llPJxOkiAfP/F7rhiK/YT18IstkBDMdz8n+Y4tJbJ5B2dcIpYm
mGzrM22mKwJlfUNURuICkILBtYNUoSN2HZP9yCylJ4l3WiTkb5p23YHVLjznCqfH
ggO5iv0aaYfBAUmyrFlMPjPAXMU8jY+pE4QTBaqffq2HEaaOA4RTgwlrXSm1CfjW
bp2ADECj1KAJO9svWQnLz31jnQNl1lz+5dCtOqKhkgVGkHf3RmiXKpsjw+MIhB21
G8A16vnlA9LFJ1lo6ULBeTO8/h0fymaFWtVfwYSflN1PTT6y57ZqWlmd2Ldlt2wf
fgbgPCXHjmvOXEpTdCsbrlbQ2SDnKWbRqYQlhWyxTaN2Wr/ZYk2RK1vyO1l5ypYa
k5+wE2L1ZtObGCkzh/t4XP6o3xFiBYpArgO3Y8RlSPwTlgc3AwqFZWd5kRDJ7ugY
AjCnKXSXgMVK2DuXyRDRR3EF4QOgi2ualZ8mYDQp7saJttAF6HUFMbmrfAVqnZKJ
8wjoBehPMgUUUllGKDQymlLybhH19WW1n0492oTqA8ISG+CjFh3kcH9Q77HswVHT
wVgy+fJiL0MzKTw7LyEsVFa8Z60eLxKlBZsAAuZsxMJHRzW8tQ+m0y0/uybEW5OG
kZ2zx61bjS3qDwDpZ6ReUPIPcMu8lJTx3ms3AdhQFkH29n31rzd7xs3H6oHbhY8G
ZrVlxKYRkcHEenSpcjjR19/sgoAlpQfWIOeM8q9LGn0u96pTYmtCFc0OtEwIc/IX
mANq0/l6pbZ5ArRCP943y0/11wVl9P0UfSBZjDiPveSXUxIQiTrodLbl+mLUWAUe
onjIRtXFluH/Yb9F5rv8JVPyo1HuNIpIUswaYKheXKm2QlbtlBTaAILfX9CTcQbF
Cas1/KRLdrhUAkzWrNy94GUYl1OLOpA6uxIVYI9l2RN2PYaIRUGh1TLGJlcn7tVv
lGRR+3fcEBhJRLAgIo9qp+dHJgbE6VWwjNMPnUOvg/+WE6ZIZMqdNRW2QRy3gkUw
gUMdouSu9O2zHrOIgF+XuTj49DWgDecdqTnKNekqasQ+Kp9BlRcmXXrTWE/x8GxR
4r5qIRVWmMVFL82MbQnCiA15Mj7b4gsdvPN+AUis8EPNDK/8AlOveJe4kBXIMtwW
dxzP6HHgGUSjJ8sf9p7gau+t0si4vTwxuipr/Wa6qevXK3a3RozYQSP9dnAXCVL8
ZWc9Jfd8gdPjn8fGIszo4iHV0lAa/HereNjcjnS/Lt5HBtO7Wt82R6HZu1IIKoFP
Rl0p9Cm3M3fj2U2U7Hwb04aTwzciRfPjd5G0mwZI3cJxn3eSYBpNUDZPCyfT2yZx
qZdVURDS2lqUS1vm/TRgGN/GGnze0EJK9+ISsRRBVV5TvrEgcNexmiotVychbnOb
ExTLSt8qolYHxbEB/dfpI+xqV80WChZ1LFTRLoudfQncXgX4htjq7T9zuN5BxG59
Bjb3R00RTSupA5JKGp9iszjVPw9kbzVzXkqXWX1gCQ5i05Cs3w+s3SSGbcZ1+RHL
jZGJBfYOtvO40+eq0ApyG9yVB7T88n27x/gGNgOx9C4HHukKXW/t+VDbuAoruzB+
aYsz4ex+bNCjupnYAkfgOBig19YLXHNdpMW4Sl79VLq6Q+hhJcatSsiop5X15ZGQ
LuYW4XUODXRPqEq8aJpj+Xvx/u319Jy4WEOF3m8YXKTp6f3uL9rOTbV+y4zEpDUY
wFNQq7rgvZyuv3Vcf1BxnJPXTUfdztOpaqukjGXwXx7HNRzUPr0wcTfM4gDLNM6u
Dx/Y8vfC1tMhR3wlpF2ft5Fl/LEitF7nP58Cpwsvpza5dB4JB/+bsVmPs4rAO760
+3Frff/EeAXhILDH3rsQXCFHABLY0AqJts5Yyj0E/DJ7SHbkfMTgNthy3ltWH62P
E0s75FerEvd6EqBhxLfoBh7WU7j8xqvfjEQJnE+4ys43VmKeDRDvf2atRtR8lJvZ
MHMn0o90M2wISy8T/N3OhjKnbmWDWap2wuni4yx88hEjbAzU+FNr9fnZhd7mpiKo
Pe/H8svPAnuy642aqNZvcMnJnk2oYOq+cT1hkwALncHFuD8DC0KNw2VwYdoz33ex
4VTUpydTDBsEdvS1nEYeHUtDMbO0KZTcvEj0JD4kHNxVBaha4OqnqxQL7/j9qprq
WxWGN3DUTSQrvSit374D2ooWbw2s0B2b8gCW+xo6o7MM18clu+TjJ7buDPQvTKqh
HVZktOh8lc1vU7A4Ab58/9gy2MvwXVPgyUsgHJEvE0z9okVNNsIz66683OJwvrj9
Afd+2HHhB24fANeMrp6LVveyKRF6MkHCTec/nF4PytnYz3kNx3Z4n1KWtZGpCcRI
sSB1JDloPVVQU/zKFm8JehWVrr0u0HUr2VoGLhbpytMyxLRHKqeARLTQhEqSeL56
/MFD19V4uiO7Br41QcMSms1xHPdCoF0kyI1ZNCJL8T/w1ZhbGFSPXIB1batIWtFI
f5KoB7JVt3mBdH/CkjEHSL1SDrAUNXDJ+n8q8TUORrgkfXCbVQZHwLZNBcIeYYXi
zTRrzjUmN7o+Tl4x1JZj0sdSSVjOAQNrsRvwt4C6yEfgEvuxg7TzpjLhs6W2BTji
Z1kxpFf0yMWn2WGlqDJg8sX6N9GYWue9ePKrdawGi1OsinV5cFkZ3nVsM3QddaVd
U3ZT0sMnzatcQK+OAKSQ4RgxJNeVG+aRritInuM6mZeUgCx6mIy5Sqv+uyS0dcJk
6rNsrAk90KgPn8dEKYKJITB1MaSgrWQfJWz5+n9OFIfaXF47kBOR24ALpWFwbFbN
qbvJMiaf2lni8fFPhSnDaQWlxX+tNXyrx9/4SexUyWtE1gFtGwRouF3R6qFUJc75
Q2xY2/hm01oPe+Ao5bM+2IqShwmBdBXZqJY74KQvP5V9TtLp+2ciyZg/3Ddy96pX
r1VyP+NGuHMdvY2RcGJalHehxFLcB+5FD9HL9c7gYp/6xh41YLMTB5Nd0Zs44ems
14HkALL0LOZghIyqUQFp846O26pYLXXuB1S2i0KMUkJ+m9aKmBCThmeRSGEM9d1Q
s1/rMD6r9/br3vvG53BI7Q5LPpLO71sQFkS+J2y3H7LFR/JFX3ZYWHs+PCRjdzYr
+61ldX55/H3Zch+uPwm2K8mOo7HgVnoJCX9zH40bqWS4cOXHEXgLrxWXxZJamgH1
sprdBQJmhGb6C1Rlj3Tn/1X4IhUK+ev4iG0M5xCRO0sgAYLazu0JS9eIIIoOVXkw
zniJm/dNSbxEDXlYSnL3SlmN0Q9RA9Mb6a3Wi/qmk1PmMcNGNTqjculktBJ5lBQK
pBwRan+LNY824VanIh5kLxbWTuH33rae0g5Q7FeqY+PAtO3vkon2hQ/gRReXqPh/
9egssG9KaILxdfvVhB8WetEMpie96uC4kBG/+f70gJthPaW3AqLghHuIvYTkwNoI
Szrpsdqyt6+UUYuXtQI3HOwr5LNuBUillU+4IyD4x0HXV/jYxa7sdy2e7BvJozs1
i5R6ryFLQGkLKAFGObVwXH8es2I4kV/NG7YkzkdMjqCsuo5wM+a2Ts5tGyTTfkSd
yoDMUcQzK4fp6KA0ss/ZVBBdNdbsx34WO/oHoGVNMoQ1aeZwHL1kta+rm7XD87lO
p1Wcvg73hf8Sw3SNv3OdXHKpnhyzwmF9R1I3HiTZaVWnIKswFMbbx6T1USrv/3WA
WKr1M/zeu2IRVEUlZ9RAgYY8uDyKsU37sM1UNIiCoXRL6nPS+aVoJGkivMi4VVnz
ZoBV528EhG1n+RKygzT4NBWwjAUNGY/eEC2kAUererk8hlf/qHKuQ5ToKtPfsKVp
LfJ6qiCokyK4JZt9nFbbyUkVMGsqhL272vViAxVmxRzPPpSOenkcfnI+N+M8Hgor
QptM68gI50ISVmIyDZeSBShUyFs1dqnY4GJHnz1Ykj267UlFWbkJDh0u2jolZuo9
88PDbhHq11WL+Yudl2Cm62iuGCSdDJxKuGnhfXaojhcjbFrzGvnZCVGA7drj5MdD
x1d1CY/yOkS//+iDfJ+TXwTN3WWvUtcbtPpOQuntw5kVjulirreP3HfIPftw7HsA
V+krHQsJAy4Xq8MVD521h2iJtj9FtVySRK37iaZOdQYF9WFKZB0C/wEVYQ88FGPt
fwx621aPb7MB4MsKe8C+0xfW2THe3SvyTxOHKHU1GFvC+v2SicLNGctUmg3B67wx
zB2lc8KwxYnSLydZLVF4igKc2F6wyi5wsmdp1WQv6gV5ncmbMfSvxVzWEf7Xif5e
ImiOxdOJJcYvENh7BoEMq3bxbqXzqqUNvf/WRHSUmYAUiheLVLMmm8G7MIZgDwU2
rEl0Ai5jaVmfs42A1PEGlI3rGQW0/vFbat+UVFKiVfzegJs2/52Ohy/2lb8N0BUv
hJRlwLhC18/0XmLiCWt9WuD4qhC7NY2GjKBChlDGSyf7VVumflosPNej7Jl5/BGz
tCPPGwTyPJqkXAOG7mV9toLLRVVuGFmkNnApYGcC2xiWIDkb5i5RB7ULdx+l9QrZ
mvpJYBo8TBeJWDbuA0jYdKB/b4zXk3xUA1AJyKqfTdtSAKb5w9jAAdM75kBxLhvd
0FrRSe+fPHFhW/Ijz1k1vxRr3cXO+eXym8x0lWriCn8q/grp82qBH7wXgIuWmf8Z
XPTDNHRNoTGfnBb8kw6lhRjmhvnqaIQuBm1reiqddrp1ov0OqmlpOqSYDlKtCzzI
ZcI6JhtfNw2j/CT+X2OFYP4a49olgoZcHSKM1Qkq7N7lZoVPNiplu3gURG3VYAYA
d+xBAa3a8N9ulGvIJR0SF6QRPBVf5XdHDzYvKBTv/Lc30c7SkvP+n7xTtnJKLHS2
Bnh1IvTFiZbJxPPI0jgH0CLScNm3dzfZ+rzIt0IzN0ZFOcwX+FxQeRU1+oFgaTJf
3kcVk3UQhlKImpKQO7u8N4VsftwaNT+2RY5z0vdpwVbBCVAm8JWZmKVHwNG7vd30
mHsHDHnMigsFRL2JSfEzNlHSai62+TUVyL55cyhbuLqWzmuNLDcf0uMrtNJFJkj8
+jTQRXWdc/NoiWrBbl9bgoOFr8PhVwMOcqtNYRo7dyM6CQ+di1RKeOu4T65ej9AG
Dnm7PJkLVXCuTPdrvWIQusJdKr8DVc77sc8/eOTjwJpJnITRRdI7HizdID0CS4vz
9YV2Z0mLOSUH6oPcHypfrq+9XzpO1eEwa5KXINGdLsGfMZxBbU9QZk8qGtkhA49l
alXNueIyo0cJvFf7drZFeThGFYW5LTTL0pheM9NQmpA265W5E3yRMVlnPHRlFTmm
9pxjXFKOuCvRGa8gQ0DH5JaLQhwqSWXaeWdmMxyPM3JrGyUv65oK/+p9Z1eFjUe8
Hf0Uo7SAhi3t91mTvGQ3WaolfQiedTnWJgVfxWhfac7fkdzweOZc2EgrH2vBvjmg
JZy1KfHftZtw8CJKxYNDaucq8LCBBO1+7TcRD1QobUlzDbQgIb0oF4Ris/j1Gx1M
8PaN5NXn9mumrgSOm4yKEARFRhDgSdf4p/acNIAayX87tMq6ljmtw4QFGsk5IiVv
ERPj1+7Sk7tl6hVIqrId3RWfCJ236UoOGD58p+2mDsIy2j8BxIGV3wZS793C7z5G
nw3Ym7TNnIYj6zyMhb5qp/skeLI++Vuj8L3JoO44jEqfKHR/vujVqpC+zDdF2hvK
VyE9vNmTsG5HTbw4cGBEWXhtlS9RLXxoGD5R/VAItMh4OVTQtNhZV+ugUEK9X7Vw
wnICrqlvSC3/CbMRFVjStaT1Vhhc64ew3VE9n8zap/Rxq2CRHzG7HFvuImEtgvL6
4rofU3vR+Hl9UAt/xY9G4NvmCG+41+bvpuyRGEdjV8yRhwPMbk3Xm6m4R8pwHUSf
F8XhM7ybMSjOJfaFLmGHTlsHrUDXFwBKWtsF1S+eJOGSeAJ1f0kOpXEYnEQ27eOP
1VLCBahkX4L+LMQJ/xq5uzvTSLuhmWvOXWgQUUw+kX3NUISpCjpIrVyllHHSliWw
eFs7sat9xi1TGYA8s6uadBWOpy7YEZvk8ZELA8KZaykRUNYb31HTgQcyLOKJLCx3
OpImW8TPc3CZL9GQZNYXVQOpqY/8Uvhic9m1qY7bmPkT1qski486ucCrt+8oEWgm
fITlL0QwGDdFHkD0vlWGbNze9voO4AwhjeN88T3fIsM7l1+Ikbo0WvEWIUQ34u+P
jLpnMN9n+m3mXY4reyOzAtMIyP2asBIts5QKc4hlZNUA4+7mJycN9+G7GubcQ9LV
hGji8lbWCB8VTQ+VL4SASu8US5liVheM0H1hOSsisS1Syuz+Fw5AnimVX2HYp5Nk
JCMQ2/tbLxNFpUmwSxBzbf7RjsYk7zv0XdoyMx6Qtq1LzIRAkeA+2H7jYH30BfTt
J31vZYQRIYtA/l9PRVdvqNfRx+wyI+oiWDuuxjAMn4Nw0D2SXZQcjKekUxZPl6oO
lH3Ot+OpnYE677HEmQQUyY7WSmHXea07SAkIF/tOC/rmJ8wbYol0gD9s2posmNGN
Ijqpq86IkDQyUbQ3utBhd5VrBMF1f5bc4D7IZo5/OmJyxDLklBceLyUGmmhppZZT
vdVeXEqIliKdmfuqA/vGdda+5VlTxhN0WyCjUGqapuvcMKVj1HYawjgbOvv/zEJf
iN/djQPPNOreST/CwZr2FQw4OF55m/y5RipJ+tkJh5qLznRrXwIbrmKCXGLh9h79
dTnaQHPJk386vvXNbv6ZRNXJKdAT8Wxhc98yLT/Y7QRrU4BX1ENgPsKNc7uZ1DBj
AmaURQQ0E5nFL5YxqW6doN29bq/u0FPc1KmLYHF4IBNIPZHMcayVlM6jVxxMxFwO
XcUfVyY8PPNp0BvlMm5MDSIo2xC3M/udk18F9BpXuhlL4EKBIkjNZkJrr89Kd6iz
i1FcFx/ejcJZg0pMhvXkw5Joi0OPf1/SnSRSMlJayBu8uSLA8xSu7N43yRcSN7Dy
FKPmUVSlmYK0mIp8uvIR6Vw3QSTwkvjJTtU2uF8CiFmnoYil2+ZPSrXwoqcKhrQH
UnuIgPENEie1X//AbnG4uxI1VXzgDPLxdd2rO0CBtFgHkTqcpwihcc4H96+s2ebV
0MVy9T+Bs57z/pJkOnj3yJjH8oAn9z2IqbSCKLj2qIMD+M72d89Jti3d/boEI7yL
sDXJ7mSwG7J+Z77OIdvSDQ4XFJwII5TUYsCw29WetRrIfDg4tlQNQu78e9IJkkHZ
SgwDX+goKQrpnobmxK3SU092sW/INDQgAWeqVbQqM3oQQnvgRTdt3CMOopKk7Mxm
KWJotGKoIr10OBqKK9paOIh5VbYhAiEN1tK76JiYCDmLZQl677dph8qr0osx7deX
mlXHRb4WeuWh8SWncmYWeC2wsohA090xRdP5Pve5DuAFXalYnMacBqE4/BSqAq+3
ONCHW/D+f/34Ulpl9xW4YZSlzrLOADRxsioMFIgg50e8JB6Hrf9W0eGgw2y+UvQs
OXRoFA8b/or4Cy7YY+9U2WRSBbBNj99LTW25XZQO3XOoJCtAhwrtf8KY2ysDKTXY
+1VyK2ZopvtOdnwOV5rskyX3WPS/sVg7H2s3R8IikRcO6+2cGpyFg1BgkMmulReO
rbI28s3PH7JUyX3Ox/NVwQFyRKiWpif0oSKGAzCyKnZAjjsNREDp54pg0tljDZh1
jduJtYCrLcMiek2ck6FGAwYM1wZ4usWkFVBWKtmZD6OStB7pLyHG82MKUvvTfeRA
AG+rA/A+3powYA6BdifPMdpCtRXLekwL8qIIygA76yvRqCfrbjAxhwDTs9JAKzrJ
1taY5gVFrAAOWX8M4b547qObCtejvTGf6VWbzxaPpp7us0vuQFwj2ur2rJOidc6u
xUMw+yBq4ZWj2gKEnQDFvw/3KrNwhR2rtPRkhL/GJSGQD8LkhQiYOVy0M7cK0pTZ
10bt5kleJdapdPPR2/6WF3COZjknRKzD7MkPWIn09DOBqa1AeNoYH/qxc87OshzQ
5JmYn1MceNMxcX9KNHJdvoagT5SNIx42ugoXFkoRPwqmFtMKoQU7AhMLO6biBxY9
47s8lCJlu9h7zwjct4Evm19gLnSSjkzDXfAVycAFPWop6lHIkrO1ooLp2K8G1GW8
YXwPXIVUSJejOqwlU4RcmrfAWL+AmdWI60WofQXJa8JNfwvV5flQE8ODF4z/M5DY
toKYbi8saoGNKhPIMqqJnNfUBmV3DUgOeyd5RKEiAWjl5uuEOSaO6Z/4yIP6LpmE
/LTZrAxfZ80qyPq1Iywj/onDXBmkNzv3UzIxYpXVRv3ybD5VE31pScH4iGQM3tz4
9jEexs+pKGS4Oc/yjB0tRGIbVp2FgG3+Wcr1LmyjUUpa8XmWAHBfSCQMAfhAayoi
XU47hpMba4c361DL2pTwNWskoGZdnbcW5Pfcw832ixHJQx4bMmtS/IfEfgYhyxU4
+wZ6pf7oZVgt6ht2lcL+7g8967izmXSkDux4Ko3niCrl5mDlk1jcAw5qXUKYtbqA
I0SrD2wlaXaKAahmU7GCKgr6Cv36KfqwNtGC0E8kJq9hIZQuoKOm7LDadVa+j4Gk
FRYpUNlb7GZuOpCgBJLHYjBrJfbx8tgWcpPM04/DZ9kj4o+kP4iyS8ildePRFb8v
ehCbeyOWt0sbiJcOIs6/r/HrvOWUMP7cyxJDaYR9c1mvwZKqPlQwyfJpzXAuvsTt
PoZ3W04uAREQJ5csgVKafExgf/fJFvZUgyB7ksPxoUuy3FRn4cmMOaPhsfMEOW3Z
8wKv1DuTU7iiBG0wKVbZv/aPr1Q4XT+eZVjLpRaV0rK8bEXqo/pprD3IjlDsfiIw
PhKieauOLstg6UbG74AeBpT+rS/qOsg97AnP7BWTLSZTeeH7dFbqBpbaDfIqEzdg
XkwhFGZNcNfXRJJ3UhYavKZUKjJwPTk7rt2tn6i9jk/RIepOrJ1Dy3btBMjZqYMF
XFJb4HZ9TAnARxQLgFdJlgenm1vhiAqg4ScXW0xcCzSuBYTxrLeUwxgNKJ/AmtkA
AQ4bmpxIE3Kg39nyid2zx1gogcVaWTc6UVaVnUqmAbcWopLDTX2+xIdJoxmpthwI
CIMynDR18lrE8SVdUgXW6vgqbpd08pwocC47OJcfQz9T6K3O8tAbZZjXQ8TC11yD
u++Jp8Tj+oqIll/lKlD2hexcFmCXevFs2tr57eYkqRGu2qmXalAFlnJb4OJqB4Nm
WSCFEeHOOZI0qAOyNf0P9tczFycw1oNyoEFXWsXbl7Q3wrKbwcuZYefoQbeArdM/
P9anpCIq074zzdvX9kryxzTR8YjRgBSL7jJuOUdH6fCyfJFLmZiJHqTG4jgOf0DN
KbGXKkaykNlEdaigFk+uIOcPOPK8aLKdBu2ekCNiYdyvNpj8Jcm+lCb7dt8bRFOQ
IgDNEnxhpKZT6I38w1r2MnvGl6mxux4gLE/YHg44dSEqf9CgLwG18vj/ovYXlhVE
thgSpUyJpUJDOf78713ub+pkZ1/eyPv4AwPanp9DZomgO4L/OoER1VGkt9I3bfIX
+W9/t2h9abpqMTQMjfLX4wl6722aYEliDk/Iad+ovMF8hNtomphjw7HW/209Skoj
RNjYl64mziNqJl60yZ945tFLIc0enDTioBCgMjPOOyw2RbzR/qhHcxi5ePh6zMnO
I8AlIKF/BcDKMgUR8lPBQbf7OxIF6Bnf5zCg9c8uE8kmg6SnNSmCrQAfGv3+O/E9
uuZRHWbLF7fCBZpGmtrCIpGnTlKHAf2eVGwVb+AKvT/KQ39z/QNSpHTendbUuIAu
Noj5G1PIcsb5Hdv5KCG00TpthD1MmFFAFT6CaF/3AKY7sTIlkfHYCdFfCt2tjkk2
ro+zXHMit1DXUiGX4VQ3YkKHj/ZSSTdtJtrZ4CzZhkyB1u2OVvpMufNd/IP4AcBU
NvZPuXG2YvHZWu3eSEJq4cksctbBsd43ny6vYbv0oE+Bwti3UERTBTY30OAb/bNw
1qeCZtPYUxY80hOwaHKVmOWlG1JELYC7BQM9Yik6z3afoSBdInNd3iPbMlc3eMs5
duAxzLaeaa/ZChW70f+QaCfuKtmwQ6xwIt0IfNmtWhbVzGz/idB2VL+tsJuVIjar
bUwtzREHK4mBxWV0SDNjpP4oXQimoghlsg/z2U6UY1OOIPjSYagSmxi6JmSDfOTQ
0wdDyqCckpCIWhcpmVM4K6b592/jy28Ko9zE0zmjKys2c5xkOj5mgBcJzwxOQ5cq
xqVzPYUTwVOeC+0/JUZ5sRWnjdhbbgqT+cBc3r+qLcCgZwTjT1YGYd6L6xmGh0+0
kZI+RQJ5wTXvyaUtS2D/6VAj2WmCwAJRvnKqDdl2Mt5bjdXcWJqp4mZIpiBPMMCg
2sIVjZMkny3PxYF9OzJRBsJ+p8YvFtDPd6sMBT4EiFM7WPfBAe8RI8re2GMDzjPt
weHlYfSqdsjKevtDOjNT0hkG47lC5tH5SPPMFOGIUGIFoeoCfst48N9v+mx5PWrs
cNjCi3DD2a7exUyb52meZIizWgqooKr4MOTnp1FwEeSY6toF0QOGa0Y1m2SLQzHr
dXTlMCwDImBelsLXlrdN44libCdP92VCQRl67pjIeCpIriCseTWmbZ14RpFrgG6u
46H+oqA5CDwjjgqKmkINZjUAx36HCKOj6lkDdp8qDF9nklnomuf9q7wH1iIv864s
rzSicTF1UMuGhhH2ndhMJdaEYHOuIt9UwY5VyeeNTfO8JwoU0TcN6MMY5b0yjeCk
wOMkLBgzZJIgmgvyWXkl8ZoFwnKorE3lNO0/1DdOcG7slYdyI0aBLfhwSlDWrxc6
xFwGlS3JDAzn9rOxtzuU9G/XDHgixR3bK8f5aHqqEZq0MmPdfTD9ps5lp9WR5+4k
h/lSSffzY3jVkGEaRnnd2Lhu1C6cn69HpmlQ6i20z3KtTbRiOfTWUaUOKLjsZolF
djmzrNwAg8bVqHSd4K/H8lLJH6im/3RAk86Xff9vW9rB8LnhA9GYI9LLh0oJmZec
ZO+FYUGRVOn8J7Jy/z7/7UwJka3y87xKJOl88c1Rj2NaH4roCQbP2ifmi/CG55g1
N/BJBB2SEqY6aXwSjBgsSnspKy39BK77ZjGnXB6jsulcW0zn7fy/4nopM/ddTpIJ
LoF+Nzu7cSXNjyVmzg4mIsWaOWgQcOMewiC1NWKzN2YiQ3P94NkGs6WHVebokjLI
ktV1S/JX4yXjSAE7sFAgRvZlkd7x9mo8mlE/N22ktwJKbKGFmJFu82NjY3MfEsrH
3Dqv3W60kx5s7QDExwEYAf5qRP/52ToQwO2Cq4iVMa+B9E6JGi1VLQvLv4ulzx8F
bZUbY4WV1hYBwQlrMNjy8AfysjNGolOPARGJcvf0E8UzjJVK6ppskJKi+J8V/Ctl
yZYdHM87qVOihrEoSf5/vE2+9bkXToyyfG8unp/oF3cgzvm4lTXcbmIVp1boHpwE
HIVoUbOg5TKSV80OSann1lkzji8Pms9ZGWY+zciUb6W55gFvJUaeyVxFiDWFGLok
iCfZJ2FYoBOGag2pdiQfia0HV42Hs3CvkGaeSVr5txMb/C3OFpOcbJbYQpfdHiCe
mPWxOMCtihoHIUaPmK6drYco4QE2b6g5MfyIWJXR85VbWASHdVM3fKwYG+oGseHi
qdahDwlmQym7rXmN7vsFBDuPcNJLNtGsZVcfGdgR8OZ1e6BT1bu8N0iHAclLv5rp
6zsn4aDYVh+n/ns7Oc8foC4muDQ5aKNovYqDQFN+JV6LXCLWJB+S12CHqy4wXOoS
5dZmg4odkWNxl1AMu+f/Hw1yg58BplJwyR2ivsnhVoAV1QfIulZysVnh5D16c6nK
HWHtX5AEJU7XWmPwU1QGk9EU0RZNhOFl7Keyg6blo5C1E8QSPGcuCLWn06Q8MYXI
ldZ8XUBWMCHdMd/68hcHyEgdOPCwJ96Kn5KYoATHkKIyHze47AcY6CmZ3lhwt8Uq
G3XirFtqNhr4Kpx+Ba4FbI3ed9d7wjmZI1HBFCEwAr8633jKFLlaKZY+x0kdwXpi
RRswuzuomPVCSIIskhWQT7T6PC6qRjy/G9du9QLimpCZt9MX+b2EfK3d8fITWVSz
a9TvnPy8UZgoirKWSdJTbdBM3x8kDJpTROlm9aWYphSeiFk8Ji3WsVokxMDTEAta
AfD7VyIEltnRxhqTfPoCfi4Vqzi4AUvtSCcQrUOj3PeU/qFxtnRczIxHLV3rfbSD
XWVDIpwmy/0TUizThbuT2le7nyTO6otPlJ9zcgnAmlw9mcJKN9zwciECkxOOMzA0
vV5lQbX26DAjGuBQQAC+LA9upgGa3Zct/VlCrGTXEUBxujRSfKix141HGN/aC/wT
XlHFdVRb8Eu+MVYA759E/QMmUJ3zceV3SYWGwb8cqdm8EAyaFJsgsilYhf9dVNMN
OXLJ8TcUZ3oQndUtC72VryYIYWD0a4agBCLqFyLKNAwhnOJT7JcWiKAv2K7yJf3F
sFFpIEHAFb4pjrWNNhZDFgw3/9OrkyL3+DoMM30rg/SsfFL7azyL2UUK/5sNqrX5
1+GSw/9i3QzTXwefC4xhpCoiqhP/AE19N7JpEHcOtuR6a9YUlIOkgFk/Yj4oeyoq
KHZGAA7rci5lSWhFOKHoDs0SnCx+LJXuJrln0WSsa50TagxDAHLGVNo+N+zpJHg3
RuPyNcSF+ET4yRwerOdVv3QN5luducAM510sZHzg7jV5KF7CpPZ2QCJXn6kmWOCB
SgbfuEVWhuyV0ZCFmb4KvNeJXWLq4bLurA8VQi8xiegk2pQrRhTxtkKXTIJ3JjxT
8SVpohP9K31xLGmd2W6ujVooOvO0hy9h+nKGHbj5qax5Cry1hjqRIAAiPwpIA2uR
YOmwnm+V627f95oDgOa5lRYHfiARdfidovqXNJn3CR1pX6jPfme/mP7hDsz1q7Zx
6hbbu52TXUP2kLr8E8NIGGJxJEiJHfEFkAkA0hWcYK1uJLrr+ZorRACpgL++kXzU
14cItqxsnHG0uw7DprVfakIbku/4cOFc9vVBm7jB3h1Rk417nLS1gMBcPTkl2lQ2
3TsG+yKJI78DEYVJeEhsNjfcwfDFz08aiUKZdNeIMvDewoMGXAI92CdP5630rmQZ
SMI1j56IZu9uaoKEFlkS92jsUht6hu8Mo0GfyV6PRUUI4OsZXVUiKdigjautr68j
7B8hi+7sGOSTV1VZWXyTl6erC300wqIfh11gzls43ytkCj1s+T7AVyR3xWMtc1R+
/QVLGnHv+rkdbJL8TUj3P3TS7p+VG/xqD7VUEJAClJjMcbO9KWuVmRwVs4Dec0I7
dGei5CwDzl9QiIV8z30H1aY/jlaiNYpllw2ToB+WP6Omy0qJNDySySiE1QGRDbks
KOkZfnPxNMaz8KF9Y9zdKRYpKQrRj/8VpMzUbfC4RLsQf1QM7SzTnhW3xHZaESJ1
AnMybW+24Zy0N9RhS+TxCVE2kDvEiUev79DznPt485IQPB8RTVhj+noutgox0mNk
/GYWrSxytG3V5HyuyE4sGlDFUMib4emw2I+j4XUcqb9B1K5Rw4lyrQeaZ0EEdRUJ
M7TZ1Uw8KKUiMPrl4kGkV0e2eNl5ggUsrOo6cHxuueuwE5LAk2R+tP85L6Q395/1
PZE6TbUHd6Z66uvauJ+Ut8pSzb9DNAu1nHP7iZhlUGd45BEXNcOa028eRW0ld61D
wjcEFbGzVVbtUMWppOe4Fkx6LBCNF7ED8byLrMedx7o9+ObBbI4+HJsvBEe0flil
EPpqHFTdVdpeH0Lpmtw6vlduVgi79LOtHzpiWQgPj1L2pexkvh1ozDj1ol3uJLfh
zD9LOTvzgoOAaqR/9owTSCklii8mAp/0glt3Wogub8jqQDrg1e/4ycO/uWpiGQzw
NKXSTaxfgxANZg0WhIdxAXSLj7Ih3dGUJC2Mq/qqNzBihMLEm+FDoBOnOq9RwL1j
WcIP7Kdp9BnxxbMBHk2K/J/Sj7JMn2/WNdiFJ3QFIARu3bE12EE4ehyISU1dl0ud
r0D6belAqHaShxEZTmBp5kzK8Qqi1af/d1xuBKCgtGD7xRMiUHJKgyMYy38h7CtR
fCXrF1lR26doFGoqPH5JjCzVrXx6AK3ivoFwVK/4TvVsOh6qMoctKd26FKH4hNvH
Q8j1NWIHAsT7o3aLU098rxL8WrgUPo4HQghSUiyrqUG73fV1TZKV2mfLy4JLOq1V
CCYWak/5ioCu/Oc/DmJ3wNIMdJ1oaHk/u0c2lpSOkBVMvZ96nPJiLL/aroVjAJVB
z+J9O0fAJGQl0KjWBMzAvKgLe60OcsXMGNC2VbPWd11Ymnb4o42nhJi3Yf0XtWWj
x5xv++0PAjpV7TfyNW1po/3jYyIoUxQQECruBDTqz+LHxZiKTGqPzLnKvp9iCE6J
If7Tk+LdS1NRmWcMQfU9Xt7YQ2RfoFMT3NHx+PAobHCQeWD36MXOCRQV502WJZ8l
UIy7/OVyY59t4CfffCscETgYDegd3N8hICBA9d2CKVuTN6MQJtAqOrw0X1DN6xhm
WJaP7R995jy4io1sGdonMYI1Qco9e5QkzwuPHdB9q6fVUViYjCrsiuw/DrMyLkk0
asoYN7TT/5YXhDcXkKnwZYmtVwG1eGlMj8WjuEwyv0Eefx3kdDTrqgNDJrpZugGg
Ke+rPMdk7FZWrrA9+IKvdAaFUgcpdkIJpGJi24tdxCMttMfPig8/rLdSAVCU7hU8
1WE/1IbPbnoMwupGcNeMe7XTBZ56Xr0ldkKh6SsJ8aq8tX0wMETuTSCaBjy7kBAL
+RgWeDTCm4MuHTtboy/W3r+JXJLDL64xFxc5bOVU41nFYhiMVaExDuhSKSSAsRk5
3w7t9HyFlH/00aHjs9/A/k8WZHwvsE1NPUAnZGz3DscIiYJl1+I4MApoVZNRTPVn
oj5mYyvcoQAwgt9EZS546tHTBLk95TaBIYqdTGrTt00TPoe+ov7NA18o8b/KJwyw
uHLKcMvqz8TlqpBviJNJIHH0vxPDZFlIJjkazLAxOJ05Li71YaWxF/KJTEQjJqnC
IomIWmPdOr7Uj5iKdsqa7GW+4Eha1Reb4lrQluGWoJknmTR+vGQ8rV9eVs4FFgKK
O+BT3N4xBoo4Yl6sOv2Jq8Zi019eIJr0DrtaLeRtawewvRJiiqP/bIm5GnuQwmRE
rgCVUzfw3ytKylsfmBcCDMr6XSMvFRttulJNEfcgkuZTREpwXZVNwFgyjKbQ81zO
FjQJPrzfifLITkdevteDAlrpa0kXkgxb4ecKjPEeCytShtfueQ0CipPtCP8+Pn3F
0rwyRVojFwiSKE0efZvQ1In2i2MUBFDTurQizZkRtayxu9PXx4Ma08tPGp/JB8Dw
uC6MD/tM9RfKEagdYQ6Il3yTUQhsB7COd9TG4Y8BI5Ixk1BgWc8HsRgYDi0YDxuv
P3PLvQFZvHJNzmIY96wMdVpr5VaXtqzOI68gZEfZDRZR2wcB5KwoD3JmGNWiLkDt
UfpdfrnSJM6jXigMtCtG41NDpO3yc715jzZiV21UQjikgZeystNf3u9H4esylIMe
pC/Bd1JytWQPpqtQZsHQxHjncZ+qSsYX6a1OQq9UXEbBGIRIn/3hlUJxAwipaTf2
JH73pT+k96wJNuIsF/yiWRy2s6dyc7nz6+vQIIg/Y1BX0FEpMJYwXujbXgjHGP4S
8QHHebeSrVbukXY6vUnohY/ZFQQdjnLLZgxsWgeWS5L6iVokhzm/7C3lwa3wyb3A
no8rY8e/KPuIqh6KzUmiSGQlAZJ17jPijDoZU3r1iaGCGajJodj9BDUr1J+7sEzt
A84GpeP5dOD5YqL3CIyjCnO3zGQD0KGVpiIZeKmygkTbo4J3btUz5ZYS/FC53I78
wQnObelsV6h6JP6IoPk9gs8CPCnkFORL7IqSGYahBn36Cz2dr/SGK3lcWU61eQE5
HFaKFEZo4qLW0gv+wCYYfKaDqAlgjGDR34Xcb2lrVYbY3aYfCKXj6ODWqEbV40cq
QXDC4WG1J/FsjuA1ILiAk8gWDUbu0njWwJvFUdlVHQWFnFFKvh8x49xnB7j4giTt
zwEKOuAl9JuWZENoObZ0Re72eEuLPcPz0xDigaYJ7yRxF+1MK9KuprcCYSM36hPP
t8L76hm2Ib10TywT5na/5JCbduK2WpwLn3wiqwqrx+rSkz3QG803FEfqxKdnKEp1
AydIeAktJhpKFL3ypfJRtcG4N2jgASM4P1HThqgdJUgOoGqeev+fJIGdOe0xOavD
/f5I5rfHO8m0oHQjY7DLei29QhjDD6sQ25ydpQ/RVT0mdivODvMXtkH+gL8VnkP6
vy59N3mC2Ir+CBRGYHr81ccM0uzt5IXs1e1osERV/cUwX665HPOnKgj3Wqvk05u+
sgYGmlIFNU8U8xiNTx2SEfLTISRf+DkO36RJGH6I+1ksVoE5bIoOWAXsaXesLf1d
kdxZQWPfnXqyz3fNZBFvYG4ZlddApvbyiZVJNNerp7xaou6Is/1vZ5+74B8FKnzo
w+NEiiOBx9S1gNpHmCnhjvvcKjEzthOu38G/tKijgdHa/wxtu9vRI0nQ3FEDpIR8
WFyMBFIp3gPqzt6bb1oVmSup7W72t8RPv6pPDosT6cS7M7mU6dp8MHR9+1I8Sz10
6e8RxRpWTmsbiTAmUrP6OtXb5KthdSNM4A2YNaLhCxxehBJZ2CO/wS2Qzy4yPyRe
4Fc+bXd74pQhJq+BMUhTfqDa63B44VkWX1pvybaUldY+aVHELgmRlfSOgMCEyeIO
Jh1J1X3C1+vLXBTa8GKoOZ41/D2MPz+955+4epsicdbCEB091XlOf7FOnm8v4r9A
eoeIwNH+vCEuUA/kxI0d50YzmXv1iCP+jwLgCA9eSs1GXG2/AGkzRiXXKDM8fdGQ
0gyG/VtLpMlA2q4hXlT7iNMKvULIYlOAk3dPB+mJbyGoh46S5sO7jlNKLiewDKSS
eea8sToz4AUSqgJkuyje1YrVwdTRZ7r2LwXFhSRvPBJ04PxG1IqtDIwwpf2sKTmT
RmihFZjCl3o1KLHj0taxD2kDrVmWmAZ3MXSmWE4EbBAatmL0D3ZTZeEeM+Sdjjvq
qP0ELLnMEKopsPo46BixEe8kpRcRyOhPiNn1Lgxgzf2clEL6BgltObduU8rHhO9h
G0WnZZF3po7GmNi8CI50pDAKMFr84+zgAhDHhI2+Sf/qMVlJQ+OP3DYOb323LYDi
nXO5XTnBjPulEKtj+h8QBTruOBbB0bZZHWwbQNHPnYNax15Ea2SWmEICbqFvC/0P
22tjS0dRUSfl4EIrjTSva0k2CllIlqdJMjf1UwoKrkpXTNKoGiFCmK8DfqthAOHT
gS1/sA6ZgwvF+7udzHZj6X01LLCkTctVRStO4EZCcRCkZ25bQk8wsf/vU0Vr8Yju
QZ1yDKAKYR4GuDTsjY8AVvC8VSWqV45onXc6sj6QVonyjdPeL6W+FeSOS6BPCNRy
WuTlYHbNbsZZNo+5nEAODP3H8COKonJVN6QyAQAoB5PMe/XXSDUzijl9BXz4mGQT
6/EMcUoU0fPLvDw4Z7LxNijPo6c8J+fPudrhkt4MT6jKZUSdU0u6oV4aVqacnf3F
82kS1kP4vNBgkvCGaj2kWqGTk61GOG/I8EGsJMfDEmwt7N+gw6ecTDdoXu9HkB1R
tpXI7iLuTZlSo3xYo+CiA8fgabn2grAdK3T4a593OoOTbt8xq2A05lzsb1gAFl/T
y/u788Ks1k9IgKJ/ui11eMXTQn5uRWppsNFexHkQUtmjJIUHD9rLKw/PaAGM99G5
76j0zunmw3VY7ckXSr4xHfdWYFO3wS2a0vF1O3eT3uEwPV9qBCNxk2PD+TEDqkMH
ZzClEAEoYtkOzwaIyINwHnv2bJJ7kdGIRZhS20yv1hQP5oGN1K7T979CIaG+QRqq
w+W18/adLZmKMJ8pUQXHuvdLFqsZA41mWmrx6cQo/WCCI6osU8VZdV4loubiHroE
jMb7nsDzlJxzhQF1iQHdVdclWfMRmuJKyvy1PyZhPo6ZB3V2KImHrVyg/rIbIR5s
V9p/+taKHWZtXXbjYsJ9+9/tBzO7Z/Qd0XlVvuR9H1XH0dj3LvcAn0ncTiK5v9gV
iqmpfrHfnOZRelUngNvgasqO++hZsLu4VOTZf/aHjJdAhelpmdBVAAdjjs8spltW
F+nBubQ4wzPaaETirZ3GGxXomtsiVCge81VoaGCpsxGW1ldbeCJdOFXJXQtX1S45
MYKrK5tfuYeDKWtREFOoyCLK6lv+8lAgfsstAa+vsUcWkHC/PkzDnlPJaQCb18gF
uLkUlk5RJiwi6S/glw1UBSNr+F4y6qtQ61nQlS9YdxPefCqUVXRVUHXqgPpw8vQU
e8PHLz72g3pj7YQXZg839JLfPpgS2Yy2bU7fUdLIOAT+074DcgdG2ZkWuZnZJ6pZ
5JK1lA861/fPw7OO6Bo+CVgqV+V+bh7t99FpapvGPLPHr3/e+EHmFvLvJwJeCP+z
Jo8Ph2UTsaDgMEanZB0Jl1HBN6fR17CwpwtxW5bPehxi9Y+Arm4a6BiNSP79LiZ/
5R8rYW09goc2mKHdSv5B0hp4xMhowsFnrhO2nyzwZw9ryzOVDvGFtTzJCA4XrYCQ
SS3o0JCVr7SjUQjzyrsV1Vntl6prVceUectzGbSLBnyuRnrZXCUYqie0cAhCGvgX
iYhTYgHz1XJqKOz2T5LjDDkZcSOqMJxHE4U9EoUNibrd5RafVBcG0WQY5adzwgIP
MRL1z/fklvRGycXp0RimC9eVzv/zDlmJ8dBUL/T4pzfikAcZqzCvs153hjTVTJrS
46vvx4vIY5iO5D2tcapbBj179mDIucmva9x1XxnNDHcLGL1Chx5hHla/8Qx1fLTe
P5HsgdrcOcJRreMCYeV9UwVtnbKFz77QOQqzw+HoROhHpZzXNRJHVHC7F6xd+gxq
lxyYd3dPV+Q7g6gwoVm6F0W7DQsxAaqIXoZWIkGmZ16es33527HT3WnEROixVNwA
lFLHunUO/sYMZyXte9FHfU9VL9MnENHLE8i4sPWYWHCWOsMZH14qQqsXOrTRCrcj
qViLoF/CJR9Ey34EM5d9h48UfWQTR3J1H0K4VgbB2zEcT/h4RCqxmsXM48nfM2bQ
M+oYdZSPC7nHONh0fgXYWsJwcd2ehfGGzvodJFfTon4bT1OxseT08o8QTBX8YupA
sDe5/G26bbkMX5JuW47OKDQ0xGAvI4KLVmN85+Hym5VluH33yjzqfrEnnieocorP
U48pg7uGhC+qTCSlM5luFOQfI43bjf+Pm1jkbB6xj22pDFvxdU/5RDIlzRJFSWpX
qS11iYLIthWs79nwZ5Pjx3t4kBOlSB7GhSYEjtL7cxsG2nCAt3xQPhRt70E6pr3O
y/YbHhbOGMWXlWYRxvHa7WgDv8cxuAJuwf+BVurKmh61EuhSnm+LHO61l0TkiMaX
Yro5K0/9JEt+OFGCD4PjpJ9amTy4bSkjxmGZQHejWGh1xlQqS7yBscHFcJ9+jvYS
n44aKHMVc3zsPSsWPc3wgDD3T4Y38gJ8mUv89GnWi7jO2dYutv1ZSARaY96fLMxh
il5dXE6t4fg++/TIvqvuOR1+8P2ATkfUKNghQi78kx7lDl1Wh7++0+vjHXsWCEYX
Ud3Lohd/6EuUoRv2lPh6Ns27eEqv3XExFVZsjN9pRj9wIhCsm7lv5SIgL7jl9g8i
YhLa7+OK4xal9v8tcrEEDmrwxr5RlCBJGENePdL61LQP3N7yJE8iMMq8b9lQBnII
XQMCS6dau/4k+S0Krr3vUw3Z2Ex9VqWD+f+ZzT6JyffIHjCI5je1/JSuLfXE3NJ7
vmPhBEcjkwGRzNxGXFXAOzq+CvdQjh2Z6MmgchEZTcfcBMNL2CwSxcgLm3krzR0I
II3A+JN4gdYOrOk6I/p/dXhjjFkM0gZ954WG4dZJ52cXicyov08ml0pKu7zImoM/
q+hMsVsqhWjOdeXnRif3WS/qq42Dj0KPlSfiLwYMfFwgZHxXozrK/7oRopRHoNCQ
M8jPPP1SF03n6FP2rWGqZafpp1l6jXSrP3biq/kkpKzcfPYrGmYDfHh6HwTDPdBs
ObXqkVePa7TNB0ErO7Sr5bOjVXHN8DGjvLgpLbBGdiIAdL/6i8RAtcnW3wM2z3O1
bbNEn9elJo9nXbEUpcgv1g/+OPZiRL8xayxccjFv0aGpHZiiMTPq1WIOozoa6Nkf
MGXlRpdVyladxMl55oNPBYT7pA3/Oyr2vtV3HBRfiv8aoplx9Aq/JuOeS0aHPsZ3
fHpNRbzjolq8vM3XVpg54L8pyvIDExaU+2fsggqxrFaNmHFehNphIakFgiVyDwsC
Be71zBcjnOzXxA0XxIUCqJdq4lw8+z/XJcjiu62/oGzr66VkjXBkoIij3eaX8XyO
cvvnvWqr8pn1fxXXsICtBvFaYdWzIIAEDjd8iKusoKkhFcWc57qUA77AWwwlUVl+
sxRZf1nU3W/joE/pgyC8gPzyEXGZNjQHQc7suCIEjXQubD8suow0/J6UJBAhhK/5
uofczDoHv9om/xWbzjqsRHgegG2IU7uzO0JZ66BA40YP8n4e6qPUm1+LQfBQpUSN
jcOSv9nQ++QVTSC0o8ZJnxR/npYCcwgQLH4ILFM9Xd6zYAYjFH5VTaRh6gucLPh1
pYUywhap5mN5hrNLi10gGcHsmaiHJj4Qx/4C9saYr99K44IBqwWIt39DmX3arsEJ
lhDzm8ZYdTI1a/tNFXgnCiE1hmdIIVagRLVNPuCeFYf5Zu2zoo/zhrtcz+owxiJ3
bfglX/EgBk2JPVv2U1mb9HxYCryzJjwCmoS4yXtASaFU39XPTzhHhRwx3VtyA5TP
jIw3cMSc31+jyWnltYeRfJpcYFZhNC8iezR5IhP+Cxbw+Oe9m4VFSUAP4ckQw5I7
y+Tdu8b8b87fds8Ei/9AegvhRKv5fhwivEFg9Anqpr5SqQnA02p7lLz/KmXNRNtQ
5Q9Wh3BMx04klA2Hn6ot86KUX0ymVg/NDvv5W8FaQN4RapgmKXfGY0Jafe50o0iB
uuZiDteKRjy8CQZPRTSurqWCH7KjUUPNmReG6G/Gd3ny1m/0A4bBvFwlvgy8Pvkc
LTyCVGGX5d4MzdcaISgtAOoJBVXggI4UMPAm0Y1KMRrsyfVfuACCCvCQP/yBdvNg
knc9xetRjvQryYh8IdzahCLmyPK4kNI4e1N4yMxO4OyR8gS3Mova20KUQxifEJen
0QsD6YQCcIdXuOzGYFRJ5b5S+VYUkiD6iTEx/Gi3HNJ/Ubdj4ksI8DfPtMMxXvzH
WM4SLN/4qiTSngcP0T53a3oca3OT6tV392td00Gwq0Ykewid4YC0w5McHzCEmgcA
W2Nw1g2sdmaKMbTyy8gLckbqdksTfa1cPIoExq4FwmMBV6Z///mXpxb9GruhRmeR
Sla4D8KoCFRMtxNytKrNAaEOE4JqpvcBdqkZ+tzWX68phVGMwoDGNEwC7QeXuYvJ
neO5Nu6NJfb0wBhYQDS6X1thi/RV0oIHiM4GgxSY7SLI7nQDfUiAkbwXzZOoqpZA
LK/GxCeu4whCRCBUHFTzDckMR8yuv26m03CkMJno7WIF2ChmLBQGWL03p5vw6KSN
yKOgSPpPD96oVe2edOfTrmeorRNGHW75zKln5aHl25TnCC+yJYvCGw3GC26zyK+/
IYSVc0+eS9OfwdGoE38iosklezpH46MXMANfmLqrO0QXJ+4gVatkbKJB9Uhyy/Hn
/mCFd5vL1t43aTClRHjhJOP7yuO/g33m0WkaltdLvS0gWIAZaIVtFcotDGZAxIdR
pxsJvF/4kUC6JwGUV0UdpEkU6UkD2lNPJ8wo6nw5SV67HfROW0dyKFah7pa/chSc
CD1v7I7GvEBvweOTkeCb8po24Yj3w9AO243VhyzpzQNPu5H9ytbPTv0kLfItAemb
FKvopbg4GMoPqQaLWniDLgvRR7TN01QHPmG2pUhujV0uqoT966KCwacW5dIolPTQ
3EA8jGqXfDXVOu/Ep3o22flIjx5Xjn4a7d0FQ1w2cuUUIxyUuXREYb5EHFvM1yZ/
ay3mOHgcRWG00KPETBuQ/UPdp7QJpYcjyA7Q1LFUq1/OKRZxva330zWtbTmt4eI0
2BoqbZXPNgpjvLrR69iD3WiDetJMf0ERnq3Xln+oRrQTS9iAHTR58oTAvxlOWssA
KeYyzRhg3Wgr1LtmkGQufKLiLkhDdiwt/YFqToRQLps9xTOekKPInypcctYfUSIV
d6kaikqvCfaVlyXXq+3Eqsz8QICTbzmqSM+RmZVyiE6+kTXVcv/H+6rqL2CZx14X
H15X20+AqMynAjve+8djVF9cIcoBru7s/G1UmePQTuhTD+soc+B51dH+WmdI3uos
EGOg1co1M58812Wfroyk9DLGIMSTWzTlYYK69qYKbcj+TVxnb+vBh2YhR2gRaqil
NXtJIIcp0PQyGmwKJxlLq/W5xlGCWhtUTiIlt0KbaTWoZgi8jNALfQrApgkVhfQ+
B4Pk41ouUGDMZYsxHcR2myVTnJfGTlTFbo/su3XFBltsXdK4s+yrftk18W5Iebtt
6ymlDuFLH7PtVk/ryqYxlGWCBLIljGC9EUTAtfSOcbtM4Si80RT8GDXeTzpmjcZ/
nsDr2dUx0uE31jWiB9MYIG88Rdvmfxr1Q+LLZoR+lBUpZBptvV1aSyoaYiku0C2c
ULs5WLANO9iFKpBV9C2SenY2bleLsnWL/6MJAT4mxy5h8XpAqCdSwIlQCmlBSlbu
yqQxdvo713tVJSeDy2gSYp641WnuSlYi9dYEms5478nMcyAh20h0YABus15aJnRq
MnexGiHjMRB9Wrf4cQv+7FJ3cG7fMpU3B7LFo7ZGBCx6xu79XujzjuRnXx1patf7
068SoZSwoO/LfMQPMXyPb0qZDPXIuyJ0gPINKx9rmCvkcLiFo+323akZp56HhpRX
DTIBsajBaKgliZRvPudyU15Nn5hOSeKd0jiGMUgkkzQ+NrAzB336bT+tAVdZomE1
Im+lj33b+vAOypqpPNO39TUCnzZqACRvzcU8vwolfPC+WUIwYm5zGpgVB+s5Hg3x
kDEgquz37J8LZY4U1g45B92S2enlMDuad9EuLZusW7nQrOZTJDl/RhAPFfxtE3ER
23qxcg+r9w00ErGAvGCQtzWnyBea+aU0olWNLCw9wZXnuwja6RxKbo+fGo2Ukxv6
48zVnDJNXBgioFD86aDkUxru8A1RmPjrYjWrVy6xf+90o29xPuyLZD4pHzRWzprd
6ZCCg9pYygJrsSnDIP/Ca+xB8aFlm3oE2fFSyyHn+Ka6EFUH+QF2dj0MltdgScx2
peAEChZrkvDjW4t6i0Ie3hjRa+hiz03ZKI0B7O0MyAx7OQQSpctNHzXnZYujZc2K
MydkMxT8aztJ4b8fL/7DzAUqvrVj9Pz6WcL0g1zBsRfcS+2Bv+X3/gjXJYHODPrp
VrEfvrud8dgoxzzu5y1WO9EcF8eE6/YcKEuf5kSa/xYDLink3qkNXM23Vs9sZRHj
IIWRwSJJ6U/42J2TIF8fyDpJKZ/4bL2tJJmPRC71n4XK4T6rFKNf/ftHkahF72wR
6ak1l00Che+wB5yq2jtiWxYemFqT0PMgs8DLOic7MiIWN9GxH5m0BpOjB5BazHRa
tqM8Ym/R4E9RL23ZwLxoUbtsEfW8ggriBV81/J7g4W+O0rzZZVZko56VYfXLgWCv
felWFJksWR+w4YCMjqSwUHB7lyMtW1P6iCZnPmj6VcjrlQ3a7opITyUKJp0mbmty
UsgjGg2JbWELSzBlp+aGUQcZZ1QftcrNRnctWIf8VoruG/7sr9ObfnKz/ktL5DWM
j720Nh0N4NRKX51HfCLJaQKC+QDJjdTuc/dHSid0HJyfLsKzRBkXZ10UfB22/1p2
ApOeYLFVbe2tRYSCerHbL4QEYXawVlr2/dbvNTcdAoHguSG7iqj3c4/bBX7PYAS/
8bD1mMeafmdjQKWS7q95CzC8n24b8gYj57GMPU5B7Vn5TWmf4aZIwTDGsVQlQWD1
qJG5hHnP0+mT8KepNKylyGdpYqrGODmiVIWNTdxdyv2afzmCpSEUSkFGUfiI+YTV
4DdDcYnOLdYvgvMSt4BrCPK6AL249s7KfjmZf/FzxdAJmHonarqu6ZGHnDGFZBT/
6adUt1wPvLyLQNntRXiC14mJq+1tpRMcQxxBDhqhIILkWB3EltlaynNtdCGOE7iR
fR5VPWeOgAu2eH7iwwMkpAaaNZ3+RiF6S9TsWFHxseaEtzYhb0yWLjEToIZAIkZV
M/EovorW+qKgxZB8Dri/o//GCUTU9i2v5ajeZoKQLfYEWdgCp8ZjifwO2aKV+Cjq
XTc4lU+KnDLxSJa8+oxe8DNdiWCDyqxKYIg9D63futa5HXTqIff7KIodvfAc34vB
I0lxDl+2orAYS9T56afiD3P40lB++5TGXlHlHyWLWbeHtjsaWxt23WcJdRV/3LbC
GZCrF8hFY90HmdVOAI+mxlf/HXwsbU+uvaYRO098/tCEYoTE131ksX0ElAoPeos3
Ncz2jrCUPa4OnoHKKKuXDe1BaF8lDhGMZJ9nARxXbJtxPKHAkC/nmREUs1mloYdp
X9g6efIyNygYOU++Gmay3ZZG8ljupWk7ycAEf5S5J5wqZmmPFuFHrX2LG1Mdnffq
UMtlrT/oY6oyBx34i6J4aAem9LN/LghOXvVxeVztD0WT/ubacNaOWWXbUjw+S8aP
rlCdgOdrp3EYiNBJOkyXlEn3ktCmrZUeHxhvetzIhxNm8V7OcWCmIv9CqNlpKTUr
XwaEofJCxkjL8s4tnPcR1tXudzPmFiy4Xe2T4m7Yk0gsesIm565cyqYRWrogSXSP
K5Vsy62/OuIItnleLhMRbD3Ha/EK9mL2hvGGaDna8SfEWcxzN9c0HtTtOkcpLykU
d5vZwYuthw+ICxhSNgc4uJT8CdkZmU58RW8ohdKIuH/9DTcnehKk4I0+ZhM7SV2C
iVdgYIDuOn4LTJ84IGqfPRSM5yxXHxrjJb8wh72uaCF2vORk219PySTKz51lN63q
+kSXH4fXhHDG3bxALKvF63gveYZKGITLJJLbOfYx5CoZSQTIb4m9X5YIOppnUCT3
QpvSu1GLPLQVhquE8UyShlF65Aw5gDqLK1LmrfsZ/sWaQFHKE8VyG52VZazCkMGD
hkSzRrWjsevgHwzd8DhWrxl+Oio1dsaVeo6I4z4WwrXnBB2QDooNlJZepshe6vqO
6U7eFZpefXBBKKsDfCde9hZCvffUnBT29TGA5XiUySt58s7whW7IT8RMAY7MZ7Qc
41SrfFsvIse0IkEu5MoGx/Rxggx7XmjXqlZzdNE+vv3cbSORa7JLP9ba9wBsE8Yg
PWRkTilcl/v6BlYfCJG12PE6+McnyEd0CP6tYSVZ4nE6msaVdewpYq2P182547ha
IYQH+4dte55wxfAfDUX/GfLHX2zJO6QKmag4oRlhz+tbl6Mxt3JrS2vnybOCfjyt
MyXMpr2FW9vhA5nG0ZpbrXpAa0BNvxyrYt4nc7HSbv2xiwCvzjubNIblyo2FvxdK
qLwR594oUc9tqukHBocqdJBFyGwBHrWilwN+kYl7gpqbMNB7Zz7gs/ht0BLvYMtP
jWZ/N4n43ajE3e+wLIdzGt3OyJ18MBIja54rqDnDydCv/mk5il5mD0LkvdQrRFOt
ZzzNMtiozOrNsBfXuKBvQUw+WldDb8dpmncaBP8AKuDaZqOkDnbQLJTn8yC7WrzX
NIDp+IjHRL3MjkUMxCX4DOpX3nXvQOTls88WhyYFkU+RXyDxuxJuEqjsDTnlUchQ
sAOWnke0hOcz4rIVMoRhvu2X5SlM70G9MpjdchsI6FbB4SX8tW8Sv7VuqTswbr3O
qEf9kLz8/vea6+GqoyitN3q/XCJgtP2PqMEin6WjIYmXJy6iVqHlbcGzzNQE80Ro
M/XRVgrupXvsNCh6CnCl4/OHv4iSEKnW+k0t/DWanzriT/4xV8scsPp3vzclMNHI
3Hd9yqCYCPLkXoeCThGA8TCUfc0hJPd64HUTkWszXG7En6fSJ9iX+jdlrrH6WJ5X
whupNvKE+PNfxhsyodvDTjyAKzX+DMWS1JzNLA8nHYw8VpOkpfJNjsp5DiYXOPBx
sQrOFxOaZv9onEdtOa51bwbgI8fxxQcT2L5umrHCIgh1Ge3ZUQ04VA55SbpmOZk+
i5kiC9Kqj/pvDtnjSgqMeivmyngxW/K8ifGOn6UeoTeXMwnlqN6N0RjjqgHvaeKW
/axXB6p4r8xZNhHZQoDx3h+UpnqiqQDrLmo29ykVRlF1d/KW7Zpm2C7zNEWUwW0e
kTzJHJlZQqTfBc5ZblPyFhscC8EHeVaMPTXiQfUBju6XJdAgllHYVnIn6XRJNPZ4
PMjWMPoQm/WUMSh2ki9sScQ1gbMVLShHgpGKDMuNio5oJWyrk9hapxlLvbUaBZns
2qojhs/ajCqSIsOwnqep1P/ZPtsaXwv5skeUvr66tFKOEIIi4hnCzyCUDfEAyElB
1cqrbAMLUrXExYORM4e8LKMdMUkHD8gBIUnv83Wp6PszlsQrUxdTMyFMNjrq8kV0
xq9iLLPptDy55nCGOOHfM4rfkqllS1ZYmuVjOZsj2Ab12b/yvfpzrGFVOm/VJe7h
Y9O1FWSq1IB9RfEqa80sniGX4QwwtWKoiUvVx4xrE+zhH19GTyAjQxJY7mYUJJOa
dhgzK+cr8KCdBV5d6/8RMF/qseHFQU324S9JwHQ7dDkSFbs19o3JYWNUyQucyevT
y7uB06ndq5yVqU5/7TpKIqD8TSOBQEnATdrzloLnJXQ84IPQSgvlq4AuOySLY2mM
ViwjEPwKgWIA9kd1jVhJVWjMdZBz++ceq2icImNjBHGN/8u7q2dbNhoAhFRuDeSp
snB9Adww0NvUotYXL5ZIkxBuwyiUcp68Fa57616581ZKWXD0d3pfRyeyUK9fbvmr
bfKRZYRnAkDxiVh+geY3rgGTS+BcbpG8RBUel1JQBV6pt145G7Ov0NnnE1X5/PGf
wkUee+aaeczv+SiZVRI2sKY4UsKAxfm1x7eUpUlYV2ZV35J/zrF+IUI3Yx6oIYhN
kfHdsl2Q0NAu0YWC6VW8ZeJWMfISGvk4rdHu6NhAYMZDyzbcOwKJAMD2P/4dPJPQ
0XiZO7l+Q58uckr1FHOAUGRCEbMkw/PkHZvXCuCS/pNmHW+jh+Le7zohnB+YKBih
GsdMR6pkGL1Z1N7M91liSSzjM81HhiUQjqjFLJ03VkZ7lvuG/aIn+IvJkhtr5Ije
2XAcsqGQzKqbEkdovmVXXe3E+nCyrjhqRER0hbeDwSwwubWPw3If4wPdOwQdHZKK
8QWli9Y3PGoR9oPv+y/DfqgUBG5DEOV3Dhk+VZpa5Pq2otd2caEBdI6xbOCXTuhl
VD2NUhpHF7vWrSy0oLa1PGCHI+/ewoLXYBlEISBcIFtIUv+tzf6myqh/Ed9keya3
wpzggf+8W9PW586hyYBYJ7DFo7WMJGXJBXBB4e0iHVguuqZwNRQAQy0BDRhzRI81
JVPuQVBZjtlbRX1icMdqZH0OsT6LeW7lJuqIh4UqWchLOSRl2Bt+OmygKelqeu/U
D8hNVUAYyIH2VIsTaWpevbRTn4HHTfBV9VsMNrFyFdbgaWGc0xwFHHV8uvTqs+iQ
lxbGjjQVsGFQKoIZuV1bkjCiOsTPMIyus5BszFnebev8esxuz9IpTKrfCLvYMKWX
URG1nFNo4PjyqEmV/KTJ7xzKfCKCR9ako36bp/8ddd3bRQt5ZteF90PA7fwh3k8E
FKVo/yZmHk4JFc2kNkuXD5DT0lnEbCcB/4sPfZ0YnOKKlUzIODd1OAseTNrhoIIx
Jo7BCbgZQRHEyDDosrFAi1HHzRinxW96x+yYghLT1V9zVQkO3Q9hmrC+tKJ/jagH
kKBpJNCaUZ6/FUVMhbyHFnNTvsQYU1uQlY/uCWt6OgT6Y71fbtlXgiVreY2Kk12w
/sJXQrNDQiCGpaUlK+1Iu2AtjIQVcB5zkjcds2ItOldGZNkbLLyzaF/jHYsHGAgP
yJoChKJYqreBNmDdlnjTlecXm/Bmw+u0fUswqUVUf/VuSZGCBe+zW11vkkWWGUg5
gCS73/5yxn1DqlSdq6414x3P5GPLFDdDomHSDDIoTB8Vv/M1DGUhaxkYCtBw2pd5
89Vtu2CWXhvqCYPvcgjyLxRhmw/ZYXwvLbAZuPsCiJpOy5iopyoJHV+m03ghYpdq
DiGlRJgzSqu3NzPAy18IzUncB3UGnFB1j47VdlyAgvQQzN0jfacpoL94i4j3j5rh
Nl9iKSXyakVo6940IGgr/3W9jMUWfsN7p7GJcsqdTPpyGo/Z+llYEF0wZldSQf6D
Z0RdDSpYhjNcjXdX8/+AfT1qgDpHKhaZXxWOmP+K0R+jFWeB7IAi8mD07GJp0+Hz
Jpup+0eci21LbopprFNfk914wsuIOlPeY0b7+xzFt/hHvEI6f1nq6PGbcjw48TOL
nEbAh8RHCp1Irp9qxPwp76ScqbZTP+9LrWHiluc6VaEqI0/bfLP7TVxC74I8rQQO
n61Uya8cAmZH5917LQAHQToakkJnMiIUewvq0K3m4SdLK0mi5h3rpetHTmTj46R2
ECDVL71LhtaSPUhqznr3E2EGqkdRb7GbuObUjE7fywQ8Iu/DlD842kOgZn4gwu16
/eucsRXO4vcejseiVJhR0nWzMFdNGiWaDz2aVZa83bVuP9iru/Hq+JCfg5NR4s88
69NZHFZTR9CqYc2KGndpdY3gwUkyrxZDxHIMIJLE8S1FnI6c6wr2joVLWVF4shM5
a2Go6cAPNTnGJUMMt8BykkeRBHf6gm7pfEZ9WHO0CGMzkx0zgIq8P/ZmUwTbt9OL
6Nb8K9+DLab2BS53qStL2HJ0+wWOgmwxlklc5t/8ILAKvyPjVNc0RU7co7FgvqgY
bpOnDwLgP2Hn5/y9pkB6fQr+Lh2ii8xAwp51t5AhU1Ls8obWcpop3HMKVD/mAEOR
vI3Lk5z0u1jINHADqvJRpQC5rbupWnNcy6hvfu0Q/lyasUng+lKxyUBMFZZtbAAs
xypJM/yQ3QiXVFW0bycknluHt+STJkJNl8ZTAGbnsTfjeEPzOJ5O8zaO8aHT0tIH
HhuakB5qZOzvN8bvIRd+1GVALo3yhdFQO5CL9csfaWTzkYDiesAcajo3kWZSSl7a
uEhuuRtKSeo7jtwgD5yASDEK/VSmgCulkOY/3fEPY7MCFwRaZx6Na7hlH9VbhQIy
8+yu0GRywig7ewBp7TzTo2cdiyc/Qm/99vh3IJvfluF9CwErnzamHtefzKWu47PZ
KbG3Xeu+GPu7VcKONuznSUyvY+9krl5NauHFRih92kBxjuQs/HqsYHE4CYpiBbhv
uuVzAuu9LfGz1uU3ycJg+MSty9ohn/v3863MqDASSI4a+Jk0TiaWssiJjM71Qwna
6xJsIp2/aurrtALnk22Qtp30IfGH48kFM7hFJ32vMtbiiuNIX6ay978s7bgTvQr/
MXI2cQoNpGR/Z+/3yvdqQcJvhuYDu2NLtrpnRmV4dDqxZld/JD3H5V7P9U+0g8vU
T/teNaOEHpT3Th9tOMXENnsVCuHAbvfaF/gWJWc5ilo0oVMJ3PC50N69oR+PamLn
+sIKPwGxKtE9hYO+QY+Bb2jl2eTHpgwZF2ZPf+wNMhL1KRjFv2RApw0Y3mzdTgLz
i03xWNnBbpA0NlalMKe9+RY11GYCeBvWnEdIl0rDxEo4cKB8MQQW4s8y/ogYcudo
7SuKm9gwN/NYnPvqN43kf8c0FLwEDDKeZED75FZ4cv7QCIvQbqjaoTDxzG3o4pO0
4bZiiytJ2iOiy1C0tFPJtq+8IPX35fEYFVAiE7z+7rYfbPqRHdt8YoKrpbRlxkqD
pL/E5xc+u6uoDiA+sY146stdgdqa9XQvwsnsEn5mDqjhJLo7qDGtqXM6aystnal1
QiL1BFwqEHRqqn3BnvCOmsTv7roBtxzCwW4nZeKzAb3pTheGCbHNy9xDO83mxr8P
Ebliw5WotdFdMLSItpq5sYWR64AnF+uXqR4KCDDrRY4L0SHhholum8FI1nKEJ6Dp
Jv9KvGhJyYDDqfiHs6lH7d1+zOIdUbxw0SR+5ZvYLnjZ/NC5/fmwuoiHkmHiUQDk
dOE7lkhgGZp74YDG7vtWm7SW9We+4/S5mHYolbDKN/RvTPqfks3RgowV7ZFiiBit
Sr/23x+E4TN9YpK4wrOhh3L//gtUpF9F10ZeTVO7EpByCpGp4WQdcN2Jpdf+Uha2
0MOyfVGyxEfKF2lTwzze5WqD4FnDwEQ+zRcaumWOIq8PywbTwmdMUnfgrPJCaLjP
0nJJsB9JruzHmike5khcXznmLQ5rS6KVl3hhnYOKGiMMRH+ZULdIB99GvXKs12Fz
NCp6ttdjiqB1eNCcaKBX+UGjrE4oQjDS6kz/9aoGoobso8Of2EvmNAF+SJ6Lczxf
PZK2ET+0ssMvqxDdzD+3cHJTnIMERUsKwYTTs3b4ljfqzE0RGVf7XPdYq5bqHtx2
5EeZrjsAFUbH8ceO81yMCZclKXnDjyHqa/Xr15EzTzwVBsFyApe5OqtKSJdwUSAw
BJzbAieJxXOAn9/iLphRf89k9QKbs6/Go/x2rf7MCZM3EuY831r3X14PRwfQ99ij
PZ6a1DTNVWiGsrQchCPkRCBa6RvLClARfPTO1MyT0vAukFhKpwLGaleHEdGucZ61
J/dR8Wxa9u8JfEP2pBhK28715vt9piCevHjHA+GQnL+O0D8AbvJBD5kc49HZp4fn
JG3o/KA5tJFt1Q0diM2tlMGYYV7pIjOCS3tY9qE7lErWnLD+f+4WwjnOCrcXcVCQ
KGRZaZYY3ZDhKhXyQ+wYvGEOWRFU2AFweEuAj9C/C9dwAx1K3p4BcbPegaO/ejsw
554Wx1TUPwxU6ReOgKUmnzELBKEpQ1Q6o6gZ6ZkwHmpSo4unlNT0Ym3Kziq2V+br
KeEzzYOg1rdhurJwmsemGfetXgrlLebN0bh94W825cvcvhUTC6NKbwGgJkizU+k2
/xEDQGL6tg9uExYaZF0MIefo3OFf9CkZR4n9zOjN+cpg67WSu1Hwt4wxlGxPOvTa
cEAuJZGzkpvj1yyUAQax31NmDZp51wtW8AfiGELFE/UTMlblfd7/8g+XO0F5GuJM
G6Jnaqk2FHfenpcjKe6PesamR3MZqjrMrdNyT3HXu19avYUe299Kqz+smYzY7liN
gth59GF+xEl5vfJ+MiRq5Nge5vudsGhB7lCXDrbl1srIuf1/3w1dujwsP7XNPzzu
G73B0Y2Bvx0PkrAHSUdcdORg0ibhW1y96lun87ivdw9fjxkP/5Cw1+rBOBhYE+kS
1yWvVtLGPb1KaVvl6h7UzsPY8oZX4JoYctkDbDJKtaTA0GOEDeNquW5OU2C+1zPZ
mNPueibqoa9EiKRxU0Rs6pD7GT0mEedlBDQCjfwy7eBLEh0QuOhdG3Z2PAACFuDD
AoIemMM8xkFZaks7tSYMcViIMzIyJzBNwdxeKmRouhZ3GrSe49Teb8sqq75qGe4f
aDVRxj+mevD0RW0bc+oXX9T1DB3zXNVGyD93Ju7BRTVkFhhUIN5S0rH3jRZk87/9
k5SXuW+emj6CfHilT4QXxSfBQoUJCmlLRmCgPKj9Aa4zOC8rk9k/2PyDUdBH2LRo
plFcnEQvxmufFnMZi7n9t0IdJ6Ns6v36OowrET37Rx2KB1VclSevwTSIlV3pUFwG
xL37oe77P2+9ZmIeBWmJ0OMfmvO0emIIhVi/fUwRTfyPhtN2PPWmzrlQBqrOiWUy
+crVmWYEj6/TH+Fsbgb2siDfIRTKvs8JfSw/qQATtWGcVTEBiAddEw2otiNQN5Oh
uz4Vz3rPE1BCTPTUum9Pv8IX77AS/1etjjRYWrlvrHqPoaHvXi8EgqZydQVXd5dU
q9S7UnE6hs4Wz0I+V1c2nY2ie5Q13vXxkhngZ+yGOxCZePvFnAdlgnygH/wEF7CX
MyhHWSnK4hhNfA5nQtH3E+CwBKXNK0VU0qe4etLscFlfIJu1O+uZKNHkEOaJ1bjy
Idjd33LP/WLk+H/qINJA7U0x6V0WWdmi3fB6xiNGUe0D709BZ24wRAuOTZGWQYOm
UmGMvuyavueVxXg76xjEmXtalaNM1yUrOkPVoSU6hNYs4fxexyX2qVKUx/0e9a1w
fhKY/RIYc0kpFivuI+UTiVjAWo0pFq9PucuhCr3WHpEvkF6eDoJr/5/r7sKAq4Q+
f+B8kKO/BY/o9mydjhPKXeofZ03b4cjwmyQkiSmRzDFYoPF4jHFtaT1nYwa9PmTr
M+muK02u5qbyOjeHeZXxaFkia038alrGJG3dD3Dy1rbo3Y1bYyLj41U5azDLLPJ6
yeQkrMxpnnkR+YrE1NBJV8WmRFF+3QuOjWG03gLiEjhRRrp8/RCpODWS9FVbOPGG
tV5QKJ1MVbRSeoDjvSW/5bD2H1V7jAducZXIYwQpHlxr/fiZm8of1AP3sIpN3N8k
UQjLtdxkA4sMtgfeJafW9MKWlMCT8LHv00agIcNyvM2qewDcKAwrWJf6nZXWltAS
RThelSjYpNlIl6PNAFOG6aAHC6/9ecp/LXrZTm9oK6IA3Vm1QKrWbA3YT5m4ouUG
DbSO1jiJ7hiwGcij/F8e0dNmEHQPVqPZ21ZB9W8HFTye8numwiEI6CNgK2feX1/d
RvTz0cSKXgOvV9Px7XHBfS6uB1NfynMgYBu19AO6C5DDexmWdCVufI1+LvovCEWV
TLg+mfT3KpgdOSOhs5GHNsydJXS+qr88rERzC3QzRDZ2uV4ZsYManwKMxO7b6yIn
h8vIdoJFIZOq1Q2xLqbSFFUr9yAkrgIrdIXlMCAzmM7c+IwgjZwCVxSJLkKWdkK8
hZn2OrPkN9QBihYLGLVlYeVVsSiGPvLdznZHyzXtYuD1p+etjNRFKiH81k39HdGv
+z1zqtrZQNp5FQZzl49t5SDcny+sTgmZNPq8HFjXnNfcPS8iAOAhc2YWwa98WZCJ
pAeHOGcecP9xkGjqHuoqZppOlWSnr4VCkP3I5kgH19rAwJ50Nw4zVL9ffECjCa7F
uyAyExhpP1JAqFre2y7OTnsSSq4Y/1UnWY/9VPkpEr18RjgYbs6vk/q9WWNKXvRj
JPJyNccENrfkvna1crvjvEy2969imZNhsj4ASVa40K0f7HE4M+q0McWfs4Hhukv0
i/fvpNiS5wGpXBuuOyCI8WcZUUtV6yTGMepSdo9Dq4GzlzgB7pBYFMDy7Htyxd91
8Td4DZE7AqtY++tVemGh9Ymono0ILNfYmFjoYz6UsLX5blekAMyAgAgfp5f0UJAj
AsWQmoe0e9lLqirhLwMtTILsQFiuGPA+SeJ2kYvlX+HLXppymRQ3THuI03ysfS/4
P3oUmADQmvr4yHw9bZtvyXXKHMnpDPlXGn5OJuqydFLC1/7aTpqYOe6k9LpBwZDh
wVKtnX+OMRYrE8cr6LQccaI53k/9BZhkcjjYDa3DnmG/hjcdvTJ0LhPgoUwX60/6
JCkw41bz7ghNfn7/pWgBzWwKCJAXsg6BGIOMpLszkhilGIbqQu4FIfw9LYZ787zF
pXyGQqCyDmQGjCFVUUsvH1QIHANNnEwgKZrtSPyMfIYKhtYy5SIJtHyRNKivuI41
wR1r/TaEGbvRzcTUuDwmrr669wbD4Cj6DE89ibLPyUtT0tHdVRmSb/Xcip5G2YZ5
7PMzwZWP+TlaDgkzkF0tmHAbYECbMw0QK8MiyNOcp8HnsHZHdNOLwwO5ndUe02aw
bn4FaClD3eqcno6yGYJ+Sb6b4bqrlkHIAluHF81bhzgjf1nGtXgFutgwE45JlZke
oVHbMJ/EbWqndxyWohpeyvRkw988kvmY8ReBsU1aENNfMgl6AH/h7ytXI2EPLg5K
dgscuInAUDQuPsELVgtk5Zi8WCEwYd3I6HhCNaC0GfaaK4w4i77l+ef2VygdEGt7
DyyJzJBizpE2AxTWc8zlEteCOHy8zSqwHr2oJ8rWX8/OMCG4K4oyofAtuXuQ7tc7
s7ERYqNHgmVELgX9+K2Ees4W2chcF3pmdI8h5nOIb6IIwovVUTKa+NPZxqz/6L4a
e92fvHxJrQo9flW0grlfQrv8JMlftytoTwM682fFe6SLq2KzcJU9mLMfCevVx1EF
xKezopCQ2Wip5afdxfE9NATFWAIsv4ISTyYKso38AvbnIZcNsvK7HPevykosAm+C
W1D6H7QuO55OFD8UHWeylAdrG2euvmEf+Dj6nrx0p2gz5evXiEfACJ5Yf5fnayi6
JEgk51Z0yU0wnuiOHHuJUGR/oabqSI9urlNj92rlfzSCIy7g1zpUPNvOEp9rlkI8
WuWejD3buAAixzI2At74mk8jDWPqCxGZvpODbT9tck9anpZq/MWhg510mTEdP2Kn
GEmC9Cq9XwmoqGx8YEH1ncstod3YXyjMv2ILCe5Z2Rywe6P1XSxA+N33gvlRNn5q
uBIIUOAhuxmteoXj/XzITcUOnC1NyeQ4HQMK0GHxtjZx9C5aeu9RK9HFom5z+1ig
JTRLd2pg7pMHV2o1xagfwjaYX+M/V/IsT50FiIF25xt5Ee05CWE6qMP1eeFlTY5P
rJhT3g9UL7Qo0TZsW1aRDz1h8MYW/XKH43MaPzMyN3fxctWHM34JmmEe/0D5hcu7
09QGMTLkUoDy0y15M613UHuKjotfq8QGfOl5fIglzxeX3iNU1Mzd4Orkp8hQtf2G
MR/NGAOTwWPwDYBeWXQ2rm1wNt0Wwfv2fIM1aJ4K5dxeaCXEbG859Mr1xActf4nM
CccuN1S12fi2Nwe+s+fqxmFAaD+3TUpG9T2LgY+GJZlGKf64rmDSSYLIidPdfjWS
3ycLMJDeMmnE743VPh/t6VEYnh0Zu0D3deeCjrwjL7BCzTZn9aRevcske5TdM0dK
rsPkPI8Lacq4iVOi8BZz0lE6IyukDS4iIG5kmIYRMATZgsMfqjcCnPrJjRuhJHp0
iv5GgYDQCXDD054AXdTaMahMZ8p7QAe8JpF0bWfGcOu1WmqSEz5seoxk271A+kD/
RoCHSCKVsx2uIZN03zIEw8p+E3NBFQCNPf0dZ7xcqdk54E1whbuQuYvOy98yHe+h
lTzKGL8sEJDfhnT5xsAwaNeD9y0lEbOc8XxytHfKQo4GCpsKAi3dXG6rbd+Zzm7m
ew8rik5ZU0bOW8Bxjr+sIunU1DjJPdDeC026iXvspTliY3+USeahYgj3rI63wVXQ
N7uy4ldFZHxiUmZ58myt8xSIcsBEnv+aoJ8IWeADiSU18jOaB5P59/z30zp6W/bB
22veKT73H1GFfW8FoEiJAF3uO/vNYSoCL2n9RiGhS5K+RbFhs65XdiF94Xl3hG5d
prE540Kw6l+snUdi1dem8kn39BbfGYysa6FOGm+RkmTLLHdVVJ/SDkQf/vK3MB89
Dtx45yuJ8HcQ9L71YkysrZxpH6NesHMwm8dXQsFTxMpvzw5CW57xUwPrpkab29ga
LcoZ9/9jE1JloUsc2lsLd4tin+aR5LJ/lulJ9lHVMkL5Xrzu2DAkT35ZjtDfB9W6
BfylLPvNKRPBs9cQC/Z7I+dIUNi4GiJ2vcXe3wmm5Sj5aGg0/ILS/IzARwdlbB7Q
V5z9iGqQOdJrIJWxHVUEkK/JOZCstoabzkEWZXb3z4DHKJuVus68oDm1D2/1iKFi
8dGf7KFt6Bo+0gcvfUymfU4nUo8d6TrHdCESoPLjivs1+n8PrT+hVgBmvOJbLB9s
asOuqzKlu5KCHOkiyCRjZIbFnkWjnH+VNyVR0qYIkx7baqvtKH0/GPsVsLe3SXkP
fRy6s4oMKbV03dzpjZTZ/hXy246ZM9lRKFUweZJkoFl/NA0FLDRUflsGXSezqx3M
jLkDt4MYQViIvZ4O+sQGqv8yRniLyaMU/Y00r4SMGQpQCTv27+aMOAsTwT9hbgGV
jPfP/onXGt2BsouH+VsMHAf3FJS0/MDByfJhoxVlK20xLAvqxAD6vDhBxPdjm9ao
qa2bJ1LIgC4Z8YbEiqxoxAznhByGzCUF0AFAd7WrgyR9bNr9FDq6Oq/X/kQN7AGA
VQ4mooHE/pvk+0A+7KTSkMk2aQDF4qdEKJZiH6m/nBrw0pijY/TvOuaflBhptW7Q
DoBr2QsHcD5lyXjjT/gYTFhShoZSpLmsaYTrQFmKEdba6bZBwa5LJwRRvHrf/kZ6
ABRwtsyaBZNMhT7wZ39nplgBTejpDsntwUJEr/OhW7LcR8Hqb5YgqbkLNsRvqXjP
LjHd1i9gw5QroLZEznNdzI1fjWa//LKEw+xzW3xTHyR6RsIlCDTgsrUYHJw8+9/1
vTXlew7Cc+uznaaJUJL2gI1CbHXvD1u6x97vv17fVCvHFuk6bDvfMW6uoHUz3u60
pDjuF7Ls57AGI1qjIfi2KXqixiguuvyiqpJrT5xWRQFdOpTRZHb5F/udoaZuxshH
kwT8rxSip5NF0iOrGg3kiJgpQ1g34qofmpocS0CdRkv5rbcc17gJGFLKc/QRtX//
tkV/P4yY+qEgfsVYc0eZRk1H9EALHSDTbmGgy5Mxs25e7GedNrhVXSMh8jQ048Df
/aMwsnXn5N+TBzrXv9LA/RiAXAhGEAU5oKMFuWkj0m3jno19zdmVn0NYza2UBhD+
X+ugx1ijIOiCn7wpsu8rhU/4te+4Iw5VT3iKZNd/W4kbuM5GfKjzL7xBk2YOcG+Q
/Vwf+hPm4uAnzHhD6LWsV2lZrjJGMGDfvIvLDzNrR+O1gG+fPt+PAH8f89nVRxn/
FYgoEGP7GFeuU70OCLwpTSLi+TAMaGWShmMqIUV1Z/GxmSnIzg6EE6Fd4J+c7FL0
9d62vOxFZBXzYGnGrDajRm3Z3SBD5CWYmYMiaYB2ZuMiR7Tl+8x4PQF6nOeZC8tq
PhsJhceGNhzIM2Zsf6lmzXV6JBwrecP5H0oyISZFKS6BeTmqV+B6F6eIsbD+2Dkq
Es9dTK0g42tZskJCiGv2FZjkG0nVIrLMR4FzEk8iVy6ZVo6Vo/ONciUE7bJ0S5cN
73/oxp8TMwJ9whggp9ENRmFC0vpUsLrajoxeSTE3mUZT7nQX6hv82uos/Lo9Hrkg
tuDKt/kmceSHI2ZhTqS0I+IoAWGW8lJu2fMrqz49DrFwu8JetXsQmkonTay4eWfs
o3iZ0nSCzMHxmxVlQTjPxIVlTBYa3yJE4TeYXbwFJJgHLymUinxc4eZSry2XZXgF
YZQj9NWL718n2ZapZEM3H4GY/FunaM3PapvF4M9t/383XoyjAsmJhh86TV1p3oli
Olv0JwQ+TZPK0+ga71UI/fnz0Ibr3PukctoSJyDBjYMzE0GNaghD35JYvhZY61Op
rtSUyBkszm8ycKOJgknNQ00OfmemOS/AvLXcw8wOVWjfiTlXBaD/iQzNoQ1o7ITB
WdAWdmgKzZnzSuNasZWG1oD7QusVP7HmOLwxrU25qIq3fqSDZDhsf97SGqbTYNHk
BbzRG9PQ5XLiDHwDPEs4+bstn2pOXS9GxasXujB7373K7mZeRDXqx7J0abA9FAg2
ccC66TAjsWN4d+f/EayIZSSIcGMeUsXpeEV0/pUQHADzFuhffK6NbfbiavQnXkkN
dAFPwF4dhB5faouJNGZEA2iCoGifGHi0ji7ZW8oFfMk8T4BS6+pXWhF+tu5/rghl
JhSgV3S3ynaaoMToAyH7heQfm4QRXGcOYy1DhOPIpDPDaEVv4E+GN32gl2MPltxX
2VMzw8+g8w+Cy6sWgsPpQF/PszC0I70JbLjhy3a1+CNLRXzphRDUK++26I+4XOdc
AaRwiH++WzcNSrpwMe5tR0ORY1Kx0v2oI+SGo9kCNVfHMk5Bn+hctIhHiimFANve
WaI2KQU82SjUGxyzw8mdzqEiO2IOF2YaL4rQ0s3Ng7c/1oGR4q/IbkalApNi6DfE
8Zgnu9afVS4tZVQ/Lb7tMhmdBph7Ssj6GOV8atAzp2fGbrwTWP2NBV0SS0anufiy
2M3aj5UtudR8TirLHPNPNEn589bzINdoRZ20TrqTq5PVfbTIrDqWGGkZv3ponV7m
1PeNZnACcdIqeZ9Xr+W75f10SW62N3BxNBIHiJBiK3hK4n4fd1XiR5Ajvmxylq3Z
kjPHV+y0MhQ7NCODBuxECCfv65ET9P6cXXjhfVDEYkwMNlvaFH5tRsSi6sQYoaA0
32JiSGPhX3UflKnhtSzXNG/lE+sUVUXOiFzISPoV/rkPOw8XP5XfQZoB5Gpz7aXY
rlKA0yeyjgdE4TZ6layYAEySuHA86mlkBaIvlHWMUFiGQlH+60CQR4/gmZlt04su
yYjo+t6dtlLml5Fw9SUOZWqMp6cw5AaRvOB8u428FsC7GWoagjp50HpaQapTCs+7
b8+6WdgFwfMGlgzOOpEuW0hE/eL+6JVUn5l9VGG6Fc9eZp4xU68j/8C7c5y2yIlI
UMEHMzN8oqXLGguB9gwYLZZ/9Xy08MvNBXT0mg9jwDBePUA9JlGPBs4UrFyT2Thk
jQVA9Z+HldmftZ2apWuAKunNzenRse+nggTdCJ8+WOhJo0LroiCmvoeAlkKa1y4Z
ZbxmwoqNezbMo9LAW6GNX57qCr4GlxS1kg5eF/7jkijw8UzOQhNhfN/d5aUzwfxC
DLJJyaGCaYtifAwxlubi0Nh+/9I1Lo08lIwqcWoZmeUs7faeGgc9MCSQ7Jj5aGY7
rqZKdtDr1rNxCl7QHU4xwoWdditS2SfjPiJJ33PZz37VMi82bihOLgy5g12ILXxW
epzriffGM7IowtOrLU0wOTWU2u1A9gwHHLzJkxCDdxRfW8fBEz8cqwUlyczQnnr2
MFWPuIL+BIqJgwu3jr9mFCY/s1Bbm/Oe5IBhSjTDC7Rr9Q8XMsW9npqh5NAMcEFM
Nq3GKkBWUoUW0P15+Oi8nZFE2VJQO5Ipc8qKMUWutuLTSyAX9v2dsmqFsi6PbFwl
taCZkSu7Y+V21dBteZ9+QGwETT2lbMcoBEu3d5jaJJB3cnDKl5Fs3EsrueRRHhuS
oszG2vgi3i5V5AAv5TwNfDdtPYWfjsJaJwtch+SpSGLrB5eh7rz3hGmr3eW+19Cm
Nabe6Qx0POsqXD9TeBxtaIuTlphf2wP5LyahhPQs4oMRxSLMHAhN4mSIydex0XAM
tXvAzNMTLCV65/M4LO0p7gcm5EYxcXU6Oirj691SEjw5rSb9n4hI8uHpNg+YvRtj
aVeoNzBUBJzRf6wSoTwK/AIJ/AHSskMwXuSbbCh2AIEMuMT4aTi5g7N35/3zf4jN
hkmf7vXqh5OLHQlmbe3eJzIhBxa/1hR5NQFQdXlVA/kIaxA3aG7B0D5+ZBsm9HfI
+XyjW2EX0lVwZFnteaIhdtbKj/wHj1jPDO1oULD28UfYNZOy6mkJbLkAE1UxB4Ae
4pJioDI/czveR2fHvAFl4peUs9T/Va/RWVV/HGgcDdIan2mR2+iMZ1zuuFBu+ikX
AJ6gHPKd2NmUPTB9odWT2gT64uRhzx2ShSMfb6+WlTQAO+1ccVkgw5/dSQWl9UBr
KF8DnkW1yGw9CAZ5kWXG5y2d5gUGL3vYxQgPzbqIdmThGFixIcJgLWPBp5Lptksr
+Bef8QmYxQi0ynZtOXIU28a4U4LRZlYopADEwVWmtnjNYHQtAxEZJur9z5dyR8WC
gdtNEwG0o62cdnzUn+wbfTrvbhN3hFJmdg3SDK4qKU5LKm2mwLvpskrO9yKziu/k
m6h8hvtbqe5dN/Yzd16A19Qq70l8dUHCkP0w4ETAi3Gq4AOj5/+cOUVR0dtRRpUT
nkDk0YnCc1FuHWSdhkVwv/j0BDcs3D4bt30LSRqfIxykuAxfZIAJNLkpAMXBkMoE
uUQSIbx9Gc1nKRMaUlqypFOXXK9aSKpMC8GmHqmUuE0AVw34fKznfviUg964hCax
WVYkR6eo/5Nwc+awrn148Ip3VjHQPgQ0ZKOJnP6n8qZzTvhdB/+ihAPhhjzBpBJt
JU1scT2MwSeZ/mJManKiNYZKSZ4F1PLfqjSuiDWT8txB7cJ7kISS7SNB5OX5POlT
jGgPzDMfmJ1zqNFD21frrbFiVqIrbIT/WencN+IU/eIdE6RyJsmO4e1vAkdFO+yz
Gv8W334kFjumcia3gsrQNMDGNb/A1ows6R39KerMmpXbCmrqNRre+UmFkXUbUkU2
W9LBHk2FoaWSiBsI6bflnVMFfpKxMbx+6Cblm0EbKX/xcrsRIGlKfc4m2Yxt2y6d
/4Fes65dCQLnfuK7WIAvE3aDwPdFJvyV/bn4GKolgTBbP6T5l1RP57bXDUVI/vcX
sWRDqZQ0IoPidXWovZoqqT097tFxzETG/QZ+WPnUT8+s4tCzXYVuLVpwfSO4EAbA
iXXAms9q8KpXicHD6x9ioMRYBYYtXlq6nQaAL2cnJJGTUi4q+cBz49UrLq8vY9MB
x6wlMU6pAUvBjLvSsfzmR/UYDCjDhPJkV81QWQSKrrJwOWAJksYl7AgKTInGtGjD
g+ggOAB3k3Rr6kA1UoMzhfsmnJKnZS5lG4lM04KN76sj9il6yJDyLrVd0+ExMNjG
40Uey/FmM8QRLMiVsD8LmCTfxzwJ8PNVoforL/erwQqYCgyDbf5R5/7cX4HmK3nv
/De7kSgulnBqMWEkLHvk5WgLQkuERPegzhCKtfqiBeaNwkLb5Irg5E+Q5DLlQDbB
lJSVCoz23vHuL8bpu71jd6Y/PjPEgID5hVxVtxkAdQOSCaH9SzYw9P3YhiHEKdLC
qvyVSij26cSy4S/aQPblpFNBjIusZsEArC3K5j6lVibuTNU+ktmvm87+cZLkyz8o
8fyRo86FLqxxa0+5Z5hCjMG7SjDaQ3bIWykM+TlRd94XSuZQnqwcHT71OTxH4pPe
sYdn7OKDmQCfNzfCrYC0p999/BgLe2NhYvnzxZyC5/hs2PdefdXpc5vpvd9ORr4m
GMeEbHMTMI8GhJ2jqOMSVI/RkYcFmp5fyLOWYsbsLVTi7buXf4V32l05P1foE727
cY6MzWNPpifNC/GJikzmqJ+j+gud8HYGsq3SnFNGloEal59tl5dmrnsGkcNJdd/v
3/pbBg5ujJ9BZUGD1SS9oAx/QfV7L2BhElgecFMBh5B3PyJK5iMWVipP3nlMeo3S
IFRQVRNi6lA15zMaHLjdlXlb+7qV9S8zW9/M9ruo5/cBuq5BtItqULSXOr2r+7qn
YasWcWopV/zHx2G0bCnZUFMqq64f999xAHXbRNha4OSDXQUXGQRkWFxkR0RUzZdh
4TRE+l1z7dsQVpt1c8UMg1wF4AODLa89xti2NxS0DNrDRxP8hBr32k/wfV/uoZsh
vgTkte+cAs4VLN2FpEaaBZqi4Mz5MQZFez0yo13QJ/lj94MK7zSxpBQu7qJenQuM
nh678RfT6g6s6LQkPhNABiUwoFIpY70FSlW91eHzAp7ug6wpate1wXCfj6iV5gYd
UcfJBhd41plKGpY6Rx9I1zVD/SL4hbAQtKYliIu42wTZN2rugjpZ1js6l3slkHiq
eFHKP5hOPuoW7qr0355DsUZfnVo8pdlTJufzFbPy39B4JfQNkSGdUx/RYt3HoTow
ZIGC+hfVKedeUG+h2WOzoOlTdJD+87tDjoa4IIggoJtBWhv2c9aNIzX9cWo6Elrk
QR1VauofHpKKOX0GCAf9LxvXsgewsIfPCvLG5Sr+xVRGpr+sO4vwUhVE9cNCblw0
oo/+VEfHDLQcf4P1J1PHGk3Ejy2xwybSFUANKZ3gGDRKLjSAkq7D4wEQpItKhpTq
mNJozBfcImJtwAnIguHM9HgYRgDsEXc96SFhr5szmMgOxr0fo88DZHnlyUo9wUQP
+43qYfMuzI2+XTlNlrRkxKoyQjz+3GKADFPQoB47yR44MRRQWb7tn6x9IxRQLqmI
9SOdSh8qRkqaZ0UIjkB42dQ2lEfITgiOSXMrljyRHLoitd4XmBwcNVe/dHCjD9xj
MLi5Tdm1eKP+avsS2gnmjqOZLbEF/H1yz9M/nvfnbGaEsRpLiK+l8qWXfjp+UMDh
3kAkcDvRj9TMDMpYeNJzDBqYfftfZyQLIZsdA7efcKoPqyo/H/Sane+jDngCM1mn
MqQHiN3iR7Jv4BSUtI3YQ+b10u+jkR+g/EyXUT4lkW/aT1M1RKxKxfg8Ck9/45gL
TiXRXLcRXGjrGzJ7SDPv7mIBlm5u7PuKqVIY2ksSNQD9vHSQ7EBanl5dJdnJ/etP
HUBd444W5hrlVXrqo6HjCn1E3M8fLjyR5bv9ZDWrNV85TJ3juJ+7J/MbRAfZef+e
ZPp9t0jHLkHixLF0QdaIXX4TKXWljcC2uguo435VRJTHtDuNYGHjnw4IVgiTG5K7
7dmnXxz98zRhAi7eDU62oMPZX2pCG4yH818qZe/yH09xljtiV7yFHwp82ZKouGIk
vtpMhW7hCDO46CeUzN7dYLcAt4nkUPOhJty1RlAK2TkdHZWktosFTJgwoi1IDiFj
ald29wFm0zUP6nqu+t/iBFU270Ar7dLts+Koo6k2CSaNDlSO8WuO6i+ddYUfdDPh
yUDHIjFilTwK9KXO3/OA9R69Gudt+wX4AAfvV9t/aHIdTDqzSgXpULepgHktu7uj
4NEWaaUxyNQcl2WV9bSp4COMGVu3hR8lwH2w/eJ1jBc58F2eLaJGI95SHM2eNC9c
4Kdz+nOxddbsEWYvlXWFbfPPmab6zFtMXYKpqNxxazgIjbvvWNMwwTkycs7SNtlG
KzmbNMaCwWhG9d3AUOfcoQ7lzQU2AyJB/5JXiIiYW6/VN3J9z40Gjid+wXQNzTl+
pLDh0Vg6HNm90+eHO0LZRy9cofW+VbkBVqzAzbJQe1FHYU0Xni+uYyhsmTgB8T9S
q54bezklIXEFCZnoL8M3md+/8n+SB0kd8HT1n7kav8qrLvkBbmmKV6Bsg+E+M9yx
jVMuourjQzzfMFgEyqbZJ3RJYv9vwqAvA6NKrCeKv8nhPuJWn4qW8zyHbPmsNOi1
BNFHlBcwdKoysbvg4bfDksfjNllxnCnnexyzYAKO0EmVlqLFuduiaX14pA2IrJK8
MReaqtUxd8sw4oqV6fC5FZl2Kmlb5Qcx4ss1cnBSUeeSFgL1Cm8UTZkkCBY+4tiF
31T/mT4c9IW6UxYjrU/La8CgLtotytv8BiS/VokOfyh2SX/I7ldJ57O9F9WzzLGw
99Ok4++sRC6HrdyI2a3CA2LybMs113QadcR2qlGpoeY9jQJfYqMxSY9GchFirTh8
zatDmd4opNqfi1PODxErMA7cb9dVKdxKlI136mVXiKwgqcmCKPw9vWqP60y//X8I
FefDl0iIvTNkLveHfr+8iRIluH/yfrQUgaUmU0f09yKI+jDuJBxl7GGxd10V2lWb
eNokySnzzENU0G/E76sbrhTMG2NaIFu9ZcRDdQfMX9gctLKX/UgNUB1Hfo/okVv0
lWf7jomz0pR6fkxEvyOH0saJCmianLfHdUs34zwiYolq13DntGStHIItiV9elYg2
+BKRY/3C2T9X2H5Ne0X6i3p5k3z24E+ohYLMb4WtVzzUQPvxdcJ49j4gLnS3ZMd4
3XQybhNA4eOjHHsBg5lgz5qTJSoOoIrmp7a0fIw9PvvGSuJOe4yVITrm3nZzOhTJ
Y5MTVT8uQqxJ0dlx4hLQlEWXiffqZFfIJ0FJLBpFaGRBhGLNwRxABAkVS/aF/lS0
ilfedU9GjhrSq7OGlfz0zAN9OB8wcY8xAeIjCjHc9pZFzuC8a1btAkg5zbWubbBP
aD70SUJyYbpVZ2Fdtb0a/cm/5b3hv/dGdS9rcJKLDzxDFypX5QVMSF5hJPIwqdwU
YfLwr1IBr68unI3/JISHOqc6KtkOR8//qKqAMsyTRyEm+QPGwIxrHCA6r+7GwamM
/l0UlZmxB4qrsRrA+A59g54gTn46ax6QYa+0IwJuFGKCNaL3jibNeiSyhtMTa7mw
2alrdLNT/MNATIrFPnmGFmYCq6vQWtLVsnBSRwsnwCqr1pwgQIo/dX+GdBuO8WbY
ShFSfSOaLDB1VF7ZwfTe0bM73yUfhWLYw8p0QrxK36N5M1dQuBqY4QpcN3jjrVR+
DMNzNWB5k/Jkv+xV1Cd/kW0Ot7ARyDQSA+N3mvgwosyzGINd4rawlqeeIha66i2U
Kd4Y9RHGEUNGGpYr/Wq4/FVpUG8r9ApB+9LLBfe0FK1f53F9GfOyqsq9bH/HrTif
VjyR2naFg43ysoBNg7bEdSzzCLYLOlxslvvpjYteQ97E6cMUS6sTqEoW732R/cVG
Pfifo71dM2Mj/kJf5D0iqGsTTFJ6o+KBKI9g2+ZgLsPMRP698Qg2Mcz/9nupB3AY
zKm7wLhT2rUzH0NcQw+WP9dtlMDlv8NPHBtJ6kj7g4YVUk6UxF3PTdhS0CWaXSzZ
2B7BgCPt5amcW4CjI3ndeo/MqUlqQg2Btgjn44AqCICokuGUuO0uM4BeUqG8rIQI
od+h9JfhiX0JrrBftSXh8Q286C64LAL8PhkdKzfDO0qpYPBtWcSWVdtf8js+EKaT
E/lpjbDgw+5sUI0XbXc2FeZc2ZM0rEQ2vX0Vsaa20R5xTQYHFbmpXegl9R7BO91v
dxht8Db6VWEgmIoi4W/aMOWPGEKbeTcnmQ9Zvg6vqTgElIiJl9oikWkvCyMBiysV
kXEHDDIWlMyBNQTV1b4nP8WhBLsa6xlYA3Xu6yN1coGYWpvJlmVtmQ8UPnTVlKkd
R775fzOARJ+n4riBl6pFATnnadiegxTaY1ZE2tkGT4fZSACASTjDHh7cLp1gi2I+
UpfagsiyXkYKHu0jBdn9sGkxai1GpiQDLYGS4Lh45pQ85Ck+LjutRS3FmBxTeAk3
eqnxK1Vl2mWq4V3fsVUatHC79otSyCI7ut0HUVHgP0W6pZtoKH7cCBPFLWeCpemJ
jBTS0aJxny7T8xsHtvniPWmm6UiCFJoA144YERArTCGbvZ4Ky02oGHxsxIoj8LAQ
4ZJnsrGqtlLlKHw67c826Kd28xBr+Adazk7kMp/FRB+4saF5o+iFv3kb7cF0WKcb
KUf+Jrq3OSHAiWc1kAz9N4cBel2YojTkH6wrbyZS4kd7jqpxw8AZMXX0Iw47yE+d
sDIGUmT3N80rRfSSkxaSN9taFBkrM6FkFu61Tnj4DaLbf0yXkiuQ9nryNJZNiIgj
Kyc5UxY5uWttHuw9Mc7kElagYalCsHVpMSO3oVimvoMLja6sBQYJck7cFyt9W1+0
6l7uUDPWEh+Uzz1FlIaSFNEbtp1mfEVWA4YvXxp5Qa7Rx9PKpGNujTYArDR3En5C
1/aMWCKJp71b58C4amffEiVT2/1eARpK9SGtrcZtfCXubf4tKGIhrfl+sRNpNbw7
aawhs+CPOY9vjcruC5H/mcTVN6PFKZx31iEsVhB1LpSzElgn4p0GbGmtGnyb4udR
fMwIiMrd1oF6AehpXQDmR8SqApRsheAFLwCa3eMzzk/vVke26jBIxemXLTLnkbEf
g8DkbqKoLh2YEnSx3fAGRjgpCedAP4lak56DXogJN/b41Cgm7GHgySoXM6xoBSqh
UZLiciHBVnWSyI48RUoyIcoQE073pz0zrKq3U8hZHZLm5AusrqzCTQe3YZAUOQdz
hZSOP7lIhxsFhNZLLJvjTIJlwrMjXab+R2s4mzrklLRZNPj6NSJcG0OngA5nEcvL
kWIh76Q7BXdCx6Y8Ki/zdNC0BCS6FHQQKoFNxrDg7e+EH3AeZNC0B7ZQNeLJUwZA
7dgThLA6/CIQvhPf0fd2/pGYVkH8dkoVp/p+BSZPpsBacU2at9SAozk2Us8Q89gi
0b7hXxQnrZYtWpwVVXu/EVwgdZZmkGyArKg/u8EGEHOs5ZgO8tp/deEXUWcpzPci
OBQD3su1tHvJ7xaCSmYjgD4+CjTeO3T8AReJSYjsPZscrBJP9KWMP+aLoGWEHMGW
6XY3rtqyROgxnYSeZJ1SvpoVaN4JodehL2MMSUoQuH+HNQpKJWP1WQUDADkB34Vx
6DjkLNv4NMkKeYiAdvgyG5syXSpIkKyMKMj8XP/1VhbgCj1I//t9K/Ktgji5ExbL
w1Ui9N5d+GO65oCuAfcnfKtiNvY4bTleICtfTmgRzNS53dYmoHh5/Z1K38yY1uMg
d9B1uCepKQd8Nfza2m4BYhRv0v1qfE7XRvQZDlceJ/aMMGpKXTNGr+6TKPnuq2mn
y0Q/uSfvClUbuzbog7UDr4TFmYwFRMy6ee33JVCADkzU25zcuddi/XAU2DE8PstE
YAWA/BsmLvKki/rRNIGHOcWr0R1j27CpWNu2HFBq93I+txbExOuOmBbu/LT4m8s/
1Ulm8I/O8WaQvcXF86ztfNIU97rqGjVEw8fRXvtmwzQ0BLVRLziSfF/KmnvRN259
KIPkM3SQUKiBimcqaezWP/Kyb/vTLUcCvVfPW18RAjNrbIQ2G84gMaIFI5VwVRpW
50nncaNWmqLywBGh9gxjL0ih2dTIWQWvRFQSjfSNGXqynSwOwvkMi77alxDO3mx0
ewPweLy44z1JNjmoB9u+mu+3U+YTtO/ZAxJbl2/WW0tU/TizYA8KqoSxPANdRTYM
yil9Jb3mPRAIm0c5lnyTCYXeXlLsQ+aPZbhve56nibZhPiLvDqnlim8fRpr0QYVe
T0vwWEzM/erd8N1wdXi2Pm8DQAadvyASiAFoo4Jefcvjg3rkGr0Q/Lteda+NK9aC
2njG+1upmuYt+so/lJRArJAXbWTTvTooTe1N4+3BOXfvGGJLVmkMZDJcZr4vyjN0
AzMqQBklptjh/lX+nCFsQCf2fbOUOsnLoVT7bHWu9iALKlL5oxXbjUJBU+nqeL2t
i8ioxoDhKgYpBE5RImI2A/6QCutl095TbhkVept2VfQJXsAKcpBU2nzDfqBaQ3aL
k2fy6l/71qI5+oJp7dORR+4tDj2I6qy+C1Vgib5q8OHuIzg/Ex+y7Ny4hUreLJLk
r48G0j5NjcQWKvMX7oG1U7v91RfDijTdAepmU8TOIzIhuxRtMMjgAQaRzb1XWZHb
/zDS/nz6OCKHi52CoVRACSeDHX5eL1Y1kHjqW26pM8qoDk8mQtzJajq5iKIiNotO
AJphKPOVwpzqpL1QmiZ/yRWSfUiiAkjR9z9xDiWtsBBMlJj8uTR5dVMgmZnOIhl7
f6d78DKQ0C+6Xhgq3/1SzFiXkoCpy7X7CrRmSaNUalv1q+Gk7wCC6rhbTqEMWZfI
2Op9y1r/UhiEkoe5jO7Iuva8MaPGyKyks+1l+kd15havQbI4GaZCDPNDS5u1od4F
swHY0O6g2EK4z4TDh2ilWDu0MRKMofittHW6L9PBcJkLuJ42Gxr0o3KYJ1gjVi1p
Wixu25KMF89KwD97VuxISlztYJFn3kbjnEbWoQB2t5JE+jvPaQQsxdHQ9cL+iUHO
0JgkMgEhemL5jfDfSiyrVyLYF7uyotbKz65wWY411J49RcHQNXjPb/A8jh+Wqawk
/D0hIqQYResprwj5ULDrypqeTdr4tyFEOe0tl6u/FH6qq5bgOux1KdsXrltZXtcQ
/AJCeMfoTi4ZCX3mURJJxtXuVpACZiPR4+oflT60LeAraOuj94DPMik81HzCSUHW
QryqVsDFdyRl/R3t4SQAoCBnvbD0dZ9UIdvzqE1ndTK++EbwPmGkm8R5h0TE/ccN
yf2o5q3mXXjQNed9Juk2r0lQAioE59Foq8m8iMkYb2tCa4v6oacYz3uQYFk2QVMP
4uZXM22BAlh3QFcezuJTLBnUTAYH9zGOsoXIRTn0N05792NEzxiGlbxOFCohyO5b
z1hoIMKnyGW15xzPFgNPG0VN50bjEajVdHgVeb5lN6wuc6nL42kwo2DYHsIvOod8
U/sknY0ZS69av56E/cEGbjFiFOHZR6J55uefJOi6TyloXKnY08bCwQ1BafIHc+VV
uzEliTi5B6WMSROo9jXFtlHQlWAbU5W3mxvGYuVlp30U6+xTrfKVgDE4sUOb4D3J
Woo544RpCl0v5twE7ExIgcc0YnHBWtOYu/zVGdC4kARY5mAP2Fpi7uUIC3LAQ56p
06719afGMXHoW1WSttzs4IstIKP9blRbYbv9Y7dY7idx5cWgI2mPTUDCHjIasSLD
qBtNevNu+EDA9bpltGHSgozHaNhG0EJ4JB+AZ+H4tomKtfa87H+U4ZVMvausLFSv
aYdG+i3ZmaxVlYUMWP66obvc0UHqyPSOBc98/kTyN6w0PZAh7LbmDIN36IAJMXUp
ALxJV3HkEZanp+LPfRGfwNz38PbC/K0U6ZhxasTVvNNJk+3HFU4O9suKuFazhd/h
xSMzkrxH8AZkPwACB2QhOcCHbHRwgTcgB1VyMrp9KjW9hItX45NFEUcDgCgBsWw5
eB3lXVYpNHsV2Ik2ewUuGmvrsDB6PFchudL14HG/nsidZba+P9GLwWEgW5LmEMeb
jdfojGF4YL7ZVhDmhspjU+L1dbFjd0Tfco5CAIKkKWOGHW6KpmiFHZU4Tu1F2kkP
uF8UI3NskIrfDPoxpUekWAVdsQWabLixna3fpQ0jUcZJVrp8s5/sBdM7v1KN/O2g
YO81XAtBL8GlNpjElWVUA1oTihIiqrm8y76Iy0eJAgOA5oAu7v3WBMwtTb9seD+y
ZnHkO94Bz4xoHwN0CtYHGPW0Fr+s8Ylcrwfzbko76NFwtSZnYK1RanT3FUeiPIhx
5vUmghZWPMgAxll2skHEGzd7jXZ3CidWEdPfRdXUf/DkDMFbyD7CeaDgHL2hmLDO
hB2HdiW3gF4XjAMVYNazM2XWtkRnX0yhTY1LSlIHWgvb8GeSlrtviIstio5/VYW/
MDqJTXoe903CyPzh1D+ASHAw6KHjpMjxbtu10nis/B0ICKQGiLuIWQDhdCVDQAAu
8BThvEkvdklHaxRWYwPSFqagO3oB+bN5OOU3cLwF7jaGA+5RfFdhq+P1QbeSZKvw
zobwVkofWzqU3FZ6I/xyobM0sh8Mk8JBdnnw4OXjB+UcXMwmbsWd8G0YbIYlPAqV
wWX2OOcqOGBuWGrV6PQdCf4PaImW2/z4XpF1P5sdt71qfP+GEU2mxP5tVwW6wKvd
KUMX+dQ/+Zf5fvI8iKoCL9dBHseW90RsAE+Ayp4mppBC+k4jyVaQjdx1XW9i+mA8
9nF7YST7wXgn0Zqwnc7UnLvT6ZjnAhRFpJ6YErzJJRnc0owtoqLQXcWd3dXSgvWF
yRyBbb2zPMxMJEX55rUAE4zpg5ou3d1ExeAos+NsMYe7iXiKf9Kj957lQ2x1ArB9
8ZL+eye63tCsk5v9qUYqNvg+nSTg4P7tuUCpAl2pCbKQKOdHw8cd2qOSpJe4Cyca
Q8XWvdXm58fRgMKShI2n9WKZWFJU47urjS+385OMyBVY5AmtZKST6fo+NMbySDPn
Tm4RBCt3jW88h7gomGaqhzpITAjnmYme+jGbCy0JF3Ep13e02Wujq5itYz5HCs47
npDZQ3TEz8KIvz24H1Wf/9XxeZCtD5dsUm2bgmyCFE/YyxfMdbBitH7dA1bP4IUX
bfT0MFnA9zwp5NDXAFfiar8UtXTKKdTRANisA8txrZVAiEoHh4vGmpidIJ4XRL1t
Q3PGvjq7UVrkgWSCqc1dN8tS1ror4U4OQT6ojZ2Q38+WDv9tWmtVXIT1zRFJ5ylG
S2yR0eiAX9KD/5Ls5wDrDmeRDS59X1BDIV6ErCjTFH+72itP/a80IzEO7oh6/V3O
MlouOMzwKggPw9nUGYqbRMfs8HEqvWGihFOAdthfRq1AH2gYiYoZeWsyIn/2k0kQ
U/J1+Ayh1g6RDNgiy9t8qmhPsLU2JoRlbyQVxaBRV6wpo7gwdp5Kf2Id14X0aFCn
UzL8/DYpZKrl7I0VJYOvAEALUfm+58Ww2BvDLQTzvWWRtx7J58xPNt2k/axxa0f5
gzmPpUIYY5Fi7RcXzvXsz8NQlcufdWjatv6rhRKIva3hqBe1P2q6uXEumwb+Etoj
4hignpzwquVLhS2i8vSxkjBhWwoQ3JmfnnTw4VJgp7Ziqph3trdQj06utSyQv0Mi
rg3f2tjc2asAEKoqNaeTV6ibSdMkHerH82X3L6RkUB8kuOtfJbb6e3hVcN6DjjhJ
krICtRN0ahP55r7TEBV1ZtmLapV+BQnlCP3TZrnmLxbMCXFDPk4ds0P0AGT1z7ar
Edn/gkTChX6/Ry2LtZTJ5hNllffGnb+MDMx0geU1U0zwctV/FgkDD5Kf6E981y0d
q05jjBvL2dt8KM2RWnkG9q//S5Uofh4lHAd+x449OPYicB6NDsohdw4vxTWQyMia
W7X7PVV/Vvla7mUU32j8lfFz5/Gbkag8K4teIB1ngl3K49DpPYQocLRJkA/O43FI
PN1dFe3OwVSwC3BdZb8xOxClThLs6kV3UD8AZmK6lPZVT4EroQbGdHuYGp9zmwSU
A3UsMhiDzXEFL3TaK5+Ar6Pl5eJkMjpTfMDk5ytAXFgfUF4SglctigM/DWgYpl7C
GBjipElCDJZ55M0WPU+xLJnvAXaDAlHLOM6Vo0Z/T1rtOoIz0FUSI3xVF2ZON++l
uGXCA47Q/+AKnVgOJQAFtk0VyzhWxPqyZnVd3hEqNvoTpbp3tp0vJeA79U29NuH/
JoLbqrhXDyVHraJVHyhGAy3hyuYuQS4jCkypW+fgvZQ0qIkOxvXsPNhlX93CCsDJ
WhNW7pRvrqKC2NFQSvaajNStEkFh0Th20nU4TzkigWLKcdd0c+kLvcuhBcyErsLs
4og+FZ6pecSTlTdDXp7kLuSRipi6se27BfEyYonZrBdesEL1trMFalN3z5vP0On6
DUXu482+fFxqz/vVqkah3KdEgFZMykC7tmxca7hEpAO0NsxIThPEJYHnr8j9V55K
DtO1Nb+oowcXZYTU7wnkGdMZz9UE3Dr4vWYZCrWV0bI9YkBeKNAfS0/48N/11eZW
Ct6qoLsMyWDtW3ClJUgJhyt4CcRKEUQk92BeF2cuZtIDzjmshQi5xUNp2DKBweqL
OoSThTsNVSSYONw40QpqcYZBVj895acgzq1uRtVbnwftjfhY+VZEB2jzeL28Ixkw
+97DC7Rqt5imCyyc0l1wQKnOGSYaUmaXOCiD23vzrLWzQx3TmP38BTaTZYaRFjWm
k0k9uEAvEf49KO4x7OVCwk37nCWnxSt1akzVhRjsd/SNnFvvn5nIDYV5Nc2whbI8
qic05z6MqEBsjt2f83pGWIkDauoPLEsA/v4XkDPcLJvTkQbvbTyAFTYN+vPOwXrt
jv4cHjABthkEwqXdOBrRtxbbaVsm6p37XM+w8DQdKPEaVzULss8ibj+60LJgklQF
ofZV17s10dPYmyAmyWKGujgd1Yb0pdPhFQGBMVOc2fYQqfeGMtlKDlKC9ac389A0
foafs+GUDVnD1bo/bOsMHQQpMJOOrata7JaQSAfahLkujFmbxErVu8wh7UBuzi8W
stKoL3j12eTfyyeJ7FjeeQ1ypiBiJ3jH6RGgapQqkRFbtwB+nt9Z0CaI3yWlVzMp
m4aeZP8n5u/ROqMH9dni00vltLiPKOI8mRJKegM2lgOl8S51UtIlEQMVM0h4Eizg
17foAPDRQBp7YbXaFh3EeZlVqNy8/7qy/UmhaZyhh9UzNnn1Ri8nQUpMIoYd+et0
yNE0jdovk1C/QjKjxSdBIs84wJzKXJT5dt6NmuoPUKBRb2/aQfwAHZne3a9Bb0DV
XIKENslvZXOR+A9/Lwj7ry74tm0tUlFb40BQHhgtiUSTawZZ3NmHUevjJfoXETeY
Tx+vDDXon4Aw697PLKMVief3p04hCLnF3aCRqhT62eWW8ZuCFQ548z5mUnwlDxRw
xuKpjBCjmD2KMz7whzJP7WypPVfD+rf8BOI4SE9Qnattczj68FQX7pE9Cb2P0SOi
G251TakciztJDNkb8XqVtj8pE1s+9EznxZaopEGexMIJh1O2c4KGkUUvE7Un203C
XfV9ogG8GgR52iU49S7d7908DpE622THPhHPhL/2t9zJDpgFpzeIhMWqs4lkSAv4
GhwDYNvGhWEUsbJ+iB4lg0lB/Qo7mnd3YUYWKx4eI5QIb0CckgOSMcLb59v14kTK
AEUMck16kjEzMyxaTKd5SvRNyAkgUAQffDimakRm/XBMBZCLTcu/ngVwooBGUKck
lfNurnCoFZDeS4dtQhcFpE52wFCwb1RRY8YyMV/MMeBy7PNxsZLipJIQ1incAtih
eQmjzCnGWANSEnskedNbYPUM2nqMrMx6bzPLGqJ9GVPuK/ZxE78F71987vFJQMuS
3GoDSA77aY8NVeBJhJ9VbN4qSvHdLTlfRo5RR3j+XGCUKiE3J/8ZooGe5Ha1Mbjy
dqY1Z8BaKNFWD5seFs8ukXPoDUoQ4N3Es9MoHWVmuW+Jsd7vxNnyjjY9kYbUs4DZ
AJCIIJh43EcNf3cknnk6Cn+s/p6os9Hc30Q7DYpvyL0VkEWUcXa41GWEEQ0/PfRA
qReSNToxBjS9Uq0cbxi0lW6SnNGowk8JMAGmqirdIy3idxjoF/+SbBaU7TZ4NXgb
ixVmTo/pvWNcbopjlq+GZrSbXxZA7TRA3o/y8r5Yoa9hguNSfowU2McaAtFhbiTG
GW1KSB6nq9bJNyB+DvXtd94ZIhPcoai1RRU+ucpQpxveWDDx0NeOzUH8uHyH0/TU
n76tQl2VJ4WPUV2Idqc7ZDmb4Fd9w+dybgUu2sBWEUC54U0FMCzncpCgOk39AxYV
JgrBp3meiBWpRcSz1lOImhNDGg/nG8OQu0GZYSW9SQDhGYwbsQEnczebKCM+QJhK
4NfBzjhEhY3+YRmz8vMW2UEMHss9Gj9vbSM9aWJb/mlb69oCJQhx39FmccRBBc5E
Cv6uFj1h3Iwdvmqv8+3drxy+02kcpDKmvY4N+BQbxB2n6IE4veGPYggKBNHnbiB8
E6j5FiqSI9GNewBPccaRZuCLeHNhKFm3iaYxvd35gj752s4h8Sn6iCvS/YrsIj8N
5kZYzRAn7cc3HiUE7DzUsZX7AyApAaJPUfZtXbo2y3sfJ/9iVrjsQ0/wmlZcAeOF
pIE6Rb4GsWUvIlZTF74u59nfa8x1GZsv4shFEajouUW9p7064pXi2RIkUIFQ4kAs
Ph1nujR84FCfD7HWHOO/1NhNVdJ5fzeLUJI85Lq+KeXKUHgYtos9LbKZoYs07Dud
riDVjHUSDFXmdUBkRR1Fdo+Vu8sCf13DC8itCxlJMAyr0VVs+mKptZoFkSVjWSnl
1hYPNwBtmmbaSJEjS9angyDWrpzx3D/JsCWzHlH56l/KoMoJx+Dq2lKnNgnUWNlg
Sm42/HH1NV47maDICxybvFBNlid9GaxNlQtyddGPJb5GvE4z+hAQzLvufscHPqFM
C5M87d5KNlrysseA4nLjRkm0P7zNkmuhwrA8Qsm8mee2ioGHymOc3MPIJdEfuCyv
STcwUVnIAWb/iiTd2hwsFSk/xUvag52BeUVDyVmeoVJVIhLGHteryr1qEyLA+/PS
Pjekd4TD176TRkWLZwte9JtOtOB7VW+11IyuIbPoEFwy36gc5XWXVKUfaSF3K+PE
Ev+97ghORqkI5URzLmTZs49jP1RJrPSVtK3uimRJCn73/PrV80va26UbYIA4gGYl
uGH27gGpQE5uLehYp0lTh1qdsEB0+R2XVbXYkQVjE1i7/ki5VJkq4Z6ks8nnU6aS
0NRxQL+20RtVhCArW8y9xMa6WQNQZtfEdtyxGM3MStSpCnWftQUEWLv+pCp9J0TU
9YTnBhyLFjyfYF+ybvNvwgBK8CuN1ezr7hdBlFMdDef5Q/ya5syArFt5NQ0tcYsh
G0DV3q7EB+bQnEqXxilx1aBoagZynlXs0qfKgIt8xtvTNwubaz7TssSg3dFnE6E4
TeItM7sLZyRJMplQio4O0RFMAQcCVyQMv35LSL9swlG8gY5AxxfKRKgH1cmHt+pv
TzC6c9DDzU2NftCy2wtpk4cJqixRw8DRQwQE9n0/A2H7dL693eUVWcfsOX5sueWc
hqkCjAGbLbdCWlEoscBMtPlUW2HYIrGqfOpV2xxlrEWRuOHnFYTWPBJrtSNZ4B/S
CFPYLna6SvXfLedJ7wmum+4iXMfTosrRK8nHQH2l5nGEUwfErbfB+jLw50QALH6q
eXQy00uh2MEZs9kjLWvd5EcVQfn349cflqcn5R+0ArERdy8cGMXcNdoPcMEckF4K
jGTncHLNzudthG8oCeMsO8N6p+JAMjGUUOvjpDYXGmkSBLpZp6bBfZPnUuomAIY9
27n8GUYFPnc2omSK7L6m3JzG6ZFu3eZ97WXleBNyGMjTA/hQw6bA9rFvweBu0s8l
jFjIb3ZLeJ5TyxPQ55qV2FAL5xCl+o26kCOZ9MUToj+NbMFV/n2lJ/c3t2jU+V1w
/nOyPv6NoiuZbSLqYyzPnwgpp0IbOZHJdJOYYSWkoYc3X/6+K+79qMBpxORxIt4A
lSDfZqoY7O6HsKs8vt9HFWWIot9ytvIiD5BGqu4+mQrkbLNjC0C4EZU7MJctc+VD
0xp12Qfw9tojWDEmrD6q4gBMpBJ6WYUAQ5GAdpDUkC3/+I/vDKzk+riITkQwgU4B
8ATJb+daBglQCF2w9oRvF1qp4iyYRY7wZPvsxk2Uol7KAT047HA8Llz+m/SmxL5i
4nQdV2qD0BfpHjwkSAWbtBAn8v2ZrOTSNNRNpa1eJlTOUbCZQiAjqWoRorHSQWT9
husSMcFWOd4HIAzQQj/ICYuNH1hSQTTS3WNnleKdThEapeByJO8Xj9KCSsAff4cA
sIhBiVzTC29kDwyIWOTpTAfTgrH+yjmjemBGfH4xLI7TPyVBzUQFWywqoy27gXVc
/XRgMc3vkFoHp+g1Nt6CLjWcMQNLJBUbOC2NV1v+ODwXVmPtBR5se/14gWrZTe0F
yOMDQRKRyj6hu8B3Ol0hvwmfdW5VusK5vQeQ8ETOvCDpc6tyxphNX5n5/kYvYCjU
J1Phd9OdGaQcYPU6YErWgYldmjiZEW+Fu/JCo253YBI4WcOadFFmQVIz3o9O+wZQ
9/2lKW23MsDHBwlnLuioTKgNANbpm9mOICNZASwSihPcgzo6vfsvjd3y5t8QcV1D
yXf6ZFIRP1A36dNDE4LkRJ5ZlYIJbSQeYSTVkA7ATucmU0x5wRHK9FWn9rW8a/Kt
P9vren2G/lUaq2mxdhA0EP0HXhDnOysVxLSfH2YbOEV/kcek46d4CZedvMfdBLaI
WZg7nB1g2oHOg3/333h8hsWSnskojRQYHG4qIrjawF/9kDSdaAMRufGGhq431Swt
hbPqU8dLzcVeW+T5YU+ws7HYYxgpnKrklxL6Dkqh+Hk9tMxtE6xjm4xbeIeUL50U
3gKOOF4s41ecuLRjxWti8nHLYMXf5LWNgWVniGSH8zlKRvhy832w+7eS843BWwZl
+Gg+TNw4lKtcZn78rYNQMoodHQ0RFznI7358Ce+Xlz6h2SdMe+HW+N02Ug5MN3EO
OwlSKz/nt1P6vEbr78U0XjjgO/pGLgWMLogc8l7fDIbehIr7RmK+XrkPRYZmnzk9
Kn+HNGFaPSj3FGSX3A/5NJwmygVbpDNKAwvPaXvvie0izs6Ag4hN0T2nZU0P0VsK
eEgqnGzhixymTMklKK6WCYvzk7ajChcLHfytpyZ3uHoq4+oQrE56owjg382mPp00
llNbUdZOQDbNEMhYWuMLvxA4UTXKWRUbNyU3tVbRCi7f1p9RmD7KDKTtvd//nWTu
EV5csqJYJbDU9y5VP5NmGbKEvy7zxPYXRHReis4uzLt5j8BJ1F/P8NTgUZQHp330
BxbfeSR2GGNadVNdLbvFP/URkRzZ6ZvBzx6M/L3qMObJPOm96uz5qK4VMX5STaBW
1qztz9lnivJUQrE2mQTp6//XwBx86Xwr6k6DIcD/DLSBAsuP86v9A3fMgZJPnjQb
3CeHD2yHbq44UD0Nt73+KRFmFfh3iJoXHdJ8GDSI+11W4u6URP8rTEegPp5TXYvZ
UWq1mQCNWSMKvqIZB1lp6A6gMqTsf+X6BI5EA/pBB8Pb2ozoMzrGBvoyQUH7WH9K
MJGquRS80OaD9XZZQS6K+HSIbgQs+G9uA5NL+7xlqPbyAzBEbXu0+tpBMRcclLC5
M6xwqxKBE6uxL2aVZ4lWyjf4c5oLCc8mgIkTqDC1vq37fN0Qy+49BJfTzNBSoot8
1Kc9/4LFxpp3OscUYpHWkIx8ifjKuQ2TJhj1yc4x2FLAEl8ntRp4tZjH+Ck4nasW
E28LBlVKhfuPfj+gl3FqYycvO8W528rQwsZg1lTOzUQMOZTIZzsWNOtFdd7Hp98d
YTiK4wNXMUKJMbKctUN1nTqXo3taDYTYPw1s0McTvrdLPnDd4SyMnT8Noga2MkXG
ZwfSaT9r6cbMKpOVGQKqxL9e078Yq+4oxIKoxgKEhpLXxf9lUU6bUUbUstRg1mZ4
h0nfwEstDlkM6OHqJHlKEEb+X+JmNAa7ifEwxtLWkefhqkoLyFCqoz6WIxQazqeq
HwUY19WKR84MOCOqcf+pgIV1Hsn9LlH6rtu7SDZp+7kniEsTARA8JCG5yPp9chEe
5anzkaag46zqR5oetAsCmBt6HH3xjWmbNJbTmcj1DorC9UweHzMWkbXloFK+ra4f
8DkJ8qWqMe5RUnTnO8vPk/dEpS+GpSo4G+IqecJV2jJwc7aFMA5t1FfEczQyEFw3
nVr3HLX9IFtJsQDnC7ZmpqdTjbfFIWnYdKtDu8rH0mEf/d/Fl55LlgwreAHSrgPZ
yYEqBpy5GdMBPzMoFe4ZI/T2zrp8QgBedTGtejD6k6Bgabizi4ofvrrgtw1jVInP
dclowIcguy5O4E95HmJwhacaAYISIQa7wSbbWj3IkA+GEk8GU1XKJj6BYX7FSuzA
wLxS5DvFfgAE8WrGzXy139Atz2rqSmmmxa6cNFlibJhFeLPUhG4nN7N4DrX5pNsI
BfDgd1hE2MdId7+79F4tkJFEHEESZmkJ3NNXixPalZPJP9UoYRAN3X5teq4lOVjc
djlRiOoBsTfTtgdogJ4kmOti3c1hVvd8XhHxCPp3gLAk8NycV93w211mfZ8wyHOB
QFFtbrFvaC3KzFvqeN9Ho98qlcZ1cCaO6ghs1QVBpiQrm4YO633KJqLndXqC6jtv
58yWW9ML2OVq5/pzz2J0nEZalU/b9/4wgXmr1125e6yH227W3R2vKnmXbRYpwfmv
DYGqbzgiP7VJtoZ9+jsOmfoK/wYs5yNl2ijc81Rz8b3QjF3wInuaHrfD3ZMnGdFq
q/SPHXjn40uHyB+0OAVvLFDHhp41wHgSGBiYY8AZxGe4VtRVgXKCwq17moIgsH5h
TOR/uB/P9waS3ARQDuFxvHRTAU2fGPW0RDH0J7kMSdbPxdhWpzfSgejZP4C/ZmhB
V4lb/7t108yPUBops8YhNaeSDwiGaV2vfRBRaUjEohFKpNiDOVAno4Z/V/1D+cDQ
deNq7FqWXduP/KrbEe7ez/0eo2H235+ftzoWA8P6o0k6dffXm/BDCH984AYkFavA
JiJXV1uQDvWE6IrWneT/wD827MzjF3KwOaOJRdgRSernsI6/btxLWaNVluamOTub
TNQwQpKtbeZTo5eY3B1Z1DG/apMXnniePZKgfwpx/bQMsWy6daWdBNDf7FIzJfY7
Zg+1R2d7p0T1XVgCo9wZ5RR63HEkkxyfCqeu2Ao7CKtzDfjBrI3i3GCuBOWD0f74
kmKejBxUexsuRxGWStBwisMksQf7W35LRWahOki3t12MaNmyxzHMSUfSapfDmUD2
8zi4fJU6tMeMPdYjzkIjOwxVjAPxSYN5lWRe/D/eaJLp0V0uxlQM83JQeNJrNzUk
Ef9O/YKVCuva3aUWC0/aliZwNbgMQpeK6UE6nvkK2PFWXpvzg88IjvBJCU5LPUz5
iwXgpDLmr/nUwbCbay5gVFbp29pzxPxEUyj8AJmmhvV0bym76UZ/dBWuUInZ8OgL
yPf3tjvfz0RoziKjt2MZXs+5u9+x0hs6KdBHyla7WjKr1n+Qpu6zQgZDmi5A8VR5
sllAIe1zXS5CI/EXe6t6/s4x/MPIIo5oagRKtytdPmSU87GEr6BiznDUmcsI8zkV
fMbx5ad6OMfS1LN4rcU08mCenMMfmD4Lf2TXw3BuzOXjcZ8/HcSOoocTiXAERGj1
Rg91ZWYKuPIb55TguNUtEqIcyW3HfqUPEqQrMaTEwSe0jR7phYf2HRC9y6VQCI8U
mKve4mPBLnda8lIUZz6GNw05B9oQXfhfF8pGxB6/mo6szFcoQEfs1SA5fyTdJLZh
P6w7V3SUSrJAERLQF12G9EDDeaEqZhL96rz4Y1w9UzA7E1IZbMT3gKKSgCBVxBVf
JZyAUw6zZfP4Hln1xJuiZyl5V/zbOSYb3p8DsQRDWeAXkyWhHbyZz+bm4og6n/Ly
HAUJirLYE2+9bIEpyHwRwhTQgVFMY7JyAOhppkfL2DQGQBNpCs5V3zSaUhKYw2tU
2pKMmMyE0sFI8BdtIOgbUj9IISN+87ahmJGxJt+yrQ2PQ978D6s7YcThq5MPYeuL
LNboPdah8NyesN8f9JanDgf6t2ONlR5gWzCzWMLPo/2b5Fzh7IW3b+UYMxh/z3x6
XZAiRt5pFh0CnH6Jm1WWpXVr0a1bkqSiN5pnOpcvHWdiijP9fxKL0Z5C9jYKzo84
piJJCjUon1HYiEz9y2nDova6cZsFCHsFWAjlNWG/7WAa+9gQhGN0Gb8I81kb6/H6
8d0fMYefHuRs73KVTL727vzviFoVwjp/4wct0Fd/seeVqhEUwKTMf+2S02TS9tCR
/GT/ODGqhJWoZjbj4imYT3giuroPtVq7JiUwu/+/4si6k8hSG3EWJpRhYpdQWrVX
KEo8Hfb0HSX2lNEL3PhAWYDIY60QvcOX9DzwRhAvKvQGSqzUAFGqMeEmi2fa2MqK
Qn2cEhzdC8SI4Upd+2frbUNoUghmcYlN8lCJgnbswJKA56nM9Sdk0qFHHYJa9zwG
7q9pfsXzEdqIwwH098Q73Og4uDQ5C9SF42tZWNNpgOe3X/4mSzHdwPhKrs9kQs4K
bchzDwgNdtUil0BALlFSDGyNdusXyfKL7f/D+PJ6qHhtoNmoeQd9mQOmCOImHfMV
lFxmYY0UFFNEKqZz8pypcHjXzoHBMuYpQKUB8+NBxGnMat17qddivzPYeIjR3Q/h
iG7S/UwZjm/HDypTf3YoUowGkxwefOJ6Tv15Ts/PNOou7uWysrCeUlt2I1L3lBS9
jEDSg+HcyfGpdbEBrl70jRYrk2pVvu/yOTYUuechoOhi/PPrQoBplEHLZOyN8Kyk
UMdYwJWq8Cc8H7OvOew2ZcnexHtsstuu900wrGi7EMj/vUT3Vd49oPBYT1RUrYx2
V0hXitwpyzO6tuLqHKaeApfBo+6oEnS1AslycYOLlLPIVJGZLib9pgueTiu38Eci
ftw/nZdT78FRMHPaFgcUzFHIpa9vaZ7xWWE6giK4dPsNeQKApF0pfPr7JM5Jjhnd
D1DetEAANkDfyU6xNhGq03iqh+btSoAMvr6TGf61UmgXZVchXTQ/s6I97nV352ti
esNwdrMffg2YDpLLpwMJza5yL9UqfLPX5w3a9YBsxTG/OA3Pg+cLpJxVfWZjN5hj
jIGcC+mUtS7oqA/+YfaZCjwWTI2k9KPc6z72nhjx1ErFmTF5r+rZwVwNuMbKHgms
1/phViMqPKwdNNxwbvIdhuVPKSFwEi3ako6wjJsHHzNFy/HXL4B6Zw7hGg25yqV+
6FT/ymnmRrwiHt17186V9OzpTbY1lDDiIEbFzzkMFRtU6EeLRtMkrUxbKKq62EMY
8v0TY0urzNfmdHqZFCu4UE5Wed1wex1TejMQybvMmU+8EGFFKkRrnHkNSgvhbAY6
zjk8w1RbaTFgYIoWYOHO6Xw1c7Vd0qv02GgnbjqlweFKZBNgO89p39H1jVsjIT4L
SVsvFJKMnLOxcniCeo0MKMOcwwacWrdTpyq1rL38Emad6KiL/b0Z1wr+bzhEqhIa
tcdJv1hJz81Yt5L0S2ETpCyXVyX9E7OSv4pQwwy/Lts2pgPq83EkV/JR3k1ZRV4l
129vwYoVQnrv7sz0FbNKRIkFhFkWl21Tvuj9Nd9hOHnclPCPDWK7jHCvAWnC9hXA
i7BHfhgnaMEi8IynAWhwkyWNIJDVJW1Ej4XLJgAbjNjUtiMEBnGvD/VZ4NLOAoVT
Mb2+Fa/hwZwKK3ftulfeSkAoTFpm6MargSNm/GcCw+JGPY1T2PrdyiW8gXsLKoxs
NB3HEEXgyXjvttJs7FmTndQXirnPxxDAhQJxpQOSj+ndQPIxypUvH/1HLwX2bkIb
npDwr/qSTiC/P1a0I4dqL8wc4SWaWNM711QU0msrqrZYd0qvX7yHn+Emjh7W/vZ8
cOxwk/0eSPh/JmP4gzCvaxNMTtEjOKJmBhAFwe44x+QHoIddUSB53ZFyGdBZA6EN
RPuWjvO/rkrJ3Rjez5sNtMdDKhV6in5+FfaYTnurTTq09C3SB3VhLHNPwGJEJ6F5
fWOag8rc+4uLZ1ytsh/ry7FbatAjnUMIBGztqPx4+UO27rl4SiFqnxmHS6wK4zSi
E7xZyeIbNdJRPm0rBKfQre4V6xAJHoeKbPxwn2/kcga3jEKm5EHgRmlZ7AfG7IcI
rz7rbyhs8Dhj1tpvxpFsS0NXejFPL7tQYVtDDuvxt6SsI7ADeKFzMidNIXLCPvE6
4mZZ8iY3fcExVqF+6WjsIz/fCAf3i1XMLLbrRU0L0dJpjFhItJhWdx5TzPNczK1j
uUsD+K6evVDwteKSDh2+LtVPajArYpGbnP9nF2oy+F1QOm0VWp4WPXyKCraglMVq
NIQ6u8WWjvfez8ylmBk0qVhhbKntZkprMUVdy+4UDXB4XgJYF461d0gDUL+62cw4
IM3AcYNAoWXeICiu/y71RGpnhmRqDJTJWtv4GYdlgcBbu/1eOyDL4zcwVsi0KX34
oQyrFqxdPk4jtgHbHZF6RSlwBEto/591UnTs0VkfGv+/yg1dMX0CyNPiHNMCYSl7
+ZK9koCuFzlJM2MTZ0IpUmYrMdNVyjKBy83xVdjmMxGgcNAlZwV8lD1n1vXcqK5+
b9QzfxwW7AOjH0x1apgsdqjPggSSihEbCzKkUPibD/AQ2CtJ2Cfz1ccOENJaLaGk
sseiZfPytFBQcG265plowYmqtWZ0cMnfBWo+gfJULIl17BSWPNrz+phsgR4CfKLH
woLePcGWHAMjrKqyCoW37Hvaq2e9M+TPX+99eqZA5eHjiqsiqgbNkZP5CFqzwyj9
Na8rHJUF9CEtrbCepnxSmImk1qiz+6hvWtN5DqZZLscjK0p659/v3eManW1ghnU8
i3vNeDmmWXOLhcQywcbwKsm9WAsxJ2ih2hae0CEGdknRf0U8n1traSbKcZJdjqXA
Kl/42tbWiTV3ZBdoTbiG7ySBJ5B6A7Ru7VpxSJidZ/vj9RGzKMvkDjF9GZzuOMPr
Gv+ukTLJ11c9TEXsGST2p/tFQlHssrItrZFW8uUALS/nDqHz03CCjc81vBV83/li
eRsw1PIuYXhBIJZueQJou0FkTZ2sQmi33nf44LbWyKHbxluoosdiKNr3DWqtOm6y
pCrd0Hdjyx3n4v9f0hhWCq8lt5hn0Z6HfycrjEL7py/DPmbDUyzHPj0yJqADOa7B
ccM1nYzWBkwyqd9webwLqHC3s0h8yHufzCibZz9LJPtQuHaWHLkevd0Fk0Tw2SUm
Or90VZBCE/fh5i7bp94Ouc1gFLLtZPhVEzYFcp1Q5S9pbLK8pI3alzkr78zcAGqZ
8IjpMZFvbILIcTGOYiyW0ZQ9zAQRMmeG2FvrtcnMucL1kx5zssfYquDTtskjd0Fk
wIlK0lSy9t0GIpqJoCDrg+siSlvzHHG6OFIxdEkXJqklMb2lThTR2sj6PtNGf/rA
uNiq9Z261474P8OZee6IoulXKR0W9LVi3kGktxFKKNoL193QvxcV25ATxEmHeEjF
qIparg4/GvcSvOUjBiHnTJ5w6gswJvTS2KpD9zsZ8s16Yc4SY3ft024g9sle3L8y
IBlp2jyUlwRN4/OZR0KHMHZ2lG6cateWxaLC5zjmMem6PnLLg5uAaEK2z9TRlXxk
gQCLz5W8OTVnJyM12LwNjUd279Wp2EjGG7tip5HWBJmObyPA6DmJCiNQUMSwI0P3
JvG5xVmkyTxEK2o6DsBeLKyQmNSoETMheFHqGLyOPZmw5kdJCtlG47VYoAjdr3ks
0tl8xhjz05hKbXNOqOxZ892o5R0hA42pm+phSxZyvIseHqNhev0bE+6DWLqUc/D4
voUfmHGLcF80kSaJXvbrzryt8cteDXUc073FDYJHXbKo9R3B9cQhTOwVegzlsn2y
DATJeOQV2tBA8noBIeQglLVlFoBrUQCNLRyNd37sJ2Dk5iNYGVOJrNCD0yIz46iP
+Z1J5pDUduYYYsKL/A0Q6qHiEUgX3DtPaWjtPf/OMM+ymNuVsRz7HbFMCpM7MARY
zgBIfiEh4a17NUatYOvNBBzeYQz2xbQqV/Z4+KYvoa9H9c/idj1jCCVFRbBr4zuU
dFB3drCqfWmyqGlviHwtypP/Dci9U19rSgZPJFEtAqynH5Ndq3mIkqwa6AjniYwz
2nJAawdimcJXlVAyNz72nUh4jXqk6rLGCAt1D+0WY1Gy/4nZKiaZG3Hp6t7o/H4r
d2Rcc8zPeLQ15RVvEW1xP7E8C/QzcgHCYseFl6SjnBvPBWBywFL6qRTynljQ2p9T
skMiigbNKEDR7kh5x/Un2dbmVFqSLEJsC9NtOQxPF+oiRa36v7BUFWQH6dJYzpZT
692tUMKwHjB1VECmXF9toPxOJxj+8JlX9VRNsFYlZz4JmQHWz7ewAfY+FS8fnlZk
FfpwXV1j0dG1zouj9g64RFLKC12/HwDkYyn70uiFsulVoOOwPHAxxUWWAMCeq3IK
JOdr3+9J3WsKgqVfqe9C1OKS+lBo2AmEu4vQf8ypR5eq7Hr02A06eVqiBl/PMNYQ
4Ksh6/n7wM3z0aCJvKZu02bcyLtUo2hlJ8g3S53eCT3ewUEenFvg/XPTCCCh7y6k
/SMHqLPVlVh2oUTP1K35E0EQbs11zl9cKpoFceHJkwkA6i7p3J3r+sk4r9CFUdWg
HZvcjvKqYZXfx5cDxvy1Pkp72/psKYAeiZ+3yps0QbNwyHc1I0PdA0/6x0jRDJGd
Tv6RP2pUmNNcXtrcWAe/dsHg0kAxnIWm6lYO5H/WBTZl39+/QAMDaa8U+bauFgfD
wLZdElCdrWDS1c7+L8X7UJvW7GB7LCEgI2WUyCdONg2AqLLkd3hBNC9Q1Xpvd5O/
qc9Aj45uOeUqTn9mJXnd58krJx6DjV3PFxPio33QupSP7Fxl3v+1I3exPsSntqir
2xY5ssziA+QAriNH4oEnlDPf+ZnGD2pHaq3Z05jgS4wgqpQ7c6jv4Ip05VFQSdai
IrXIACQbhfWj3F6qCBsIWTT6cl6VXv4Ic5eqhXojElKaTohm+XwVcnIwzClFJGDo
4HauLr8/nwIoSPeKLnOJnbv+EubU6fo0Hvfwvo0ac4cDyhbmvWkOrY5g5pj6b3be
vFqTTkibBn8le6Lzu5t4XNLPE8QgvtZWu7aJWjWpo4EKRS4idOe0DGrOlZkQfFwF
3G3Ap706evIuBJgP36ouPma0jOfhl7Eo8JXZMHQFWg61RTGfP+XBzuUpo8/WPEac
XTo6+KjjnbYMJ8yJamVEhqubj1l3bcb8J2OZ/hng/66W/Ndl4MZSAJwQ/0zaVhrO
Fs3dHe8hK8bCeCVgFSruNb1M2KTgel1Wk3ItZTFVt2i6bPTY8f+EcB4bim4YskpI
LL9AlWXD1XeR482E/M/AUzUGWmqAIKddhsdsdN2jdGCeLoI9WPIj7/oohEEBYmsK
hW7GXS8xQVpXi/fWMPrAX/bSTafHoeQYOqjYmq29vhkQYRwAbld8881ukH/dIVwu
Iv0qZVe6vM3vcbjV/m66oyOO8WjF7Sw0QARxLA0Jzdqs02QJNPzjyN0EcoTAwTLM
UFAVpYBbeleZF6+F5ybErz+TqNMhciMrvLSoXxEsMCm2MljHXz3DzNcNrxtErpUF
chKaAotwU+4Q7uAaFWBAV6lii7wKCeotLgrgytZIzSYABrc04YuanfOQj8+h/PfT
n5HqGWrhvywSBrB811OBARnNvc4f+TMh9/K7JAfA2hfvf2l8jLfX3WQRc3kLVgpt
GyrXYShHriz6kx8n95Ca5vA3Q3cKCGP4hq8CVGBvKCsDkIKLSI3J4PoBg0irA5Hh
NWYCplXhuIo7dmpOtpH69Xo/UPSP0rldTz1/bTr/CGCaDggtUNucouUFipd70mV2
C6+p6C9tI9Tea5QWDWElf/wTe1EXHGe7y/2kb7gMpOJuVX8ApTOnMemfxbt1S8j2
tgrNmjujTG38QmWXbe4m7HWdrzzJScJXy4oMhgZI/yFZvg47OznFsDR3cROAwU5e
4YsU33WDllxQ84c3mPZW5IrLzsJJotZ4+eImvDb2sko07h80DSFqMCD1f2e2e7cG
XInri9aIIeKjU+qvgn8JItAhH8TDZvyjMn2hzkl3YGBHuJlrDMfCk6c8piw85Cfm
OtKH0GAuV6eMtkR63oJrj9qiY2vBXc1Xbyt3HLCzih3EEUUXxjqKSIqI5FeTBEUH
9H3m+vDznxrItXMmzMOAEwMD6ArLkq7v3Hkx5ZRKwFBzsmT0kUhVrJOxusr5VMzr
2rI/YTdPpH/+xuzpQQKhSuNuny90U7JrZenwO2XIr4dXfnsjx6u13Lrb0IIMdUrU
K3XEQJARlv5XuYQ0IE7VvyfPvjq4DRAILc2qQ0w8bKSiCQVktZAQpZrwiMvlyCG/
zlnqY135KfeYkvU0XUxcNFflWRkrN98zrBe2Hb98nrT4N4YKIfbD+xZg7ssrCsSn
ecyi/tJsAT7PjYs4AfuqA/dxLuuGeviqXMsYtX7XkEXHRBooxvm0ezFlL1qQbqgO
DnFL2H/eiw6dMcF34DH8j2M0AqcpCrxgPUfQzs85pk6g9SD2j91WQXankK0AHk95
YEK0UkvvfeUEp2AeKlPPrc1NvJhf/jxozLVrf593kaOtKjKxvxLowzOC1xxzVnF9
wxmouETzbZy740gX0ZTegSjuhkj+8oG4U+b77JFBVOGopJWBYyjpk5svU3Pgb2LB
64Gvd3BH1kFiogp6UMAYH2zDL7oeIK3wvfl8ZbF2031Fh7Bi/fPgDhabkzNXm9Vu
obFgfB1KNoGnh2Ez7AMj//WEBXSsCXoAE39J/8WOVcbVRufBNstDMHUx5RF8s4ju
enw+TBdK5o2kQ/zPw871sh53o1t2cKmeACcGFgLc8N+VeFte+MeoKbhJxiHD9V6t
3xfiVNVVu0gLUYMLY5XiZF2lDDPIM0gHYfSVSSJYqduNfuAIiide3FX5DAFr1kYN
tWvHgKPP2kF2MrKlCKBeyVRv3g7ED0dqMJbgvXWzN2NqveFg/lO2ObSflokW2pd8
sRZM3JQbPAihsAPWGjiapnPWlsDUIpT42Wq76fAzLUMO1mV7Y3dLiFEuEPqNvFIW
W/KbmXyJZmgrGWon/c3vhZ1w6YvldYDecA1JM3kyE1baKLinZsUdPGzGfXY2Pm79
TKMpzUFCfvEwhVCepwweMcHY5uloMYfIybloFJVq2BuBDyirZ8yJnhSxMdGCnMfj
PGSWOZRZtdxAswUPslTnM9YSWnqzn1JbntODIFa0aCa1yAXsApGepYYCjLy3bMEd
0qPE3tuESLWaden8cJJJxGW5izI53Wna09ntKjrZTPIlQ/8DMouucLLuzNeJsLAl
BPZuY2CYLT6nsg0WrVNwU8ykW9H2HamIzO1wQG8B3urVrSiS6sai88x1BzssHh5c
uQ+TrhajraeexSdUNq/2IgyZ1ilU9aR6Dq9nPEl6ucCrGFLMsL9VXuYJG9Q5m1gK
NGZqNXyPx5qqS8OlVmfMsXhbqhHprVznOE/X7XvvyVGbvHCySB+oEMAw5A4Tcdgs
8ibjBmMC5Dbkuyr73HsmmmY1XpMcT4MvZh1RZaGC/xrKmLr3FNoIP7VY8+/s10Sv
xbgznfiL+g8gBDi1eVjaRYWwx5Mhc9sUeiy9WcylpmJ+1PWFBZESAybaDLQL3uJQ
MhMsFnUSlzVoT6Rf42PlbdwD6Va3BsbI1dnbPnqzyYUFWGpul75uLG45fCUdmTQ6
QNXAxhKtPLoXupNmsadrYx03pOJ4SKWz/InrDp/eCVECs/pFL1ENooheLaqGD2mv
L8sNSvxMvjzBqJU4Tz4dJgwVhITls8h8hGLwrKG3Fg3E3tEem3for5Ove9rN5G/T
yIYR05ZanGg3yK8C0a/hcskmT5NlBq/iLblzzsFHc3J7Bg15lES69EJVAiWkfpaU
EEPuMvQJPAXTVN8TaroBFJNI2qZBylztHrtOcXqE5vKSIPBxU9jt6ydmu5hDF/OP
39TCEjR3n2+kYrxNBUnWZE8p9gtA/93ocm/XcodfxG+hq2/bHE/bH7lZqLQWeC4P
xZtB0UVjPQWI27LbZ4V3Onhl0DNFCD8bzAQHJ6zVdRdKc4S8jBbX/eoIVshyWnnG
YTugpBKwLiVcGrMFaxG7iPloB82ZlvDUAeOEXw85ESt9bhXfTCaGzzwAKMgQKbjV
msQ8pqxJXUDSdtv1PtTlnTJM4hDnL2giF7OPshVkdgeMY6JiBRwnGktFj23Vzy2i
LBs6mo7ny8fUk+AJnZ7pGT4KDWB8YCQQa/r6UhOdbtLLBZAZD38CxLemiZ8PEDmN
yvQHzHpMvEJybVVrEJM4eQM4u+GSaqzedCQ3v2kXFF8bRVGHZX2N76GnRe9c1p6p
81/sU1pTuROHRKh9Olk4PEX2C2Pc0GSq8XglaPPPwOXTHH+FMb02Jf8PFKR79hVs
HACbYAKz6P2E/rj7DymBejTr/DhVsa66uMFwhxRI2x2Pf2y088mcdM5JkiukK/j2
5ODibn4RfPA+u8jpqydxSiHhr4Stfv9PlvItToFRKbF32+lxRiNVYh242VPr6zK3
HnhTTcWv2AV65SRcbd/3UxjryB4ioy5z5KgDVEPaIaxc6RmZsxPXK05QpMUtjJL8
32T1jFGXffPoCEcqDgZOFOYlb/al3spytQu+5GETchmtIHTc8m+Y2byHS6t7iulK
cof8As4wERDvihNyaSvesyu6Id2uNLPfC1K6jbE88GCz4DEnmT/1JqDxa8QT9U5K
gQ5t2OZjETuFGtUstg4U+fE0cXmZlAK2TIjQoJpSYs3MUSh+0jMOxzI8D4FDkLei
JZ5x4mmjgQs3TWMdPZV4/V2K+lZiNtvlChdnOm+BaOJQRHIRf5BRKLQUVmDoZx/f
rTYSQiXLRKZiRuWVJLWJ1THEzTaczkYQaio0Pu5TaR4sGXCBWVWY/4ZUN6ZneGYX
k1GjcxkS5/YQpMmTXE8Ap5c/0D0Ko9Tbpy/X5IAjVRoR8Mk9h0IWmNl9J3CjijLy
6Z/1ifMMjR9keve6FKzIihnrGjvNBn8hyfQbNWnCw01ErGwdzBRFLMQUGIUpuyGt
riJWkbSP9VtoIE1kwNmkOttdN/nhlLCkUjGLsHkNq9X1wruSY1KTOty8HqRDNelM
wF/9A32q3FuKMgjqUpcuHgpMYYlay2rFHP2rmX7EJMrMMzQ05OP0fJIEnRViAS4w
2N7gsqFMZJChFpQOjm4dnMLRv5mw1YZFB0QIt/fmzSCZd8kBaVGyf6Vg0ybB1w4w
jepAXthRvzP3SauM0LWFQ75H0EUG7p/A3XKCpy74grMUMyIIMrnzvNOJt5dSArVm
yryPIfv8yUlirMJrEg90+TfPa12x77kx6e51tGHLNm1sb9QO5TlPIx/HebL4UqII
VlXJgrsCE6US71mjPr1AicL1aEcoW1MOd2wD20QT6MeMI2j6fc2R0QrMZJw19uYd
UGYmtctnnHs9OTDcchhKzmRlKcdy5A/vZgf3oaR/oxJaj7EbQQBCzAtdyiGNpnXw
jq5JF6iaZYeSjaOdLqKcgMWNSrgCNOnPwXL0bdoI3po1oOFphQ9l7coZ8N4QRIEN
TrX9gfICNQphJjJjoD5raHgRHicJRjw/KaFKlb0NvX+3CbphSY+ldbT5zW6e9DO5
7dLw78lmO4cV15iOeNX44Vw84Sf3VJTDFJD3b4fc+7/qyT/m7gUVZ05pldK+pRac
3KAZcj+BByoD9reuorc9qycjJZdMT9m+HqFCjNR5AbJNIIWn+gSZ5HsxNHaRCNu5
O82vnoJMBjNTHIqtUP9R0lbsDuoPrgVtfN4GoQkXE+yV7xLnpwiY1csrrtEB5h7w
vLjbzkocsygatpC0LqA9czKmCiQqbRHuHFSLMOSAyPkeiKxOrTVAmbhi1hMcYF2M
1WFA6ik6ues9T5OjyELNMr9A0FB748aL+kvxv3ztZOBfQc8jyI05YY7ARGYCJhUQ
IEIBvbrm46hRcyt6URJfyUUKDrgEruBS+yHBta2Py1fC3RBFDU8GNNhZ7v1KtSDJ
hrH+y0+KGHNQIaMwFXoL0eX4EoGotL/rhWZ3Ka631rMbkD1oiPB1nreEUDvWiXo6
vOQXQwkS9GE9niVoNGTjJhO3eqqHco3WMMltUtgV5lOAGuurr6VkhANFo/jvr3YL
Hv/MoN+xIOBK7DMknI8UWsp3eTHH3hBirxc79j6xdvlgTiEL3gq+qwpkev7O7ayd
dhyGCOOP4qYsTXneJqHeTjvu2Luxr0USUaZkrGlWspunojHgfQmXV1WrrhL2a5o9
HdEl5dNp9dHTwxoJi4CuXXVkJYAFJLvnQhdvekknpqcZrDsdpmEnLZ1vzuNfNkD6
NDGmChhVrys6g9WK43QGWR3gIeR9LcrXMe+p89rH2FaOnRYYoR2irsrq4dsGMCgj
C9vmdAo/ZJZhWZ2cS4h2XVKCxrxgOfrh/tWr+fML+xIotwH6wZ5wKokHaKVDWp+k
zMx7oEmizReKH+hE1pXkkJde8LmbBP+1QizcRQgVwIYVF79nWpPb7rFxYBb4NT2I
8b/HYupLxHyYGt4bFqT6ADEVj5Dbd0J0RkOMv9AI7BRUnsh4tjRPBAUDLnGBq6p2
7a4HGlpt97i+7blymRgHHwbOf2IfIFd6/HUO4B0I9J6MB2W/xkPOzOPW90wxnHu1
zR/F6G00VKXEqfUKJSmddj16PcdTSuAMMc0sRNiqtwBKAm9K3n4k92tcAtiAFXla
DGuMd9feCylWxJY2tpFvA2JPJwf06m+RI+jyVJ024LEEHNZlV3aJffDTZvMt3teV
b8p3oL+5m+pFye57U7dyMND2mElIt31CH0g2PmZwgHc1+46obyGqj4Nhao0bWqK4
S6xIhj3sd2p2SZxj4gIRubhaAx7da1YhQojHoRDsmXKjlrukm9z0umtqzDV499v+
qp2Uetaegj7NuPh0s0uBy1biOzOFRWdqbtKmxvdGAHxRFNCkRF6JNx8ZH5Lx5rBT
ub9cjjr2vVAQ/cnzIjpGI8Dy5iwJsELBZgDyMEKXNhVKXq+jN1tMBCBbSNDnKZbb
B5E4NU25KIHKLEpC3fTLjZCeWpJIgLCsposOYYaPfTmnH2TCdNb4MDw6MjwomXKJ
/oaWlIXNbv1TdWGcRsBlvM9gJa1aFOKY3tBpWtehWnsTdUaNOzqBdC2/0ve24Pbh
popZxaPcBvl51dHi7CR6ezTLl2cdU7ObpcuJxpB2FGZwNk3P+HyOlBxifszTWWWz
m5KqzcvtUZZ/spWQy2n1Us2q5GVKQ0CZTh4cJjyFjVAhruSKbVboyz686b15diE8
wtD6M817CnYSADiEqvM+qkyO7lUX/RQke5un6EY6TRoE4AvaG3WoJnba9KjhfF5t
bpsWGPuaWLeJh59PT6DcCnvvLi+1tcoXvEVW3Us5AU/XQ8QdPDGf2fgQg5rsfJT/
Exc5CL+1BhFm6dA1fL2FT8MPlzz5WWsLrjwVHaEgI2aa+9Dv01dTuDaCEbWhwVfS
eB+ArqugF5VhIYE9ntt1383AfFRC4YrIAwq1rfWX3rmiygjQMTfqWXk6bq31CN0D
qwD/RwrJHmsDELVIgRwbdnGszHVJUN7JCD4SOZteHQ5q/oDERFWm4RsemjljRX8e
vOlZjdc/htoRgUSFXDBu96kWVimZwwUdNQFZxkS773kwGo7yLS0SKre9kYJIs5i3
EbtaAgiODzb5urYGglst8uzJ8vRmp7vrXED9vnGhSAgQgB+Vlw20kIxO/ycaeWcK
qTutsqNyiWBN0plmRgZDd5fzLOpLSDuPGS7zKdHneusQAiIWNy0YQ10hfhmMtwNe
buOfQlynjHjy25bNqlOI/8urk/58fJj0F9Q9y6CiEYMVmYOfz1DaxO09AWLAcI1L
FPEF2THbPq5mbovvvUr6HZcsO6+xQVmRjtSD0gtaCwH/a04FG/7aLu1JUoBxGnP9
QPeoR4jmMhXbMXzJLOv6Ky7/DEk1+4J779lLv57S/QvIJguvAft43ro8vVwymHO3
aLnXK7PVH8nFLTdg6XEmR6PkhUJe1iEZefWW/t89yAzrtqWsK4neqFCPLQgHb/rk
yykKS/kTcDNs0FmyGBrBqi6mKn1HonoOtnv7pnTuN2umKHxIt6Vfj3j/Fy7yxKSk
26q1xutzsSc65Bh4io+Q7MqzdDc+TPqIPL/SdhMeteaf0pI1j2/H0+7o0FeGgmLH
Km+0T2W3hMP08wDLjr8nhNTRzYt8ZJkgNFkIIVqY06TxQdcxPrbflON1lsBUfpWp
h6usZ7es+bvnSB5oNqb2r6QtZY4gZd88WIEYN5WPK8bQT8PTxqvnLhz1O7TTeaW2
VLxrke4Qv5bvzk8JVZAHa9EdPfHZJeUE/x5pUXuRCAmOS0NaMBbDEMhUNljP8lIY
/maLDofww3flaD9ub/O2QNg7Qi7amWGjg6SMc95iNNI/rVPSD6KHrNtdwrg2BxPI
V4BM6QwPQnGInNiWNW4NaUZxqaaCuzUdrEGSOU3DydoCVnqtT8VwDRqe7o2o/ebX
4qn6ylIIsQuBHEm5nH2FgWj7DnksihKIg1ij3z2S3QHVLF2CPsoYxjrQXVLdDSDp
yUQgM/g/6mhfj/Vbvgcl1hZojpqHmo7tl91DH3rMc7o5Nkc4Jyng0UqYcyKGWaj1
HfS+PFH2XOB0FIr86Tu0XXCfM67HZIXIbvSwwz+/MhgcEJ26tG6wiymBSN2fSXaW
XkrQtiuUwOhyfJur0U4HOng2zN2Spox8SOeslZ+oo3dxvlkeq+5aNgwVt5562v/o
1vmeq8vAFVAE0EoLf82WPUAWcgCOIJ+MHD5jYt3ysN8hVfO/nwR4rpia369wakjU
ffwupbJNFiN7NS4hVB3byjWbAsELoBMlHNDv0qDvkM8AUXRjqBpAelyZ4I9Xh9JC
YLmAnonBSdIaSq+jt03ZmiW5KnADVkjLV2UelUyvH2ElgOMB/MroO9+4PLKGmkwv
QdtLbSgmgK3mtCtpDngG/k9K1ykmn7mkLRN5o6jnXflNYjhGpKVPdMIHiAAyj0Ak
nGOz4jf+tvzJy6XkYv4aJM/q8UZyokYx2dUDfrsQseiijErxooO47JdJtlcWEMzh
T5FIGthyV4khhN8e1jOk32M17Xc1bRY/8ODXBUtkJt45/nIC8YHiohCiQhxmbbxL
0VQZ+atLN0GkjNGFI+PJEg+kYN4Nuy46dqvQ72tfwkKb6yO051RzWmBNw2XMT2Kd
xX+AlXSx83FSgZN8U0avtEGDQC+NPuJW+wlyDdskC8YvmOQxG/azK0Fe0b1YqbDf
j3pTjHB6du7MTIQQVOCU27NglFQ3gubYnyMz5lbjkVM1sFqPmbRUCFJqFp/TXEGP
1uniPls6u4txUTvFxU8FGqjuQ6AfE4gXm1vwq+oXMWzGtuE6tuofFHXNWLZN2XPb
/mqyWkppi/gTTkKJ1QuCfBmWyJ536mfbaLYrf5cltzIzZcmtFVg89gD+SKIeWyFi
zPVlJKr6U0P+BXh4HJaKunoZv9BtFy3azmElVkIRzlkmaeescSDSFu/CYWC0fTOq
M4BFfL4/rHpS1NIumfg8kUt6uuz82tLV/qqiN/kIncPwyhAl0RHO5mn24q5I0y5y
/94yjPiFaHRdp5IDmdXjQJadgvMjZBGodlQEm9Rrg+Nuh05T22qlB8T9HaA5OsmJ
KrEHBpOCfD3/aCCKsw5ykkzOtoeJNbee7zK6FMjCyskRo1m/BlTlRyEHaAynTJ4q
ADGiDWsZpf/N1c/AO12o09psCU+KKqSGBeTppt9ZDyO6HGWx2bwbym2lFzUPPaLD
0sIyyWpLI2qt9mFi8iAwfQGe37dVXDFPDjic1bm5Qf+jF2XXqPEKMIYLRdKIVOKQ
0zbFRbUlFthRlK43YwuqZhrjQgDUcHAtE4skqO0JPmZJsfZS4G+TfDeZaj1TQCOe
1O4X/ZiWEpNbAtisV45MmuHhn28YHSixtqaUtOIwehqEwN+YCVQdDS3fXq+c54Io
1f5jklI4Fnfw8ldLYoJDF3NgAhc1y/eiMwpHaoi4D+p7LtAiH2vBnEledBA2CaDq
hzGFQYb7tlMmjbrt60pIBRw0RJavoWjikD0GDqkXdbtnP9p5PvKmHWh/Bju8K6+b
2bnYaYcxnaPZ7dccVwSegQ8EogZpY/OojDH2F4CYcvcQUlT1ON0++xzRxhx+CCb2
c3GQfjkRrHFjRtw7zZY3J/phYHsmgq06j4lEqe098GGlLWEkWGdmgDxzoQnc5z7o
GDzP0iqEjuPBMGs1XbAkS8xfqHGf2q1ZqpUfJWhZsk+EjVlL6ASaSYwHpngDSTVZ
T+39u3nHxcmcR6vPBBf18keNdY0BvbF8181CdDFdV8a32NsgV2e8nDaeDB7DwNuj
tjftDeFsSBRl6WNYZFgfn02tIjYlw3Z4rjH8YU26WoQMauXaxkB6NgnJuC1Vgqft
PLvN16SG6pSdKjGGp9qcDjNGbFhRoKpRhhhuIQM2lAD8lzQlK0oWeaj6LXaVmvGN
aGSgThdnqEsgmBNQ23Da+o6RGkntuRa8GFRGNzgG5byjNSqPh4FsioOGH7hxwb4t
idTlQig6aqXJ/93azxEKKingBmxDpec2t02dpYNy3uhSDeUfbF/u6uylZNLWSPC1
fMcJcIKOazMGiO5fMw1sFYHeZTbqdDIZI2jyFSL3VC0AF41wc8EgIg43v/QEa6vq
B/ul7pkxW/hSeexQCl70BfViTfZgCBR/XpYoM1kG6M/7MSlyEH8ai+K07VhXZ7nV
wiuKToWIfdq1JDV2HZK8rjTNtho6seUDhZUYwiFiQcRvINrk1Ifrqc9GyzTYTPLT
cpLrD0dANYjhYSUeUoPWPCxYvP6eTeJBS6bzF9PqikhNfOXxFQV6BxhsiIEPMzdp
cM0zOkLFk5GYeTGYDEaJl9x1nSnufoqYoRjO1cDGDPVK/F9cv6EVqp4Dl1RCCyNR
c7xEBGTBDkrBjy+CXvaU+UMZO5zV8vxnABq7DcCZeb8TGCiVapPKgTdhVRETTesB
gyw/2Zo79WUTJPg1HmQ+V5tgt1yzSM1ZNgaGqEgHMHfiIU7FiaM+y2yD5e+uBYiQ
viUJfW0oOWgFeKkcoWuZyIczvsC72smpNAiFSs7jO2o/9TIGveJnqKPgs/3vm+l/
tPJs1bN2fPX3CACYaexobiRMYxb4g7jdGdWSrkYw7r7Kb+TPje2wAgdygRK9XhMA
ByAtnFvdDgbA5XQElRB/pOH/XrwH0YwzC1CbewaR8pS54zHP50jNtdUiw3NFYqVl
K33D2+uV9+dEZO+YflhBNkZ2A+aCukDdZ3Cx/yW6etM9nYj+GHjswMs9CeTx/D5d
ToB+JiBNe531G12RMoabp5wj/pnVooOkeo871ensgUyqkVIBZRAyZSXBFZdmkz58
cMRrudTYqmpDvr3yBqpe6Og7nZ0zjaOlx0G6nwc3HWo38wmqt9vyUB0s3nGuCtIp
WOl05i1b9UtjRyjXcJ2DvNQyaJgAIHWUvf8rRFX+UrSM6FMypW6qxFyRoF5AEw8r
aYmjUYABhYXCHZjtzRQjZ+HJX/0ODt5PSc7tN9TZ78p9OiL/k+LiJkzr2jRzh1Jf
BnYXHe/d9bz1CKfIosPjMEZZadEW3e5tcdYh1fKcHwJsTe+tL2wHUaqdmjDVLN42
cTuhGOeQi5R4F7acOcI4/5CHafE3jokGAZyf25/llAnUjHgtBySlDQcBuDALWq5Y
fmLhB3iY5kxiZxT7QoonBHZ0TaKUQGS0ObudYQUw8faUNfjt/JNzD1pzWmgiT/NZ
0IiaTRrfn1/kB29tmS1SpeB8t+7os24h8NHd/1it0cAYeFlno0Xbr7D0thLqopAV
awilbh4c9Lq3oNL5ZBAxbmHtHs/Cu8IaFUBZt3A1G5bCkV/qmfBQZCUcNHoLb+yC
wwaB2/7KKE+xVTxHAZ7tdzBubJi8fFbudNtR5JML/w/lDwzBcPg9EzptlX6nQQix
SqB5hbQy+H4OqHQPOIMGGo25J88aVsPTFtpQ1lVBrmmm6siUbqLZP3xWMRZk+IeR
lbh6lwWmYMd+HJYO90t0S1v5XU+mRjHdLTeb/VLoea2fmRaUAQwEkqJjFjM1pJx8
9WV6rEoJngUYqw6ZqiF/vxDQv8UfyLSSJKPa8ozHo9fcP44lUmU3O729Os9XA375
mnjHlSrOXomcYc0Ujngq7Q9KSxLlgGZKo+Cl/7HswjFZKndsqaTteXr94eFcBEX9
Qpf6xpPp+ToeLmDjOzMo0Vke4RuBCTqiCwZIiug9Rfit6oQY9ufFjLCoueLOpdIE
NiWaKyDVqqYUD1nWId7nOp0sZCW1u6sMpadt/YsI1+JXEr57W9xN1vfy1eQfwQ1d
DJ8SIbHUQPrVoKEk0PPoXCepP23+38/oOLJdjtIvUZBm1S/XIWfkrtJ9ZNsvvtoQ
OXv5ahrNeVhS+mkkH+mrPR5Qa0t+IqjQoetgKnu2r7ArRlTb7bvFnofqxtY+BQDS
ecJx4wVRmN0a4Cyq8/Zbdl/BLgtNZ6U7P6/y9qQrPTFxR4vcAXNL7kMXohbLjH+z
LLzrbEOKsXW+ObqHsIHlYFJI8MlIJqDzaRw/CwU17CyznS6H/o/Q0EV/UvgOWspS
i/RKqVXbzONcfH0fPNtVNs13C+6vX1moLUQOnCOEPYDFXfEnUhuxENPLWZ4LaW+m
uaTmOIjJZOV+4vAg8WjxvGXXhizB4j8J+B9gKxlBu89067gzth0oGUnWRujAUr0V
jsAGXSjnU4igp0u2DcWcnI0bsrY4IGI5d42vbBNC7UCbY+3L9f+GIU+JO/BpuvP6
qOxiG5cyOFCdSiY6GhArQ75bJ5aiCnyCP5rkRajMsHmtvBNicBkBtgErgVu9/K2k
tDfGslbqyYbrsfQN7i210HlCyhSxwiYR0v+BjwFAM0hfL+yxsTG9fjSDlEfAbbZ0
+mOF0Itj+l4hfvtSPWfo38brVgS44wZKaKrbM9sM9DzaqpuGr/dDQpGigUycyV/e
NbyrrfvKL8CJX5jyM0EmfQVjbf+A3/xu5Y7NIi99X7/55lsKL5n8kFOoU9p0WzYo
aqGqi2/Ql4OyQHKDtsHP9RVN7bbM1z/ynuCGSq7SX9TgOOBz17gz3TwoMksRxDoo
xept9tOtcbsYpwwBSzaXBgz5+QbgEXl5U0I7ukvrAxqmiEY1uSo8jPslgu/KaPRn
dZQzb5OTeba4TXoXMyreT+FpJoFYwXyjta8NjxWlGWEkOTOZcyacRhv4Uc7rjUo3
YRcsbCNZqDn+xHXXlT94JZ87jy3gHcsg/dbsiYVH29ETylV6kYNTRHCafsQmmmvf
I1eyf0lBwQXD9dCDRKz5DQ2kT32ZGRCBmiGJbs7Kr57iM/2gDCDQM2pOwOMeG0k2
bZJ6nOCHu7n6KPA4TNPouISb90SnFLZDBPpNMKOjdBQhhY4gnkqnCyCd/q0kA9Zs
EQe+klrDKaFuMFLzQtL+O0e+bysAy0jCrHTHrGu+9GT+RLZlj68MR2HbAhN0/vDW
cM4CoaP+ywyBQCU/cw5qW7w7q2ew/HhGNfZIwfrA7kh9br4ePwZcL70fOuN0Tyfp
ec1nPuqxZSCXcCnVjcDSET9WpvtKRDKkmyDJMvipmHdaY8ptAmOLWC5IOwwsqLp8
1Ii0rlZxhUM3jCbemGm9mp3Ew5dpwY8FQmYTz6HMWGDIWQ3WLFDyrJGNTd9Q56VL
rNTxqM+rJcCJJgCNMufG5xJVWaIcuIzxOjQsk+QQCEXkazvIa6+vFI50g/8wH/o/
0sx3Ui4c1vSNBAjbSl1ebxIjt4fYIGpoiGgNbnJJkQthWtiHghQpWVlq5gxALCPT
Vr7FUAPGX03vvKSHGFyZXGsASHo7UhzUsuG75FPjxfHetHSuZCQMknjUF4YHEzbh
4HyRC5Q5x7FctI4tXMCSpu7VI9zRITmFg6Fle3wn8GlMjh5C9rV/oBWQZGmKe7Zg
ILDN+aKgv9itR7QunDN7C5kjjMkbNO8lbtGrXMRQHEWTXCsjuN+72YiLGqApXKg1
qpzIq+LjF9MmmAMddh+IADgsuNouxGl7HbF4TH6Ky7VFImaTDnzj4UMeStPEEMB5
hklmy0cn6kzVh2n3DHZtUWIWFyKY/0kikRxiagTvmY1RzWTHHYSWNfUWKvIOkpxO
0+3ZIwx3a3zxZGzVlzebwC9TDgwVAr8aAQR5hKBs+bzc4BNkBL3vwSUk5l/bVdtz
iubXEDnxYpKhKaIyrup1yXalVBQOfLyzUutL63P+McYSBznNhMxvbkmReHgl8IVd
KRiGSzAb3FRjQ+a6KpJpRd7WL2U18L+6bCdUdVQJ5P0hGHMXVqnw88vezWfScjMd
3za4ALj1kyocdoDz9hsn7K03lEEtXBgVvwxe3y5GQXRKDXmPqP/fTmxB0kaA/J1H
UiMZgOt6ga8g9NwkfqKNX25CPSgVYayjNSvTFY6dpLzJBNOPa88NBQHNlfB9Lhi+
RgeO6OBwI1NjXNYBqzrmbUB1FgR4aTfttlksPjQ+s43Vnvf9YpIPzijS5I2piLmE
9QpxB8xqgqUmjO/ibz98+6pBLEktdsl6oUrt7QwiqNTRsn4g+ZHCF/qdUAg8XOZG
S+UKGJkJSqt49B9OCBuKh7LtM93M0Fzv9Rd5FfHAOjcHE/KLwKWPIEymCgkqVWBH
44N4ZNbjwmvtY/t1bqJz2rwOgL4UTIJguDFf+0IKkLBtnj2IdNBNYsVtlJn3x1Pr
3wf3W9TzGV2Cbp7DszoFKnTAcl/rrCHLfyhz+FqCly2o8SSZDC1lMcG87wxJIjAc
XJtYBUiWAKbzjHpieYqdDt0NL5zrYktOHDMfpSdwOkiin+6nZHbh483A9aeo5rnp
OUlWxrxro6sKIOcsqeK6/io8MAidRFGQoqeHNvaE+Z0OEVXRq/vmXcTFM7qWcHTU
4P+jr+em8TlyAroCy/Glkh/utK21uuqrI6Bu9BocDgzUc95dbI0nf/6Yqax5KyNW
dcC20UTLFeuP0iW0QnVda6C3ly1PUghvK27BhCkHaai9BgFEaiEQll5QaKz43+vG
SXsHVWtP7/qsKROHTmbQLSbGffXBrLLoJpBNjauGSOMl9af26mt35+gm/yBV4IZ/
rgU1arRv1QniQqrpKYlW4pjKVB6sqIfcZZZRsQQWJBHebhrvuylXAtOoLdVCWIGj
MnOKqnbOU8qz3NkrKsIkJcyuV/Jl8XOxRiQ7em5iciPS2tW6mebKNdtLyaXeM/dG
tti2fGbyVQWoOKsY24Pl+DCVcPBEAX9odmYaAoMPKNhS00HlT7n/WXr3fH9Yzz2Q
xZA6Azulzj2RS1XGeegfFwde93G4B30GCvRldjEH1Ekp5kzfkJSfBvhst2V7LwCH
k2sEetCOZSBfa4mdkBW+qkzF3lO45JgpEWD2UfOITrTtDanMt1lDMzWs2D8FNJAt
dHlbMONskh/FKbJw4/X9O/qKNeRp28aw8ne3BDcUCv2+3MYN1e61ggrrEp3s1tr/
pmn3Bc1SbHoaC8HD+sMQ9SfISUyL1EGVSrl2VLwSM4AaYlPXARg+0KY8hUVdaf31
AbVtIxbzAWvA6mouRPZMt2IOJB9DXhW2Nf/G12dnQXaX5fbOWh4kYnp28wFO5Ndf
AiO0suBvCcb46W7UV6eGNr9BWbvPB64tvSvvchypHK7SPSF9t+Bii0kSgG8T7qxQ
0MqkV+0wtgfpJ6O3MnH5J0gBUBrdFJYT09v28AsDokNuYrV68nVhYKYBpIB4g9gR
VMCsQaqf8KJcmnOTb1rp5ORCta3ZynyWoaXcU4h4pBCymP0XfoNrjQX5WLsBf+M8
yZNflXUHyiKwwSi7QC1FUa/CC2PYYokRnxkhBw1rPU8Ptm00ME87aGCIWD/cT+jU
DBCaxHzOZxrKvz9emWNssxbGCSEJJqvkcLah+37ui4bB58oUBoedWQLdizcn/4hK
ezNaHrL0UxijQCyvPRtjivJbcPCF2h8HAYt2cKt4CQQ1UFhCCxaoQKfemzAX8F2A
3LNU11Oa8YIt/zzEhhwIzVIKgT00GrYRgeMpg3U/0KA2Q5LY870JlpPRvNPWh9mx
BCsUkZzJyL/EGbcDsJFz+0dLK02iQ75vJlrZkENWKVwTGJljL5XiWEwGyMfuqys3
z+yrTbaA0LEFaLx0o7vjBA2PvkXyQhIxanwMul3LDy6V+YCpMTa1sNEe+pSUBOQo
kKEVp5IcCuc6SVVvsQaMCPcL69BcZhJ+EZZd74quUA5/psSS2j/5hzFY3zyis8ba
24ujH89YuswnTtbyR5M6zX2jWs2mbi+gOzIwMEmRQBT9yW67wxBJnfe+36hcKs1k
kXvrnijncowB/vCFFmr+G5AbcOZ/0/Bfkpe6GTKNrT8esqChlqYK93kq9mzI7NKu
MgSpySBv+UBOXgfkBk2zl2RoM3cJyc6k2ydqURhhULZbClHnsU78WvPJRdWtfDSe
1GT+pp56wHWDigZFBdVkuxGyW6vt2SwQODa4I5/5yP/18EWqraJ2VEBgox0ONghR
PZ0khRhwGyYSRtrUOEHltJey/o8N8AIr0qI2CcxvDQT4Im4yLwLsCsn/zpkIMt6G
gSm9ASCJ9s2my3aDmnCT7aJjzO1C6sYpIgupQ9/AacA8RE/yYbNT/Hswk/ymlPOr
vdjZ7smw+REf+B+YGicwKhY38MfSP6sdQONordb5l1/cXSVBOp1pjdEyudVzk8Iu
lXa9oDSXYs7jrxPfT4UAwToeEtFTO7UCBoW5JjgZPIuhnx4ylwa/KkioiWMWPSt1
sJ2TjjCbFglLB7NraMCs+ia+VwDQJdpryPNPZL6e0axraQ97fBu63uG14ntSdsKG
uXAwgSFSAJM8UrVfPfUlFOvDTvLMAnSulmi0zNetvUoXB14D8uoF7Il6SOVfKvOL
aVc0KfIMiF6ncstunaTkon9wraVVxpuxaVjDNVIA+D5YsHXVli74llxa5KlcbRle
PyvlZv3bdCBXFaob4vjaAbeI0POoQu15vk3PGqK7nLAFchML2rXrUosQRWXpJyqg
OgnWfDpPTF4tZZj+etezns5vZeMdR8kRi8g+p8K0e0W9lcNC17sXFmp1eVEBNWtF
fEM71C1A9MMzJBAuZXvZsQWSbHa3OXF0ggccnbhxoKzA3UYyS+W4OCZ/oQihdRiW
rmItiV6GNwfDFgrHGHjf04dpuBGzX83LfkbME0Kn0GeWK5o5GDwFqjKojmoroAT1
xqQn90pKW/0hJbS1y2FmxEB3RhS2pIJhcxln7nD2ppRaLJVIBvIg/mceFY12SkDu
TmS1taSVmU3zH5q53ehYQU3sXRoFAsdNUMVfKrdFldPM74Z7TyYJbpiM/TGul+v4
RCv6Mx1gPVAkTnk+YhKtKupobx82mOd7rucC8YOvWIZMk+ebXMrxDSLeNElzmmTs
EixBSZ5U7HYuwdr2QwRRqSUAAN/R9C1yNWKjJ2FNJEYPC514LFrjj83yRjMHmnnH
g8R/ZRa1pglpwxHsQrUxgchSDdgY0jpCrN41VO6LotGFe7LVKr4P5Fc4wAoqKRFf
u7k6e4xTwvbUgw8kx6IPZ4CBykx6WcRXs5oK/RjVQBYtFLfVrrZiZ0SdZWRppd49
074gXWMRJhQaXyoDgNuWXb3W5ivwhvjZOR57d691NoT1MuGHJ6puQYg/Wh+FOj4k
dwvuV9Ti4r3PwjKuoobnqaxhzYBDcH9kh12McCdx+nlYS+UpQRfpR2odmffjHT86
/sCN1cbLrSqYUB83YAztOHM3dR3u459OzX/PgujwTb4tnZtXrk0BZo1hj9HAL23y
VdrGZHYy+NoHmhCprX29whbVs/EEhbIBP6v9hswXtkLc+yHQkO/QbgtVNfeEoVKl
qcZxBwseTBEZCGdmD5XLcN1Q+95QzMUToe9tXwNx2GZAZhVG7KqkpEg3HpPu+1ic
q6ybf1fUbeDav6q4cTTSwNudKyraM3KYAR5l/MGCzPvXoe6NAL8C96Iq7VvdLy3A
jLtdIXTiPqa0cYrpW8eKX/8AIZRTd8Bt1KlrCg2u639isAIVRm6B0WA5YMo0rAGb
d3g/eZq5fLY2w9xYxjrBvCs1fD7Q/LrMWpOi2+f98VwN41IwkujHZJT8SAhbIgLi
vmTJrtNdLiKEzho71UVskP2CI2G3DLMjLMkmACzz6XBYiNgIO/onQs6cifghHKNM
vtvjrO/CJq8J71VNMqCRBrPweWa3/9IBlwkc8y6HA2l6DKZk8Z/pVP2w+AHnJJwJ
s6VkEXztinjhuHHDYXMVCdJ3MeR8/Si1e/CaLxHN26NxYdeIZdGmtBHXJLVpRnfj
zBy/eCAjy52iD8kznet9D0xLVr6efVMr8PAGPkjNt5EGSJFw9G0fEm4UT+HH4Bko
Gbo9vBO521KUnUW04JCxq+0PVxn8ZhK1f8+PdeOyg4C2cS7yoDv79t6QeErHXbU8
aiggUA/iju6HhQQ/IsS6xwRuz5gIeNB6rMXJNvZe/h6bYYEuCxTcuTkPXFesIVfm
he5WaaIGWQeavuBkONvZPx3EezxM1v8Banwd06FgVCLNt04KK+KlQL4itVswUWhS
9wzxgTXj2FNtsmmrw1YU/AbU5No4aPSge34ECLH0+5Ga4FQ0xXr5D5LXssl8PLLT
vax+fsYMKiAw51512cnFk5jasI/0Pk8CX4hC8QqbkzIpW0hvnQOhnnozOq7Jz+HD
BX+s4p/2EnBH+Pl0tS9nTDuGoXFPVqwnLmE5ZxuZC8p2NMJ0zx4K9mE1kPxQh0NR
ZMzgnRttN+z5JtzkgIc08ROprVGEflKmZ9OMlVfCwqgdnIx1V3tYGnddz54kpAGT
YcxkdWsKYTgo28Z68fcYW6Y97RZMjkDIxsVS3Diu9MsT/B3Z9I+742Za/L2DCNzS
zeGrMk9iQw3WIgi2+irpLcpNY4BVMWzE5QUxPJqpWIZGhyNGFSiE25g+PKqbrAJi
PgVzhaqG4yf4yGvF6Qcww2inD28oycEfC6AlNL32tkPOek+Zkd+HqueRZpggGgqu
c5f7mPM5LOyUuLTJlt2eM1UCAGGrMpiV/RUDnsmysKY5E1fcpGQ5Ws+jwqjyTm3n
6nTiQbMaq1gLdJNTaZBkPZCNRINOAtMNgn1Py4aQB3XVgrXux3gxrqQA3OU59oRS
U38uYL1z6NVXFZ1w5wd1vNtUKvXJghuTTFlfsaqklP+IxJ8EJZvZ2dCJzrpYOYlY
tY5O9UH8rEnR9pzvolrcVL4GSQNbFoDbw6CnYlyZwvtIZG2yUw5hqlL8xt/JVOou
Pbj3lBJB+jznEI2b2DXkHnuFsvCPReeyjb34b4SSAWuhfHeSlJB8P/Okvw7cF5WE
sIQ8SiZtEd3RwCzlaX0xlNNzzGW1CghizYxxmtgqyuJyAwN5fclLOtRa8iV2xZGQ
/iV2QLXqJG3PfCJgkiEPFyJnzqba3MPBbeDKefjae7Vnu+CyM/51COrMkIcCUen6
Slh/KGxGSHOCt2Wai4lizAKRLAM2esIs/9T+NA3Z19FAksPhVXD6NOIDpuiAnBPl
lyILC3W5CwGZL5/FHwT18YaK3IBVxZjyL+sAxqBvAARqRcf5SAZYqEtCubSBSbD/
9pyIgqUT4TL/ZcsPv7kcCEmwK3To0fNE78miQsn7WU4qVLpXUQaIM1K1SmoIYiTP
Pe13Dq0yF65ZQBS96tA9CLejLZa8mLbvhJjqwrJVeHQu3A0+7O4jDh8ckZ3DkV/k
5QkO7Y5dQqfiEdY5Ksc747871L+kuJ2o16nzSY7nIvk4vSDZ64iguDqCkeCojfPB
ZrIBYocyoNOKx7gcPk+VSgJF1AK+LtFbsSuqUtDeOLjHW05D53oE8p/Ren+meeq4
ZNgnkI4DJgV4Qodh/8d3M6Pp3d7WOeG6UPej6FFxIYrNJk2cMMcLkmX6bGRr0g43
97pbcd87pnxAMmJ47MPUGteaHq6lzoPL/MrfqxVMevN8qrbJ+EtUbUUrM8N87d8A
Iz9Fy/wf70zaqXPe8mJpczShHktV9blIAKfUM8rtd2Akh1FWOYPEZPKDG/z3d0Zx
P1cbB6ZE5EzstNlB+wlqTv54GjD8zXEccWdoSw90ELKClZ5wbNkpN4Bn1DB9dllR
rAbmT9kFsMXuOSlV2w+Fb2dW4qorlzk137llj98A8T0j9FfXOk9rLv3bckeZ3Kco
61p/vvH2xHYp/EzpRpJlxb6hzsWUp+mhC7Qe1RQEQtzgixZa5Oe9XSxQSWzZ2ZnJ
Sw7iE12cCOyfyeYabWPNsaLFLJn/bT6XJc7d1k33w/kwcmKdEG2EDJIbE7xyvXJ3
E+wPj2yOIdaRtCdENsVknBHMT/wkUfP+GxjCMZ6i8C8CRZHbAryCk/uGfSR1AC6E
dPG3CCWs/NR7LCAxjRCv5GHTVM33jC6q2ARInZ2DDNEzsOu4JQD8Ig/7eLET8W3v
h+oEs6tg+TrfOezUz3b/Vv5ABvH39LInG9wMZnXj2zKXVW/y0OYSAPM4kxkUg8zm
WTiY2hjCtdtX1zjqTLvk9dCUSC+EA92vjknOYt1VGo4Xi4gzfZ7zolWf58V6Db2N
fh7TCMnyVh1UxVVYLmc62rB2Hazl/TwINOilMojySeFf8OcxSIYXfqIaOekCQCFu
V1HYP0QJ1n7WFmTAJZpUyCzjPvww9MNWTUBGqzqrvUG/pFrbwC19xcJuW1OgMAEK
3L3MB7vqQ3Cmr3OSFA36iXOim8Iesm8BR1ByX9tTPZWpjBTNP+GvgiMuxzgD7DqN
3APZ9ebX/GGGKMUrK4jSyF+3bs2ve6JL17OnimIjHIMh7fgMvz3GagXUt9Z0nscA
eXOQo3gvfZZqIJFUPqi3iSMaImuCzBBvAJ2rL4iBreN7mONISSPAS6EbO5IvHj/e
cVeIz0veuin1UasvVrKWyj7pP/KUN8RP/9dE84OR44vdczwFkmLrz1DEwp7cWO6I
Xb+S6ihJ3++26hDPp7U8fEVbtaG5LSVzsL0RKJuB3RJpYkl+EqQDTHxqSbiA8CWy
tIOrnRKYzFxoO24GaWLUudOrfJZaC5PssBevH6S6cdnr/UH9KhadPbDw6n7KYboD
s/haj3lTzcb7mgW3NecIrApng/2XXj9kpa6jM1Ka5wUUTuLdHcXaCnd9cMzaDUxx
fUump2IsuhEylCDD9yib+DgJ6S5ru35kTfIupj5NQ4/vZK4IdN6bDiNhWVFjBdZT
6T1eXIPSvbPN/XKFTMwLWLwxVa5XUojjZQy/GwNhI4q6aZ04PbFk/xWAqqsy2Op2
1tAb0NEqli/Y9sM8Yuz7ir1XyScYhkT2hKfJanSvzZjPpR3dHS2VWouzpYm4Oaxj
Qhd6VVviHuIhOxTGaKd5wHvUdOOdRroTaAB/O5gWWU99i9j1AbudzM+0afg7kmG3
e7zRXzDw3wOrRiRpx2zJYKI4KgYYsket50DNkGj0b9jomaUgvbFGlbY0cRvJ4cfj
JQJyVmbdixhvQhsS6zDrJfdvjNlWrvWIt9Qxotun7zeKbiPqQB0fQpDQYa+eWFm1
CQSa04Xw9JgFxn85AprYJqn13UjbZA9OsCYsX57qECFIyVhXKscqcVnacfCNHZyU
r7bER6Yq8id1pxLMVybEe+z0j83OEq3T7/TO4GL/pAbE66KKQuBXtA08mzhSdC+F
ZHVaNW8f4hEGpzSRzcUhERz7fBwz38r1f/BMcGX9KlsCMsnX9m1fWcBPkdrg/x9l
9O+oZBL/gHJmax5aHykCiYFy+9Lkn/WPNVgVyADC86dMTMwzCYOg7H9xLulsTRuy
6lKBtPwD+JA8R2dnOC9mZ8bmgrZpZCpLuLwSKsxPPr2ddDrcTwST4eLkfCwPHOz7
2P8nYoh5tTS0sO0D3Zg/vDJbtMnZtLvAXdUwL1VOSOf1TB0SO6HT+5rm05BYhuLu
Pq9TXsA+ekEOqFIc5L/t9bE5eE5o96C5Lk0cD9XjCWCEmx20oYMO89JfjAVbyvqk
XbeSWUrpMuX/XqwWEmOd7LFNGCvr+LrM9NJ4FBrytpo2PsXf926aSpEi4gey2Rza
AXZLHxyghEXyo3FD/pW7etbdvzLQQEZsp145brwr5HV+1W6/3wtiAOncuTE8BK7Q
aDpOWaq6Z+zawr/3HwW+7EgmrW8GNRXpD6Mj+1g8F7xrPOcrxsdEi4EFwBnDioKv
B67UxR2WmUSbvjKiCF1S4UwTOS6Emks53jDBwpTasSlQqWNASsCxJ3urlWSpVdQP
B/ZuYgoMno25kW9t9JxqoVhoQooabz09hmT9ChKtDdG8cGtl0xID6JvQLFqdrND+
ArGlpbQKfr/3mQ3e9O5uXFMoDPJzL9aimq2gFMRC/io6XTIkbPGi4ypG0e3Cha5k
RdMOtUU4t5hU06xriH6EuzJVyQUxStJuRCQvmqBHwB4zYOch1BWC05kimWh5MT5a
IQKw3qURx1MmaaVQFQ7ZvZ6w07CEORXGit87KN9W10Xx0/r11xPk0uJqLw2Liznq
RjVglWJXSTwxQlu9ZDcRdr1Qq/NMgThxhIejGcPETBFNL7HFxc53rc3S6GFanJ3/
+egv0aKw4TTQaNLcTUGD1laFnwSmgTFR5c4fiF6ACNkh70KESG15uCHD6u4mzkFZ
ddcOJfAfyZUQH+JNn4o6SSOwtMwUz/K3O5VenLzxIA3f9nEFLFAFZsu04JlCsByO
9hKQoZwG4cr0TKTNceFXaqXh+9KVd2cbCXpry59WAagGl9skyt+vJOR5aREV/oyF
lYeNjrAORtaXApRc+VWr+mh5vfMLpY9D9bv5ulJBZsI7ArqfKJz6ks4bcsPTXfiM
QfUNUdGCI+Wjt5K/Sh+qQkWwVnDtVb5xEhEQWyqJI9bohQamWZ0WTeZnOEUCTgLE
FLsyyi6NHqcm7KnvjYgarcVKfVyhSJ31Vmt8jjh155TTx3hj1ahK8+RVGAMp54e6
I1oKzqti4jv3Y0jmMAlIO21CowGW5Krta3sOSkT7I8cm/F5NB9wixFnJNIRztjKB
MTnE+A/8f1IMsJfoThVXaVj0hfkFi0dh/EecmcvQeF2Y5rAfUcoqFFpB2KnaqgVf
xkM/Ze35Hu3fM2jNbOKjsWvPqxkL4kDEau4uIpiLN7QHZhZ4VDQGNIXImEgahGrN
GnSKWSR+5rcaUnJvI6OtOMNzgxgZPNCZbmeb6MEVKc4saJIoLn+Z5aMnu9Zm1Z3j
El8nbShEPk6fdlAMDHlSOVRQiRCbXxuY/g5BwUOZ0KWeXb23R/v2SS1HKSFdXFHB
1DqaVQ+luhDSJcW4Kiquyk0Td03Dmp37QcEf8/3Pvw3FVuO08gbCD5rquyUBFW/3
jF2I/tvrsC2nsy4/8euAm0hCOx3GjUWuNu4x2GuYPGvtJd9Xso93fCm/51FZY211
5VmC+Fb+HZybTEvzLhniZXw5QmWC/tC7LJ3g7gAVYVT9C6EgzB3RAgMLmK1+bJnM
v9RA/k61yHHbojbAH1g+5L4qvJCSqVMAj3fh//hX52EjtDkHYGbQF3HAalHF17aI
fVlrQg2D2IE5Vc6jS7520GvMm1CgjZgw282+D3UjLiPS+yBhEmWSjtCi9wqcqlP0
+oa8jeSkqJdYyks8fLC1IEC+jsPr0JhYloAjKKdfEcgCOfSomc7lNB64jjrdV2wQ
7R9YdLh1cUW6P1gGC7csDa3Y49Bzp68DeFlcOJDXV/ygCZeOHyMRBWZwxPQ7G6dc
Lw9lTvq8N4BsaRQijNj3C5F4queDOxtzeqpnAPqaM1oumNAS9mZb183ydrBICP+S
n7LMicvoBW3nxASft60fdqkrUB0aKFbB8Of2l4A0LR+Q/OCMKggKZqUUOL3O+uPn
VUWjG/93KRRs3c2ndaJhyx0N/3YuYcq6nQn6PGTBQjLkrD3ScRbqhtz8eiDGb2EU
Y1CnA6Pmugn39agg3pCWN0JWFKdynVbYQsC8K+nfGxIAkNHb0QUVw28Ut4nvdz6I
6NnX0waiS4cabdSaBp7cjeyzqNw9enN39s/QRbxJD6jZAIt7uDh44vDQ1HjZoTcE
F1gW+kSY4Yu+tFeItPW6XPrdQmLdsRf4AKVJmvTEBLFdBYtu8isazxAOcZAi0yIQ
UG7Y16KwXRVleQPawFtSNOedxzwp2iujI/d8005zxjYJoEOMwCRTTvQ7TQe8yiwc
iZwPJGhoZ6EDLgvQZC/SFr2UiJP4CicdlZ2kic8jrwA13zq6aY6cR46lFFGUW6uU
u/DihdjnkuAPEDDko1mnKWE62PxSetUmT90Q3NuXzhL+Tn9Xk/s6XEnoAWLvD+Bh
uufoZITO8wHe8Czh39VMwfujG72AmaG9NtKkUIZztkyT7Fw14js9qfNF2JY806mH
cK1fMEsqMpA06hSQct64nkVlxNtreGysnb8p0Jpvvr2L5+7w9kk7vQK0rsyPqmY7
l+IrvDdMwg5cE9YnO302MZ55xRBwzoWpuwGEqKFZFQLMPAmXiOkU/Axyb+I71j44
p+Yhtr2gLRq6FCtg5k/wGvskSfUaR9n0EyDTH+2IYhEQ77XOw1p3J7PuMGpl7EAk
eoPytpJhbnFC+0ncU7XRy3qDe7lbA8VrKUtT37jH4a4sMDghAXT/QMUOgrdx0zDk
ohHVMGMCeqo0Q24h2rXW4j2zC08SddzDDae0DZgTAKEjz/FFn1l3UiMMI//15i3a
iwwwDJE8GQ11i7y0isOGpkWgAGgCSLO0fK32lILBdRF3CjkBfnRnEL7cLr3KRXbB
cf7xDafFF/wIGakK+RpWjpudyFWp3AVrUIgSxrO+C/0MRj/B8SPOZLpdh5x0B35S
WsszAYicTo0ANsF8/X5VKjFE/0trkYzoUFc4O7C+jXJvKdiBr4b7Dsd00lwVruvv
v0KzUXxHBmSNtkVvRl5kSqKzb8klFvLc+1atyh4Qv8q8oDAxMI2Uy/SyFg3uYCoR
0jHt2zHmCE+YGrEckHNphClfwNkQXKYt27ivEO4ZisywHjzF9ss/bxF9bzLfrs9i
3ZT87RoILKBx0VPrxc4zhxshPsBAP0iXp4HaI1kJws5JJR8MEc+lWX7ICRn9MIiO
itxDt78HncW0lt2u+KwfkocGquX/d3CGNT/aG2IVHGWDAiImStWDrb0lBX3faNh/
KmCMT7vkp2vldn69pGb1vTgum7Rxgi5xGaqkBBoCGISA9FGqzLCY/4C8YxWluXwb
ns/Fy5AnUwYUpfabN8vGA8DIhzqJpLJA6VEGfGoZA5UP0nSCztkEigIMQiELijLG
qLO8Sc+zU0EJpjEyChAAgHlyAniaZSXfXExjh8f5Jmd28rcKbdjqZImFz1OpvggM
V5F3iMP6jNzeTYlrPI46ntvWo7Ga03DEUDoO1KslcWXSgwI2zeWcRbDzSK/s79SP
isdLnj25rXwjkKSW2Mzz+zCuLjUUwU7IHWYv9dNa0Ka7ZCKQn2uj/O5GD97QR1ae
HYcpzUvpz8cuog9IlkieeGFnfH9jK3Vd396+YE9VkA1Zun+sJFnQpyGvFd1QMOMV
LNIhjzPEv4kPE4QqAPqqEUmM3+8lVy7d4Y1RZmnRatyKnXJjDwTb5dn/ah9f/wiO
d61aUvLXhfjC06p/k6C6rGAQUeFX3HYuHaCuN7E8KP5BfsLiB9cllri0U2RQnatu
rWduL/fBAXw/ee0AcjIIOml+6vofXREaMAeRQEb/YqiirlQYC5IMFO4hvgxS8Ntl
Fo3S3ThZYUfZwOG4GzCEKw9ClELFrEyY5WDyFaKFAZJV8Zw4k7WjJIuKfBqiov9/
g21Ut7Ic+29VmKi6OGNo/DKgbW8FVkH698SJHL1W7JwYrT+OR8HJUEMPXqONrGFQ
b4KSXXBejkvIWwq5ab67Pjy2fhPzcRDfs/HR4nA0N97VIX81ha5+ct01dQHAmqqC
lljuds/lmFJ8ffV3j30y0Rkj1GYtsLPpCzSwbepiV+xWx00EnR+b2v42brwvlQPE
+EEHhFVX9QNdgJo3QPeeNQSI+SMeJMKqwXOsDJc26XteLHlHs3nBm1K5vdSJY47Y
hkeP5xCZxLtrgqKMfimRlKVmQCIFYZgeTKb0wr3IRDUQTxkJGnebIb7pNXNowobz
1K1qtvNvMNZgJkr2xr1JbIvMP++Z9tb418aBI2WULsQxx4JYTHvh2u4xij4yrDOv
+lFf7hdXwvNDMJJC6TqSIn5qzPxlWgvQ0GZy0ca8lu6zfkK9PF6Z1ZN+0PJD+pCR
o+73+t348VAgM5aK1AMU31BeZijoxuKCdfwTri2cPM3eCVv5u82EB/0oJU6XCkpC
odD1FbqRo+ZGkRzbmg5NP9jR1/aR354tArV/cxwxJBEF97DznMoEBBk9K13eSo2U
olRuqvqxWPqCxK15QjcXGunUEMKBAjk0SIRYMq7pBqLpLwsKvhAs56Ei4hZYSFr3
tKKno6EakZjnnIupcYH2zARY89s+apdhZ+x4zPq9QpjxEHaptOUbQH3mtRo/Hr5Y
VugMAco/EscEzTzRcr6ugy9yXh0GcF4mgdD5P2ywzb0Bx1lxhzjW9wmS//WPFigG
NLEiWgXQrwlpstkQq5UocXNBNChqt6K4zp/4IApSA+K6dmaNHg9hTCqLv4mzdWpj
DgTjb6Wy6Q/ijNOKTVtoBIlF1x5Kt2UjIl3XjLw+uMJWAllu2gZDJAXXC9oXq5FM
WNwPcvqyvAs0D/qXAqlDYyh2TCnSvVR/QfU0F7lyS2Is/wwaIyi01OmIbChDmOLY
AG51spxX2QH2IEeegfGirvemM13uYSw5dweIu6lWfRcYzc06k+Ne7oGw+YB7y1BH
Krl0B5tWegaqP687xAUQnxUrJGcGDX/4i56AxCHPtPMiefFX6hRyP7dQyAsMwOWB
g1KIm4wO84m8G7AwYNqw1trH+yyQHsg8D/3wpNU7Jl21824nHnAYDWAaldcxlgWr
Rio3bIsz5m7NaFv3a2aXip/LL3CvhaJh0Z6Q3XooVtuUU7eQ+BUKDgHGT0hrHped
AHUAj72qJSJ3wuGAXWPe7GOOFD7nQ3PWc89Ny2zjcsAU+J65pbPL9cSKTkI2c14v
UaKjBV7IfaIVaqYqRy5tcLOcqwLoWB1V8K2tx+2ebI00oE3PQe1+0B546JrGmWEj
B3bX9jkXigTwb6VXgqwM4tCUZmQFnZlVzqlWQ3Nz54k2/emMJxX6LZWBLkp9o+1G
xXNaz7LuuMUEXPbCy8OqdLZoZgBN/UT0mD5ZP5TVW6Hd0F7VkyHpuCt5fz9J4wQr
cYHqACui0JNJwDmCNBl7LcYQ6RzFVAponWCmZJRrPH67iaVipkaY71UJfK+DYNWl
iSy/wNWQ7Q7yZ/ijZSuFpna2JbiBaK402d5e9woG2J93tzOFg9cgD1gUNqcw6HeQ
s0ZaiRwENBglMzXtNijp8HyOD7plM277Xb8rkZBRLxLkR/IcJq3dBye2AFyuxBn2
boJyS0rendDJKS/OoGGkpl62KcYpg9joL9f4GbswzrCEoGNzixXcUqH7EQvM0Mux
P8Z3BKBKcHcTZSvmyt7xA5XXnNnCRdkpePCOx4t6TS87SAQgoZ1N/i1aACcOkNfB
uMwzAYP0t6luM1blhHnH7E4OCLwhD4QVhhPtMekP5d+VBNi2Gaap1jre7B7Nyfcj
Jby2oCD/3RauQr60aluDTEXdxbovp9BJ2VelnfqQEl6muJEXVqMZU3ju6ByKrIl0
2J3zce4DJe0zsMYNTZrfPFJRcVoJH3Dvi2i1cpxCZ7jP1DU28sKp23LyfgmvMw6+
8QanWB9ks6SRR7W0i8RauhwZcsimoRPHbdXOTnJCvgcu/5szGIWZjCjNncP9+1d4
pRlgG+Lw+1rdIHHQflfTOuqUXkQSvrk7tcH7vamuiR1e8BNkhQokeDx8KkrqFGWu
JV6zVLRHEc/3AaJe1YuRsgPqrxRov4M3ivcP9BzIU0Li3SYxyfmEQqzMc6HiAdh7
f5Ib9ssOPHftzs43e1zHnWtkes1zOkQbRz229hleO0/lh2Roch50tPyz7tLRDj6k
HuMUmiLea5AEbmFX5oZHfqyjOB+ykqXHj3LS9AZAIEw5Y+67kLqpBlUQTuiRtKGX
Nwu8v++48cScEWT+Bs+oWCYEwL1VZJNxKVJDkH/YrXXlKaCUcTS21LuDU8HqJkk7
bWnNItqjDPhgM1TEYG8AFd4wNSWfTQGb6fmrVe516VfQXxeTc9MWsKYIGpR5D6NM
KghfRaR1KKc9dBXM5IcTdfgD/1QPYaNyOEJ/+kXYIi5J7hhd5a9QcK+iB/m+IzKe
pRsUFmCFOCO73L1qic1CmXPf+S2ewfKqAYo62siNrZpM/yHrB6INvBd4H7/yxvUS
nGPaXWLLx57B+xJ9R8+gPAe7VI7ML19XxdV/QC7bs3fX9Oh4K4GefkbVh3Vg4PeP
36UlE6HgWmVvcgNhQHCPhbjhqcHr9nZ16UKb5wESOD4hsVuTysoNV5xl1jEZw9T5
+1wbavWm1dyn22W3sXLWnjjVXOMT4qcQUFZsEZqRkbok6KT3m39U/d0HV1aMckqR
ShyHcVL9eOXqiuREQKDkTTjbI8X64gXWfRq2jVz6rm9BclPrE08KelCbhOMhd79D
leZWY6io7omzQAcSysVyAIHR+iZdMZYI5H9e5AEiAb5s6Gu5u6MJidB1W6nTlO/M
5ZC+x+bnjOH6mWKvsVQ7DBOvUMpfch/7WZx8+zb3Or8pV5CeK9t5RlIaUuIQPA5S
a5NelkQ6yAzh4G0p4inYDzF/zD2OYl9AKZTzJ+YDdROqaLciWqsHP47Nmf53t7Ry
OytWIFpShwBOvsw/8WCeU6pHBfoG+Od97pkdMm9epyiiUAU+qVMdhgPas1cm8cBL
UiXxwosJRi++ze1Rtr6RI2fHLbyoTaUrCVv+iY9+bUtEtt4hOsUXA2w+EK3t923f
lZdz5id2rh8JKnLS7t7DyD1vo9E8jyeUGya51i3Lc/DXY2yNKeDm/OWdYhf/28TQ
Cv0n72BpEiFOycID2SAIruTJkYfLlnDj8nYeNkHGKxrZIjxWhqlWeWdY9Qv0V3mN
f+j9KThsjhCw1646+w6tqApqQpoHP9rWUe6/JGJc9UDEansX2hWlsuRMWyDeJwGz
q2qIElYYkW42BOfX6hsK8JBU947YP7MFxbd6TN7BQvuoCd+CFO23pNOw91GnOChB
rKDdNBuDiM112atf0G3JIcjx9BL2Ehgp4I35hC2iaW3U+2JAkWNm+qkqAFPf2Gfo
2C/nVcXtELhhRLGT0NYN+fpjkVGPrY7hTmEUtRE3jnA1qm7unrkd2yLhpzEetZiG
7GOswF2RLxA0gEQU6yr4OT5oFAF5QdGbbcrw29mLDcprSTP4wW7AcpwFMGASzdHm
/OU03/8YjTBX2o8mhcnQ00DWElSF7LugYgEMMcRrfukz1FxsdJ2w4tkMkVHwPHEN
gVldjTHQevncV8i2u9FQLH3t55U6kft5j1IsKWZ3D9JRfOM71oSgfrl2vpsYdua5
uB/0w+GHgvcyyMMIuRnL1X3S3TUcw3IAYDg+kICOVcMfG9FJ7RJZTC8rmPtUNpVs
+e3b08HwD+5K1atWs9zg9VpbhcP84sXuBxv11ZCFn+RuFoG3abRgYs+ll5CDoRx6
nozzAeBBA91Ann43c5RmP8InB5NR/H1e+pyeJCfTBSO9k3Xg4mxQS1qoB6JI7rdd
L+cg7rjDWNVFQzDy2wCk2NVH4a8G70iFeJ6oCYFRhCIYVMp0A4kgaFN7dQKxQpC0
c+uVzo/AxDKDsEZBv5gS/tm2xXGVwEV92hWl1Rq/mC7W9ujM47blTIZg0hqhedp9
+1Z1bQPkdLeqzOELMl/NXsplUukKtWYUN9xAC4mDhyMmeZKP0A79TvidFVKdtQdq
O/MELXdcKwPvqyGn38puLWzU8erbozB5bhfEBWHSs6c5re5TRN8G19Xe5kpjCA0W
JOvcPvAy5MlKlDj+h/xMidh0NdGpLpEDa1CJ4uyV/9LiXohENVn21AGciO8KWIpF
tgz6n25FUh97xlDgL5y5CIP7duhyEGRYyShf3/aNj4Wi8pntmF+CHC5g6V0pbwuZ
vqbLNFAT4T65dq8CtvIIfhAJjP9UAaYQx5v59EdNhYcw6RmBTvfb5T4rKK9720aU
RgbQQCc9qtv5+3U954Ym9Ull8P8pN42JsajVME1JYZem1C5oLKd1LWTbvlAo4Oc4
kTdfAF6pCmpPxXLgrktp04IeQayES7nhKsYrO4BQuEuYMbqW+wlnRqg1JRLOsmqY
q9eAKxlIQvCABZCEvDqim9x6UbHhzIuUcFfyCdagJvV+w7WC/qpRDgZOsypHIX2n
2ZVmP1qOeCx4+4A2YMAVAck1Cj/mgRDFG+0x2G41kSzL+chuQ4B41cCoYg+UoqLz
HB9lXZpk4jvElEKDeXrQ3sNzlpIIJPgHh03oeBhsMWN/FSlAGN/kf1edVra0gYEw
EDz3nnY1z3ZqgVLVJwKWDTpgfCRFltFvbLQF+VM3blEGn2R7iSwueo4lmpHc/xzV
dDw4NsoWuH1C/N7RS8byIy5s4I2S+pBbCxgo7cCOKgI3gKWKMu8pwFl+UUscr/+M
A+Fw1v41XTkNVpbJsEd2sn80XbbskiZcDVbecqR1ZwFsyWehmPgJ8Gg/l8PxF6ka
RYjXN1zrKtg9yyAN9TwxkKg71PFqNQ+grwsJoeXu1LdddMQ/kuBGlPLBACkyhbUi
fOLaXqiUBHO63VdiZf8sQshD/UAL+ZTopxAfOPJ7lwJc2Bpzo5fyr/SrVZRJK2sb
y1vbLNdOiE1u47AOjceA+F92hxIAwplY7fULiykUNX3R27/WIgxhEdUbQDhPqTGN
bIs84Ok1pVSfcQ65TAW6LJI5MX/lajZd7Zd2RS0kpBRgLenhMZU2nwX16ecDt28G
WlVRtCU2H+rTOGgu/8Zt+43i29bV7imHsiqVJ8gQ0gqBAJ/BcKIPyhaz3sHfVzAN
1QCoqAQRokXmflMxArXzthQqXO4f3GE+um6+9hwcjdrJ0ADdsPCZxgQHhmPgF7n9
TOswD0+YFBlzx6q8/wn/ZaQXFN/SY3EFt7zN+mdggZFqolV+SWC91P9jDDMBvxan
HoFROgVJVyz1gyfE/gestXxB67DDVBgETUiE6R5/F9+u6BRUtsQcrW7m904367m5
+HADasw+5DqtxhRr2pzSi9egWo+p5nsCcCZlCigk9W0hpMgwZ/HWyDZJRGP+AI9Y
yeRbGMr0Ym/t/EAH8y5l9MwzBivcLOmogAV8HYIBvuVFqb7NIcDD2W0XGxqRd/P1
bgNa3P1t1HlBq7Br1Ge3OPFc5r4lmnWEZbHOfEeoigvBWXvXcAfI0ONSxofKTTxs
S4HYuegmK6zkXeNMW3gXT80gur5bUS4N59GBK8Y0sIHDqFzQy22fL8hyf3punApR
wysfFIBOKxC4PWQTmKoWkQJjQQq/YL5R3DWtBYK4pv+C4Hy/pld0T7PkplFCvXS0
QpFlty+IPaVezwIYb4V0NJiVTrjOLIHHlSSeCumMejvXdydcrPsm6cnTNOdbOyQ7
udkL4IB7md+cATwN+hDb7lteDr2IBACD+KoSbSgcp6/zvpvSgacMXu9HkJR8nHgM
nTo3hQPljXArB8qTOlKS9aNW3IeGqa5sTbmts+WpY9RZDouALZMNfCwhO7gJATLH
2FkqbgI5+Td7YO1eI1uUbbswWZeGFlgFnhawr60u3w7/Ll9mPm/Hq2iwUTDu0NPu
fkZVytX4+tAJRoKzVc6eQOGSkeTZR16YqnYA+6GF8znHSUz3JV5HffguSIIQTMn4
cT2lGrVA2zqxS/FXnH7otI3TVq0HXrgSK2rfFxBUcnb/ZZtCnVnZ6NR7AXw6xoti
YMoKBzdaa/ySX72Ps25H3B9PjBOVOaw38A+ealmiYoIVwv3hY4KEuJ0C+kP8geIV
zfvuKjUrL7516NFE+YVUUCPUluhwjEOoGl7W6RfVSrXbOprqvt23ZI3uyHHyCZYL
dCXEaPjvbPA8L9WGfwL3D0k6X+c0DNpyTmxHd81zoeTduwBgkxMhFkYfU9ceOyet
CgfbL3MdkbZpaR3J/WSoHJCLyNJoi7nQDN+21Ek1s3Lv3eWnPzZ8oR8S2bMfMRhn
5QyLC7wWhOsizaTPE8CbjuRehAuBx8/+XUSVqtUh3pCW8F2D6upU1aQuRuC3vqPG
QjZMZiA5QhtiikEPhphdNAq85+7GIPFRz4ZS6tGfrprao06pKakmSCBrAbMZu3sJ
7q4I83mD5Skr+64ZBApstFQNbYwIi3latIFXWhrzfSAD1IS2BPjEvmz3cWWaO/tw
X+SxmSdtsG1pn3b81S/Bg6s5jJtCw1QflfIehfomqMmftT/3qpepP2BVmk1U9v4N
t+BCmJBr+V8o65L2Vy/RWuHPZFqluvgAjHR4OgLpC5nhgs+s7dEO6hQmJlvVBGkW
ECAWKQdgTVJfniHVUZKU5LxFoo7kIIdmjfH90eItsVOhhaqTIwdNh6vP5Ou9JE6s
uStYN0W+p8KWizS34icpQmcpjWtdDWDiRrs0pNcLJKSdLmgL0PplGWSGlRHiZ820
vvFlWbAmWlqIyF1VR0IdpwGCp25q4/lfhffG6mzOjGQ4WOPxJ6DJwkYy56ptmag/
IGsVHeTAP7AitHn4lBnLNHOSFjOxyfzZrqSR6UjoUi2xzC2VL1KmpPK8FZllH6st
22vGzpq2KaxpbHGtbjGFkh6XoB5NaNtMJY4GMgLYAI5CBTVxhqCL2M1IBuoMEI5Q
PFFqPHZYeHYp1UiIdhr/xaFXDTT8j53Yv+Xuu4Zbjx7onnS6fx0YrLccyod9AmE/
F63wEy3JbJYmQ0gNguwzczf1VNWSFSlEjhvl1+5emhgpuY5VS/VgUNtMSjlJV785
wWyAOxqnjylj0n7AyXWEgHwmCF0rbCded4aLIO8DMRf05lCDvY+EmG3pM6aiPvPg
1iHCLPhwrkZxMatrSnBR8AV5QxRVuwNWLrlcpd51HKzKS2V+tshqFfu284Ws6ZL5
0VFayL4KFXFl7+ozs5Yqn2I6K8Zl4Yn+Ql5eNPV0UtXm8gWLClgjebL3wejKELVQ
wFGnikWCKt36oob2FB1Y9rBziR1QSovYse/Ivk3m5MTNrswVJoXNB9kgv7hxeDF8
7p99PL6Ip39H1lTH4Mch/Go8Mh5+iO9UDMH5UebRfsAg8R4GF6MZN3FhmjePpJzZ
MQW4zKkWuC5eg/D7m9CXxUiiXmYTfNQjMgT8ehisGkf5FWpbXQxrSdcKz2kB/iWm
eKoeE9CnmPRjQpz/Wn6mfd9Z9nF1/z5eVJHovnwtDvc/744ZBiBJr1bvrRi81wcL
SLvtIT8epy/LuuU+QOrEVHthwOkQILs4GsvHyGZHKN8HXdjg0NVC8G+le0rMLfmH
qtJzVTEOSRgbt0Ahutlwyy6j2yYdgh/aQaHrcHc68GryUX3UTd95p8aFDO6+v1O8
PIW/haZ9uHFdahcsxgLaEYJ6XfoSE81beHaM7+rsKln8yh0cpy0XUYMDm2NYbpQm
qpJBeFfTgjEM4MGoUTARXVE7xqYrM6ZYQMPwOTfJYkRwT30Nw89Mr5UqjCGcX40T
Wgmqrs3TYTIob+bocb/1UXMPS1A1ERQQm8bo+u2d7o+cqlrrlfPmd1OxIJxAcC6T
EDEO9WYNd6a4vIo3JVwXCyiBwnt6MEiRIBuBYUMCwArPOi+D3unRzlDCe6PlK6HU
Ah8lv1Dy1qZZH13aI8L/po7wQq2fZ4M5QvANnxy0tKRLIVZw9uIZSHRLehGKGFf7
H1mL3ApMtSas1TvLpCAo86bkfhhN0YN4LCkR1pkZRBwfjJUQq+FPNDp0uLVzCyUn
s0dwCEiRJ6DpZ0vaTXpDdFh7F4uyCCKG/lOj6uIuaAsjWgOCkkpy/Jj6pw5B/McN
+JWH9QOevUVKIb1iLnn1P7kOmnN17tyOVBXCuDtxhjIPlM/86kz+/o+w7b5l2dmd
UkOWISLmHi0csGJANcVoUenL7FXP0kE7k+svuJYhZXNJLoYXQ+kQlPPgkm7XSeD8
xmTcypOBERAOgxFUtmjJjjbglPwZhaHv8KxbAnrtgc9dp5snD/1z6kxKCyYG9oyH
OzQpJVwuKm4j/wKv+lMGwKslr5fXFhIoKqiNsQ5nPel5NX/dR7/27SSJo5Llx5NJ
USohgqMbpLcF5xpTssM/ows0qh7MGAglsENXplwaVexSChF78uKp2GHJdC4v93Lp
gwL58ucWP4l2T6JqYEEZyxnobeoUWOVUPJRvJucMBnvu85KdCxoEpEXNQWHXUNRF
A9rVv/o3q8ssrT2rCY1ZvxCCNuipZfMC+sNZn/TldFLzLHpqQPXQC/23nI5iRsdp
D7sGsFc4arGfETL8NMuLN3OzcgSfB8doE08sZu8Uen2BNmhlgp1IfQOMw9xVUqWU
z9CgiFulIyWRKym7l0yRwNNMpKrITX+9ZVu5Pw8t9HVBnv0dK26o5P42etbjnr/x
aW1aAKbClvDg57m/ZNaRv/Mb3JVfLlAYOa3X0WROEn2sQqpvRNPpb4dDOw9fmS1j
pfOyxHps/0uL6JZNuNcWPJzZrS8SylOszFwCOjlV50YzUq5UkuxRmeigNkTvC6Bq
SJ9Wk9RXp7UR7uz/wyMpDPdZU6E4zRkGeR9bVzPxgzk47c1YSV4tFN6He6txJs8Q
zs4eSxxJ7M/kqdanxuILCR6Pp7AsX2wmFvG0BY+v/t1HwpJu9WzoYhlgJ2Bc7HWn
SMZj1jTakSXD3d5GJQZN9xRiiEVRcWnOWKmjFQf0bC/ABtWbfh5TlCOK/p+eWaTI
KkdStCzvk54+IjYYD9k5imb2jkUAlJsn+MoLTMbbTplWP4QS5Eo20EZV4er8LSqA
ug/JcCXANyCpkZrC24QlHLTABin9RNGmKIevI/GqM8CyID2KfP8LSvIvE/hrcVc+
wXfbgWqMjE3qU9t7zZqc9ZY3Sp+tZBNv5P9WwoCKbGROfVQiO5KBbT06tMdn3DRY
jOFSbTf9JVCXaWZOMOux8s+f8sH6UQJ75cQEPDBTvnOaRmXioEf5j4joEMLEDIf/
8tVThxK/7HP9OSqpaYCNCfUNB1SFzu80ZnR2YJy9+iA9+MqhTAZbaR+97+leF7SO
y0RjiiGh5QjR3gDuek371CoR7O98IbaG15PAZaYkHN6aQGgBiseJ23u4F2cYpjSQ
sHpkmYudh0FUJ29p8luAvX7/SbsQ8yrdcZT20c+1ZoOO+OCZT9neNdV6euv1v49n
Hky05fOUeeTyLAl2x34cUp0EozIgkDCQzeWESWGzC243Eij7m+DYNVYNXlcFsh6u
0V7AJBLQI455mtkF68XWkRBdtjwtweeZeGp/YMdtVhczAMdlwgiHRRadLy8blU2X
fzYHYNaQ+gHmysIrm2CwUcxDh5xAlGRn/54v8twSuONZBvM7meu7QFY5E2icNRdm
WNi+Hgugpw7LfhU91aSFORwwIIh2bRM3wb7yCWw05WRszu1JF9Mg91cxU+Rt/QbD
4Y3RyiVdr/tiguxF6V+yzKvVTSMjF2ath2TpdyHgP8CkyVwpLwGznbqFiH51Veb6
wyFGYB6As01n2VhY5xm7QZpONTtbNLDcFk+mh7xNJl3/jZ5D0zfMdd2HXLmcS1/M
EuO6RJ6dI7ztcWqA2NGQ09H29EhxdfCnRCw9nybVQLn5DKVPUOSNZw93En81p2xW
+UFZqmjS7f5vxVKfXWAvneKcyj8cXf+NvUrAxIo2jyh22hcxMHXkbFsnnbp/oEej
f21SjHzqoQUkehGyY96RuI8uX8qQ+2QOMwYpPaXGY4u0hkrYO+tFGf7SNJSEAcWK
n1CeGyguH+8uZCWHOugNQ4K7kkqT4hC7Wj9MSHnvxfie5VqHhooodXvHTXiqAwwy
4MQS4533Yrjj1kn5+IbGYq9RTPn1toKrjFZ0YdjIDMx/XpuHKJuoBk40NCgLImKB
SNVn/sKYY8SwAlJgLyaJmVmZfKSFHi+l6MQVUCgwf2wwEkpkC0bgGDMr+wIDNphI
YHYBPSMNNXxu5tDjXJtvE3O3ATg0+1lybPI4fGn+YcUpE8foItiLwP9+Qlim5Wg4
3I7sclus4wUwWPtiShpMI4jdbryeS11XhkVQ4xsiEkQZehuQmG7rjWxC1ApZii3O
6qbAc3hQ4imD2uOr7tnX4z9CgP2F1E3Z75ivPsDYZSATTjLebNH4B6Tz3P69fP5S
eb5h1l37YyAQsaeR6LjcBgvWX3AL/0GymggBPvEH3W5bECRv/RdlxoVnvYhn3UJ6
Ex+aVYZ/8MWzz2zesRXOAnfk3bbqEl/WcJ36lsZf0HR8TWPui54sjHXcd2d9pDVX
jGeRBMl3QxpNoYEkUjYaE+jFTFPWn/2MEIZem+DYhmaMoIctE7WjUYvs97tMg8Rt
PLZ572ZtkRjXvDFoWidebJ3OD/0uyokmr8g7tyebbofJn9iSddK3l/ejuduNDLAC
XrkYlyeb6R22597XywyayvcudPwA8WH+zFn1YqSY20nh5w1do8fCoqSNodh7MrZJ
dTMfgjxRS6rci7TfSAHTl5yx6uFvXeQwfSH30HKk+1rZQB4H7cZJmI84BlOVkf6D
NIQRFt8sGhJdIM7p+HHFvlCB4rsousdpFV9SC6tSPGNHySr/C0+pNDksKOSIrMc6
N9CprDrOP/X0+AF9f8XdBaqjSDD0axh/B9b2w0kq4aoJigN2eNnK3jJhqtSzJnpB
6F3qOEOhxbOxl9mn0TKv/2D4dNV0DRq/muMc78oS6ZG/F9mZdbr+aPo8I28RPjqv
NS+fdOU0rkELXH1uQHgWIggdcpkL3OO+gr1kn/Y+YO28znODkOed9MuzLb2cPrEx
3n7EngoatCHKAgRvnmFnhTBqmeIkrk6b3gmrACfpvr9eXVV4fbe14u3/818YYzXH
4ugSv6K519upm5+TjvfJqlVUcce38UuwKrzD7gDR2uWuTVbUmI3HQA4q1ke31jww
1B+f7VS7B+zgdccmdcwd04ybGeikDTPzpGx19emnlBZ99e02UPPiJAptIekTZgn2
QhdsvuJEJ1di2gGQk2FkZVNXlpq/QUUJzqgY6GSzH66066sHZd2vOJu5X5k+85c4
UubzPUpdzpibF+lOUglFZMlghS9TDzhSp6lsQRmxj4iP3QnJlM/ZFL51pVqAOvY2
e+aamHeCiZil4XTDCegANWywMeunYCae9sUv50A5jSXFNQoKaXi56pqPnFC4Ezr9
QWqv5r23mFAsJgB75wS4KtdgESzJc3Zy2WusQeeOTA/kYnvm2L+SSKV5yRYIFzEc
P5qyldzTK4ilN0Dy1O7P7A75mnNDJlzricL9Ou/a7tK4JK5p8aeFl2WjR5JZO/f6
K4lhX+D5kV5F9JH+sH0OeKUoEH0clVqa6fryBUZoQBC5chbxIHu4hvaQ+q/66FWQ
J3wyVtQT9KstV1cosF4aPBvEW9cqGAAND2Mwdidn5qJ+9HPSvru9e9AcEqpKXJQd
4JYmf/lEDA93Cr2xu8eZ7YU5FBXCILVphmg4Mtalb5YuWge2Nvkb7ebCl9x/epBO
zdtviSx9JyqVjKfn5u5ZtNk32P1nGUrwd7AU/A+KxVN86rKGmVQ+uffjG/EqvNAo
Tw9+qEhF7WUgBaxN1AK/trxlbCIXzm6JN/btGatESHgt7U4023rAB37yXLGkI7yJ
kf/xTWm5SrzbHWf2g/mJd1pLIlE8sxi47n2CjGifg9RaRVNk7mxmke7NM0fQ48nq
qg6ShSg40qVkatb2VzFHv/uzT8EdxuHxhTSlR9S2WayACqpDjywkmM6Gnq1YgrhM
rTCJ46BhHD8mE3ztwtMUIkr/+yp3l9woUCBPVaJYd7ioCBUhFEV22Md5r3C2o4Oe
CbKEqQKheeXm/KioRoX7q7epVkDePPAog5/pJrRkcPJKiO16w03wCbJZztnZC+Bv
1t/CZJfR4hrA1JqgnJAMJq3j1tLwDp2cCGYylz5JV3JlpbHBO3jTOHbnFt5PF10o
wHkjtZFnEZmq5s6Pckn3e99i/0DZEDAfCLnkQ35Da9AWKdpzQmDJjISqRx6RWNLD
82iPpQSKnXJ5HzHdJbGnAzdgpZKmSybebW2reTHMLtCbq3Sl+0tk5lWPOju8EvOA
mYJlwSPOpXJ2kqkznp3tgr4LnCO36X1WNPDVolY/YCzc0G5ZD2nnR79Am1bDOYV9
oulmfAATEO1fVXeHx+aQkdicxnzt21L9HvZQZlTIoigQUtRj96SbnyxrJ0Oyx+Ij
LeHMTbCXybJMOmk8yN65BI8zaSwtyfhmQPnHe29z8fwHmbPv4qUHAK0/GKmR+UQV
H1AzAzjFWSSwAr41zbRMGvhqzo4qM1T74p0d2SPEii7zeybFpyOrs7im/I/IOLmx
PwHfK+rXmFMok+Id25QjNU/IT17GA6TYyLc2gUi7b+pDSXuq+kr21rhOQw8t5gPV
xPNU//A1SasAOLYfTAeZ9CwvR2fyM/yVMrYcfplv0FOvwiS7WNC/RCEmF8WO0bgL
jKtTd74guhX1Cg0jGKhgfN0TFmlyF1cva76zmxKG0AUn7mrvMuPnkpuWo9ljMneL
CX6ISez+a2yFj84i0tTw7r3wrSn1GqYSePj/QaY62yKl4Kg8Qw0krQi+RRxExg1j
P9wUx71uXONvFVDKgagpnqGUMkiONhjj/TgPQAuclzyQFYvhn5oilhORb+jZP98+
3iMqiFztNJqEmT2O7Cb8z6VBNAR0+tYVctKyrtX0t4o7PubNslnZK+cfbkJjx92s
8alGXSKOHZB845CD3SVun7cKrA7AAjt+lnDZyNQHCf2gvBTtnvfjCmrHzUqnCZ/B
85ZbF1BpAC5xzV4UDwQ5L47NMDjUPnrc8CG29dYPFNWXrT1NMoCyuecNqVD7DBkm
SXnHrLH/a7mHlSov2akNlolwiKGuw7PEPFVyVCbIIVDdoSfhCvo+XLOxupktzYOo
GG2CuohpQYJ50HeXUZByIzNsWBaoHpSR7E2P7MNAPkYgbEWnjYsBFZUxJT5zXoQX
jadxwwb2bYgrexflYRUFYDoOoNe5DX/GPAvCVsWQSQqfxc0fGWxRcPT3ph+8ePrv
Q1jc5KXzJNqSiOYJDaZigdh0US021IQ8bAwN4ZoyomMOo5n5g37569AtPcTLwaxp
kDPK3dbrXgY8Zm+mT0S/+FP8P3oTpRs72kpV/Hws73Wxh9mH/ZaQVBP8yW8GRkGf
2yN0fR9SFCPvB0YoswVLh6bhq5+MsFkAW9FPrxIfl6X2wedHW/C8+/PEaB211vPQ
bMVteVpNZ7BzO4vZ4lSyPLkRoAfrJFRSsnlAzbXERietl7UPNXRo4/FAdBrm9uc9
qSI4oxvyCfgTxpDStZebm+yAEC1QXRzYNxeED4BePVD0RDXq3sZHJf7L+HqZ3rnh
w/GkNJYdu0DT75kd7RjDhso2msxKleVWLKSUKDfEIHYwqzs1mbKS+kXmEi6D9fG+
3hAzivyTMdBwxy0TkdHnDlDyS6AUiT4dQXT1+I8ctZ65MbaF48ANBtXIPsIitsHN
LQFa5t/parHxQTUyFaPqqnBTjCOjetH8aCHfEF1uH8WPjwskjY0/KDSrUvXnaP8D
7hVFblmVbEXFyjtgKg3nzkA78a1swl8oRGDkOe8WFxaYA7vpthm2HT6q7fnnyUa/
haq4rdcLrXM1avqvzngNPWyld0JlmYbJDIETonZs3VB4kgMnkjfcBgOYJ/mQSuni
LUtDX3cXw7k/9LTjewVkqvlBl+cc4SKxFNdr0PXmOei/hOyPWKeyIZq/rlug3mO1
vkhaIAJJI2vtus3viL+0ZKsKkei5wWnTAvidvWH4KQ6rTw1iu4ErRi6Ql9/3O1cQ
tZNHusDwU1WOYv+vwDtAVIGecwKhFEXbHohnTR0EDyV/kh7UWxKXXIAxI8zDOBCO
U9v6f97XGIKP9L4fdrrssYWLbrtblFQEhwxkgPuvsQf6RL0K8sdfkZEy1Lfq0J7E
ZRl65P7+KZyR55hRf8RbecwsMvveMw7wk2Bi1eOuiEjaQmVrFUIhQxoxDCJpYQIg
xsag97sLnAIi3pjMGKI3fuCXp2yPWynzsvmYSDFlTO92mPJCadj9ksMUuZ5kHl42
eMSLZC1jKLIRvB66sogUE0+JJhZPFqoMWg0C41NrJWRyb0F6z8Zbg7BqnRqCZaLh
Pgb7gpNpeFobVva+97eBDTg+Vubco3BGKhHYcB2wAEqumyhZgt7XAdHhddx9Mzed
hfsusFHwmbwAws2CP3lW2YNA3EBEmOMjQtedZN1vzWdfAiLfko73IEfNK1r+OuL3
6zNRu8Uzs+BwpRN+rKKirFg9mM+cpucqsJErKK74FI+kC1UEH7qCk9HEvZ9K1Vrj
vIWX9Vac6ViRuXdzJ3J+3jse26mF4YtQs27coijFyAkMi3EC38ST1fz7mis7ivdZ
onLbqT5T3JQo5OXX7xMUolFemYQQoiFQbJJjt/RSLcPTvKUVc34ldqU6Rp7rcNRt
ZA8hYV+kergGWwlxqzLEVkOqW3Kaf6WqpVezfx4rGEgJwEM03S7G63TzPHHOzzG+
XZ9fgZmzzN+dqQqQNGnRqFoYBS7EwKJGPMOz+T7pSn6EkoUyEWvJS5d8MBya/wpY
ZQuU+5F+Sb8DrpOReYaHlck9kQCET4RoZh8/nIY1S2ouwmGB0zm/W/52kQgwtVqu
JTFOTx4aT9gS2cytTqGbxYez88fHUxGNcFDe9p6Qd4e8ighDtbrxvJXz4WNixJ+h
cEfDD212H0eRaQ4xWutIiQC12YQlk7SbkZRIsA3DROfWVgjXMY3zOpKWWEBScHm5
VpCSYmm8vGbhYmpp0p41e5jgHATdrUlwu//T/CCxxJNUnGxZ9DP4zZaPjJWnQxZH
2eqega9I7OGskO3ij0dkKTTxru7hlepoh0Ihitg4UA1seATRlfS0MPfAhGNgK/1r
W0w9gFXIwEImOFGokej2xZ5cLsaPgpimqWturuHEhsYxQwAe+5C6moBcZeMrrz5/
ed/dUZlzia0nlNrbD59ssfFFD8yispZJAnRZqon+c5RsupqbHSc5spgiUM8mjZnp
eFNeX6qzqPcmi47lNa8doU45El3riY7k+9k2ENZ2InrZYpSiS6Dv9Mx/P8yEtbYx
a7unJPW7gf3B6DyC2Tur1P9SEev/Zuo5PbzzfwJ9D8tbzzbsUk5J7xQjPTwZu6RL
AKVQWPI0CNE9OwLmTvdkfPksER8QLsgEU7XlR8GQmpdLfgjBrpirpvBJGopFwf6/
zLbUzYL7c0gjxpI//3cJjiuIuu3YjbirIcE3Yyd/195IVZa93Z7tC7r0VBFk0ymh
S9WeH809rAcPcgkIvpQ962D+qANhNoLYZWv1pS/WQ1Ds6XSrvz+DnFCTKfrTEsrY
frDjQugV5KB3k2A8ns/WFk09xw+M85Iw5jzbMpvT2ZJ6ye5sSKOMS+S45fEaa/MK
w9C0F1PS3JBYJLdsJ1EZMlbILuVjVAKeFF5u1d3622JyJK9vicw2PkVtlqSwaLvx
+eBySiwN4UlFn76gnEiOWOEcoStK12z0CALOOeV48ua/I6RySf+/rwugVjiSQxny
7Kg7CqdhqzISTvkKM1qMdy+vXypkKAzIa9VUgVAcm3/KLZuT7zME14o2g5xzanFS
gWpdmNqTC92g3HWOGuGeQuHPZ+4ok273lXyTea4E69IrP3N3aivPkt2+dNv5AVTe
WyBciDaqmrIATJbpI4u+fglQ4krgNY8pWbiPHhmfM6YUzSEWI2aSqYuQ1KnTVrYW
JDBNWcMvZWW5TbBV1LZUWXydZPavwqyN4noP1/bo+PtdubsAsy3ZrWl1ExCq1S9J
prnjlRY/vd0QRPg2uZgU4oo9P1+2nCvKCfxqGs+JbrIwiwCl2Adn3a1Jve+QWmqE
mAAVbeYntv1aHuvCxgn4LLbgvl1KMxKenPgyKo+5sN1sk5gUcA9CoEiE3mg9yoAT
rlY4aXMWPBIUMnrOAyeGCO9FDrkkRlyvk3JMdoqEO8CIZAiJhLJk/FcuuSjMOzor
9u9bDfpMoEV9zkUGkXKSWA8fTsWlE7B907I+6fcnTMGloSBttyVSAIbikZPLwdXd
F1t1hJAQSjg7bgw+WLZUBGFA2HDdiOCOEeliBssMuy+QmFuRHrVFAlMVYsRSX2W6
SLbewrRwTcFO5R9rCi32NipHmLAlt49cM5Erk4WAJABGbWTMkqwCsN4D1kKhWo33
MGMsR+ZlAL7pJb/9sEINm6XYahcZuBvyWW5vTXESGERJFjRA0zTMrRAbWv6EiGCh
i0qNDmc28Fq9XTWsgF9zegceKEl/EJw2wc4bgPdgHkPcO9PCL+QZ3uzU1kxjY/FU
GUeGiF/88L80dsCKeg4oQud4ok/0Hp83WxdmlwMhWvulGqaL/jlZFopXB5IyDgEZ
m08CG5g64z2sfQnIOyOsOK0ChtxC+EB0P1GdAlAqW/WWr5pVU3df1kKxEFy8cVmu
quUaZHL8WNC+ISkEUX87GxiafOuxhVG8djczzItAw1BI1xb28Non8StZClZJaFSG
dWQymEkfGCboipplqXex2xBcaI3jvmhaDNvj3HPiXri3+mud7Ir58aES1aVoc5ka
bj+abrpee0BSV8x5g+QI4hKNLwiMQ7R9Yau/tEP1Im/Uxm26taiyFrAgiKQLUwvH
wFOkgI9F+ioUZGoqEPCmDr8TfErVclUs+qxCuf5ABVseyNp4PYrbqFkHnURUb0tY
YfT24pSzAyL73z78ObMBaHNNd/0PZAJTrItIawgHrkIRMvMscJZfxd73irlC2bUw
pGaicFFr0C/uB/KHGtdSEr/Mb8KY8JzCSgE6h+9IKHF9Eh9EcYNEdyhrCYkDzlOr
YZidvTLS0Yy2luX26fneBShC9GY7twk1xV6XaNLcEDovgXQsfhRchr3eRZ7hJU6o
gIpFXYqofKP0/3Bb0XVsP2fR5KIAZ4g/ODN3uTgg1W4oLblO93FiRWagdgiMHJaL
nOQjoBBIM/rAu0XBfrL5cHXoOTomHajThViuvufZ9voh9ySgbFcfXOTu0D8GbUMw
cwrulVOtg5tGO6Nxo48z01VJt9h54ny9tG6/3sJLymfhrdyYb2HU6libflIGpYhJ
0oxcwaL7i3CAk94ePbsRLnygiX19zy2wH24nHlC0zSOY3HCx7A1K5083zUtOs8+I
fWHD54CY0txPs1COc1Txv/mXR9z5TT05eYHW3jC79i1p/yafIrVjIJV0JubsLoFe
PSfEtkNWuUu0/nUwh4uf/m1Zk+o5TkLjWvTSJ29jwAHdLz1dHsT5ugRydeelEf3Q
EOa+hXuIXdCcmokqoxejuFPPRh081EN9bpH2D0DOwcKTps277MVH/uWkg66XNQva
TRSCZ+mI5RMgRQMnnfIFOapRn7I7OPkkrHsYSwoWlD0vH2dFKLKCzRJYJ0VhWzLA
Llgq7DbA3RVhckEctDj4na0gihSCd2P9pDdLh4EuDHILdKhmsloGwGAXgF+bpn63
G06DK9eyfQA/LwozmmXKHESyM6eqsR8CEocfy1T6PLU79VhQjuQrwVB+QZSBVv0L
DHlGKdzlKVZHCw8jWaS2tBm0MNGAHU9A6GLy1p6sCbkJ7JarUa6R47zIF/Hbd2v5
smwokQijuaBubZE2tEVQhUm1uVGBzVhoib67Qn+u4VN9m8OrAm+IDmUsDaVq/04W
gmeEq1Q/WyoDEXceZ9sXgY+8x7q2+Pk46WS9g95YEBUHGak8c9hg3mGilJ906XyC
QeLWQy97zOEQLQMowZxFhiRSw/8rWhQGktmzWnJLjn+s0+zwhZFXWWMahTew55Gi
HYd9ohNR2HP6p+fTVV3DjKMPbEXukR2MpdB9hIxMuPhbgzLmTd05zEiscGAzT8qP
6gF4PvqtsgqCVtXgJ/WzfWAFQwcGcS4MyoNp33AyGwNrPiTVKSBWNGUruhS7MY/q
1CnWu7kfIjVPffzE0yPTG0dNr+lomsidZJ1qgCTGxftANiI8pf72c0oh9Cu0DBWB
ttkpcH/oDpj3Agh4VxsF+dFOIxdeA30RRgMSMWtoZ8oiaUGIYZNf/Tc7fUDd+AaV
iHlwvIfca3JV6FiH1vSEAseDvdOuo2SHvg5uNVAai1KtptaHWQwCmnH1Gg5lkqN2
jrqK7w0GU4756RT+pbmXlUJHi31Yipnbp6SkdAfCD2vA1wZde9LeNCYYTJs/TMi6
PJum8BynpKoajNNPaF0uScohIHr7FSRMtZ8kIrSwL3ZFjLp3HuK6Wv9uJFWib5KX
RoteBhhnPJarv8xLkB5xw8E2KuUJDvELyNJWcWaF/tP6rPeTx4x+aMBaMSHFNhNM
+RN6lLau6GX53OZ5P3NXasIJqO+SWlTrRG1pK496z3TIbS1RGcViTYlZ7zjZ3aIs
ZQeZY82DOOjb2vs6clei0beEtOXPDJr/CXQwMH6jfGVf9E8ooBCQG7M6hK+he/Sc
jNkusx9wlu4P/gtYPJPk3jCWGCG1c6QGTCnzcaJrQ2HFXidWSonKMYVKH3pxvlfT
dbWmhIwKScGxPvp7IOe0NZNBCDwL1Py2ovolraFOOmXfDsEsF+gbl4R9zuFmlXt3
dgPWvl06fb6cz6WOj21OyDtbwTAfW2pHyQ7aVWF0vIEmSOkmB9OsiE5IhqdKr6w9
hZLQjEY09VzurrGBEMq7Op/ezwbVwO8Dk10RhHovFEkP0jk/laRAHYqCQY8EIwqe
PP5oGRiK1JxBF0QBYxEVxNcRu8xI+jAgl19qnJo1/hyzM6Yab/kRRvfKQJn6c3w7
9DuhvgPNHHy2t9JzUaZxXLbrApCzvf/4iPGgFxkpItfdPixEBZ2nynAiW+TFaPtx
Wn7T72Bj/yEID/+BZHqNnhY7bDc1IxxX8o5jcceY10eXDT1sClt1cjGV2knjP4xe
7S7YgaifwyFXBZ5i2eqw7Lpj9KE6b8fx9tH2inT1Q/SAszPmrVnCUEZ5NUpPy7lP
dmmSphkcSVL8lvlMCfynvItupm0tEkoO3zcB4pvGlVVHfUNpVwvhoktfSIx4adsK
rkqwBL4NG0n2+J1rG1F6kgsRRz2uRWFpHCR79vp05NrBizLlqUxLW05TcFR2NsJN
4eiX14Wq+A5po8eUVBoSJLNgYx66kol3hqJBE1BlZ+JAyVxKQi8k56/2IVhkYSPr
Izy1SbfgBPKdMHWMRYT0pTKjlDvtqiBQqOQO+dr0RgJ8LPHD5AfcuLwGTmMVPjaT
a4wy4TLQ1LQLuQaAgQuoSNoyq51y6cflQC8aN8ReNpUwnCw5W79CXxPF7HXmQqoN
v7M+/IDQ1Xo5tFa3s+QOKo0Mj93OMf0Fk6IfTWRi9MZrhjlJTXTozWkiDhpxEH/P
lj4bqVOxjLgb57YgfQ1ubX+w+PmeyvbgW8i0c2ADcV1nq24wcI9MzZz56clbGuHO
7hOb0AWWWI3Yb5Wcb/8ZcaWr+/GEkyZLKn15SOZOhBghVrZUKbM1q9QobKGgo5kT
2+FU3x2i3lwfh+ndr0YtxZLpooRxBdPEsrT4Fkhb5Ve+i5z7ubn9pWJraAvlO1Em
7dev/5XP0ZnA+qqhO/3d2Uqz/B+y7YDScK8WPB3d+WQODUIIwOtQ48uyIMpAcHsT
ItX9RfjECvd+SDJfJ1jZZpwTMoM1ovjovgBhtKGgahRFTS//rkIhC3keMXR4ApHD
/AHUYCaZ8GNKtoflzrWDlkYdopD6ExcP13CmvvxOb0YOC2YEWSoCbFLg1Exu7+bu
0OLff8THMR9P3Fu9Onhp8Qv9EFkAiwW9yoKdgSWfbCC9V9C4j6HbSln6ERuvs9DZ
P5mnU+osylzqGyezV+S33YjoojW2EuCuXd+i1VbSMuBdUyfpgXNo7oLm2Evv6t8A
RpTZ0kKLdJtKl2FP79yuw2mauKWl19vF6mKu0qfY0cb9Dh/7OLCvwSm1+UdV47oT
z+uZ2Ey+XamCIJItvntTXr+NHXLUzJskE97sVk/J2h7wf5VmNfi92Oui383k3xDS
8G9MmkqaqqAdKmI4XRAxDDpbe59LMQCaioFUOuZFSxk28ZRH0DNuB5OqMI1N4vB0
rLaraJz+Iq0lepsc4DL5/iJmBBU30F6Pl32RBlQoyuFC526WCDBBmKCCL7XGDBkI
cn2nbugYGZiN9TbN/iVXoFiSAt3zypQPPl54Ns91yZUWNAyDpdk/G0bTpH7thK1Q
SF0X9Nz4ilttG1R+5paxUSZe4x2d/1GPWSIK1l8xPvZybMUPd5arQy9QDKVKaixU
dskrF0yGvUl5vi9+LLTO9q6gRIPjyc6+gLAhWFVrdCRJcI+iGeNMsBeKhq4I63H3
6POTO/Wcab+jUFaKQ6FFEQVtYE4gDqUiDYFrNOB+SjDs3c607MtjQGsRKF0uQaoF
ukSTRJINRHPY38C1Kb3eOIy52y19Neh8OGJoB4m0BQjJuXm3/dMnc4egCaVKxFEr
tc3GEvA1CMT/DRB6Ars9mpRd9JHyLUFJYazjjoxINjVShdK+MEp32tG3k0yETLOl
Jvfc220j9pLuYYnWbFVcuaUFOPUeRzpdcTBXgIb4UJ0PptDVf8eL0pHlwixdxfgY
zFYLeIPAVmK1kaIe9mcTdjqcnP1tTeRA+Itp2jLm0zE6OWrP0GYeWwSi7HtjWktn
V4ZXYjNYPOZCjrmCxZVlo4ZbfdfIlImWbbPzB0j13o+wMNSOqiKKnrgN51cbKN84
3jqEnHJFNnmmWrPRz1iNC3m1wdQw2C4Ruboe2RRKCke8uIjz4L/z2bXLo+H6H6yh
jhFSUIGkxgWokDD9NvvOiVuMCXcvy8OkvShgF9TqC6GAB0KvOrfebtjmXMlxiI86
G86E/FsCE6wXhOYic/X15N89iVRqoXPFWPrvXJjlDNdpDl6ycqxbVK//AVvfuUvF
0RohkFbsVq7aan0i4815mlD71tQwTdcTYzr+iAq0+JJ0Y8+7kwxz6xCZX79mh/EX
3Mn6d7AFiLy43xcmjRDd1FTnAyUmOnE1VW/fUDTfTfeKaHtTbEUwTMdsmJcLA8CJ
JdHMdhU2DNmfeJclzQKvGFV/C2nIXfsd6RplwlTaRQWZRnqqMeiawv+QIIZdrCNT
KfcSG/pwzJvrB8ENSg07Rom7UdfZRvl1akN5KGYCDHOr1bASXWMQunEAn6tuiGGy
5Pw46GtS/SCJiP0ggl1XxYmaKsWgvzvkYYOtTWtoBHt+36aw8qGKXjOZ8YYDNILg
7FQaGIcnJ2WKIeMozstj2v/y0s9end/RHUv+E/tlQwrrOIFlYnWFwCLCuN18wjJD
twm6NfYXHrb0Cu5iART1WF32t9lLH4++1g1pQzFcJZn81jFgPgzyeOBedp6BtTH9
7oDSO+l1NpbnaL/iEDR+5V9DJZWvD/K5co9L4Yr30fnNFMEU7yJ8xWAYB+hCnEuG
fyhRFIA2fo8N9UYhVp97430zqiWJf3zG49wzhjgbLbLgLzlCY7vpPRYgfnKOCKLj
McT3MsIyhKbc38ZGVZ2lCLjnB84VDbyFsth65rwblzOuAIn/BFBVUBOiHct2wJnN
+lVi0VTcOVOpr2XUIR9eB9k0+8jbNcpU6wNY2Edxnt9eFNqAjyXn5F8h5Sng4+/s
umMjkqUqz9+iQUbZvlaIis1y3esho7DXRgYXYa3+9ORDwQYJSwcvygYsqjAezESE
2y2/LnI9VV55JpNSLBAYa7Qocu4PAok2i1rJwSA8+FUSK2Mo+GrfJ9+RJqSQ48tH
dT21MBvfM9dY33amBaYgE8u3y4CP7GAxhTIf9fV6D2B/POyj9t4yPMvgmH5jrUnW
K9Rw4iH8V1g63WCYlrZNPh0MipEbzHNPEK/Xdc1wIOIfowq/9uNNgY/q3XhlX8jc
ft8G+yq5Ie+DBzfCykIAuX/QvQL04H5mhCrFEhfNVUEc8IPBOlkR+EOrbucLwduD
SVgCUqzxC6V34mjqlnImB3LG/UP/5EC1GdrEbWA22gdundJxfsHYWQl86tLCeR18
5dPLkDP8WkzelEgUPlTJrExJc7I/xRv2UPD5ejsCFRfUln3qchhg7KhIvWWJgm1+
vLQG/wHAVEiqMvfTMdGX4y5h0MoJwJ4C5Hi4MLIGVUToyxBdaTvTL/NjL6ujOWEK
0BrMLSlU6/m6p/qL8ev4PPVNe+/alSK2sfed8X1R8i0r2LuKDeaT2C6yhn1TwKFn
oSVicmz1Pj1D9dJSbkGjiHNruUQutd/nulzxSIy0HnuV5rWsaZVbe8IDhJYKyyvu
v/BdNuvw1cTJPd6rYvl0yLvZQJwNI3EYDgq1qNRlaRGtBiUHIDLcXEHd5g3rfB8D
59Pe/wrrxUNNr8mdQ849X4xJ4vYWsqSBzhASWm2dKEOkdwo+Tf74aZ9ja4Cn8u3h
Tcc+6/KTZzm7SUPBxpk6+ueuUzVpxPWTCd2eALu+m4l6iF9vCrmp0yv8IYzAr/oD
vw8NyHc7f7r0UdDo1hIAR1VI2t27p+CcDEAcvuYfJi7yOFb0QIAI3B8yyO+zrGb1
2epbO0Xdlcp9udQUpH1tUw3Azs0BswG8qn88bbPzY32gRn2az8vNYhd10kUf76Vq
v/bPOG6lD/qs66p/hjjV8zo0+FK5M1v9fTAtvwDsJ8ru1guo9MjXMnnEy8wvPgDu
KSFwtOhltMpNYcxsPY4twstMbiWYuafzID6IgaCTd9zxK6USfQsDti9D5NB17dWa
pfHrHgpm5lFJXRbzSHNzIp4hHDmsSbsfnZfODCGHyybIY77AvREMyR2SbJUCzDcV
dpoDbUEw8LhlMDwdymllSM7kvUaIWGJGn+rEN2LOscP7lcqGza5fMQe+jcqcw/ei
cexqJFXAKEFS3tioRe9Ai8V/fosvzM+jN6OsUMhBv8FZQilGJQe4XrnMsFSk/9TI
kSz2rIGlenmMqwoOrsj4HsznXMTSzzkQRuhljoh1Smwgbnjx+jV427smxgY17UC+
FMaKIO1pfyMxcJueBtxBONUenTFOUqny7ZgfHLw5pi7POD5oOx4qYH+zLvWUMPdb
QkKFSXRZaGlIJzBAfUJhmJQHsKY4M3EwavC2DOe+NwF4foeXVhcwKCwZPD/Cpm74
3Fv9YpWqx0lHFFmfr1A6x38pKRR/t7qmJUlXRZ4zRum3s8THcyzKRGtEFFssL3Eq
lEJM/YRXCapgOrcfH9JzUHIaoVL9It47O6YLSQ4oSbVpWFEB5Oc6JzBGdYeiljEf
Hb4T5tHnGIuyYZ6d+G/CiqZUxsR4qfuDUzp6t5f0ccOSvcwqZemSqNHGZW1SEX+f
PkADshLhbQ6Op+DxVf/Gz9zBL7P4+C/ViCqFWImefmVuBVr2YCyAPrMBoGZGeaaz
DzFVL4DNy0ZRHwUyZ6B4WfORGeK2aC1sWgl9VRrjvM6iEXqAXjW8PwXOR7KFRubR
3wvDLRSG7u2OUYD3jfoXND7XfYjPl+uWSkpNjbAPKFkZvWauH3Srnsk1TYmN+JSg
6VrtOXDZUIUXw3T0VMS+rO4IasoHWHkd4BEQFwFQNEvv9wFRswQIhJMXVMB0J1DT
RUxLE7CZ9OnLQ1Btp2BuoYLE0tlkOAsdJmXc5MOB096rdLHljoqCZKU7yZajIAt/
5914meRJmLK5tQeNT6RBBrK3jXaOb5yisuwC/r8bkQl1WytNNq34CEiqkpoobUhV
qs7V0W1nqWhYgSVl9wEBkHEz6GNLQqEPs2FUOD6TrNBatSdcjrUe+mTACqK7uqCq
xXkFOuID183UrVIuAqTa42iGePjrglONUNJE7VZGEIGvXETtL6oxU6AjMzWdqSyF
EmDWq7OdSpI+2IzshS76Ghn9t6YAfTCmMK0eAJu3kKZYwA8sN6dCmfFqU8fUHiYp
8WZnF0xLbHW4PBD9bf3HaCUYUDd0nSIgWjeCIwEk6HNJcaMjtAnyn3yA8jRDwn6E
7rXCzpy4Qa/ns9fqfRNTcG1V+ME3iFuVY3y13A2h+/EmvByWhjbT8Mbs+6udTQrm
cSkk0sBZiMGEUnXRUUibu6bDKlNRuZFpNyDCpisJan4nbiZIsNJaFjTO4fRgsIM3
Ni/u8ovQwoYlxzcFB4Y2shKGj4uT+7pnqxoHaY+PqpPS1/73XM2YrU+a44mQEuhF
NSOB5gmZVpSbXgkmXSg57Oc6TIJS1Dk/pwdSi3TBGVB9bxrsaCj+CfG8S4DN4dE7
ianT7/4PqMKrI4t7r0JU84FmBeo2BJlnh5sbMMwpFqZy3rl8vNGKtxy8308zlzxF
fdvclaLhQMoCZw75iDp1OIVYmzRnMNYRnF2aSA6Ba5fKe6Cywywx7VNbxsjPHxww
pQML4NM4UZ3s9dEjcoKo/2Fhc6wLbdBqvoEwsGjIHvmdnd/UtuFY3+Fc5Svr+7G/
qNCLV97q9H9+pEeeaJoGkfQYG5dYBeGZSC/FsRZlVI4cFPP9Enby6bzudWgfA2Rt
e0ZM4KJoFI6gKhzhVvkyVpUAbgO++biUJnh6xBdy3m33j5yxkW0tC/G9gSFvlLqY
Chfepq1bVrefkwN9VKqh1vJgtuGajzGRB257zpr+ZG1a8taZU65qB3Syd3EBvWT7
CCmOMFqBQcdN4l4zlxV94cCuoI1ND45B06ycL4WEugeX71nUAiE+W74Lv/fyVqj4
B6s0uuQQigIldtnumXyMbo7qQ1TnUsrksDTH4C7aCkCSauUyB80hTa8fC+ZqPhAE
5IAaXq/lAkwoNHetkcGBTAqQRIr/pFEektE6KM9ZQLa4Cv8AvYAKA0xbGMTSoIil
Wr1CNQC1T7mm3cN4bcZaEVp51vdQAJ7lYHKOFFXzgER1LY5t3+4uan3W9Zzo/EB7
/vtMjj0+DH7N8Hn1uNlVkOUHo0SEhteRPdzp0w9u4hRsDH3KrT8u2nrriTwYV06t
VYH8RIGhfMClfRb1olp6jO2YQl/6OhHWJxogHRhtrIpVRIB4q7hd/iRQU/UmI2JE
w1zmVZINXMd47E60QAb29Vz0/ZRnpPFTolcswP16Gw3GUw52MGRLdrs6fhbzBpEj
P3xIg58BoirOql+otEsG2Mko/TtuNIRGQTKsDC9w5KQReOtSFy63deWjELtlnQ1B
E/de3CtHEE4tlRlu4zqvCvg8R/oRVQSXvlA33FrkskT2EQxtJcy6zBNvbIeixB2f
4LCTZsa47Fja72QYZ9AosZCVzJEM9FW5vL7Jt0jQ0XIT3FjqGyfjgjoGbKT6KM3c
jhFasl8ooIGtjqCKn49CPb7h3VEetzStK/miUrNVnf0SzSXKb/tVjMJNSSuuRo7B
DZEh7Pwi8nz4LVIyhj8pYeMNKsN25XcCLi7GIa7XpFLoFPQCQW7AEqMbjEHNAxo+
2g7OpiL43Cgq7sp7wP45QiTyO/I1u6k6x+oyxaj7RC+PNiTLruxE2OkoabsLkDiT
R1c28/EEFuhQxuMsCCw6W/G7ABU2Cv51YY+dL6yWFyHJjJtctMxzjjUHWnpxxtSd
eWBqtsSnNI2wQUkpY93RSLFJTEKBvFygNVvmuiSn9/KYDHhfSs6K5xr8/DsbQvo9
udL6+Z3hZvyM1rH//RDiMyRdtZQ8ATlftHVGYNWJam6GGmo5AHufXQ0qkD5WmkRA
oo9Y92KnT1+fS/bTVhdEkOEvVQ4hW1ecEzofizxG+/h3TJ0aIa2Xhp5CJfEIAVsn
s0T3rhC3NZ1ta6gk0S/+VJP7ulhQngqNjKrT1H8TzhEcWCNrueSOxw9GTuKf6WpQ
XUp3heswt2P2CFqYQq8v/xr4PakAWSCznPk7b99EvjQAqISPZJk3TWTDrfAGsPR4
cjncx9DbGjV6EfNZATkGuauoXgziDw6rNYnXbYEU6Dx1UM4mE/e9tfXtBdrTXcyP
8vtoVLNgYBMaPFovpOlLATdNlgYv4Qywop3m+0mnfHXZDQhtN+iaGxl/EVeenVTe
kyfSmm8x6wrnc4y+KkE0X+zyg6RSE6C5eoVUxhH3F5QXFc5AO5IomgfJXuYu2rZc
gEIk3TkZn5ejU29SLEJRZq5LCw9jnd6PTGOZoQOw6EUYvUOXbgPTBgQFGwzssFqA
4L4lRpdPbSD9Qydx3/Wd/1ijkyz45GE9LXPNfbfilCmBzj+MoZbMAHIHzi+sDY+F
CrI5QIek4USRXCq/GYoo/0Xm6ESDP8IkIZve/8b3woTOy5TjZeRCsMa1DIGIoegb
I/gOvtnwb1L6eowHBpiCmBICk0cdNZsV/Yz9gsxmsOGl4glTqX0sOR29R2JsnuTg
0MZ4NQczDTSdCCV08EvtkH9133LMC2XVxsMoA52yL01U7tBA78xoaV0GFHcHn3c3
l86JXUhGD9/agc51iUq6EIBW3fxz1CTJvFjxhIgeQfXoEBeGl6PWQ7NsHrV9qQUj
oIN79/CNrPOv7s0Hk0PNYGcurO14qzzIVzazKmTaI6sUKn04Dhtxqc9N+O24tUoT
/fiRYf7V/mFcHhgq8ncmgHa4SffknzSfMMG/65TJK9zt53hsN6skxuMWTslwpRD/
HAE3DHrfThpzKUBatWuWR5wwFsTiOUhosCJuXmzFD3dftOApzrEQAfuBZWbt6RpW
DlvA77Sbwlxfxx0rAYIAD3BaKjGWA20nEvdCQXvDOwZEc5hVlxwRI9/ZEIHWP3pG
hzk8iQ8rhWsZTUctp7xMeXWbyONNOdaqGF8z53ySOEzI5+ATi05HUpA5nSRCL7xR
4cLEW8nDEV/f+oTNFmftmtF7wVn9nAP9zF7z4dfta2Hw8ITqI2XC9Dk0/YJhSOMQ
3jlMdealJ0NGH3l7F6KDO8PdQRgaWqSOAgZjl3hTy3RozrQoZXLG/ybcn0Cqr/Fh
alcvVp0+Q/Zogb1fU4p82b8PFwn7v3f//3BN1tETmLxf30oNoQEP2bZJ3V4zdf6U
XseI5RpmLPXKMtB/Sv7Bpe5/VNX6QuBdjxKl3R9Qg95nXgto7r3gUiJkxrQ3Cf+b
cFIa5eVGIftXfeeumrLm5G9LymnSrO7ErXoNJF80SeuxHQQ7cNYiMiEMZFHOB1fa
YEB726wmTpk17YHBhSy0s1MqwHK9vvuoOfQWMT0MGdyZPPHN31fCs92v/YiyKeQk
4eEgss/AQJjCjNRh+x/FW/JWyD4jQAz/9ztpyUUYEiq/f9srDdMLfidkddL7aEol
hznThD3IVeCgQLfYC8/Ae76esUYkX1J+35AeYcaL5SPsq56g2CULahVxAfG1QpNE
uP27YvCo8UUhA2CZ+qnN5j30oKdvB7pefN+n/NiTn+osxjd3IizW5v+BpxMTCGwZ
Mg1dcNc1SGQHsqghB/qBUFOwHgFqwDjXXPdotFq65K3FYfnYnKWys9z8Cc4yKIPy
yvHWSLoHdR02+OtQFG7xAfL2RQbfRfiX76OLC/DwWv5RyqFopYCzvFT4Hz2ZhcEt
Wd59q4hyh83labReGYGwEIW+tQlE3Rryu6Ly39JiZ7j8tbyBe/5Hqut8T5BteSnh
CaYCoJcgb5g1IRsQ0ljgo8v7ofCU1ChXA2kmZhuZb1Q8gJwC4xD3EFB9ryCzDYZG
houkq7FBJy+wliayjs6Yw95kHLhu3QCb0U+QQD+oFQlA0JJNckhYpFofCz5+ynz/
Xq67qrRfLLsVzUY7wlW09+q247yrxfnxqEl8D3DIbGk9Wv5BkimQZauj7tOT79xJ
W3KfULOLjvDWzFFTt4rqef+EwFuM99nKnHG64fBn/r/wiOCXOaPbb9SxPm71XS53
h6fE6R6StSMRr/u/D1qLkp+3ojXEmT9P9McxYJIHkda18YaxSv65Xqai0TGFKWks
Gxse+Rck66A3yTfACaKmuCGIhmkGEvQXydUZrlo/sbNl5hqiC7dHYfvfNQRWPoFv
0R4rq7GNufS8NXnGGnN0VGm5MOEjITClKd3gm6DQ8spSYy26jiUMXOH/QYio5wnO
pAOcc+R/txeJr+GBoVF8Y2wLYQXHhaFXqruIvL958gSG82iZwWHN5pimcpWjeFob
ZlZQijRsPy2FhEPuNJKFx3R9X8yCLXQN0aylvKkOO8xWmiJ6SUweZMzjgsU39YjR
esRhIzjEvePPkOPuE9/p9e9xpjWewUkdY0kz3Fgka4Jq4JB4qqqCt+QqsXcFr6rN
aFbsyjUbLX+TGm8wqgcRW2Es8R0+XN8aboPyXIEAFRc5C1w4Vgt4WJKRlU3+qwHF
YJ3EMPpUvhESKI2JTioAbsb+0aM97LvAMmqeUPKfeISLeTu72rnLoNXtwDwhapu1
F3HUAlancjMSJnp9Bv6nedMSmG2j9aKDLOu/XC964sq8mkDd6isRxtA0sJw/OIqE
Nhkd7DTwVyy1UeeBwCds65Tqy8TCbrDPgg46bNJMEw06gOn22s2TcN/nr4RAo1P2
Vs3jLQlWgTNjk837UXJUYWXyesxuLTnIuXkYqkY8IQ5PFKL0FSGU50zpmWh/35on
pifHJ+c1aEJSUHttg1YIr8qKRTvIFVVgWKjfkHwlceeR2ym3ehksVKT7KS20riZS
A0jOx1H6DRFQEsxw9SMuxXtI5KZuv49Us2DyHn6SK6uvNiNyE1uDExUQl5F79khi
tnMA3XiYDgBrrMKQKOPts7fFS7tPGI1K5J9WcKSamEA/mgqau+ecGJzm7N+KZOYC
gWAUp6PBGnx99/kUQbnaJhZ3eh6fCsiG+obUaIS2sC3MLlfrgdzbhUmAk8wsNPs/
tP7NlINYW9si+PS6Ws0AffTyrPrvrOaM8rQ9Esc7RZZnLj+LV+lZjcywstKoGocA
7okf5eF3HFKyiRpVMJEfjh8bhC+Ht9DxYgDREN41lKuiXjKvIOkMidMZAJ+yPSEo
+OZHCN6DD19ZiLCjEhftxw3ra1z025juMZpSix3AXh7ACyM+zx0Hf/ajGyFUjsDL
XBzond2LxVpdooFOeDWc5ABnwaQ+74CnYWwqw5GDIRBm2j53G9itgEP9xU+MijPS
ShyflN7jSxaRWLVS2288FdNf9e6r5dMxLz75/TdV0kAVePjF5zN2x46ows5ZpDLA
9QP5N+ug6RnK/TAYsgGtFBj0B2304oEMb26ZauYg3gVHjcavaqryhXdKB2joetda
GxWkOtGWWOF3+AAhukBNN5agK0XuS6i61YpuGCUka1L1h8olvJ5V/m8dzhZSQhrm
xjbYwDZqBaUu+EXy+dVLDh94efvhkQrNWrt1YCUs+ymBn1q+D7xVrO338IwU7R3y
r2A68VF0YFnZ2MoM7EFBHSkhzCGVHAKs6hS9b7UyjZE1rjbNDPQVaDyd5qeHVn7q
mhcsJ78DKfPcqkBEJoTYxN2/A45P/29/JCbA9N3XhtenuYLiURqm4RAhEEiwdFMO
NqLsZKgscsR4sJcVDULeZAG/1+8C+bS4bbPnYJ0XW3mL0yl+1cHhmcqUjkmrHfKK
8JOlstB1DZW680IIF3MTd7OAF3jyKyjfueIYdwsuBwHoUGpscGl1KMe0RWktMoKj
VZTWQqqA+HlbALxhd/3A/80sWIME0hMu+D0gGUZE8ElOthvMM3j6b0aXYcVd5P9p
4Dm26SZMIXMYx/1cki+cWWSw8/R4j9n2PJOxeJ0TDDzewuOmrkqzytmqF0LmINWk
kz7zuRexPQN1cW9KisXZ8/xe+okhnqLHVI69+itk3D7mQjKsWxXs/j9GkTuye/GE
oqAqDwHgqnHSwbPtI7sdYJN9Gc3kJZBu3PeCwgbplFboE7+3NtHD8HRGCMDQgWmG
6OLO5rSiOCRqGdJs+/F+z3vXbLyg4XMFfublpbjbbX5PwRmQck5q64vi8YDGhZK6
e4AHYrRE3n5lWa4i/u22NwT+Mjh+MLlnepoiIhQBfkCHpyGRz9x7c5Xip7oKXfcQ
Bnefs+zuM+hxRvhPjv263aD5iIL1xCPmN/4pCoGTQ25A+AQZ6Hkc0Pcjv/FmycuE
SHRDjuZgBe7D4VTGPgfOZCdOSBkmrS9qNeRasfBB5BSJJ6DjDkItvabPn8aNj9uh
l0pxsJde0qmKsluCpXgbDy2q+FxabAW9vI52WeQZRHO2qz1U9gYKDStJN6B1+0n+
ZMe7cvb0AKkqUKyHlSj9ebOM9GWFjQ49eMxfKhcA7NOas0m8Nf2AWqMQqxkvKp7s
Blt9iVSBPNYduO/Jp526oRF/4KfJMVlCMHbtSV3VerybBaqw2ROuJFBAGOEO7eqT
261M8f065KnnsOdCEUyzfeI0BUdWw7pqpOgZ8lP/GJ5/qqKOiAOqkNPeiWqz3YLx
a3LH2GZuCP7z+mV8E7lFO9d5hpwdcFk2+PCKqAuQsYDDRPOHvgl2ZzDTzYMl86pl
COUsMUElyfFr7e9oAFcVXyQlKhmtfgATeQkEMF5swnwrAQE0CGLpIRZOZgDJEZZ7
QV7H+hZCAOLjkOFY8nlr5h11EsvAFlPxulqos2RlqqGxuJtag6DBGwkD+BKEg79P
caG2ImKwUuBAH714OXCkqBHuVN8/svDuaB2DWbsWgC+rV+fjNcd0e8Rh8y7Ihh8G
lX0Wemf3w1F4pSneJFYQPIqVZvqje58J7t03Yyqs7UsvTgKefh5aTEE40jUAzQhC
W9PyueJA37MEwRE55Fh+rObJR27M3vPQ69T72av3B+28JK3hKxGRbIp5YLNKg2G7
95o16Vk6FAwebl9ojcpfHvQW3WjgskHMYJPCsCOmv4x3eJeOIVrfs+PQCl8T63D5
sZA7Y/gCnCYgteT3EQlW2MKEca8ZLzlPdsIYUkX/zFmPR501VjRY2JD64ivS8Kc/
rsa8k8pIRtDRkyHTm5L2gauriFmrFkrYVzQWAQgObU/ZMV2CfIWRNThzWmXVCVJy
CWq1ywwvjgRz1/fRM10YQmaLvC44fht+XbpkwBV7revAY4JMJdTF5n4IqqOgHo5R
e+pDcLierm9p2kCjJ4rntVzOkVC+rJnczvSwvzomTo3jmDc3WSJUUoLcovbP70Ww
Sq6C1xq7jLCbmc3zkIbOxAB7wuUBQm0xt18d6BbuzYeWDcI1USU/G8bphlPHO4+5
ox3UmmtnmAI9NVcD/c+e6xHhXAbNQI970pohjqZUfyheJiVm7fA4dCc0ti+G/t+J
hhuz6QKbe5R5HlJOBpwTRfHsgGSEXl8++kOLQaYJdentPhWjGm/Y5bybaHMVo9QU
2bkyyV6Jn+8k7QRoG7L5CG72iunoe430jpf+wHbHyLI6yDeqN4RXtRGPv6f3UzAY
8NQJdOf3yBdG3sP9excGqQVbHf2GU5cgOrb4RrIlvyW95sOh2TO0LJOtv2C0z659
KLfUZNzFpKVOinTdho6hPdLogijvTxo952LLP2QtcoGiJc+nrwLFfg6qu3IvTcQA
zOIZhGxtKowX4slaGeW3YVAgMmIV8mypP6F80ejsbfmmFteBvgxvRJRkfe6iqNO9
yKh2ozcVq042956G+049fbLlvuc/QZjaN/xhypBQCNg4uKekke4wdSkkrvIDPsbI
nBogR3wRtNfFjsIIfNXYikTSTgtFs3yeDWgW8Z2eE5PNvZ68rAM3wHMA3MU/XFpI
sXUV0G8K4hBusqVebl2fdnnzMmvPGEndlls7EeDM3mMVV3U6D4zvUMpTf2uiT3vk
jrD7zXFHCXasNpRWpIwRukWRFhkRa5kOJXbjuxi8ZGK8Gwt7rQL+v/bip0uCP+xO
wTUCZfejtRhC6n8ehab1sWpIVE5fDP+0cwHOV3pE91JA3CkgNoWpCkX1nMbH92/d
Vms5+sQqiDp+u6SMikkSN6zPWTzc0/SZVq1o9lK8m46QyXPaeerx9nik6serlTvB
pSp/XyPH3bzZq1bFBu8hxkFGn5oCPFTB9QRJUvMXcGM6jA7BzQaExwSnlGmYJHwT
TShcOsDP5MANVL+kQymT+Z6Q4Hayf0QMdbAdn8wmTGL4vT9CEhgCp4YY2NhdS9yW
/x8Ku5UpjnsY1qBbKGMgH3xocM92H40jxF7/bH35r7yF9RJntreijWIqIr3wRfFW
i2U94pxEyoZabAL+/FM+HvYU/7s6wQZPU+k0fFzOIHb58z599nDJH1NZjS17nDUp
85cez9FyFt0nNiDkYSkdzjOelxZi+5rHgb3F7GcGGMPIJBUZaukwnaljYt5X+GME
ovOfv4aUHvSoquyIi78m03Rd+jcA5Y5I6/VU1IYvNbDcWbrwB07gDjXO5twSDaKe
wwI5NplaidQNSawKvJYnyq6s0gsBt9Kj4Gwn4GdV7NvhNTOSMSgMRMuLc2xIgKz0
af/QWH6ko8baQbyp+Lf6ljUzXl7uCNd1ITCyXz40xnRg6MTYnX+poroD2ofi+XGT
stS5AKBEMGm9ah7cYOFobgtZ6447WRktr/iJ+5ghoJQICVCRRg7ltPij2onFNfip
GJ/iOL8LWqqEq0QKIC0NA5MYt806Giha6ipbkgweuUfXHRYS9y0BBfpJAoybJzMy
NfJYrZTGLYI0y9vMJCQGBz5q6wx9eka04rstgOPyzDg0MS8N2nGDy2dRMeqFVIHx
WhkYyHXAisHnPSU2OOm2UV1ZPC/pLLiCV9UU+3HLRXBVHmuYJJaPpA+wM2yZgjPf
R28bJxD1QOQY0UFL7DIbc+sMgwohBHiTBhG/+Y1uY8imcgswa76hIM2RN7NHeKBs
yRCMBOZUr1IJo8NOLL+8oMvABuOYvG6RxbJcnHx/XQpXXNBqKNAUR9Pk/6BRRVJj
nIVTMbQ6LZyM4k+tu5J+asleIW1pglj2XdHRZ/0bnmb8riIgB6doABoPfqIE9WWq
OLKiJPz2XkC8Z/mupYSeu/a5DPPLe6Bl2/Z44ksZpmRxTcrXLLntqAAqGvojr8WY
aK4m+mTXkgzAlvvSujxG7Cj2yA8Ct2HmwR6/uQpA/Wa+iacF9J2TFNYAfItAd+1u
FiurTQv1s7BXQJ+H16RMEtwiwFYhBryBi6nMZF/+fa9TEimg9PQ7Z360jRd7/sP3
QzjNw7EEscEAL86uzdxSyo6qaXVVDXpAEmFr3XVlZ+Z+eFfygLrFPyIaSQBFXD52
BC9ps/+GbLyV5mEiRgE/3QcBFz6ztQXpdzdhvaFQ+BM7sbxRNmFKuF4rFi0s8PMd
9NazjiMnOZXzHspJ7JAGzpLpz58FvxR8IntfE03/TLHE91KWhZqNEr7t/VxgJAH+
B3Vyh+IWIf2RI/HvhDtVwPTPg5FaQtG5yDeombsikLQOreaAgTVVQXkZgZ2IWstP
Kx3fHLEP+1kdbaQzgln2dc9vDjC9iyfTmVK45+lkoHshtIEcWHc1PXje0D8hAvku
wEC+6B1VoZ9/CW5YMVcg4D225RMcviHvOAQ910q6tzTPx7oOmaAIh96uvKM0qi51
NB8WxVxJQ2pShasPV44ZUU55FAqiw/ICIoavNktI7CI5//aOCKIAessyfMrD/y4B
acRhCNInp6amXjTmpOiOhdSkyg/uxdnTPyZDD2WXfaZJmspMVuzN3xEw2RUrH1Jh
FtAViEvi3SAqbmLzCwiDWHR14/D5a+L63LOM0GjfNOS1OQ6qf5NjsGsS4ix4sbyz
Fv2VvGmGVSsQ2LSsK0WpGLIBOLV6ChowwZGH/2ByZlWiA0WDnleBBuNIEZACCEj4
VhxTjXCY2kAbWDYI3y7bC8XfjkZqP2MDus/haYYumlWWTs/kyWalp0A6WtxrTM0e
pPDtjUwGHeyQa3pNv5B8tXhL7vMUO7og7YFTbF6HrsFuMd7pe5rJ23jeGYaBprYm
gln4rR3EsEYjcOvWGeFFPG1JpMMHkItP8GmVouLoOtCyimjOfBO6HB0EAWRqqjLa
/F0yVuH6RNdzxweyw+0AymQz1LmIQsSxtybOVrSDopLDHyA9kdMhQ6pvfbo3JMoD
vPA4HD6DhCrzm80lTXuStZUsvPsVi5IoHgQO0GZvLdcYFsl+29yET5Xm3GCspZBP
qgifFCD9vl+I7VW6DarIuhnx5UgdfO1gFMc4nlNYYY1cdfwJK6+e2XjtbFsjQpKi
MtSECCbuImDO3SKwihAhSM00Ea1X18mAcQKNCcdlcdf6C4THeT39LumI69m2u2j1
fHXnCfenq+zIDgXzPQ8RcqG/GuHFIb9aL8xAMhLq5Uo/qZ/YzsVR1CGpMVLLnd4/
OCeb4DH7VcwFi8pjIKYVeqtiogn9k7JRn5tmsGwEksS75MBbr+Gyr1IyDzCcBQ4L
rkJz48ORw0ujTrx8GnWf36nEM1jGQIixxiYh0OiiDBuWWuHNcgLKwcWPYC3Nom8V
EJWat9BcYus7DhoGqRVEN9tVKWjPQFBSWV0d4xMZCWdw65YpOnywN0nhV6kmrcE5
7iMpSVngMgODpEe2OZlcfi17QgKeWoLFrjsEcZI03ssAiIZfUPcBBfUiQa4T2Wph
rr3TWCxpdf5RSMHeIuN171nAWWx0hM36JVj/5vFgq1UyyFn7hKuAsIU1u1aUugAu
EuiRmsnxEi8KIP4NcADq72gf1FX8vjNaP3yN9Wozf0z5/bJphbw2IL3D7d/R3dmz
VtMTS0gGHwWLCuWb3huPzaHvROvZGn0pOwqJIY+vj9jmVo2ctZoi37eUjngyNVig
bz3X+F2wwOKnqMeK5d+zknIHXy6+7E3T9FzJ6LYfHScTxJ9hDgkTDazIqgHoR8jZ
gvwEYeDw9sJWrMZqOcLRnH98o6LvviLcZnphEFrNVJVehn00JpGncVGt1y0TFJyA
jQAcqQtHcETv2DrvYTup6YMX/rG8xqva1lwUdnYKnPvfU1HNIMIkXo1w0uuHhjcp
LfXIVijez84HWqYCGN7lQqZciMBy3maPhWzBEA37gFVOY0RuLepK4rsbKJtxmvxo
fidEGi0LOYEHo/62TPTcq8WjK1/6gQ67WjGmYnxwOS694b1za1pqu0Rp7Y28gFu+
xalNmLZKdFbF+QSSIG9iDEp6fnddPJHc0AMiP+Z+rNnvDFVBRjsKEZnTcSpVCwkC
7ulNLvI9TOXuiR1cwmc6Qgk2ziiM4l3BEf8C2LTPfRo5HF8BOlmw34hPdMLW0+/o
6Xh8DhPTSX6MwznkjeirhLAVMNvLIwfU7FAxPJaEZ5JP9KaaK0GtE66UVB3FSmKZ
OYpp+yM7NZSS8TUQDDUqILYvuHkw9Qq9jURh/xevqMVoQMBpG8Qhyq5QTAlfYUpm
pO7uCHkftiKzFKlXxUP9NW0Z/HZ2o9bTBZaCDWsMl0bd8AGtAm35WfuSpJVlIPeo
Q4bGeFhzQu1ijZwbfRkvA8IpkvkthsVz6f6qvOg+8xs9AtqA6pNmePtAqRwBZXYm
oC9rjphi8SvcE0Yu5xPeC8ciRBS2rTqTT1mv74wkNdwujbsvSlCXq4Mz0w85VhUS
D2d75guhDiIrFSiMcKdEUo2wMtYCllI9Qgm8GT5zXLWiHCBQS7RcxbEJxazI8UhO
Zjnme1itd78k7cJvzbtUpTni+BzcS8FofohkYmgsm7sOglBImo/nTTrs3RBcWwnG
tjZF8TvDbdgXNH2CeO06yj+IswsJfQIZDDeaqNVuIQOT+phVnVo1nFPd7taCqM/M
+jcafnbSsUQZYrOEWjZRv/hdYgYpUz9fKhrFjKmV4Yut73grLSSymjwe96JXhHMZ
9daKOuinm6YurNpqirWnM6QRevzhr1T53FgVSA0vAdcmMq21fwF1J+ofD7qry1ki
QaF3pjttRqEeQZdMAe1frO7syxDp5+3ObUUt7NUUNWD15OmY8STlrsE/UdFAw4N7
WQn5qkJDopILEkB/mAguPZZlKRezFPn6V/Wc63nF1VDZY2mzPbQcTfGmVZZWJ/Wx
s2NKwzU17rOSdWNrlPOZlyLylZdaYB/pcsFiPT/Jt5r/2GrgmQ0Tden17i3eMG/3
DjmQEbkldwyBQJODnX17qnMyjkkkcXY5DdmyvpqkT9QSrhvgRUlkduCGmaPnw/ub
/NwCBwWT0XMiv55fhWC+XlhRBCIbU79Q1qzEhNr3HU8SQG4ajacnVJvQVksBalY4
aiIazvhoUqQJJsNZxe+krWP0RevNK2yOZFJSiO8JtbeHrSl8SfeeW/+8yqWlU8qm
mgqTZv12dvuuHbCWrwgIX3i0nLL6cbNaxCmW/WsCi352S80FADYeAoxvhwrUOLNd
LKKqs28+7ht9WNaWBHWkC4vLgQpnUYEKydhT9JpnWBb1YMTV+q7eZxfmt1zuciDR
QNmd8Kpgx8l33I9Soh7HK4CmlrvkGx2A3YhrZdCXahIIFuzxUsWo3VjebrI1PIFK
7L4cvrstTO3A+qyuceoNC2aRrGYsPMC4T7qD7doXZDUN1gxA6GCdk04IlYcgBPS7
bNlPfTXpTfJcPsvZIo16XRCJ7+1gyQwC+oUnla6Wcxt6B0oa9MNceXySxQaE6y6/
/w3l+nCS41rnJd29Y6HnvgDwgZfpmhBUcrNp4qYLerREoB6QdM2HN7XDI1frRx3i
fvaW7WO67JZr6SuWPdiUoz/Ai96DArXxefzHmppNyu1ellV9R6LyKtkVxYx9m53K
o+/na7B8S+/6/pTFpto4UVMjDIyEE01hjoOsqPDOeaW8IJmuLl85oTqbyJnd0khK
bRvpBYB8c9w8On5FndeLUAKuK/YxFXi7ZsMQ/5dVLwFMI/z3jyH0jUUTHrf/5AyW
hrV2CF9MBrXAILv62dqVXKT/wQ4fMT5rUYDV0Azr9RVFJ18VVJfk1xDdwyUKp9I6
A5hqtoYZPH8iFR179LdZiYQOA/Dglpp18RWTGEVw9cKWaMpAYWK9m8i92L71HXlC
lQ7xOmgsAFBtE8q7Yk/g74yK6QB4um5MbusAIzGfCzoQ6tSrz5iwxlMVBY9ycYZk
L8MbAD0kBUxU2lLNLQLgPUJ2HnQ1RrRft5pOqoErQM43V8QTD+Bkafhn/cAC8thQ
hViCMd22Xxp1GJNR+OoPil1HM4Kc/RYzlJFI7w9xjWSrczBgLUUObd+CHHPCRiiH
6QpW0BgNBAvRvlicE2KI9yrm4ulXoCGgB+v820XcWOjIpSWVDGhUJ5M83gS0aWkH
xegwpCt4TRmYr4hrDb2Q5K9wxIodwmHVk2rUIabackyfdoOLO7F11mh0HILt2ovD
F5+6mbUzzh5lNQ0vpba/gFjYPuysZM0xfiqpFq+FUt/GOGaMcaYm6305uoMKryFA
HHlVQo7jacW6nwKMO7GMhn/5o5BkwEaNl+E1AglF3oNvBhoXwDP20E+7yD6m3RmR
w3aumhm2CxV3PYzApc2j41tnzKWm0cvHNKIRdzpOMFJLIlZPDVbyKU0e8Y1Vhfme
Czc2Lz+IYDrERdqh9Z9EnJVOwlYSKZ53+i8XwzXIEKALB4zdMUvQrHp+H7aBcZit
+FOtAK3SqWzwEmOEchurR6n3WAHBrMgnAljuSssRb4bqZ68w7rS+ZF/VPxSYOP7e
XGWVRIjXGXybUOJVY66qyFZ7FLzyKhtBCdIVVuoQ9vIQNnlWNA/eh3HNxSjpMt/J
oaePAO7R+HsXXgsKBuXxxx0bCzxkS2z/sIgzeCLt+M313ZGxvxv5steb31F5JoQH
aMdD3vmHhtNDNSzl5bLKLCCXe2ur84hdSoUxyRAIH1kfK9+4iUgO+eg3+ItTixoD
bVVxNWoj+DHLbi+lcJqioE9sTm5ATK9CzigF6jH76WpMlJPztsZnS0LKSUmK0l8O
aLibFTWbQEX3+7PUlCAGoXjz38ROfkpeRdOWsBVWEvRA87V8tG/6R5+SiyRYZzhp
xh7aY1ve2iExNZBPwJ7ET4PhEvCSlatDwdDLfc9Wh6elLToqq4Vh/WP9CaOxM9pd
EOvrrtUqG1e5HaSc6nTVYSO15bHYeiK3DVyz3NMeW6SkqjTYBxeiTu6LMB9iavD/
REvUjSGusqPTCVM4mkrJ/qKpo1S2gxEVumsugxCDqjU7ZIaboSGZ2UGS2YINYsy8
bMRKVJAsagePwCMIUDXlwqNcVs452lc44FNgKnjc/niCxDjRokdihoGFKzK5ydUJ
9awcuI3vChasAxqLsPLhUCd6cxDLP9XDMtzKHpFk3FQISosJE0BLTlFghf1dkFDn
/sB72ZHN+LlS9cWxQytg7xbuol/0zdMp4KNm19u99aMz3FJDr3UJMkxWgtyTCRgi
aMVw9A6e2NLB0HHU9RDaRptWsJbT0XWqJnH5/V35HfqfikxBidHxLKH+aDP7J7sZ
Yn15l8t9eYcN2uhK7y9sSfPYNYvp5ozuqSX+lPoZ8/QPNdRyH0QnzVtNA01crLNS
X7Pyf2Rl1seuhWF/PY5snura3a1F/ua36zZU6PUmhDW5ZqSsL4aw02Uqn+NUFpFW
5e9CtGOyqYF+yfxliUns8ytzvSciNU2X3JGV38OHm/DY4EigWAbgGC1dupquCtS+
11pJMow3EZe/svyXPxgL/4iTgxuq03/+69UHQt1I3ItR6SNo39iv/dfDZPg2jqUF
iHMzYyQe6ZkDmFItMJFepKjClfoovSNpNTtA/iUFr6EQcvlhjVy4pUT2zAKuJ9ZW
1EIrP645QY1TN+fG0VDxVjeDhQ69Kxbr/GLI70VFuumFnzTf7sW3wGsQeQft5xSI
/DnQy9v2CxFvUNA+pN7JQH1/mLxwkvMMzjeCWhNJ3LjYecpAuPakswHNs++34fEb
JaD3BzwGqhPVN4FUXVRVwtOQ0GGzE68wqe3d9R1qW4FHushOOn880HVnN6VUB8Fe
Xf12NmGAJ/dPZFExA804xaKULiaemB8xJ244ruTdL00Kv7c/aI9PVfkcAChXQTZi
SGa2CgbcTYNq0Mo7zRa0ZMfj0nGz2PfTCtWVd1cPReFbDsk4RxKJopo9JKVefy3g
sBhwDY2eF4PTEYwGwsRsGLgiO+M6XZ75iIdjcHAJtSToqI4I+ww/g2YUvdHsqM2e
MO3Y0foRypWazjKB5Lw/FPAdkZv9lQTSmJGLWXfeaERyBzBfI/YjuJdAdt0TNMCx
yLR+ZmnIolxAee3LLbUMZwHtl8HtTJNQoKgFSoWsJQhQjHHI+TDQWPHktlDrxdwm
yOf01hpuS8sDPjpk83/6RkCBrhqyHYUwbQe4XiLBL6fd9TLkZfw4SwpoMbe0BkFm
PZM5rKMk3QdHQPjG1FvxnoddYtug5ln/sWNVIN0EHb9EljEbv0hWpCnBohewjBO/
baT1BNh+LJsywkljoLmx781SS8e80TXCObRze8Gzw7tAIyOafcj3FBr5aqa6F0NU
EIsanAuVUriPau3EC7VmJ5BNrr2xVuwqn0a+TGzVq90noe+bvOv7uBOqwwokSvfX
qSTX6IWhAD3MNgjjyN5SiH+5ncd7xwetaV7PFSCJtOteCxByvXsRqPuiGTAl2fJK
Geb29ghGIkRQzsoKQyD3j5u6JmafajYfZwmz/8INxBoHv2g7npQdXxgYzCNnAdJY
qEGclBMiJJ9zqO7PPyw68P4NdOtmapqLhtFiHswza0Zw6Wh+kTu8Sc8ZEm7WYggS
2ro7/rEPbzdF1X/NFo4HvLMT9N3YOY5F2zHuOBwBaUiy3fpZbSQ1jLDC9GsvvMa9
ZdDefe8Pb0WZdNSr+4bj53Pwp4rv8es+ILaikfxjEmr+4tFIQh8kX3e/gSYe1Lp3
DaOYZneXiXaGQFjW3Ml29upaY9L2/OasZCX/fBC0rpWOiJ9600C01t2G+Xadxace
Tm3XjLyYSwmum2QBBNDNDMyp3VgCZRS4hmuQXznTJZA4wKcV6rqquaDdFw5jrj0S
YJ20ZpgqxzeOJC4mc0TtA43Kl9dajkIxbrDW0oZhvplboB8bxIC0mmpcTuUuRWlu
amAhM6GFW5pq9hYK/j2D5kHe8qgFbzj+b4ZSzwMb0bj50EqA1NMvB1FuGLvybkBo
nwJ9dGfEy0gR72hmqn0vIIkOflPbUPwBYHjx9moEeiVT7wktEMYpTvh8nZf7/6MK
tP866zPNoRRDA7UypYs4QtU1rsDKnDK/BYGik6DrO3OkLL+J0vHALT6jHcbDo6B7
I0N2VpfLN+wve+SM52CxXhPyy+OIazRy/bQfLQvfD56H97UxxV3U4BJbcQQamBlt
UxhG6TuambqmDFhw57+p3+GjbM8MO3dWvMeZaLvUM6zS3Tfb5f4xjHYuO+Va+4qC
othyGGz0YRdzr/pLasoyoq19tGG4kBEnCIanmqH+ExRHvpALw2FBePVvaLSNzaY3
PGhvmQSHRl5rT2yItVA6SHdYZBmQTmrPGnzj47E/+VLIWIPJZPOCcSRaxmp3GBEo
fhwBxUO6uWgLRBPxxmY3tv8/1M9tGNL0XZg8o0CViHS6wo5RCSlufxnU5z2FSfZR
DNVanaI1LX7BFDvtesz4Svcw07BlYz117svMxkNlCRBkfcQYmuKmoP/WaoE/VEDx
xGW0laurRAdvsQBl62jW8wlwohK7he60H9f5zEd9FtWZhs9Ofpu0hcJcUiA85RCB
Nd2Ta56YvaG8dyDM6DaXr16cJczJ6ukR3sizW3D/rcyEYiGpUklzdRhF/RKzTSa6
vNt5u1sTlwzvPUqjockDyivNPMjrbiWU3reKAwQ1qo/fB6kMw2oHUMmLiGU9YwN/
c9JwYoq0T2LnxvegHDytps3imkRC0KeszQ4KnUi1K3xXc3bumfmlFltKMZ4FE+qt
qIpGNlQZgg2t7yPLFHOtY6LHKCCcgkvSIPXrq5/9xXmc7CH5qosj4RhhR0t3g//3
+HgnPSzMcN4qk0egZ376daaqTTwE2NUnrqknp5oanD45lPiPGU1NSzDxkIooD4KD
ii6XJS5jCltsNMN8Hd+f/0Mq5RXM9z7/ADBd2AVhqDtCz7fTOqjyVctkcydNOm7w
1vXKke24tgg0NoYKmnPXM8KVE7BGenqQqjnuorWSehJCGfj1x5PRM2vBtQ7dsfj4
gVJRM81HRwvHykCkCgAy/sIvtrSBuzoBdTJBSNzMoqyf8IVfTxdMMqz0rSeGDlFO
SBhV1/olnT0yubMK4wvGiF989S3AvhAfmFhDMTbLofiyCMmcmuKzwVvvURaP8VnR
yFiw1rNI7NlolSLrAhfcufW/Ax9xNZwYYysA9ub4wwLhPb0RycjrALIo1LpBO8Xe
QOpZ6gNFDOnfQv4kk3jaHesFi9PdpCuib3IASUS0alwXLjN6+X867gt/YNI7pMRC
xHYL7kkUdNFeW38aJXd2XN715fa8GuLZ8wMKglLunJ1FXHaUHKwE47VXTG/Q0oxE
35XHOszFig8W5LLioZV+NUPj/UqufjK/UgXvXjPHkBg/ZrHujbyhQ5gQ0Fkx1Iky
8uoTAd0XQDjOf71abbAvXBoqIIoYPlt1bwa8deywRfcpmo4Pg9XuxgMD9XgPJMT4
tw/amac1VgDO4ye34pQ5zw9fnhpF8hMaB6INOmDUoIJe4bFXm2EJpAQW83H2j5YT
0njWzaLvqD8T7U3nP/KyXvwo7pK7KLCg5plaIPxFEtLxLYESnN30Mui1fULHqFGT
6bPwxAFR/e7bg7WWz4dA5LJYWPv9FtVQjlUluYd5EoLWXgFPvK8g65+nddK+M2Ja
CTJ6UDxEWJHRZJ3sKcoYrSOTgjcupGR0EFv3ws8htS6mqMTb/hGkCuR9OpftKEgd
heanoyNxW/VRfvjyJ1O13R3n15SpCa9UW/qcNhillo+F9bfYKJBdmGgWM795tQ08
YlAwp21TRL+EDA8d7BgdcZizkQqA6vWgwlMd4EJJPocrK7y+LK3DH97XoDn9lcYF
9o/XKtfSY2GbAKuFzDAAckzcLU4scbnNAR8tCr+B2gHiRcFOZlW57qkJY4TTMr6E
UP1RPMyYgdwro2+0Lj+BpIhd5N+js+Roe0pvTFLb+L1D8M1/t2l3PYJTV9oWVo14
tcCzO7DEd5s3CzCRUPThHZZaOuZZJxBdx8zqdGaS6RvFGa9rSMgibIbXw5Utbkap
MqVff7rsAJ1RkVjMMI1fpCP9HLE4q4oqE20Dd6UKQL47kEEU7tyv7uVFgbt39Z44
YOcYtKsvPq+LDBHMaaK3l3KjBCLel3hN/tlci0tbWM8w02o3F46Ixp/hgj0zA1dn
cFaqZrpGpzxTLLbsGboOazHdl3DQx10WGt0bdS6xH30c7MUuinb9zRwjb7t22hJm
IIOl2cJfYuCA2GuCo1PiXBuS6v9HFJ2RY4By8YM8IpFHpIid5de91X557854m5Ku
4JsBLTvQ2KkXs6t27mZNlIw4v5TYZA7dPZfAsPqEoZnPfxC+hf6meaj+luCBxTvo
FUCg6Vg5VKPshXruJozE4waeSkVlGoakVv7qDaw81l2GUYtKgYHlE/knEUC4sL5n
3WG3kSC3oKrFB2q61Xbz5yi6SFwtbIIDqt+9l6O9YJg5ZHII/hKxwkGSj1BR+8H/
vGMI9OrqS9b0ETR3aUPJ87kv5MCakUkJMSgNyC/ZGgUJqjK8P/bNR0TxEK2MLaCY
wRZJ9c8XiZzHYuU6wuFKjmKXSMHw+WAqZNSaP0YdqthJO59LeYiw6YmyFaY0GATN
NgMtaGvHx+bvf1rajFs2vc3QFUljzBHeK+rz+VqQi1H2MxMtj3e7CxPF87B8JXGM
FMmkFf9DiwPeSSTct4AFpE0O9PY67w9Z9Q3pN/Uxtk3xuG8Jr/ud6H4yFmPAeBXT
WGCzOLjNhudVtsYGjNNaqwjQ1esgZrOkPL3eX2HeS8v1nXyEg/xJpdWjdXYDQvua
AtzCRp9kzzFxjgZWx8LYOy3pMub75PGhgqcMLa104y4Df9M8ZQMAolYpaN+H+jxe
Tbymwk4XifKB7wSOSXvyKFZbYOrbE+qE8xZFp7gASJuo0+4ERDV+cNo4lY8Bz4uY
rxiL2iJAZUQa/Hw/H8XA/11C5Ds9ppNeTgphX6smYn9Oci+Qix3iQgPU5uqG+FUl
L94YPou+2mno+BB/8CETZAvQWaL2t+siAIhvPxeziY6PzkL/ClxgiMkwCKW+HWQa
yFMp5efHXeBLtwv4tsAJFiGDU0z7PRuGNdE4vAHDZ6v34ZghDjsPKvSiiyQXpZxr
7tTqXFjPjKPUSMdWXBSit28r1yPyIksYN1w0Bkb5l3DRG4Gfek+w5xgyybVFkdJJ
wWcnvG9mBXblVAsRBHptlwAJvSoLGBzle5engFwb/oIO6Ptkyv0gAc6uoIzS0rGJ
W7GHsRKeEumpJqq3S4XaY/w/qKzRAmQq/UByKTAhprkq20dJ3D3ntEKMnMgYuYhm
sKhm5oVsF6akDuBwrk4bYj6xYaXEfPlTDz8BpjmJDmH0kuVrtjiDM8AUrqcn1Lz6
S1l1hzU8M+0nhWxtAPFnNI60mcamkcaWCtPJBHJvsreby2ilC06+gkevgviKd5KJ
4puCVJ5wSqmkUYR0LD8GJm2sPM9BIva/LhBfAy2V6scSdxJv5JYj0LHsxMINAv1O
dW+Z9PqtYyFzxrunaFN0qTiYp5chFuKyYgT91kxx9IbeTaBrWSmGSC09S+eKVYtD
tp9FR94V/86DNXxJgy/0HwU1LJiwPiD2KXkNkffe9064Dq3hNi+yhlr5HAsPr3sK
CEnywq6WBCX0SRXGvXxUhYiqsQda4CHxVcLMUYY8r1/d9AFPg+1fsWJFRmdoV878
pF1BPsh4CbcshSpJ3Koixpld0MQclk7iPyC1mw6vAzMUAJwffXDauI+Y4dBb0rRn
K3c2ceJzMi+n1JlbEiMn9N2Sz/2bjnCSa6ZajEa0/qp5PBbPLBx7s4Gc6/1Ef9ET
V7Gpb/Rnd3vCYEffNdVKoLlX2G4uEslszPAFdJN4SIWsWMBL6tdYi0mBgLUkd4Nt
lNoVJaOwkWM200yVxuui1mi5kAz/czpV4IY6s0tbgSuaxMruZl0EsruUrn7jPeRa
68m14+oUbqgmErdEOTMHBgZF2xA5h8o0P6n4xNPAX+ZJJCo416n9gFRgSjGdD9He
uLhCwnaRBo/1L34iGWy19uKEGLhpiT7J3C1Ky6bTE9Qt0e2bUvw7XKc7h1N/nXAd
Ito4h87+9ZW51w0C+aGGDFDr2wT/ScLPzRp1+6waLtHcR3nIF5p/9G7Mq32P+0pL
2/wGJpiqOXaYQSh1rlP3orsbA8NegG9yAd8CPLDs5wCk+VBYwi6cFGPrH5vsXOYW
7ITqhnosPK/vEiixIPGPh8aIgyDwY3nBbsMPfCkRGuctPWAIQOycsfD4OjI4bPdu
EjzXDjtxurJ75ujzJga5UcbGIOjeNHdA3VoP8+0XZQsqVk2Fq+5r4jLYc6vHyz43
IL5hGh6YlBqGHu9dBpVRC8PzUHPegm4VZDvowI/daKwujztO3XzYOoouEHAD41mo
a3GONDkpfkmFyV9TbtCDJIyq9qrAMbZr3pJ7+HG6unlfv3IPwxN9LPSCz5lzwC9h
MeMM+nTFF3GD/65LYq24pa3z+tDafMTK7J1pJIxqsoZCcwlCFLh9+hHONXVdlhYT
YNOBeA1MiLMXWlani7MlueI7p/zBTAC8ZRqRv1k9dDaWglUmGzjSPiQBtMyuwb/j
sbuoVthP/dx7+q20kpsHoXOG8mPgNRTKDWC4LHSkCSK7TlSNCu3nsbSkKguGmOHG
Qp//p/Gm5Ncb4rpjiqLPhSMJG6iXH7Zc7qecF6stCBRyy3AdRvkzU4MNuOInb9OD
6TNZnJxWwkcARrO7o5uqZyQqw7cCUrZxRwScbnjzvBl1941ObsfAnkG6unqjrANA
CjGOed2Ls7sC9Mfv8irr8xY64qke8dM+uKC6yigBVRH3TrjsyqCZe13LxJIJmH06
w/Eao4G+ehnKF20FysUlKV0xgEuRaw+bPhKz3LWt3UxeAux0apdyhHy9oTH7154J
OWj+x18TgU1c1tv/5lDXn1fwh7ECHY7uxikg8MoipYBWmOGsA/V95Kq7OSU7c92h
fiJl5RtvffENBi8qbssWIDon3n7AhSSQ8BoLrdvbvJ6Q+AE9/xD08MlMhE40Chgf
cyeO8i8sJsDokN8h6jt1lw2KZcAAN3+al6gzdZF8A5yxyYGavSJFR71yjAu3WENh
BuM9I0M1kqa+0K1bxEVppv5iUPb8AFQDv5StdAI31DJMvuTwh7oVAUoQ1bYWE884
XX0UMfKV07XWXDjVvkM7Xu9HljZqhIWyvoXQb17m2kvRfNIB8ztuD++X7h1cISe/
+j8LJb3hWhr6scHPXqbK7hhE+PvNKsv6hFLPzoQFcdZcVZaZq5jDhD2Jz266Z9XI
T/D2rssU0Uj0r319ZGJdalBMx+n5LrYvFr2w0qEqJ1IjNdA1RrKMCilD1GEF3yuD
u9v2PvyLsaKT0D8KrhA3dLRMk579a3xLYqFEbSevbRJt5Yb6JCcTuFmWknFds0YX
xUHxNWSjOZXNaFBuYRcNT0CzF/AGl2tKRfInSq36bJbauQpxXqmgTE6iafYHUFxH
PxD6vpPJXwARgEz7gaJlA5fp3vVgDIKoNisipdnS8I958jNQhNQ8/suxBgshwyNF
Vyjie2sn12gyNkeNXgHrT8gwqasBXA7c74VxYxeHCDpcFTXZRUiPsucZvs+rOcqF
dGB4V+WWkpkRW/5VdnrcRJ32knfVgpg0aQNzVIKenXgZl9GwLW+e724uIkUsodvJ
OkJiaeuSp9f5acqRljnvyeqELwmzh+VQLX8FBgUHor4nYbvIq2Xf/rsyaafEa4Ml
O4Xx2exE6WRHxP73L/oCiFc6XiPehYXeI08haZujiwmcvWf/GnZIeipqxJSRudsB
dzy/B8NKkaCasRiwNeyG4qYy1rk6LWcpcX8UBueBkwIQ+rP8IZPigaIKlybze3gZ
UMY16tdqN5jpsp2xqVt+45H3Db8VvDFmCupCw8z4aRlSngp0VSL7BN/XNgnF018e
0OEPaFHMC2ibeGdI7PWf4Xn4QCW9vqSaT86UZaYp5REfDNXobfof/R2z723+eK2Z
3OvHGrS09dcLJ+7iAETXgPEZkvBL0Sk8a5yFa/9hLLrTQceQSjcJbLVHRSZIXnyb
J/JyPz01jw+hUOmSj8qZ7eT+1fwJrKmQLhsdTV38Ja9l/FFPu7tIdMMPce7BQPA6
Ix4Moat38IAp+5qtwA/UPi+VrrZeSJVXTBfvxC2Kw2RFXIj/qHmP6gP+sWbLm33M
jWlK7tqS2Kcza8kwtcNFgtC2oLJ3YT3cagi4wZo3dJ91FsBCzFYdz1ci0zCH4Mmj
ukNhsJqOYhDO0f+iuGOfNMFMRcNDU250SfOx6mWiedXRbrRkSS39sYX6klswVBSD
szubufiCj0aLpNKX1YYLVzaWHIkE8JHP6qZk88VTZTB3q/Uv0TsUuY0CV9UJME7I
zEn/RH3zfOmlZwK81lQPScNql4koabHwduct5+OHD7QltaktIt6e8hUNQkHix3DU
Zas+YeXN1KtpuyHyovLVuqWX177R+kf2Af1KJW4+tS+/Zf28BeIwOULjmi3uYFmm
6UjqtIF8Z4TaiYfxCMkUsnom8iykTSkmqIAxi0FBB1GjbNeBcb3gY8EsDYLe6GHe
XcT2TuEf0C2Mrd3r6qB5OR2l6BNNA+bkcfd4iFLK0B+VLLGD1xIHXiAZgR4hm312
t1V7zmR+mY6F/ZAKDnm2Jcp17mqjcyM73y16gmggjc/hch2S7Y8Jj3x7XlxvBMGW
wCWZ51gY9swvc4ySr4WSDbEHw9c8OJKt6P+aWlM4N4pJxDUNGfc/du1cc8Grmm2H
lOPe6GbOCcGjl4+KQgqORqkoSIf2ercsTJaPEga55tfN8uFizN/H9w7c22PGpZzj
Aoq1KFwIIWbHkyGboQ6Ha6GRcM9l/D864W0kt+kazIrnFcnKeCrhn4xkHBICz9QP
Porya29Qhc5OCvbRlOD/0t48T8MnVEM4BKaEODufP/PN+hZzbjYFfuRrfEaxu2Pe
dF78Ct+JH77aPWA7MSLVwsj/OoVz0WGbgedxWQhHli/zzBC5Uh58ae+OhzZFnpj4
uSLSX0qcxkpdnXtHTs4ivoszstVQ0xYpJQfY4cNUbJPvxRQaYCGeG81/rngnJ7Pw
UdduylzzVNBk6M78KRlMmsb3NW0o8szPF+Vp2MLQd+DT/4JmrxHUvx5Ly9TQIvo/
t6vK1BJqeOLfd/riOYAef+hIsQoVW18dw88r7OLqVQfohPj7EQGMPh3NuZQScMBg
HUPzu1T4O8/xCOJGZteQYEnto1Zick5E1cAx9vAU8GmnwzPjk3v8+F1aDfGOThzq
wjx1zVdylaZbs6elpby2dzkiYA9KdfRqR0Vo1O23spQPxEvINqYlJ4uNVxc8bFC7
foiTuGL3uPn4RnGR2V3daw9YcKo3ixLNoWTizLRadGic9Q2/zUi+0RRiPTCepu7f
zYuqRvM36R+ldXVNCkh+jSFgmtPBbsvBvmNZS2Tt73tNznpbyuro0suG1KmhjVyb
vEIvX6R5wEBFPQlv1jXfpqBzM+0wON4iKiCVl6FiHk0vLg2F+euNksP4UXTQRUVT
N2ojtNc+oG01dbt28h35wM9Brq/StsEJDjXuKmuoxQxajZFrOT2kXjWF+UPQas6a
agyhd8/6jLGthOq5SOwnSL0mtiYqxiC0bpiWMACw2GE7ShBRjdb9Obu1kmTVEuU+
wfcna5eKWLyoASvrPqpOvilOg7r8jqcsVYXLMolRw8QuPiDCyrndiIUIeu5rPc1a
kNeybXEe2H6Vo9NWWzHegWbIXjCXCot5w0tvfpNqx8R3AhpkoWy0lZlafYO4+dHH
lc5l+gbmNoEAi6Lxk2erGQlFsnQm3GRpjl7diMfJhsSDYzHV3Nouw/jwXoPpaOsn
Xw1CoVLBtIPKbmyZ8gGkUn77OaOAVgqPJMMkDiNyb5PICwz1muUCFPM1I6qLXib9
1xeedES99vsftnjD8zWcyldYS1DaUsMGgvguAfXirEDo0Y4YgK1ae8b85J+7Wnvk
49MdmHT7+1M4+sFpOKMxydN9bM5ShcnJRNimcmEL1gw5ALCMFUvmMxhqpOSLPpkY
FfVyh4RGjZg3/D6D2feRSaI0r1OY82sYN/eRHG8oubic9X7Rv7uQSdBrIK7uv6nB
rcn49LBI4GJqjhXy7+J41EoV0I8OpI4rBhcfGMDR+ot1DfUxjdtevFU1Y3itr1ps
Xs0EEGIbctYFqpJoRAk7FG5NOmzvGsPf1iP/SdTPto0YYw0PTq6c5l1+272QpRPj
SLAOv3H/T++ojWpUwEcDzLiZ7jHRM+H9g8SCrG6QyH44uYF++lQdTqbbVimkN6yO
PLrICR+gCbUMdtOp3w5GbehDru/AXQAVE+lI8RaamPsWap9D7ftwpj6bkxfqjJdx
FG+NxRKRD53okhAuqbaH/dH5GYRWm8+YcXyQyQuLVpm5VWUxTzkIGqYBXI9xL/Qw
wltR2w+N0ULPidhxxS19MO+sM8IrdOsiK37kqHiph6qKmBUeMLG3NFycNXvXBDer
LUoP92oyjZv0pr9s0foyF8YDXwcPyBmU72nGu9V6stMS4+wqdbDgre+ajII6d8wF
ml0KKcrEkfY1kLw2pN017uiVVbV3GBewAZjpftSF+Hy/WhIZshCdZJpXxfolKUHr
s4/wdeTjOO2Jw2wujQQa62SqALv9EtpL8sHINLfG93xEL038zldxeczo/J89XNyJ
ltmFrd9+uI9z/2XA3G+3iX1troFDtKs89XAvRC8behFQhaclnFl+/UKkNCvBDYNn
GpTOm3DgelYQ73Uhd5zOdkZ1F1GVGJKuQp0G8eNqGHZD/eEXRFWh4Umve0qyaGlJ
H0RkAIK1xFsK8mqot79kMLDI1xmrY2rpClbyQuc0hlVkPF8QKxUWKWu/t+M8G6TU
Mydnzg3QY0iaA1rmT73LmgL0BK8cxIqusKdbByA/95fWNjQHaIYv5Ak9FSVll1D+
pyXx4v8TO7BxFHlDOp1htQSludTHCrGFY4b+M0fSfp81Xg1G0sn8vLPbmPRMXBmZ
PMvQhplP5DpGiwVL72KbFITC56F3H+FCrkmAFi/zlmDUPYJURdQINnssYgaI0N3x
o215initKudNzb16hMOSfIGTD8H6grQUVo5RaPJDhGrWEntt7Bi0DJpGfR9sg5xr
LD+Q/8e4oOmAMU0myWgyZ5Bn0IGco3OpwgPyRp9eQUhqVmCRLuUwAJ3aHfND65Hp
Hx5ZtS1tbYNvMpgk/fuy7nDODqfGu+ad5lTFXYyVoCb3/wIvsQ425ZXxfFA0equk
x9MIiuEcRwPA1WXrvfL5H6mSuHFDbzNHmXCf3Eus74+YVi56jmOJaW0c0txu9A0p
giHpnEBP5tZSunQntdQ2QrhBVCUM8+DZZe5msS4Mwhu1OMt3L9ur7JfAOj3HdYly
E7Wae9LzSdXmT0jmZuc21Tgx96knSbxQ6CV2MXDQHCPqvoHmYHraeFpI5cdw5mxL
poUo8au6+vB0XyLqkYi3P5Css45BXWY4igm5pKNAbQsXnmnik3g98LlwIBp70Wrh
sPgGzeYzIhZw84hVIHesS1naCxjCEZhy3E9bEUJdl4aAdl390rYPvRXgUuJ0I2ZB
4nxA721Lm18YdR+AUfg5AijlYFyjnzji73OvfhGM0KcjDMNc9Vo+Ga4LHN1aeegu
xk06JZWNlOtKQNiGRNAkD2DkmEZtKO4+wZfFu7d9JpYA3JNBOOV+wwyi0isgV2hm
nNfSn1NofPfE6tHDWIHV99fVcmiOexNIeu6CewQjxnckaC3854gT44KP7SZfAhcW
DD4xVZwGvquAzt0od/q6YDF1JOUYXnYCot2YnoixUKeHANC+u62nG+NkdjsAa5HY
cFLf21tRu5HAARIRnqzyqNDnXMZqGDUtEmzXjsa87XDGn5DFxBkXlMHBMO2yajs2
Cz+xZUHMTac8ycM5S+qH22TrVnDYHvAeoi1seRaPCCAJ+aPz/REpE6ODt0OJVeUC
wKkbkIHLeGP5Dsi1sI3ElyGlpkFwue+fMXsOHACsjI4QCcSB9vOcVOEWrb7HqykW
bAoo4tflUpG+SudQ7g6OBWAqMOSS8+FK+aUd+mxXmoTYd6wv8ms0tFLzL6CEsj+W
ftJGItYFitKT5Q4EViEbN9ZcrauxssRAGmKGOk3aaDc5fDUyrKi00wAmyTsYNWZk
db6wUXHh4WJorDoWwtiRcTP1R1UJMpZdittWHNOlAt2x6YKPjYw+M04hNJ+M4sk9
cI01X5p/24U5Tasw4tMMNtWahUdgytgTA7baNqn9QOguxS6qNSjjBPyY248/yGRr
V+1KEMtcI2ATtg9Xgn4my0QeJSRk8mtoAs8020rhzhXPayZS+QtYDnJhGwSA14US
Tl67aOb6aWcPjrR37TlLQrOSvnGJ3AG2UP6AixB3ptyxByBhb50YmDyAe3O1q5ST
0kKHAd1Xu03kj4m0PABssb4FDxPpSdyWYDR0+neEGpvIMA4D4tmxKKV62rKBjnoa
47X6HyPvxKxYrPbu8NhzvbEpqxSxXetbYIfZ5VlTk3m7g71HLA7G72fA2BgrzP2c
iDJXTEnr+J6M5Jcs7vMipsDEp0azZqnkm9b5kW1LDq4VJEymTvogHU/qU8QnGBiZ
8i1C72Cj96ufCzMvTWyT1dZVT8/YvZf97cjr1JwcU3M2bCXFMlgBXxOVaP1KBj/L
wJhVbnynlmrGFaiuf8lMuT19A7TSZE2X6G3cKUdNwRbPXVbAM7P5w/m9uK+QRgAe
DYXhAUbVF3e3MIt4tx6oWDUnIznvcVcsslCqcdBKec8PyqxOUSrzfWYzC7PI5cjW
DuPQJgvN5B8szwV8dMKlOoEiR4nDwQmmDn3ckD1jBPvhM2JsOzWOK3B2MtLDbORd
JYjAeyMGmwusaM1cO8LyRILgUhOI2mQPPIhbzEyedx7D2p9JlNkjocyC2DKoxGhM
nq+ofiBshUuLr/zdknJ1hD5SxWZGytNwhk9qECVoXJEu4OBj0cF+woK3jcaNdRpP
xUN0gZ8M0EevzbFFsdEX3aDbVne42keUGDdJh9AONVhAonkWZf1ze9vgaq6kRYce
R/57LUZVQC1Dwd3U+Gw2gggar1JYqpzSvWp6KaU7Glbo7Q1gAAx1pBHOgazW2cgc
rmX5QR6WIdAkvJyK2+SgtYmMZ1adD4X/trQmFDeJqLs2CPJWX7kBnihTzbM/fevo
4e5L52l+gtlSqOI9h1jUSCc1UYYOsypkJ65vDOo7u5lpMNCzjlLVuoKsMyCT9d9e
ai+LlbLZAyenC9vhMbBELhhByvGrSIVVJmO4kE8FCe7meh3jlWYgoZeO6AvIwUlK
0M0Wjc6Q5AMNPT2S2pEkDDGDBQFFrxnNj82zaBXPeboPUqHXsYjigVhcMyWWr3Bm
Oaz7SKZtK2lRFlaUgIK8QPn5KCUJ/aUITvu/N3bQnen5+Q9YGFY3FudaO7U+uv4Q
NW+wY9ZyaJmt36DFtR62hkbt1hZhnKlNaEGN8cCwEnSy9NLR4oblZGe5jVITKbYk
XfnwZ0QBQJpzrj8ryp6z3vraWRbCQCF1LGXM5dyMhNP1BqzIimfWdaN3RMQCPDWn
btajVBQtkKJhyAlauLG83W5ftSTatlFRG5U3BYAz69pAsJV6NuRLAIpYuFAkRiaF
pSO7tNYiswX6hgsm4jh6MNtJ0tev8D87HCwqo+bdG0zk2J1SAJHBGAitju30zPwK
DdHIJmM72Rb0bvtp9M6wNWdhrfOpyXop3tt13s2EH359PQ+ET8l45qubugEUHrdD
iGQLOGsW1MVkkomFN5JUMPTRwelyHzphpFTOkVTUoOwGEbPO3Yb2WaSp/s/GjgCR
OR6vhHGTOP0zcTK3HcDOVTs8IqhJEyAOLaDqKLHx5ifd3W+zczeYsYJmvNVnS9iD
C8w7vtgLkRRsJ9TAE3P0LwobYkMz1gv/O0pRunj7nF9r3eJ495UaaTsASqAqTT77
DMggOLMc5F2r96+nvCKNSTVmaRVdPxT1tPwm4b5q9cZMH/6K2FtCs8EReItVKAS+
6A7hstOum+/OKwn7bOLgXgd2FsKHuOcFEycONfz41OLb2pkap4wpV/hGgJ4QEZbh
PeS8X+8qTaQzkVsuy4JOtnbbtbxpOiNtPusQYuZ4NbTTnvpmTX1oSv6QvWC6yZyF
00y1odrzOtN2ZCWOpqCq5OOXV+FtPfEftdh7ogyaJphtzThMPfUZLsnTqAnoPPOw
fMBfuYBuwwbRct8iF6wKAEQnEJ/97elvfdieiaedttR07yZugYA7nU5F0f/ppBdZ
D6gKmLwqnHRv0/t0rhrG/rFHjHQmPZyB5m1D1Jskenj61g9M9g7JVLocW2sxaBJ3
vvH6MKbCC+KiPdDMeohUpQZNJg2UzMK1qXbV1eLv4Q5RTpMVwNqFeo/QMEtIpj8+
hkMsg41qas2tIgRHSpW2m6CyhNMeU9LYiQ7uns9buJlIf2F4nJxZbObi7LPXN4aT
8a3DsMTCjdMPzKdfj/df3DtXpWTSCLtE0FqwprtLN6UvRmTQEG5ieKdPKCV9RAUe
zxWo2MLSLyzfAEQDUKfDu5RKjmANjcpzAgQxwfnbwiWZ4GY5an3iK1tProB9K24T
2X16eO24WzJkHfdwm9g8ePHR5e2nith33+duPermEiZRbzVbGjPeUmg/u0ic/vS2
jvoOu/4YOS8HlblcnOOHItpS49ZwWTa3K1Okxhl8KDyQptcX0/VzQkBnePB8fhGV
CmvJh1H26FJaBWCyWPJnPULKWzAX1NWrK8c1MbBHc/l5f1cPQycOwGekMj/9xST8
x8gtt5/R2+yphfY9OmVx8/gH/esPGeJH81/4W0lCeBlo9j/ayAki2hglcXPDV46o
1TDMtBjl7Uf6Nn02WKJ/R+/mjby0Q6Kt3X2ByHF+krv9k87S7ng7RZWduVFp4WhN
/V5UXK9MkgqFzWIq+CK15aeNV1cpAlZpi78TUSuICBnMZjy1rf9nl7XGIj8OPf6t
JCe1SwiLflsf6936lq3XD65KJ41sQyd3UpS99SrXNw+TEdxbj8dLVYaEx/h92iDv
sVI3BVGb9Bvy2rgljUlLthOtQJ1fWV7iRc5wGcoYvmco1kt9tgP1HEFXMXAKhSk1
Ak9ZYiblp2JMLor0a2hAsoWlOY0vNfy9Y9CbECoQu4YNtVsSnM71s+COTWkls5Tp
4Hb9KVC23PooJPjRMI2rQSfiOi5BAFtUAy89sbY5sGMVMPci5fxIU+vUNfyB/0B6
vy2GTUiFXu+0ITlSJvD5WZ9Ua7/Vp6gUl+6UooqUIqE6VT7TOFmqyCKQ6vrZcUNK
x+XZN25cvqbF9sVwPz10IKa4UwB1aNfz1/lgHJX6Zs2RsOhyiVpQkb3Z3mr054dZ
SSU/3IBXko6Xw8pbRQVROoNVzHwm40GjW9uPfaRxLuGHvqZMeFYwfzKgTzxjU2nC
u09JWCDLj+sROoO9Xbr2bmHaOr7X/MrlWrW3+6OL607HDD73OYp73MZoNpM8xtPq
+jEnImRf0ygbapudyttzjQ5SxjJo1Uj1x4lx6VCDUNVVvEHrAwNhKGG7qN2BJgX7
pscawphFptidfWingfMAhcyIInLunsV+8UsWVjvW7MPk5YQnPjQJHR/4eyG+JxUR
GEgJQpmxqPr8lfN5zDC8Rc5SH+jVtliXELOXlEb9MvgqTv8XN7JAFfGSShogARO5
MV+I6SqWfgc+aowEskob6Vo6xJ9kPI91TwL+yw4hLPUNDnMitQEywRrNyu6jJ5iz
b/5W0dJHZPBrixGDeDVTQP5C7ug1FbRLD8N1c6+he3R2B9yh4pnLP3PrTqHkcb5r
1Ya+d4ctkH0aATh4K3bGXm5cLzIQfGLce11+wSqBbr0AEBBCThMXpMdP9J1Q5bOl
1j6iEI2CfUNAETQrT8rWSDKGWlPM8bd6s1qlMOhjPdT5hvYFePJP1uLNw0nCALOx
+3GI4UI7FK6FsrxKBFrX2pf/6Nk7tokynA3jgd9YjudS5i29jz53rwVqqR1/MFYG
UKgXO+6aZVTXkJ5S/OMs7hmR9Xa3AMNRTpBg5kICIy7/SDlX2+koDVeL4FIZFITX
HCsFkppqG+6Z5bonDfNzHKkGXIWIztJfK962+htdX8nuOySj4ajl9FVJdMfYj61H
ePQGWhSBK4hUegL4A03TMyl4lp2INv07HLcTx3dTd+Rl0GapoHkosE7obaVJnUKP
C9oL9SlpZVS4f/6BxuKrWe/gKIWFTdCCM6O4XmPgXBHy3PRMpzD4WwXD4RvTFAmp
5NL5iXKf0owf8lNRhiVAMjAj9+dT+HKisRchVT5giMLph+0GKjXHVodSJUurUVO5
Fbo03r9Ygjan8O2hfm3HhihlbE/vkNJ/nV4UGBhRns3UWO65TKIKaWW2jcXISsMM
c8SpcCHiURXpehjWl3XBzYPqoIs63JfoQMchlxUarYdFBmq8YwqbSrmU+C5VMBrp
82TjIos69K6+ztE558UC7IfRFD7Xs+zaxI3uhqiqEK0WRe6x3DCG7GjRdnkDFPHX
rYdMT6aRDRwbbAJYVAA4kaHoO8N7UDIRVmHUHGf1gPDcFp6thY1HLI8fsXawzwcG
4EpzE173dojz6oRc1NriODJDNn/+KgHhzB80uMyHJZKEgG7r+0bdLLe7cWxAN/nG
2m7rhB4OshP0tHlo+7rxNRMdKxh3lruOmH6L7I9hFbAHtmshgRLWHL8eSs/ZeNC4
1feMKCYMKBjCzHADExYloUw+y6DmBzeoImVuBH7CaLoV/SZ1iJvKMAjBSAl1krmU
kVDxOC1GUudizJOnPgAnoNTlNKg5mCvwsWWoBmKQ7JUKDB0NwMLCZcYjvC8H6BwQ
MxsSZ3Fgtms7BxWqAwj2KRqqywpPZQ0VbGvZe4Urbs2EXnAyo7/teVuJnuMRuUy2
QO45EKjj6bYv6oqPsQiWEaDIOoRlmd4bono4qY4ZgTFhT0wiHfHJHGaD4DbXlagZ
3fGpZP5e97lEE+e+OEvVamZr4h5k270xDpXOC8Dh1FIR4RfFyQ2SrkfKuE72XBqq
brSIfQWgb9NCuij8WAiaAjbVHMRDZqJauvpl7CBbGB0kmNyRjS08KRULmWhsthVv
nWdk3DT/805lYK9DHlnYbeoDG18pXmOhnKRwK81TgGk+KPRXI1QX8oEI0WvbmLpN
lOwvSCqJCAj9mlbIm/wTDiEth6ra6r+A1tQUo8/LGZQ87azK8CnT0iGLF/s8CY6L
2BaYkCvN8EaLpEJQ8hAQQBAFq9YV29fXEV8LARrJZvlC5KPQvdKkEBIaCwUnXdId
llxu3uzY4hF8uFYrbjtw02pTb+9xurfF702bruwLtuQeWOwvyTHclJ2+0RukKiUc
Z08eY4K25TzyiprQdmaxo/WIkIvNf/izHkJfSnlacGC0hd54NeAe0l44/VvhKb4L
xDlLZbdWnxZnMGi3ecHYOmF8uhjTYvnAQf4oxLcuRp3bzFA9SkesOjXjKdrSWSEs
kUO++J/yMcenoSzh2eLbaQbpBDosSG9qcO8RF+CW13/tjc/zsThH26F7Iqi9B3/c
knkA3koj6J7UyLxZNIZp2yr8HQwe5baG0pOmWL2RfT7umvP91QbbYsx2O7vs3KHZ
39qiPDe6ytTzGY6vMC70rHs5UMvIRnf7K5kL6Q5izK5Iv0+fS3Mzaxp0CdZoy0W3
R60S9MEpUjSPFAMQKwjabXxIfCBugUIkzTo5jTdhp7fGFX6YFeeE60jRX8qkZ7ut
uqCiuLiidAHeZApdNqoX0g9vsYSRfeA1lQTFxfcfSnLIcA18nibycV9He3i6Q7CX
K1d2fiva8/p5hy9ySm45kdvkG7lNlx5cibPgWCeSgJ6uljNOEemGmonLX+LE/S9n
+IWHTUl/xa5skEA5/D0ngPR3VUpPSt7Zb8zHiGyUZ9DEickNAwXkEmcm9icF7FK7
M88xuSYuNA3RE4KRGfVKy9CGYi3+xiVMuELBPwcc4c9BSgRFI8vMBuFJa1JqwY6l
Qr2GxwHlfqWJu4f7U2AyExBsutLGdVkAtL7ilzdQRrnckADo1jhwhErYO61ugndd
2KOYB3z44sjaVj2gZ3bKvGO6SV2r0Vaa82bUhBTH7L8geAeNe3pOAxCeEk0ZPeo7
APCMlcemNn3g86IMXEROBN5tLDDC+3we6H2vPPFMQM2NEM0Pb5FS6hR3YmhYUWcR
7fP4alPo/E/e8NDXTmROkEMrfviXspUzppt1fSQ5FYLGMZcj3hN+YcsINdGnpVpq
3uxHOZqz/+UqSvJhG0Estrf7FPZtP4zT5ZfdyOi26Je0e24gDwKYVvCDE/nR4Nou
WRQJHW9JJ3oTaIV30F0gZLx/BG458MRSKZbGa4y54XC477ga/zVkx20izJRe4eEF
za7VB8+rW5xwKNq4gZfO+ivv1PcotNjbVrcfpkJeSLtiJs4Cx3EBE0C8Mzy4pDSK
yYepbXoeSzWNcNH1e3QAUjkAN9VbevmmAdVs3GsYmPnowXDVN3CQ5gq8/dHOITKO
BXCmGCzsk9safLt3k9aK+R9l13xGK+d9N11ty1vCr6nH+00cD7/zRpPXmKH17A3z
Omf7fDOQc0eBndJTycJUtk3twXpivlRKoiJPqvuyeuhlE5DGhU9Tmrn60V97h9iT
hY8zuhzRHq5RE6M2Cdo0m1E2RSsY9Q2X1b21NVs3KT67ZUqUqFqwb9w4sPM5FWQY
hnpPnSYLbAL7VsvjGb2ZmNmrJPvC5ZdIKUGZIys+4H6LkdwVeA0/ZXeEF1ggeRGX
e3fAy8eqlRsahQnfCfrbNY9aPHUnRTGogfsfcOk6rA+lCGkmhE0NF+689J+keWh4
nxLioB5AzUGe3lTZYr8aRw83yDXnlH7/NX1/pdqbWQ7uIm2nZsojAhny+w/kD/lD
hsl+0x8JVmg8YObFAf2vswWgDfMky7efA6Rk31H/nQbTukBKTB6bTrgSxD6uaAl6
iOTox1RIH13NFwwalophfTeX6t/Ua3vLpSoY15QAmqV0ifJ1D60X2p3V3rntrN5l
llrh7cDn66fmpp/nS3Wvrxg1Raj4xepixb7dF4UcsbCxPZR4J3uhKumaBKXzgy+l
aSLQBdhjOoc3w5CGCmguNl/f45JeapINmxEwGlxRKYurwD1AWNEP27Qccffws6fo
3WVpM3VwkE/UTz2PbzxxaoIDYJ4duJeOwdbzyCBSab45LQ4Adlzc3m7KCIBOp9Xi
BdA5/z1TFn24IDZtqESIY0ETBdiutLs48nHgO0Zmji8oXJxrH8sHOdq0ImR8avb9
muX/YHCk1iCMsNU1SmIjlalUe4dIxAt3UvGobQhYSVNJD+BJfe1wGgwfCa5TmZgK
MZY81VUH+hn/qNgqUR6j/awU+6gqoZCDxhvYOpVwzIj8eL9UWyhhweHRHA5xrMDm
JRTXM7pFV9BxTlQv3XrKRwq2zAPnd4AwRSVnhtKDUZKvcNZcQJqciCw+1gEN/Utw
pJZSmFrk2PT/nsPwjoMSUkpJUVrEijVHKaGgjrFpwG55GFJS5vOjQ4x8kKzlXQkY
csTRMc0uvK0myz0wAwohHPLBrBB2HhBAbuEyGQttTp08vxGxdeaXCLGIlPXxNfsk
kYdWQqCkOefGzniNiK+5gPu9NJXFEE9xlI9RbPZwua4stw9KZqcgidSgnAnWLpju
GxjbDIPNevgB9aBMyuqZ4S6JyeTRvtc+QPNWBPhRzUO6akB3X5a+v+4RnBHNIaxU
Bc0spAptoCpF7HENmdQL6+vo6Cx/XV8FAvu4Fulj3TrvFtWc34QvvxPbpVi8m9/0
bO+MtVgOREyNT6zJkAmJFu8EODDCouYi/vAoVrUrdESVoHQm+L2PI3LNm41ds1Kk
Zu9OjL1ih4N+tO16MkwX1IFB/QxNjYn7ZyLE/+sf735WXhS9sDKDEQv+lxGAPVB1
VNyC0XJkUdF6FbjTE5tHvkO/OeRp0/nzw+MRT+Tur05ysEVlSAX5zKTiHEV2ZIBH
2pScRigMXN63/ohlRSz5FbWwi3tuyb9W3G1Xa+8yljuYIGwZnfHxz5lgTbL5wDba
qUQ8/QSjFBnM1LxgZUZJ9HrMcsnlnacx0PNQxL+Z0z0igfsCQt6wG/12G3d2evmn
A+rfEaipzbdZSzXdrRBmMKsUdbvJQ1BQaNbpU61eBtJssC8W9XBN09WMQZbiED0K
DUGhF9qvWz+tAaOeWLFyBulTDS0a/Noxy9VJr1GI7/EeCguqksKiJbsudU3zcLnZ
WxpaEWCfta2xT9fJSFTJfS6X+B0rsFELL1al18HKKbRlmNtA1xKOQzmpzVoxJz8E
PbZN5ovsySNBUfLNbB+WSAbrYQuq9x/7PHdVOIXAag5QQhx0TRFmhgPVGxYh9yVW
qf5OXTfFh7/7V7Uuy0Y4+dWqlsBBBTp12fvmSTgwbgiryCXIFwwZrii+pp2E3wIe
mYYTVXImwrPc+/JCMAXhDJCY8A+RGL4gJx1EddKfwg3uZQ71Lnslpa2XYj/oYaHi
t/nLkMDsHxNbCh1jsvjlJth+31v+SwFxM5IOTGl8QWlpadbCrTAuyPqwEdjlJQUM
R0k6pHcEjHum57XabLJLUpuMCALU5JEbp6oaqYwGU+knVEvDb8UHac/gND2sO24u
K0rPbHY/kp7f7wR/K3V32+8aXucqcJgsLLxNfbJFdXWhHU1hnagL2zMnjacD4BSK
HUyYf9Vf2SiWH4YaQeQVi+WferZWtdziDd0NwXDx1zto+zeP5JwRCY/bYAcB6ye2
VcDAZses1+vUXqSspeRF4p7HhQx7bh/pojsFozFkJIrbM+9xXxMdMzqNYqwRWZ8x
zHI7zxRBM5jZqulzUkVUcLTKbXNE3pX2y6wUuH61YTmUMV7UZNERi5MtZ/6XFXxt
gSXZjPoU2aqhW4KVj8yXfBs8o0eroQyxB4e1fDAz4mHVltk8fLVZQI00rBKJi7Qj
9xErU7G3VbzFOdWXbR+6VM4hySx7AliyrQMiXLtyV32aD6tXRSTbGBXmQPhzTWmr
YQWBpK3Jim8xL70MQKBgDPYx6ff9ffoZzd0TcmXw6qljZLT8KMj+mXdbAy0Q8Tn8
/9GoGs6AvL7IKiaicHiwG71a55hjFpaAUO8rD6jHly5OATabtqlwRr1zc3D1uJp1
BEKefvjUCAmL0DBKAMnJ+6LPgVatP0NVhslYIPOqoTXzs2gFiznahc5p1xTdsNP/
3UOayIwsu8dsRSo+X1vl8uNdMnBXrX96uJlA4acrz336W6tKYyWgXToB3mwb4cPF
i8ZzuyjVXRqZzmv9c0Lb+cvVif4xpOJD6Y4mP+MIQD0gkiPgZNwsK9GqvfIVc7Ms
yc2dtcE2HEMEv5HtHq3Ud0AlgUd0lUarwHta9DkurOL1V5McdkfVvXP82qvgyxR1
vo4vFSNWpXZf8K0NM3e1kxOvpRVS104tZ5EMgrWNMSkDR3CgC/RvuyeBlM+tGCrL
0fI0hy3v3R5gtkLdrKi1cM4xmG86l9/svea/Nans5riPW3Gg40iRqyZ7I/hqn1rk
kDGZuPM55Wf6SLskubijZ63Fuw3xQt4J7vOEjbUYOW8qcs3jdjyl1xSxF6rGbaM2
Jo0E8Ubo3vsxoim2re7HPmQoYM77FJFQijbYesBYanE3NkZf7uIF0yDoneUIbRMn
RM+yDgwAWPvtCmfhWxbtV1QtxoFncKPdEl58+ElHLdeV3/7wQ4LuNfIZIP1yqdYL
Nl2TGdYXnUnZHeDvlDyBp5TE9AjyPXjP+AKgYG1o0Z022wUd5l47SGFDNVtXEdnS
oYHpKF9V2CR6s5jVBnrqyKzq+MYyzMIQj+0qomh2sIpdlrJpU5hPm85PNw8hzhwT
DTQKjFaRzshm6MMUO5OzsexT/n6JJgtDAG4edqc5Om88hjsKBho0BWedNsCXMd2i
+8TjQBpK5Wos5rgjaaCIIuNdyDq1R17cpGaqNMdhCTVz3joLNsXCAKznTIEqiKJE
BuomIpmv5dw9mYcx7BX+9jnWWfjKq/Rp+0Z23+W0YiFq/27eu8QiUVUbN9od4rnS
f3HEBHsjz5M5qSIZ750zesm1h1XCtxqwS6K5KoUwFRxnwSJju9LbJFchbcHvuc3L
k26LPXAJJ5S3vvmH/BfFrOoDCKxaLO6fKYXzgJ3OPfOZUyuVNPQybRzw9Zvb0ERt
BQ9sPwGca0SxawbXiTcW4VTC7b4vB9q2GnSF70LjugcBt+bBnBabLYXHC126Cx2g
aiX5Lqkmr4VgiYdJV9Eo3TwYGsxaZAu+4IzHSGy/5ccN8OsZO4zWYjorQUuRY7e5
YtBfcNoy7JAAPrbRXcDHwOo0/ua1ZS7i1M9JS2AJVjOKNHk5zc9JWfVumiRU62Uj
5NELKyNvBLc8pfiqGDxdIOJMlw8HZaN3YhuV88WSQKWu3nYOChlq7yEAvzwPSSWG
NThYNTX2xGeoyUR7qYZKdKVClhtpWLAxiZi2CQBKX0FB0NYQiTy2btvNhuhiZI9L
qtxfxnNRCCofJTL5AKrX0EBEvEBmoZuDogFNElg2ih4VX3/MfknYgcWSmLDi86kC
nYRUGhjW6uuQCGAkU0Qyztg9FhQVrDPZLmr+FQOoxYy2Co6dcjZ2Sb50BS42acDT
9DOOYbkaO3n1fPn4OzLIS70gpwvCNuXXLPyAa+rHkvnDDOT8c2z9uwx7qfaKWDsv
dVGEeYLbyCoH5OTQVSvCvd23YLimhQ6ZG3lnHN87WhMcd6Z7wuNgpoJD+/d9Dgmo
qQLkX+MGfLiR5koOiogviwbHj/BojoYhcidjg7/FRDp3MA6RYQRNaSqi9+4k1p/g
VadqsO/U8wsiJAwlSDDuv6668i4FJgVyqNzSRqiApAJS9Rd6TagE+Tjcw/JGjo42
DrC4CVNvEQtnAqU1T06zpmGYsg24Fki16Nc+tqTZ1sfT1X4HuZPerZ4jPKalF7DV
AW5qJupizkfCKCqW27ekxCUEnvUHCKTvAY9vrSIWNl59QzEXcI6zO8RoAO7jWnzs
ayMRqTFFG/Y++dTgnh3sPyGfwO8K88ZDf5OQ6/aspxB+RBdd1KSs0lJtrP7/NTa9
IqXH4dJYn6qmkBL9UBOmJPBgYzp8r+FWmhlu6rJJERcLjtYKQa+KBfnOqBz/XZL0
ik4qOP9KupC+Z2vK13l0FPfH1/sOfBQlTXsVluqHU0W9WcDK4M9o2RUIN0lvz5Qo
dBEpnmLxB2GauAvyT/JV3iMkhBjAwBn7PwAAX9VhrQ+trOkaI9jG6YfWb7lerF+y
LNCwYPaa0sjz8PzvA8mlK1rpgZGLVaTCCgXd3pqv9HLZWZ3//Jgb6Tu37slrQKGV
KaXnyLjiPcN16qp1EXa/08H+kTUAksjlbKKBggUVyZpqJhowrGNCNDohwLex+q91
UR/VhhJGiV80/66dZi+9dlnzQ1aMxgCgMgkVdSRENESRhqUyt1I/ho/eaJeHp7xX
lyTK+2H3+sRjPzpWGaWVmEp/rK8H2+Z2s+kqvK2zFTlC0sNGFWCo4W85di3MOP0p
iWE+/ulgjYHrytVjaGGZrCLx1Mx3tiPiZqvhHx78OBoRVp69C1NpjmYQd/pVS8QL
yvD3ZF5whkRUUkI8ljm+JhnjPSqgxY/mOmUm96ZdT+l1v7s1PkoyhqxnCYlWO3bx
uf8OnXcZ3rRKF53E+HOVRVaBWCaSV6XL0kx1c+DQUuEOjB3+UC4H0una96+6+LPK
a30ujo5WEE5lK9D24kXD0xfrGE4JSAKWdC5tbVeqKdAn7tSjvwL1Rvy2Z8N5paD6
fwmXhR4cTw6FXa46OEDU1exjDj3R7eQDZbAnuyZ/4QUl5TurC5kn8GEF/78f8TMJ
86VUWBurqhcU57uJD47EJHG9M7Or1KjW1f/NaaMpmiFNKliIHvTsxd9VYYDZYEFK
a6HsASGpeq0W/ooPa9XyK8cVVfk+Roih+WbfMFY2ZbeMVVWlRMmJdwh2GVV51ZpC
zOe3Apl1I0Fl9REiJL1kArmywzIHUmvzWBjgsYk1XvW9U6DP5hzy/ah5FDICW82O
mdZiOz91OulGKi2RVFU28zLIcQnREEA6QmGg7yO5NICY8Z0v1t7oWIvl0Nl1o+wo
3ghAo2ka4wvbVPYWyD9uwY9XoxCmRBSCm1n3BgLZZAnu1VYhDdN02esu5FutmhNn
812h7rsOwIZI5xnzv3fqnXAq48YU+4Vk6hVOtMp+7Uvw9VyC6Mu5Gl/9FtYMt6kz
jBi1PVmxf0LOkZCU4K35n2Lgz2MZIlY626CH0/UNUkGVRezb6RTGU40FFTh8ZJbS
X/XSUYPq6pRVX4q25mLli6m44Z0usfBpDPdeHnrPguvx8dHucQQpanAHOJM8RGtm
ab4GMNWECwYoETwP3N7Vs6sdoQSftrJ6tJT8A5LdI+qVzFvKKYaaSacT21l38ycJ
6NjZlC8cOP992MwQkYPjqEl0eZz6BV7uzLrmIo57G/8SPAyS6wRV2RA0RrPMFI6O
12uyKyOJUWasQlNMCL/YCGh67oGGqvRMEy3DC4oFkBzgYigFKckMhnDmajZ6a7sL
BrGjRClhGnMtmId/tJFsw3rpBXXIt48vtS9Qx+/JJ2aiRArhyp79hJQav0BrzgEh
coOYfUXFvS93mncYMREqDjYrGK7OwgrNCzc+ekSPKcNtF4qcFgkLmOdoqAm0o/gT
dXqfOL5smZTWykwA0XgNH/H0KhXJqWaTvSDm00wE9iGzzU8NN3Xx+z4Wp+I4SPU1
CVnwnVstvELc74IlqhsGM3Rpr4PEnmCBn0Nu9ACf3og/8hVzMPNVup2LUrG9WsLl
ORnNy99XDNxhiJXPvobAN60ramLKTxGanKZ1NY6Yn2x8WUmYN4+hG7mc38vsnyqu
guW0PqJiZ4NKvoL8heBJdhSRCWqw4aeWK5puTCBxfCHIe5pdRrPGAsnLsTlOp5Vr
bEuLQPOHxeZsp3n5kySGCGT5xgUgcsNg/CdQreUoRb8lscRtZJWqAcS/hrLrLuWS
Z/HqyW5f3D7DXj/pX5A0z+saZWQQz6L7PrF9etGBldrXDLkF0IpgyLN7+TSbbOjW
xg7XIjHYZuWtbBZeQupkdQLDJSo1R00OJwCM8hKnnCTy5oCr4uE12Bq/coXZvuJR
+Re3sILawQAf/MnYrcv7G7HYuLq58LH7oPTQnBNvm52NWBXYkpaprJYEtbV+dUww
NM3jQzwHRlMlhqugeoK3Q3Rs2dQl7Xdkt0paqugHgHcRfsEEH5nnX0TlencqRbFu
H3g9Hi360nfkCNf6f+Y3u8AldgwxerMk0uysbcSDGj4z9Ic7vDNK4p8tBydNoIPG
1ZxTU7rCLrUycl1OGD6wTrOq9NVtPZz74tHf3n8XCk7kklxJh9MXBWEjLHBqdEtR
gsQe2ukzimlxhsbHOPe7XMUpgdI4YShTJkxRTF1bB+/iNMCPMIDNYBuEVdsXxL7S
KuyTjPqDZb//HeQ7OZgURUZ8fyrSvGqg0TIQawaULoZskEiV6V8nNuKuMnQnxoMH
cHDmmQlwmJQTSEa0Nw17FG4BIqJRqFI6YDZ1ZKjtMdYvaDZYvJwcvg0BagfBFwLC
ghZnOW1wwvQjRbwI/1BcAa0iqSXszfZN75n1U2ZkozaQch1G69qBPZd0FlWt/qtc
4xSjpZZFRLZLvxPhsRO5OdvKxP0LyNR19a9fj2zKPKcwI0KjQH5RdtpBtnUA7v83
h/emOGsBLcSamIKW6UkWPhhfG2YRU+54rv131xYJzevM4G/DyFeA1UElVEOi56ds
gZ2TGuZ5/YLlNZxA8dieYilI7bIspFBN78Z8q08QNxn4elcn+KIynBNu/6TEkQM8
AT57zzWlFDd4xNbomonaUOAZIoMLQ59FNM458kTPNSrMyroIbYmQSqoneCxZItd+
N/XuiOczK2iWq+39+oiCPhi5Cla4DjeBjyphMdBrFEsHYkfp58rDiwbCgY56peVM
1EmaveyMOzv6cXc/AAWtEh3osqnofKu1gMvsDqKfqDJPh+6qf0EGGm4oB3GbABEP
LKtRph4lD1I4ecwKOS5KoQ3fCTFTEQFFXVhLimBC7TJLIkkhoJhdahY6zoITCHrH
0mmiP4hIquw1/lxSALG6aabcYkrIjKPqcMw6GTTGs3qfPXUyDu0BZWxGEqgf2Uif
Io9aRjMxmOJnsawAoNlzlhk4BejhOOBIzcWL14wJmBGY8irv7jpYG1278kNGYIOA
7Ma1+D2McIqMVKkuBmAv5WESWzuKC4r3b2yOcc/aVVZXliWqjvEKVhxBpuoLWtdm
L+jQxs6lgilctgcJPRju14asoY9Hj9cD6S2x09T2fu/jBZDgBfwuph8kSOhU/Tn0
90ocpVUgkmKc/hqT66KTpAyIIGPjnyLODtu+clHoAeY3BJ1ATYi5S+rRKuZdKb/j
bbuJaLTggTBdUsXBeVe2jLbQzVY0OY/tJUKC/hy8oV+FgLgFQk4bBE9aEuX9lKUW
NTIUe2fGdk61rwUe7KJafCPcGoa2SMK+5VzywZcPH+wbrkdmjYMAHJEraZxGadpv
3AF8BSpuWFwJtrBHhLgiAmy/Fq8EWS8r5KPeiR95AR4PG4qP4zWEA3qda05+ZN8b
nXTfxRa1t7H0fqOr1nKLfWv9llyw//3T0IyYrQq9KhZ+9NVkC/6/ity7/3W4jJWG
5BisK12Vt5ThKuhcgSYe3pWMkge4QHK0Sc6G3zzmqWgsezB+fV0Y1sZFeL4s1wm/
QrYmuoIEAsrsRYd+VdndM+MaqODhsaCFmwoVujqpeZE5NxFbzOF/J4WSguyfUaML
ity1OuTWqFeCWCwtSJHwuBABdToVm4WrWjvR6LmpmMnPcQgb0RqZil56RB1f66Gd
zfSe0x/7v7Y+c0pajqETKfboqIWVf1JhTTnoBVq2Nqq6DjD/dMHqDQWbX7vk614L
h9LYnxpqb5V+X7LvkOnB7BP5wXE8TVoQoPrn+/wLfo5l/JhJw2gsCMQVCG4yRp7J
E/37kA57dOVkb5fWF8paWpNSMB3oXptgzB+SGwi7zI1DQ+ydKigEHPt9DG+qvO/A
rOV7ymLdoMq8arPMVrMk7esK/auxqEfQRIogIVf1M49turXbHCpSc7+p+g4nsIoR
tfCYZPsaawYcrKmBO54rc9HgQugKJdX8yRII5eEuUS81Jd6XZDizJ8yf/WGd27gj
L1uYdilpIr/b2LpdFEt11Q7EwGEc0G6HMdckSgHqoqkor/yHFrK3z1ZoM25xvXWl
VpOGcqJcxJ7I1czwQdaalOfoaAT7hzaG9fgOdsqDY0ILDkxCGEHPh10diY/+3WpA
SQ7WGVo4SN58PkDwl7VaMNPyCQ33QVledLl2uS/PVLqMTZ2y49jA/mQtK1m8qQ2u
Sp3ZTcE2omMihpLSGLL8Y100TSjWtkjCrJUla2Ank/NZVCcnILmxopLZSjnY0c9d
hE6fl3MwQuv3PKc9noSEzgHi33BXTgZ/3C7fM2HRkI+yy5uwoYI3HHRdSf4S21h5
FpFHtyts7xllATMcR7WPDSWVkIjTPIz7EvWOI++IEIQGQSO7dXXO5/ffg+G7m1+a
zWUbTdNODmfwq7hRjoQsQRRW5DNX8/sjlEk8Jndl1s6AoWayUvOAkvpaYx4QiKxu
FBGZbpAlNkz0TvfmMDJmTeKkIr20bTvmN83Byq+EPijRAP9s9w77Lb4/WUaXVTEy
+wsz5EttCt+QrI2m4kGS2rd77DTjGlKuhXAQLiI7oHiYwntOXHDfCe1cZxZdSq+T
pbZrQyBC7VSKkE1nRIORItPR4svonEhPQB6WyOkQiExq+BNnYr8uJZt7ZIcKG+Kg
7/djqmdnPRTati2iQlQr7uJKEUskSsR3Y9k9xc2J7I6SZPjl+01S9HwUSQavAY5e
8mh955mOeKdBHVeAYmUe9JOdW7ea9Ir68dPTj4ByrPhr4SKWxkabpBZbSPGlcTWQ
8ipOpPu8NeVA0lGUOQeoHMgxrE80b2eKsNOw6TSUFEjB7pDUGkb+P9O8GxcQnE04
TE8s087kJ1jzY2pBnERw+8D/9UX/+sMQiR0omDzkmcYSWuen48BlQmHAXqv0KQ6f
rN4O2dcyf/N/+hjsJ0NMtsGvZGuh/A/UoOretd5rXoLNoJD//LchApbqgw7U9k2i
kqeebtwcGb+WamYXeN0wLlZ/cRjeiU1UTl6o+FaJVm5QnAHzfc4Yb7aNg3AFpjKf
D1QVF70JUNkdWsWP22gY3uwftNOek+liKe41VCfU2o8lf78ckyRgQyJdvods8yoX
Nt8Djvm4WVlPxj1C1e0YEbAOHwCg3tdGXkARVf66F84IQrMLsXr9/p6GNau8DAmI
ffDktnWiKeKSSN4Clbjuf0Sl/5cnhL/eBz33BwWHWcVVfPEiFjzLrOxfe1rRRU7U
AAVVbjXrhusL4/46GL7OQS83q8lGT8snCAcgdpFSGnkF8W0DPRpKxS6i7f6sJ6tI
SIeu9UzCMQ3O2foXX3gJ8/oFyTslBrAhrYpijS9AR+MBIQSJQklbD++axu8EmYX4
OncORH7GX+jW3aWX1mxvCuqIvZAkswruujSykHptB2EnwnBOIs3jymkFcGkIffyO
b0UKSZgGaKUMi9RIiOE7i+BS+zPlWCiqY+SVBkH78wA55Rxt9YFg/C+fQQ2xyDOt
wGPDBjil4f7n0YQ38cUE3zlX0fZ873Qlp8NWvJu60mVgt+nYv7rvYBS5Hkq2hxOK
EOfbF2sMLxaWf8J/KmeD0ezdThlZ2YpmvT0Ln8wJoLbhuKAOZ5NKlb92vpUkuOKR
9X4LFXN8et4NYzlPJNiXT62PE6zHIrK6kdCkI8JxRD43uqZf+F0vgE4VoXULD/Ko
9/ybvZD6jKyDr5Dj2YxPeeSRbOAbjI6wB80ZtAGe2K5dHwfo1j38UZgl1eKJM5Ye
KQrQKCt6NiEyA30MjGnWzye33FOrHuKrAFmC+GfbplZxoS9YSEi+ahzBS8gAauMM
iXQZlQklIl19dTtc5n9QjOJtqr79HYKlGXHhS32/jBde43tvUV0I/EwQ6PfmX4RQ
5czvlFd7saA6pEirnok0nwQdcZsB6x+qOB0037y0LcIv7gQlwNKm0EmGvIeufGwm
j3mmE6qsLSduQ0NgN5sH/IQ75j+dyi3ur1OMNkW0F+x2KAtHYnpAveH91JIcd2OT
kUSzMwkl6P5bUnad5kiXPymUv5Pjzbv6TnCTSKTINTy9r0LKWjlwNEDde0/9t9SF
Untjc0NeIkn2ro+POoC6Jxvsvc4lZn/2hgaKenPrNEREjXCP0P36CEreEYC6NwXl
HRmrkFxihUI7A3uBON4FStYCLC3K5r+Qk175AoAjUh9RBK9DBXlupuP5GaTkWf9Z
1Xiig5ukVE83rge8TeRPm5af8gHe95JDLy7w06Zi2LL4HyI2aasl8OgzuQ7vtsAI
ajQzPEu+zX6y4NMQPMqR+WMHfN1U5ugc+K6jlpW15uH/w7F7o3vYtiBcWqLoO9kk
dMyP8NzZ2DBrXOLgXMtsc5wzMc0p/OrEXLZ4SpbkLWyT/zYAWkj9ri5JFbIeIjX0
JOAmFBaDoX6C58zDwk3gxeALycXvMiJLnUg6hUiE7C1zlNXimpFtYrNOyCZA+5Dk
44qDVICqzggWffPJhxgUYC0DWG3KXa7V+HJMjczMiY9EgI+eGjYPNfIaJ+GYzazO
s115cmhQ1lQUpURruhWqLvZb4GHBLODJ3IX6qohqtogeURmYEFP/llswfY3E2Iok
5HpluAGW2fdOKFI9R+/8kPrSpyDg16gqMBLteJiu645pjYar13cXNXkfGP6nX5Sa
AmWL33ISWjGb3pcA2aOdG+e2rreMx7UfjlNS+XGICZZaUmezk5OQ82AA8HVL1Io6
Q8BZInfbO1vbJdLzpe2adWLwo/zr7hfGNKDkEYZ6evK0LAz23yhWRVFh8tzLorS7
s6auqug+aAWJUVg91+WMia7OUOVdV4wy8TmSKqc91pZICS9htyBXunHSl0Mr+UvY
P7QCvLxlqQWuLauDxbcHa5e5mdqHy/vAJ1Ph+ry0ZapCf1lG0zD4fsVB12bLf0do
oLywmD/NPPNmfIDLidCUQH5hJH7+kN0awTQV1EUCjUjIArGiK7+PhZIJSf5qdwG+
U1OjhOvEpXW2eh607YZoI+AYsSAyqjUwctKa7c69jFjj11vKDxD7JHeQIrO/ApFC
TlTpbtSdeYgwYLaSdEo7DfukrmQNilIEhEzh8MURuLxpwTpV0yofbEDdwmzYeH4S
EE3OLZz820smqNJHsCdmE3uzLuTzcoqBFWaTa0lIgiugNjVeWD9clcEOe4gm6sbm
DZwmh9YlARYn8lyUMiN8Lg+x6QF5jskxoi7f99AQxKSeuB+cggEUw9QgrAOm9qog
DMJBXr+WqTbOw82P2Qs7ZfdoF3hzVwAEHsfqbw8I2RCLobghs/7pj58PRcV71mf8
ZZiNlK6rioDASUpAWp1ynIk1DG9nw6Jgjb4vdp+hQrrMQOs5bWX9gdQvWWZ/eDWi
grcxJTL6D9MMNn8y0a2zBHiSkJU1DwiGhHP3MWdaw/n/sa9+4+T16AZqgCdkllnA
hZNfLoY7mhH7efCYN4l1zIQmR+qjFrQCYniXGMDNphLk0xYGtYR3kgJ9i8YoUIBI
wwgn5QmLziVkyokTDTf9YopE2WZn5ItZblHEY4m52TKVwNHHlWYwOl+r161EdyMH
sg84nwXlLJbXVofFwSvAig4MebuCUPKuCJ/+H3AEIH3rrCYKZJBUCSL3fwKeXJiZ
JJx+l/fLyZyAmAQj0nLxfE0JDj++Q9YHSKjrv2LDnJdYQDO7b/p9nA6/9+Mr88FB
5w8SgsjpkrZX3A8MjfWPihcZCR2yjHO9ficA60SHpeX587Zl6wJjyHicLpoW6dki
Ghg6jNjGyss+0Eic8uD/IT/uS1WRuIxtDEtpx0EZI8/zLkSAcxaCiODefNWylIOg
ErvwKIzK8/8sRFJkSMtUEQi/i1nsSNNBx+oeTIQqdPSwkJXZCf6s1El/ILb6Epgh
8SWFkARLQ6OHbpu31cytz4WVA/0nP46YfzAuDN3ceKrX5h9I0rAcqNNnZRvlDhzc
V94oPMyx1qAsUxMvZKyHHQI5NSRALcV32IeXOos8cxcpBy3viNPuEgyxxir67EYU
Q3Y0Y5OyZBPCYB1rQRHEvmcPdXEH3GziV/CK8K6PuEj50enrYvK6W9MXN8Pe1701
uZx9ayS1aA1qCgutwk72u626GRuIJv5kvdWbqeevJsx38O2Yw1B1bUO2rB/2+qi6
I8naV7GkNcgqG4nSmzf707/Wj0XbLBtuioZf/h10HsSMZ1rxBOEYYfdBRrjsHYxu
3c5XHcfCW4i2zrgVZ7WTvfdkUU0P/iZYeh90AAsxgJF1nRSvWXJET1TVbPOQt9Wi
1U00/XQ/ywnY8JWNcLtD0+gRxu5/B0DMwm7zk4I0Vo66XgN9BalCLRjwPw0wDmU7
zxvkowLakIwx2UNEwqwGdi7OxxuMYRocHRe0V/4ajdDxwOpYAO0wVBmVQXUKs6QY
QwFj4TokoN4qR+UoK+JAMazFR40xK7nwil0yJOHoMMzXViSaZ9xYXpRATVlG4y9d
t+0I+DGydbiPrKqwWneGHdSnPJSwfNsj6Ba5VqPkARNxJ19XvGaoF4AhDN6ezBu+
BrUzWwkoKD+/zp36qdctVhKUP8Sw0oVaeluwjKmPwp8A9HK8/cgdeaKRzw8Xvpo9
HYlC+QORvBeRfC/Y/z2v47pmxVPSSrvOPjIV261D83u2h5ec1QmlPv1kHEClwiZQ
pFAT5Qi8figGHU9Z1Gxq/eugfkkUsFoB6oxEjcCpn3cnvM1wvn33awXg9Ml2qGCI
NyWkDCYmx6085EsH+50oLZgvAHzmRzEi14AQeRqb6414If5+Ob7LB33YxZe0cHyM
qfSS1QxQAw+MCsMeO/AZybQE7rWoJFFkOCC9iwPtSIF5Xc7a7as9RklaSZA1m/q5
6ibvqezYiMiWtYxQBZawdnfTVLWInmZXxdk/DH+ravHiQgMRM7uVE+pzLQBr4IKA
Kq61FwX2P70PGl9oPodZnnzzCCV0aDvwOYOElCcEFfPM5wEW/9JQlbcUwWk3YsFP
Vbmu2W7At45P6awR5uwfiaxmr8vMsxuw54iasYG2acivLb0Ijag9M6S3xcWefku4
migvmFJF8OgaveaCsyc/DFbcHDjiYc6lKTezs5d573NkxFMYlAa/Xo0UbyyqBhgN
y6rliIcdUkqw5EkjOjPsGTD08ojpZdqb7R9euu/5RvwS18tEeC1I1Ip2t7YcS7fG
/NvHVjNpreIDeq/eJujyhLe1YWf0TI5OvC89cSpZIi4znbkygjVF5ue67jkzcBNk
xUryWC+U14U4gLepNdFdpIYQtvZACRHowmNuTTnbBg2aUvMD+ZRajR82SsXr8ftI
QAC5yG4nImfbWFqmxDB2f49RxQRm4ffrshXXKcIB+qU7lCnvieEBeNRBEok5MT0X
Y4vuNq9GzG5Ft7diKXkXwWDMG3l+UZST5JkiCjhkXmuVpnilQlyNrNYilUjnpNdF
ndpMyFO24V9KNgrjaT4fKhAzyThSEogpSz9Z/zmsh+eukZJ3x358CFPwYOTRN1Nw
n7Uk84NHrzFBU7ZRz8rfCcj4+vALdQA5RZEMpdjOQH4oHzkYyArxcS8TXGlme1wo
CaQmQ+Ri4k5waJu7Sdv7+lHx6tx+8s9h6n/ZReNymkYrsWqGEO/X7eKGM30KLV5v
A5PR4Eydc6XBXvn4ILykUjTEZO9zsJjL5KUpyaB0Ms3mzsOHIBlZ6InP2d3xkxjI
4yfVm3Xjf2Yc0k5bu/zww8MtavaX4o/kNZXPP5qUoFod6OVS0VP+mDEQcJCpVDyW
qylzHg5/gztoWWPwPFp/ZIb3byiGt1xn+uEOl0pSAfNnG2gZwvRd/sQ/ZVHmAtcf
R+Bi3Mr+hQFlanN5E/7+bSA1cLnKJbSGNz6UJ4nnaj+vpklC+49jCUMmgv5c+4Ct
ItoYKgMg+iW9XpjpVRQCjiPewZdhXoqWVgvUXsFRLBr64pijHz442RKzP3yDJa4m
eM01qCWksBcMakQuSPeqvA6KQg3rv4U4RyZxgiDeYp8TS48iFuGRj4D1zdLMAL/H
tKYX2wFHhiMjhSoEVv4v0WIXa/cPxc0mzzw5xerjoUhwp4Z5VTQDqupcJv9EIw2i
RCi+wW0aq/oIxoHlExQaUIv/+gmoFl2h2ABNqfuwsY+2sVZ80KrEaWP5AnkqIpfV
MrOM4YU2uEdHsKPXrbjGdNrYbATKRR29n/SX1e5w/EFT+z8lstMFaXopalvjHkz4
/QJluXF24Ad6pwesUT6maN+PuVsLn+Fh7dKUp3U3TXp4nJ9bj7aPgsqT4gDD/tDR
yBjrlCm7IQPcbSeRZlj0N224lwljVrbbGpeTBHnyt5AJApmgyAjITf/KiFCNuu/Q
/NrXEwXhBcO8WBhqniDZnKrZX5SbQ/xbfzKo0InkNvULlPzCU6XurluFdoYW+DDb
e/slS2QMxX1h3HlYIAWWLuehjpO0wexClUOPnaSQgzqY5h7P+QR4H28WB9dkC4yM
cyZ82ms8MFHzYcgDbHY7v5OF50ko0sneRgGzS30yrsWWCza4HOn6OE7BVP4tG6Dy
TxDnog7Ele3vYKkg6/aYg05s46WxFV84npU7WpVobdW5INsu+dOGOjm/jn2P47V/
YyyyROlaD9DkrYUMy1hoPyMTYz0XEH9s4jxiaUOga8EMKjHzkOuo24o1e1KVH+SY
55zKS4yNrzX2ZuFHVIWN6KIg/5DdMoK7ZP/0caA/HAvYY7lsy3oDpwkjulyIqFiK
HzVOiKiPhimkQksAocUS3Fp8RGQyp1/5+zozhP7bNlCpIlzHeEObk5/9gA5Lw1Rd
QtTGTMwQDs7vp7GMLhO9BfLeoHusTWaJfYAXK1CYV06o3ClMmEQJACQnCKiVoWCm
A4BRkOQJmKIxeDApquxUfSYlpEHAUtr10qpx0oDRkg7SPzVLLeeviqQROvdOmoEb
5Jc7Mx4v8WmLENa9lWXwnLGwuSXaVXdQAIYNCbuYDUKZ04uJrMbE8tvyZShcmAff
nyJVEZMHSTP7WdhJhHfM8zgnGNJb8cWgEO4dByeISfypuci20N2Wx4FMTkjyfeEd
7VzPUn3jVqabj7PUxkl5hmIRmHCIcNKd13/hQ0fMlrx5iAvmkQDhO0pCrYv9JAFV
E879o2FWiN/ZmX7UVqSpmb+jid9S+TEp+hOOgEq467Odbf3AmJmP7Uy/E7G4j+SZ
id4cBSOZWh7wd0jL36q34UNLGwcQGEaW6sKEBZf0FWSfVqJmKSST8m4yugBZ4nzj
XQw2leBk05QifLQmy258QsJolLr1QRIekc8lfY7jTBX6/PWh5P/GHV3XkmFLbZmD
q8lvdCNREY+Ta+3yoiy1UC3a+IVGnZ9QuRSmLevc3nR8K814bG475C33OiYErGh/
DgD997ArWvVZwRpRrp8Te/6ZkcN6SxF8pg2+p2tqxF/QiCiH1AjrQe8JABWZa5mj
ohtUOwwztg1XCcnbYxsPWbkxmoaABbmOgb2SsbJ/y6tiOrdCgFelLJTlLPPoTCGr
DQDYG8LJR9ibXSr4HeophVGslHtoZm0lSL6hWyBXtXTTuKxNLi3MBagvgP+w3uqX
D/6nUeknrdCg/S1tlu6+TurNehIkZn8BtXddf/5G7zL6e9602Yg8a274lN3ZXLrc
8G9afFR/0ajTFziweJLHNbZAlZaGXS8ooVxpammvf8VdS2x/yGF3FEUfNZqMWrna
3m+lcG9S/h2DNMQyD9wCDHxDqg4NmgpjL4DYufNpXSs6/RYHDeHO3g8xBevIKDQ1
rwwOW4VqVnXRGvgbFrAWbsjkKDYwTy0H8us+sWABfh2ElUoazdqbDDd5c5bq0qV7
qkEbDM8l9sYoun0eyy6m7BpkPsBQpSuaN+Nqf/hJEOCnrdjvq8TNVcPaNQm3YTBE
MLNp2BOwHiuLGaj2AL1omPs+gMFLyZFTQ+pSixgpMhzlGTIam5t1amMiv/7AoW0C
uEjQeCLGIkJhowi/NK8i8VE9+Kis3Skh62vuyU6uxrLH84BSd4+/kby9MfVq1hJb
L8FRuUk1QLZXDo1dPv+NdUGw/0T8KFw2SWzrs6lBJZwbrMd27hn8jcawaK9pMOx9
kNEce1hUD4FYbI31PjzMaDnKJQYHHF9DZ8wh2+X5k61ck6yO2kdCKiaoqdo8+CVD
VX2HzGv4tEq3cn4LN4wX8MigzrpfBSzR+lluMkky4Fiqbw96AV8jmiAUuVEyjnD1
NYS9Q9ssMmmikCIjaob6AMkfdEap270OD3CB8ia1KNGjcdRpdEHxH5xmGTsKAu1P
AnWoAV/3ZSx/M8fue76a/hS8AptBiNz/FJzhwdvVCqD0ODhsyfXYwBTxqa2ZpZJ7
3wULAkXtYHTwlQr4VrZPmztgEpv+kVMqOMNYI78Sk5eW49m6yO1ppWB/K/n3eGvs
0D+sZxJT5mUA05TMoIcB3EJVaBGlc6mBhSWAni5aRqKJUNs+iZ38Kf7bsdhw7RGS
wM1Xv3TYrNTBqmbR8LHUojUiKf0EaAtPrC/DAiPdcgpFgSaikkpM8EE3nexQptx+
WZLohfUKXWR3IRWdWZ5Aa2jbHBiER1tH2FYke3Egq/x71FVTGuEsxg1EijL+CZkj
ej/+m85SIhECDMQbmHc8EGodNHMQTw+uLG7hcVE9ondyj60q4W3m50Q3djGO2/6L
Kn2o2IZQcpqGLKJe+iNTGaWLyvL7Fu39CSTAum2m4TiUAk1NKRYDrPk/r42mbar8
qTtsaozoQNdG8aofFQ278kvpd9sWqAjJiK4XoJihaEZVeiFy2qA9R5un4e1uSII6
5haSZ5bcjIzmAagt2Zr9QD7C7AEJs0WgJ3jNiv5aw1IkOZ57bZab9JBHYgHaZAby
QR7+alRiitYAdPevMkVBxKVV6sNnvH97NBISUAz4lUcVPoaHt8401DTVfgExWSR9
IHArjcMJQzHbusZJYwLTpbbAHfqsU24HImd7rblTbZE+OEqjfUrUmNNANReLQLHm
AGLc36HWjfRWPKQMFjER0uXqF57dh4p/fqFcrwYw/ohEQ/S9RIzvUZsuVs+TXpse
H2jJnWNcirzRo0oqZ6/Qv8MeMKiAly5JpWacar/COterKZ+1FD/WbTOy4rz6rNZM
qwO8HIET+JWOWeuTRA0CJwBb1YWnhL3WWjNdT2f9r0g/ln1j1+zrIf4jBtjAYmz9
FjVqcWfx9dNwukphpKaNNM66d+TPJh1IOkyH0VXYsjr9qKYk4evQ5DeKpmot+uhB
MOVkWM0lDwTVP48Ye2kZACsB9ZoGsH0nfW2xIeRznjy/RNtIF2f4dt5u0Zhpojr8
C5Lz3FgsOWyF8T+eRJsIOUa0lXlk5EEMvAE2ih9NfReyRXebU81j05XbkO9r9kkG
k1o5l+CEmyedD40cYaE+HbQnFW3I0zxTaY4SyYGcJyISH4+/Y8/qAvOOMMigzP7B
6snYbE1ksa3rFl6CHxyN+fTPBDqmgND+HwPGR44Ggl5FBm/SVg7/6ytM0F+dPhNr
c3DtZs0/2x4zciDvZ/uzZjiI885RjRVeLQpqDFb+iqfkje5mxm9TK3ujn3ZR6vrZ
xz5UjK9vx1OMcLjtOAL8PYN6N/s/2w9rKdgVJxIdpf7lGimwhHVPNhU+nd/GBjjQ
Q83Qt4CzUDeDQw9F5t/DSYKb5qdjk/yrB2a5E+EeXeDrjKdR+qy7WFSgSL2ticFa
6VmpuyU+UVi4HRi+ZJyJOYT6qsXgvjrzlSh7GPkn5VF9rJnFJ7eA16Q5M+sk96jV
jFw9l8OVG19EiA1aIuu92M42CiEg05ibN3ApiBd6xv7NtQ1ap2RuRnSCpho5wrLY
zvFhA5/2KdS0jvN+TEh0mRg0688dA22xNIqWAH3lLog0dTGwRdAH/6epvKK28Rt7
xyWQrGYRUIrjsdJkP17SgZwTK8I7DhSFEbh5Jc7AF+ZdYXYNVC2vgDe706sAxm4U
VE7CiLWQVzD3iiO4Uh8i235Q4rNg/EGhypiQAsWEW6ziwircMWhddiht5UgLXnS2
C77ZJB1RVQoolrt5hzsg/LKIph1EdMS/KsB7IMj+c1L8E74/o+5pj8pqoEIH8dgM
IH6qQyA5jd3pBOOog+QF6sQRbIeD9ct+7QbFQQKHOtEWIpe4T5skrvzlyqSJCPB1
gNGgrazKHvawwckvIbczOcVSfSUx0A8shDTB97b/vxzNjsZzROMgT/+r3fkEIAOx
JH1cDZNknFTK9iobemMuVhIkV9D1T9TwdUXUJbbrwpQTE9/dKwu53989MOrq1UlE
546+EHyvlIYKY65LYjGqV1drqPbHhDgoaQ/N/2J5N/Q0FlBf/7JbGwJQBfIUhgOw
e1XADtldHPScHYj7GshdGlKdrUGd7naRN3HUPNAc99TCVNr7Ml6085lRQy30WqLR
+uiJTpW9GVO0wOmFfJ0QGHCn6bRmc4EaPwK62J9XbzpLrKppaERDEVkRINW84eHG
/LTSW+MjBBM4VufJ6TfiUpfJmf+yWqN4JQ91I8yXGzlld6yUfHGHYk6RiOuUq89t
99mJNZ0F/QZzVgJ19nb0hbmwSvqV8Q2z/0ZLaomoROi2vYMAq4cpJGLtNPDvw1LZ
U9RSDAOYuLO8NdVOgPy1Gj2mj7mgoYyBrQBKtg2Q5uYi6hN+Sh3gy1i/Gb6fds1p
FRctjBqERsXea/d9vXz4kLJXj3tOk0ArZBifCPqDhMBluEdPyLWf92qr7a0qRBbJ
Rdr621woEY5aLI0C0lnRRuZUnJeNrWOCIUAVmN1QZTw6zLBKB35l7s3dGs+jw5ok
N0Ve2hFlTBdOLrOPdYZBfeRh1+gDi6wLqHtPyzyaCIcQqQP1+Rxo85d346PWtPLS
C+El27APvQ2/ptJ7K+fds+3PMfv3slLO58wJQhyyQKyqvGQNlUBDejZCHgzMkAdi
sZPjTgnC9odZ5VLps4XDtEsLVjMwvIJHBrsi64kyKxdFW9f2Y6AvLaF49dVkwVls
jTteVcZu32kMyH3KFMilkQXnVc9oIgF3cYipz87KKeJaRtp5tsuyUydisH0lb36g
oqXn/3fBMvJNtf71KqLEyXYeBOY+49xE3K3IXenpz53hURvffATYVuQh8dtinoi7
A/514UvFko45TDRpJHjrbJ71MDcFaUlxCR5DObYrBE/Q+ImatidfjQmz25qw9aLN
TrUf3/PG5/IbG6BeXuKaiD/h6r8EjGHLRRp8wle305O7onWoq1rLGbWUoHpFAW+U
/EwEDeuQJFctw8Zves4/2cmSl4IdWt6wHeyaK3mXUMY4GTAkeVJg9hGlnMTXPccC
ATaGX2OwvO3dUYHhpHf2if8wdv3r0Gh5n/dNXzQlaFIwy6DcZsqzgbUAYiuwKDfV
CmzZVfYiOv86RQZgJ0qR9U3bndEFy9NNRkGZS3oyoJ8ifTp7FkDoiT1yvHRRuxHi
UcqQNtaNTOHXnrjoNs7HFDckNXgribDiC/eRI0hW5THZ3jXVqpGE2ZN3rSSWry3o
T2bSA/KgGbD9mrE141dYFjKzFMLzKSKiVC/5hEgbu6YX1p2o87YGo/PkEaECBEzb
Baw5ySxw1eyqxzvMupz8mtxsnZVfE7Q9P6NmYatizrh4Hrap4ME5rkpxlklnUph9
LG9nENC4QxAA3PGIWmEid7+IQgja7jJ3OEuXn10rPAcjFT64LRlR5QJ5szRwuQlg
WjhXcyRTa19QTfBaURYfzMiobWUGg+n9hAOpoxOZvuQP89+f0vK/A/bxhI7vekE4
CpdfZWzwD61YIQAvAyM5fYE4bz62WlisQsvTUS1531FwlaLqbSOOsUDuix4Dt42l
6OE+s/7YzPXuoFv/yr56fZ07e1OaIybVnHJiIT8nk8T+HZfkPiQTArT78MKET6PW
bKTcaIxuQp37UtXDbT2TRcUU7ROIB9OfeSBwnuaP1P5VIi31U5IJGAo1z3U3zm5o
8AivPr8fZBEHnWKKLB+pdGUbWzQGb0UXu9GYvZkRWSlmxBS0ayg5pDjGdjxC+PaK
Z6W/N4moG3H5R+irGyw1U7/CutNNde/OfaZ7uwx3HhZXtfLAfzq13tCZhR/1m3xw
Ym1+cpBgF2ufkXHkd60PcX+2zI2YjZLHGTrOIqsdLNd/py9tfmY7KMMjhhD06myu
BfdkyIvb3cKSCjAYLrjgU3ZLOEKmSOv6ZFFlHFtzKqSWlpwutEh9jy+NjBErx027
YI09a26TqTZ18Mv9Db4NrMW0EdMOorXRrebj8EKpuTlngmY+IJ621zIvA7bEslr5
oMyY5BdpSJtbHFu+ixFbMjs7L7Ns7QtKROtIQ5DV46OFG+p6ytli2BgX8Ggx/4Gh
2dT7X8WpXsRtRFUKD6AHHDP4LZdWYTVka5w3g9J9MeA8vK4TmmkNr8i8r9sGoW9z
7Upgj1IAQKMPyj6Lg0EGEc9NvXm8SPd78AV5cjBDWblmYY3ex39ODLXpQRSRkv42
1OZhjOS/xv59+WkN4tkTmV6S04/+oGV/+AfgwUdstKJI3c2zgqhZEro8BdejChnd
lsBr8qvs0Gh+0uMIrd/s96cZp54QBN2pzZkm/XBbz5b52MKxM3oiUMTIzBps4xQd
tCxdoRg0G5UYSiKvub35JedhOdV3LhwjatsIVevGyz8wYeQGvPkGj2LHSoqc5eu0
khx11Mo5G6Z56MTt+R7cUYwoEFbhDg3iDxh39EFG+YlG2N2NbgAFEBpiy7nlZVqy
8oZgKxlSfIaKFedNCy9ScR4LKucrlXBYN54xCHIaSQEBqAuYKbZWxAqGLTvf+PwX
UWJlRwepgw16hFyu2NCw0tQjKA/X4HuOMn2OZo1cE5kkE3XzCN574szy4lKDE+2Z
3T9z/aFcU/mOLbNIgUHE+ABhsc1rTHoNS9kYXIWn5Kpv6p8lHPsViREFI5NWf7+V
/G8XwKocAmsNBED7qby7j6yKrjf/Wk5ttDJGtTbewDPUbKxYgOEBgSIJMvWsX/TU
60XDRAgPPCot0XmkFDG0aMBsQcF00jUEycLmb0vvtt26cXGcrLY3ouj03EDoMbyK
z+RWSo6a5HdPB5fF9XxZIG6At2CaRfiAUZozrGCkdKffFl8zC0+VEcb7PCxNDnsu
nsjyl3Aefko7SygRvsDAlJ8y1G4t1mCvcf23/WE5hoL+uiOq/sTZDVu0wTxnkevG
Ds/9rubwH1V/TNdfd1OmoZv7jQ5JvWbHDQ4o5JbsNqZg5xeaBt3fUPVuQRcWsSOT
j7/0tlIbfQ/6TMbrsXVxkQqnCXJ7SrnENPuV7/zSryG9O2zmBl9OcfmiRHjz+wSv
Ot7jCoY0q7lWFrVGUxhIwpqs8dbCmrFRmxFpwUpnz2lFCTRjymSlYsQ6LNXfo52q
IvCOj1mTI7vjVJQHWztqTuqBY7US/a6Uz+bob0vJ16z9u2vGofEbQ+b5WLfLHdNc
GX7oLH2Ti6SO1Rz0Lv1ctZ4uN6XtlrEkp6JfMuU236RQfdKtARmCCVUjv28Dn/3+
wMqFmo+TZr/ohQ7i/5BN0PjcIiCn/15n7gD2zUL9uwZrBr3rIvF+HC+kDbhcBeU/
R+mYpPOQjWZLk2kjUequh8Scx+knzW8CYqBC6ve2C7Feo2ZRgv5Ti/fAbCLNScWs
sWUb5aDqcw2mI9yeJA0OgXAtTVvHl3GHGkLXKLcbyxUcS72V1d8v7TVbRrMdQxBl
Xvoxay26/tUOtKFZYk8+DPWVbXmozo2EoQZYpFB0iISqNkN5rk4H396ZH2Vnciu7
Pyc4ppKUkfeunESjRB/KOXz1rkUolKsF8NDz2hkVpA9BxPRh5bkpmxnIdSu70LGh
K79GQahWlsgkLSxsns1UIdO/CdxtTSJp2X7Uqie1aGJ1R5auCk3XBjH/hWCT9TkB
0IxZgC2N91bCETJzL9YSwQGnlwnPfGc8MdV6hCXTieOO8nHvmBl7vI9WPCZRu+TN
Ng9L2rLG7qm+19Fs8GZHe2U+YJyR3cXzQtHgvXimZumMLpy7Vb5WLtN8nyp1fIrz
xX5TtSoX+m5WBLtbqEHPd1ePtQa5dvXnR9xay++R/X3pNMqZQtWsgc4AMKUbtCxj
6XEgg0oGX1Fo4aDlHQnDxA/ZlYyKXuOCumdL64x+ip3RKoy/DV5uAubqJ0KgjCUp
lwIVradvrPO0gNc3hcFmSQxFkUYdkeeM5IiAEdbdKldOyPUXiqzKfyIpc3DPdW/g
o9KbXFmqLnMDXkVCyHpfmXn2Mlx2YvPu/ANMOMd/yPE/NqSRYcR7M5KGQ7TLvorw
9ccQ7ppCK4pWIGvZr23M7iTvOnTRH+bBCjSfHVj0nKGLLt7JSPe2rf2E5EEJSSX/
BOkl3MHn8cZUcHhN97XWOm+kC9u8jH0jwEQjVSsSl9/ZpscyGatV5g7A5VtuRFUP
b6m8djHteY/UI808lokCMsgLDBDi0enHVULn6Y5Opb2w2GNHp52/vw+zYJB7qRHl
84oLdy+hHzODXaO0tPJkrQaFxToxLvsYC8Oa48o/zCaq0xYsySRojjvs4a2xzfTJ
EdlD85P1b/KwZOuQdkLxdWO0uhfDDglAGLXCyjGOJ13cijXgjx5OwMSoC1ZydkuL
LKui2Xsh+SkjiDtV8HtgL9R8jzRJwS4gxxcjEeIGdgaeED0ACyaLAU9ALbmGeNo4
6vFuPypcGBXTzj8e/eIzvTFlqq2vyMuj9HFromj8FdfXJpEACm6cL3K726JfZ9Mv
cfAfqv5a3IVMkdeWypUO+j4jJS6NZ9TXM+r6scqzz1FMRNMbAIfUu+Ryawu5Nl85
5AgnaP8IQg6k1X7m0bZvdq5Iq9TSRkbmiPhY5lTbzMgh0IUoZIRl6sRhBvHfkk4m
qGiRVFcHorNicaQ3yaseO7ttK1C5x14WpF28W1qW13/cRMfbJmH5rfMUukKuHgbG
Id3W0e8ThlY/PR/OJGtz1SOvmLOFUhcWZCYM+3Dp59BSJ3ylOKpghJ/bjTwnkKJR
54PSjuCD8qgW8u+Nu32KaqUWer+o3O1mXeljo8tGA2NuR7nAEMNjkMeOWsvLI+Wv
u5YCtwDomrhnxq3PqhCNN259WVbCRNc4BaQSOqf7rhU1JiAbsD5ReUCT/EYROGai
Ona0OXishwM9X4CvWQdgQDTA3E1EkeECIigV0lReF0U0fOFLcibXnqx+OC8i+YwT
7D9ZbJ9zgL1bVnrDscER8DMp6X4X/mvzltxGTDE5BCz56NvxNgBeIf8XzB6axWRK
JZLmF0bu7VkjKCBleM8XthhTyMC4S67hVyrBw5nGgwRdu3CRYPv0aIWeH6sUBcpp
byNwaqwp+lsK2KiLVEJnsIN3T+aWAeVY/7/4wdmTDl4YfBTY8b0xhlCKeLjh08MH
gJd2z2tVOS+HTzhxE0HWPb6Wo1Xn8WVHjXxOubymGcbtE8t2getfMWtfr2gs75wu
GynDBl9YA53U3cAMWisSw94WbfVStaDhEK0EiPYDof9G/FrjX7c9Sw2FBDwDEJVn
xhgzw+H/obPwSWLyi83MWdQrr86xQ5qd2gLM+BD+RDMdWHYLU1wDkaB+T0ZZ22y+
romdbiCIdYACVRamub5g+3qxERywTq8b7EWAmwgPQZT1MRQh+FOcIyfMldastW8K
LOCw0zqGwgHDLyxX6PqO6F437KZSjitITIxyOMiPfZEJSx1D+INy4El7Pmc8OEaR
9/UlsvOdyxUxMILNoiVqqUup8arm7ESypMRF7fx6MljQwzLYVLtnOzYybKZOhQAp
V3TJF8i5eGfRjitJ995DLZ+MR2YPsW5ZHDFeGZlGqIO4AF0NjeThRA1s9PEpWv0y
obFbtG3p3QgQfE9AQL10NOLsxIIUHagxptUmnxJId0v/YhiQ0+J0re5DewuTDa6B
tLrlncpK3BYSjo7LWaVJJJ4gsCAyGQeMX4KHPk0lpnqn5aekgghfP8pNe6IQcqcJ
AfZn+Ugv2IQH8nGCOdPyA85tWqatbAPsU75OduQWAoSUnoAZHcCgwRUT7Ly1QirR
NKl+FMtmohGxShKxZYoWPw0+0AQvhhIjUYN9Wva3u1NK0Gm99VSC/EKKlIocM3vj
n8Fl/BNkV/11LkbFgnktxk2yf9RtFYftjRfDOugJWwiEBHl4VkqY2moEZSwdg6Jz
V5HJn3UatVCX0B35dgwtuGRSAQpKwUb2u588YPx4omAXe5OOIhAfW7nF1mY4tMf1
Ne8zwCrfLYt25H+e1wydtij5uJ6XsmI56FlpuXOFc/peurZWHiY0bn+mwisE9ft6
/7HRvxRJ+cOUEmrMQ6I0vGzLT8NKC3oj+itImHsvk95Xg/oGs8wfjhUYGEihz/+o
+AWE0OajHlsZSJrgwUwGmR+M3uKzb0+ihYciZAe193/fdbl1AVBJGn3K3Dj0LFHi
uczt7ZNhk/d3rGLgcIDe+V1zrNg1Yy3UJH2gilCIiaan5qWxr4ZX9cnyyA2QMP1T
r3QXWV1smUGWTTFaCO6b8FxsCgx5Eaap6/tgMV60T5lmpoVPd4w7Mqi2ipUORtKp
jHZatXtuCxcafj+V66jhUNoc8SlK0jdjuFXNhYURJgarGdpyy9PtnvNsuoq42wFT
l3nUqACPREF4ezIwn7U1lZ8/Qyb+9ZmLLzehKIemFQIr11jLrtSJenyBXOCsLicr
RKAMvIPrUYDzlNtcHwP6Lo6iDDq6HfumfsSFaRYrCdBxcZSY4GWGXmqtIefUBA6J
mnxs7H6J464MvCvcl4p4kcs00Lwc1nj49yhjog2ya1MESwiMQUjDX1RCS2HZUPGw
Iq5bqTHwj1RJIa2yY5HcqMQV4uxa8zvjf9L9Dj23ynT8vySHlkFGdHlwrU3xRIZ9
XqkpmeDn9Yrirvig9hhQlXVTvEWkqghwlr6wAMOhLUqulznJw29uAd2pGXiGzOgY
hSpSUp6OXQbxdinJkoKIEuH5nNh/vVTxM/cySkpZadzpgtxzbIP1IyOe/YRd/JAa
klJcU5DWlD2KdQbCicMBu4uaHklo6mlacz7124AmF1KrnVXtD6O/69dhCrXnjZUk
Pw4H58sCxVOtx9k2HCviq6/NCWI0/7yEKE4CDrQDY/6ZHMY7FgT8UZKVoNx6ub5Z
883jyYcd6HlrNR6KjeNt/p0MrCy1ClB0Lsxop6sAN1VBp22U6rSgc3qzR5uDBkNb
eQ8AeS8mtbzP/TmLbfQEU5clyciL0joTgD53Hc3jvEbx+3C0yhYubESWrzGE2cCg
Tyr3NETs/DgdVAi5vh4XXy3xsjyC/35c2Uusvfoy4R6PNLZAGGmcD9Mqpr26/nPB
R0t6FGI+O4Fm5AyvzAvMpdO0BS+ssyVsvUslqDRuBt3QRPt9F0e2d42gOpuhb8jr
xYeHaZdrWKe7bdAF3GcYl6dIl0hfSg3u8YdgKoR+PCrmYl6/Lok5AoKl7hhcnPn/
KqtQ4T60xROX1/5tt49AWCkZqAWVBSEOXqz08eeGa3b26+GpAkZ9XoVYRP/bE61y
QmTOXzP5wFyeqf7VzBmghkEE+qW2KqEm3Pr/+U49r/l8ZzADXcYZOwGBz3C8SlIZ
ZIERlyYmAHfGh6ou5PxwM8L+nZiXm5f4jIhvsxnq1nbdUvRBSYA3XQLgW6JjMk5a
Iunflp5huu40Oyhg0llTNYNff1MtDv0zaZFBuBw6BBuT4Z196lbKFE0o8Nfgcqkh
baKzWorfFmStBRhJ+0iV15nOslZ22TkdaYVu38LEsThF2ZhaySo+CGDzgcK0vuwM
V8k0zkuio5md1E7+DAzKmJDwQFwpt6ve/NiHU+UOI99gwzwuD511bzU/l826rY5x
8tqlDrygqhdYUFrVZ4o+x3FkncYrfkzcd4e8YQ2Dx3Tuv85dHbzLvgHjlXw+Vcni
JO8aTalWZMmw0CYYLOHsbB3LA8/HcDdb136dSu5dG/HRCKI2r++8DunWMHokZClo
vho21yE3C/A7fQt0aslAFQu4oSpM+S75xGKCRBRNBLDX82Phs7odz0t8JcyJ024L
fasrlV+FeQoCYVPJxbeA+o4z4LxxC38hJZhjM+U23Xwo3v6KUT5i4VJmKF+juxrt
GQin3qoUCYCTV6FuvzKKW7nDs2ufbvp73/aRv9TelVf6YBKyABXwLr/YbqSNzfY7
WMqAqMIDqxKgrv69UHCTw4iCajGPrU6sDXZG6WXJpaCkidLSNZqCB1x+Jg7oQ/Gr
dfUTTFc+VinmE+RsHd3EPRdTX+SOQ0yiaaYYMfnZJ0Riir4tgW97pSB6dQvhyugY
+miMbQ8GbESVzr8cfpULyxZ77ftwyUPXXNEeHt/tsxV8dFyFCciRCAMkU9Z2SjJn
BhgUuL/RDiw7/7DgEGbvwbNP7+Y9ZyWZTf5fyflOBRpkMQ/9bGeeYI7wcn5LQOAQ
+QT8UPGC7PONa8lPwuLQh1XVy81UvdNn7kZSp3Md0yvV8ySmoVUIc1Vf+yGDtnK7
YqADyeEwRHPeNReWduukX44ivcFSPQkVwxMUjRpfcMJ8ZXCConxie0P03wlDaVWD
UhNeL1iCXLSm9oj0cbGGBoBPH3Uab5QUy/EQlnhf262uecUUEIqudNj0LR6OdsCo
dhUIxuy1tTwvnh6LKahXmSrFpEZduFAOpHR/iZpvtDT6I/kwX9gLuMQyRG+p+8O9
4eGQDQAnhXKITuVp9ALG2Lb/RQKO7esfJ2dCD8g2SBssrFg1VmXusRe/lbrQsVii
/XB4LN4DwfcVOOYIdZcuPoLZ7Dxq7yu147FKseJ5QsGq+D4h8sWeWx8eXPn44IuS
qdehJIL46SVxdp3ZwCWk66ww/WjViQfPRvUqcvMw+Hd/guhrosaRN2MUjkSJUu37
NAH90lq46M/wRT0eqLHJ5S5osK4ESXP03LnfbLOecYLwW/SmHwbYPV6yfA/6Cmdf
0hLCqUsiW8kaFK8+GYASrxbYHe2VXf/DlKYfo/aYyZEpnPPXRkqZNBo00f4mt0oc
wslBfJH5JdXTmgDhQEZNRoi7k/8yKaZkQSxncYsZwh5nYPxqXaUvzNbkZUIvPNOp
2sUIb0RB7bwAHmZ6gmuZY2ei7KYigvnLMbLxrz59MZt7iA4bGVo71DMX6RxRpY6U
6Kr0rDcFMboF6KMTpiMHSEh9ufE/l73od603yHrsba8qIFiVXZE/uf6PQXi9GWFT
dZWW2zG44lwYnmX+h7HDZuMKpGRS5J9TZRKQkoy1ExzcmJyr2Y3zXu1WofFi30CW
McRqUh1XTSUX3YEp18j4oTz3KB+e09/m+dZ4oaOJtgXibgLBcJt93uuQ7mziXSNV
2IO8M6DWpEA9noy45MtGt7foe1MgVXn4y7Ii4ma4EZOGcyifZk1Eb0ZEP/A2t0Kc
jOi3S85Q98t+ErUtCCvzArONleOV+8dE7RkicOqkYwgYIWPDMjsfN8UjG6l5zRus
C9zd5WXQq1fyIemB2v2iOv8RK2nC3kQ/+ZQtH2vNH/2Jwh8ngiJh36S/qOO+nTUV
aUqQaBOQ+NjXxo51VS3ZsSwRAG4lZuRGBNXpr4CuaOHtQLjGl5WgoFdBh2ld17ku
14ycj/dtF+ppdjfdA4U33OfIz61+7u49zR+fYVn7/dHNw/1Fqk8k+R6FVz/9NvI3
x7kwSa48PvNttYjt+VhueTPRCloyOx1cAjRXmURRcPf6gOacmDDYLdHiuL6HPt7v
WRfhpnt6+gK6RP97eQXn8xc9rN6hP0/llRbh1+phOMYHAsW8bgR/77DdDELkorJC
u2cqa5e70ABWXSwFwbV3L40CXCfbe9VcPBTsSS08g3Vdo/oxPOvgn5QH6Ua/Doxv
4aTzH0ZUQJ4RvPEWC8p3axZnUx49/cqgxXr9VbmY5ZJYCBnL9Ftz8ZFyV1Wp9QW5
JeGc54J4jHw5BUaNtlM/yAOGq/gG2k1gT5B2JknEjFuv8ck79VpukYICr2/GlLiV
FUDIvlXppY5tHPE2PsFfzflyQT5ka2b0RIaB4fhFsojvRxHFZVT1MuNaTeAkPdWT
Vsghoqj2CJ/JFO71bsJIducbWBJsWuVfa+4SMJzLheHNTF+qR21Um3/1mhkKCamw
w811I9DNlKDFJkF7+ZEhS92w04ZjJVCeCWwQPVEN2I7BSo9Y81+EtDPzzJGrcTqb
tUISwz/SeKRHN9AEJcZ8bpggK6SfDjrFTDis1KZI3UOMNBqyE8eOJoJbgUKraiWh
Pgjw3wV+p5Mjk+IU7qrTWBccBzhPrtNeNIYfQaiVotw8/Cdv8EM7PeuO/F0Exg/e
sR5YLh+sl4J18zldTqe1VqdJ2UVxB1H9XfsJhXTroEpN4GPxw/HNx40qLN+a9bHq
zAwsbJ0Nf0OmI5GCgwX4pu9F0r+GOTIvyVESdAjI8lL1xbsZe7h+vP+5p4ofYh5g
dN7zsz1ML65Y+XP+VmTA1gaW2i5lPeCpbBrEVowdmzSSxFfEx9UCt/pj7nTw/pRV
ihX0s863GmEfby0lA75q6VnF7DIv9eJx4aKyQ0p6a53ekA0UnfDv2G1PmkdL+3ns
lHVeEwnT8bKqE9v2+xOgWEUWAmINvXgSzV297hOiOPJmmv0tW0hFwrS/5IfEN2WA
nP42Qyu8WKtvuLocw6yqFdZlUsc56OqJ4E8eNSlP8XY3dJlNq7LOmZuvPI5MD+w0
ZJ4ImvdTEaCiGIEyUBYpL261TgNZrPev6q+/XfARt5mRU+S4QEqxF8ogx28hHJ6G
XAphrWxgTuWWO6nRE/B5enPio/8iu/pV8YMPNpqNfS4WCYNA3KTCnP6Saa1tApFJ
udGLoUdCZdnTM7IMpDO1xCoPHpR9QoWHxU42ReGXQCPKKaNiBBhCzZkXcsI1HfS+
mOU8vOi/JpUvAuCfcQeB+KDxTTQSqBmSxpnQkRmP5j62ClzfVIl11ZL0/KRIPPli
iB+JMqu07LgFI2x42WT481ol2prDwqekzkZLThFNXNhl1YNCR+vIPcCvMAU2vPhX
5P/96F0ggVa0kcF1ZB2L19sSZbi1DUYwKfT1nWTsE47x9wpqJTUzAc/6p5lLfYcA
tJtLDIwtuVh0ER3cDIYrW4w3ZNGbwVnqhrLpbkWTh1hai4wCm3SdL8Cu3J9qW0cs
jSjc8HBzylCqJROh8+8J7Zt0nIIY6aCSsScKIrk1tqTDzxsPWIzuPIezD9X4vR6s
q7hDSgXwxBlyw19IvoV5jkOWFZtx+NHi7Ufkt+GT2+Y664bWvcE437zbOTWQjTWq
vAS/JMzxGSXCyHF9pNLmKrn/Io27VnDe++gRig3xcqh5ybeAe6L9e1Y0l/m/mPyz
a5uxVYEyJLzRFKknKLQHs12jzn2sotjPUNqmpn77beWDvG6i3dnJyoJdGKd7Impt
L9gj1HjgJSZE95+X7uLeGB8LFntO/O6n/Mf7LI4LLbBGZf/lkbfKDZQSWSI5hXes
gEi10aCTw63TvHsz1w9wEylz8jWR1zjWt5EcggJE3ZDJu4Qxf2q/E915/MTZBGVU
rhx6DoWnD4QIUALdGW3XoC0lFY0Wo+CF8+grxS+BRrPS+CxPvQNMpPhvWxL8BRGA
hoPZqppQRvEIzLvM0JpbqHXBrOBwrM6cDebsG3YY9ksfBZyPJBIm+zSIfgkoIFtW
90ruNMCyL8bhr0NXEhEUIIR8zU1Def/8qhaDLqgFQjKRErfm4jc5GOHBh72Z0t4g
Y3kY1hinDlXn2IIMp3H1XaoBOxA7My0Z7yKG/hbYNEFBsucgwyvTGmwz9YqTZy+2
JH1aGlAvAE2tLg6H5eoMg/XrvEb7MtKmYG9v1lY0VF6t7tEgrs9LmoBP9iYG08YZ
4H9Z/foQOS9aXdDE+yETcsIWm1Emh7Yq8t+Kevfp6jsc6+nv/W1S6IolaJ/pfb1K
3lfmjQV7AlMKlTUd+29AbsCtFO8DzVe1p1KNdt5ZbPnswcy1qyGMkPHc+9TrqqfX
rPVq3v5V805Wu6wUJTStDzLT5yqz+CwYB/krCh/HsomMMPsGOOi0/g5NC2yp+ldK
8IGFP/G3ALtGQuQisadw1ozVDoIR8eww6M6qnVgX7DhOPML7FJf0sWAA4DtoIKCp
YNqGWj4Gi7Dsce3R0G01o4k91zEzn8FJaPqczDVrw0S4pJiRckfTw9Ox2QrNRtdj
GFhfdPdI0hvy9kNp0CY8GUzJCd1aQxPyD4ktnc70zLjl9bgCgyvsR4dwnGv47xkK
ZH3rRn+frLazE+ik4j/dQqNKBNeXPh9/hPK32j/8s+MYItke+zH+g3nZtGAji2rS
1FyyWUDgzgqM6Afe507G0WOlplZtNdldIdk6LLG88KuhOVf/n4Y1cxMEFgYDKY0L
HjuERS+h19vBC+l5XpEHZLyk7i+23FW8pVv88R5eQ41TrEwHNtjz0m2SZiHCIZEM
nCyNGZpXsKckgYuBLdkvttkgVe0SQw5cxFc7LXwY4u72d6bB0SsU3wpXr7cDNfC3
e8UAb53+UpnC0S0sfG3/0ILoRLL3cF7Ri+lXjXxgUipy3prSUqYKwjT6dyLEu/D9
x8FfmatrTExFenrRHgAvKREbt1i9391lc8oflEjzFt0m2nkiWPpuIdbH4izK/Asz
Usv3Acvkw1YikyysNvL3C0yZiPq38ys78nodKuOFuFn9046FvKPdP++dJfnylXzG
FhcEGbDYCEUTTeSnYJ0ExEBgR5KKsPrYLceVHEOXbV7WE8So+B/us+yTQ1Wi89z/
qRD51IbFEG8yNrsKHxJHSAQJuOdF7lTEMsb0XbbJtQY0H+UIXrnLOak30Rtma+/Z
EBKzb9l4DAJty99QbAS4tlqTq5CehlCVGVhRQsQ0xCP9CWve4Gj1IKpwkCGzziAD
1WNhxYM5HZdJxZbVHUdgTnjMoXfKobGAS5Qkn/Vn1i5fjUD2RW0bV/8/dCx3vdsm
sANO+RJPQQFQTafy3HeVeHo1tXzftyeNQUG3CojpyknuLeL5uqlJPMMaxWxISAyd
C1Z5D5P45Ar/4BiRs1yiTn+Z/gkDWqORHobuQzNHzfwrkXVyqpSIMNpN6nBSacMH
bEXRWnCzjUQ1F7seeq+IwhEjiMPsS66L2D+HaUqNbOqBO3a7gB5iBzfbxsARTnys
3qExgR/87QFSBKo7P5HmSkmSC4yHeV8xqf8kbEbZ8zLsW+iLobqho8HgpHE8VE/I
kzofmbVp7uo9cyp7nF5xDQ1yjUWqnw1MGhdSwd2xG7iF9SzhjQvuipQrw7Tf4/64
dobKGeHkSTW7Kj6yEp/UOjVLH3RtQSJATP5YHhGw3v6WE4hI3WSnb8tm2a9tMIkw
XpVcETKmCXDoiNSWgN6Z6kFY3kfbQxD19dMkLrALnY6WUDgCsZH35XnZm+3q+Seq
jUJWe9oOrXzEIGXm5VMMZnLJpwJdonL2Cfp7bFTt5iPGMZ1wstmlpMk5o3cMyTZs
bcf1DT67Ka6Tz7fKObMbf2Hy8OXFrmPcCRGe9kWOdwDRzBVyL7XUiHWpWYfQV98T
8aN+ZhQntrX7z6XZSappA33pzRIBPV3+sFSIQh6rKx/bFQbzyYHan+WCZIqxCuFY
/eoHjh2x6Erj85uGmc7Y3GhXuJV9tiXhxujwxF3dvtMgGBksITUgfo805YVt6tvn
K1UgfPmxCPxbBRBRpkOnEc8lcNdhDgdMzrGwjE6lWl+P2MlPpZxOPj90nYf202O2
jzaOSx4OwOXsleth3ZS6s/hDN3K4pqT/T8vSa4sE9KDaz/DAGMnElkLZDxDqOrB9
/SF7gHATwVjhWoDm8JyaZPbD88v1Ij5UcX/DarqTNnLNH5X18+5KzlsP27aUC+RX
6vfwkssfVpf8PxtXEIa9GL93+M7g8pv9cg9uPVyXNu1q+U7AEkzJrh7f9M/ZFENR
kL03opbCR4MeryykmGaBS5OkEvJ/GlOu2eOxrXXdJFSBaFmvwT5hiSubllEUmcGJ
VL6+jJYTKl4gj6Ijh0/cd+qGgmxJCCStKutrS28rJeivNxQsvc99RS/TC12XSSPB
7m/KeDj7TL+4cBgbPA/le+aCP2v5pGEahSQXs9khjXYpg+v58cBr4ozmZkZMvnl7
m1VuinF8WXO0xBfbcoKPA2W3Bxk/DJoWWfB+3C1zboeovddLjCImt76NXgPOyf/E
8kI4qEvB+Qmm03NTxsoLfr7m7IVDhozDs7lWykejjN+Cf1J88U73T1k/lmX+uAor
VIzJU5LZajng3+TzvpPPVrojz9k/0OvRf5GgzDRxBiUbQ9+ywPZttKkOKpvmNdU0
hVXTrAYb9NZNHWBHj3RDT9/cWgFbQtK+rftWbSJWlkDqmT5j/Nmo2GXjJT7ivaBH
6apJ1zDqqIODFf5eQjT9xRkLK3Ngkq/6mcr4ffuvoy1TlPC75wr/H9I6vNP2HOip
e+Snp6LtYPaB1S9ING/MVzgokH/6MyYJD/emBQbCd0GHTxNGL/T4UcyvVGCS60uK
dlpQC8/USZnLn7jPKwyLgE8UL9/lvBHwKbpZuPXQ8QeKeI+Hg8pmKp1v8XChFuvD
iO0xZjrWodgqWNdQi2NVvVNH5dM5PQCSh26yMp/hEqu1x7IgH8yEa8Dhn3aEzHUi
QTZxC0N0mnKT20VfpJJPQvkHggqASp03Fvh9ut9hxsxQ8FYyKsHaVVklQjBMH5ky
sO73aDOCQCa0CsDK7IIl5FjZ6lw1EtDWai2QgU8Dv0b68yheG14rKl+2lSZT98jS
I/0ibRIkF6094TRkpwscFfNkJj9rHiUlAZLmgngtmZiMHi59AigAkkgi9O4LKf0C
qGmF1uWBtui9bhJCS3SecSx89D7GkMWisTTutE6ZpzU9caAR9oxJxL8lQ0VyvDdG
wi5HjLxscx+lMBfnnpzcU6MamDssre67oqfpMV+pcoLjKXRUcuj8zDsOm41qYKXQ
74R2/yl+WBlf8Vtko5Jf7UQeux5/bcXks2tLFH6z577yY7JVj3JEpnQxmUYYxZYC
CZmQxE82GAx8huMcO/cFropyxAdWjJUKyZXr/WgTtPJWDW/RWs927dRpEfZJZu5E
V5SaA3Z+U2eiCk1kQWSLu18d/eeqrSmp+qcPPPzbi7wq6kLJGyqCA4mWbYmHnu2m
wlp2JhFDu5pxhDhUNdxh8PwSxQJvKZmAic5kgf+SVN63Nk0TaYA2w/5ya7ZUkPME
GjyyjxGqTH0gXyw5gXrrB4e9W6vkz1QQmrCvbom/iQ/R3aMgGv7MOlhtXvDztTHl
51QlNBXlRkmA3F2W05XJuUSL9EqxyH8xqHOxiJj7TQW9JBHr3LqXPClxF1zfI4LY
Vr7QMMsKMNSiHMuvN+3+Y9BFZHwe3JgfSIo/eDLID7ayJKChKId7BLeut06nhT1f
dPpfwgi65YwVYtQetHy49o+dawpDogzlnwn4PnhYQD6WgF1cPn/pZ/+2PtHEqPki
Zmp1enf29WNbtZrJGMkvL1OqbBvLbhTyz9f45KByViBw+btClHgXOrebzWFt56EF
H6GH/kT+bk4wgYTOU/oVjhk0e+w/RVy6RYR5xlCsJ1rG8S1gRVwF2ufg+qKj7fvb
4w0iHh0Z8QIgIB9zCpuEYvXg9qC3uXsOWgKxolP58e837EeEXoPfq+P2qRjrFgoL
clCZ/SoaY9Ttd7Q/fUoxIscUCeAoTHUh5cGerYtpqJbItZn3wpVUGRro8HbRntNS
d+9MDIZp7ALAqsSPuuV9un+lHQ4TDPIStuWt+9tpGN7ZyCwdfYdLz1yvnbu2HtlS
yhZDNUPWduVZwiq8qzGV9PvK/nvBJlP76AYza3IyAKeGWyC4OfRqwRuVKK0gW4k7
VllBn/U6xL7uzRK1yMU0WKHa059mCYLAusez243u0cYYWF7kb+AegrUWVwpONsgX
SOfRdVbbmL54vD+R9u4Rmb+1JsALXk5jUiu6Qo0dLg1GDE4b4+RtRA4PUrE+fXZX
y79cumVfHloJfFmgXLtyhw67iHLsZjWcDGYSSqBQHlruVVj+w6c7U3Kq+BdOLGIu
GUhbuKsP/1PU2w11eWC9z0C0HeQ3T9oKtr2Ax4ltIujOiPNPJkVrp4X0xGcRVWuf
HhYECT8s242nfD2n9qjb2NNptlCIdi5JRcwUyxH/KacLakrkL4EFg7ALD/ubngu0
rLnQCf+EX70mPwyL6hvPSqEWDEX67g0nCqFXc1pNxWxIRsxGuNfpVF2S5dca7ZUf
omEtHqt6bIX7X+ntrTq1+iSVOnhmL3W1mftjKwkGq9xIpTyT1J7zJJViYpCX91cQ
AGJS2lpSPRxx4c/Cphr8Mv3cVgnugXye/UqDCDfyX4Cn5oTv7LWuUp7QUX6679dX
lYFxd2v4zXr8FPLPkE9FnAaV4AdbLdgbvFVApBmHRRASYku0vZKSHBkMSYMVFaxq
Nr+M7d45g1DaT8kO0exmQE9fhs+No1ReszeVT+s9s+rK9NFJQc7D1awFe30HOpzt
uvMU4yyfgE0871c0hL8cpmnYtoz2YQWDhsGYh5W+395NcQDiSLNeTPHcx6fViEaR
v7ItpEA0Hns40CZPkFPhRo0aAvqYZ/HjFy10XTA6s6Ansxo9Xy0T5CjB1bLv2ZPV
vkkVRWGFc1V8gFzyjJgbHfai12hpDO4s4EOFrIlyS7U9VO3VwqM1WSK0mXoSuio0
q+6R6V0P5xrfukuTdPXrQ/q5opMcYHpJfhrR5gtxZRKZR1p9wEJNybN3oLUHhtEb
sKvuTCNR5b7oFFiCQmkBLlfy4JkY/bCPNQsVIWmS/yv9hz+zpawA9NqwzL3+Ty8N
CU25g1JLL3gn3eP3GWNX/EoWy8HHhJ/IwBqfRS050AOcqV9nXbenrcbqKAGQ+k+f
dXz416YZDYabIY6aIOLHUUr5ItWSDnIdn8AM0tdzHL1CP5AepgDuyEke1bh4H87y
R3rEo77kECeepaT52Zon6M6pnKUJFVbqoDJOZ2BxUsiuRD8T+9hKTZn8nXZ5/HId
iV7tMMpXOgOMb4197OYE+L/faS2IO5qTcO3voc1PBMEesJeQqUdLBtvueJKgOF5P
V4v40R7+Iis9WcCWGD0UBA+QHfG2iuv42xGsbKaErAwYJTQQKwPXENwq7K857MWO
j2ohKX9KIgnhuUzNI6kGvn5JQaMQc76ezY7XSHlYcUlH/WHrD0TO0jLJHTfTnpBG
7m3rfgVWlh7/jd/TBSKachZOotbta4Xj4zbXCytOhcuvUaQSf3bsaOwZHvrYjn3F
LwPQignzeFfhaiX4d8DVrfi20AoXKuTgugvMu/BX6S87oBDFjuovbtD5C5S1vEaH
1kf66rdUrG+S/4NVOl9alYgcZRuEtI6BVJ9/AtRhXPkhfkcl/4SKttgBOHAm/per
wl/Pge+ktsbpw0ajHQuZJcXBs/tRzC8e8g0LxIgNJHqijTa2HcA1dqYxM1Eq5Q8H
wleh6bIvVevREBgQYihFq405j7aMDxvp8/f5JUILET1DmiVi6NWN69PxyW8ZLEGh
b+qr0pstFQNqO1EwxGokEPhm6fhEc5ixd/mz3O2SL4DwSACU+dPlw94BhowfyW63
FI0HAAqQ5mnqj5SHBbF7+X0S+ATPYTsBCmLyx7hRxB5DsKMeaolU0IxSNHxqSA3q
7FsowQw9E56xWFMmFJzzsPPgOTMpMYB9ce7MU72OY9JzYzLW957hVy4eqHgrg2GR
eJCgI3fAbQUD2b4v6awJU8Iu3sGEVNI+Kqgw/nb4Pw5cUJRbUtXoS6O6EPTrUnAa
Sb8GIDj3WRfHIOYsDWk/b606HCzKqc9/4N7qEdJ3rkVtDdCBglaMHdqCeymVHmNp
Di0qc98GjLHyoR8tBYG8n3G10c0rmh6CturZcEXSa+/R90YmvSbXNvoKfde1nHfq
ouQLjnRWZp1Kyud2iVd4+bueSuoAKGoeJQFW0k3w5+MnUImaxiGqMVaqQIobRwiM
S+uPh774BP5M7c1x8+u5w6VwC+7VXdEl9SYmOH4DU8Uc8szL8XzOCJhONshPJBs7
TfEZkvtlRkcOTfbgs0ashW0Tq4q7SHwMb8gUeHoxgSrxzx1TdaVYMWB9tFD43YBO
YsYbdy+es+tlTiknhCGn4OhMUZxKAX1Au8McMS350+1nhRY/EpkZmFC48nSOeFWO
60QvxC54NrOJxbDDmRb459nUdjwUt58fpNmQhAhS/KCyF8xnrp0ULC20XDjKmJYQ
a6azZrh+qa2rtyLXkjXmPNcKgM7aJa1x7fZqQZHTu6NuqaDjloFIeqlgiaSrXPxm
b6+lM6xseEuDQ+iPWdzsB0hM5ATiGEQrYYEzOhPiucc/R8uM/smtilqPpw+c767r
HzZ/4ZEFk1qDLJ8apfZddLYZ//GEFzs6Yv9CJYGX+rY8U30MeeuOskH5HMC1nNPu
V2NAC1UABILtXVmwh9W5Rrj9J6dG0inIPhKUJaeWbxgmQ9CoE6a21CDQJQLCvMxC
GKsuS8Yk0ykybm25VK0o7PHGsng5bUPhK46q5RrZt7LVBOvDBYvHo9dsAihMF9Qf
CmuoU/BS3trfqLXp2FDTQafrogdUkGp70+8civZLGz4OoWikPOpuDABmHUxAC5xY
kt++MtralsEdIdlOnuAU3sE0wKmVPFtjgdqgMKhjo8iMJmmZkHYBGV2middB4uzx
Zg7jOWMG+v8go8oEQVP+ldiLqamHkGlzYplKGjcrctrV82Ppx35kAAZYqtPNi8rX
hzJr6hFPI/otwn4/2zYmFUA0ygp4Y92atgJlQxb0dnwb9ETQPR2fcBh8+5OCTsFk
sJOYgmgCKPHOJHEAAJvv+Enu0Xddo3kKB/piQlpuSAOi6LPVG49Ga27MW0VfVbNU
cpS4iGu0ElldpmeY1K863LycyHgbgyECWpUc/1Wn6JDCQzC9E8t2Cd9XOF0FD+z5
lfl1WfDarvXL1rxC+IT7VSuHHONqxlQ+q74f3B22LAI9ctABgcdgtBWrzyIQzqn3
pxJN2u9AZvgu/ZdCMLLNM5c7mm5OlYDdZq+WtcL+aB5OwmVwZ5JpJT3tuWDPjXOh
3F1pLbM3lNQTSQe5GZ+5rEDIYQK6FnxulXI+SSTTUB1BrDIbMUZd0zW7wagjUxqd
V/3uVNpIUgSLt78WzV3ZCoqDjSB0qla6aXCXkFbew7TBXF12WtTZa9bPYEBco88V
EPg+YXXfx6N2jiqB8ycWQlhRsUkPjV//PE5EWmGfMlERSz/7FTb1kMXxKlemCV54
/myqVSZduXBr+VU938BHk3RoqbT6N1GDWJb8gVUP7WqFsOeUP6lCnI4zOKPihBSp
Ry3wt/SImafs4i+5n1gYaH72zREX+qDO72RvDk5Qi2YiRTSxBbolAycTecwbBOBy
KlpGaVHR36uuXpkEQdeoEyNrqzQG1dIaLwl5SRAHWXHwPiKFoKj0n7WO//3Krhlh
yAKOPDbDaiQW1hV2hvIfQedoWbq9gE++QVBasgB5vUdg9nUztxxwcX3JSz5mSxd/
B6oI1Zc5/JjPPuvehcH4JtRFZFS+fFMLlG6m8iG0NYsnxX149++HoBfmzU/rf5S+
4Leb73PvJh6oRRHihFbGMYZWVdErAzaYfgqhP1WyZtvAYEqowyvuNFJL60piVf0f
6bpVoxextD2IN8Paa0BhQGyh2K1j3ZT9Dt2u1DX2Ux5aTKiGsxmXYuyqXZbOuc0y
3PlEFLVhGRZfpEaPp2d90oWybKVNO5w3WBy1Hvu7zwNGzWbUuF2cFZi6mwa3lhGR
tGGqH9D43WwX9b7svgG8RcHNxCclcsheRMI7y3rM/ZEz3OT5wHm1ShSK4pAwdG7Z
ZzIgn3CgLXgtcUuWy2FXDlogX1KUG1Qjpmf3i9iLFhl1AxXzC30sfIt0f37fl73Z
AMIlRzjuQW9h0vJeMmo9JSb/VrBirvGuIARRZmcP+lfvT+87I5fQ74KgmNzwvwxs
Zo1PhWa+fJpMHiHlvTsvCH1rvb9sS9zfiUy9wM9f9R3Mqh8Jmm3p/eIWt2AAGIEn
QHkqD+MOX8NrQ8L49F7EqjoFizeC31cOlfeF2v3zy+YefDXI9SdpGVewO/wWkDlM
DhBFH75UnHBCUyZS4YjlE1mGP87lh6b0LrszMEcJeI9ghhMum6+HdNr3imldzpPd
bczJcfEuY2xTnGATPhrz96sJ4R4CJOLdmRDjkrY29WyIh6CVWL05PEZh6C9AT3Bp
YcMWrTgUROyaNfjD5pGVSEdP77KLrGSiDZDZj+IHQfChWFC9dzpF1CFjpRkBf30z
pFczChxOrUvbYQ6jTbNsgFk7DF10sljYZ6H2KxMogWPGIe0oQ+XaA9zFsud7/gec
YDvczYlQQrx+JIhvM+2uDX/bL9l0iFdsH4W8O14HRSqDkJw3Uxm/TrqXPGc4BEyM
SsxSh3HL124ZH1QoDqPH0iDvWNgqc71tujhI/1V7BMSofykx32Iztz9S9LU4FtDD
i/jDNsI10kTYL8N+OlhZmrwt9cXbI5boVCkOR7MZ3tQI17d3ZNU0BlJf/0m03fC2
kjGyxYNfO0i1NekGCO6/LDWyjVUSfmtka4rJ4lGoL6DCR3GHcOr4P/yjjm929ycV
oapvELn6nKycPFd0KzeKWq8ONuaZAu/bFso+msQCONKG/90GoHzcBk30go4uh9UV
B4rfK1iDnE+G1Ex4jyXy7L0Z3rjCm1Bu79r6wSHXW6eZq5kus2SH9BICnYlCI7JJ
WoXk2/DwCYAoUomZgDgo4YwJivDGKdUnmS7/ip5hZEF57f8s6epPmUZwPuuLqk00
hFahpkTaHl5SqcnCV1hUD54rkAu931y2WOXibyUaN226zMAj0dR95aHflTukBv5x
ZVvCwn/bHxHVxlqxOiIXq5HeVAy/KXYkJR9j2gjK0cbbzuWpD11MdSS/Zpz1+Ld7
KrvEoR+RHcjhhyotIJWiWWOPxz9i6gem+ZBFyFw/kbBm0I29iBB27UHYel4f/SMA
hvXSMLojA8pyPt1URrzRABe0Gka+ooeI89mXZPCiB91UnHgQmdTEMsNzqTkd3znK
3EEFaMPCCMeWrkfZKGIuaTrCDGTWjTeBxYkoenD1Wojz9iaVf4sEeOVRtjvVgDZI
gtE//04bCn8RF7045odvbZ0m3OPFnAjqZhKfcr+9Rr2X07C5PoKrujrPG1/OZ6WV
WsnCk1UJHo8rIwZJLHQeM6YxUDZLX7UnzXaj2BVlyTPJQgZVPlkBOi1V/JDs4qJ6
Hn+IHQsWw2UqrKtpdzRQal9WRnRhlsg2Dmtq0GRuHJ/frvZG1YEWraOrjNHDV/NM
1Auqzr/3ZMBuinfpZZNXtjArebRrFdO73MvgeG+uSyK8HXb9HoaZVcdYqnInnDs0
OCflzVZDeoxw49oh4H3Skm2VWCu+m6AurGueidw3OSIAWuU377QDp8cD5XNrQ/fL
oVIE9oy8nKaYSX3yjfAxqQL9/0bzu8lSlimzOHI6vB2HJVcBz5tVCj6/ft8pCpte
hnXEwHPfGXq+a6kvdiDZDYPJsYY0DKlmr/kgI2v8AwCOYviArgX6N3/U91/JZEa+
AS7LyWBf/dYlHeZEnXUm4FwpvBRinbrVplwAzkQzXTbqmq5GtAxcx28jxBrxpZvP
b8cYqRaz7+57fioa1pmbWg6rE+jJgBTrye17mvTh/e3DFmSpBTRk0rmuThiCE+I3
QraOXhMyv4xeM3v1f0Ye06+M216qK4QAGqAg3sGXijiFlILN3sS5D4xSOrgh+kiA
TktV2fXVxPHJSYv0/0GBs4R16RCCVXTRzH0pwVcxhGgUImw1bQHs0935RxDG9Jih
ECPNDaW6kD/NnCiOPNRd0K2q3YXnq4NEiRrf63lnyD3QgxI4GR8M9Tie0+YX4Gnf
kvW5KIPbEFuhJcwjmLQuqr4JiXktC5qphHnMej3ry7mUWfTOLCLKmc9o8DHF0Yvc
MKdre16K/eDKvZW+cyoEuTGbIx3In8D7lAeo05td1SepL1VnJpjsTltjBkHWudOT
xwxu86f+fS+WCwSRuPqVMSuG3+dU3XApRdsiw3uin8Dh4bPijlQ+ynvJBTZ53cDK
nICh6B3d0btf6QzEFCOA575/0jx2/TpZ6m8vO5e9qkrbDAjxBRxADNgDLrvxsRSs
aPtYNYm/PyFK3hwiBpCka7uhyVfoGQfX15X5X0VKh29GG1C9VHTSa6V/JU5NU46N
wKukBeafrUKG8HONWFEQBjBD4aKKmqSJ7myy1vaykE+la/wVw/MjLlkzC/sIOPuo
dZ7zlGmnynHc3GTrcAjMOVXfw6GlM41jNBhM1SkQzApAZq46khYBct3skP1UfulL
F+vE6vsMGTfsNgiu40h5OoVvCR4M1r/Zdt+F2D7BeBOShxp5lFrZdhlulgbJrsa4
CoredPKFx4rdTRSYPRcI9AH1dNGugsIm/lrtQqRkauIaNF3BhhrCXOzTSlwrH9RB
Rsj4+EbzBoh1BRfgBMznIprHR5lNZyUhxxw/G9cG23M2mp+hiMIThFCUCgH8hKgu
XM29Tgeh/5qAWXzFub+AzciFgywmJI6mXQmSOYaBDcx4Dy0NER4EF2mKpR9M6bNn
FagpYmgAnFSLV8Hwt+M6RWNbhXOxztAolWfLwBNOAOoPz+YvgPhZ0n5tZaZ+TFi1
4I2MgAEFdNzoHfv+HUR8ug94NMRv5jejO3Lq8Eq85Cre2WLoKpDh23iUxB7/sdxN
kyhZnNziWRmnoiPKjzxkvBg9IA1XSbjARrs7Q+5lnkB+Yse7IRASep0plEv1Ze8U
nP/DR9fNk3u5aqBgj57YJ8xzdLQDKrdnN2026DW0zIJv7KK2bf0IwqWk7QP+qiS3
sp2EjrqAN3cYkHMUYxbTAv/oC/12t/EF8u+gbzR58ADR5Ax0J+YCj3IdAeZohxJo
cJXvQd7LqCQWfI8vs/3sPKGoXYy+EnuUhPFGBhWqB7Bsy2F3024VJUWeLni6uXOG
ggvcWDmeZbjjAxGaG0Ed0xnnmR4doovrox+7qU8vVDP59nC8oU3StG6yqr/dfjKa
wFjC6y7owUzTvNnbrTiqwkpBaYO9FwbAutyCIvYxVb8GNtgho7PsDuj1GNg+s5Fj
XycfQURu71l/OyWcbcJvlV6x/J7lYWIZASHxwuN1bv7geLhEEAGIeSYoIjmpS0Em
0J7h64hcf5HpTrs4BA31uwNXrSg2uMSheyU51POL/C6GPv44WA7GM0i/6b8aayoe
MoQ6eacWkyAVmWE8HECouf9FDiiVyjP6+L4i0P2NPBFesIYIGVx8QdWx9CwD10rd
SAsuzGnaGIVGp7Jj1OrJT5KfAlTmlBh8E/qerS3//BotfMI1I4WH9o+09n4a1V/M
qze0tbowrx2fvmXmBe5SUyPrJcTmpkwk66kNGitfTqhS4bdd4M5D4HgDl0S+mbUm
/DBnBO5itIghi3lktYr0HRjHTXXtTU0F5LbnchD6MLuo4UAZQ9/J2yLTyumVFLl7
sLkMotvf+TuG+S06fRExb8A1fQNbyKyN9Upb1LVfPdU8Eq4HznwChurLanUikTor
/8zwTQoS7ET9Ooi0cwGwKZcWa2YgcLC8CIDuxaOnag1XIE1daJ1RVBf6uLAW9D2V
1ib9Mwo7LbnWORvUJnZRXMvgR+uMC774zG1Y4Vwa6W0ivo4s9vovIS4iphs2DTOI
S/hhQ3efYytklJSTyob5SohvgLSxOC3j1kH03TUV6Nai3q7Wd2tqgbSmtc4rMq22
QAMuhzdnat4Kd/EugJnVEp0JOg4B7yUqSLo3eosRd5xVjDvFparJQO2hALzXFEkn
a4QrdXa2n+1Kjm/PwuLKliqa9+r9j/WIe7RaI1LDKjQjr+fOKYWnjMJurw+43pFx
aV0FbgsUqnu5l/rk4l5Lh83ZfwWbEBv77WPhOOqFfF3S5Gs/X3XVPSveeVEuHWBk
6dFe0ltFaZ5w8WNj+Gjg+SZpOcSOaHBMKzk6bz1Zljz/o19AgsDuDQzm/hwOeqQu
gdRP6My1m6F+zDWNnwdwI/XOB7pL/D/P9+qv4yXin3+pBKIwq9uLJWDc9syhpPdQ
bcYjIwG/L2OQl3iuQxl6M1OAjr9Be3P0wrJmwu7zu9AQ3DHsoiQfqJw3avUJuT+4
Z1ni3ZGTctPrGkPhvHJoZnwG2UgM3mYOHN7tRF5B20wKDB+0gZNig6ipjl4oseOX
ou2KhuRkfDhy7HDdtcSpT0HeT6bGr4ovwyn+q7cyAUq5FsJEUxA7Zk4bKLy3F2qm
UMIoNZ91J+IpXVh4MWpsdaXE9q2beqR4RArmlnn1gcKnPgwIvx59lFa3tmxuUNOf
4NLjfUz4ssej4sA/WM+hBFTXmsbqQKxF50/g32YEJHvylh9sU/lq5r4wwSVYU1/I
nXhMN7rLk1ZiDKlZvQ9mGZwRZXtJAJfP6rFnWn8wtjuHvjY8kOUF+YLG2iEaqCiH
uJuIp68Z0YgklfIoJIrJNq2fqUFaBqkAIm/1kAPgswov4Ol0gXBFTsUsJGwZigjf
ODSp+BgD8gG8fOSNzdo2poUxMIUTHAIgTyJaOEpfCPA8GxTMC1px8Wq3pmDz7Cqd
MkjMVN56QcxZSvsWxzhBS3/921gQAOItsLaZLKno01OhqfJvNhkZdp5GaXx0E8Hs
x+FvUWaVcL/FYPysEC/XSu0JmJEBVKVsUX2FYv9m5frUm1qhMhWd9nGYpRKQdoBv
T3WdNP+6oPQzE5hOWFbfqV76LnCKLuFtjxUysCii5WM0N0Mf7lzoIKUjRnIvSZ41
+096q+Ut7Jh6sJuY6i+AQuf+azn0C7akvXzmWEOxPpO0LTJ2tS/E6m+xF/08ljJm
1KBUDU0Lc3FrhEqUHnW2vYAaO38bkWiicBoC3110eg4ygxVG97u9Hcxn0VOXo1kq
KdSrdPzSqkfpx5POBC8+IzaagumVEB20tFAQWinhLMnU2jlcU+PIxv0e/xIFiQu5
8R6bs4eEendN1H+fSqKQsOYibK28l5ErPjA9m9l8YOhdOQOJTjx7PTyijk5oK8uV
n2tkmOfAO4GPlktCMP0Id2xbGgCi1/WUPyY45jWI7Rq4SdZCVlrur81On/VtrV/O
PiyXtRXdr5aRTSeBtwLa85k9a51IhVxFxS4LCCnbLRfQlaMaJptIkJrY/wbN05EK
pSbTdR29GBWT3VVjTc6kF9SVsxfYegwTARjitg3xPOuGjGcHMuWCyyS3sDjaTDqr
eu9Xw6NFa9YSfpN4n8T1rs5q5SH1yY4pMoobFWGbAYisAipxy6tU6UpqK9Lc9yto
E8gK8D03GIxK605W7H0mjdN3KrsEkZSsPxI+L/f4zuOc0AUAV7tQ4PGr2b1UeWrR
9kGC68ooKG/UN0vmWZb07v5cUe3xyRAAtxf08JiXubMIq8BGRxaaztwgKYw/Qz6c
8ONr9VAtqq7HyJi40YVLpAnekC4M7UNsIvYOORvxHWwQRl9dQ7CN5CjclqBVeP/i
Ex23l8gU+GPd2/RTsJX3bz9FfZwWAC+gApZ1aYRmJoD3c9JjxMpKoy2DaHZcSUZo
gmv+D5/BASUHiCgjjSxPKumjqIEiIxvR59vG+H/2UNjp7G9a9UcT1rBzB/KeXlyh
wUJ5Tfd6rI707c0t/uKg4HqfMqGcPhw07QsiGxW+NzZFKsOJzFsLCYUC7zmhVkLo
qZkfgn+Hec0ZA0pfVtW9GcPYC77oHp3Ju/THHpNdzDH4uOI16GoGLL3M+TLS7MAu
Ov5Zqd+yvXRwiocmj/f9B/C2c2h8EJvpRpgLydeCtAznv9Bfi/urDWQoUdKfqhOz
5lw/+vpVQF4qG795XhxwiYAxD5awHIc4wFlYbomdL4nYSPd26t6K4WceS6ja6g/o
TDnXFCPJOVyXWV2E2PUOvwi52s2Lm/S4k9z7jgbYNCKtia6/qRMNOuWSLt6Sz+4c
v/oJ/vMtOPnWnuRJLIUY7sg2kc0JqpIjj4XooaZZZa8/yqLIL2y5uVq6j9uUeTPj
UhYoi83CzyRyFcXMFNZBjSHjLQRMdnf8tBidWR/BDkiF8jVNaUiLz0m5tyq1QkkZ
Dpz7PPmjjcg3h7zTOJ+dgUAyKQfikV5eESFV5cX658KhmnUHIY8kwPlpJVOGyD7E
a8Cx1n6vFwQmdtXhP2y1p2fdf/64exe2p3vfh6yys5VhL3Y11S+RFs5N5e5cfsGq
CbQmrKlvJQkrzMxQhtPo9IyziZyIj6bil4STo1B6LS/6/GglcHTqynt8uFNdz1sb
6VZ1TtlwcrPA6K7D3veR6kJZeQBqvqBoKcqQEwbvvJJrNJwKcCavwbwQ6UABS4Qv
wMVEGR5HFGg8eHNbX2vAxW+b4RHl6zo3qUu3X+VOCqTk+pt8Es5SWSxKJTjlWOav
M1g6+eM5FMVOMgz4GC/LdhUdI48xYXPwJfGjjwUZHUx7meRSh4Ty59so+Pcpa6te
4FcJbxOmCSWz7RZVQmUrdqzKA7rinJhjRRoJu5anElVpjuKFP5RHZlNRFvsweMO0
mnR9RSNMbyOIVPu5i2ubj/UOC3kPj3KFjUyXYWE4X/sB4QyOPDFanKl0oKWmtz7B
qQpov1TZ2sYzunGHP6G3KgG2BGWoZJw01sY+jDn9OWW9QOcunB49tj95OJYRmzLY
6h6Qkg+7R+4reo9JJQYz7a/SGV2bWkbJX26djibUE2cf8yQbJ+WJR9EyeH6rrijR
Ft45sOQsrx5ofObMhD0WKaXDzFvPCeXHp6CZzSN8NdmcFLNX1V2+tguaAZ/4V3sY
JOkdP6w8yrENVFlcCJkcC7p2KaFH++3CMCn+wjf1HBbxdDyg22cu6/leRImVOvd7
nZSUuLiICmAxmp8O19T6VcfTbxtrsgGP8F3hazzz1zmpsOGq2tjmnxqffCEa+baf
xEMYwMpgXNRjPJbTmeIcUS0k48/dWZocY+sjKIn25yEMmL7LpaNa9JjtB+oNI74O
1DGUNvz2krfS3p+8CnmuN2eLihScix5kneUf917D9V7zhNWe47JegXXN2YU+j0Vu
OIxmO9gakXhhdbKOXmbDRDSVP86JHMIJyREIuMbn14kbxTrIFWP4HM4Q2jMRffP7
Eksk7mNKGJokEr80UehTRkiDfNmlV1EWoqWhOk/CfwpzHha11b4xo3QwUh47nh6S
cbC0AvqstZN467vrOlbAEn8mmMB3UZHAwVIPSauxOjT3EBbHFZXRAsVDy/esjQoC
HAS98Ov8LF1hR9xws2LjV2d5TXuA5+skqNkDSMPnXy9DYyXX7vEAVvTUj/2Btgwj
bi4uRr8BMnccnGCk67dwDLw40Ixic2oCAtjlHqgx47tMkS0T0uDR6EbsPF46pSML
aWRcTxWpA50yeqk/ctvoAL9fDjgX7fM+tTjlvs6vxASehYkZ0BCYQH0DxS05s25l
8FypdqvYm6aG4psJ4cg9sSqE5fh2K5EdbNPgOeMGiX/DbGJdKKyl1m3M1urCBG+q
wU/pg0ubR/l3BzXWJQdbvSqChr2zR6E5Z96ZAOe0WdYlPueDGpLv0bme3q63ZJPj
/lDOUBs336TM2B9l3XL62CO6Wlslei+gMD7ScWjwTgEoRHukGKzhczb/Psh5NPG3
hzT/HeXWAK1L7mYUMEO6fqrJO6jx10WnJZ2b0Kj9CNk8FX0fQHO3z1MWQ2Ki6kAI
6aLKVJF8XkEIev1fQ6SGvpNFMaMzQN0KlMjIlWEz6reJjbn0D7hR6baMnoxPYgs4
mCayuBslGHBBAriBXOTtJgsM65/CLqOnWJ9ziAtOCi3dWSYT48k5cAiexSkqcPw4
il1uAf7I+FV2W7yVfUg/llSHgn6pezWIdjgHXI5hoO8ODtMLKGPez0UU6j3K68gX
KcBxlvqnTEezOfdhZJeCn3ZRpaspQ9LSijvBkTAmusyIAIAvLfmP62i5zrcAdEQ+
t2Z547wULrYxjPkJuTkn4iFcsHKZJDkCCWIu0YdcUgkV3Gg4C/0HxBPTUBIqhB3G
PoKNWq9UXA3PapAPFbxylwX0w+NrHELjOY/e7LKKxHmE7+gEtu9GOvgrsTg90xVw
OvYQ9FJs20gz4bsnzc7c32xZ8Uu/2kcjGAWDvVsGPe+na6WPiLnIe8mXumwo8YdF
n4MwWKR0SZc6rS3MAeDEsFAzZvzGoQ2FaQYhD0A9kBAe5ldg6L3HhZX4w3HXYaqB
aZuW7EgsDbAmKuUObnviAVGfIKWorUbde2TFzcDcBhJ4hhP16ekQmT/hUHjNRR4K
7l43gKfjhXe2Rc+jljLy8vp7kRXZFw/NnILhuo8sS+NtyTCGn5p+aAddyeNsuTJE
JkIyFmpXEabCvwq6Hp2pTQrBAS2PoVDVfinkutfxhvt/mxPFjvtmTMmjniMPJ6G5
qOP/t376/sU9Luh9nwi8pjegldCJxPh7R9h6fuRKc7/DzUTQJyJzqH+1q/MB/hOe
HiphNvEzmO86hx9PysFUUkRxEdAZT/bdaVdrtbgRd/hy305Azh7bLGAmU94xDtu7
tJ56CD6Vf9tdGRl60lznrloOwOOaahxpd81aEWOyqUA7CkeDiTbe463fP32StzmH
v9EWLJzRCIPQc8xzXtZ9mLa8q5mAPUpYeLuV6Zf0z7qajDbxwiZ81GlpdP7ll/jD
UVjL7r4vdDALgVd0np3Yrv9ibONp6qpVM5OCRaB5sFg8dAA7+FQWC8pW1mYuLFwQ
14u1BkPire9UXT6cWDiu5uwAFTH9BW9YjzGGI18k522q/akZB0pATn1KmSLm3koT
xx0UOHTk+SrVQMq2rKSMldCfKO8Bb4z5lb8WI4wppl/PitLde5Jr70TY16v4BZaF
AzKN2VhtXYIwH+ERwinAgpFfJcl2g7hdjut4zEXPd/aupC4iJRCN2rs+AkotEEz+
LDmitoxhQCf+ZueyYxm7dO6LDs9TXmoFVdCe3JZAcxhABamDTsmvjj8JNke3rQjl
CKk7YZIJGiNSNakfVvnPWuHfenf2Y6ONflkObhWwxw7qygkLw3uqJl+YzTFmpY4v
wTZzaBnS3fr99WMzn9jqnRqKSfoaW+lY1YQ6ZmG3eyP7WpqlaHmBMREmu0GPc2Ry
T4tEJptUep6Oje0UL2dOPqi3RZA/Y0YF/Y+LAY584VrnnlyxmZyZOlHEOPwGu95l
DloCSEO0aqqJDb62CMEs6kcTCeJlv9zW9TywXX0NEpdM5/EGTszexq19QAymfnhM
QpCJJc/mVUzlMSdDQeEt/ZGQRdBFUUh7ZJ4VCHkTOv1RljFpi5gvV6JbtOezA2Es
xiggAfKRCW4No2EgMqnGOwWpF150L6bRHgamLlnyl/sYGB0+msxPadtcoqCwnvuy
bq2VgJSkNYZ639U4qxJToZ7k3DEPjrr1c03y3YJU5Rlt4Pj8vO1J1c70yw/0jX2K
PRYr/m7Yz/XIqnUNuZ7qyOP7B8NoY3n0NLEe+kGF6twXPtq2uz8/hMuBqIG4lBmB
//MnDr/p0yF3j01Eq7Mb2yV3QivMBbOlg7YwRKAMJ9h8GUmswY7Bx9M+X7Hc53RL
9yMPP0JetUHGrTdS3d8YDvPS2FnwdRdIjQ51rQqhYHa6GRB8ca7S6u8O1Q44sXV0
Cxl47d+kmPA2MenygEtZC8LvJhKsnzvMBkG6d7UYGpdWfxuSM5r8e7mIU/GrzhSA
7MbqHyF+OKLdSXEBrY4+8mJLHbkx8YLsCXHAzhZMnTqToJTBBaDevXEwh9Ugdtcc
TYKRdlFXOHC+0PT7uI2eKjMrxECou0KCmFgs9bpBahOSzjcixuRMPVqUzYlZqbMt
iAQpDPPahuJKpuFHYvW8eyLClFnSrjqcCpbfROGKavfZIZQaJt8zzbyPiS1x5JLS
3RnepGf87TXSmDEH2ZeLRSaorYV8kgi7VtA+50RRpo88qnq4PUXbq9UVqgwAGnRa
Cqiv5Uxn+hluHKpK6qG0Lrf1usl6PJXjkVo9RwuQz9U7L0R2UdNvCLPtj7r9Bc/K
MOZKfSzSRbrEeF8SgX3caJ3CDwe7q2wJAf4K8SNQ2Ph8XxRnvo9KKkbEQFs0hWhV
XeHGwlPLEP4aaKbC51mwIOypTYMH+oYAt+9PM53Qcfn+DMsKyzAxu1L6ApWypuSY
Ffh1SxAqciPGCMw6R8evdivu6A8CBJukpa0osxsObyaw5oQE2Zh/f5nFrhth9dV5
7jdjXNpAg6laNeoZ692Uo2ZriFTrJkjF5vlopUn6TLHPFeJojXEFZqGlxME/SVyP
HFrj02nNnUj8/N1ww3xucd+s2kz9fyiWX9Mh1ZlSfvnahEnV1uc7y8p9ruotC+eP
M5Hb+licE3Ooge6xAQG8A2oUZOoWDHls7YN8SLi4/g6rRw8pAKsHg96uXpxuYR3f
zRDGD7v9Ryh/T41SQmD81CDes4P1Fo44V04GnzlOCxt1MFemAvwyF8ZI6fTpSLdm
Nd8j9eOPlMJxWMNn8P9f/NIwzYiGDhyI/DHZyL9pDVL0sAKvzwXeubXTc+7kh62Q
tHTIek+wzn0em9URqI4UiH+pPQt3b5J4f2gLNiQkCx16utKtLOfwbq+6GvrYJpd8
yWRKFvSIL5EX4LryLUV/eaq/fN+6fWGgTY4iu4Q6CZGfhhoZVG9jYWzUIn5v3y6Z
RX1g9+LErdPSsJoF9TQxmJfikQmvpUooUQlMuOZ6MwI/j0eQXewlYNI/ys8kJCYk
OucstoNSCjO/YN5wANMkhzpcY2DRcrj+QY5fVKMOQHSHTq2hTTAF05oDtWut++IT
36sezQpAqtSWHXM6d97Mao8llns2HKpKyQ9uvUMzLachyf5i8gfOOgjUC3sIapXY
Uf8UwQWmwBXR+QGfCnJTFgdeOo7PuQF2ynIblJf4QQxtyiQdj2UtnQnbLUmXi/18
e1zZft8nN1wvSAOxvb7cQWlTLEz80s/cDoyi1H/9eIMQl7PVWNisAFS8oNEmkg4W
5844xufqcy3IRIhhpvI0NLt/aN7y8pgdtVnbwO6ZE5r8uwrlRhzm3xawH0B1D+za
WUEwWF3Sm8BMBfHzTl31E1JsDikOR8Z8VfXNfK1dS+Po9XdxnHrT2oFD0siSQQil
qbfretjpYe5/CHEpDwg7HSxN7uWTtkg7f7GHvFI5o2ej0eUme2ORbGLbwPUI0fPH
HML2HXqziipXHJiM8G6qpInKRFwjuG8TG8hndOdPfdXTlIM2ZTEl3OMjHJVvRhfR
aAI51XZdCcK+tMnu87zTeRLHXh0Nq73HPhsfOE0dljJSxz3T54qHUHjq99RnrF+R
cSVM6TrTMUElEgVNr0uyHx76E9DqrpNiZjjpNOmMgxLlcK46XQB2MrgDm+NXv97A
1HFZI0KHe3yd6Q75P3Ly1Xi25p3+n/zPYtDjmkGiV01RZP66FJ/3t6GgIV2iEghy
2El1V9oWXPJ6HWOdVDxlP+CqOKnLaQ5fCTq3aWEG9cIie6wDvatIbu0z4GfjVBV4
NVdo5wCHTKwk42tOFt+ejQcof5oCslqm8m40qK1+EDdIhsuNDBrylnJu7wPfLaSH
KKv54DOkrh1U4JBaIowMbh2cKg73iNhtI3i6ra3xEeRKqWTnsb7+Y+3E9ToE9eDB
TprMQ7xAWyb0lCRwK6E6NIwbX4zh51rI8wg1H18x5wQJx5oAeRh6rUm+QwpqaFyp
OIdgfVKtoB+pN8hfEWx//8hC4WT0JpKmPOFrbCYegZ081k5TaqnMoCz8QF4wvmCX
gIEPd3yXhnL8RcZ2Yac7EV2irkueLb9Ae+9kheN6yb086aspbezkDrBC/VLvMPTM
nIyTbbKS3L6FP2wPfIiqXd9AbDVa8Ik6c8zyGdqceMSOcUOCF8N3zIAzoH+uh8om
4XT5uuWYz2AU1gkw9ZWXh27NhCgD0lIHsw0IIiH0Ch5k0LZrdvAlDo2Xch583lMQ
YWpRzTjP1M61ANwTvYLHFtgVd0a8A3qSKcPjtdpKKsxpuNCzFswgavLIP07Nk08V
D24hbiGDZP62+SVNSNvVZPkXrcoPd66BPqkud1AQH0TXhGThPgoVuwdTUM3UQFe2
Ysn2SfHMKFVBE8Ap0yi8K+TU9BfG3R45Tns6V2qYpg+OHuoHK7kwrwQcLBvhLwX/
WnUB5ytETX18KxaBORl3PyPOHqJl2lHsjUY5UunnnBeDFP7O8dTjF97FoluYXIVw
sbVKtNKQen6qJ6+RHGY4DR6bgnCOt+ttkkTcJwhzdqLvWlIOuTdEm+psq9B80E5F
uO4GiJ6S/BT3SYs6Ipwzc+Qytdj5P0t+ibe6e0q3rjhQc8zDDJGuwyRxAkM3lquI
EKbJTL00cQXhtxKioZBcvI/dYNZp5h6lshfL4zPUYc/KUjvCpT2e7Nd2CTQ18b89
0AAUsjTfMM5fxEKYIujNgTUmxdSWTh54y9KVhrrkKpLedsMtieUuj8OfTHk0jbV0
rTTm8cA1lVuYs4lLALX2JR0KGBgIydT3C5XLrdd9nkQ8j63A0/ASGYPSn9hEqT/q
prsCxY/8DK9wJRSicxqbaVJafJ7pC8iAZgn4m1UMzbmbDWmGdpy9k/sCfyZO3ahF
W2KOSxMmt8qO6O15jWWpAWOBkn7M1mS/fmmb8mtIpTDyV+cMoTWmtxWia9AMSRz2
xgTwUhTn8CEvsLND9nfSq2OPN75EYIcMc3uDfGl6zgaRpWZUyUTs+KLn0Tm5ygjE
dfAcxEk4xYWfGgEAmU5f6LP0I/hq1jcI73WV2eED45LewI8OsrwKYeKgDZCukE1w
byzpfzZGX6+wfyZHuyOQZn2i0wxnXtvEKdeVntlg6uscWnUMDGOYUsLWynYPxuLE
Zw9cF9MQet2Mlvq0nvIJ7b1Jv2Krzp/kTBqjJywnWiDlfdsgkPmumcTvVL0l0tqp
X3GFkzzuMCNYvV3u9LsoDXwcbrUekZGLP55qI3mI1J5QC7lcnowjnWOJE4KhwxG6
UBHkFDFaXH06oG1bN6wwavR0LGaKJVOBnUnMvWQldaq5ADhh0sCwRTpJPKM4CLCK
hNonUmfGMTRsdMcQqxMU1xLGyLf9w+x8dDYLWFYTVPDCLFI0xmfsxUCaT7GbTWbC
+67rxhrw7gxPVp9sG/VSSaMhpab6n/ZcNM7/Peqvy+iZHOSvdNYqlxB7W+Ce+d3+
/qw8U0ZX7a9aBHZr1y4FHH6DTC01/bl2KnQyUU9Ssxu6gSgRmUHxL7y8Q/H4Amn9
W1J65DVbPimCPEvjSlBy+J3ob0j/z9zoQa7FyATTpNpqpyubAEDB3lI0Jz/qW74p
XQxcftpwfyhAoaD0NMyeTVJ09Noj5otBZcAKz8WStJ8gD+QkTaoKodctVNMur4jd
fxBL7R5SNyXuEdBUwngTIw0el8NI97oPaHquD31Fvp7rWKzIdUwx1UjfpnC7W8MT
1xeKxymRRMSsrfSGbWMX5siKVBxs8NwVEPgK4Q1oJOY7gzp1j3BEbYVhDLVBT7mB
2n6uJcaoVb0spN6+O7L/GKPA17iv3T45j/+bSc/hdaAW7X/6bK/v3qw8mx+TNkUe
R2kcO1xt6QwiTA+s2MbA7Fe5k0bJZNain+WzH9+BLF+7ZIMRs795XuQU2OKfEVDL
/YSl6pEdGiLVoTPhZvs4e67Z3M8SUF5Rzaa+frRZsEuCbsW4/yZOLfwgHy9a2xvP
sLT72vp9SrOBrKMRSMeQ0ljzED9s/M+sIaAv/zokqagR7cUiSG9F+QfdqIaNvC/R
J9/3eTyza4N9dvVPEOpfmrsgAyS4HOqXQ4RXXTIxqnZh+C/8cSFtsqL+qaUe3pRx
maBBqXUEVaoXlr+QI7CCry20vdZ507xOU7ndZm+8gNxUH0k/oRGQJQASUEkWAwDx
OzbCAQJ/WEK1XnexKdM9OMPHYmTpLbVfRrP4nYg4zP+IJujvgO1oXTmQK1WOKRzZ
Y9fTANvAGow0S2WAGlKlTxKmbSesuL4orUly4pffchXsQQCjCCF8BBbrLpOOZ3JU
WektH48j0N0tNPQ4c5TnXyRX3fmvVGfPSRJRefhg5Dg6vy42J+VpteldxcaZhcvQ
lvtAxkK06woBhwhVLwSlNZVLz03EmPr88P12yRgY0B9CZEH4MnK2Dch3b26Eolx4
duLzyAKLxV2PA10Qp0bVUrtXoFL9oBaA/pEBB8krsR78GhQPkN0iuv8/ZgN5/NGs
aqyuQB3Ln2vyU/id7flcLuw1eAn0ZwO3cMiUATyxA2RvuXvl+tMd/7L/YFFdOqau
+gIYQLAxjwp+y7YQGZdtLQskHSFsKtRdFN2N78MPY2wgtkuaAoUeLbxjXSosx2TR
DO0bJm52UW/cOhJXbe0RyqZo8I4kysDyJUkgCk/WsvvJ6CMi9UlGOtM80QYziSr2
1QaEzcuiSrPGo/hS4sBC77s1oUzCd+TgsNbuNg4lCPDnJldC/uCTsKrRTFc0Sk3m
crinA4c+IcWZY+bOZMbk4ZpKBQ+Dw7JMHpCDaSV33L9/C3drqndxK32ea7ciN6Q4
BlxDe5rrCMMPypwJ/IkL0yTYFmHmuo4tMbWiG+t2jqyVElLfJuvYZC0DwdOy7I8D
2VLvEZmRuZoFB6v+h50H9uL/WeP/8rnevkxz1pCGfWFhLSMhZzLTX2p9lJ6ug4Xi
YrAD+IIzHe/2HDtuv7AzlKjHMcEGYFIAAaIdFEK9RwX1TB4pSe/WUdUImnouw2FJ
c3pv96wdYHZ/5u0ADi0vQqnZ57pNhuZPtP7CPIgSU2ery5DvogvupEiUrW7WiHUu
CUCBHLfvMZoTHq1MCBMzfSqdZxJhurLao5nmlSpw44CQkfb27yoK4YMAkpfszqRH
g54HMNNFrvESrYdJHxoL5YessVBPryIYVzVPrYkON21uPSyondtSO6w9AVLsGHaw
nSIJ64hYApC7KKoaAizWg3EWKfSKKF/dpoM3JnHTtzBET3JiqOvoObN8DXHdEcNC
aU61j4UFiDqOfBxZhKX3YiL1VTHWT3yyMD36Ub8M7lLZ41mIR5WIf/nOn+DEZGFk
U+Pt3M7R0tlsLqnqNhkGgCm6ZOkgBhcbhHPXsK8CvtkIahhuDuD8AftrbtqrFH2B
oHD7qHQR9k+pCTyL0t/vp4dj1wKV0gQGrnWuAq7aTGJvFgdOn9WPZ4e2PN69WNcn
drkVPsltn+fjRzbYZvYM+yRy3nRLiq9UU8qkdOm1PQwAN3FHYDvHobpslWGwz/ff
8EMVXWtMEXoU4FHxjUoYzEotmQUzRcAVJqkNIRsmKOOJtzP5A/NqUFt79SlZ3Wqn
mNKZGNE/5xEIBNFekf+O8t7xkhvfaBjOUcJkrXyx9yypnmwPqt+pKx8mbFEllDio
Jqm0SXLflAuHUNGPCtudb3NXOky9kJItKykl4YFJ378KNrKkLihyS1DZVF1o9uQi
Ln+MTx66QoUHkvlvqdR+IW/RzmO1HWf4roWjZbfGtRovOy5e8npjXOC5erpDLmcF
MzNQ4VWjpFRc5soTY9UDH9Pf3Y/6x2fMzNnbBjopP4jA62TaL5DX4+GtkZjBKLFM
xfzBZGbs3kFP5G1D17NdQjpUfYoA+lfM48EkQHomGEfcymHjkmEqIkgjRfKtjG58
2kY6u/FWouJr6dr4f5yy1w9g4Pmxb4WaoPs/AkQ6ribsyVkpKrZG8H9wXBRk4E5y
EDTSdEjO4ZMnzICoH8x8mwEq6Ykx8tJhV23RRTiCy9XhBizGflfvbF7UTDBDYcrc
IICIc3seo50AWyNvBTkA23mNiWzadvIvjklRiJnyicsM5KBvJJifqF+eZhWF5cyL
djtQiUt7F5qDdIf8/yRIhFJJ8uxKfw+DgVxi8g/FxoVkKCP7+s/XfKcGVMwHuv6c
eFL7RStCgR0u9Ls28pZozcjT9RSkUItMs+Bghknl0iWdJwqYF90pj4TD0ZuUzXbi
BAvjL9xRpdWWG3sdoHsQT2GEtx/EdHGtYjuWFdxDqBSMedp9vMiX8jQLZwsT+RPp
KGgEKQ1U8ei0lRz8pYGfGHWdyl6h6f+V8DxaxnkVdiZgf+vhuxzs9M/MHHhPXFNr
wp8VWTtwYFbVOsQ1nNVE/1VnYRVf5Gtyuv4FLLGCPZONOGJyIxyhx1Tib+wleCoG
4bJKc/AR4opfEac+fAbcPBaQc79V0aXzlfvKKtUoK0Nwgx5HDpS3ppCFTtIskVlf
mgqKt1jVZUhp/PuHEqt8LtYSI5gT2imt8zmjoO7cLVax24ARD8khBzeo4IYN21Dd
WSuOFyAPZ1xyVblZ4VJHCnAgzUxNHYzEICLEoA4P9c8AhWBAFnbBfaw+Nb/Lkmls
AghGt52QhVoQWPl47y/INiDvu+mtvg6/PnPajyuIUClzlF1vwjRoIlY3VgSsFzMD
uj3AEizPWTxqXmre28twSbaGQf3Cc2AzZsodc7RtNCI5VtmF7fsaSaD1N7U3yMCk
46PIqeJYvHnta6Ko9kFjMppDh6tHkw7YW9+U9kKXVQBMfCfrZIhQhl7mwbyxhknC
loHtiPZi/vA714XoGRdsYglNmejgUQ3+75vvmEBFmG0HvRCMswfh37DKp5zc9CLe
zkXrjxhbqDS+C5Txr//9VYj5tHfYFzt5ahbD4TyecIC+ka/fGm4EcdGicMIEZrWU
xtWTiAraRPQfZDwqPr4y0zxN6u8v0IZI/Bc1mMA8DG9+vAKmBZrUKT1hf0qYlC/T
HcvFuTS7vMFJBmYGr9vAwCMAe9kL1W7qWGn+zt5s0FeLx2lWMRwy3EqRv6GNk7uz
Fz2JbFbvfKSo8uCbv3V9aLIfKERLSun/5JgEC0M0nTgimVfS5fDMCbkcWfgBhLHu
uY2HrnACXQMS++ekLsX+IIvGkxehFPWGlV1/+p9gBo4yw3thlMfUK7S4DQne4g5C
BhrTg7DJbbcay8ZDdj0YM4wFpLcl5oblghKqY38FRZcJIFRip05sT54Y1dfcjRzM
s4mLw5r6CKmASBHFzfHg/NOln2HvqawEmJCc69sLzk5F8DnYxKUh5ReOV/tBzImX
2EzVsW7Q6KZGm3X8gZnn7CSXsHCaDd1aCa9hyUd3ulnL1XofKyxngCi07X1VCbZd
/HexW7cDGXYJbxaSDxbz8OULFX0aKNvJJO4ETDzEJKU+LFBwKCRR7jrmW4vjXfWn
arbWZHRPrzCCpuwM6kYBDqoeiQO198+VUiFFRbu2Z+3mzmdXUWszYNUwCX3lMrgF
rmswRJpyE/Vk54lTz6py2I38GOGQAOLegBDRByJWQAzfePkGaZGUch4nkh36BTnU
2nL9n40GtzMuv/FFSIM4WYJpkFVweIYNip/px4o2wtAhs44+FXbAuicH8gO33XEn
8572K4+TtoPoEo+88yeS5xfeLmncdSZQ4wfia0iHP5NRweOMndrdex+OYo4LN4lB
H7StZDtBKcrClmsEKpBtoABqJ6+u44kCWIssa4I60r/qauj2/aseNYmbTfg/DnoD
KdXZCdYQ7wQd77IiQBQ25wJ+y28C3pWRbxLKO/wTYLUV6jXkgxSgsXkRerVOBU7V
qxQh5L8aAF+1keUXI58zhEH79BWXsO5y8Ry5lLsmxlA//vkVFgIFQQSCVeWV4UCi
ytzxvB0/TnjjYLPU3cjOR2LCGS8k8VeXIDc3zGzw22vjgp6WNiXWc6h1DIBM8wbN
sQYsih6uEItCrsDJXY8sE+4yVzKd9vV6Z3sA2HpBl8Qi6v2Uqc634TN4i+MFfl7b
7VdeZjG3p2HmE0Ro5ylXd6R5uHVxRixj0Opre3l5XIaZjjGhOXQdFD21tsAiXTAf
3VmrWPBk51Nmh3Hzv2tZxp7fReUhn4cSMSTWR1KrekthgEiMlbHNnNAiYs8ZhuuK
1FE2ko562X2hurOiXYcvj6Mkfo0fi5tecjG6LOcqJGIz0mbqgYfX65tvG0nRNWID
gOTNtg0nOLIstsLIaIqsoumhqjdJkEdBZ972A/fqx6SVWb/lj7szH+w8SJjOdM9r
hKTJu88n6JrJXMbZh71SQOr4bIsl86XjpdeiRcpfqC+1uql8IzlGDhhWoEKj3H5I
HflEoiMvdRGgb1JYlU70iB2fcSS9/mpSKdm3APfSSOyjoA+w5KVIh8hG9+9bV+0M
VkgDYt1FXWKz2kOJLMKo8oMhYpvbri2LSJazP4qJHDOZXaLeabKC7HUwQRFeaPpC
CIaOd9k7Fp/zA4IQX7k4iL5GtQTLDk6pPjXmjr4X5i3kff8JDU76raKADsdK7OJx
FIcfna4GqmSzSI99hlhL8E3iN2rnAx53aIstY7cup3l7Os9wtU1CFvtP2g1Wn+ti
yeoLxvb48uhUPdQAlP87fV2F+l86vRiLJnCJuA2rCHD05QuQXZh/gX3x8bc094s1
uu+L9s9rPYF4f8MQ7HE3TqE+lnPSrBSMtkvYKrK940ZRST+GUZe0LtWr8pqH0TEo
9cQUY5jQnZrtM1+oc+SOdP4jL4ddmYGIchVYN9/D9Q4a6WmLDEzWQzLH9SBrvIOG
YRaUMU95ir7pT3HxcWZDZvDri4HsnpwjP+RMzvghiPT0THWJcvoTv2DGzhR282hJ
Ue5wIbHlRYUdLTtFVZO7sCZk7+TX2t0gKOuDPbVUc5rwsJQodP0a2nC/1gRu7QF1
kOECnHvEHUxJeZHcp14nXCKgkZeuLR2Vk7EW7239/HE9tBBY7MheewRtnmuVqgMs
3ahrTuJoK94601PVK1Ci3b586Cz4ubIEVGaOYDfon8fVb4RCR+UFpZ37d+CAhMLU
L9eOSYazmZ23Vz6VqASF7IPBaD1B9C252JbHVtqIhXobKFxZgzwbySQeaKWnk3KA
zINcEwzkvNCQ5V67FOECq7xoLbLX2bnVu7QA7H9kP4QdQwMu/96D9mSOZeye2fiB
/hRnEUD6XGjrLCzKnqhpfZC1FDKRij6rhnqSC5TWJfoJdWWjTBqce2jdeqsm+R9/
i7ZuIrgQZY6/qnTZvhCkZApRHqPBHZublmRc47jF+gGQ57zrSQ8qc6VmmfdBRsLa
i5vTqYg4NgeFN91rS7EEEwFVE6iql5glAPKr5YqBpvoRj9R9+cTYLaJrzHjN1Z8X
hNobqehGSwyogDOGNPdNOZU8JXXK1bPNn5hpNF9MHvRALeGg3AfFUFgujdJUFh+C
IjAGlGbjUdKbs/r+FtusF0jnM9rFI07VJR/SjtzWsx4244fB1m9Uw86AVPzuywm8
3iNpcDuYyXJs6vt6EPxuRCXrHqDSRs5hjO2pUm8zx2Q+lX9J2CQMhbLh9hdzOzrG
kww+79a3NjNdlvAKcwyGxI5rILOy5tK4B27Imezn8rkts9q791pfjWxKIRbhm85X
RzoEw5IV9uVi2uLRcVCVi2rBMbCW7W+1UlUnee/YOQ0XezS0OFT4zeN4LrdJUG+e
rVaD3L31E06gt7E37K6VVWUr7xyfmWdnNUVbat4BRd3oBRj6wXFMCHdozAEAOeF5
2SXMHALXsldVwq4iGDFUWzDIYG7rLIJmo+b4Zpw6PPXHYNMQbOrlRLwPhC4K0IVf
X7tke47knECywcY6hU1PY4MHvegzQz9AUTbL9mL0YQaQ2scpvwNiiyqLmrkmP8tS
/BsFLOEXj+AIEOcZa78vbAkfuIQJVZGby1p6mG8V28LJRe/zU7frzlbtMmY0c6L/
cVr4J90HJIRAgsYYKnfzO+/wz4RCtqsqw//x4obq8vpDQZqJ5XZljLDKEadxPoA1
SWWeqRYc5lfw2ae1KXtzV1wGCKC5JOyIK82KjS3hMGoPSDe7IHDMTFaIHcu6sF0x
MCzeWK3jkdsO9PDzJwSmicK2v0BCr3WCUXoYXj05xeqZaMX9S/yO12eTbJjVlN7H
X/eSTwIAZkZpXipl8CPh762OyHnv+4wASTrLs8XWwka0UI7oXxZvx+Y6yFSUr0OZ
aB5Fbd1HefvyG9mnJ1Sn3jZtO/EnBAbOyg6q8IuoFbyF/dADUfnB1s8vw6Szrrzz
hx24+8RWGSn0Y402/lD8vBDD61GnWPjPas+tU/Lb46RTF+b8e9qDqXrBWGsfavix
9+Xf5WpAseNXRu7MPT6yzADFQYTGDXGtjTpdbqD8XmXSZkIpaOaJSQFgVeRk47mg
fVscjMKmsG9jIuxKnA7mOPEYWnoy8dUlz7EJKI3btXmhDI2dP3CA4Ji7yXhcnaw3
EaVYHEMYNtNB4pIH4DXpUTWt402InFQ9u6SIZBhZadykjzH3/5cHH4vPU95naVbZ
DSAjIVjTSwJu+Gw95hwa+AVlHiArDkNL2x4grG1UqE092mc3XJZww4Z/A8LahBYy
O/2inSp5KSk+4OU/gOlcFQtevQLekPE27z0zGka8Nr4/6V6f3mHqILSVYDa49/Qh
IlT/FOsjQyLt9uTwJHqwvGOCARF7fTQqyvLBH33j7hzwrxLu5pyBdEnqUguD4POA
2IBvv5wTpXlF5igve3d/oQ5ZKI4Ub6yHUbniXewbP9ISzl2iQSTdgXylqTv/H4S+
r/c/7aR99flPwX8olVotxINiYommdG6f9rwXg5kt8x6IRUFI3O0TpTzmRQ/lnr1C
uiw8azn/cW6hX6vKFcF/RRnEktQFuMkccBOk1t59FrgVcl3gB1oPW6xtfeW4v8aC
TislHawH/wusnH4LrPewYPxmDFnUPp1vCxpr792Yk/8KvZtFTF9xNTRe6BwWmLF6
i1bj0JQHplTAGZnRODH5YY6f3ay/wHCaw9yrxg5ZlhlR4X5KvmU4AMp/10MW7f06
DDvHMOY03ewYhc0ujJgfIQbj7S4pKsHmIt8OPXpIHwGnqRfTqyCFfZVBE90/xqSB
fhv5Za1Xa41WyeAv6284CB2BN7jntiRCMRUsQ9cTTGfJF5LCXGGo9taATWre/M8M
T4ykrgm/dn3mqFA3w3irSOIr6tuwVSAcZe7WR+wi1GuaKJQ2yIJgxu19kRg4TkGb
A8NFuTw1zbXQp+shzxowXcb7vwA0avKdCuS+qeGVkDdRFtzN03Djb4MJlCEvnxe0
P3A7VDIIq8dEWDjnXpGiA/QgkJfa1ag9JT+16jYMQTa76aUIwCge8Azvv+8MSV1w
Tuke/TLRAjUNpIgforhPUuvMJCXUlJBXaijL2f9Mdc5YbFmvTRW7qJOOqP1zu4NT
DqfuQLTUQuAzY0Yq1Ebm3OozFkCjZ3DKXJD/0b6a/MU7HvD0AQbzZVYOlHyzAGS4
8NDNWzFn4/gfkExES34tktN2QQ63Un/lxY6SxoXurL782arJN03tYU+twbzD7OcW
MAVFGz+86xESUD1xnWJB73M6B1RPXqcq+UXTwMNIcK6YBaAv8noVPjl/DSpaCUUY
uUhc6YDUQEhB3rZgLGCVIahgm5gA5/aFCC3FSzsXbZvGY1Ma8xRM6gAQ/69u434u
N3AwjY65HfaNSs1qe5ZclJDrCqp+L36GsNDiK192BI4azRVTudS6pfsgiG63fjNL
VgrlRBqFf7tp8A4QJLTc+rGDpu2iqKzdN4c59jh2bYvPkmPKrzC6d8N6ozxsPhZ8
32LwCYRMnao5KmSsgnp4rkuB+qrpuB5wgt0W5Ahu0D9ra8QvfUvkajK0CzeCpSgR
6JVHjoPtlYV3HjHQDYZ+z2lGq7uuUe+hqVUMYmF+zWiWt5b4hsAbvU1MDV2IlFV2
uOHV99oMbzKiJu6aTuV7/y1iDZvpPxBE/dZxy/hMxAizDXKzHgdzLH3Ij/u1yQcY
drrjcamEQcbae5otRWzzoax6GQfthbT+ss28PTcVTXhdoG/h2mWkCZVnVsuyjddP
3F/wwOxl0U8YaIQKA5V6BrlwheK64/QaLUo1DkTtQ0nIVe3v25RDy/svWiVIYZMP
hTiCZNamZzvrPAkrJ/lxcRipgNzfup/rrgeAg2yY5MBKBJraOIQrLrpnYx0OTCym
rircQtSIbi/iBxD7w5uAJzcp+sQUXWXtKpCVYrTmeUKrpsdHXOchGOzy0mXMzQea
sOXmC/DiBtHpKBxGliv5U+bE+Hjpcy1rjIxjmQUT+RtunybCexqiUqpp1wI4wsef
p70ae/9/thKc4eefpmvP+oWtiQw9/HeWfIwELBfPAS+xZ0QO365U4H/+ad0QGGXl
yFvgSNbyevCiA+eDcwHH/S4QiIDqoDGqMYbvsmH9r+7hm4M1/d8P64na4cfGRgzI
ikORL+egD5sBcAT/MH4SofsOoWTHuvC6xOG5afPhvo6Cr3dONytlU7sGWrjXnOVt
K1lDtaT37oJYwdXBe5Fs8fKhNdYx1BAa/rgCgoxGILyo3fK1nLXfMA5BP5rLAH5K
Grs25VerTm5MAwW97qrSu23He6AUHmxx5RRWPygJQx29N30oxsHxEZNfPhTslxtt
9cdM9kRbHAP+rYf/ZhZWKUOrj9ciuUxnqYQuwnHPibZD9RuF3grFf6G+pSlboNYT
rbYwQuPwsrihy6LgH92/RWqUUU4EDIzKoryYnO43ko2xx9rxX/nQlw5FuiBQmtvI
1HJ5sLrRT3KJl2CJCuJdVC8yr0mkVPk5FiqWVlrMqEwro5/9L2whb4uULoZGwH4z
obl7OniqNJFAm7CGLL8FpperwJ3uiDq9ws1k4kgRhTs0V3hkwu1e9YtHnB8J04Kw
vV6Ki/vMUc5jEXdJrZp+t3oJH1mw+rwBgUPC5MqPf99EKs7tNNkfAvB1CA5oE+nU
ckGVOVTshzl8KBnhG0YzP6JLZ/uZ873DsrjBr382MQbDOtsSYCHuMlnG5NJxkKF0
8xf06IOga2Do3iy0rgKXz/xFi1IaZBGd/cZyA5++3ZiDrA0Nhz3ISbYBXGubS3ZC
OdWoaglc7sZeaqKAl4tcZSdxiEt53n7w1K5j8d4SBYykQBAlGWy6m2iQGdGO+xc9
B61wMjR4hQlbAg84I9muexdCIB3yXpHxjPLsWqz1eJG086fts3zlaZDUMc+ppcJR
WcWpPvjjMC7NjvKTV2hNkyKQMXGvnBUFPw4Cp6UFu8On66khEQ3n4vDr/iTOw9hu
Nuh+eBrdgEYZcXuqKdE9lrhxO63WFpoJKP0JqJ1nSn7JkUzSSzFzyrs+a1maq5my
1z4wK0fLL9E/hom7cURZkjePL1PeC3VF0Kct3HcrzGI/uJYQr7qsz7rQYZzXnNDQ
9syB01eMVtEjB7oJ52HTWNZoltQstDYZLCWXKbBCr+hiy8uE2npMT1OhhqdjjKu/
8LT5ke8SGC1SKNiQX0bQOaMXfxA8/H+4reLWb+2tfn2OvhZNCKt25iqKcd06Y5C1
r0wA+bf8nMEtxVL6k1iRk0g2pBcrBfb97Y+vPxCNyXF8P40Q+qeCCdLu5Y9+H8vx
gljPUSnFBbwou8dC4xOv/+ZgvIsYEm4N/ImpX1+3CbEK3SCFZTortQz55KHxoUwI
/RtpY28kpp98kMa6lBVpFnVxNNor2jdUydh+XRX2JKAMv3Pr66XAGGZ2eG4p5KbB
YgyHkV4Um4UZdy5VCVvzIBtp2YrKkMyhsDdSx7hF3NBFHzLyaOzf/cFdDm/Dx2Qg
k+BCCVWIcYkl0rdAYwVoNWiDBaQ22NRmdpELP0jzOnmbHzsBC1qZZB3gviv34wJX
+9RzZjcP6daeS6aT1gujIvEojEGD5F3SgA46Be/tqerNigHXPwOK66Zr2tYNgfNr
HG6VoweYEXhUHoKVlS7XNA0iyaaUYsSUMdNzI10SpbteYOWkq0r/WkqSFIzGbyCv
26bHqZa8UMFlTBIgkgcFx8w0il/6OGRhaO5va1mhht2XXePHriA0LM+905kd5RtO
BTBGIysseJnalZBwFGyA1q0GIVtKD2YcwsH1TJ43xFHZ/ZvTGvgSOUQKpHkdsgjW
ch/xpy0uiN4gGvWDqj5V6RWHSPAX5ETyA9WnCuC4rXUCTWhfQK6S7mckM5mzDi6U
hIl4x56bWaDc0FN5ziTqDtGUGgWdZXONgRaNafzD76IMbMleV0DLpQKaUcCeJL+M
IUREIPOru7hPMcVTK5DYKn/6my1nrME53acxhRdB6vCrMVOjyEXglEwHYs3qbik2
b5vSF+mqPBBkxmh0M+1vxjFbudOXwM53t3Fy//vlpmYMqFhd1CPDGNAHaIvPpOEE
HmnSb/ZPLDv2T9Bjl81KljeY56xm80cFEbOs/XV2xeJImGI8GWe86uIA+4HMIRHb
ZXr56Fbeai50+ZCQJznDoXkBE+6p0fp3+FUJGQoUqrtHbQm593Wh5VIstNHg+sQw
TDOtR1g8QhjdNyN+6YevPoc35DX6GSP/gdkZgk3EHpoS4jxUcnYDK95RMJ1ghOTe
Ase07+EYEJJ4zitQFQd0L07cvzuAEGyWzqR7gSWFtP54W9aHrXEHKV37NNGhybOM
Nxo5GJ4Ib1r58vx6IWYy/49aFTGsBtPGGJh5A5EEZuw5XhIBpJdKLU8JLTMgf+3q
zcQcijak8rflpktMIf8pgF1fhCRH4d9lkouA6CQGoT7mGWX7Ic511ChTveHLaZxn
1r0cKXk5vfl1pkIbd6TWWRJOViDFiqmmk1nnzbBTH9ZsxBnk6C8qEQ0xu6VkY7ZK
lCInhtUSI4Lq2GvKQr9Q6Xu6AwsXfVC1drbKcRXHXMLY6GWG5k9ATFKWtZLCB1GB
nI7oUtIL792aqth/K4R6P8nvsAVQEK4e43ZQ3Rzwtvqkk/saiTeL0S4yI0Ee7b6/
ayD4luYzZ8ajajzUSQA6hPaqLUDHstn/gxgkbPLLtsF+qddY3ufv3WYnFxD9mTcM
waUQLPoxy564rV2oeiuV94T7/8XmdS4h2AoJ3AkHRWMXSTrkJGU/Ky+XUkctrZ87
LZSWpqK3zU9HmoQLNav2MLuDbaDsRVMG26VBOWJYVEW3mjS0ETGXtXOmypcd8uW7
p3JFig6zjBNajYJ5c7/kS0V135eBdF8UDniRM0z6jR0479lStSUAB568TIHCnhjT
inlExCueK41+GS2W6lb5TGn3TFNcvPjguCvxkVggc1LSY90yi7QHxAhdbL3LL71I
/hi4nEAZLP3KJ05wbyZdXNGSQJSzKkgWvbU38C/XHBCYFkWJGeOYKdsuGvjqWj9R
i+Uu80jbpwHklkBAK+PQSxLCEwR/7sPHbOpgX+/fCsl0EslZCGlKxor34RWKihdJ
PnEvpG8poEhLJOtOn+R/cHr670BN3H4S5WuaoyKnMAhkL0Kub2QxGAP5gCOpYYJD
n8MD/cXW4ZTh4bPWFBNBcBlnQz/o6YXYD0VhRMaw9cLovZ/0oTwh5PU8Mv09htAb
z4j6BpEkaNkIyQtpTOuDKhe0yF/+EOvTmpJ/sekJzT5oML00OsEKtSAMSa78Xvkc
CKxunszm4EKGndj1Y1o14waB8Qh0AhLSOSzRMwP4pzN2V/JVqL25aIqkaRjZsYyY
pG/dOCGFBbUyfVckQSEcIVHH+1j30FcnbJupTxlppDefwkgtyYJcPHPy2LUkr+vo
jHFi9BedNUl4Ld+gqdMWwK+Lqx9fQCCkW5ofd0W839Z32xxWqWXjPENnQS4VfgKY
elMQvswQx6uc80olPa9pdZnCbLU8PHJ8GHwgywD39OXX4ZbWqKGxNUuXWkxvhDpX
75v9iymCENCGcp/8qWBKmRUgEkfi9D9Ju08W2nh+KdXYpKOlMbwe8Y6DURY5k22+
ZjpU5/wOJmCKbbPIQr9i8ajebZBgZsjPq78DnhO+Fh35fVrpi2oDvy2BopWrDt4m
8EVWiqztXmLc53ZCmLj3p0H5m6im54s9FLXRtvGj+yB5EKvA0a+r9UVs8X0qwNWS
8Cb+IL0P2iU4ADOc05ziTImswNqNrZb+714fwBJ9UPY+9Ap8HWlJ8u+wYymmvUHk
qTi6dIpk+vSDP3JkN1OBa1fZOP572tX7nWNWANvqvddbqr3njaEydK8JUZ29P528
+wUnq4prq78bsnZ79ZeqQsVRDDDAeDBDEj6NmRrPpaWW6YjdHauGqS0DS8GrAdTd
ecS4+wBVQ7I3J+LljdaHyal7SrQXmCBUv6St6hE/kTD1zwDuV2CSGqKPwT8M36wv
Bfe7ZJ8A1C+bq1OHkk6tv3PsFAbZO+xtcU7SyXsx2D0m3b4hJKY48LeZR/liCDBE
cCCBVT+wpPtX47CuHLo1UeF55Oy0Zeu6nZude/I0gIk4ltXI+OMqUTtOQ0Kw+qST
Rk14Hb1DD3/88v3RF2YaURr9I3KC6QIJlxwzXv8jLmQVxZMNyABeKwQh/6v6GquW
Hyt9Ec8AtFQAAeqoDUb5+VDHO6JJEpNta2/BdfqHHIoWGVRpVMDlBuY3mflcgujA
VS/Dquvei8RtFZU5xQx8lLJgsHMM09xFO0sGtqsXDIxbaWU3s2NTC5XsDxeXZrhM
Kzw/2zIWUzYTYjv1nHW9UiMEdizfczJf/Y+m+0PPRqREtsu7trCWuuuKBKxv4r8j
uKy93+0mJr4hrQLEnfpEN2Mj7T2BXKj4ApDwNNOSoY6GOhbjf0tcPTEwTG5AiuQe
KYdkqqbSBw9yM9JN6v6QfV5gh9aTdAfLcszAMg3a7IUlhsnI/7QZvz3Hqs9rMzy/
e/FRg0lZ5NT9XwE2E7/o5x1PtDAAxN2Xng77o3a+7rBE0eIUBfrW7xNXM5o3TK+4
7ds9hluH5pTmiGDcz67XVBbBpCCAT2EMk5SvGeg5EZYKOwNGp6kym6LrCJM25m44
oJC5W0SwwL+tArq9oUVEEBjHiMe6qfUspgQI4IvcOKEFGFftIgj71RpTazCOsGEP
y/qnTbVEjmTbqDfgdyNSJmFbqzXeEQjKVjknJy5D1bFm1RpyWpaYqg09pYH0BrGV
Gcma7yaCuwIwpTlz2+1xlRSVMoJvUrdr77VriEu7YZthlnPgRtta96Rywfdww6ny
dJkYAQFlMMiGjpOibpsSE45tgD4Wavfqzz1T9HIB0VggxZuo10A5PdiG+HvIToG9
PzqLrhQklP3/mAU+X5cu8kSWGCGQxt+oM4gmJ3fbD5r5bE2lrCSQa/BPEyeatBeJ
cJt06pVbDdobwTv6gD9ITSYILn6LAFcUvFjTwM3+AID5C9pYGr91kZFzGfE+26pz
Ow3vrAdPEeBnFLZ3NzagwhP58yb2WE4rqTsrRevIfoiqjpnFliB9q/KIuRvStP6c
3DSWt1W4v73zUR5hTTHtXOY/cpryq5IbKg0S7zjuVSLIgfxeCHvYUNkI5cB61ZMO
N8I+TdKsI4bcvpNeVD6A/NnHoSU0MPYNBjvweWeeaUi0XPv8HvaengmGFerO9DlV
3jJCns2EXYlsRJ207jMNqZR4+vqdZU5jqVD4mNGU8UfwaDPuE23j6aGg1hHyLQB6
bGiZqWvVa7DIT0M6mIw0d8klauRUr5G4EGFjIqDBMRDf9MrbYX1GubtLBqFjSKh8
ekYSEZYMg6Ry2lCITllHRUA8Lw4OnUOhZnfjGKtUvR3Uz4zj5MamOyIsEquEolNB
wHFQrNm/k88I6ycXtS/iFZeREzgZHcpzxI17lAebIRyTfGXjOfYwfpdr8wq0rXlz
kgNlsjCzcG2dpXrH9+3Txl/JDS7CNuiVcdh+moDGt/73W/BeTOd6OuAgMNGs/0od
t2gmJx1qeYK2ZXNKcCObd9ZpU4afIoUDalvpb5Nn9O6nLO6lu6STLbzSgRTiuyfE
Fb0SvwmsY1wxi2YPYec6CzKEFqPG87VH/wWitTGZz8P3/33fGcaIZk3tBfG2m0YZ
TRj/VWMRkRnFV7D8CDPEEg1+3ubF5G4X0cUThC3H6N82WGpnx+9X70bQyA119piz
Pfcgy/nFs4plicZKTl/Jsa7yySQ5pzHVQxQT2O1dHtH1777MQ728JaMKtS6k1Y7m
JYsmb7n2vc13mRI/bMyKtV+havioBGLkaX/DwEDgxeYfJOIFcKJzh8m5R7aLdakA
CA2LDg8+3qKj82EMfu2wBNTyT03JQUc9Ri8pAv0p6XJEjWc572YxU+eoqpoE129t
ya9nV43tP2vzL4l59wxRWcv3s7Wf4BVjwJDe7AM4h4i40lb6sDO9b17hrWc/L+q1
DMPZpyHruDeBWm8ZX/Rr2CPw+BHOwgo3v8R06gzp+cvcjPVKdReMe9GHJ62eaL5L
UQ6c62pMm4CWhEeptTZxYj+xM0Etf4p4Xb2ZIKhf7b3CF3NgSALOA1Svb1kMSlg6
CJ0xEjeBFX1MClJMGRJAwXUrE4+ENiaPmaBbNzuhcFBoEqho4QI+QnI9Z0MAfn9c
EAO6pu/+mmvI5v0VsEK6g5JSS4Ho1UkMGZPDjVEi8LwpE5vxtH395QQJsQdYGlk/
sy6bZExFO9SMoihxHjfDTTXyfRSwEVBGI6jqEqCJSEyDTvyNkReJwxgjlKZL7yq5
JEnAV/aGXyWe2pHiNE8YWSx2yKdzdZsPnFkm+pkLOadtVdc1G7brZUhjgYkuOxrZ
DtjcP/xJfQJnHBQtscihqRbW9CcS8xh4GzYw8Jf8500X/dEcXqbji1PJ+uvckWvX
V7+y/YNrT6fsonQLwAmGMy0Fg1tFPoUmiw5qszFML+xt7+Z+W/0Hl3KlgkqY9hOb
8MALCyKtO8uA5w6pAbGWKHU9Vo7uFewgtlKCowE+nridmu7z+E0R7eg3XLaldDpY
UAlDmj/Ch5ZtXIqoqjq+eqZoYm4yEAcNOZJXRQUgZbQWOUXqHca8iR/d7sb6q/9I
2ro18vqLv10isyB60J6m8Yco869DliMs/HemfEv7TcQ2VcfezJcy+h58z7DkVjHO
4zBdryz1YaArQ5mYNPBB3912il1zBUUpO88LK41a3ann+bWJ28J3z4W+k6KhdEya
lfQ16/yV9rDiHcjmypE4D2gkbuN8ygw/HfNePgq7L1miF/tXAdBLizQn9766/7rL
SEjnnnSrTh1s68ynmMRiFOZTpmG4NEHMt2SinzdYNVpGUQb7eDZl+WvAsLo6Ds81
xW01InoAhHPkd3+8Qt9NpFPig/z6ZvaDElFMoOznQawlzgBYRlyQdVSZRZ6QC8GL
AQSZxs0hXex79etdrJnr5vGm/PDcNtUc6az0N6Soag2npErAbMbMd9O54UMkZxOZ
GolOQVftsbG/Dg+ExvaTAiBFEmKNzOhU6mgw/uHUII0oBKIHjlDkiSb43VxhRNSB
KHeSdyJh1JYyREOXqvAbHQwXaoN9IilZWMx+LJaMSmBGSNu4ve09ooLZFsU3AJhT
AkzCc792xjp/bpT5NzcTI5BM5jIeSMmikcg6+a/TzDjugHiVSEE+MPW1TBGbfOJ3
LVp2k+aUCD3YD5UHwSlzXE3lGW53ZRcVJRAsbrtfIIi8IxTRvk6k6bLQq/bS1MR9
0pY+tExRwUgsimmQOGx+42xUPTkFZbYlvPcyxIBH4tI2IGJpivnTfniOF3/f/BtP
GxlWLmUse2U3nMTpVUtzr7BK/vpKCeokp9EKKg6HUXrUeGTwTxcfHP91As9V8mVH
pzAKZkb29vZk0PV0KjV7UwPYO/JtYnokdyxAqcjqTAruGG8fDI1C7+y4DpwP01Wj
VjdzsciOnuLCUPaJ1u5nYuCxARqrEWENHBeP49bZU/cBknLQlGFLOHaJQYaZjw+F
+sZmhS4ZhB59VI4JwN5xKlLyYL5VzEyLNY3YNE9Sxj5yec1FOY0mbPxLa7i2zEY5
9KjEYtL4n5tIiZQXHMikhHlnvFOZBJSgsJ51r9r7yoiX9EH8Pd946u6doVSp6P+T
U3RROw03az1/W0hsBQosrAOOfbn47Q7lO6U3JnpVpSe3jQdP+dvC0LquUk626wxQ
QydTHT+5yPHE9FOlGjD+6eY9zHyxnI215LUNLWGiWkyP0p0WV8XkFkNtu1r0Frf8
t4qCZQa31IlmDk1rApom4bmWQ5zL7kNA7kEknxL4A5ssYBOqm078QrKu/U+TJso8
/08kKnPXaRi1VgUACocBtHylvpfZMvmnjlvyuKPcD5WWECN8Z2SeK9YCklOnohhj
GgK5oPMMRhXbtfCKx/NQGWFy4vH4C65l5TYTAn5oHySfwdTIlB+hYrVEp/fKzjEU
lv+Ho+GL6Npj6CRtM6hz09a249VeDzNKpcK0L8otgNjOCTNzUWBuam47RNKNXdXO
KCAR6Z9pb9Yk+xiUuqLrkQZYulhAul2X0lZo1dcm7p4dqvzQ1qjzt8u5wPTmJkM8
wrlttUAhrD0H6M49Awhx9AFeu6gR12cuR/DQi3qB6A/XL/8vRmFrSFjxVoJz1DbQ
/zEbWX9uZBWE2EUkcj9WGvLK2ISw4N7ZLMdD8+NiFiDy3pIy9hSDXo4m7xmGACnl
MFBMK7QjxL0oy0voXyyS47Ma/HqYQYES9yG5gnYClnI8d96MsGXTrDH25mMmHVkp
tJOxdQR5ntyXh7l1+ddd9d28aQFmcVMYius7Z2MzswPs1bQR4ubcf0ydFDPyhOLf
zrMUeKoagkYyRXOWd/TdQY8xX/FzRd+1IeuA/5WNn9npe5k8EmlNS7DWKoO1Fu41
SEpjEK6RI9zAPKt7gCcCGIa13m3B1/r+J8agNNJb1toHUsnENJ9wXlA4d2yAmUCf
IwuKAHs9GnvtwLY5F2UpHgMiIZNB8eUL/vYrSb4W4kijsuMf1AT96/W1Ur8qcSoS
hYXozNxW2+y145Yjax/tqg7JkK8jwzXdM7cEzqyFgAHPSM0KYHvZaCJ0h0UIdCiv
BEKBoiEPENyy3W9ziPSEKmuuL2Ah96lK8v5z36g9wjALUj4N4i6rIJJoB5x3AEuk
vzVo0uJn8M5vDtBoHgo+SfnHeu1N8UuCnTnuaosXH913mEbLj5b82QW7YH5woFa+
bm6+A7xps4uqWfQVAQQm2sXnyocYgaNHWLS3odpjId/KZqD26q1s6fXnN5zDmjBQ
QrITZ6ZCADFNGgPWGWDTFKbwBVq3aKJDC25AFAOvaWKiqeOxX1dxu5gSPf3f94uU
ytexG6mi9RfIbGmopBqDcQPbTfKQJhbFwbPzPDs6Zh4b2yuHEa7jLA5Uo1u/hG5+
PTR0APw31ldhsXG/099/s5/o+Zv5aWBeOa1a1U0R1RVuWG0y9nJfSQUlDRo7oCVL
AJ9YUM7Ia5pE7NLhqzj7dIhDTLUj/tfYcwpkAlDNSSvFkll+ujLAm2Sf4bAOqcYv
whJ46lx4c1bWxkLLF0bmDLWwuHqqOm4Fs1ihvLwwlH/39wj34XJZy27AeZRTzmRG
lYzU8Sc0wV8QfmAHX6Re38wLSbKgtZLPVzDubXw6Ybbm32aqRe5ELYIgcrP23BY6
HWYe+1OzumJGIVyK7iRc07z/9d5Kd1H7sqWIwQ38O6NDWL77ntWvBKLTfSXRPcQ3
hhrBTBpraJCPaIq0QQt4Hc94wQP7ue0/bNelfngKXlMEgXa5YGdoz3rU0gD5svHZ
IdPO1Yg/0bEWJWOjOJpjiKhlWQkVdf5vyGf3QAcXPfYfnvO7IWRDAOZMRhWTLv+M
VTFfJGsNpiBJbiV3DFIARsdgSJS70/j54dZK5/wOiBhT53nx7MMMBEB3cneJb85w
im0LOBynI5unQjQq1IUlhC9+3AJnYbHnF9LaJ04uN82YH4PYuwd+vNlD1/rQXow+
WCzuweLtnagNI1XJbndmh5QLk+c++BhtOAHGmpRKzU8ck3tyYLfTYMB851SihpwI
/3GhV0+yqJQaqMIew7I4pHBxzccbPnRehThs73Crin1suWOZsbxs9myslDcOFQ6Z
oXsw6qzstzzE1XJLpD953vdT9P+kjFBv1rGvSu0T1Gk8aHjsKhwvIkwPJhpgs97J
K22PnSgtYLqcsvWzbrOXA8WzYzF1+U+6ojOOVkdQvk2TEF12YzApYMZz6OtQnlW3
VsHmo/mDAAMZg20d8xYB2x73Gv3t7CRpDgq5HqZpI1ZEtwKqSqx4uadlElCLPdSy
w24hZ4xxbUK90qE8zRywnBrIwxEVGBTqUB36myvnXYK3Ib3FhHZ5wWUhv9mYJe8t
3MsyrnlvtuDzIQClrv/kfJXpFMMo3wdoK1D7aNUm2Ye5X+9OYj+ukTHoQ6a6iA2P
UcCiWAiHO2MpcmmtfK3e1cSDFjjoQD4P1NaKV/2HG3qrbPRzeCeZZMwGO1BeWXUK
NU6dKSWh9uSz5KSZ69NOw3UY0LaP0OcCRv3zve4M08EW9D29G6CK005eE+pSBO4A
jaG9v7EFQoXyNdMJ9kIum74E+WMg0QNNxTVod2yu/xWva1mgbBEnteae4Ro1/Fnb
+kmeOO0GKlGylH7VaAO2bPYTXJBYpIqZo0R2hgOcktnC/XRHxMltJQuBHpbGKHpw
Z4zo5VjF7Bm+iqX7A/RtYLZVPPAdAfj4VR/P6wR/yF4UxhIidjmdjIw2VwYZnGFT
Se74u6Ht4bJNeCJx4L2mZk+Bb1Rt8HeRdhk1hb4YUMiiVUnJpCjOOv0hqgNQ1Mjs
YNsWu2ZbS7sKKWW9bR6KDunEY65tY0Gf6vj8ztlpzT4QXXxpNLsx0HGBTsqJRzif
NZml+JDtzLgbvtCxG7jp+IRRjoMHNB3I/MVXodFNJ+QvmTOUuRYETSLYOjcFTlld
sNS0I37duvg98d1Rh/2HwBXX+P5yoewTQ9Ly8be96Hoetra2KLviLhvDAQ6Vs/8s
bSWxGaDkuhO8/ThqURrOMu48h9oa7JDoheoUheWFt/JwwpeItizqxuosFRagB7h3
OnI00LpzbeG8kF9L7D9/67tYfcri7kNQtMz86VLJPkikBMx7kcalLgVVIq5DWVul
CwzrEP0refjljWZA7UKfDlajwAlExg2NGRwD1BeOoPF2YQOw5j20VvI4i8gOzBG7
MbR5cQlQxE7P3FyWGZ85jXK+gRZFtzX9wdl7tKCMD8I4OhLiTryzVdJGSTGw//wU
DB0ObICIwYj0xsBExyeSSTjla4j9bXHYJTLAiDqtA2NY3uijo+DLLlr4QGDgec58
4I9uV6a4NnKnVI9hYnBH4lF39O436qE9BvZ7id/LUPhEb12PvT0v8DJKd2y032aZ
9Kl1UkAt1oVnw5cjD50Pggeb0RJubdeXpxLm40kCKM7Lo/njX4lPdKlpRw3BBGIa
9DZLDDNShSe6+GtXiS6ALOloTEOLBExzRO0yr4JmqX0r/64vKjJOr5xD6htZSur0
anTK2CjxOD1ki/hM4ztGwwWbzLkOySa9PVPdTOQHuJJ0Pv321aazXTbBV7VLpfKj
8BZqhK2Q8pyiepx1j4zWiuSwJtPnEKhcculD2cfrWuxDoXlyIUBcJCECIM4UUv6f
2mBG3M6qC6oXyuJRlwpU8RvJvEuaKCJ6Uhf1Dzbt/KO6BB8XitD51EiB26aRKaQG
YdedJfHFFjEeKFfCF6jjjXraSIMsrtIQ9cU5T1gJggvespui0fZaB0/fRtq11v4h
ihlYVHnHY3tNN9i6pVdNjX0fcGLyVGzZhCDefM/pGoGU/wvD0TzeqUN/KOXB1tRB
rgcRoBiPKkAeUUqlY/10oBwtYLimzv23INoW5WdAOyJdXT1AAv14J5G9lwBRFw6Y
yf/pofS0t21qHyOXdYzU1LrLpc0j7wIoXR+V/LdqxNicdNTvnDudm1gVibQj//Zk
8ri9f5GGyr6MqqKBjSHettl9rK/oxmjtrvAilY/qzmea9XQCDmF8a8RnkAPDSK/h
Vw6I/1HMk1KKmelHXm9mzA98fXcW4e4qY8tCEDpLPz4YfTmTgGo4LEoAc6v3nryb
9+qlxrmNkWoSHLSp5j52UMlJ8NBR1cv+2dQ8eKp1bzZ6SxQcrru/pgUYXBFA8p1q
pl6L1Hl6dJMuxGZXdeuwdAD0Eim3KfoFuC4jOsN5wSB6BGd7+zIjSWY5itYHymIn
017645sFLl3uxPk4yFxxWRc9UQDtmipEPD6XCgk1y3HgVpyPfmsZlq1H/x1ot1Rc
HsTrGvHLxw2UH/p4J+7fvWpFrSTL0L0Jy/bfqYO27/E0BuVsP0zXSpDwDofZkJ7t
OHbbgwlLeR6AXfJ2Ndg5fSYv3mzNaN8ViJ9eqBxe/OA8NPNy0wlOZW1Wogkqfgzk
2W7gVVtAxIpWjT84Gnq7m622q3WdPOjn4nwQF2+vG8X7V+GS8P+cAZvJ76uzuTAf
RwffjlhhD4k4a/gd/8muWWmUBflseMDu2xVfBz00hQCXIFxgSoboY4ZqyMFYIyqL
ga8UcGwr8C8ZFp0vo3+RDFeXs7W3roNqnsgpm6NwVh2LNWF07ob0f7Bn34Iw/y0w
HLdRc9vW/GBZdPcEkcOHag+2K/gnQ3nHqdz61KrsRaFmBCTIgPyRjuyf8hd11PI1
l6hsc2nJ6nagApp9RpGvHQqpaAggiY/gKUJHvnGAntTIypT4BtE/pReQiqRnnj1v
Cb1aZM0/Pdp5kgOAK6F9CDhq3FwIIj5Ipf6qSKprlm+sT8aaIoCul8s//WketF9i
guME8OfbgeO7NgD/iGupgO6xfdyceddQ99YGB6P7EXgGkfhTgE4ZSuunO8i/MeVD
DCNCP/iYEcnLs2aroAnCSZ7IfKyU31Clf+Ynk63+UHSnEcK2wdFSkRtuSHmiQ+9t
A7m+lXQ1h+154mkdjF28290eTjSQK5+OVHdh2x9m5dNI8zz7fn3EU+aaYw46CmyU
jB1dTVWjEkazb0j3aPHEr40Afda2cCqHKyfa7f5wBAJ0/vkL1sjvLzWFXKJj1+s8
rIOG50WZbQUJRYig3mP1dDKnUzoX7+Zg51bFVc+/HAPgbFo+MKYcPPo26Ctvctgx
U97l3Q+m/T/of8oxoFcOXG0cIwVVDYoZPPJk8ZPPuv9LJXxhRV7tZtUl1p7eBGH4
DLlGStuyeoUBGqiXebMwbEPBpNSoa3kDwq8gskD0kyDE4KUNedFkD5GyXNkLH62M
4pnI4Nc0f3Fw3DhTLtiLumkQ8MKJqbjV4cUtkB2DoUy011sAVKciMRTicB5eXGF/
JyYh+N9opI4LYM0pKBruofpL8Cu02aebZJG7Bvbnfov8UvqwIN51xEwp8gH/zLkp
2BLFDmDR+BQAxJHzQ7QLD1SruXt8darLWFf427EoULzL1IcIhCfF6nbeMH64qUI2
K6CQjphFNnZcqmH0z6cuUtqbH9Q/yGkYjVGzDt9Jt5kbaLKqujdHIhK/5KoGT3Vg
vyjDLim+uXC68zovCi+d0/LfjAQhVAAYJ/fLnL6CRfdGlYZnVHaPO2qgheNH/tKt
lANN3Jk+eBUEIC2FDNH1rrG7TVPIkEAEkOz3yMwVZY2Dgu6/eTo/vy+BnorSunq8
HTWtSsA6Umcl3icYFcgyFrMbKlr9WHeGGzg1AO7xchkcj7ZN6W6QYSkf0FSFDkuU
Rhe855Wf3jqg1ySbnYOx7y7qoty2sZNUOrg7n4r3yJ7G3GMdUZZYT7oBZxLYhRow
Gqy5i2uouwz+5meL1xPiTI3q/Ozmt+lhVTFFf5eeZt98c0ZtTO6Gu66+BTGr0xku
a4S82xiVnuM3XktbrRTldO9y2ivoQL3ohiVY8KQHFjsuNABj0YkfS49ay6v1/rUQ
DLw6tF+Il6aeT6hgWGFxSqe23A79NpLdIqLayNEFjYpoSyRPHuGiPl6Zf1MofPEK
mgpGGc5u7WLVYYns0vyBo4vcf7TT+o7D/DE3KFbRrP2mKJSLr2TeMJJXshEDFU1s
FhuuidAp7I+0TyTT+A5f7qK3RNlUIJSSt7YhHcepMj0u/nzKS8E1GGV7pNBsNC4u
+N8S9AWFfEu36LBIewsbfx5f68W4qFnZksTVFH8nwTOwCcjkO2LeUt06P0+Urfzm
R3dFDvogj3zxikQzUE5LtWarHPV7CW9mFOkD2IsPT3VMGl7fa8rIZ8w3SAoNRTF6
rPsG3aJzHlZ+5aepZynYPKHQ54oMBgmKxnCDn6Ywe4T1ISTor9xgHJgP34OHadQI
AsiIyxrMR+J8nfZ/fnHQyizCJlAS+zlr+YJubwGLvLJ/6eVSQCYT1QvCiIbUUwAh
LWwSbMajFh7vbN/hBOcLpYuRLz5AXVuL+2GaymiO1SKEie2QDArArAQv1irSPOU3
9W53+Jgo/jjU2ryOK4VMw2Z3zjDnbIkSBRPUoxp9V2CjthutQtdIxwhcAuAUt92l
TPfAKcp4xjHvRaqekXmKEulIuKAq1F8bBqEMHjaU4Y8B9WV95DaNRmDjeIqkUyyB
KmSUD3o5ryV6H2XdZs/vTmVhDD4EZapz4HPx64JERMP0LOrjWD5kmLxD+50BKaUa
3EO6tkpREi2vUOSv1LHpgFK5seTE+4lyz03+kN3o748bS7DFp8pbs3qjvCsw4oJm
PuIfJTrE2wbd8J9HcEoC2fo3sHebqSXstAizkG+HW3TVOLizcGZMv7bqNszGN12c
jsG+LWKR/oSJwgYq85+3HsgLs64Tfyx+3vgfLuOP+yISQyBbW3DBHqcaeIxrGnYT
Go9wumJHfxqDmqlEySIuL20ywX6fi02hN2RJXMiuGAbFYULup613+SO10lblfoUD
EkYR4gIbxCaUUt1DzfVNBYJwcYiMammYvELYAcVXsF+Iw4fTcONs+JcTy/HDswWK
0wkvwkGHFIklCqKGgFHnLEWMRFu3+Sp8XYkTB8J4c0sNPG3MC6PyKPw8vxkDCN7L
HYaYLItV3VCopQVgKQldx6a/veX6QSG9utOAboHKsFEmk/P/h+nY9vaRboN2Y0hW
LnOUz4/RE4nu9N11fsiFfuqiZIQZ85HlbcOknIAiQfarrgNE9tjoMgceU+PItm4q
giJKpNbaHVGEpOFkwJqqDQ5YOZZD0S+XNdmuCaDBFcfI5fBSNtTRULMK6JmIU/iR
52WjOD6l/vgCqhIFCvJFo2Pccq7yBjeVykTXD8O/WBY0ptyJNcjQQA2O3VFi2mdy
yjY4oMG7XLQ3uX8+Wd4FaG75Cb5+EUeCKQbHmV4XTWDoFMd9xXjiKZywdNSxhcoZ
29TEKYo5+C4nirsUDOxVY2GLWwY8PB1BT51amWjU2vm5qOsg+sF10tjW9W9uvy4l
/JxCecnK9Qb/CwU5B6lnZnb1m6GgPlJ69LwMPqJKuNmE6Xq+lhCGnkckvpRqhL0H
FAc5RpKTsJf5WzRLYWey3C9UaYb3fT2LZ/VVmpJHcfUzOwjQ4hy2hbwWiMGQ1+gu
88QvyuOFuoHqYR9jURuS/XpJ0iPpi1m37nCa9rhpPksF+/7hFiNHNMYaZ59REntM
vUCLH8kAroVr878Udfcx7bkQpOWNOEW2ONZT3glokuMxsVc+EBANpm/a9rKYYRks
g/UP703zXXcUhMee1eWMOcs4tfX87uu4JDCVsWI94/vy1aRda1qkJgRkrMCQU3xM
yMywECt3OFRrVL5ciHlJPBapZmCEeMdL59JwQxBX4ZNQGV+OP0KA4kMEjzTy1NAx
7r5PMk6vyKrLv/xYPaVwK11lg5kU118lH6fmziIGumnoRBPTjsAYXMvFAIRmaTUD
8GNyxxYRWBPK3R1PfQqgNtiJ53wjRdQh7Oh5je3AvvxNDeOitMa5GKcwXwqx1PwZ
7MEbAGnDZqUG5tWYYtmeOJooHNzD/dB4WLVPGH4y3fxuUlUi1d8LEMncH8MecFLs
8CKutw0fZ9hONKrqzceghhE9pGLPckyqZQjWXiptkICiiUOHYf1ndmIT+BjCEfoB
saLygsQCBbGRm5nF4NDfSit3+zHH7PNySn/Hmf6m3Gugg5vaN9tIRNAIboS4YrZ/
APZ0Hsi737hgqwkej+Pq1sNVSe8jDMdZIkejYYuul9KaXy/tt3sznMzpM8X70dtg
44rwSerjsQituBBbERXmcwDdJqv+YLzFM0w5qZEZKO5ghavwdOAOhe7NZOaZbhA1
rOIJDHwH/+yjkjQwFZb3BiFIivkm9uTUvZa0EJtHzk3i5Cow601glMNZl7lTGObb
TY1PuGU5xgIaGk/aQzIAZl5bUU3Jr01wSv6b7yBIKqct1PHdHj9878V1K0Ed+3by
Ub7DpC4ZEaB88rOL94sYsgMNuyg2rxgw52y1od02rIfKtx2iC9/2LyXebiZPVVHh
VdNkPMFgYGsLQ42w9iDfRTlT7DOi+peu5QD3hmFs0U9wCWF+0/xQ+VyjEE1EEOti
F1aH98xH1+i2AA7eIe3rHDV+Ni9rqVIoz6OTLZKlIqBzC2Tg3GhG2PVab4MkbAML
2YPSYIF8YV5cSMOWq+pgOvQzVOHulbprdu22RH+hOm1cO5Ge1UzK4ED1AnGq9G6d
WRLlBLskkyMJHr3dVtiO4eAOEzwYgk6QiGUu0IYA+8t+sIOkcT9tmRE7dFfA8LxO
9dhCK7PuEMPp8g0RnZxBP33F5qRJe5+F79vq3VzmwRGdk24MQ5IZN991H957yPTc
2TFLoC49IGpukSICeBV8U5dZ3faFEJtVIsIVdFtrlhZC7O8ev5AC8yrpthJ3qc9/
obRXK33tFxdGij58jUZM9HX9lBOjp5qhKnp50sn4gCPMyRAgRpFgx6KfemjkyWpI
SO9Mex52GWD8tpMJDNmhrY/ZFNHvc4jI29IuGf1vxEK90M3DnZOAIaFEzQcW04xe
8fNzXQum3Pp+i5DjB6ll2YwrowwghDZS1Upj9x3hwKk8FUWoJOOAmQPSSy3/0WmL
/AOBhBUf7cSXNK5hwQLvbIjDsNXbVUaCKnaesN3NAUjZmaR1tdwQOO5iqu0+Tgjq
4gAV4TcfOLr9ZuK5iIfODNEkLIxSUuzz6N8EygYpOvqYiyg4waNzbXmm7sltLeaX
WP6cj7r7F/+xkjkVpDyDDQI7ty7yuQq6Jmih/hTBAbzf5c7VeNs04TY9T/CQFuGd
n8lG23PP5qZ0Z0DULLQeJd/zbWxQi6UzB+qh0qTy4USSx7F0uy9Bs+/d9iR/lB/w
Yb5pVTWdZqyYzar4NT+fjNX2tLb7p8GlV3vEOyU/sArh4SxB7joAbo/vU0OpsU4q
ZFjup+zpApbp+Tcgpx5yYmg03tHP/yCzA3z51Bp22xvf96g4Df8M7mctY2+kJ9wr
wDEqhkewGqWgRVUJKKZU9wH9GGAYkcDuAaGvBRPIc0sylpF9maWepYnouD1uRbRV
qZfqa7ioze18eSTty40ELEj/FG7esjZHZtVx2gHt2zvidfe9r3vUczdxXZh0rm0p
bG55WVmL0spqkhppCA/CydlRLmqlbOV0zj+2CyiT9lvyND0Qo4Gtd9Gw4RiDKXJJ
xwiYCFF3lb5R5IVT/YImPKhsWtRQYJ2q+9zA7KUUGhHAn+kXphElfiYKEj8bgYEC
R3H6NdNsnGN8fOL+FKaC3mnl9G/kXI6kndYUXicoQS50ssDAnSByqSpHwfPNWEL9
bgRbXo8qD5nNgFYt3Mh+0BC1zoCB6EP9GciZmyijUG/QeTHE+93qlWgXabGnO5cC
xIMDvX/E953GQ3pUXl8Q2LuJahpO2Zol1EzPfsyymXa8kQHtH86erfgp34OgwlxJ
5Rg5oS1v+Mbld2b177Ln2L8XQkvPjhTAdI/0pPsbLPB4l/gITVdwjUqwIpsRRt49
2tn99WAzr9h+T9jkZqBSxgPg2NqGhzfBZu9gL6Qzgk/Uxzc0w6rCJUCoSGmw3U8d
BedG+cpXhtqc9i2yDOvQ4BBBRqBTEIpuC38BdGCV6Acox94876kRHhnKs2x1NLV2
vxwBAK3L6JZbHpkInS43rf78ILa91wG4BPYsXUWJiW3DosiG2+UavNELxDqDTTm+
FgX74HTDHk0j0YJgCBbonN5VLI/kNeObYEaVOV0LOTmPKyCGcq4OyQ+FRM1f1ziI
danhX9vy8xg/wBEE2XKccIo9BANqAFm8bJZdRItjl02YXB8I932SsJ97w3THvIyt
EyePv/Lv+fIpMGkHw/VlZcQNDuBiu8GHbNPLrkQy3WMLt/VHBB2KAB8jVbMe+5dy
6/waN6Lm+tcC9DWKmPGz3d5AfHZCFGwgnjEyD3omWIKscIe8bPobHVo2oDY4UZFn
7E97FamO3y5hoCdi8Ir/GLoaPGwwHG6WGmAweowEKP4LqlCfdgRa8xWaYW+2nkd3
XFR0651HDmqJphdx0bSKXxspVBJBxSfF3gUAxWhX7VA6yYLO10Qtn3su2ZZN0VMP
65erfdL1/MsMIH1MdkYa5T6J3ASB5RazZOYi1zMwqci/U1575MOIi77QNGpsJmOQ
Ifs7wFR2ns+TG465Z8l2w8p4kbuCJB5skeJsJXnJFJ4zpO8/7cVo7OFB2Xrwx9UR
rj7quTr0qc3h4HGhvqad91QKjnHruWYDSDwqiQUlYhJgr0WiqTYI9FDqqI2CzlTy
mZox6RBHUVwfgdLiEvvZ0S5gYjmanox5J9lgGLAVs1GY1o/UOETyeDmHGR0bBLez
/WbRNgjP8q53PaHT0vLegfkkkCJOkfsJOJeQT0qZupMaR+uRHpT4MhfuX79At9ld
FkBTyGAfqtdxQr1mKHZIsUHwtsPyuhH1q3uFc7IjgwdoKIHIInvv1pT9i1tJoYjf
zcIEA3Jo7kWBG0UTwF7u4bBpFY2WnelZjVypd8QJg5ZRxPvkZNOIWTf93wfx/9/4
2OUlsP4kFkmE4tILIuzh1mxZTSYA7w4PfgEA2QRxR/sK80hhLq+5NZNJN+BXC4ZI
v2VGBDQOiECqo1RklFrugp2Er8LrqB2/iCbZa/ZUtNuzxGzN8Gbzcf6zCW4T02YM
vJdRV5En7Lj8IRvlo5j7evcd4ZEmfOctWBckNgsRkm+Tj5S8Piu+nTmf5cQRmzVD
yjynjhitptAEjkq1xCiG/jS2mSDho5pxoM4AgMmqs92R3+1xMQy3eMaKmkzwcYS4
ejTLxaP0GR09VmTJz+22WQQA6YeyVj2zbabTXF9GCEGR8dGTAp4zpC2bXtAWBVdg
rPwyIbieX2c274Q0pBN/j9sLM7jgVJWrdq6f9WxyhIBSmBm8Hodu8vwfTzB9oQR3
9yPaKLNOvcVZR3HMrvMD7Hqt9yHYJeq3RmCc6umu0LNgPQHk92GsYpEAMaWzxQyQ
ZfLL1bkyEj7MoL9L8crmS/ZhXrtGZGq5P0+doBNxKMQWJCTPqqk1kdObBrZXEYW7
nxfCpmUl8rI/ibHZJN52fHsec1qrGbr/5GcKqSSVuQ0DIGPKRhqNhx1JzXbzX8Vu
ztS88/fVZ4L6OOxI6cFbit2dmhQmiZ1eaGCr8exzjaXjEbzensb6ICuorbhEwXcN
g2Pv17bdGihWgvf43DMMdq3Yx+7yveSJjvqmFgwVIsqyTXis0Jd2TNoK0u1NaRSr
kd/1RoF83jsA8lGHTNTu0JOzMtuWm084t9O89X0PD+SY1Bh3Tdv8ac0jVc4KSSxv
QpLztvcozBTf1DYkuVtT5gh0WQ7BZAD3FjysHEOpCRIN29SaRmNN2goz4+bSOqsk
ZzLEuWjH1hBIVgj/D5aDFk19B+xj5wihAvjyXs6tVttBaFNGm/tIVsucIbgKt6UQ
lKzCSZeUcty8UwjAZyqYUZJq5zNDxbg5jpzaupHVTIBY9VZC71n05+qcRR9sVY/N
PaqQGfTNVzzomdlK9YdUtuzAe68qEmZU8JlUHDsZ33KGL97dfAk2eSSjIBfJWI8s
5cOynY0VuI9AG3v2eB3se0Ezj1Er7E/r4tvBREj11uLJgTfk2HVJj/ktnTnYciG8
R6CIJPOA/Jph3RJRJHy2By+0/5c4lcSOgfP3ekGgdGk4WKEzlc6/rSPZbS88oETb
MSXpL3rN6qFL9zTRrqxdvpO8AuT12BfTxPED8p3Ob+QcPU+94uFEV/YqeFXBwamV
GkWgKrun+zSI6sqTRkshsntfI5SRNw/PSRU3KVA+m1LMcwq+foiQyi0+Pe62WcAj
QSdplxYE+YGK2UnSRqX6g9pjCCmymNE57N7k47mXX7G/ptBaC7xm4wzMz7lW+kCJ
XbvMpWyw1DExCV6bxSAFGdDaxU8GTl6WD0z6FONx2bm+o7N2JKVMpfk4xnw4mv72
WPMrgxr5D6ypgyjxZGIIoAYHL2iTsF/E8vmweRLx5PZeXb+A/XuEE/tTd9Apcgcc
tk2gb93JMEss1DOQGj1GKvOOldPvvE+bwFfO1SaqZg4+pngNPnsz1ybxTqUgnUlq
cSBrw8JdcrieMEUqmj1vYJY4x8xJH3f9j/MFW7RfBbXaZ7g2FoUpconryL1JLzkc
yUfMgmVHqb8uXW0FHMWNprK0zYMWBoMgEEBsouRwzOQmC01k5tiDRNtjmM62ZvwQ
MEjH/sBtuFjoKEbrWhwksAjk3noZjqesdSBGBnOmiJjKAHm882ZQmVmDSTUIBaDU
dsqr3KZ02ImwdL1LqkRuiz2VDiT43Kn47WROLHZD9o5vc36osxlzfRjL0ie7Fl+L
p5Cd5/xezyLm7OEn+JbAl0iBG1g18Yk4Xmx+GAtwNotLnXdjkuiC8SXimDNvfzfE
HUs839ODFoRVOvpfIcJHHm6NMCEgbYb7pFebffhefVbUoQQHFzeqO1ts+dajJq5A
bho3clWD07EuH0sX8U0Asp2IT+TgAxhGYTFGTVSRIAWCiC2VqxMjhXcjZ18ufjUW
2iVjQkkF64LtGzVjtpjcFlH2459oUqA/UR11zOtjabFyBd9JZ8hREcLFbwogj793
rc/KJMHEyB9qahljl2cMoV5c9W5EBqloMr1Iw62PngrPYLOeIJZaS1FRSYV+hUo0
B9Os1ZNNoojgPDdjnnEMU/A5iG5WjvynDURd17zXvEprywynfg1PKTqOhm1hMlcg
op63J0f2bma7IuUlIQGSBhCZ3CYHbXiT8MM3qcZ+qNtevPfJIK/qE2eL76AizxJ+
ZvQcWDhH6xyVD+m5S90m6qpk8depjuChTh6PIiNWeTftbCuhK7PEE2pZvP54oAjM
Ba/2FANOU8s/b/9rEYPuywHjY2RSDcMpcMNCcqWXptR6Tfk/6bp2T+xClyCcQEe7
ugynh4VT3BCaOvPG+dNcBc2byS8zQtgiHfS72RQhHTAVMp4cP5JK4Yef2hRJJiY7
SE0m0LCtveQV2LbXUVDGiKhf2/h87WpQkhVhPzahrKezvPYOH67MnQZ+lBkbxPf9
Z0uVpOgityLPTqGblKSp6QEh5Q9xbnBvnsXCsoDhALC5V3vFlmvUaWNM1+txTGEt
LjnnuwszTAFepqimY3J3OWYkbeh1TpgKncpJfCyNMzKF45PkzcZhsGZQeAn5Fs3R
SChvHHxCK/J9hufGYiQzPCCG/XAQcCN24wc1k0CXexuBp96EphmjGsXJSAJWtjUg
22PbfeyzvGvkyzCED2/CwsZFMK0H3MUn2r8pMhG+aieUpRcmFzlJdrYhiG4TuGyc
zxz+XoOwgQHTQwi4m3pRSeVS4f98AfVzVrZIL+fhu8b4hhPXN7nb+7LReOAXJ4gc
j1LLxJowIz1I1GDiW6j4VPu+JpZDoejq/fR1Pplzg/ZPK4K1SuqwVrlwvht2+m6J
w1VyFrfiuB9WlMxSAqKjnsawltiHXa+Ij4iyS1w6kNy8AH5zIPcgKv4cQTHze6qW
0NVsp1nbLfcflGZyTo+nw1pkhSBzvbv+j1AzzZtAlZN/mU8f2oNGmh9qL23lC9oj
4NAGBvEzwn0AqzMTkwxwQehXowWwDqMLBbzw1dFQAechYSoZeizF8EvEA+yvxRpR
cwpEky1heMhybPUvIE/BHOpwFqv4mWmzpyXbHs8l+7u5ArYUZzy2JuUTR0DI3pGR
lwSRixYvG7IjbDRLnqfKPseSDaihuQFuvbx33zNNxwQO48LzYLdb8PGnUIIXGQac
kLqQENkkr29GmbKVT2w8ImkzSiwEymuu3PmFdZQWd1GScocYv3qxD/cqx796iebR
zBiWkg3I+RRBoDFNSdB2YGHrHQoqOdNOA7gNl9mlnIQMzdoctTWXq0fuskuwCBH3
YeengvdMl/wkiU/oFHz1enP/ECRNBJhwqmphvsaPUj0xH0vi1pwYDP//R9TxXMt5
jRBLlnMstdP0N8fSd5Kb2wuU4dv/8B6HcVWQcJLltsrMG8n2z9o1iMXODrpjnh7o
c1/U5u0O10mnXDlrkKkG0hHLjSTbT4A44q15a3t2aJvMawN+arvS+doTL/7hSSV3
OXN+prJ3fE1I/WLXC0tUij/ueOVhK9UH25BxZDxAZeQ5IV/YxSdRbU4wIx+d4Dhz
2pJpJuJ8DunLOVw0Az7DoHkieGAnnI3VzWyS2JuJI59GJh4DCwxh7i2AL4pJ0boY
Vs6OWLOWrMY5A9JqyYe9xq5wpCZKZzArb8FLP3yyNOVuL4samyuA7jM5R5ktBUQH
0kqCfHjPj4JUXSPY1BlDAg6WJdAZQWxO4by8OkbmAOW5q96vjOx8IDqxmGhRWjHA
13cM0W4U3fNwWkZOvnojMTWdInT2VUxJdO7eeiPQh3YxiqZ/M4qP0w42avTfSsfA
ZTqpdTFeDZkHQORETfUfP2FB3U1gTjv/AFYqa9ACynsNwi92XJVQk1WHIrdkh+ga
BZ7PTqh5UGpclXNxh8tAg2yeZkAtxth/pUXBaPRqKmosoiPpnVsqM8Hy1c7fkD8M
HuuE79KJVaAKhbrh9H/rp4X/wIb6EX9Hhk286pSoU0OLDtWPQn/pQtiIEaaC8AfB
Rpbqlfc/4HNoSxUv5oK57a00yiiZz10qOxp2znqxky6+yigbhIpnjyFIEGgaXJKz
/bvkYxZ5lfMQ7ZRLr0NBH44UvDqk1ZH+vuTiQo1z4LBlKnUSOSpm0yNbwtIfVYnr
U6g/0x50USc2b+C9J04DYc4tcF+ehV6hUlW5DU6s14hOVhgI6G8T4rGlKtEfW2t7
bq0ZsIlO6JXmhmsOguhEUPsKAHQpXJRCeoPeqIs8mHfe0ec4ea7ffqti1pSfWVWd
a32Us/+TEz9bWGO1tjt6VaTXeQv9a+XTtOIYzkuqcl+9Ij1W9KU5Z/J11FqOneSE
JfQ3L778ZXmMu7jDl6nmZCdYB2BstptNo6ADNxd0IwiPUUqAvAw2Ml1BaaA3RO8C
VDf5UPCLxGHl/1hEUEV8mEk6Rf0lf7f/1Rheip+VKDIcgZi2b/1dx19AXcW7DQOp
v2SAVbfHlI+yTfP7uiOWJZ3FvtQMVLdE3fT5tvYv5t7Q5EADdXbXbdgwlNBbCduh
xMe6z9a5XoO3ODhptN+TdJlidPYEpeImJhuyUPL8OSM940l263sikMBVJmwNGfRr
jfjCJSnInoqY3kTHuHCO5cyEJlH+teho7y3bJxnjxaV04jeTSNaRNSrx7fb5xn0t
c9uxOYkIclyjKmipaFmi0ApSJO1jUTc9cKH46Skao8V8EOAe8eSHrGcJm0/AYnji
gFIUQPAz/89d5KkKZCjY/b5OXE5WIUXH8VXfpB3eQSTIP96bHFMNkAfOl6BQWX8U
lwpombXlHbmc3S1ZrjA1V4LKcMqkYcPw264t9wP7UOFgkHzB7X1TZOU0Y2ibtvcx
qM6flxWyWrVN2mKJXtzBHd1q0lkx6o2QxujBlIdwHfcf2pmx3kqs8V2fEKMXliU7
j7xvhiAeMhROvIOtBaF2mqBYqUNksTtn5ACaITGppZ8Ju4FEXJoOh5yxQLD0GySi
TgFd/2+HUiqHSfApLJpdlSf04V8FrEj+fJzCrrHnu31wBu3yO7lZH1Ik5wEJ/ROn
rJlG/GJRoMol9CASpF8NHEISmbfx/hG62vg2WgThuKr+OXWYBBIUKpdEoKQaZXsW
+VoXSVX+DYY9sbBj8JdkL0LjXGf04U4iYYqZQTriXmQJIyF4+Yec6AYsvL93t+/Y
L52a350sw/9jx6Qy1mL0LcUX8+g+Rg7n2H32tiONqgqqbeeP47RSIQDhp41OwruK
wJ5dmCMBYME8Dsc/kfo5ADPqNk6rl38/Y/XQ3nKcurQ5pWzwSAdkdBjQ7gqMh4u2
BKx6b4ZtZHRW0eox/oMWjMz5G0Sf96n2YRgaBcbT0tQ+DgYXaH/FeZEDK1IkEHfe
/rGxrhrTSB33BhgzaBVnulxl1S8ahrTGjSrv+a/ETtfyrQDgleI8DSNdqFnwTQSS
LbjaETzgWvK8EeoW/4zLdzf1LAvePZwqvLL34vBfkMnK91RZjhW1zOwjwSOFJJ8u
tm5ob9Vq0U/0ok3qzoKGD2+Sx/1ULh8eAHwJkNKCcvL4irQwBth7FZqBXpzGEeUO
dlzkEgvTd7the+8brzfbfV9gDhyNhHqwxUrU1mOksi71BYaPvH/KitqOaUbe6R0w
A0D7eLB1INodCaSgeXB8/m7H8tO4/rbM+HUAlPZLMJm5XqPOeIx05UwzKIJpmmlc
7/FRbewGVoKBj6OJhNt0oh5Z1Al+yFX6Kh3mL9T1AHrtx+znqzUS0plcmCLzfP89
V8IyQ52QSpscTLsQEURVbt4/hf3ekfTIugM22DIVDvI0fDWQClPsv7RarpzESfUk
e02I8WB37GC0Q3BjocsrxbwpuAAsv778BwZL4MK9nZNTZ3nqzUrKSSAyvcca4qKf
//l1xve90G07dQ8cWBdV907cp/lySQGtUqHD/mWY+C2lgdh3r/a6UGhY1U/2J28O
HtaITp7PKS5T/YPy9/Qd4f1RO8lvWmjo+7fsdokRe2gEuVfVDHBeK3h2y6UMMi6R
KpXIXPHhPoz/FrnbCyGIhWFsuHd6PqCBb2WCATFUPJjf3pp+z2/dtSDTbCjx+DOQ
IMwHvPf7dAPjqcl8Edltu3L41zeman/EIbKUO1MWOmXdQ9G4abZ7JkyBFl1oLpJL
LQzRg6bkpgH5vGlnK8E6FSLoD+i/qIkJaXfWF759rW48m9ctGhiu32gHsVSLBLrn
UbKKgHDYU5cTcVMITnF5dxJR9v8TVYd0XxerMxzc+hAuabZd5wloLB2zVeQxBXGQ
QOmg/32YEZTC11b2BqM94dVMhJwBGhKZ6I92tfMpWIJ2wSYPdCk1i2li15iRZxGf
cgMSI+Zah7UTyhEaJoYPulPJ6YmC5JdVt0cn6wMUWZ/bSKaxGt3ag9HZ6kmv9Qyt
Ph9DFvTOWdvRJIWMQDcegolIYnjkLdDx/IguS5SUztjU1+0q/6/eeDqOihGJrfJy
QbyiIdIqi3jZnkNWrQe5xZwT2CVSVNTlgtcYv1+ARMr4gV55pWIOdhtvCRb+erfU
ybTlXP4+7OCXFKkPFrdFvi7PUsmIjVqNder1gUzIswCUJUN11LTkhkJTr30ojfay
hhk3Q55M5nGgEE5PBqiV35un6vK+fPhc0vsfJvP3EJSaI31XJTSAsQgO1tap/pq/
w8POZu04XFiVBAwIPHJLoSIETxOurBJsiY8ZubdjzG640IFw/2t5sE0EHgZxDGLM
bi48rbGwmzenmXBZuMWFaWOqUmkb0J1THi1ZUpI3dERI7kEWqGPXuEP0/eQCCfeZ
lAJtHTCBvIm19KbAHIpZdTM5Pm4MpruNvveSoJqBsThOeOlJUWg2fa2R/dFlDNSy
4MuG0fg9JmMjwTlgT5ENmTXoXfIpV8EztZXniZl168Y6xhIl0EgGj+79gWjKiVZS
YALmApG71Vzm5BSoU424BRvLZTHSDlgmahwirT5uDB4raMphGhBej3OYpWNzNVmD
TBW2SfBz+hRCwCJUcnjTS5VqnUWOrX2ZuLF2q9PRdfu4wdPG823OTkvaGM2SBXmR
ddPUY+Ruz6pNUcDRJzh5YgLj2uL8dEXd5zh6ZZpzzVgBtWtt8Y6VjZ5ghoTkiew3
n9BwQXM1zDx/GyCS0z3H3ZgaKwmgArlWj2ChkZwtJle2wblZ3pr/vas2D5ULnVld
bUVBsJK+E2/gHd/TCVxaQi9IDyA1a5Mk21dzRkc0cpsO7Jme/qBYHiffGvS5wItr
ddCN2u3bVyrHEwr3f8mQBoyGg1ahuy3dVBItAlEybyyrxz9NRYIGCMy4PgZ3+6wy
ZxfIyaOZN9b79mHaczOJ1rVeAgDXxO7pT9jB1/JCPFvJk7tVq2pjms3WdPnrKNVI
SclMEKCA5MyfgbkCbrmQAY3OHQdvi6lVZHo+45XSj/tmZdDB3Ir+IETMRgkMmXyD
6IsLER6x/70Sz8wQKh+TUPR1jJqtja9rKjrgt+4yZpNNtExeKD/5qwPRQ4JE7gd3
TfL5pG2YGzqonogwZJtpkNYgoPgFKRJNXUYFvKmDm6kvc2OLwhhlTLZYPxhrT2UB
sO6ZQ9+fcmX0H05/j6BuL2CIoQPrNubZaFiIfsCKG/MNanLXMWIjztjvC0/WXwiZ
U1MerftY4GijUeByQNmGJflG2cRPpswCz4dwLGH/Q2vMCwtJLPH1692xYCBmG3cw
gVE7E2bTTTMLR728l1w4fRq+uA1QEegRNov4yqIUqE1FVbzgmnLtzu95wF86Y7RP
Pzde64RDy0QRPEdqru8XJKuQ6SJsXqPHloHK47xcYLn0LBe7/g7pfd2Mh32AQtKI
+Z1SR6X3CvlMiCUFBu7Ht7UdQ6qV66Ge7RwOIwCFWuoY2zg6i/xCKT3Xf8UOzm/Q
eZS5ci392wguQIOpezy35SAYJjnsOntQDOtiuV4E0ugJt79x1v164yHS4tE6732I
YTK5TpnbtHG6RfBGKqS9IejNtBy0cSP4VH69Lbyl9+fpxqZcwJybJN0LQD+aufaQ
KR8FsYByRl7clAE97g15BmFBEV2xJH55wqb/Zvjfm4NV/xJ3fjuJ88/Gbu9zZtkI
yDfBKvb9clQEX0kpiYOuyBCdzUWFqpm4a3l3gShSKIs8xsjrYD8FG7O8TMTd1WLX
KpwtRdvCqrl4M1jm6of6nIPFwqpDK2gRDK/5u8DdZr5dI8w25PNpl2ZypCWWXCiz
4lOIIyrjUpyTqdtF9Zf1EV76EdFEGE6XOsSLiwhFyMC0avQYUEjw5Q6elEhQqhJA
vw9XjQoX++Sner/8vKdvbuLezIAexc/npakswTQTwO+CVby9s8vg+VR2a6CIYc4W
mX+oDIoSO9jYnvEfkPhy0TCNKiY0zcFVZeMxQkIUZ6fZGwnCd7h9Rcz+X4wb1iHx
V/lAABDExh+iyFe5A987hIomXgYmVqmorC8+djc7SOh/amGoXkEGsjJ2bjKypRuU
cSC3Ow+j/tEVCySnfTZ3iJEotH2Pxif06KR/HjQJ6oHEBKx1qTIrS7r2MnK9NuZF
1AW0HhAzjvp0uXdJgUV2u+pC7ok4QFMFEJ3hjY3XJsT4VEsOqzlmo43r9RpvdOv3
UyVwHaRsn0eRHaXD60AYaf+mbnihoRC5TSoBVagZ3VtIR9fE/dKu2YUFliomz/20
IW+DkMVVMhDjvEh6J1x+sPLAeOWH13Ti2UAWWy3ohAWhw7AH5V7osBkMlVMLrc+N
uOwoVi6ihG1G7bmuu+kAbVwW4ImoPfuOQx/TMxhizAoSPhhzINrZ36bqPiOqqoly
6XlnxphY8jx24HSntYUUR5OVZQCF6DvRAv7s08t5cTvVvnBDm9+ScgMNb4WYmWtr
CIORnXAhgNfrQ1zHUSQ7lfopGpFzO+DiY2Ig7gcS7SATf9FSYlqwc3PmjEFfpwGB
W4mmL2+Ri2JoNTsKMI9fxvvJAIZbuxRZ8OdA6RPbrXAN0NBm7AvLfdNnW2TyDe7w
+9ag/486lNCfvPNMeaHsfMTJ4S/scVOEnQR9LU2KdF6jdqKFJ8LKb0NN6vr+N1Q8
Ww+oiF4N+hFA7ZcuCbFQhMV4OEkZULaxk+ACWW8TkVnGORr541L5zTdeaZxmDaR1
mu0UngUqifCBN9Jh7sJ1MVUIyEv00NwnuTDVxWsOGGDhCTShVFYLL87slBSYs1e8
1nuAVA9KpXk65c693NlNRRuf3BOTGhdwl4Om8LiOpwGVTcJfT0uty/cY5WWwyZhb
T4S0KItKdE091D/ozqzuOJRD0wTRhF2hwWVVjqGvH8TLlQpg/RGV169JVVlyzl5X
+gc5VOOSMw0XCIMwXYRcvCMFMn7qLEl5ZZ+q3pPj6ya4U+PsvpSh05I1ebJeu2T+
WLlOpJGaggcuIfD3GbmZlt8UmsElMcTZ+ZgW/0WC6MZJlEjB/t1tZbd60e0PDpUK
jHtqeA1aqCglkz4txYKEkBqW9EMXOdiHyjhnyyz0vAD1rJTzoZNWlEHZeNljYjrC
Le0yT4QMAIQCnCXxxxPUh/HUo8a8lYIop/BkMG/T2CPtYlQC6HtWL/T8pL/Mf59K
WRAGkour8tAmDFv0vAUDdCQ6g+McZbCzhNiyL93HkYWlDCYJ+40pznjCQ7MlAo/b
1dh4vAEHmfK4YMAhobu+FB4cIlTD3Np+1TjuNwVeloqWz6WXR2Mj9dXCj5F4/nGi
v2kVwSoxWHRjdv39oGLupHY7eQBsKMCMdu0vOmkYGl0UUYt6Mq80XiU65vIG35GN
ltAGUY/VnEQTWyfedcmrdBxwtkgtEoqOgsib365TZVwC4kiS6O8OPruu5N01NmNa
ReP9DyIXlBrnWFj5B21risuBG4BURO072a59OQRcYpuVuU7X9SRNp9E5S+D1KhZE
g1E7CeEFdI9/P2P0RYq4H/NLRDpg2FnIsVx7i6JZFDTvlDhX5OuZ+PVp9b7dKfVq
9cPh7NOjZIWSQJxX17eNXLCMof4HuHvKRVSAx95w7rkjtS1UFemdZwqQAa9b8xlA
4HrG6GRSYJlQvN7Vn4xGh8iltaIrWiC1fUBgG4EXTRCfg+YGzfTSp4QZy9/Qk3gm
9RJpd56UAxedm6L4ZZJO9ww6PCx04ZU4YZJQFWpOpj1kKN8xoiHoMOZRus0PmRwt
1xBcvET/b7kZ3rkrybNkJKOhTTbol+t6OTnfCb4f1wiz6fogkQBkxlHOeu50F6jy
VewXE0uvQMtwtYT1X05+dMO+Kz6j9cPQ8YUPlj/YkJQsKgYrFPbt4wikMCMGjr/W
25Bq+0XVnD4B0efXisdocv9W1pJwMQvqzwmndvVKPu4Ww1OJdSLPnCpngvX7ciNx
Eb1+2sYc3WA8/IyBFbX6Pdi+4bd4UWV/+gx9zxi6scYcuZgYEnpEdFoTPiKnSXkp
qCXb31wAnLg6S+kBPrZgz+iImuhH5UN+MwUpNGxc39s0ISIcOZHq2rIVXoC0NGBB
uhqXuUU2zOT4Ht1W3snEcvK30mYEyTdm32z6gSTZ0F2TIUm4LE90Ua9xcKN0rHJV
IQREd58PqrmftBXjAtyicHqXXedMSPQDAZuE8ZUefn/Xl0Sp+WfUDnJIrnX7zwaD
BHz3FfWz0G4S3RTQciY6hR2s9c3/5NbzFC1/NGogrY7KCCHhauMydK5qrVm6I9xp
q6C4peWhav42iAkV0R9hMTFUp9wX5eCEY8jt5h2YdgrUiCfh16qQOYILX7qv+Mkp
LX2Dsgn5ICvUDEizJnQUTvj4LFQ82ZKhWtZK16Ju+XC4tstyvV9I+z16JMQGvA0k
+XntuvBFCc9aBFHt9oFjrx3ASRAgXzBpjf44CAq40Vje3dzl/QqX4VjRa+6vrjIe
wHljOIBvly8GK52AEzuly7qAf5L58AW4vz6JufY8R+VrjlReUAa/G9M2sgpmB9PP
pIGyWcU5T5/GGg/HEUGPbifOoMMhzsFSPpsOcnpflf49PAZyUoXACUhiPTcLOg+V
YMakTSmHGdfytbOs+HB2Nxga542NVwyqDjgPH9SNOdCQ8ewJjdln1kM36Q5e8Iho
2nPmDWWjyZlgsXSXdLBoAKKsn1oBdvvu4bYKBEyEXTxFDY3kvvE2gOoe6rI+gZeQ
BDz01BF/0nOu0uTslpqoZJpXg5iSjO6BIhgxPoRyznljtY1wR2Xdy9MhS6Cms9YF
NUOgn1qfOmV1znVC7aM4cy1F7+cYuEgf1Z5tbyIcM+p5nKARktXLYrA+24W09iz8
wPLkxvDU5PoBHmffkzjuhfzHnwzOV673K7+16iW9LjMCRYcw/xXxrEgnnBSozjZE
l8eEECS6tSeWHXTsx2B0fOPAdgno+0Ohaf9hlB+VCZJ2XSdWVV3rhB0taE+a6ibb
8YPmU8RkM29zURN/5OkSxFzobwDnUME3cmCB6sO4E/uOmxDNkWdmf+fsKoYGZfWU
6jgpOXYidZW0xR7dqQPvOh9+2ip7+exhtPTT5di2HOSeeFzAUTXjRDIdmVAzeQSE
2byofKuCt3V3Y79/5cXdi5e/xJZC7BePEDmM4Y3KVBGC8FD1zMYgvWcJWaLCqEbe
qdbYh9laBmNNQ8JdNe8rsPmGiiOTpg1mCcROoeHqHN8FuopWpNbJkiGROoOIWEcG
FVCRbS2c5MaXdnC9ycNACXBQ4FITXfunAL2gBoTgqQaHE09cVmHjkfGHGO6japdd
2QSy/6+EMQlqXti4eL/JVR683csJG1zQY1IpBON4vEl0O7Ln9Wt/mw30l8eTwBEy
KqZjgRZN50CDBTwdPn7J30/usO7G/M24YYfYCSjnME2AZVp/plERiHkrSSwwIFS0
Wbhv8jJ7mvCxf1y9qIEReJwf9WmW0v1eZQOrq15QFncJfKqhcuqgwa9cV6g6yJjS
vnljA/FtyMPgXy+HRqRcc3+1GBXIdgjcc57zlz1buF54bKuV5zP+CQj+HmSd0cyS
VMuhhlbmYMm++iXHkXPYnVIQvVPrPochj1ZjNUBr1pmRA/N84HK8fkSOkNRmPJYf
rhs5qTZWCK1rAKEUQrffFm46Nnp36DtqRN9KmlWRWqnYxU5SFhWiizVh7ODt1Rtb
uFEGnfC6GMUCE2bxiKOczilp34dc7gkZycY3iDhWaa7x90ZfrjVk4IDhI56o8W+S
5XZRkr04UjF9AmXAnhJUAuBJ6Ce04jmGR/k/rWPM+CsDehyKxI3QXIh0pHzgAnaN
gDRRamJg92SClEh87TsN4K6SNxP9P16S/NyBdUg5G0ReEMVR+aP/vx9NV6kChRVu
sAoLNOiZ+hlYIYXY5qx2ct96ndTMzeVt+PJTARnpsN0r40ackZi+mQgA3Kr4FDqR
f2/5JYy35W9B+Zasn8X0AskgI2W3NWX3WT+7IbYj186Xd9jokywbCSQWVWJ+0DhD
nkv4UpQGFqsvBIvHL+wJhLxtYenE+GW07RV5lzDPCtqbSsYYtCctXCRYz0Vk5KwB
fmUkOmhe4pl/kgCPXwludD7CV611WPoM4alMoylfp3dFRHYAztdIp0l0S6fcoYPg
a0I8qsWGDlMuOkUE/G4ALLuGfbsgA1kPeTrZdk7bsCjwmz8n7jZHfAy7Em7I6WFV
bPcOOkwbu2vQj8YOFHxkyob/KpBukuTgwUcnrnwlynGFoili0DVCqbQ8F422gYkm
0orIASkVc6eo9GGNMK/8i/ehHRH9To6FYEHyuIw0WU9Rl4qjyky9vpeGUfA3L9l7
UZFkBYk4+Hy6Wy4KfeXLwVkFTEzkxPZ9mkyyXRwsUlpNGlNxYyfc8j2px9HMI62a
DKgT3pAftevAXOentHvi8cSuYPINrwWgJNzXVUXDX9LTyy6Zsqq2pJzHybhw32Im
pYFAiRPibI4rvhBzeJvLxtRzi/FkrPHatLV5JzxtBwsQqUgWbJapgiTX6x67VeS0
8sJ6TzI7/G7fMz6L/RQ5QbRplESYo/Ic9+4Tevf2frt7Re3H/SvLmmSxv5Q8ltdn
DEBXguG/n2qs5YRguCrwByrVUy7eKxu6RWEM45x905k/CdhP0nSzBQ5RQBAqtY4j
skHe3FNbF7MaOYXgSWvy6U4MqqMGH7Jql/j3ARLxcNKgz19FnBBbmliO0yRAVhYG
n4LMlOA7WNKIcrnb/x48d41gVHUi9XZJzURoMOxswuKVC8kMiXYCtd+bHuqdMhAk
c3swwAH+CZP2B2ApOuzfvYQTAZOxMHAFRUbVnwDAQ6vZfiRfSp2hocuFzjwgF8uZ
occbQwEPk9haeoVaTqNAqNHQytXwBalOMB4ElTGMtpyuEngIue/2oK8bs2/HkdEa
Ij/GMqK205RD/UO62XLueEGxWwM5odT7ygYm4HE73Sl48uwnf2i9woyAnIk94GoV
WY1YnW4n7zmFg0jSMSEfaLXBYalJWWcqcdjrBgYm80qHANeGNKX/LKpYFbS7JQLt
XzSnMG3hgt0Kpkk42IacO+XGlVyFDK8HBawbhP2a5+QOEbyd7/FbX6eK3elCy/Js
QR3KxKtO/tbjiOHy9BHt+oVQkw3uUHGyVCUQzJlRygZEMaMX8KapNjMLGzXkAqJV
AXDIRJJVzLz+m3Ds052SJRC4nj/pckCb/ONqoWfVVFVTk5YmhRg61HiL3TQ36NBV
Z2v9vsCwj/xxvY4MVKBUZYRYYZljaY+C84QjohlQIXg1l7en5CLTcR+EAaLH0T9O
nS8DcwiR3KyX4FByjhQm33bkkr/2bZ3n5lII5f0KMJGUuSVKA8t1PeDhKxvteSH3
c/b5s0WmWPnOPpQYXAcuF+Z7tSL6xi0AeBm6PsAjCfqQ7IhVW1RT6f+mVpGM6SQK
v4IgXr85yzh9GNQloEEBNSBfwgbLk3eG1BYXH+SOup9mkOR7B7dFgklwwwb7uozR
4ez8tku9C2I1Aw8BL3fSayMYQvCIRxN2aF2Aahlolo1yAJN3DLqksuMpcsgofSjL
uMQQLQS/mG1tfIdwDIphNh2r1eCD1YjFSzI8CSU4cvzetNyIGK+90oP14QHgqNg+
QWvRRN/SFZ/7T5UjIKmJXzUUGLgV5pBNqRjrR22WwsY5LLKlIQTIxu1psxpAMJ4Z
JwhWz6igAxk2mGnpQZ2pK0wx2IUgkYIJMrJeVToPA+X/RMKIODPGpNiHe8I9JeQ6
mGopwGKjtflm0CCdeEPEputhHzcqnFeMNYrjZ8rV6GUnS6BHgUcfS7AYMSB96gMp
No2KVaGPY6oHGdAbiCk9QUQr+aRElIO8aNqvq2iRAt2RuEbwis+vF7aN0ZjEChEZ
O4AtfdGsCGsdPAHC3nT3DoQUeaFAzfavUABOsL7EAga9hVt11JAkQR4bXgrJVjhu
1SuzIdGrw0vuMlQtUZMYkYwTuCdSokDhSngwdA5JCdAXZYwlRobs0uW6yXMZOD2p
lLaXG/GRNspeEBMr5ea7f/EJZn4A2swuHTCvMKwBsZ004W6ElhL8yNaMr2O/t8Kh
CXNZa3/n1lsEXdTJbwlsP2c7HeDTNVF4+ZLeOq5hVbX+Acf8ttX0fVmtjAfDvYma
c/q3ZW61T9VNDbRyNCo05CozQ/j26aqov6CJdsR2YlZ6ZFAmqvUAlAwy7Ox65qsw
MB4VmayMW5lcIvK4K+5JiiSuWwD0xyG7UWdfyN9kpyZOIM/MFGnovzx5hn/pmb6x
07n+9MKoUrI9oMRIxzpM07pw40eUjfytGjILcje+9HHwRrnEZnZG7sJ271gWTifc
q4vipzlvfS+oaF0qAj/dwy/4STqYxodVgAPezsZ44SVKQOzC66Y0olEStts9hJvm
Z2iuRao6FrtCmAjXzmvLbrMnCcfIoGFqZf0mXjzc/HROQAX4nVDoG3nzMZdX8y+L
Ng5U5os8LalvN6ddJ2yxUc+EeK9UwbirBvosETOghh14qYBR9KHxAYAMfguBWi1S
H4Aza0m5R8mwFCWgfFl6M44GpmyDAoeoWna8ZSERir4qse4qmk93edG8KLe7U/nA
1nzroHQ7LbJU5FlrMMwoHAek0OOaerATdDHIum+2/6CXIdUUiLQFJE8NMskE2tPF
idJj8R6givess+XQyUm6S2J7Qc/+rcgJNCB4+5aK53+3XOESrbrHKTbSxZIE8oyp
kcFNpLjSdaTRuxw2jMOUIF4jtXL6nyTUd2Sdi3gJ5FdUCz9GMc42WseQRisXuzA6
pxeCnqh+gvMb9Y5yvuv2URez4r7sfUzfrJ5zTx9FjllUeTP38uHN5nJwNCua4bHu
HKer2y5W6HQ3LDZfo3TS7Yhyg6+9390K/9Iqyv60F3JzVazf/kUQT7zCPhHkYpJ7
O3lBHnxiMHTsnceMJhTiClwmzDc5e5tyf8c4/PRaCN+q+N0WHeOvR0B8yPJw1wNB
81OFSCyKbZW91+oiGx4klOh7UwCzMvC1FklVGUwwESCANmsWXAj68SmtSdvAPiWy
sFmPvDBOUPLj7Ae5EfdbxL1HNmtDYAgJJK1VxBAzAJX9gK9Hs1YfK5qZNVNnbv/8
AJ6aLPkXVyobEw0QITLFzMFK7NJee6jqjA5U5ewWFsKr9Zir/UwBJ8YsptPJ2Ua/
J5uu5+m3Yc0pRQ1n5owUvKO/sFphrKnAo7IRl5jXf7l4oXD5rk7t2axTnxIqBKIS
+aNvnwP3KTRTqGJSYyqmeDHg9KVrOF5fiW6N7bf6GqZ4gvLEPIR1RYa3QOWnwX9g
ommxSH1df4DnatsHKErFNA+z8NKwTLB3L9xrxBpssv+nS5PllUEwKyg37xNivcs3
DnM6ggZc2WT/VX3MV9S6p8N7CnLjIRMnfiweqFF72FybVF1kUG/UEzQGm9MUvP7l
hnRc8PC9FEwF+kUJ0qtv8YdrFtfGAVqtyKHiD7d+zErk6/cyp9ylfIEn7QInz7zf
VJMAOtjcp7mNlmryAC58CrjpvnZMD/qPrLmzKK6z01xV4/GLyM0jl1uLSDjlpstU
2hiuRO4a4OBSQ+sgvNF7UHy65p54SO5fjixcAFi7+6L7TlSQgsDWnMDu3OsFLJVw
EWwz0GTL6mDKhY4y/iJGYiZT1ue9ieLdBxcJBRohSBP1tDvPmyRlhCJtO8l1hQTB
MDQY6D+5+erNqQGI3RAQpJ453eVNIWLBEwfa4CD+55ghG7M80oNnlTZeE3FkJF5n
cm4ztd9dIvcu4HjVX4X0DPcsCQp1ms3NfDGZnBT0qoNnh71DIv1ay2hIVttMbLNE
eo/hYNgisB8UPz6qngQAIu4ENTEaK9GvzpmO9yYEZ8Ly3PyC+6KmXtsI4eXL/Pap
ioS2AjaBkKu5EL19Qun07nx0bs1Dm6NfyFyJA11L6RHIi2vcEOwFK/c0ItA4GJRs
QEyth1Hr5JAiWwLuDBkIdH3BLwlCdwfLQ4vHldzCShFwn2+Khj2+FpfXR8PA7OA6
iLrt45L7UpLl+cQgbR1R+CGBZNNoEVFYTynxiMOxO09R096RrFbtASkEjELSouwZ
WFmcSxoSLQzs+jtoug3ze4zY/fXXOzUSL+uee0HIUNBlLNItaRjC1cNCZvS9bnZD
HCMz2KTVZlGrxW0+ZQYIKJq5cuJEmuy3RP5h6ZFl5ueRWnMvNROBusI3r9nUhsht
6aCunUMTwsTs8FDjV7bJ+ezSYoDxMYUCHsqNyAaIB8Ur1zk1TrxluYiMwc3devkr
Epf6bvgFPpRN4YQb3nVVMuuqeHlJycN4eQFPvkMIQ50gZ7TwCjwXds4jUXBZ9cJi
xXX8IZ2Bfx3OXxL23LbCmxYEUJ46sG67e2mEhyuHkmN4o1x8RqB39WnSNUZnu7I0
hmxRMqGHQAQuC8HHIIdFbuBSda3rcGs/FXAalXy/Zn1E2bsZmX3jpVEenbJHl9cU
s3DzF6cq6do3F49lL7O5cxKIFvyGtl+mGQlfPWfXLhUP8fz3EljhnV5QLY23LXFC
KzWZfh3WYdmg+oZle5Oc6d2nyvUEwyGDJIFxzJu8q6atHTV9gT+e74vlTmmyTws1
EFnLLofQHZw38PM/anp2eQQTlfa0RUzU+8T5FTvldL58WdPiEVEG9CgmLQQE//9d
jIBQNo6F44pn1kHFBm+TH9NDrfXSG0KplZyOQSvG+rlZSdx8S3/01RRcBCVhN/3B
U7Mm8d3MwZGeD/wikUCz/T8YQfz8WCQvJG5AbHwVA/Xkvt0oxSSdG07BY7AldbmA
Fq/KweGVoRoWgkGLwkRw697DpFSHJ20IXWPoKhtX5zbDCtn1uMoO+Odnzq/o7mht
5lSFjUsp0tXmKuhKYt38doNBmQWNgBfnMCLTR/wcN1kzbiDmDuHwOnJoJrurrrDX
1T4ZJa8Z41SmfqeOQV7sBtuhB6wYiidi8DDXkclf4AddxgsKwwruO79BckGDa4pW
VOuu2+7Wp0jM4Jhdup36jJuq9GE9DcuDpJ2fZwICtQVS1GH3632qWEpeHDKuOs2l
qKqnZuZd3s4X77Jtz7V0D72gzNXYeW3otrUMHQkKpMf21tvUWmj0ZiWVIXd/X0Uq
RZ4Dd+6XcUtd+OSxOs830O3Cr/j3PeZo1QPyNaI3VRNyuZpXXq7nNQE29S/VWKzQ
3vY2yAVlDrXJCLxwdHcMQ/9eJbXpfxxTpYQ8iKr/F4utfzExV2pIQrXbkONUQo+n
6VKriah2kKJo8pGk0O3lnTAbjn3oazt+TLvN2xuVZimOON5u9Q67zAZgu8ng+A9N
LwLFWu9wIbNc0ebVbnzlGiGO29GKJ+ZmUVACzWveLl1eIKgGO765EY29l/vPFDEV
f7DQ6ZNvHHTH7gfr6YQXbKJ0BMgkWqxf8XJl99l4QxWdEwX29LesbagHkcvbx+Sz
EFMQMMmAkouzLSAUHNxWuTcvNw51X1xSxAQixM9jrxlVRUc0c3jvUpDBBZLJFtc7
H86mHZZSV0V7kaJctIjrNhf06KG1+K01zVtSwCNURgszvwvNGKUUZqq2TxQE24LB
2UtvIlUB94wM0JvU2KDgaTJV5RJj+N3NsHpELPMlgWxvYZfRzbc6JyIrNIydqKrc
5E5cJBiWfL26vmPd3TGZ5TUciILiSa5/IMp+UB7m1FV+0caKdLxT03+OPT5uSNDR
5hU5ezDmYXCCHlFm/xsTM4SePXcyyZXU24t/IwEtdjF9UFzVvpcxW3I/MshkOBN0
+shJT8gzQDGSTTgFR65zXB3dHqju3lQaV7LWNwZftlv5+xX3hH4EaxiDw+w6WgyP
9yytvDoQWV0WWFYNQ6pOlSOKpmvP/OIYvM70JUzLM7CuqrxnDYuoaljarjGzsbQ6
TnHedZWQNPTs9+NQPu/wKwOv/o79wuK1b2Isdems+b3XfTXz7WPglBNkzvRQSmGX
ah00g9aHXr75hiGauqw1jT7FSUaEqvgEwZ8SSX4uV0yjLfn48NY5mqG7bz02OcBy
CeUJVcuFVEVi4TzyfvjWVIUz6rSqLRfVI1NsA8+1vlXABK2svQa9XKbPu9m38Wf4
IqUlHdy1NgCAoRVIkXXWgnIQuTC8xHmgIEdspX7jlaq4iXgPNC/RMfTrqae2tBtw
SNCpyyrL9KEzT0xQUnT1dwzbHXP/d0ngy+t7Hvgh7hLsdtBK5sZUzUuOak7WH7v8
Hxn4nxHGykAA5GcJiF22NMRXi0TH930rBGgiF0LIf6dGiKVjip4adsbfqGYDhkZS
ahlHGtEXXmETHCNjJUO8rIrLF3ghY5Zrnb9NNWcMLgABKhrIzGXIf4kjgUDLAQzC
3RxKZduZAdKasuaOfEO38wSk0hwRMQWKlWQfOWGi2AO/skeZpAKiBtVuEkI5f8Cl
3/e1uA9G8fF0kXxv7R3ZjYP0Vw2sKE/Cw4jzBw4gKj6S5VVkcUExYpfrJrdEh0qY
d0ESH+Zkkdha5Z0tevAFkABuaEzY9o2x+4b86iYtYZXZnE+LNIGVzcJwnT92Kd+B
1706vwgi/o4ui+fknBKplT+KtxF6Jj+aZzrdtK8FvC19bU+IN3p/c98Y0GzJQGv7
Lv8Wm3n0672N0E2+AQkx6mmTcPH56pooAbpyQN+Dyd9C3Bz4U7Z/eep04AioBjsI
6YZZaNuR+vsIglxnx3+Bk/NtQpKA0HHj+pav/6d5YUN7N+oM+2ODNUHI1iA6zpsp
ncsLpAdBVlZGoNazhkSetlMEJKy29yIde9mnJjBXZMN1XL/DQtGVZsgpj4ebx4DU
P4iRDMTA7g7VdSNic6FlQrSsGxBmTVZya4yrYHUPf1/UDKH5oc6BZ7imtBiIgGE+
mBHsRzKO7AB5UeITpwZtzxLP5TJNyslPKy9fbey1XZ6fMqGoIz2EGlFmIbeoEWhW
+78cYw+4klymqVqRLUmSwy0yU4myu6fDcrvM8fr2jswR2MBOxQ3jDiH4oOaJX/T9
3TBiFStf85Qmj4n6UExK61cYKWcUnrFjKXCHnvoKpdJEnMK+R3QUUJGl7EApRBon
mlK4YH++rkWT6vsK2xJzSm6fCTVWFJeIWHJ0k7fweTEEwh0J4mDhlVOy+BdhPe0T
Ovo1bgQ+nZ/Iu6ROW5BKEYRasDX0zZqcS7oZ+HsS9Z18FTeHe3DUKjnOE4lrZ9n/
FfyCHgeNJpwCI1jmDyKuZ/meajRBUUg5Rll3feDvXtusgy2aJTB53+GIaDN6myb0
3QT2/YdnM7KQssTf1T5PWureGqzR9SDBpFMoSWT6TQCNLS5moE3Ge1am0CbgPEX5
mpAh2w++tyCXkPkBohoqQ+rqLpReYZ9RujFl0kOvxpoQRjyAgIiE33iDl369NVoj
1xBUMw2ZDN0BtzOgY7ie71ljlDsd2PIz+Q+2YZl+JFj/x5HLzM/iJyxfPGZ5OkZp
2BBFgx3AGv/dW/GkTIPyJgzwaxmsQKc2j+2ZpDHhbwVSEEyD+aHLFO3Y3PVwik3S
qxY2IU5Q5/YWZab6YYvBlwlo8IqxExkbOpbxs3VdE14j8y7IgdmaIRg4gOoiuO4i
+WGIpiVIAAWeY0vKcP8+YnBNPuq9kUrCxiVXrteW9p60Hwi8kexQ+sqskz6oi8A1
ii5jFtGA8PNXLMYPWXqyl8eMmDMKTgNa5BStGEBLZ7Mwl2pSQK8y8bCoza+U6bbw
lntQNydy6AICk51zh+ooBS3ZpyFF2lkyl3Me6ceDo8uZKoO+q5YMJL3Rv7TDYM5i
hLCDa1wYtHiNtDtcuT5/jp+6kxreUdi+W9quZbNVbnDXIifvhDIxyN273wSnaL2B
zJ03ko2lznr66VTBuCibtWba5FCEtbdTEWqAGCwLftrHI+cuy6jxfQW7Ma9TIhZt
l3pEyQehxk/fgRNy4UkPXUirYzuQvPgNbD7aEn/HzLjqyCiIxlNQXojNwybBhC6W
IDEsTKsvWQurVvWG9rCxTFvZMpa0nUKLy0BzyLpOTBa9CA0Vl6edqaQr6ux+zP1Y
gkThS65zfAUjUAMzEnPxYSOHm5ZbZFiFYA7Dr3+yoIHFHGcVQu+bfIMQx4Ad1oD+
W8e+EJ2DJWaX9tzXRsOC9cUyfpXXQhUD+C82h/X5Q+v3HxY8Yqj7aS53KR/7AVFW
qEAV81A0OF39WoOVpjaKcZ5AIzFeqPGUjm3OAJUMQWBC1WYptnZ8B7LdcCocjVYZ
K3QIPaHmCs754bFC7G6WzgOlUxz6KXnN82y/yw4xlRfdYcyq97zqdQhg80x3Belu
mlV97giw/mKwbtpol+9AmB5AsODj4WSi1jN7RSo/kZnR1yheaM5AyUtsIl2C4/sb
uqXaZwYbI0ajLMDDuVvZHNC4NgjEe98SOOC2FXpKYlbJzJ44jMIkohVb0WvG5joc
cIP5uy6FsIgJCZQAz9R1DCcZumckENdvcmW6c6Bg9Vkopx9cvjTZpmnKahRU4fcw
ZIqtZP2WIBPS74Z43BAqQXdsqFBA6pgz7cxS+BKM9LmUPMzX8MN0HUVZ3TrbQKmC
3HbJGbrpnBoyIN7L6HA+Bko7Hp4p4//bXiLakOU12ycplDiFV0KJaKPrS0EY8aYU
FmxKS+UVUfxNTJyR5pYlmvzBeIjBD/ftoPDjDk6gWg/L6Bxl71bNJKvfLBWiWjw5
+cUADziPSdCxKsBV+HlCofk0W2JSZz4SOb76QA9JkhEDpZGu/Yxp1b9VW4M8Cndf
AcJ93tRabcB+QHGvCdNPLTU3BM0kTA4hvVlOXYTqns78bURsnJm9IhVLySJmGvvc
Kzk/koNIZmwsYpsdRSzm3MP8Wbp+2ofh2jmhDONrFhrEymiltwOzkBHjbyz3faEH
MIq/daHke3ie/ABlIyP44kfG04nvSNBskqlmCKD7aS8ORahTgfnqOQyE+5/zx2V1
FFI/HT1+ebDemD97L11XTw6FAv6zvaHiDC9JTYeCk4UOQOw7QrCF9UfwQcbjKkn2
KxOyAVpkn9313xsWZSLnE7Klfdb9cWF4fivsNuy5z+OKqdpNgf+adxRzWqKNd0RF
+SZwdAgjBkMvYq6NOoZFDvBJJx/keLXSEAHWeZNR6m89UPIftTRaAUezsHqCoTBH
nGov9bV5ycq2lN/SlTqQxjupwEQ+Cn3afFwV0kzQsJ0Ua6NlQEWDPmZ8b/2lt01w
0T4cYceAMCPWD05W/KsGI1lwSa4bCiNdQHnt2IW9xCpw5uR0c2N8GVurC0jQpiqv
aMQh7XqULSC36eLvJPfSIQtTu92z44oucpR4wxwCJAfvpeczCk57ym+/z3x7fmBI
syhnvdA4+PRmAwriw/6FcMtZzw1pNm007EoeMnnRNtAbjEaok4vfWAfb1FWISPSG
CUjtKkVqFjbxTuSPw8e5VyZIbN8StjUE7Gz6/kcGF+qvE9ftlaA0IzZY6N2dAlkF
7eUi97Q1IA1CtfviCKxyVcEEg+JHyEYjJzVPxjtDVYDJDZPFJIF7T348JokHGRqz
pBi2YopxnMRv7WLPIayb9Ns/7Dd5O4Qd4al7WdYcBWfnACWh9Ts3j4ZNQIQBmNbe
lCtsENU97+Ff2RsS4v2Z8CM/DeQOhgT/KS0EgRdHCjpMWOD7z0SRtKHGUBqG/+1N
648BQ4n6o9s0pCE+T9Xoh1S22wpuRq3qgdmGwug26HDUegRl783brjzHn0FNpxSz
ALUT2MTn95MmGYAnR1s77WenRV69/Jght4Ld36QXIOFbUzMUIyKF/o4AwzI1bvqq
5LXSr3p7RFRvOeqfINvu0k9eBl0KxBKjqZmVRD3E2e41rxJ4+bk9Ib9tjrRnfqiB
Sa8W2Nt9wGr5Wn8uAXCZSow6q4ZUFHVI/v0RmMiDUle5oz2KvtlNms89iRL7Cjrk
MTSDImh4LQVERfXGxAne0rMtz3PHacCzNJSjM3vH4kU5dNN+qw2Fb6WTCMm2mFXY
+9mggxxD4eJovPtWMQ1HwYOEQx5YR9exGqCqh8WHvwpN2y+pb1Cj902HBhLK32c9
xxugqaupA4CeIGWYBf6X6yxaMhhxioBWAwahOpYl3QT7Iamn22RnU6r6HzwBTBmo
sZWemLvIWwQ+ut9m6TTq5kKE0r/W1e7LTO9Gjx1+3I9Uzyi6trifVWRdP4EaIHe9
D2EdTjj0QtrH1fp6EysqRz71iFj9eWkWfaSRmw7dumIDxCeSBnzdHATFiIFMqlIm
s008Hjjb7F4gQiA+Mlp0d3Gr3bSXuT2ale9jh+EqyZeFZXvmUZd7FNvXWZsWWB7r
HqmAD8f3ZBDn9jJxLavZKUu4IdMsRkGv2TdiVsC67WrKk/88sul3TUQzepVufp4a
E4W/5gJ4a966nK246JDS5tbQr6A5t1tVpUQ+a4iD8YZirxdhaPf7cfNo/IQafv1T
8wX2JyxD6iZpfJphFmK+3dRXVlhV6DAM72xM0agPlB1uuhs/ROqbOj7beOyrrXNP
WJEASSVnGgzR+dMItP3zU9x64YzWhgQ9rDtUFaMHbjeIGgsqPBIJEdyVvRUNDbND
9Dm04t2eiovD5koaRDDcNXgYLF+6etbpIw94Rbm1vQEkAftIdJOkArOMd6I1TViK
qJ291Z4rnk0pb7UcYedyhnw6W4oljnvVxEKFHJ9o5ps75jtW+O67Bp6VzI5rNuGz
iMsWHr15p+bq7DyO4HoH6i/R3NgmnRmVyZqR8mSqCo5dyx1lxi5IB7WghEd1apVw
Kf43oYypzEYHfUy803/pml6/PwAMnRxum+XsG52ssUTePaIys8X5E+bNmSs444ZI
dmd+gf5nyPVfHjm13Vr7yDHznE01CNyeq1EkQzs5Qu415KwPOJX7kfnfrqD3QaUo
jXFheKCFxEU/Un7kX5CMjrehS5shLQ+NX3e9/tUq0tsgD2SZq40X7Fqyd085vvLX
PqrgR9y5KVVMw9pr3KMnE4F2RxIU/jL1iDhO+3Rz+iyFSeO4gPLSFFX/MRS2rFNU
YobKNK8GFrxAXaqsj/Z+DjEPHzBGTnGHEYemHR0Ei8FfEWv2ONbkf0Fh8ACv9sag
rZa/p2XhwgHjeWvsvfUv4WRCEteUVJwmXoUvD4I5N4Fxe5eerq8E7A9VLGFvY4br
i8r2CnOQOeDcSMFo4xfbqei5+QNOYriAr40kvaNHPBeyNPeHFeDXaMC6aNo5dYAD
r5FUrz8X361JodJ4iv+2JpbFgriFsNqnZwqHKkXTFMUI3LvBweFbjkOT4ZgKgq/T
G3tl/CU5+NEGOlMMy9v/mryqNua/HhiSIgqz7K6hc9t24fBIXlVuG9bxD4ZuMkc5
9earG7Qu/hf98AKabLb9439u1X/tRUir6/yIHTQ8VJuyWlvl3EtH1Lc360K5bA99
U4RwYfsXW/fexL07tCSHSwdAYiGpDzBOFR0vtcM4/1yMz1GP13VrFfekywfiSrJm
2ivUuqAdQcBStOqM88TxaRRJW5SJ8h7UTDfoc0ENIDmQUs4D+I5XT51sQTVOxyqg
fesfVymQUKuiGk1+FrgQ7Jb8x4gxZcZpql+QQnSL7f+CN2EVHbpz5W2X7kdzWnoy
6cxnVzIWYAZQDIS1FmM54AwO7f0+0Awj08KPpTJOa3FMVUjdwzTFjhqupcoDsflD
aaDEYbaixLdrSD77SpxlA/v46mCC92Ge6abQATOp6MwtnGLAlY7ZrsBVHrND+kh3
zWdDgvCAiv3q7tqALfb+/YKuZPFcPs/eYsUfHS4gLGvBwfZI9s+WRmAuNDaNg5vK
v/Ge0Rf8TIctccG05966gPdngmN4pS5hXmO1ltMFeH3tX5KOXmOYK2fKviVIriB8
J6+xT6UtBuofX2FgHRSHtSio8OkKdzSdgJzAb/LZjMZ0G9NfPUQE2lBgcgZTsJuO
nhjvRLsPnXbXAs2nfizk2lD8tzId1+uviSY3q6py2hHmPbgsn5t5D9Ayhj9QlY7N
8FC6PINvYCrPGDr9Fr/0xFv+jFSz8bLadWoczBUt0ltIiisdtzYykhwGGnhk9Zpt
sJH38JsdsjQcfa+vlr7l+BhSYLiQVufEWjvAovrengVjnkQMEufzwW8BX5Lv1tAO
/Ecpl/XMGmsh4XBkeaZIYBOTYzqlZiRNN1jys68SaMkNJQFv3lkRh7F73aUSuBFl
VBXy+K7K/SVR6/LgvbJuc4Bn+lDYmmIE5DJI9N7CmU8yxXG9uYPa64qMPL5N34hW
f+wD23Oi2/Ke7yNiwIuoByi072mY51u/5B54p1lwowyQItYjKA38X6DumkZ+nWrK
lKRssvMhHbPUWwLLlaV7MWj+RnMwEoCNMxGIcqaINTQWIs4Ex6Zp8HDS2N71U+W9
bG47veRGc9mskBY1auVO5+JmjS1WtorYL6FSrUJNscjD4eCPuY7TD30v7UkxzI+P
HWF64fppCcB4euEXYyzmXpUUXV53ReVc6ZdSYH2CIoOEBlEBILU9gVLtAbI4sC/i
Wvu/KiVB74STGF2ugxIMPw2L65HX/ByuBYs5ll2BzABJMbVQlNwopINspGlupatv
OzjmiqXlySt4g+Mo8mR/kTr2qw0BMoYFgENMLqmbO1hqXKNFof1FMr7mv7bPHPvV
ymy1AItwD7ax4Ez/OXvglQa5Bn1NATRNZCy2/MWSvfD7aAheXTJbzgMTWltJ9Y9q
AF0VpK0zu7e9A2GczrZNBcN/+HmNlPXoMrWcYBqu3RtBMASID7ufePmjpl+T/DHy
gWAIG49nf+Xsma2k+e8+pJ2+ir8hrAGMzGgswPLXZ/swSNhw1xioDbWP50zJg9eH
qkoq7U+Uxv7i/AQPHQEOOmMcaspA0kj4UFAPdVSQa/QFg+apnhmj3aEsACULdQQm
Ge6QnSPU3uteVpZRkiVYrbbbvN8li+UkY5Tm19tpVjtSX3cDzlgXeUZpfcHLpb6c
67j3VSn1HTmEGRdr3j1eOX834FJb/NEA4hiqXCpxiyyaWpDFovsMT6wtWVBgVBEL
UtZtJVNUtx21V4bjd/0lMbaY8HCfnjsxxkSMzT7vCI7Q2rS1aMzBA8dVa58bmLU7
QhFKtTHNHMsTHRuAGz2yGjSV4U0nBYyLTTM+gErGiO/bF0RRLx8CwWvvZ9TXS1aO
qA5TabDAsIi6iGK4/fSBq5UJRqOVRHNqbDvbARKB078gsR2vHi0HeGdh786ukCNy
PnsP7MVB0BttjBEqAurJMSJjPX4Bwz04+W5V/yRUTmNClTuB4fkcxLxS1lMHLn5r
bMTmwINUoY3lLG1VVslQZIFPj3Psk+d0SJzMwziOB52/ScqzluvD0uUkHP2XhjBe
LE8q6ykKKSj1XH1xCrONNgT7xlIURv1eimnpU1ksUhni3bCPC7EbzYLcBwsen29K
VpJLcss7ULi34ht1l78lpXcKc5BiV2Wjex2Mh3JPT8/XJeBF6qs5UC17SnTvaORZ
tCKeuneihx/9q5VE3jzKyu4eT4++RUnxSfwGbtOkBqynC2E4j0tS0ooKkBdAVLoB
wFSowYQ+TGCQZuVJp5c1pvr5xVC4z6dWlHaPIsZIlDnR5+rvGZRB5R/6lswc3Aqm
4xH86jTz+ty106gM/flvL1inEuSq3lJQfo+gZNhHt4Oq1jEKJ64iF5GE0wVMY6bZ
36j60+pt2XZDPXS20B2YzDZaMAqt7NSZz9PCz8kH5+ehJePFoVeWhIzk63CT9B2N
4ZVBx6vw58UCHiq0glwCPwj7y+nyJAVRg5vvOSrm0PBqDh3HAg7E+iFVeJn3K2pU
HmB100LIf8ET9THhWnMZP+oEM87pMGa1P0uakbHj8Vm1HAVeUp70y5izYegIlKIh
WQvOC8/lxmgaSvkvMYJveKP+ZY3kb7bQT3UVoQloTTXe8vK9fzv6v9awIUpQvYhb
ORuHB9Ilk3HKV811eeCetrPYhNFhApQjtfwrPK3BjpTNGF9MsiFm8QjHfPZOqeaF
4LZRNXt2VnQd57WINaRJPDmJlADDZ9wRFiIwn0Y/m0NyLYOBrqrcs54a6vWJPL0q
YI43WosK4rRU8eOk/glyWVJ/gNUUI17o9FIWz4Z1WKIAIqY86PXtQHDQ5FeP43pP
thhlqQM2chNT1MsRdUwIHVICM+Evhn8yTta03UFRdzniBpiJgXwODF1XZhL6iwi0
7c7XKOckp+rB71E/DXl3hWBWSII4JEY39iLRqhdunlc3fC93K8j2ylGZZW2y+7Op
hbaVkgLlwP1WcVDj7wa+hb6/Zd7jeHx1fjJayy8GlsA14T1fRBThDG35FQq1T/I5
6b661ivOK04C7vyXxkYzqUzIxm2q+Y2v7+oGS8CxiOG6cAgKcqmbztyVbjNaQkiK
NfKa3xRTeJeaWwrP2aHqW2ZtgVYDfz4J79oNm2Dtobs+THBCAi+b14pc0VCxmCf9
Tja4DnvSVcWpXocka91WNNpTBNRTyQkkX6qaqPM9zTE/TB5Yke/Gs9vQMmtxBUmS
KFATCkKtFJp01YxiLmV59JrPpxFrfUt8rV5ycLgYFIib+75jEQVREHXv2O4aisO4
AFvKr6Pflrww6iLqy7XHYrpKwuOZbVCYyGv3S1i7iHCnmqsB9AG1aI4WLtr8Lq+J
Og5wg3MuBEJy5GRBrXDvwxenV0T6vUp7kfgOHMX18/1qMhl6fFVGu5TvSfh2MO6R
irdlpTb2x+m/TF3ag7SmRSC3OR17KG405rytKFaUQsKRpV7o72eX2SeEPgPRW2GI
sa9F1wrEzmJWbsQ9BffhbJq/lCBW1dV3xrzhYMdusI0QRl+OzntJejtM6RrDxn7f
wiXxYy7BXC5gA2aWF6m3ncLDa8un0FWij+Pule7EEhndmZ2B9YwXcM9jDQrGbhzN
MhJI1EHWas4kcsj27nyxHOIxANRbUM+GcCx04rjGS8PLUjK18jp+QUOZ6a6egaqD
hVNNquZZcTD9mJOP1FIGyAhBzL9SRu3/n1rTNTHjIgjLwTpdu4I7J+6aitAWguR/
ShjwY+iXfWWIG6ZMi6DdQTv1F0+rqgvi7z/SA6qjcWKPqguEdnlKSQbPu7OWhu85
ExKKrcYLQ6J4dc8r7Bzuom2b56ubuxnsXlhpaBFt45RE8Fk2HoiJUCcq984UQUMd
5j9qPPt1bxkWRDkH5q+MgGM4IleyD85KkkXeQNQNyLqqLi7rRXnAPxBt8u2lvOC/
KhbD1ECVCa/N3fH3cBKtekmVS6kGbKPPLm9ccGquSBjO34eadfBDNfFWVi1qh4FI
kJNEzZuSuAiMd2A8PR8OCw90zUoEREAr391g+ABbROR1dpw/M58wOuI98U5anJww
L3AmsP+IQnDAI6fI2uXG47td90SE3TMY3CMU8i9Pme+cawyLAGcp2fp/jUNU/lrs
4jeJDnUxwch6/H7aJyZ+CJ48UTvXZgnaEVJ5p33BHgBb8MdIzT1HfS6Mz8agv0TH
EMHMmhZtF0/xeG7nbzDH9oYmuKsDDkByoRD/OQCDu7U9Rv+11yvrqYcihfPtxIzN
kIWbg0BzzTyHLFrknCUnBZWVz1zXXT4A6RuFjxHCxL4e27hKeos+25D3tsYlFQiN
EZgW+1SeS7OjxbvwWQSIa1neGgVqfFjLBHNVXrttSpLefDcLySIOqcgA4qrBUyqB
JfAth7p1TeMCVyDTKXkqIMOoU//mWNHl11c8hUcwhJRQkcNZ/ldISRa3Xw9NiAGa
4Rqq486YWhVl7lGYK8U13aWUYeT6LKa7nxDYKXrGaLyBOp9AvR4O0dhI1blPZAH/
z6eBKayIIYWvyu/J0PtG4KjVHas6HReq1lxTRjCW5edmZvOD0YqQxAlxvBHXz9H1
uKyieKGTn6D/LO4EcFC53ImaH+ImN1Ig5I2M3EkVR22qpBIKVihGY7P6djdPbJHe
f6fgbF43Tv6fZUHqLn/fhozU955q/ExFPZ8mcUlzKYEcq94V174yD8qbcwjVhgjc
vID+L9s31hnj0mBQhDfvu93e0BTCjze7ixsi2jVHL9am+AnUucIYv370WP4r2g27
sq8PQ9/N6KNQlAEeRP3nrFeE4VjCaGCcRCHwlkJpmDeO60NrVkoc9OhoNtziFFhl
9e4VGbXQRUHFZT7+oiCDyRsdvrn2T0pdqeoiFmToQ2hfCah6coaAvkB/oV6mrehS
oFRaQRVfFRc4X2jm0CpxS8UFvKgzhDMJG8/84ZeiujvyXMV7762gL+mgckLb93jX
35lpr4MKH/IxNPVub+IBMjgP6elq7936sMVtQMVBxqRpd1Q3lCQFZu9stXw2Hl2I
87bPHMZh8S+c4qN5s8CnqjTjTTKSKrGwj5U0A6oHGT2/E35MNDa3wRDpFMWG6jlZ
I/5S6w59rnhROvFXXq/mbZB+3zA0OFMka6JxHKp2fzl+oXhIcQ9229HqS8MVac5s
FDD/CqDP0rMlEC/7WTocNm+E8DXtRq+1qTtkimonZFqDsI9X1PiZsRqIEGn6lJ1S
Y4epjOY6AzdOHBDk2IuQhkfDG7gxHJUAmY0IOjaWlDWVio3x9MfrFNBjo50He5kc
fiVWIg7zZ5X/7sOh4WBL/2bQgSmOcxxzGQY4G3gsFkDlNOfpC8upb6M0miBLvb7q
hVqo3SUs4m9tYGULTMRtAyBxKYoe/23gBWpl+UOG+hs3f2QfPZ4a6JGaMKo+C3dk
6kcZ0+VtMUcYk37ZNKsEvDG6wuTOnZGF6gSwEiWx1HRq1IcX0SaQ1AquiXEdylI0
3Neb4HWQXl617tlLAPaMoYIt5Juu/8u7EUpvqMPiJ7QnXKZPlHgsowqQV4HYs3Kg
fo1KpU6Fw8SkoFfT9Kzjc1MilCIaPtMBF5bqp/ItcYOZcRKHuCUQFgX45k9NKEIu
7hJ9xHzc1WUs8WnQZJ2EBx9W7lfil9w2QhIFNSH9zc5lqb+15DQCDA1mUS7lYxdl
T8Lr557vX69dsMa4R+MM4TmmKXO1GzTQ6WmlgGunN8c9e2hXtozz9Zls3Mu9sbGH
OnAxqKHAQmoPqKaXz328/+sxeAAk4MNl2+0SfmpDJCRD/cujI+ZvK/AOne75QOZ3
J4Smk0tu5KGRXrrr6G7aYALG/BAhEMnxdAVLZp5lIN2hSdUz9vmwvrHIdGHMBAiA
HCZwx6WtKmAjwnlHIRm+T7H6DKBkNv0vqAPB6LeSlE8BccOLUneFw0oFbl1l30n8
YmNfbl2a4JfuKVFYeiwMSQtPdH7qWUauOmC0ro7LR2mOysHO2HIUNOFGRcrjSTQA
qBhRpIUF9XCUiBxOrEJVAvOhIJMgy3HOSuUYFPaM6ILFnotGMB+QbOzGL71Juy3D
R9lOF9gM4GH7H07FiSieKQuOC4pfu3Y5N2D26upWqYa2it4tZYX3f7e+5jSTJ/sa
N7ogSjOR0tAnPij5Ti/J2NvSXAyK3/YuVYv6stRC4PCVEQe50fOHrx8DPg5OFNaB
z3OlPSnwjAP5+JlmJM5QYE2lZ6trYiDAB5PGBMLxxbJmGpTWp3v+BRTONozl5DyH
FxYZ6doFkuFj0slY98KLpMowExBdxwK0wa7SNimf5J5TuCaXXzBle7/8R9kXJC7a
Wn7UA+Q8lO3TaIpi/55jhM4hiBwVVKpD+uNC7wI4HyA1amE0H4xpmSDxW8hwovJ4
/EsjGK8sVBhTvBsTHlMJeyT8LjMwoDHYL4LyRjRchdKE/qErldcFP/ZKOsJ6wYjA
4rj70fManShhC5kG9DGEkoumSCZ4y8AXkfo8OfGryvVgTeoM0ZaJwyYwpnySMR0A
Y05SyT0Oor6/UChtxnYNYM7sa5GCwMkpUtySzpYaPfhkLFjaa1wRl7HRQcQrRBHq
2z3Sg/GV8cAr3H6ODAagf8SssdX30kLpTjMpEVHmIHlsRy3159d+fvOqT0lk5lv+
3fu7fkKeabiKcocDul8ICSdR9XxKwbGOXez1jdw7cLOuBCewzUXYEActL5a3xad7
LvHbAxuxcKdamL8UWcFTv56luFffeOd9jwqX5oyyPGKAA9R4MBCe9K5t549woeE4
F4En5P10tOKPbvIbenl85oi4m9ujn2SKmL+g9JUg6lcEhFy7qtJRqY+ZhlosCiRo
yicgHvq1o4ggf6WUKTMHqNcmsvjgxKmKDQZWAM6/UsZzR8EXM0+DEmdsAgCJo6eY
LCKE0R0v3wMse53iI2KIBehPBHBhv0dfieEMKekZG3TojePbYV6fm5ZP6ObiOGDb
8R2ViLTKNfl5cmWQcrYglXAa7qyRqkUPkIbCC7lRRfNMWs9IVx3ClGPxt46UOWoS
rJ0uXnXJP9jhDQSxJDS5pAN93GSYzTXVlpMxvKOiy/NywVYsxfzlSh0HNuM7GA/Z
URJcHyjCybcuU/ddpNehDA+OSOK8G9wENqRpei0dzqUIbJAM2plRmybsjsq4W/VL
X4K+XunXDK+1bYOaXjRI1/vwr3OrT+Uqrp/RfAHDarkDG9KHNsy0OyleYIr68ysx
XpLF7N30MA+xWTP4yMC4IH6pZR8QcynO+votklI4zgcgzkWg76DLL1e5yjXsoJ6E
eWhST+PjHH4l8HceGCkLcvtYVF4cqy61AR5f95A2Tjyy9N9BjlHrO1jRwdM/ACKM
fVVkkCXxR//F1ZL+Lqj8UyIBNg860L2UOpfXhaVlTBzW6znSZDtMZkJ1Fl2sacha
2esNWtd3EQmMK25DQOf6sNAw87aSl1z0XC8WV91n7RYbfxob2PDn+ZXW7OrduGTD
Kf3pvUs9bRkIBAFh48Gpi++aON3EPo8MG/+Og8xsx4pP3hH+vvrHP8LH/D5zR+Ad
pSZsHdhNl7q2PLJ17QqCv0dlGMJEmAhrtrq7UVg4+TQ/vhtRmUV1JrIjurpE0/nd
OEf724iAIMW8eI6ZaHOWxpI55NWnOyjtQSetViZLaB/KyXTcZnSSkT3kKZf3mg1E
ddyajzYaALTDwLH2Whp/tqHD8VK2qHaNlAe+9SpvP/7uzoefoP1mm7RruasbgN6/
PoY/7kiXiwYkS/94EnzEJJaBdCXwFT9lJ6D1ne36XEcdhCHbac02I8ZYlSTnQk37
xMUoN3eLzRW9deGITozR0kAVWkSH5v71H07/TanWMibkHVBgxEBKkyCSFAvW/4Kx
MfEDgiOo5E0/ky+hezLRYPZxc+/JJUMydeoOY3boZC/AZbhcAxVqlGKkoCy7XywQ
iyPEQiuNZgyhbWHy3Av1PvsEuARNa96Y2C5a+6CuWaX7urTvyquoBsfehFsdkp/Y
UILoRQ8TTmCD7CJopJbTVWZtkY9mmKcNHr7CfMT9P0EgLq4bqISjMTmb6SslS4Pe
CI4gNcS2uqN598mqfWFj0dELqWb0wMIM6w11E9UMbuw4gDbUh/+FSoiGatWNwA5/
yI/hhvPHTMY6M3HmuKMnZvbfusbafZKCevo568z+hKLNIqHQf6wAEPYDMEbm+eBy
tfZKMoFgMZwNtRDZGCoIdZZGZ1Um2esgF4I7MG4BJal7SeQAf6RmRdQucMi7Bz3r
E6hcoEfZKDvjYr9dcjn1UZLdy4T5FY/0e1wPgxKOtYf8H5hLJo8ILzpQWUiUqTFx
5t5Fx4d9AS1ruO+bjfEYx4eG3tZVjyWUPOM7UjQ3ll6mN/y4gvm0f/LWRUz2Wh5U
DZ/MHSGjLoGQMZH4yeKouxwgHumgTYWfKaIvJqLnz5wPgSgN7/OShjVeLDmI/7oM
8958qMuqZ5EfbwhDBPnf0dEGupPLTWqezmJjOv7WvAPBFLu5roqKoJLkCbmT2MBZ
WBHSZZ2+OapUU8rbdo1lxV6EkgtRTjcKB+xvoeYXnVzrZAAPUF3bJc2Sj1O9wSf9
p37YXp7gi/lvcI5/aX6Bjo74mI7OcymxNYcv0IQq/sEm/79xbRuKp0NSjFfDZiCt
PEh9SqdjKH4hxhbxd2SugGovW0+bies1yiQbx0tRVWY5SHZ3TBopOz0hIZMu+2q0
updSJ6QaO0yO5voT01rTvNcAUX0n6DCB067p6abAJn7ig84u8RbXwIQr172ELojl
rhaxw4lzjSzJ1o6Cn3EgJEREB9oxCBcLCMAJTdxbJbbakZHC/erkzq+ERinVllhn
RDN3kgzykmYmInf1QY+Mx0CsyMxBNXOh7TOJP9f8rTR6x1+cq8VxDpPpFgI3AQ0l
15F71cFR8Hx6b0zrKdKnTUO41/8k9ts8mj+7hdDPj2/ayAMF6kz/HfLX6CTyUp6f
YGdEjaX00Bavvb6Y4tZeY9joomsqeWfwUeL/HyeJ69kPgz5AJx3e7G+kVpPINC6X
XBJugkj3mvkmxnAX0kgOUkssvv0IE1ppePO7okWgEb21Q+z+qdQRGJ7je0Lu3AgZ
QRiyCnBngr0rtUa3sPfxwEqjDaz+kXZsRHl5+eJ5PjAhupd4o8VwknXzkifedA7L
G8MjckWcIpSjw81TxdWpBdJSNpqDpXEwZFJCAdD4YjSZTzrfkmGBf+IpmrT2Ioom
MJjCuAbJX0h1JIRbUizhwauUoKAdeZxVRrEas68evo3nxnwK94lLPb12xfVMwTRG
a3ih7GtbJah3chdB6w1uAN5IWeyyBfPPZQ0I4vJMDjJOOJD/r5ZPgheALrs2QCQ6
sHKhZDSOyvJ96DtDN/rzRshB85r3nUFPf+f5dDRrzTXmlt5EKJQUl6d+39Jhs1V1
OIFeft66ASeWxfNu/l8Cu9IaNW99jlLzY8w+0sZc++fqtLd4/NERLaZnzyPh72Ld
EYoJm/6tHhNeBXeNiZeNorbfD6/d8HCoijE2owsDedChPKMvQOc925Bf2byZk4XT
LvuAngGVWFj1gmcSJ7F46QX2d5bYZxuOkDh1uf5W99Hd1PJpdzmPBRA8gRI9oXck
sDE9vSnQEX3860fn3k8AUf2+jvWC5VC1ZCCDaH/fbHg8C+P+KZUL9mIl+fq5kzwL
n/5P/5qQQ/n/TzujOUaeCtqqsjk/8YFAG2hzUCb3/k12keiY8EsLlu3+nvg1KO+P
qzrJliQNWLc83GSmB81ExG1+DeSNCGqzjIYdHTXvUsdUqmLBIMJRRdai4yyEmAOO
7wIcQt+fwz64VV2XumY+LXIZGL2ot0/NeURePWe+H3ydaHY4H0swvvYwYCpJyuHU
CXVWZwbCK3AACloS33uobF/eUoUit9q54P06QpK/44NlOyQrJHboWN3/XogHsYbC
JJgoAFJPboxZuirScw3FvEjEMCOw6bkrMqu+4i/cQIlVJIwEzqatWgb+LnlcBYrv
aTogrJnlX4sdGZ/R7pk3PNULBsel+Cxe8cL3f4NNvDNdm9TcP1wnqO6WBysKfkj/
kkJcAO+42245ScfHell+SgoKvq69YR8REy5c5r3eSRdAXimgWkEw4p8pnNf8cIHu
075QMrAOXu6SZHVB4D6RQ7IjRlgxD0Ke/4Y/KtOaQjnWxqKm+t5VYCWysoDJboJA
ZcvRqxSG729TdnmpTZzg/eUgEYEv3mbhzUxBMV3KvjKdRTeDh+mubRMnkRgWWMfb
EoCwCR4YRUp5EedhUF8OhYT97Q0clW4VfEwjGuY8uYbS6FgbbvoniZHBthbxgQCw
LQaECitfVg96YLeH1sISr20bpHgj2dTJwImyllBDeQlyUi/gAIpKBY7IY9Zgr3ad
kw9jjwb6Ef+VuaqNSfZ6mcLiMo0azxRG73VDuj7fgk9jVWoB9/a62Okx11DHKLGW
FO/oy1M78/Q4D4OjzdYQ7XvoSlZacO4hxWmrR/uCq/S7I2hQpfW4uY/7fLolmcv/
MeABOn1hhQg3yQeAp+8ePapFR8M/BQoRdmxKzu8uIc0pkfjnYZ2Lc+paD/vOU2ki
ZwJhSlz51p/KfQURjS8ilW32EhXmlybry9X/fZjxRI0lXIJD57ZZdYWpFA3su9ky
fRdQpSI1AfM2fKVixdHCzZJnzK+SDsoNLF62v6bIbXOhUOIh8W6aN/2OtnnEJ4Zp
GeOPrWrLtXQeObAGk/3CRfA7YSsxpLpHRiId3ryxmG/ax816UJ9Dh/jXIlkU8NDt
mKQ4eq0JryCkBplJAVpiKEJnFK+kvhII/K58CqYQFRK3rE5ID77a/zg99a/DIW7A
oM4L99MsJi/Zxsn4UWGDHmRsQXAHP6gVVAmV8GHRWGETDsBayim8JTvwt+pox+Hy
GWj7wsxwmgo0Arpp6IK6KFvCw+2iYpdPneZOfGsBm3R0R7npFW10743ytlEuLvFN
lwONVCKHAWr5JMTGiwIdUYA7z110e/iejsucGX6keb+zL9SqfQopgDgW4dRmVUBx
MFOirv9dlCYREnbgfeYtXTZAD8UIdxxcPAvXygr17w6LMod0851L7K3ErcpDbo2K
ga/CKceqOhuuME3DwtkmDmaxYrSA+ryejuQPjOt/pp8RixvwoaY01CpOEUV2OwGx
YEn2/1PhoQnPMw1FHGNN0LxHMYZiVNCsRXaPxt/gH7NaCyYU6iHCj+eUbumnLe8z
91Lyneo2qpH7pjhyfzyG/X5ZpF0Tpg+UwIZXoAGpZGXWTxqAIoQTKZ63U0CHCtKM
UQ9/2vscFl3f9ANOIOCg++lG0zKluLAtRNH055GAFxB28ga4AqdyF8aJPUQeanZK
w5c22dezGJT32xVAgjG5hPqYKKSWi+8zMROqLVtHa0bM/m7Mcocs5cvHmaNthBXD
aTaCBUcePvVNaFCj50/cbc7GcXyGQo+EzSHcVyhnpSjYK/TbeTZ4Dd2XMdSyaASS
XzypRxGfAQ1HR7rOsGP9UzZr7S+2Gm4laKAsO2OYuhBo3gNcdfRuMwwJehZHWEEE
nw8j4fV1YiQUmVzRGK4j3aUXCnnKDc8yXmBrhGVU9JcNdQV4Yh9U9bE+3E1DMlKn
xGZzBaoK3xLGHMbr5sAsuPlXlkC9Grc6EwFXxkGA97nptGgr8dlAIafUCLr3h9+V
y48+HrrJPduEC8FBTMc7jjUmUq9rIHtp+ybk8jheBWU49SwWB2H5ZX+hETiJhNWM
XbCDNReXWQ0uVUKqafiw/lHIHbccnugY33/MBFhUbpVFQ9TLSel59jUdAjee56Vf
Tonu4C+kUcz47nUHhg+ZCJzjAhbYiHNLiMmXkvEDLg+7J4ajy2EtyFfHjpfEYsLQ
ywsTu9I+H7qYxlT08VOQO+LRHZTOLqrLbHgl0oyTFVOvMN+fB7LGg9nJK1PPeEdZ
GzWjvcTRi+dvMEzhuBtPuT5PPJ+oYKIj9Sfi+2afNpAvP59hTUJyKJX59VnVa/4W
ExnLrzn3+6038O0qT2+/8O1eHJg1RRBlylnu3kV2YaiZd2w24InKdgxVeeQjTNTa
bHcZB9Dja79ThDdcM0pTODYJV+kSRIQbcO/a3cjFyYIezsjo6WvDCz6TQWLd5Mzv
4MjlMYyCUqq3BJIKp5HxngXEXWDN78omBciHjMiTGwxh1r71utmt8G4WnNDC9u5U
bUQNPHfkanpd20D8KiJivhP5JbV1Hf0/fMJAbr8VimkiDyDud8D1FfcNzMeA/RXv
Tiin83RGLoDpCUfQnPRialvCIfcrXaJaMi/I81BGwNtYpWi1HmsVymF7U08RheqE
MRQbv4PpAeY2RYozd7s34HS31rRRqzJL440XUCFLzO5hYsnR6rJid6Db7pWoB8P2
MHpLTrpiEnwM2sp9TOOXsyyFQZipR0S/K56k0B+MzYPIek+ICtypwvGWEdMj67nu
44Wvfo2yn2nl0va51Gc9O2XoCYrmXMPVyJr+qAlfXOg6LgVY5iuIqcYoelfHLb/t
GI85gT+QpX2j7UExBuvfXufDPjPNwhlm7//brodXGnAjxoCDty6q8UFgoPUDur6C
mvq8Vp3tq5jQT2NdnzdYa1IKD2eJn1b6p0nK4/JqnUAevz/BS0wecHAZNO7wcZDi
3H+K8lOuPS1Xrqidw7vBRkAKE7ewtGNqHCgr7omMDqAL/IvfEMYk2+hvRtMBM0yh
HOemGUD3flqRaLqwkU0MnNwVY6fBq71vkaWPX0ASkIEzTUGjj3OjoLmEOyS5ZWNy
LmQNA9vE+KukwnRbSEjdns/XnBEb0T3PB6J9qj+Q7ePC2P7XvDsjvb585d9boncA
GFjs4/ZyA5E21SoMVcJyTHI4IMnL9tHqRg/jCURYX0MoRw0DJSpb5q94JllSnhYP
lL6tnVdvuHdXx2ymjVZg7ed0VzCz04/2TMWxR8jeI9fNBUeNK1J30Vd+F3h2WOsk
CwLvJBIVaLXSwZRWclwRDivLSDPkuO/kC715F1tzjo+R4ap7Crvri/KxmffxlFHs
yIqIH1y+wR+JTtU1aANCj5aB3zDQwaXOrKzoilBGmlHzx/X/MgrS6XR/STOv73Oj
LpjI+NA/Ss7lWo6dQPolaQtM+KvqK/OFBI76r1cwdylT5XsFiyGo7QC+J8FxgOqT
E7i9eePbb82yrf0NdpjYVh20GRniJMGjnzMMZ8aXRkTKDmV8g1Z7rBxbcGWcD2Wp
DIwPkEhk5vTeT8iJx8hbeD15xMibxQ3o4QY8uZBfuM/YQ5N0AvHW7RV/oh128gpb
9NNE7y92T64uYzelj3jA+sixKX/B5mjqfttvZkRYMuOaRJNZJ+uU3zvd70fO0ikn
VOjY09ToDKS/7ngMCzua8XQRKcQcPISX8vHJxQV84mJXMNO+D5/c3OOgRGoySvmH
dQtWmLeSJ+hhCFmceF1zrB67QZs3YNPtj56d9kaVtkcUfXoX34NLkWPunRbx4EOI
Jbicgf0ehEU12zhARjrtdCrrsjmnFGYGR4lr2eIC5CX0ppwA2LqtWwgfmmdoiOun
4BVKWH0OZGJ+1cpw/pibEMdgsgmqmJQRaqSPYWNvY2VH4FLB3W9gfHCLmRCuEFp8
Y0Yd6YXbWo7dWgHPORcvgWUYHasbYoKSCpTwzYJ07xDYG4UjjG6jlbggyieStJOq
znBMDIfyQatLKWiZDIeE0Qj/A6YeLZDOS3+r+cpMjtGstZXaJelnJgHz7VFB+5fq
GWJpGdM+Jv2UnZG/TQZkdOpPzM2MJqqsig3Ukd+8VQ2gv0+jSX8KenPqlXSDbDnl
MbF5CVZrhJqHHTHn4DymJ8A4RMLJ3MOTY+hVmGPQNGZxZMQwXUpvCXpLVMb8qzBr
qwPatGDOKVndoqf+HMaC4B4dNR2mIoHQRDY9qF4EL74pd6SCo5LQhSJod5Dl02gP
wzcb91tFRkWEXux7zGjjOnihGRtwZeUQWCjduYF5lYVncCgj5qFyMesoTHqxbVCS
aEyuHwrWu/eXHRc4ep98mxsvQBs7Iv+tAW9MwnRUdOtZDSh6IXza5/lGkO+cJZO/
Gg4Kinyl9e6RCWw9XculMe+hTflo7HSWFMMtVeTlxL3GiFFmIucOGTsrQZzmB/Ub
HPcmxg8DLZLqLLe7Z/cOSN9BMzBs3PEqvzhETYXL4C926JWhJ6fvPwB8t9p3sVtn
bgYE6n0sSTVwgWX3pu5llhhCvGG5hapRQHy7jvFh3PlU8AzqeipKbSKuQ1EG+YMu
k0vBK1fU4kyeTAZlewWPMxuoLPWF+IsLYQrDYVnm+Oodvji1K62wXl+cbHz+OiMJ
55Fm9xOOUIuKZWjxgljz8Z6Wgq8sIFd/4Gs0ryWFVmvMVnHf5pWk3AVR3ad2Voho
MTZslyCAmDiSUm/tzkKVcwuLye9PNC2IQNoK/vI7ClmZBbJ98A9b7IfHxG8iVpvk
v+lzw7pr2W1qT4OaZVP/xHuWRCzVIJ4Qg6+DC8faSIQ1Pdjb8ecJ+F5Og8gyAm/V
qG3YmYMOOSugJTQgDfGII20XgD0HJPb9kbcP5yBF/hv8bS9t1OPDwlat33YDKDEU
43L5Hlig0jid3kEcfN6q1/UW7oxAPTGNf5cxSRAqcwU0PHM7awilkoYVybhNLtao
Xb8+uqX6IU3Qim1pGUm4A6pOoREE4KqZUxBQ21IwATo3nro8i0orlQ9eURcE7+lb
AvgH+DGI8LdiJY8574bPiv6liBSqQLf//SK3su6sOF3oQxfznct1xodk4CDFw5D+
O2qgDTTjl9OtYX8Nz0cXBMrEkVe5Tol7ofMQ1wkngyYIp6Kr8HDdZowL8Em1RjAE
gOW2QpvXvcVNmVbynvbsHnx1Apb2viVU9AhP4vsM/TvE+JTwg0WnrligQtjTKJWA
tq2oahTxoV/xoG3JcjR9m87bfsJfqQ84q2q6He4X3McQZUNSAz4oUPyeU/keE0pf
ewYIeYmwq62k/xU0KyKL0VmquMcVUQOXWNwaHPpkLfSJl5DxrBb/sXhplsqi1eK+
9ezZcekGkrYPRtF4M+uOb2nZsTufY7ReJfftRg864ebXhvjkXHVpTL2gQ4BVCCU+
5p0L3d3tyurdHo9LzRk0pzWZJLgyuEhR5SHbQgXngff+5iyvusyAKfngQWaJv+yV
iIy0+yZknnaIKaeXVuBvhn6LZcOMmTf6MK7MpjEuzWnB5CpH5/aq8In+dd28wi9q
or7OG3ljZDG7ExnZvUCCyNkiwijVBBz16n2rhpXX2vN8x6rBzs94XSMtr5sK5XiZ
VstXYis/ctSfmkfgkMKoCvTYiGTMG2qFo55DlP04WayAaEsxSx1L3BXuFGn7vKom
YxRxoeN6zkDfa0DsbXiTNAOYcKY6yMM25AFUdmxB6YMuD0GDPEehz6TpKg5wefAi
aXgjTpkIdNByAVel1bBVmo37556r5RrvWN04D5tBmx7QuBrCYTC2bwunUzSfjiLb
uQuo8AOVI5ohLxJbVfMpoAZAbAMweg8K5AcWU/gcTq7x89Yn7HUdZz0BlpTvjyd1
viqfZO21nlM9QyHBoACCGjZHKVLRUY1CxxdeZ3v4ivr3HNO/dNt9x5z/Cds52I8z
o87I97s+89+E443ZfxkO8dgLMVZsI6yzGzttDCVb3pNQugZEE2HudTfbGjeds3V4
V9vIlbRzgrxAj1FP+Nqb0MtvGzcDik5tP7+83PZvd5/3ekEpNlvV0jzZENthm/l3
R3XLtBM1/onatzij9do20wdTbpXiemyWE4QTu1KZ+Dju3NaPhbmFFPB/1JyGgcso
7A6jDpi36azG9GOi9ZSDy6BT0TCVESqGLtaL9CtI/g4tERxbEIzQDaFueAvIr3Yb
6aC6SUo3YDq50VZgg8mE+bxIgQFwQqBjfZf0UIJNj+3OuJ3kXHa7du22XChgwO8l
UD00CckJEDhVCFdyIfcmn8jaWQK4IrK3fjzuSCEJFjLScyXNwzgUGoLNtLjnrCCD
9cydZlfidGKmSsw905A8oOgc+0tR2iRf0idtr6qIyvYfBw550T+BNwtkivCMtVVa
9bi62xViibJLW6nl7pLhMB3YgfcnALCrtxCHvKugWlWq/Kjub9IZ5H8+ZXxA+E9q
Zv+1uegKttLzxiga9vnze4osv+EFlvx2hUyQTtfMqitJBCkx/hcEidritvk+ae+h
4Qif7+Ka9xjkZiFHfHU5I5biInH0BP1xE/HKw6/TtrBrjJRD5wGJpLKCi2+J9CiI
5YMyFPxs09IsFch3LIg64SJyzpdhFSTT+BDaSlxY8qPUMDGDoDyvxfhw6fFOVb+R
vzoSSeAG6QXQpuJZo0AfDeWDrHR9c+KqlaEMQynagH061A9OMjlG4Rz8x4suRLip
EGcvFrSUtuUkVrrH83AJudGmShxf46LXGeVxg5M9RyD3RmQ3vuJsIIWJXpF3KGfp
b5NIxnKXf4kSvftaagBbqpUr6r4xnE7EKLVB8qepu8v8SIATRBcP9Ab0dIL8q1pT
ZLBq7jLd8nZUhPMz6+5gYDkN5dBxs2bOm/LFT+qg0dDGvMFGW25S/0kTHC/wyiG2
toUhAT2W8pW1orToyFecx5BbDw/l4Zzd6uBrYcFNypPEKm/wA2ry2URaNCR9+zOa
tyw5OL2UIFawRLNmrxmAoFpde+JhqoFdSupjFdKlpnSdKX2qBnrNsQjqpMb2Ei7v
LjNbM8AJoti/OaCxUf3x5O440LLxnTasq1k5UAfetIU0tFx84hzKfbsxxKaRwmby
/I09QtDbyoz16dGBRlWwZeIHzTOT6WGeF/g8jKLE/tXGlyWKiaPEkCWitYrsi+mk
qXpPo4HuZtUciduf9N4xn4MVDbdI0ygNgCC3rb+2AeyBRC41DynEPLKAska9He3M
GwfM2zprarZuRl59MXXgvvdfxRzyo0v1r2DiJbKBltjDl980N8KpDCbLMYBW+NRl
tqmhR4hNLdYNm3GbA+6vBYd8nkxwZYUozOunq/LnydLapGjj5cOARQJTPrOPn4/6
D5NTy0+sMXcXPvrJjhOc/L8SHDOKZBLyQIOIvoqSh519ZJ/vhjLnVA1pz7xsjNmS
QAa2EqypqsaN8I33PqO1SNb3wwyeAuSzuZOoX7j9YxCF1+CSot6LyxDC2b+bnPqD
w8e5ibpAAycgXV5mRCRcKRIuV0NGSCeTffq/F58lR44SaqEJwLofAq+iMiEiPdZX
EQcKd1rkp2RZLLLuUHMckQAACjQzvvE5RLeNPjASwEmHlescxHfOWwcwDXwyrUFd
dArkEvF786953H59perKSNCp4Ospr0DJq6G1mkIYcbslc1dYrxYko0K3B8rh3pjs
rnV8epuQlChuf/uF52YtmKfEit3Vu37fxEihGGdklZQMtSBYM/IbvnqkEBwFQ/J9
OPvT2K3px/Lu1nRDGF1+9UTeMJeV4sdjyTPEukiDp2JFHfil2fQ/52nWnNSj2U3l
UiYyQeftmpy4yuDHrIuJ2TlNWOoMM4ybB53dsmZ6Taa+i+zBQBUTMKedR77ieCIW
04Z4pFV68LxAjzto+xrioOa4hck8CG4u3tamkWByXiRqb98BAq5DJYHQ+plWMetg
C2JS8bQ522zu+EoxqKfL/DHa/hL/Mzt7ZVIwHWDDIU8jgyy6rUrCM5Ds9WrRj3eQ
7ucysQcL7FhE0O02qa971tCDZk/SBe2mzXRa9z2W52GNLk9biMeCodOQ2nZlDU2m
CCLmteHy8zWkAe+a00Qz4Lw0g/iJ1ulyuTwid8OvOkmD9Yp+0xlyi/r9PofzQxmh
Yn5Zv1JLZL/DZX3q3fuW80/mrp2x5Z9VtBcWzqxrFHg1KNxD7cc75QH926T4GcQ3
Dj+ee7SlrZAETwMLqU5DKPsqw0o1Ajw+T/vEWS3zwRiI4uUfatGJIChESnS7G8Bw
3A62Sb5l+vBRhZ0kOxSLWAmjuzWKerKT0hMAfMlHkTaGiwnN4V/76gApQUyIWE2H
ySeRb13GZNQSX5BfmbFH25V+gsHiPwAySAj3RXwGQgUQqNN8A2lX/t4riTcOggGN
/1SPXTbyoo+zMl0BgTYClWVls/5lZvCBAJX9iSPeQQz4fguDSc1PJKCufKG+sPpw
Ndj9y19shKqBCR3/HwfuZ7DGjeoptAmqiFiPq6p1jn8OGxA2eNLwp54ckFbJFN2h
Ipzg9+7vwOgix1zjigZ4YWbKpQK89V21W7vvR0TmyKmofvHnd0d1b9R7L8uqZD5a
dcWP1HDUjtTDswAKM+hve0LltUQgekGUvqgvbwGhENpFecBm2/sMBOervB0rjkD1
50QKLPuwTNuGpMTy2+5D25Jj7qtGA/BvyiwTmfL2iNwNoL9CYEfNg4n+O8Yvssj/
ibz3CnA2Hw027eoDsqSxqcGgrh3zrr21DiLyFTPN9WEGzMCEhitrRdpdAO+6ttBt
z3OvfJKzbyY2a4mdosxJHTd3q4gdd4AD5HtwfNhmQxPAdOjh18wS54qrH2whc1YP
q2TevhV3Z2PyFL3vMjzAzRiSgqh5eu4mdtnvsTbvt+paILYBtN0PZfvFsMucGQTf
ezfllyCTJ5a6yPydOJ1p3YB/ToLfUfLRp2fpBlZrEcsS6YNUvhQLH/LxMSMSNUuD
SJ+unc4ZBSboUbnUrEsuzWJw+MZa0uxcO3cJHPQgk2/+qngDXCP9Uig8bqlHilOn
e/Mb0D43dTrxPMNwYIg/pq58feRIApHJKnyhMMDGuGRb/PG121kgiOsYU9xyahOF
fdurhF/Y6eHA6gAFzJ8ZYyrdTf0l3CsYe6p02tUmhDMlhd5gCVgw1zj7m1tIZqSq
IlVsyGlyaIMwTigQwsoGt+pUwggTQEjYfT5B/Zw139dsv4iuJbGOMKGEu/wTgbwj
YpbQaiZ5scDJIZoy6gbwCPKhJTXNhdoBDnHGOg9rZXr2Iwk6NeZFpDN9M/y4OABv
LZ3o9mrcW5TmntnY6XV0mdFTeJ3dsgS4Ty8FQBkZ6yTjGnPAXUvf9ICmLNjeP+FN
rFLBEBuNmEVBtau4NHsE7i5/YQcw0o6tBvjVqk+bZzCUmQXKGJaRaWlTRp19PHxT
5zHlHng3THzdjVtohyzhhJYgGUk5PTv9M2MzFRz1cEozzWfrwyNb0RrOIpEh7zpw
C7Im3bb5tglyptygIs6G188MDOHbLul/UZuG7MQUQ+UrHGYHEpgfGQbX/KqtufwW
4IC6sXKte987oJN4pYoYeJmb7ZVMvPm23x+pIgu7QaOwQ0FhSC8SB0wUwifVNC9u
PWC06CZ5ATj/S+irWgY0wlyuf/KrGqfYVEGMblcDhOT1/XT4B9LSrRsecEL2MD1a
rKONfVkx8jdUZRz+EBMjPGwwtefPq6Idd8We7Q73xBW6v9JK5SaTdO5NryAZlRnE
3b4wpY4ztTMcgzV8wabC5Wn76fzMyt76qq88MnVkJ3IhhjpCLb4klpymYE8c/Fgz
rrZoBEGBU1XVOPMXzev6QeTn9/yuOmcrnKmN9C0Gs14PNiOwSFvzzvRD6wBa+589
rQSQy8WPyonHzGZvkZcU5l+8SF9ou1n+v3YADVLiaCc7Ngq5qFekM1u5bmibNKxo
QI6adOGX55cfTKK3mhW+tW9TrSakfoL1QTXtEUqO3ctKja68Cd3Icm1tsnYc7plx
Vvckur5aT1h85ahSVPjC9vM9/e4VcFrXe9J9Q9W9TndWQw1yF5K7CO1v1272GwNj
QGEBoHwK8ZrvqrmAfx5YQ1ueZko7tsBWNQumz6df++oc2L3SrAbOKMyKpAcsmvb4
T3sAbmvgn7m5ths7k3ltKUB3HPpe1AxCP1hRxwzQO9z91LM7vDqEkh5NX237gMkY
zC6oeMoroe2vv9YPnittUDe+MwxU4Jw19J3CBVlq4hz0xRUW12+Jo+QEso0TMV6F
1DNp2NLeAEimb8CP8xzkFWKjZouSTIfZYy9Td8rnanyd+4VdZTU4VhGuc79nXxpD
mN+f3OPA5tHS1tmx0pk6oxAdne7z9U07QUNlpxfuNabLCk3Zjled68bpLsa/jwJ8
5DHQEJlGCODfnMscocNqyuyM/9VQHDHp+LhcXsM1QdahoStVJSexuhONmE4or6NO
9RiCkX6kY2nF8p9+W3543LOmgW0mI9WKkckUQIG9pE7rs36qwhGI+/NK+PlXbffd
iPaJJtMeONfIWOBZNuYYf5VwAjgez3DgrECwkm9Y1N3Gq/8EGYjrg3ezotzkWeVS
3+GHVfRp6lvNwBU4xnyUtaEHPELfqZUeWYuiPiMiTJmNFcQMyx5cOg5YhEJYbGYu
gLPEVCBv0xmsMO1udLl079rLGmcCejjjxR9fEL97EmKqQTAaXQa7jPLW6HBtsqXH
SUEYFrdzFj7gwQowzsTkuGdeF/sthlSW2sgH0roa1kSQapHBJgAP1n4Bz5qImDjl
Law1XaLKPENIn5pJV4UXssoOIEtbcyqMzqPEdR99kGqafFsZUR+IsZedAaKWxeiT
+6aMXabSMZ8IEbC3aRWFIMrDYdh/BMD8uDLhdEoQueV+y0HIAVLG0AaemO7+I4z2
KfqJLCdF67ZDh2rKajdQqyHe7eLOGJ2x8pHuC2R2Dq58HKjGPouJixc5CcCLYJ5x
TGQoWVW5ese+FCG+Rxwpxotagqfxpo3jVsssjvSE00FTAJ8PdD/3GSV9N/HwF4tP
DH+V3H/A7sRQPZGQxpPBQwXu1x0n9YSGdcdJVYVCyK4dLN8gm8MEVKd3MkZtkuIp
/GjZXGWxNN7oKJJmXRSqBGlY7ECjaFREF8FG4J+srhnFOipzrlHQH7SROZlltiLE
+yIw0M+oeyEqmlWZdpVaslgsAJwGf4v6w7YYnPCyVgQbS01fgjPZJJcYzFqgZQhO
TY2HHVzC4z3Px/BhUA6zO0fPUZThVYr7+Dn3NfOtMiGP9x0IGK0bnE5a8rxm4UCh
Rrhw/ZESYK0zhpU2GcdA8JDg6Xwt0DAfEs68xml8Sd+8qaGcD6zKhxNaUEpazzSZ
RbfveRL+SHKDxgtIfeWLVC+pJ3YDqD4NhVA/w4s8XMSv8apcb+aqr/gchK7udlUi
xUFdR8rkRTzhGlAYXsd7Ij4I4pQqrYjrbk2DT1+n+ndltPQ/5bh+jvl1OLJ93vHa
0oxim0Ikbpr9FPfCB6ZmCmbsMAxfm24DhNcVdWXaDepGZa/3jiyNmTIgvcfP5qww
AljLwUrsRT4F1E/OKf5qoEd0RwWmNokFiCiOMvSkPrbAhKAX/sd0QEpLXN0oOzX7
XrnIU83lMSML6sxoaKb9AHhphQc49yBYkenpDVJurt9ecaT1IvLSPbRm3mr8Fm5J
+s3/8mg5cEss8fFGAuUqgVcMg7C6p2RKh1EjQZjyvvPRs7BW4mfgeCSx9iAUEeVf
/9W1zdxh6bUHFEcdsciTop+J9fh/4AriV0IymwsY015cO/CsN1/Cuq/jtDmgh7B5
16o3L+kfoH8yN5Ro+TQP3YyhiXKpues5xe5DBqEsJ24g3dnMH/Uddv6fRRbI/G/d
jPElXV8V0s/5tMhdSA3m5T5z4KsgYq2r/cOPS5rkpRJ06fEloKc2r8tie2RvffBB
UpYXZUn99trs7yQEvnptbp9boydzio3KoG6yKPOeRcnRx8rrO5Nyzu1Q2od+BNsr
rB/NSk2u+0So0FGChOls0crwMXL9mTO3pNUM3steEyyWxFWovpqPPZzRq4ajFrP0
swsfWZVuvfqcebUwNQf5+aMzH6T/xDaA2NnVtw+QiAufJGr3DbxuyBsLzdPPfWyM
tS1DbfR+N2RIs0INxToDs5I3BED6pLKGvKs9NtG/gYNipsVQ2Fc9L32pn9ZFob+g
EPHVki347eJSRC5X6IN1d5h5iGci2wg68bjQUe93LJzxK3Qj/syvRYX5mKW2UbUd
bcOGNoWgPnhEBEgQ1eqtu9NM2QtA4Jmmbd/SqkMg/0Itk/jKweNwv8Xl+/INnCoV
6+nGbOKwZRMNKQh1AEOWdIhZxAhS6uFULxVonn0olqxd3KKJGHjakFByIJKVW8zy
Lm2jUV1YNjE6tFhN7FBO5PaLmduP32mNL8qO79w3Vu4N1+pOBVTOsi0ue8Kv8XVl
eft3Jgs1vHh5Quk+PRk2jcjOhgdyPMh0MnmOoUfqhan1HaRoAbS5UXiIDLWmIsjd
cF02RxYOiZG6TOE9XwTAPsQvFQ6SsSVQ0Hpxor0eu1+hc999JJ3ZgvT197UYmIEF
5EnUhL4HqxDRPn2PB/EeARbmR2lVr1p7njZHZvxEwFs//ZsNNw5jBrdrt72s6YBg
fNJmRp7k2j0SenuLV1SO+xxIsNgrFhdrfjNvMeuRCK852KxaskxabMoQPaKjAKJD
2c8Dp6T1cpIHwsnCkOVsZ7NhSZi+pI48dt6hvR0co/5P3Trbl15jUMMW2jMrU2ag
5TAd2zDm/uG99LqYVeCtY3ajxmsa+PYVdiILBDFbLNUhQCYevq4k/5d8h/ZKP3d2
K6bgFgv5Vr9QX1efn8sLjTk55u0A78Mm+oy6Iif/X8OCCmdBmXWkk8QKgS/RhQbr
ZKUztqK6RODREVfu6rp5X/z4Be6zkZQ3gyB17ayqMWz7n3+lPLqlyleqYm/rje/b
d6Zi8o0th9GqxkC48n22g61mz04v49/200msci9laOaGc+4Fk/BTtFVitYp4ujT0
+jMnOmpxOaAvNzgX80OdfAgJBmT2f/W9VRrkNUu1EbiYxMinlKLH9urLNWTIFJW9
/+Z8agV+pLlVc4a1uCZCXf0OM1VknItBmJvAmRbyzJ4zShS1l0z/ckp38QVMt9KL
xrdb0fEjyy7YBlnNqBGkBkS5NoPxN5VAokB3udmU91JwJ9qpVHGpemqBEFTNVmUh
dS6CMfRvZTPsYxqXl0YJvoN37gJUvAtof23UIO8r0j8KrCcUhahs6v9Y9aEgcPVK
kuDFHeVuPe7Ld8rKKwKR3qiyEkKLe81gIG2izf3ZRQVMUa/JgpOK1kIxUcmWZNjy
77/IrvW7lXwvZmzfg8rfaAo/GfkpcW8rxF12j4vaudX/WNEijAFbY99rMbNqYY25
yP87Vae8ESYl6oxWIZL4JSzErVLRyACBoyXjB9lRB3tpYN97F5jIuA3ev+xCO/BC
JhSxP0AFK/iqlvohZ1okoL87SLYR5M/k2F21zSRj9czmiORTu4PuSKY23uAVJftR
MTX4SMJJW1yFdrLkGvan8tD+aldl+vM2tXmjwmpX1iXqQu3jAJ0YbwRX6KoGEvDf
vTDEBNVD/jsX17W15Wo9ekJJQcTZy7HAf1wjebcZ6WZ0d1Blx5K6JoG/PwoqgTiF
ev0N1DoD+Ea/IHYkNctcvVhU3MB+zKHegghe0fIW3bPf9/RoUqklMNM+NfiwG7h2
Ip6ISXIjTY4EBeU5NVx0Wya5BORCfsMj6kKDVGgcX0utf5+r6Si4jXmXK8JwicB1
07O0rkQtuvO0B5xMNPUDTlKYEabjkycLkgwHUp+WkI6fL4w8Wel+EQDnZExy5UdU
QJIDFIMSlDkWVvxp6SYJD4JA0vHB0dG6vSfuXjLGVGG6R2nSzbR54mbtWEq9HC7k
68rJSTIZKPX5O/qCDNqOt7eVFSCx8o6w9NaTgPhPLdOB1DF6P0h+nDeuH0k206Zt
koXOrTaJcSd6a7yodVT9NsLKHXeYiUHIh7kDhJrQcYYenC3Cmm1sIdXwZwQvyv9u
2iwMvUKWs63UrgeYejWg9+CjqSG2CVdFzXSlLwPbMqLfCaDTck13fpE5rUJVRpQc
EBwIvdiEOQxDkkHZtqDf0YH7qN5SIawma4XPXT23sL6jkV/QiEyWMtzoNMvRFj1R
7QieW++B2tXWR0V18EuuCVLnbgFLhXB/PxXleUkQas1y6+KyioZmhQkZr1Rg4CAg
kfDHFs39vIodmJolQcp0mKJmNdx69bxS3iNaZgVNliZyQ8JM3d+4qN7SCC+MTT40
fRsJ0YQwFgidMjnTqJAmqcPoX72S/KW2ux2zcaqydJOGdISlVrVF64GywFov+pOp
kaYmZ2p0+y9PrQkiLaw604eIYdKjG0+oSpVjqrVIRZnK7A7nWFKMUzdT10v6hZ/1
3/OMGfJNw6r1yQWny2FfmOw+wO538cx6FL+2ZMIZ/IEvORP8LTPdKzT2HqeOdvYu
kqMg9vFvG1du/d4/yZ7NniTDf/9JYF/QAc8t3bKUMqi45ciyuioO1dfK/R2L87UL
MLt5jz+kpAtmiVVTg9kvq9voOwCCImau6TLAGZMv0uALtOJV08Oq5Ac7Sz7v8oGm
yYaPX68L3KJI01uY0NUxoSdoCwR2q4cZPKR+zpR4/VlyVOGXHJnjzldMo/kEe/ll
YAIxZ11SLg2Jvl5J35TACSwKJ5tUpTun02il9MH5EME4lIouzlD3b0HrZbwVbE0g
SikF+XtOhTWAqtmTOMSQ3ttv6A5GKCLKIghMi0WjRSUs+742g07/VRkG/8KfkfSQ
hwhF+6v5vWrSJetj5owQlFn4iG7eGLxsf67OqrCHK1WgC211WKc1xW0zcJcylLxb
mHED8IbDPGVYS9+2O3WA/X5popk99vG1XXdXkq8/zD5YoQURutlZZfDx0FuIrGn5
2wT+LFbPIk8L8ODtZAwMixE2fHJD6r0kxH5cT50cFaJzK+ZcKH8Nl71NXUTkOLAe
cylH4JwOosoTadE+FsKixIcOoarUfHpZQEyoinM4s8zVuLzaKAYAZBl1b1vnsS9y
igEBxJL4T8jMEwrU5gXxd0cJJDUJ3obGdpehVvv4o7fsVjjnzTRP1K7BpfMWzkV8
f7kLOqamrh5u+LqfAnBrO2XOIyCZR7wBL5U45KunuwxqGh8JPmGwFKzaTUcluxyO
pNd3XZOYNULyR1iUntMr9VLYQbhfIBS6lcpWdzIK36styD93YXCSonpCuIdw2Qrw
96rLFWDfW8OlO9/dyrRElYSzRnpx2SnOWJ8I9kVZFCxi2bHOBVBoIu+1mb8CNOtG
5UjZbW99YwhQ40QL/zZW6DsZQtUYNbmvQ9DRIftQP6JeHl2ekmFYvvUpTtGhZIJc
YC1cdp0tTV8M97yT0OaM2ElEbLJuxMlC2LInyxpUcHOpkAdfY8HmRM/A7nS68kdU
Tlbczo3p1yMnMTHtUpJ0w4MiT3w9xDfZeX3bw0dWrlTyFqIB+jY1R5kZPKF0W4Pu
QH1+m+Q+yQuirycY5QOsHFy2h8CpO9kTY/h52IDhU4KwwebLLDcZwLF3A23dke8B
yd1b0KP/s+r2ERhsmWEkbcsP4wbsWMJRaXT++FZ00GPc2k+P+aS7jZPFHH1DsDdy
5fr2y6yLdKhuO7Dcojgnk2PES3wcAB939WsGq93AB8lfJN4unX/G2q5rQD//6ah7
FymPqYWHcFyQYLBcBTw/FKwdsLmWVPmjsZGb6SzlqZoHUQ7ohA8OxbFVnopZdGFE
bc1DcxgxXspYM2qt125Uuk9dpQlCJHMVuimT+riVFWmG9ztIQRdLSi3c9Now9uHO
bkY/DfQRAYZPdzGNGa1JuFYicu6MuMAH09RRmq3iHRt+ppnQqXqu7QMkDL6hZ2Ii
C5Qvsd7YQRAEWwoqj3T1KhhD4oNNEeFzeSmyJuSSsNKaUwRgwoyJQMMZ2yk7DB+i
Uii6k4OvqCjFEethBduZ80IH1sZ4GvtQwU0dkz2/5ZDC7ppAV4huoawsq77Kvonw
Tb0iwRp+57/nzeCtn72YQlz1WG652vpG1620kAmBGE3ux2B8oP9qhte+O6MXqhG1
p3Z9iBcY7iBobMHbXmaj12FjPsC+MSvJ7hPH4pcxCIfjA7q0HTEuOi3mNJBiF7yV
yPGTGjpc/xS1SeSv/ybm7iItSiraYM9FTgvGu020dsx0SaRdlkc5hSoM9oyoQ+EG
ZkoV2DnjPzNSSlb8oUVIH3SAaxCIDP3mD+xsB3oviZqZp615XY9BfAEFlRLP8Zn7
uEp9Pz7FlXd2TFeu4fJkk0ntqtd8tQUNfJkP5wEDCV1Qm425wZe2zg7Cgsiw4ATf
hNkfguQTj/O5B3xAyxtZ/vT61R72eeSrvNbXs9XQNCIdUrf0vK9mjiTh2V4hn0fa
6vWsQAmDphTrlexDRull7+wAfxthCPeNlvieDIhRZMZ4hG9yDadhzfbr8u9ArmEM
PsMqlOFjKU3yXdufYstWgRYoRn9L8sgVDu4Tm8wzKg3AfWrJ93Vjn7ppUJwUYnjR
T7CtJi1P8M/qqorftBfx/LCml2o/KyJQWn8p4q009DyHjx2fC14uMfcLxTAcg3QF
OOJh2sTRCtDaB8857RhH35iG0ruDp0qm7/8bIyzG3OCVfw9roNFhnSm+1AHTjztt
79Lkw8qUFp3rb5VyN10AMEXDbGARYQCqVWetOheeEuwVp68bCan4P03V0aJNiKJj
H/lnIxm1KXu4Vk8r6MMiYkL7sB0aUmNvpM/iDgAFLV+Qqw/sNApT4rt24DjSEb2F
9y2O4/Ux5A0UoEpe0L8nq8VJ5MjQOenhqs3nTdY6ISp7WQsmcdIoaGbKPMKs1IZ9
5g8au/i/r/ZKLYrNpsVDJ3k452C9FTzV6uVhuPo/tarrYkJvBA2PlmOXttrWhp3g
52qiNlq22C6I6ssK5nsLrmPlt5OqLXL4ATiAwHih26WJYzTnmNoWssLRgJjc7nW0
XJml1vqW748h+ONd9XU5wN6GRYg4WM8wHkfdaXJ5TRMCTRyhq3/Vxv6RK+seJ65z
rBLQI3mlfK7xQwMFAo0fj+SX6od4UZQvOJG90YR0S3NcrROMzx5f7apfn2Z3Q/Jt
tYNBBn25Q89p/qj26g95wfWd3GyAQx7iThKeIDpz8m29rxzcV4wERPGNOl8gZN+F
O6i/y8qwavfq3qquK9CqHN3RSYJnwCriEtf7m8bsc8iKIHOxxRP7pLhNkl0l9xdN
6wra0tj2IoP1WFbiC21/RWGOScaZoRaCguXtT/VNEpBscAL68/IWep8AyHVw64uU
JpjgYNk2QYJFH0uFCKalk3pkoSVcyfSxwNfYsux+b95ro1hMM+twpAxoDoMzufsX
DMO0BgzAe4WKbxoA2OvSyJHvYoIndbX6H6XFloDzzs7E+337qFMHaQy2JLtsn+N7
+5lROD9jln0Qq/sNSEKGDEvxylcqc1eNySuqezxrlvqH3u2HIZ0pO5NUauC2ls3Q
Xn74hCrnpna30+ZAZ9G7bQXq3xohaK/dmppXkhk+5uqbPA27eLx8Kl5A9ydA6SiK
755QYMUtTe+dIEeQFu/aHwr+/ttlhOKkQ8x5I8eUKAPpWIpD1fLwnZwctR6FwAgM
f/4IBhbE9NS+ywErLBlKs9R737+pE/RC7ROb8LbVugZzz+IzSlLbK0Jn8YBGsCWc
DsNI/eYvGqEBNhLVcBS0hFF9NL7rrvlGjxUKnm1MoF/NUu1zFROaiR37mw5/+GFN
GsaCQMZqcabZgW/4RoajHGyK0nW/1GbHCAzG4Ka+4uOmo2m86RDPC8/ctGV4zpgz
ZAyyVZ9JXc+vUedVjPYUvk2NRjhv5DrrlwoWQwlYhPRF+CHmxsvVRAmwjpM3vJpx
YW8elcgX6LailZnloPpB7mXk+eHC8PyNegjiic44P6Vaud6btZt9SQT0wMh0i7iV
JcIVbz/ML9Cdk4ntjo8EMaGTodM0HxgE4mFfONHJtm0f+Z+7Lc2E2iAvG11QOFkP
OEV5b0eQ8DiT7lwoXadMrd4Fm4Jhl5sxE+Z/h9/uMdlp8OGgzwoc6DvtoC1KJqh2
3tm1SDId7pEFHlhMjI/Ojc3AmR5wfljL3JbzxThkcjD+ubFAGfCTzD81aumYSIM6
Dj/jFbWXzTViayB79beOAN1bgljZNgEK8NWnXC/o2SKWIsGoLtF9SViUU786kApQ
5SkhWN4UIw0/VoDkEguacfCK3CnD/fupE1owDvIngYciBKWoe/L67PkPyxmllyd6
j9yPVBzKn3FHdOPdcFjsL9DK7MIRiYL8o//eB7oUucG+xmbU1lkdQGvZV5ommw8C
cJmMN5naWeSVTyKSVTFQLk3CeCiK/w+wkMkSWdyXBtoD5rQf1VV9vvpfSmDWYCPf
Tnz1l9JUtOfLDKFVO2eanFdKalWEYRTA3o7W+obs6xw8cZoWOGjIJMSJKf/2eeX0
qptlb/DFN9AvzsThWK8YhZ6IyYra/QSfuihTjQHM8B4hodw+/KZbtgE8kIvfAGhx
itNG+Jkng6MvvXys1oHsKU1UBO1s+SHzO01kyljVGw+H9RctoIkZPYy81LBN9yRT
XV50oX27q97HVm7Rwtu6k7Pz3RmuNr+Mdk1H6Sw4SvsKoBWEqW5GCu52zQqcTXTS
2CrKBx+Ok+kL1xHUN7r/ApyifhEVUydMKI6dTgYzSDcHOghStTOCUL2TVxvOBTFm
fZH2njx6l8qDVykt78CVPSTlzZg+ZX3d7uZYqFwQ84K06YooSbPq0dhOMCxa6z2P
WZpzFaM9LS8gDQp3n3P1mtJTde7CfRg5GigyKE4jHPMJOEqSnXURVbBbwMksjxaR
Mpl7HNDMMJ/eAjD72g/xNUjmyH9Cs/4kwax1m7f9r7DojBhSa1Vs2mplcmTz8UhG
vwmwGT08R76kAiF2Oy/kuS39xgFmcZFKSl9bEZSjL6Su2mQbcgIh2AYN8rFpn5Sb
xTAVgvrRrECTT9aOvO+iFfmDuo6kIptjKVYHerhmcVN2rZvTRmG6Ttq4fmqlJ9j9
qmsHTfz7lLL8zBwhOphIz4FGxrC5zobaZ1/XM7cI3g7cmfhoPQCy1nwrKboF3ESE
RcD6L68lmIbMofR3gUwi1KtD2jWS1Mgk6PJSsnFK8U4MOWWr7TZBFSDP0QacIDzG
breiZS2PuUdf0kg1xdCRf8REJg1kVpmgu2RJEA/IqQzov8KfQAYvBW0pzvjdudPh
WmhvO5IQw36JwjeQDTTVbu/x3fZT9kx9CNsK7xjY+f3zCDkCFbcsbOJ6jBKTkkdV
4rrxamlnZLlc/9lrxMiLJzkQd5Ghn91qYvaVA+qhJY+rXsIpA7edXHLGmgdCzy7y
nMzAsX+q7GwzvcqJvvzLqeJ9jNm9GcYdxlFeLPI3P8zwoUcECTHVqy6KuCxejrTw
JWxDYi7/lWIEo8jGMI+jifHAjFbeyiIB2AktVzEmA8sk43uzf5KADV5MMMpw9UL5
kycq2sBc46vzk775eFRiMxFBCYpG+S7GqJf499EaiScT75bmLsQ/hb2rKV5QUhW0
oBKLCfqcX8UE02EFMtMm1zy7ZoxqE4PemQOa4QSfjS/QjmH+SXL6I+PlzT1Mt1uZ
DXqw9jHKd/409WxU2nR7jzdQadcL9M/mzzVTcUSqlPjoYs8VrjjxcUk7RkAvotq5
eIeBpCtpwQzEMDnwMpcuwr0v9+xJ5V8K22j4SxCDiXV91JJxNC69kZvxY3fAR0Bq
w9y0or15jD6jDv3k2GcrDFIBRv8TonN7d5RtFlkOEPwKYF7Kk7bUUOGC0zJqeter
B1n66Ik0TJi7nlt1CEI43m666JZrplcv/ZNMU7SmpCRGy26ROm6g+twFqBz3dJkm
pqhirY7DMQraAmMgSBf6pjNO/47rJw2jk2qbo/rZo6vMekCtisY6O4nk7Iv3XMrW
RMZMVfKpV7GPhDWHVlBJUvXAs0jCx8iAcdTP9WqgqiskNM1T686MyWp69U+7CdAk
mrRDoNCUys8cTb9MSgRdr+WsiEzZVjg6XtH7q4pEpPW66Gg0i3UV3vfNGi6CFLwd
mEM77LjsrNyjkMOsROB6JisvHUbp872jqdVE378uo7ZGZyTtfsSDt1V/pRlNL3XA
Vu2mOgPlZWs/UBzME2WdZB+6u0C/ebhXiUKPR+1LcU7YTWPDSZ5hTCzJQbi7oDA4
6lDb5PrqYqR1PaEMuC/ug1KZgCh5YG+yPKyj8qn9/PDNO9CrqNx+Eisd+aBbQ3dG
Y9Jf2RQactsaNqQjPd9LdM6dj7nhH4JJp3vHDIoV1HjYUYUs7eunjpw8QwAFZzYk
n6kIR3WB8d0jjHDAaWD0RIt7LgPt8dJFbwrR9aH/ge/XjxgAN/DsFiTzJgVwtMsx
do0bL5CHBeFAOmAY9Hf44EEF9uk+bWDbjdzmSN1fUc6G4BfDjdoKChi5jZpYwLVT
yILy4oN9nVV/xJnTgxqpDEl+m2t7r1oR4FxZ7tiJR+Gk9gTTZncieGi8+NpAy5BC
G5YAV2Dn/FvY5+e5xJboWSHCncZm0eE6MZFSCOz9XheCADTs7U0oRlzpZ4LE1jLN
eiBuUQWGxvh81dwQhCJPHZxjWJIiECQ0lAjXOz81yI1A/9HaMqE9jshCyekgQiV0
/bQHTitd1QSdqQeATpQefUBSZ4KNbI4LLJSR37K7W0WtQhkAgv/y7SIOZ1+Cx1vc
cD7hndXgbwuZgmI5Dxcjxxa/es/LvvX7CXOq1kcGDmCNOMD8VqleaflVzz80hWhX
XYPKtFsLJgsHd5bswaCqq0TrU+zYr+Lk5SsS2oNl1MZidP9VFHo/gobc9erlEgyP
zFdDJrrnxabmO9lGJLBrhxxvdVYCgLkOhtjNqyg9m2TUajJ9B3ucns6sL0ixCtfD
YYxMiY4NA9bMZTKVMvMOKzCv59F//TqCe1R8vm2a6kJV33FpbHP0gtUcnxPQ84Of
zqXmOLy7EbDKMaRybc+GtHHDeeVPuTAdGWNGpRK2lU7QOM84jPRWnuTTQqqbAfE+
qV+3dd+H7QyYzsnZrYso1FYLerI5wSKgSVUgc2DpD/RARAvS2wzlrxLYde/x6Z3j
J/YKUlSrUoxnSUAm94tdDfywB0MEMV2NaAPu4ElgB0KxWuH9jrB9AIJ3pUcAoCLw
bEq8H5B5UIaHkW2xVzFbG0BekFIMZNGX9cKKO/ISEEKPvuw6t9jnehubpDBu9qkH
QNytQPOgViL+19hAAh3ss1wPgKwwzIwTKq8Q+lvBOoQzExO8bW1FyTG6DngBfZCS
cX5fzwyLj1zkoRoiRu374R1FatHCkkpZvz89lB+HA9ZCrlxXeTFlCuQMgXRx/o4a
zs72/Vq8g9aBN1w93W2Pno0xN29Z4DGSPm7jlAA6xTLPV1RHWnxRAkr18vjpDYGA
Nbt+rUIBJ3NcxOqJEFRfyIXzwRUGY8sYC7zB4G4aS4nmkgCCIFvY7wUee1qFcNKa
Skf2WIyX1h6NMY9y1UlFMHIciKcy/sF2LhFWo/qlUxz6Byp/whCPxfpPCvfo2WMZ
Xkm2EggY3rlnF21984lJEnvS2mcamPnOQcq7q4cU46FcK4eqO79RBtRmBk6GA3lT
d+ZdlQWfBnYjxAHZ9u36JBDCuDaQpvglT2FYUtLWF8rRbqjiMiv2xroBrSLYZDJP
NOi5Y9J5RhEJ/K24tTNXhPjp1n+XDdyVu/gPqzX4TsXsMu6mmJ61V9HmKkn+rZTr
45ph2wEcn7HYmW/5VN/ZfDr2fR/Bp0pLRAM3y1095+Ci3sFsX94k7IUJDUfiI2fY
qmT8fIhW7bAiB75ruoG5ip/UUDoJZWOqIEmz+FlyZiQ8tjq9vNmnUU+bS85oEwjZ
kNJ9cZYgeI7QETdn4P9bQ167H1H2+txc0MFHfcFPlvvpVl4Y6rlxvKyUnhPbr+FV
u5SI/xXBTKtZROefg4MTfqZlUybV9k+ZidBDunOcCGd7AMW4/SEYqrS251F81Ekz
wsxn7byTdRprpoeAHYd3zoP+L0KCjINROfHWaDUhZYPUqSs2PoPQxCjUJeQR1wUo
SL34Fm2U5uAru+8ce9t6pWO6f7w12pli9nDxI2YKYTsQY/YYo+FltgSXrVM2G+w8
ToaxqzmGnLqJRaet3rsnFblUijQUmhHFKGsuRMzJbKOmdamTS1pGo62nwqo+0DVy
0P2L8BNBtHs5kq9437v//QZpb5VY4Q8FIr+S1Oe55fFhv9kf6kUrkAjqG81ZaCyc
0DHfpjWWF3tg1R5kFQeymM1UAc2Y9kSXZNZ5Zn4/kMzqrerQXu06C+8ZHMIWK/7m
fElbRhg/feQCI27C6F3Pk7ll5miL7ldW9Pkm13uFjrQ1CLvZIEW/ylmZM3ubAw4v
ad5HTbacmXyrzpiLh/vqgU/vS48hzjBc8m64pJgIq9vrtul0QUsblFQAquTahEtl
EhtmrMuNx+NjzdW82YFdhj8qzUXEuRtd4kPcimrhlXG6yFsz8HPuBH2MtRTEQkEO
acIj2DYF63k6r7c5AUfqGSrpVne9S0DPvwY6iuJgtnj5hsIsqglZItYmjaPqCNrE
YzMGA+RzcN7WOi8/lWcnlAgINQgIyc8Bd1qaAD1TZU1FxFRREaldNVGNUOiiKVQm
9dKGfvhRvrZulqTX97XVn7oBFS2iOeWeRDUQqqCHkHH4Tp0YkATU6POBcuSV4S8V
fg/T2zac5PAHBIH4O6RSYABqcyyCNPyC2IqB3I4i60mqp9Rb5xlN0KCvasY/tmx+
oVp9kcEmzqXDw4muM35xpbPvJ+l+8vUdbX+OtFu975HHeV86JU3jcz9ELKSnPG58
nf74qW+kpj81EPMqIrG12CIL7VwcqEOsKisXWoAahPguikzZ2+IILrVqqWEQFuCl
B7zxCgTfucfZmn4dN8egVKl0MD1ekOBFdLs0GvEi5pVbbFCrocJkfFMW74KBgb2Y
0xrbG7Nd8mEzNrOrh/ci1wiH/LhXSHbP4r0JcNPB6mEHlviaknEDW6PnQgkw/2Ft
Ph/DIl0qcIn2BFry720xFQ50B8vgUfm5KNq9JYlSBu9a7zXjeJmaSTs4r1nC/0v4
nmAWA14nNpCIFjKFZxLpn3VEOP230cjy5b2LM7PMYXFrl4NzB2U0G5YAHgHHU1ld
sLdtPT6xeiGuye8z1x2GwlQmNCLszvB/odeaf8bEFfIoAv6AgAbtxEOeyupoQNxv
hEvbqWZFa67jrDEBL+wdxbtWIjf6uXcOfCvX2tnw56N46kuU0NzW7CVFB8VZwntL
c1lG8VSy39Q5ZEwcokhGHe6BUkWCi6vt5q3ZITiAwUOtUPxA5x0pkzLqWviZqCmd
mJzdTk/Tj6kW5hQFb57NR0OLgJBTpuOcyTUgniLMYjaolN/HDdpjrRXQBYE8a6gn
ktvSqvmXydNUWsMcRkX7/9lR0U6et5DZEzgx2q07g1Uj2ZhJ+emfT+SNnafN+tSX
Rn4pd+Q3/IasZrSRd0kVmPshGc9zc444Rozun90472yTn27BV+uhT+a+qfzVxJUE
1RMvtC+ZO9n5gaxO4TKAuTodrURNqUU7ssoPFqb8qDkKKiIjJwab26ZDNOMlemYC
sO3g3O4ZpCjVPNQMWEM/x9GRy2bXw/1CGY5PxmZVcfO61ACzGgRW/ZmuGrr8QPvM
EH4+hPZJoPmSDZJd7ZeGgI44T3NJt6tG5PTuAG9BIRuiCqluzikuRAOqCatm/cEA
uoaYdjC+pNVWVnRGJEEXfi5zkLl/OjszOlXLicaaTImHkw4uKQ4vL9wzeXgCAbLJ
AfhhB5urL74eukPvBmfygdsvamdvS42lKXWth2SmWt0oQEvYYF40myEkQkxM9DVU
VjK1ZqBRgNBvvQv/uSUDa2WYWyxPctSZ7uwXfD1gjsdFD/UlfxJH698D2ExQ5Fsl
GFl5zlQfQXXIgKf90YUJJRYQwXHpUJOawUIK70z+Ne0ecUhbI8YKozKF7+64fPF8
9ZqR0bCmsbeuWZDM4cAGTb7uwaVjKYQZk9nBKQLBVG1R/ew2f3Oqdf/In6ocPI0a
R/Kg/EpAY1rRglIRXHTQ6uyIjMzXKfo8nG6V+YAtabwTq4t7yNYABN6OCQF0h4Av
w/GPOn4hc4fCzUXBX8JTQrQXcF+UMyo6+h0XAWQjHVNfdL3gneMImWlu1KkMuJQX
kHeX23250ngotVoe1Pli0/78seB+uOUF1iO7VrgLSLRojBrGsVn5ORIIUIgwe4IL
M8Enr+e7C0mRg6Nx5qcttNSEl9BUQmozixm8rX05VAe4NL9EbIHkbesAZewmw1B6
iotvk36yNlrtC7MQ6QXq8EpKzUI57oA1J4UmPW1XBmkEad/F9pgrXOQM5WY6qxTo
Vv+2TtBXr+hWfEOOZYnw6UyBv45GlGvruORqGytHM8TnM4EdntkkBBjCdip1+dav
MHohJYBqavB9S36m3oxhDeSL6vyjhtiZ6FyJC+kfK3EmK0yI6ftrdmIAtcMkli5x
p0rVu75f37hQZK5B59jLknubsNAGBR5Mj729ff2d/dPLrYUZeCCJwE+RMR1d43pD
AWSQJDbESmSjOpqomBwQoDZQcvwpnSB0wvU5vYgmESTk4VCrbkrVyMbq1pHEGgnk
/xqFV65wrDaE8uQu8XbGclv2Drdxo7vmGaqBIQIgWscLbVKYCqMKdPmeVvUeTc3P
cn/Q65Gf1d2ArUG/uNHmLxV4gfv4qyl51wGMyHhegBM6iuipkx9KghlN2dcGxJlE
brSsN6xwBAreikvgmtQ7TkALvmoJlVMWnXEBwF01TvbqIzTJ3y4CxqIvLjjR+15r
yyQmRFMN2WKTI9pfLxetqSrEeuLmTPHJ5tANofoOwT6bPdKTvTrTjZmiwVIVHvMc
avx5rTkBnNMgtkV3sizlUqZjy0gJeZ9dVu17CdrgRyiyqGaMlC4vPuM4QCvydYTx
FeBFd6bTb84m9zT3mE4QtRJpkEl5k3InyOozFXTytU/mhDpeeeOjhEWDwLDHB+t1
wPAnpNDpGsqfAYgzyKUn6p4EIAMXHYI4Yh7ac9yUAJ7wskTUO/EC2nMWBUeFc70y
NRzkzqFgkheqsyIQL0ImvH7qswuzdst/JKKoxtelUrROJBQF6dyWyESEaXYVF4HJ
CnjMpVGD+z8NlknAJJLX1JTTxfT0hGt08djo1aXAwRgJ5YOqmHdQBY7i1nRyvjrt
VwjHP9v3oVgfXcEG5wUgM9BDyMJxPp009oHTn1AhCBtfhHiFTLLESm1kd0zFP54G
PuuzAaaUL3AYLAHz3PUtMPMq2wjQOW1sEf7eOPmeZEdMRxauewglcUYVJsSqkCm5
rLFtYDsU5gAZzQNheZ8rdgb5hfY5YPkSlnG2RJL9jGKCyml7CDX6icZR3nvhxWMq
yJdaisMOPM0T5Xi3WwEVMIoWRCTV3lZTjWeclAoTMsVOgLq9DSClcMepXFxuBpXL
+wgMByJw76aXTG0gN+wKFzModEXBYBBNlfJ4Mk5SEDzsuhGVaEwYZRrY/J4yb63g
p/e6lFmlOAtYEkwS4kf4A07jmN2izQhqqfhHSbZsv3H+qNb2fC8aCdyYaxqK2Q8y
1ESaJGw7Izl056aUNRtuJByN8hgEl4Sh0b6KJ/6XNUeT2Kg5nS226mZ2TpYDC77f
GAezdfMLwO21XYC06wGKNOShT/7K2n//e3eFrpVet50q97R9qvPA2bPvVuNsg38e
Px7fb98adrpUEsmBeWA+jCWmFALNRRpoeEQogBK0oxn2GTcwlUDFC5TIwrQnFvkZ
Her9SiGSNCYBr5NuAgVfqOZQxjQ+bSta+EcDr5Mj5MOyvNplaH68wZr+3OTQDN/N
IHbMqj2leAuIm/6Vi5Bs+Gw6mlm+J3DcwyIk/jvOoiURNtFaOzHmWmGMBh05Obgb
17a1bdE+7hnOpoDv8N/r9RNlpeRokOFeYL7uwGJHg6wGibzGm6lud5q+9oDzmadg
UF+Jpk5QWyfe46qiQ012ogsBs7hU2iMjaYB0KLdl4FzzGZ6v8CKeFmFR60zg4WfO
HS7jp9u7oWS5hI3DnI1m2Dh9lVZZZvXyUkBPfPrK6/BjCoQbh9vtOrPvA4wrhckv
+9MT2z2PWfYR6V4iLTpeA8dEfpDdR5DFM+z8ZJMDmMnoqaKk/cnmk3MYqonCDInv
zR/T0Ki85oe942Km+lFzjOCny2HZkLp8pxOJMZncMQsjYJBy+EgV3Elq+izc5NkY
sChf5W/yRctP5tBuujWqU6nVIZ+WLjDPdBLTf5iY+VbdeMUYHQv8JuDoQTHc6DEk
RzBIMLou0JKPpwkqUkkYrvHuqHtcHX3lQw44gCc9lDrKl6RjUSkgLsXcBEyEzzg/
C9bcnBCOEq6fM02Js4NfG26AJHWe9R8YV4s4LSTndsFDwksEnm/yXopDxW4icsEH
2wsL71w7eZaTTswZvzPGNQPsaKw8qxkEbCjfKCoNr1IRud1x+w0jN+dgtPwFMehk
1KbetqKFypbfROcdQnHUiA84ANm5GiMLeef+IWeifWYafI/JAlXPnztR302vOQoL
zNM8/43mLbE5zD6Ya9jpJUA9hnLJPWeCEjAJ4XHWEbdtxVp7MbUisd21YfjvJGgO
VaUcnVdxoyzkQvx8DnZIZsk0bENd3CbOm4w/9Avx5pHnkjZWudA9XXN1zCZsjegx
32MCwOQhtT7fOxo09+auVL6I4a3b72Jp2CINZI4TiJ1qQ0hA0zSOWybLV6qRUHIN
ARIn1FGdqrwmGnFPW2rWc3NOov1BIRjLqdlKB7zEKp9PRZyo7skpBHjND5Mx6n3H
2vLlXDXEADDYaC17tXVhKjJr2EYNO2ejBjL6aoPLNvTYbt4R7UQ0WyZRDfEcrgXD
PF4Y19ADUZ4iT08SirUWrlvHIpeNJfsdeyrDlmvguCvnEcb+vDApCVjj8z1bIUdZ
U7yk8SjSA9ZnNWn+aelQVIfn044j1um5wpFBGrLd0IVx3JwRa4LmI2Am8spSxdj+
3RYBdSxKw5x0txZ46vD738sMxIjbEfZDKctdeEfh+ZQuZQTmIGiwh5oz7If6+tBR
StaG3D4JvJYXjVxJ6lTFLNYEI3/1B7mPz24L2ydvdg5Kxo6PaQt5qRFtLfAYiS/S
/cGTWP3phGvkl8j7PpyhOPDrFRWyw7ogK/bIDU76/x/h7QkwjdBRWUsuanUKr0a/
kfATgO72GRG9LBs3iuprXuUK2WH2xrPLtaolIKqy+VKkiKzQV3ahmxXqLXXuav3J
GsK53amOqtPaYsR+bxMa5ssC8snjwxJ0Q8xXfka+0xj8gaxVXQx3eRIQHZKPzPEu
CXOBAD7e0uFivRCpZk32ycS/bgyn5qLUD4oTwuiyCOe14NTk1mKZGrG85FPvQzoP
/+Vvj/0jFoIf9c28kyroBj2oJrSpKe9UZJwnR/LMls1MRRgA8zhhOMY5mLb6+RhH
TQ8gfT3G+uHraoU8xEfWk7ZVPAC4kJUo9CW1C4qoIYG3beDtpqJFWZQkPlVt6jO8
xM8QNTPf4hAeRAMK802x98WFijhuOlSAfPCKn+l19RKhnPnsFbndElJBAv8tNJKF
T9MK1wWc+CoWVp0C4ezMNiKjjuHaBKw3IFlfJ7Jyd7hfLP/v9BOVKT8Z+zzprN0l
I03VAIfaeHpToNcGBO/99C1dcxPlS7zfZJ9Wx0bn1eb3ge8Hk/MNjh3K6YTsrJb5
xllIADsQq1ACCzZpaewOJ7xWPz5sdiV7OhFiwooAZjlM15GQeI7HCqHq1ZwIVPCk
MPcpHaI+UUyQkRQFtUHqLGawNpaA1Jlw7VW1Nk1trcVGKIAZlcQijTK7XWSUue55
5lu7F5yVh1nnQjY99J+LNaqBG3h3zYiSoKXH/azXxa3KJn+HqBUJh6tszqOI91WX
JOfk4KuefazQ3wP+MyAwa6NL341YzCMLqbYM1vo7q4RzYLC4e4xUtbnJqu7V4Jsy
kfq23cYlVw1hMdY1TLA5tEw29vgHY1S9i+Jtim4kkCNjxEq9gtpNqjXByPSLShjC
0efHcVKPeoewwxla5kq0kemQJpDEUipbtmBQPQqz+LOOVfRukw8wJh3bU6wq8FUy
691qi5blF2rnSehXT/VMLyh65A8+aiVN2dJzTBxaIdGV2Hb62mvEbAUxSvRywnES
CPmH6zCKWcHIDm+T9noYPAK6aFXRUaCn5z/N1sf+U2vXhLIZj3uQa6QpG2lqJ7NR
GcXZs5AJ0NXzOG6oE2vkjLF+D98lLAVHv304v2wwDBv+JfgAFgFnXerJ7JYKSQFk
try2wLfKUxgwzpRRulpT/qX6TVjOJY12TQqYhY19bnmDvuTA5dMs8LfVm/waYG0X
foCTz3k/E8NXhDYlLP+P1DcsApvUdIkbKE70XHMd5cHihUzk5LwwX2Z8TZSYboQu
/mn/5P27l3ZdIMe99c23zMGblflj8olbdLn8Y06rxKUrPwlSUuvz+gfRI24Qn0mY
+pMKihEpsG3t7BLUlhJDUst36aTI5lS8bav0b4wouPrifLQcgU/lodFw5pz8huj3
2DGmYa/nLTjA74dMlr7iuyraj6NWAsnAHzBBgdalHNlLHul3XFAzfFnOyWDPEwbJ
MyaEc0v0fqR6bPUHImL7LrM2rL3v4j00wY6yHWje3eSiMbOtwXFFS/VyJcSoeMg0
vCdGrY4SgHiYiHkzDhpOIOJWi2aRU/PAZagbQL+64fAiY+5hKR8CgfsSzU03T9bY
U1n+gg4aDimsgDsyS/STnIxGMP+VMXQ0zuayZyyk7icEYvl3bO62BnvjJtWuj4dw
dVC5+Wro+DNz/8q1QWVHns7NJBuN3EptJU+ZlngGQqUweSRaxp96jKewyZSnxtBw
ZqO53yWLu38KJeC3S94TdrH21RLST8zuEuxfoyw2gAsOifQX4z/NTvfKdifpsudb
R1gobpIlywA1NgBI6sHfN7W0ZOMN7ely8mRk872c6c3sravp4x4qDwCsgYbDvqbR
yhQaNvEEB4YiYtd6hNgPchRGOez0ADUdVnfMGS2+Lai0YjWAcwTlgRFV/WuOD7bl
JP/oxOGsy4O63jvWQl5C/L9ehuG1nC/2q9mZ9vzza8NiK33VkLdPO+zZp1EU7BpN
iNpQ115wS1c4A3fuTuVOQ3aP4JRfIEWVGdTt3uoecm4WydRebovFJav/qwhaZwFJ
o8HXaVGFXo77aSQ44wjgw3IZ9gg5UC42J2uBgM008GiOgOfNYoQCyGmH/uTWfrYY
TZsNynCaBzEdTwXgEtQujk+Fkw4ITTyXbig9Z5gk+AlhFcgpzD/oz+UdE0vvy/Es
F8Hdcxk/aVfE58eTIXwAxHUX1g6cUbwqvAem7wO+mWmL43Sl5Ef28hUxs1JyIhP3
prZq45T+laC2ZI0UVl6FpeoybGsFLcuUdm3zcruO5La7PMXigk2Mgo87pYwuBM2v
j5gnGsGRkqxJur6isOYN7qqK3Q7ATwUktFlbdwWweF1Y6LjZeIZ77a9Jt+S0FxyU
xiOc2MIeruSXlk/4IPej47sAkh8SrAn6/9wWHjTTT5GIOLTVkuN9ETTowRVV1gSB
cHwRvzvWWnM/uiq4rFMlFW+v+cgR7XRZuq6HjsBN+U0mIIilNDy2O36Ia0srfUG0
7gCdiMJHQsD1OYT+pwNqlYctTD3CfQvIDr5G44Pc++yx9B6FDRG6jJQbMHc11hz5
YGZCsJLFqAMcuIZcvyaRbPnFzRimAUIgHfk/QrQYDkL3EDTCxpysHZnRmAs7CjqN
p8PZ5mGhamhnutQuchO5S26/a2eqpSXQ0XvXwciyUagKo86rjGi09C3dbY7/FE9I
BmLVsL1v9hs+nc3ZZXLd9aTAwzsmyRvSqqpbW/VRuBbQGXkM9OD9GwfiOgSFfoDp
oTf18+MqAg+A7d9QNIAGCLE2FmnuBwDDCzx/ci66/+/tt/e3fMGtxqaPt6EGkw3s
6a1R4yvR1wvITG4LXt4l7OkcuboRf871XFB1eaPGneJBV/AYmTICgweHSxlo1wSX
A6pZkNt6408IKbQAGuYAwig7IUgjreRcytT+0019vrevMwodLsvRkVC/xKobvAj4
DMDziRaTGqIyHkUpE7JSwkTz0CKd4daalYJoYXYQ17BmZqFRTbO3BaLifSBSGrGt
CWBHvGoSsXn8xZM6DBM77hoLWcxA3mmSTtlZDu9ANnX7kBqcIa3NtoPp0cr1F5fd
IPKbi5ebMZQr9OMy3I0KNPHXvINFfOEnbCKFMUpCOoecVM5BkxMc8QFOajFyakBh
EPTQedNy+EwjvmVfqzXayHnrtRLm4CeJ2I0lGWPanLH6fPaivb4l8fmo3yeItDou
Wl5DGG2NgUu6b3z3R99Mo8ax87CxcMtEu6eYElHAPiktvAxODJdqybAS12cIr45/
GgRAGZH7L8QUoCgCApZSrJr4zwLN6c+A0NOPGlfAm/Nc4BBNWLLJYmZKBhH/hZxH
1UUwgTqQHweJpAblk9L0CUR+GWC2IMhUCVOOnVGDm613GqxaPIuc3mSk7phnReLJ
0NbB7673J7BHkkbX+wsqx6m3XWSqhnug7eqeTPB3bH8Br1aiJM3am3GQYsEHEQIM
dEFfYtt2Cpa8HThN1m4jbD5khMtnKxXsDfpCvcxIBvrTh5qjQsIu/QQZ0NNlt3DW
pwRZeGDD1lL1h+Thm4eZHJJE6QyvNkJw0894fLHmUWaoVDllBhZZKhKH2nZsS9n2
58CBBe1Aek6PEe3m1aH6nZWaCnND1apLPWD3Enug3FGMnT//C0q72aLIAu1HO9Fh
nmzXjYjn2ic50ioDiuWd4+ZTRFE0rRHGWY7cCDiEzeE7jsU0aKFf2O+UogwNRRKe
89oviLQngCOk1zSMcNGGYP22E7zxq4ldgCW3ALULtX8dtW0L/ccZS+jgD+2nmK27
z83QdT/eGAzbzqyX/Gx070z27UAOUL1vqvWP6iHjKrreIkCEmz8RKnSBC7bbN/wp
4nzTRK0kMP02sDlxtg/mj2tHlWUpmoP1ngLCWXRCrmwN1YzjyNLok/+P7V1Pryy6
2msqKaE/uMpRVKKdrblPhp3kRKIPBDqszniLf/Zwl9fORW/4WtsUGM178ETvd0JO
Id7ROwNquCP/+qBpdICHFtvbgKaHSyG+VScMhiceWmo4XD5IhTfMyI9xA9j0pnRn
ceftS8vD0nzydh4kOHJO7+JW/nTsfeO7UFnTtiaut+N05pK2iFz1E1hB1kSgAwOm
T6IfkXmO3B7oa+NSc30bvPUmA3REJJT65Anxh4WWPniSBZkohRi85HAG0NQYmk+3
TbiTD9u/vBV2uh3mb/MgcM5s/uf358EIqETN8XJTPaxD9hystlNiXjfRY44l5zlZ
8zkdaur1258oKG1Jw0AshXpN8EjhhzVvOHv+iQZV1MwhytZj9dI+/x2kNnLZe8Sx
FC1hur6hAhJYNMmsahy1Ggp5ca4zuPbzR3AH5urpfv7ggBSO7VsQ8v4S+M0Kf5xS
wzk+mrtoxkle0/kbxpskzjDBZvTfU1xI/MEYyZn3aHby4/oYTFTlxWQ0LcIcgbta
6H7fhESjLqVNZVPns4bSu5q0aRta6EiRndCLOWXigSWhPEelzSnvo4LMS0ELJfdW
7N+rc/fLKvfiq4bua8BH4B1cj5dmCzq//9jmttSBJMka9gFjyUWU56y7u/Igj8IC
5hCH4agsYBt+Lkrobs3G1KJcFl73mlseMCUJ7v2CPtdtG23+Rr34oR6aLbKgq/I7
hyZGoqCOiTUUCHGGWn6/miqJhmjv1DKIqW1nhvOWbHrVW7osDueFZ5lKv1AT8pyP
ATEA1RM8LFuSwzWwSV7d9aGatLtbvP49JJhllZcFwdV2TJLk1cHB/MoWuucTsrkV
YONDK9EtI+4mogaBjkYeUZ5eZi6coZas6fbiwgt7Nee3X42ioTKIHqqXupUXCd7K
BEDAQOHdmxj/87PTXUlVLUjGPWj3tHDD6iS4nABL8kCdrU4wTorODgMVqjoWPucB
D5LJ/4+902K61gXfnd5At2XD/0+1Tg/c2FEpss0zkfGQTWbHlimxvMDLky4jyhmO
AVVQW/06IRGS/h2FbJ3DDZF+JatdfNUpA+1NS0tBU6GSm0bs6U0rFLTi22U0a+xJ
ur26O8k0x8I0Gv7No+JxRP99QugOTyipRwrqPuwEL9WBuNngNBJ14KO8iGZfzYZM
bS1sBT/ZvUoxGGBdFbGDL7s6kfRpi5gymNHgsyjiEfd/Cgn92wJnGeGxq5fY472Q
avscWhVrjT44e+ueQ/FGgGyEJ63G0H3XK4gHlPoHY4tZUuVaIWrqaGTWX49P2aRA
rYy6YtRng/qym4ZdV/uLPwOiuPqvk31A63iD8uotUmRZDweqYxrai+7E8NiKMotl
Afyfc9thoZ8bq/ZdASNJtO+gibWO4EGCerG4AvMlNrOLFpZgLOfhzd8Te4FpREBh
BSf2zjQD+u/bwbu1CnwZVviH66027NxrHyw3ZzoI7ny7xcPVOiylP22IGVnC5Qrc
ijVvWVlL165zU6KLBw9QlaqJ/ENlv8oVkO0lEqXp3d8wiFBTuJmGeV6DD2OjngM9
sVh7rMyfaY08ZQFQrbEaly4L1ScriB6UTdQ9dVOSTmcLC9L9UPlMMpO2bjWQiEvU
uuqZpYdUkl2II+SpwZZvsszcNITBE6lsDu0GeqIBtdvKOf9w4nUaNdMR35dDrWig
/Ok7tF8l58fP1n5LIGHkNhHuZICXKNdhozv3Aj624iZWLBSWKXMUy+bzSjKnQAwJ
9/ofW66lRQkhZdd8ktjGNxt+xioFhJ3oSwc/4HWdoLej023Q8FwASNLgvbMqYzrw
NnMQgSxVnv26YHrXcue43xsvExKFlEOlTC8DIBERi0Y93wRvj3ESMJRThJuG5WMs
zSJEKzpq3VawsVtKLES6Wdu+ePnopsUy4bR9B4qKNkuI39E8w6FMnMDG1M8NRZgf
BZ+C5Nf1Ia7shGBVty7nOwks4Pz2SXUA5jqz3FWMBV07BwFy/ElDydVdksq/zQVg
Kx/lQQmu7RdIrkxmnawiNdWja8sQdj9iGNq2a6CjIH8Os8GhCEyZvzH0NlovRSQG
e8GWqz7aruD0ulioVeeLsF7zdiEqNkD4DFYlZYiqZNmbb3QRuNq2zI7HlWKV8ECJ
VxtgPzANeOKRLVIghdGetGGJ4mwp8blf2hfy7SVvTkxlVBf5P09Gm7lAzjFi8/0h
05FVTCnftFmTNJJyBa2WdalwFvqLMdDEhlVOCwv7Sig5jKOAxnnARqy9JIC0ebc4
vy/Xn3owU+nU8fzre1d+1GcGOcINyU4W6bW2y9XqnhZiPVzl17D7EOQe0tX1rTXI
UiRrUgarLTVmYK3Mxn/6KLzWYldvzdM8FAtzAy1FWuekJ9IkVDVlHanM3YiTbj5s
v5ouWIFV/LRuLgpcHTKmsykl/W6Ws3eqp/VM2cQbapEpJ1riTSbdWYxqqJj6QaZW
2lZOtE/bx51BlEsS8+uPgrsOHHiKsNQPx/1Tz8rIRD6syHJ6gdnIsQrjLEvXFdmp
ymlc1LJ1bTCnGEVzGTBSHPwzg5kqSI6wHKBJJNMMjDOT/UNNRnC4ffTx93afMNv9
wNKaO5vKLgWEX8e+CWNPVuoSgCjk3YHP53b+VIcqi1M+WQrcMd2B0O6mbBU3R7bV
MoX28ScuF5bNmb1jvRbRnHf1cGPkv7WH7NSi10sNtXqD8Fr8ucB75Z5cjyCfOO5v
stTajviTuzQwv1VZY5BoOQQcjHLZzEMIiiOM6y80mE12RtTdfVi2+E+A1qTNDVIU
+0F91ixzQ93dmIddqjNcN5O4PA4x+bdVhbsY5vanhv6GH2zbBcrBMeB/NVG3NFHg
gpT2vQ1NiCvsfqJ8/GxTL1QpVKi8c6krkGJbfHuf7Y3gL3AFidZwSv4k3D2zfALg
ZhhU3g3roV8tRqd3GtB17mvUz5zmO2YDlPNod3Wt7eCyTLRdLAI5x/ARoqSDt4Mz
AAxgouPO1AIFOtfT5Qo83v+BODosfRTZCZ9OyqrUpCSimQg70qqMJHJv0sMElIIS
mJmYYl5YeWX/77RZpiJD2635kw+SAaOYdf/4rXbZNKSIHZP2MX+bSVO0maQarQBH
q9PzV2eddZmQGfzrMmw7C3VZLOKKeZ/wg3s6sVwdfNntrZ8w30C/DnTDFotPlCAM
L1lWjNFa9LizEZdr3diYRrWEUc7oRP3XdJDpptfnMVDe5kVx6JTAENzxYO4pEBzP
XGYiqESYY2GWjVjQOzLmGfVvnGJH0XaisTGbjwcxUHIYMhG+p8I3RJjCgGqrRwAt
QzRInew6UPTE8iGarfD2CyMWTXs3YuTGgv2lh/xzOfMHOEDhTntwZeiab5HqrPSm
kJARx8eUMZjJB7M02GBG7Br5OhYFaFMFj4ruweMEKm6kn82VFjkJ8Z9JYJ+yH+91
4/uZM6B3+WA35gXcJ6YkjNCTbz0Xaap6/bj+WOWgye/NCSns5ylZNGyBkBVRmQLW
8qBYeUHFncpRTK+FU4sZmUkfofB+h1fyw802q/k5tO/SyNvVrE+J8c7lRQsYIuXB
HkkjGENn71gcOZx+7OkHAjNWgXnj6FDQSyDtqOGy+EJ++28sxC5uQ/7CxtXnxQAa
RvBI2CYwg6gyA7pXqp+gTvO6y2s82rEtst9OVlL0ibg+UejmEAsx4NK6sUWVFJic
5gloO/2WldwYIVoWu+iV4H3tRYBxckWaIVVC5lJFCw0cz+i0dpADfsZ0XyWLSkfI
Ah9ieB4Qqq9YXNc0TSwFWKaLtBDB+Nfe4UVapJ80vbk51PXItg/cMB0eopNyGN7r
Qu6dSjkWAvHHhtBXVHkJVeaA4/Sr38b9Z8Tm95w1QsM8tMYL0+giHV1p6YRgxJhl
h027biCsgNjzO5FP42CHCf4LQRarn69wNj1RRvnCow2IX4zNLJ8Eg3Kq9Eyu9QYx
f0RqIK8CvW0W0pZKZBliqO9iepoYk3cdMAnLaQbYS/TLXFaqo/BPcvb2tunBrAQP
JC8BNq8Nh0UoKVDZ42BSobYthSVvpPivpw6z564dQEMhJyMDrTHcpaJEusy3SRRT
IeP+DkzlPdQ2+nn6pvCV1A+Qo8RBnGHCOo6I/4B3eq+fHHl9SzXWnyUng/wkZpqO
8ORi0IooY/TFGbWxmeGTPtq1hgwiyvqFGTX8L3oZUAaxD2gpt+fnQ4Ky5Y8OWcl4
0W2ZzD/xhUqkvePlQK3V6sssj1ekRYNvIMzL7X46T3hc9KWhj5nc49pyHHhTCK9Y
+laPQ2pCyTMU/UdN44QFQnGT9xVNIuseECi59dHyeQKNI6B4u/9eiJG1xZ6L7u0/
HtY2NwzaPrJETD3wi3DDIXdmAbN2CPlJZjbs2T+jE0/FmYM98JQq7GEVKUaORP9j
cA/VOYWcVusVK0nr+61xvA40U+SYpvTi3Q8Vam7jicr+48f57/cGEyfE2wiQCcEm
wa2dvwMvaPuRQLi81Zldr5aU644Ebt8MxjdLYTFguNKzsTZu/3DZIqEnU6vy+EJJ
YSWgI4sTB+msM+XIrGfC6vVsAIlNs0gjanlMcdVAZjUNYlL71rL5aKxsZ4aA0KVd
cfFkyK65ZPx5ry2C54vECcZMYPX8YAH3X1Yb5rWnwiQ+OcI2PqKX1xGu2yq4a+/m
IRyGGi0Ov3DOzXR47uk4ziTihS1mtSb9z1O/0cZhhlwQujsKHLdcqYksaYDnIL4m
39gTVmkt0l0zk7P2kjjKc/utz2pT5F4xeZDrWCs7XZ4OP9ssXzpQsucFVUnRBZuj
4p+5ajXgfCJaUgqPLut3ZTdTJwrwfMQTR/hPODxcKIayqGi6ZetH8Jxta0ZiHd6T
Oc8oHm18lqZvzCkvnDXeulC8o0RY7X1mVUjzxtqM4DcoWnc3kzIfMv0eHxpupp1m
WKitlHm+2ezt+SK+6MpPzncgMstKSXo0iAjPOms4TduBETLq7WivhFbDNzi4keb+
v7y9Xzhyq92luu2LjzhPYaALb3gMd1g00+I2X+NzZiGy1GCvbrT8xmXFOXCm9Wuq
nQN8BpX8Qh4JUiGtR2RfQlbVIaSJNt0JckYTjBI3z2Y3wvtDz4QZTtMPUzPr9qWQ
XsAZAfDmlEm/mD0BuSVlYZXDNkaHfU3O4Ce3XvQpidS4hMsKWWhQ1r0r61E4G8Lr
dg+ZPhJ50ALBGOM3Qv5+iN3CdLd8LMKWq08xjkCtPdP+IfI8/CXQzqfvt/eg4xyJ
i3mLuyM01Z70FEdhxV7E4kqa56YHME4nx2jlKYmMGXzJMZjyXMkueTlErhUQ5Y7j
2QcCZp7K2xBMIBJI8Z6dhnxp2WOby9Ll/AnIw7tx4l74v1bkxirhutvS2pASJa+l
EssSRFOIlGalgwQdldemCRqqmlNVJkXCoCHfrElw1eLq8u3U5kxXBGhNoX9ktssc
nSBE902z5M0rVwxeUqMWHc4aWPyzF6gAQ+3QpIqJ1e7AtbfdX4ZSBK8srMELhcSI
Wiec9ecQQizLlxM0l/3+1tQihWRPU2kxQtFHxS3CoL3UEqfVZkbnx7ci7CqFOFOF
MCLdDD8wz+1myhVGUAM72uQw/+tTJEnvVm5IfcLHAwqbVH3+WFoh+k3ulRrGs7vp
0Jpz59Djs6Y+BRyfAdLrSaBt+l0EAGdr8BG4nhvWit62qmPaAVZ607XuelaNV8Rz
S7A6ov6x/wZg4b6S2b+CIwmAangSSs/nD9y8vRAAy52l+CoIKMdBjds+eXTVVMDA
710SPi3CrVkCSquqHjrTKSo8zFXyASkF33+M2ti1F+vPBNZYf7k8gsPCxjOksy05
Iu4KdXtdXTJ3jKcZ/INhpvs1zkVNKK1WHJl2dhTPzbc7lFy1Yn3Y4kAgwnAOdjQZ
EN5e+mAJdiYWTPAYtBGslrB0IIIAb9ORXOot3QNl9OZXzSxAuLT3jegxOhyp7/29
bcKWmCG2At4Hnr3BSzgsQ61302rYsojpmZtipDq1a2QccemHwnQM3cUzJ73jFW1u
OYIze8JVDMW1NNb2sisBw/BLdIXwYHo8Nk8zZNC2sVmlABmzt02Cg0fhDjL+NhxV
3qCS5csz/wFai0MAptNcLunLcG7LL8EPwIGY6E2Kum1FYKSYweKPzN3uFkNIek4T
7KxaeBRCv8yjLRJtCZeEq9jNdhAzwDlYOnm1lZYHwykG4r6yCnacgeJbANAB/jPf
qOlahsh945WO9aGO4rgbwHCMuOjLYYZj91eJnzv+aNFtKtNQo9zTIl5RFWeZJ2TA
l3hTCfaP6HZPUPdHHhZhOBe/Jj9ukL6bCmAkWpY3GHKKESddsmfch9lnitwwp3D6
cFlDvB6qGx9NEzetrigDg7yBajgGLKDO50TJ1hBWNZZJz17veLtjNrDPR/ona6Li
lrIEXBLhQuK9CM0Z+6yAuCpHyuZR8ZVUJBtR710FUj8+yasw4KuFWs77w18OypBX
SZ1kB/qzQyxO0fkcCICyC2LqQpXY2t4pLQwoQaUOaMe1HP5PMIV99vY3EF6xLll8
mCdMLH1M0B+ZMdXvXyUdbA1T5koWJqroNLmJSTOUEw0LSKcjVUg3teP7GemuLPmC
AxN2RVB4tMms55kD+5YdBrVtb/hDj8WOUB0jBHMMJusIZYlW78NvdiDi5Kf1Dsa3
wVtiePGzOHBvLgFDbsdH8AMb9l8xx1q+pKRRoOa7vcbaeSuC6lSJucmJYG4B9FdY
Lslzyz6057Y6emoQqs6pgdjeCY0lSyagv1E4Net59J1Dj7+W/WcWwBm3iV6xyO7Y
OfmDdG4lnss6BdEe3Td40VMwyiVCrxUvWMlKCMbcKNXbtPhCeklCEfDDdeT4qr6j
phY1RPnrOU2YfVPP4u/IHKGt9a+l9Zs3D2I/lwLXznDgfYOhs97GmltMvxddniwm
utCB8Cy3FR/ssLHcGEjhA5nLN2OLlNVqLVVu/I9+blfoK12upLwsaKGe1ootS3pF
7VMjmZg3MYXc0ARP7CUERSzHwY6EaoA6G1ekq0pKAJvN9B6QHeVj5MMXda7oEv9C
m/eAs7h6QI+oSbsLGcwtAlo4dgBJ0dvBQ+EYQ+v7b/2fe9UNNuCNa9TCKD+NRgfB
/V+FnxT8uJNFS5Y1Rml1KW4ZnpoeSGDjE2aSNW73JyyBxrMuDfw7bZ0sk4eQKCpl
Zjgup864pTY0KTI19WRcsYP6nTPe/eHxpg3I3qkqV7ycBXWH/5HrX4LFozdOLQH0
FUo1i/i/HY7Cih6CTcVIBM5ahzlUZSetVCpgWGxaqBdPxWHjnOlf9FZQxOMqEZc8
GAv8HQDSpmQuzY1QdBkzrtrHxApprl5kveUCo78Df6h+DGJtGfj2AbXcdteH7K5E
tQO2yHIQokv3o9g6/BRLnwDLe4xhEgsTkz+pm9gfQk9LGZYdYuIBVDVe/AKlDQAv
m5wgLYBKJ47YZwPa8faLpzJf5OthCgRegV472yck+p29OjAk4ZizM9tU2XejM5Fv
zeNOd+RWGKt5HDMtpPOFNUOljkVQGh4JukyjjqAXTEbPpg/t0ctnPUw3PmGPtQLd
P6mbFyCjis4tixq35r8ghbTmHTNw1picaXPB8RRncVyK3+ntUYEkuW3znxy55XSG
n7Z7u6cx1fsmpC83zVn36HiuqKGblSmccqBA5xyXyxSWOYHDoBd0zAD1E4kMxJ2B
tgk84CG4VkqIsT4ZpK+WcWuMkcblCNgDx6zdGKDQqDXeUxejPbyUYlVvZMzb7/iG
FcMN6+dqZbl6hXEoi5yXsb7Fpsy4eQWvIODgVI+/UcQKqJsdADwE8nvpCjAGw4+z
TMLuwovg4+jTWjYRsxhYHDxHNxfIy6+Au9koBnT7+wjRaNfB/ZIsUYxF4lR7n8yA
0im6+a4kyM0MEwQnAKBoeCePdeTwVlHUJUjoLHiDABpHM27vxaJpcewJfcQXWH6K
F1W92EJvn8QtXgf5NU5ZUlfBxu8DsBNHi5ogXQ9W4dtRtYgr8WW5qtqg3+JU8/rz
ZtEy8FVYn4rh6oHpwBXY9cZP8HGi7GAzP39jKObe2xe8n+hP8ifh8WMywv+DYmUF
5//n88/z8QG7rrHOKwV7/dYsgUnR1sO3u8XHkAhRvgKrhoZRQ/O0nCnw5b4QWlX/
25IbDpOvVpaFuYrHhM3fpLo6RqDG1q+nwSFSDEaos/WjUPMxVf/2Xz/XcxsLC203
1nLT0ONBrkChCk2bAqZ2wt1TN5NsNHo7OusXtNfEwLuSqt0lulN0dlWk3+WSJwry
nNPQFvFe5eQ4lZiAsi40ppvs/AwnNdoI9C619x6OE/sKhuFvfUHPODr4CPSNJ3px
UPa55lavkK5AUxZ0Uc+lG3BOfbbjg5m4h1I93ERe8Ej0tYuAFVPnTFmgzqyUlCTE
+XoPABYIh/yFAfBYy548VvzKq3roUKKVcZ6YA1IQTES6d2Vzn32sD+PEDiocup3u
TIWbYyCBkYW5sFdUuq4aeWPONZa2FWv+EJby+njLIiQIdRwG/XIpZXP9bPF1SR6R
npISMtMaOL/HZQ1t5vlh6JfyWJ6H3xDNKa2NgwvIolWafIeBHORpM8/ZP0hbVVHt
TScwyK0bsmQLczSjgmwxuXCY+rJR3P4pf4cGY+BdxuWNl+nLX/9Qx5pX7hcwwkF0
Pd9NOdvTqEfPNsmvd38m0rLQPu6kIIfdqK0ykXzeCAdOrMWsW6FtktU4Mr/fXeQ1
mMjIAlcF5tcz4rP65Y4BSTMLH21+AMJZtEEqKITuePOEvFu4eItg3M+hCoGLK+BI
OJwsJVijXTvHlGucaglU3MxTplcaO1y+3I/n7k5cTN1iPiY5tTdeS+nBHBHv0iVg
dh3dfk7NSgNXS+s9fp5D7gcwyDKRTcEULIR+GJcziGN/JcizpCrJqyTV1MgtHsXf
k/DG5qLxRqFCkdCv9hYXqls/YSTfYLOwVW0VpevUo407pTUor7o+rKwiQHBJ4TgK
oIDwWPSDipi36AA+u52sU+SqVapjRps2Ai+KzHM8iFx84SCs2b68s5PHSB1AWdPh
vvYZKlGtE7WMLl5tNt6gvd+alW973g10NCsvw6vShsJRmV17is9PECfSteZQHfuS
hq9PV+iErDl908Ly2kyAKAloGFX1fC/GWLDOlvOTrkxAANGxsTeELFRLAURdftg1
GKvR+LbxPvs9ulYLoC3bRONKZY0ZWH5IWVE6tKzwKhM212zDPabn/l64ye20p3oi
fHGbw9fbDNpyHo8rys1OKHWWPIeB+ko/PB0QjhgLphPWq0K6NiU+cdhiU7dkjHkC
xtzEQEojDSnY91tKSOyYKPNK4G+THGBHkJHPfvhrqoTUV6SUDl7vEFtbf1Lj/QUy
obOHAd7Rif6BWgWgZR+BwgYVF7lqQt8yVqTEHrnyl+R6RiBRzH8K4xiCja3AA2Fu
UoRgEG0hVWgvU5s3xl60YpzOKhP5/3ngwptHOwXik7VCzzhL9eL08EJPJJsx55K5
wuOpkfCe5vh4P9T7sstwm3cAWbCJjgXxkWNlmP/EvQEadBhKfDuWEUVltZk85WbF
68sGt/tglQtRlYE7YZmtbjnPrIszP4X4g9rwetu98dPisBW4/YuxYLK5HZwbiPtp
SqC9Fp7NZpxS5IbazvledfFifC21h5gZIh2xWuiIrFpSUbH0mK3d3PIaxBYzmYms
YgcUaz+D2+Q6T5SEfEwt223A/0c5eyhFZS+57wJnNd3EcTZO0Mb1gLXVfVjbDx/P
vlMyPQBPOmIrOzSQ1EZcbDhM/i/eyiCldQsLgKtfbv/LKuJshL824xZ4TTh6MTs/
8kd/AR1aYzoF3Hc65g8vURu8riHx7+GGynvtA7ssbAht8XceYL1l/GbGmtrT5caa
Bkv/s++wgqP/wXrzwxoRV9qAOCn5XOaL9Gdw1X17Vs6GaMGfQSwfxWX3DwgSSirP
BrtL/6haiIp+pYQH2KgP+i+u+ndNk3ZFq17KJkyin9nkNuXpdUDM+X2gSCDLWKMP
x8S0LFtnfN/wI6t22F1TeOYBQt/UTeRUjLtFYkwz367Xl/dwVrrpGlQc+ySI9QpZ
7vRQS5FHEhLpEBKyPHJIbLCjxOwyuyUvIKY7j0QX+WoB5wi2kyuzgUy/38EHwmt/
FLOuaJ98UiQ5x3N3PY0de8Lg3AR00lh5tyv1PXogKXa8En6QJgqjoJjZH3FsAVdd
pPonw/TVMe3+Huag4/o5nBx7bk4dhBnH6k6tGEWvITZwXZkN1Ckx1rwx6iSIyFRc
BmG4DXhGp+HHgJ/NqH1vK8ckvf3uWgWEM9gzYj2MbOunPzA4FWEvwslPHDVq8q7j
fCyut47vjIWQ+CfHMo1sH2Pu5lD1DF3bbRMysT/WGcZHUgTInPEEvygNrXbm1iSz
neX4dibpfFHNOrGWIyvHIKuOEUwNv45fmuNWDZUPXJpxBxouulA807LxaSpmDAuB
Xwt4WVPrfk3RMFkl8cgKQE79gDw94rvSUOtJl4STpRxXNzOgqbUaWxVOEY6HMsFC
Co+RvHaptZzBK0sKXGEkmW5r4sNMC97exg/GWrOjX8gyXa3XP1/7CzbLopUL3GA3
WnkKHuKA8q67SsxVyjcx4T4C7D6DuTd/m9s+ZUXkxu+55mEtEC1tnHQBtuTF5ufp
Vmgr08sY+EB6NhcCTTSV8YvjqC6wbynbKxAUccrD9U4qHEqLzebdCyN1f1+51gRQ
+VREr7ObmKzOIRG+9ujz4skanZGZyzVXCQgbcZzqefZqvcgK25RVdY1RTsMFR0lr
5sn6IDW2QNtvrP9oWgBwtzwq7txbLpJ3aN/KRxDHIm2nAW4I6t3T4oM+Tjo0wVco
h34+dCZhEy9X0M00dTEQJuoXNsStKcPlkfdNhi0vSgLBMjx6iJTnglF3whc20z3l
6eBAlLXKrzgbXrvI6jY4cXqlk2Ai2rxkKu9NRuco/4cZ0XhP1uVGeUmcqYbn93/l
Aem7HgUUH9WYiQSDdQq1Vqe4517fR3NCixhaJYZa4r6ykWWgNfHhVW9tv9KdPNRq
ijUb6dANL4YbWMBl32IQTuk8nh3UIvFvijLkakXwHhYtdr6InJVP335pOwmhLIbR
V9Bvo/94n/JRrz1JQT6oS/S2j/WZg/mV4aM4NibaodTa9ePM0syWkiWDc2NDNArF
fMIueALyLXYi5QJ7/n7lEH4UJn/r1xFSnQ45Pp/U6cEfhGxSCJvbZ8lPeUZt9tSG
S0xVtSAeSxfS3b75nyuOrWD0p69c83VdzwJaEol3Y73shbjcaq0CreWZxh0GXewL
RnyrmD4t0bK4V0EcHSp/hAoUD7xiOsYUvGXQqrnPmUsUeIctX6TgHlHMPNSc6RTN
xTZXYzfBtlxNE/n3ldW+DZrtgr++gfFYCMSt/+j3Ot2xaRKPUEhHDGkLHxmeT3xB
Ka3L3yPjerd9eG/EKbBFhWlgAyaweDfhEVBYf66AKZj6QEku/jFvJF74BiDP0n7I
Nz279tb4K9Os4nccyl0sJIlJaiCNFLgD04nHlFHwffS/4ALhq4X9aI46LiZNzI2h
ZpzeHw2nHbVFoxrpINokmIueheDDAGP4WXWxItjTNofAvb7/jNSlE1hOTYgBHMuy
L0WqmygkNUL/zshbIg51+kIcTElycryPDBXWipAeAO/Kt0W7TDf+KwB91u/RQw2G
ztmnilEB5MlBr5bEe5qKLwwdc+zGJQOr1PPqUWaK0kqnuSJG2ft9dqeE/XbfBT2v
fIZr8CcL8ZBBw1RmOCpsS1nvJQ30uwHDbOwN5AupdO1wjd/tDNTdnVkJWG7tFd+C
/MZBpdfxu545XwSOLyI52kgvHa1NuvuSWTY6F5mlWXAbZ38WJLm6kWrYV+K12l1r
FsZm5b6/ayDjhd7tNFeJn8wyqcSNvhhJEhp5xoN4KU1aSzbbLCPE1Ko8al4cycG0
Kceo0ebUGw/zi+C06Ea2vkMreEhwIsfAoAeSGLoRY3lB9Q+B7hycNQ3vZcyNql2V
mxwSTLWVV6Upc3sVSHmjq73Cei/Zh0+CLeTuBaY1mJvZG5gOwQl6VwGrVXeBsyuy
sgiqMxMEV1aNxLa4ApwIdTcTxb+8qcdHktrasNhut+3f6YMgtKT6Z87uvPOdr86T
Kx2SGqBfvr0vSwgrBpL8/zvqEZ/okfEADfQifFKaLeS0G8PRGHLFnquPWXAaAnNj
/i3ED69Krw9mKA0GpdAoTAPucxTV5s3k1ziVs4ZYgYfWqF7SHdOIAB25Y+dG4Ygg
8bSsuqnIvvSk90cWT+T7Zbqpeov2K+EJlrUrvBoEWzRm/68wnmuUYeLF+3nggImK
bQ0kiORCUkUR6rJYFK8nZT5Vy1ECOZ9/tgS9+BCt8x79xWxK8H8DVPdwhPdi3N91
eThgOvFyMdsyWWwkymJbxqQbAkgkLgrnUDW5IbE7wwg/sKSq+SlBQpb+VNbiTslT
RW8EGZVeFvOJw7Yw30LDBPg8XKMd5JW/zIWnd6yvCJKbGGXch/7/akRzRVhb4fnA
GgYYIl8NlMQDNJbPD+cR1PlPPBrFI6hmUXpt5DS3k+NQGRM6irLlI4M3G5vol1/J
6j+OHoTo+GAQpUEv/GvqrWwl9+IKVGHmY4APWaZ/jX29YysAF4ygsulARPTtvRqE
IVsyOoC+XI8MUr9NUvpbUCt7UWxHrIKOaJZ/CObozzivFugKyRbsu7X/R01QprXC
RhSXd6h6ZmDNt+2PYaulHUjvZN18Fz5OOFMyTsHuNR0HvLBTb+ka/YuW5gbYNBcC
BuaHmxe/+LzZvL09QNLrtCmu/h4Tcd8031cWbWYp0LM12silPKLlWQe1XCfvnLn2
4vJNIxScOFiP1rxTID6IEEpSGVUd9dra2I6rdqGInq9bZ6hvni2V7wGMEfby9Mzr
DgcxFSWkSdDZaVMOK1svIBY6hvMtVC7yb38jmA+gZwlzd8Rgai81EBuI2QSd8M1p
+J9f3iQ+6BHCIGa5dgw9CTKUQQbETJb0kvN+smDGNKSeswjytjJ60L4bB+6fNVb5
9++VI85NdKn7zcQjf8fBtOsq/tzzwWdFJdmlJYUpEFGxaKvIS7frJxzEtS8KZOPS
RDRRygn6xu1dB5nUnuQmW/YbBq/erqlIyQEQsb1Ak3Qbo1MCfuZd9mCw2AfmXlzR
CZcanFG7fd+WBUO1AI+KnxE0qwgDfJ7zzgSNBZ//a4DzP6rfCjiwz1olEU6Ue3dI
iVbJnzlHXiIdhVmNazzbfEe0ROgxHF1CrES1LLyFB9cSfl7sAaowEdlE9kB6/fxK
JlPIr+qvxqOsAScue3Rl1WCnZ7GTwzs31O/4L9CR9OcmGR0WwccoTBWNnVW8eMkR
X8NqSdZfwBnli8A1IudPCMZMlSELfuw8hxmmfxb8WxCYdh7IDXKW9pSSe4wGRWWe
sXZlphlFIn4pj0OWdqQPgf2pHjLAEezwPvGRDHmIYgi0efQUelZocFKOI8dooE8E
CdshUUK/tzDPIScS6RjDQLIRL0RxrmJ4abz5xQQZCyOSa1Q13xBUksKwi50W8Apu
x35VT81Ey8EOWhpN2I4N0FJXGD1Bc2GCEYcNep/bRuu3W9Y0Ly9Vshdn1UrXkNjp
Bt0IPSrJICstrU4EOnHx1c1yrnNTH7MKvRuVJjQiWv7IPJk9pLblP+LV7cHIq2qf
QddpLaKbK8HJwUeT80IjsItOSDYh1Bx/Em8/DUDwZtoyC84Il6isoW2V2DV6Ot2P
BnzuIVbNGYONk0g3zSR/wE1AR8UQXwdDxeYdHxpn/xnJ4o6aWoO6lnTUD86btUG7
R1e+KpTNjJ98T763a82j4Q5PkmyxcCRR9bW0U+TIoAhdONcPmQjbGWGOY3WII9Ls
v34YG0+dCaa4JB2g7LrjqiVau+sS2PdCfOxYVP3fU92/heC/Md9JMJ5fbxTQxt09
+xVqh9Fe2lY8VYbmlxieZi7e7tJaLfVeFhIkBOy+Zro8kBICUJEXyrPBQ+J5q8R/
JQlm/gmUEhc2+aVa+ZRFb/IJ3pTMgsTSfDsBS1RwGSwf12uzlIPKR+g8BxWGpF1H
7mqIhQJvxBS6NheJsUKdcUsbjRSIFPjcb/euyJkMPB2pzoCS/7pG9PrmuKqKiH9z
pAGH3ime80RqRXwyKI986ShCtPXDp8xDv1XN9az7chxgun0FVOJjqZKXzF03itiv
uw3A4uz+NOxHGU0WBp++R61rQllMRlDoqg1JMfO4Oc1s4jYC4+JrgZ6EinNfdhGc
KZgI9Qoy2Coua+8uKJZ5aO7hnmMUY6Y2ZLlD4Ur7gBN+Het0oHMF28Jeb1gkqUfv
efhJ5WaExcngt1FF+42Ab8/jkXTJYhoS8p4ZFJ4Bz9Azo7dwUEJppu4ugFIdYIUV
3j894tWyCDteU5wFzzIZ8Mj8IZF6d5wBEsgiTNKn9DKjTKlS+f1NcijgcSVqE3xb
5Sa25QVcbd2UgTN6urN1G0RA2zMhNRWPDNg5+1PLKMEsOg+gmQPJscYs8GetAbXB
Na9jHxAAa116uj4O+pFzSy4xbb1u9Klza4oTlOQwC0Blff2et5zqihR7Mpw4JKnc
YEWbcfjCKu2+t97vDUBQlLWW49AAv1l0fRB5nuOm05fDgBvCUmr63YPEj4sSQfRX
uo6trzmXdWaheDzydTHsyz6qlvqXz8LDQBRCV0OzjiZ3r6xGvuDs799bYkaBxmJV
TZOWvzXZVcwrG67HYqlDo8rKPnQ8z9NK+UpQWcH0ncDk/rFv3n2MUdnUAkAAaEmY
T4yftXrTvfNuIT28B/XLCmeN9ROLmJsI5e1iVZOO4FNOyurJPxaT1+2+gErB2KOc
dDFtjSY3+iY3L9ZfIg2CMsX/3EfeX7k6qJlj/NIO7CfqTQ2/SDrB+oK0Y3ENlJk7
znuqfEq83fak62KYkl2oe57H7YryRKdGuAEA5FcwzBTFB2QR8CJso+YC555qYrGq
KmbGbQVeaOKFIz5ckCRyfS/TaeBWkfJRAKX9jCZfV1R9fRRCoaDNdGBbEfmXvZJ+
CMchOUGYu9Iu+8JrlUE5gfXC/355gC7SjHH/kdolkmKWWOamdVSYlBvZHTjY5Rup
UHrE5rgODwgXGBJrKAtaOCQLY0JnvdxDEg27V3b+sIqzGYRAEhwP9kWP3CjN7gB/
t7N9bY5Owx2IyYHuJ3jRAGo6ItZO33pl/fyyrBDhLiAGId8cxlkZpjPfpcR95a1C
v7tbfUb03z8gn58L2etkKTM6YAVfdYohX9rKHvld2N4mw+VzU6Es6diL391GqR18
uydvBVKNkTmisp0v0/OP8k+oLuxGYdCRNuvid3oVQgJXZxs1HA6g+E3vef6m2b4+
Bsbc0XXpR/GiLEdivGNywd/17XQFMWj0OW2YZny1LLL6kDFY2LXqdfOA0EpufTd9
S/3LT0F39XO0pAIz3EFv/xi9ZUc4BqyG44KXWIiPoLJSd4w70Fbh8/aOt0D6+cEk
0FaipcM6JieqZ7xJjlxVf6ae1yLAqZRvi7u6B2pdwVS0p1V9E4yR5FkeHuexNT6l
sLB8b31Nn2jTtNKasg5Ph6f+qMzAhaUe22XzRbByMH+D5+DRg+piFT7gcDC7q5e4
tQ8VgeTetvDtEkWSKvuwGbqLKsnzxoHnXKgmhJsw3MyQ8l4cLIYrLk0lwgwSpp7G
UlrVIj3H7+VwiR2+klmveto1/nPKXxDahpCVqmjhkqCRECGab+MEgcuQ0jB4gv8v
8w3FcIFAgD+Jjp94YxthjTEVuSFA/dyg4rHQ4Tge4baEmFzoUXGnxcEs3r5LtWdd
e/rLgzLGvPZAo3E3hkQc/MiHTJ8jPKWo8xyv6jfIyb7H0PmGe6MqgL6ZiwNaBc/6
/UjPj7IZ5X/zk5HgC4H3OCaN1kb1f7fGLju6xdAVKy2pIOIff2X+9P0aGUXNo7lS
9bxzOpDy6hFQt2J/ASbUBUfxR6fJwKYfE2En1j2Vyxy4M6qiH4NOW5/CjG5G7s2W
B3H+MBPk7Ncy6uw/zLmgJEvzaeuwE4uN/670TvlzKm0Zx7hcZW+bL+FiU6vvAlCu
Whd/F5Uj+K/JGN8KOkw8eQyUtNEKJZaOA21dcUBNqM7nevEdPeUIZDUoo+Pgt+oV
/Wu0oS4tlRXqcSN7nOP0GJqO9YbbK/wDefiZyNM3KqLpH8xTsQG4IQk13UE5zqoq
mINvKpTAe973Z9iGeUuA4qxt0WtQM86P4byQ1FL5E4TCk+N0qsNyaIhQzqrS5EuF
Fx0yCN3RTkKzyzNHKeocZCkerRoFEPRE8+MTy7V7Uycmuvm08FibzdrKgVjG87FT
uYLD9N0gUX8UOMt1xTW+K9LFz0gNZU4ITVeTKadRFQt0lq51scqFh+zjaK7l/6g5
9q6gPjY+p6cFT8Rmdrn0BZUCo014qp3vWlQnU+gPh26BZzd2weESUnEiugGG8FOX
ay8eHtLseeFHd0dlgAEIUxSBvZfv+TGmHSGvao0H7iS5T22heqWGfb60bL8VZKkS
UGrrhMNh7g8LOiT7qU2LSUZrP3qWPvVlDGae9ToJfcdx3LACAPEZ9EvS3ixh8Frd
v21ONu5zz3pE6nC+WaUIBXAW33GJNMl/8XW9jUlppmIgdvkZN2waXiX1M+hlfQ4y
EiYj32xupd1WxZl01it14Ly1sOQtLxrWWD4bfH/E9bYHtc0jug1U+jy0QAvyp1H4
cvYkkXeJaCK3lD+at0ubdYZq9EHQVdOkM5qrWO/aKTtrafk8MfL8vVHv71W6j3RX
BSnNiUnEbwR6K5y4OCSuOoQRfJ3IKeKisy4tYGgov5uBQT+ny8+9OrRsRZ1BI1gP
yKD+sal5gI6jANe/59pPbf94H/xdiOHQpbTbV4KnyvgcTWegVnIWihbKVzeX/xL1
DLrmx11J4wXvsYCYoHb9yTyZga4c65WtNbTiObANfdLFjOmc0k0VvzAvHJz6ss6K
se42TGoyA20lVc0i2C4XhMOVhx8VCNaBaAnwdQy/8J+Xm6qwhAqImPHl1uo5VZ8z
dbhfQZ9Dpk2+OzhYnMJOE+DfXDiyhvMzuqln+GwCI5mb2a9Y9zWTe26Nndp8x+yG
esE3t9uiXnobdcELiOBpew8l/JPus1jXQAdBvDmGRBc4wN6bwHjdtJyUJ++0oxt1
6thsTSjDdE15okaQB6Id41Ok7ML841RZrO0KW7sTLt3qWIlHKe3DTq2j6XDUBuJN
edmMU+H0odawbg3ob9Sf0CxeObwr+PQjUduHSAgFLAMiG0RcqNX1K3X8XXnDwBEM
3atkiuiwDmkTqVoLprzuDZC2V4TzVEpvXz3l6LwpeXs26SQYlATky+hR9uyQBz5P
7U6XQb+3voMiZ0arBT11p6iT4IfzuNpsGE/h06c9VIkvp6gb5BlCLi9sQ4tJ0OFy
/eKiqHKCbdOAiHIMmZV74PEtO+YcSX+AyDGYOaJkq0EmPg81MMGV9YV54oW/pxkl
hKK4Ie2WYbOqXGoWVzxm+/j410WYgZcMlxw4Bp0Guagx6MUCpqUzOHn34bXF/qW5
clPd3Z5PEzsSm5GWmsb6HvnIgSb1uX1aLJUj4mVTu+7kOvNRFrCX4VgdCNjqRHJb
CPTtQY7wd5G1LnfYUg5ldm451PJtQ0VhMSg5rnZapyAAbEd46SjHG+R+rf3rx7Ku
krgBKRvKnW5m9UsEudftWtaQPzL+U1JINcUoGLbYtZ1tKeaP1w/PBimC9Rnbx35c
rkZHpybczGQwsVH731Gmd8WMy6zKnw2RVpvLay4ENavaBXi3hdhBTZYMq3pRHVpI
GslLfHNrUiJRHqrVNGKs73OSS4/H6mEOENJsthggPJ9VQGYpx6TSfGDNwfLPcHf8
1h7iGnpc6uBDX1Vhn7dWTmf8NcQw8S2rq9cq0ddP7bMUKPrRCtzgSmtxzvqyA/ko
bRBOn8gQi7vnq/5a07KtPuMwb9xLfeN3kRYXNaDCMihZYFMIePGl9WMQQG3t7CJ4
wM3RNgRMRqXmyGTbL2XT/9o/OK3iwR6ryeVi9z1Pb8AoHtO2toH+S60cw4eV+lda
SwSPylpAlRfH42rqbCwyw4e2mQNWdMRcU+LXOTMb1AsxDIBCR2I0FSPcbmin10L2
hXbxyrHdjBtC/cdTgWmHdmYgPcZ51RtoG9eEslH+nCWM2KDRsjUiRqo/KUTzgJuI
pG9d7vLkDUwDflE7x8+F18yu0EtOuYia2CwDgfPFVp8JUvoG4v8x+VJ4kJBCEwS5
OypywuduVSo7gq2Wua4geW2JeWLNxqXhB1iEndb73lhmVOlMfUAXinW5zRjcHPGm
55ErtaLk8Uo63vMjTu860OU+naSSknfmbk6tVyHMLIIsq7GO7QG6JwsaWDzw1YVg
wF2y6CkP0i+PTeLQLj7YFS7k2swYuG1EfNL2qylWT8ldZQMeVWL//InfY94R46yL
0axLAOU3evMgKX132o/V4Q4JpCif3CdlRnmVPEfKf26w4VKdBege8yYJ1/cI0Flz
g2RM2UpiYV/7pPBUAFNFheswNLLhrmzS3SIdzzr4KNSOpf16jPy8o4vQKcR3GhCp
2ohDEeIQ+giDie9/O31s7LJqlU9WJSgaZfIRIkGe2d+0iVCOQc2mCDoQYP39/UMl
9hSRauoJqkiPOjo2N/GzOIOh3ul1T0XuHyGdFSZ5da98WAE3OIBJLmhAPGgMYy2e
JCcyJlGK8Cavd55l+a2E7y4NEpm7gHgicEd/1tnTyw0bd3VhVmvvsRcUixDHbDsZ
Lswmhh+HOYQc94q2XAf2PIDG+IBk9cZC0baqaYov8KfTo9UI/bTinAAySyXxPOYv
GVi4FLWydwNXmKrtmXXMg+LLIgOeuBXwu6e+d5gd5ZsofWUSz0KAQvfiUlKryWnB
ZICPSdlHvce6A1qwaDh/YX/diR08SWWGbA7NMkRVE1MbUy/Wwbc5XdGbd7lazLue
bfNlR9ATsAvVm+Obt7g7C1i5RCpSQFp+xa3HREyxRyLgurI/l1hkAuPyuhF3ojvM
JJDAgL3nkZ9yF+ArJYeN3S18scxhhW2R0NbB6N6eHiblF7ONljT8mWVRku0ZO+WM
xAo2v9Zu/IBU41DNHcN6VvC/nN7aiYPyrfGinxLUwSddSW68JIapY0hzICZI1ruw
i2bArra4MM9CTK5q7AeqkkkE20OoQMusAct5yIlH+AC0DwPN20rtJAQrnnrSMbNZ
oDhzK51XwIjFMspzXh1EMTwFFQPaa5vb1z0OJxRtqHcVaP9gPdB1AGAnb4xHuS5t
NV1M3/7KLWvG0qDGttx9EfNI+rFiXIlIIdgFfgLqIm0Y+vAky0veOGkR5OOwa12w
PljfpZI52H1fJGxMthyYDxwV8bMlUvpX8H2aCk5J9aeN+/zReovnIyfr3wcnyzsm
ab4DTYs77/jZKcQ4uzF3OLvOZdvKMAztxptyaVzDSHfNwQuVJgXmazPyXCc+63zM
UqdF70K8uxu6zrOcxg8LBdp3fcAKY+D3Nal95sxX9PzenVBlRGyrij2MF3Pq+uJx
qrwdaiRANL4ROq0jVRd1nk9HCNiiqf2rB470mn52LIK1NNGuyp4b5Ow9GsxqWb5R
b9z6EowcMIX8+iLhtfzcukhOMvK78fDRtMqSVXZWqiu73HDG4NPZtJYtNJ94ZqUP
lzve4+StFgNtM9JeZaIP31J/aqflaXNTr5UkVkwrqimC/ZE75NzuaRUux/2Jnqnc
JdSTTuqTFOOFCU8dwydLfEBRXlmE4EifD6qrYgnnokgGFqTYW788OV6P3VPqEoem
xrO6m9JqikjsngYQG6CX7I6c+8F16dVRoOgqmW5TvVT1PjhjH6tKKW6KPL+C27O7
0bYHYHg2oZYW3Hd9U8079TTSmoDa3sxLg/tvceIsfPfzQV2Q3kuYadGKDJOt5XgV
FDDb+bVVJk1jwcVsdfAEeU1WlpyQi9oSmttm/7KKcWaLk5WZGTCnl6TLOh2Q0pYx
vSSuwNxa/VvgvT+gJSYu+SG7FDc8ChYy3/FOUd0UR3YStWYNrfXUqkkLf4pkfNB8
1pRxs881yYAA3LfIlCp5yWhtXanIfAQulVkK4uwk6ZsVrVzKlBXKZWQI7P4r+Xp5
/Ut5djAjAFm2v4xQp0aMw0ZtPDXainSVcwox7JEKtMCO3yZUkDLUOcn6BZP0zhDc
iPnGl5Ow0guq5pWxDhnvlwZ1z/8K66yEaMIKv1O6QW40YQzMP7ivMx+XmXsOBtQU
DhiOmD6wCQK74Kr4MqH91mB1j6CBqjBfHfwmUIjeMOq7t9Kvf+iVPHVOxCdbVeKW
pbnww9u7ahkeGGGMFvay+yhMv5PGTfqXus48RzK7drlLBlmBaov46nsfl2g8A/1h
rayDu7wD5+joFOAzDpUdxqyCAmFP+cNHHrMPJGKS3VtMQ+SGu1XY0z8TkbcVqczC
n5SEZSrq46dPMoSbobpAku5skfRQlqbScSKqmSWgxQMfJ8SCRrqsHaP7yQp7WTrS
iqWj59oZYXgMcUbMv1gg9blTpwj/6sMrdzwyVpucBMvRlhs5sY5IAur+vFbp3zNn
ua8nPtZ+lcDpxDZBNXkJz25i2mIvrewe/CXLvF6JxDzWn/cISqvya2VQ2hIT11fk
CDij3P1hf76g2ZfOND+BCuMtb2KeBwGfWVc/yiv3Fd6y8prIP8lJMdMRhsogo0Me
uv3PSWrz80Lv0T/3z2CNIfRUfzloWQ43PMwLjSSbUUZH4xeoABoNwA8vL6CoCHTU
da7sFzY8vYHq84EawlAmUSzGWNGCuDxVKkP/2/KFJSkxfS1qRkmyfcFh06V9L403
FJ562I5GTlIQDY2rizPXCNpaXOPuZQu0JQUbhdijdWjB3TMC7Zx7fWKxnRkIOzz9
hTMyjCDsVKWj/EzkMDAqqh6PloR3O+643FrXxkOmzG1H0t/IWHgKgM9H7rcsuvuH
nIxdXnYfixdY3uDuZgUKQ2sXjOIj46FYLALeZTdPavWj4/7uk2SJ+l22IaPxMy2R
bXB/le+7TGcQ+abLhAQy2wsSiWj4RFoNmKWYCZOrDPcQwcL9iZaZ7EhvjmadfrC9
XQIJ2xMJrxwTxw7GZZbKfwIsX6CDjxrc8kjZ2sXz6LdnWUM9tfWjA/3SyMpVhpHW
a3J7S1//aIOoc/z3aAOWszGLsq/Oz/jpxer5dyq0Luo4LZGGBupavOSv5RTppJqk
usxVmErLwyx2FpP2BKqnc4VrJWc+pbyGV9gewo20usvAkQcbC3TcruDZVIZekuPB
V6Nsm7G0hwX9ZjJ3ERdjGlmpfutr9EiP6H6/zfBNNQCftsVqcGxok40QleXDIZV4
m7sXge+0GFs3jom0CzUA4DFnsCSWmoxIThVCyqSKi4C7czvHu/+KgfjO5CbiiM7Q
CLDm4wP0xClN7jWbAt8N+Naz+n+dKt/chRuNnP5MuJRnf82wOhKQGqp0No3YCMFf
xxVdSO5aoV/mn+5/w0miQfPtWp0woFLuxFDkAmdJg94YtYNkw4L5TNhVl+45a6Ke
JgSA0EEqdLefCQ+daZPZ0MNo6CiLgmnbwm0d7ybOs52uPwzuQTMk0jNYhLCGfd/N
/XwfzYrwdDtPfWoIEqA/Lm+oU1H6u8PJyzA6kN2e+cp7aCSEL4OALsAY7b3JwP2D
OhkHI7Rn5qMFrpf3f/XNB/Q6YMPncHkNKILu9q0djobjA/3gBBMiWLC6dKbLIoZG
LqgIpYq0rcjy/plLLe1kf4cV2Uao1VvgMdw36QUP26rZFjFyQXD4bVImsiUnFLPQ
wxgyTUjyBoeZcCGbt4tmVUuv0bW2gpaJ3cf7nLx3SCS0pDE0hwbY4xqZyCb8BF3p
mJIfLsbXJ7xelrEduHx3ZKCUCfMDXtSyCAAarp8angl62FVRlHC0DQey/20NwwiY
LoZtnG0D+Pxo6IDSPF3Rl2ffDxmuQsi5lND/1Hat20n0SG+4FGW3QL+w3ZMflfxp
U2k8Re0l1t6d1T6FcF/A6KuYibnaBFlNyw0bl6WQfY+DxHUMeB1b9c+EqWzT+IS0
cxrJI0JS2WUprMk5ZZGMFSa80upDQ0hWciNul5d61c5d1mKtd7JfGbBo7uJc9Y+y
HBz92lsx1b56SMx49/MU4avaZfvc0XXHZ1PexbVI74XktFK03T0ExA4kFaGQaYWk
IcmEkKcoZlTE387Z3iQkKhIDnO8fmClcIQ8x8OceHQCKxXzCQpkOQPhO/aU2iP4O
BKc9PAw2CKuSj+QVOAe7NFjPrSpKWz2xL6thEAs/lh/ijacd/DKQhfwIR/rsirZn
JV0Lio7u5zbtCfiOpnCi9LnOn1PqP6MW8Ht/6U79YxhXbZtPyICIdzgJ+aw9zPQP
/EyPGByv7SbDFOEZnwVbiQzbx/07VIq2wsRUjAr1cD9tFcXSFQC7ou3GeXjVFE88
4/eyHljG0xb03JgwSmgqzI2Lfl9PS/Dlid3JbQNFztZ4cX5s2jLNPrTvmVS3LGz7
IotDiPBKEBs7UXTct6fOEEWvyBfleMMTP89AI9yNo89RwASOx+3yMTc2OWCy0Qfr
wonXR2V0I5JgotTq0svC2Y58bY+Krr7y+hg0Bqbr2313/Vm+c03XyMDTga3Cff/Y
Cb5SmuGXcCrEH9TZ/iF05QgnQUK/FSA9JqbYdaAuwlREVHtLCHzr9PLKWeOpPbyz
7lZ6Eh6YeTztYjlh4tA97RtyoY+dfWCH17zfmQff93ngCht0tAgWc2Im71M8MFjV
coYlF8xi3b8i8ZjAFtXWFHjuOtvZ4Lpj7bUqn7S5lhZWHjwYobPYzfaMu2rfyRZc
1HluTEesOlNiZtHNITaOmTXZX151egoATc7e5kDByeeUjlWGhaKPfejqihHb7Vdi
V0v/8AEO0GNtyeVSvF4OTzlz/RmFznpKGhqkWCezYVCXESOJRICqRRdUI5Hgnede
OrPyGvIBgfTYD6BebzfQUdQVRjhHvhpqagNOTMNBoRSxtiaezTQR7iJ5TugvGDUr
1XpoQqcbFDm9RTYRM/AFyjYgFPCzB1G+M727osT3tagsQX6Whf9KXmsrYQZXflOM
qkP1Lrv005dOq1jQaVaPNAdNqwqQE8DVK2Jyhif3tcNs9Vb25G7+mQkPj/7BHBau
NO0HfICSEqBOb6LjNlQAv7pDkhFcqcX41ibRUCHEyHlWgdhXetsx8mv8kjhPfVfy
ZkdTSuBKprfs9R98uY7yjp6o+P531UwmUjlnSVAL5Y6LLRlk07bR3/UKK2QfrFMr
KbSykLvqYfbT39ZYLv/U8Wav6oHG2g+7ZPwElR5zuknatoDHyB/Q/xCNY5le+oa3
jZJmZ2FZQyC3o/apIWPFwVCgre+YK++EWHsIL/XpCn9O+7yvluc90iX+PcPKTdta
CXuWt6cwwHdpLcPmcpLB5D+0BFSSR2d/Bb1El76q/dHbcJF/U5r8GCdzpA2+SH2k
o7uIemfqB+nan2D/mhS+iHn974veq7p8+KxnHIxp8YsdAsRZfW/3cm1HENEpVVYy
fF7CX+LuXZvZu2tm/UhJv4d+c6462FIoQcfEGDoG634zayecsZVLrpJ7OlM4UDbu
8rhYinL7kqwS01twI2vb5VS14rhMdZIc09VoS2zu9NwQ3SjOpYxPGmqc/127/6A5
ydQT70i3VNuqE+hciQgWz7sn3XJvF+z2CM0zSY3EPdQO91UgrD1pMuP6Ai582yK0
x3fjO/0Ek6txr6DGE0WkkG4gViznYBVV1CFx6SnQGL95dYdYjN1Dx6If6zx9rcPc
ZwP9KstNtCaH5G6hDnE63rvBT7UE27y01Dq0vDBIWuzLld/m/J1vo7D/wbeJgaMg
S4gj4fLceqxe+qTje3uxQnpBBWFSL6gIn1NTgYIEJXQ5wYI4byLe5rJMnWQOy/uh
cKfcxM2rDMMUzKJlYY3WWXqPGVYugpbnLSrChEcMqjbeUKXZTDKUn9Tbjd/xOhrG
Q+rdZ1BclZ44CTA3pc/gSKLw1AqpqXwYplXiE7Ak0ahrG2LzDASPSybgb/SD76II
i+rDq6eB+AhX4yXD1eajoxTSSDkLOKcYHfo6I82s+MHhvHgqchr0oS8vSgJSq6/6
fn7TdMOyCIh9H4kdJNe525QhzVMrcg8ccFizFql1QEfUgbRf76ZMxJms2bcUYG/S
YjnzrIZ2tGE3oGzpPo8/Cl/75W3uwUdJ4vUnVNRolZ2LgE20Th3H+g47z7Yo4l2a
PsVvKNo1JhtEudJOmFnriH0puXUp6T61OyUlSP7bWqBcJPH56pb1zLooTMWpdmFk
BgDzIiDNOAaoq/PR7MmzAphrEuB9/nSfJst+Gq16iKpV1Oeoo0nnX0+b9IL+cs+l
aPGpUx4YUjhsaeqzjVAswGL7SKCFG5hGtrTPwELwEoNiM8uPV7CfH0OSBUv7+T0d
toHVqdmSlJDsGPjKvQiTlYqjf16rY8eQWHYPa7aw5lxhVF9DlYBNjs36leroI65T
9DSTUfJCho5alZFp6VJklhTI2VtboYqTQ1O+ZbqTUc0wV2uh+MkYW6Y8Yv3NFNlb
X33B/TCX9Sed8Utfm6eOEHuF1BjLbNPQpMWD+K2GYrqKmxkIaofr1DbvQhBiNNe0
M1L2xJEhtQCtzcobiEPzixs59p55MnjRaN3hiFx9m5s1fw8QeL7oux7drHf/ITFP
PlWbHRual1QxJDZtBVcOPakJiHtuYNRAi/dA+1mVYmQqz+txC0pklA4xhSjy7cA0
m8jFG5ccqT5mliwm5Cd7roGLiEDMpe58ExlMakFQL20eXSWSQf/RiPJ9Fpu8zChm
nq1ChCJrm8OG+QZIajAz0PnFVkMy0Y/2OiCtkjudIJ4ggzsaoF7jW7fY6Rv+1z4w
U9un+tIf9z/snsvI5K9Vw940S2ImjfX0iUGsb+qxqT9nrUFOlZdWf7gIMTeC0iGL
VWHXPmnioNWtnPx2A/3jfDaNRp+Tyg2mSnpge7xWTGe7rQIGYs50GwC22DFtrV6S
ysAj9tOAchTJE6HGLLRXRM8mvRREK1yDTKM91cR4pdSzc7A00R40OD7a0Rn7/5xp
0yISWM1m8sGsxQV7fL0+w7tGZRJ7CmzburiTDr9C9GHn1CM0jiwL4SRgEy59/ncL
FnvhRh0RcdEVTzY8QpXE1zapjG/75/5kvs7eSG/ywWCOPiqIEQ0BMZTy3HTk2qIM
/VIz4RY3d+APfX4yI3D6vHHovCk6mVRGrTzRqSupkx/U49ENwUcNw7MJYm/i5wW/
6tnHxueCxH+TQv7Ode+HglJr0xJV6KjHipj/OakLMT20CLakEcxCnaQEILhXfsDk
8J1bz/xuFs/rMQpAhBA34H1k/5j0FnUGoWVlfozRWA3sxDcm9mGDsxXavbsnrixw
Szc2+phcNqaV6bCVigPDqOxOBrirKWcipUzzkLQOZkTuCvTpkx6gVS3+vOreVtjC
ROkFoBJj4iClJzeuffGaMlK2rcZbuxpuQFUZHPg7Dc4KF7S2eQScq8BQ5JIncuWg
X83MXRp7Se0MIYC0TmqbBHYsMns4Lnd/F78IHWDOLNe4GZQ26PeuXSUSjlq26Zha
iJOObtFcBlZK/vvC6UuKt7ZSGD7kOqo6HuwrDg34u8ULU4uvzV5aP3H/mUItQf3a
8mQjGPGH4MaR/RgXP9ICUsoVfm8t96EI99VYTAfW8a+uwwG/uvisLccwAmtQ9zy0
cjVA01AiZVKTXTbDYST9dCnurm4bAEXpaFrhSanPo2eyGlHxbEYQSYYgd3r51om4
Jq/0ExwQhr2GTjXkF+Y4M5vjevadU2W5vWOsbMSA0/wzHClPeHiOX4/76vWODFl4
JjP13lxBkPjPnDyywYWxGArW3u6dy1+4z7+s6zsB7tiFM/jwg9JNyuUIJZ8zZqNs
UGo87LLUGD3j42TakOcaju5shb18sKz69y2Zcii+LYvhso5TxHxgEz0NSzcHAf8a
DaG7TcIp2RpU+0Cl1EQVsE3+YRpiTbGZPIWd4PkyNhirbgamTUhJPdHeAcYh2KDp
O+6M9p9hRJVLNjefqjjBAJy+A6IWZtKLbVFxka4Kb05Cj6w4Di0SYj1Nvwq/1UhT
m08IZ1b5Pay7aTrLSUDrEccZrWeRHrsGxn8PKi/9N5UxQMkMw2pvdweZF0MbB3Zn
dKdoq2s5r+jwcKvUaedz4sxlRUoNzcSw2uoOVwF5Vv56ME89rBd0tghAdyuqF6a2
ER91yr4SusLYN7YaYSc+BRDhzNQH93PEossusZFHEu5gmJ9fkoFmf0MyAUCHL71B
iBwsDRy8vNzcxoHd6aGk4lS3qT7hobw3s+nDZNw0J82Yz1zQLCVACMbYwtC1pgP8
KRqaArwmHUBgF9VHrLbEs8heWwkrKxzusy5VY1xP6L1CWdT9kiH34ZHhs7iyWvzJ
ZWh1Fxr3V1fDOVpMChgmiEWUsC3XIE4F+keseaIwrN+FBcvrGCgSaiBNebv9Zpxx
eNUQuOaIkj6KTNxrodBxiXNPtej0cFrOL9d+/DsjoiEVuZn/KfZfLgdXS3h0sAle
SAKxgiDZAp88INyy6AyhV4G+QAWmR488QH+TJkGLKpmab2fmV4kvXqfopch8C4HS
24v1P0iXmTYN8VzLyIz0KT6zMeiy+ftSsXTXtEkslbrlEC/pOxUOdnkUsoIGy9wr
jPwFhhSMwyGr/nnkHrZl5pH/QsmRKKKRqAXZZiCvYx5GnReeLtYj9InajdvX1X4V
De47XnXonaSd/mBE1OjervGqY7jSV1e5Po7pY+4f5q5MD1MjYDhJWBY9bttJRaMJ
l85zjD2D30oxrpFg9RFio6kDfYl26lAgtDTt3F6caU9HSTWdUgg0iZYjH9WoAQEH
iRyuKvor9wAC0GOr2Kw1obHcBr/zbmBzxdiKFZ/63IoYkBCFk5Reh8tCEQ5vBRwc
DCd7DwaYiVMiIAyeqZ2UMMX+5dV3x9MqFv1+yYSEaRm81BrnGb+F4qZHSAJUPWRh
ohfFaAAsw0nSCc+WgsAZmNAAg100zYO+NYmQok7W1a0GBlsxN/EcQUL8eeWhJyla
OpVsDaWLtgMxK+QJ7WiNsl4hwMpiCfxs6/3pEzxCRRyiwFLOX+YHUaIDCaJXkMY2
zxFFi2Z0dvQuLLU8Hl11Swt7hdYDByJFpjbfmvkveaAVPQld3jj4SMyzO2ANjLvN
CIHbDea69PAFPvyCxidrbYpFP97dzRukdEwSIfMeb72W4xw+wZRnW8Zm2et0tTs6
nuYI6wWkRUWCl+SauLr5Bz/9rVt+Im9g45JDcehKO3Anj8ZKnN2xeu1RofBvhPoA
PN6lOnyV3I82o3pIm34h5KxtiWxJuAfSZMG1rq+0KpkWivuDcjP+RX2aQfFuNSvX
XwQ0I5ePy00LldsCd2Md6emrGW6tZtCdMkQ9GulOoULgWQjhq9Bd0joZGVJmReFa
8WxqMj5GXPaBX3Z3fcmoTpp72rFstea8nGYFkVMnJGVl1LjFFww1hOwTBjtAhAP6
2J/xHDS4M+mdNNgVpjxzttzR2uh4YFsyNjmYrqf8sJWdUTVvZ0w0GmY9ENfYR/3T
o9MgJsBFkTmbMt7R78sJXx91bDHd20F7aWwj0omcLCzshZh/lYCJ2LsLy0OzxUfY
3hfXm8Z8KENmPVzmrkXjOg/vyIe6GhkfBTk41aGD/nWE4ho5zRRsILJ4iHUkXsWg
IsIVccn3SI5EcUCOBQJ6sX+MUaYz6Slyg9k4SRyZN9l3zRja/BLygXJEkqvNkmDL
kvAjcbdVIObQicYQ4QISESJOYxSVf1ro3HRnnxrLdHdlNvQOfVe2WB8YNWSd/Izm
PoJq+1z1XI5uDVGSMXxDMbhz541qypg3UIRpbaG/OIauBRVH0tEqpDMI2fAuUV0I
CsHE6GoTz5gfU8tsTM1nobvG94wHoBj4GWxEl4amoyBvWrVqTWKo+s6pdoj57aUp
K8wfEcAYur0llIQALu95u9BfqimIWDggGkkxGc+rBnlfGt6xC+hMrtu75gRvTaiU
ku3Hd4sOCoY5yTEQN7RbWJiC/Zzi0DPrOxHjYmLU36YZDSg72kTfwnlej9PWf9aT
lrp5ZPc72ZHehGkO/9oA3vonpKSR4X2J6xx85csPUpYS73ObSnR/Zg+fALgmWyxT
9uT30UkYSCN/xaQmD0HUsonnm/6Gu/nnyq/K86QwS/zX1pa0+/Q7eDAdPM58ZBpW
rwjfyZ1xCNmr5JEARw21yCQ6ENgXxUs0URzBcoFM6iKQSf9Kw+Ki52o3SKWIm72Q
XofI9VX0/GuxLxMRmZ8j1t0xGAzF3LC058mJUlOifUeZPmYb6dDVSE6byMNjX7yw
LukH/ljS6zCNPG5bC4fFURzxuzgExVLjZmXengDz/5GfqBsoQ1TIQO3+6UN0oxOH
GocQk+Idm/cfFeX3rF0jfZ5XSLM2VP56DEdI5myACxtGx13L7XbAkAljultULHxh
Ra6V3p4RmH4rIzbwwQO05hjVB79uTZprFVGwduUhC9Q1cIpvXZyarqqcjuCj9o+n
CdQQtV6B5LMXgYjx6ASeInkzyOYYExcdJWue3Yp+yA3viHN9qw6m64o1kwicqpLm
4wjtg+4Xyr/l3gEM4Hde+398Lqlv0e4xlOuBgiia23lfjA1VQt8zpQ8I0hmXWgxb
u8GHb7X4Vx6rsRpIAdxd6/CP+PnC2Qw0Sf2h4ayIKbEto7TyTiaQyMDM5VcVt4dM
oyFb9PAle1vr2I+bjSxB/VX0cUebDCA5RDOzaYfAHkJ3owwzos6/KP2je3Z27w1f
7Tw3d4Fcg2QMJrdNugAL8C+KBvHrbjjfXtFMvyevEPXpDtE0s5c+pn0PstoK0rH7
dlAtKYZhiauOvEA/4unOyfy6N+kTlqKHNZIex+ajuahix1xvHXyWCiu0jr6qxNW8
+Bnkm14JYUACoGrUmf8JL7uQbsg6Uh3YsPPi143pNbwWI8JGk+pX/siPEeYFBVB+
VXeBa3f4cEjPieW9mGUMXaYm9ZRbPx4COzugSVlgQFRCOpuZRpChW5X0AuTQSWiz
pkbXkXSrO+nxmBnA3lmqRwQ7BSc8fydJ7Jv9HPtEz8PgozbfOa6/V4MhltXdghj+
B+cWa+bUwt6QhQQIK/g1jwLcYUllGuqJL8YH6G7ep39AQCj5N1iVYM+uhPJihgR2
OWVTcRFwgqAkOfLpAcS9oekc/Hs73FYIY1ryLHIHEr203kZnOOW+pOgRoY6idTuM
1L2Pe0GGX+m1fGE/If7Fuzo60ggTO6jlJUd9MKv8YRfwvQDs8+Fl/l2R/J0nme+R
rs9i2A4OCJ0cXM8tdmZEgmopCPduOwh8dSBdoR8D+ORBacULOCjDt8UafLdFdAqq
D8MCfQ6XwvV5HGOovlbvPxC58Njp3wgy8huyo05tQgjcwf/meEfb5HXnOHTDT8UU
WdkWrwpnMT36cljQZOaYWfgt1yNEGx8qHemrX5tTB4CHQTebGWqLvH8AQoxUdvEQ
aYdMronEteNW0OhCchei1fddJocQp+GWJkFkxX2L37BGgdu5C7UVptMyIEeThUXw
aNABnX0mhxTHrN2Rynm4wxCuhhXH0M9lIjz2vIji9SPbTIS0Dy8dOt+a276KOxuQ
xm6HayFNHMLqCz2xd+oOV1f946e1eqthcSRIWUBJViljSz3IAyIGKo3v8gzn6NZ9
CNJMVkCQKJUiPrlLwSiPijdhCv5Gzg5q26HNRAtdgKUDaohiQOA8R0yQM2420Hwh
GkI7jVRbJzvOqRFAffREqYSRjElb0uLdH6PytNB6tJtctX9GdpTCuXNyztk8gJYp
7NQTQnZmaK4xrDhSwlaZiloFg7W6+eDpqwVwTaJVqrcaMaPtitM42xcsLk8GV18K
Iz6namvqiKcrfhW7vTEFALaC5XoZDigE5YMI1Dfy4tg5IY1OQ6rrALonwBngiJHP
cRXOm8F+g/CnkBKCxC3s2/cXIYHt/3JxmIq48bz6YIIWzlsY4yDXPlElzpJBimn+
CwtUoku2Y/cti5a9R1RoVkWRZYudo4YWlkSLiN8EgrognpDLN/Vd19pbpGSScUm0
H6loBRAi+KqhgV8O+lp//z64N/LQWMpKCt20U0y2ljAFKKpxBWZf2vaFM/w366mT
PLVSx4htpWOYu+tUbmROJJ/vnmoLItZt9hr07Q1VuCi0sCdGN5iwlGM8qMjziehX
4y7yObbzuzFBzs4ZcT90WytX2NGxvp1xSNeOAq1K+ZEhLGcil7qgHg5qX/1C0yv2
1HbXK1cacwki0NQShB7QHpuRmkQW9UooI6KGmaxBkcke1cpnbcFEpJ64OmXaupPx
unKYE+J/zXO4y4kpQKljjfCekk8hCv2EwBtzspkBWhg4LW/2ntvS98XP19fVIvba
7mywvtx2gr7N35OqnxbMiKtsSFDGmUBuS1NADETyyYR1+LJ2oZGKH69WBhAeRxGz
r60FCJQwZrq5SmUM2YKyo7TNIfB/DpQf1vaCFdcHaRiPhrYUjgFbKi099Ff/aB3e
PltXMmwh4EkmAdiML/V9yWOYIr52sFUOvgwRdlG6DA6yrCKylI5G/1lCOFpoS8z8
qkAsE7usfcBmnEgZsGjuF2FYqdsS1my4gGVlH8fqMyK8cB7SZ6+T1SQG+TCRAyrg
uuoToQpPNTdcfmo3QRzfrGEchMamSCTE2fHy13o7bQsn+2etoA+wKctijQdXHFPB
ZlRkjixYel+VLAIBbBMzR+/zrGXOVMjHMi0LIyg8lEuD+ciYHvbFTN+DZ62IsM47
lMQJ9zzRNFCYmKEn3dbdmvvTHmZzBoiykB5+w739JjuEBSXnKmyvmzpE3zKiUUTl
vdbfGqtgaSyd3HKJOBsWauo/mnk5pJDtFVjOHKPJ4jUPEOMuDhMLmV3Uew21NJq9
BqFvNtntIikgpyh2Lom/WaQgRzh5BifbglHvp9ujFHK5vSoG8CRsIYskjQjqMymW
+QoqSGuuCkhBngyRlry0mdioL3C+rQIeZqV2Su5WnA38YU/nyhI4/1lJR49xnT01
zWAS7SeJ0SzjN+bOTbClvNGWJsNECpTIq4Eqrx6sEXjKDlhx7XSgKaXahdG3pOk5
RjR+/kej/rI65JPQFcG+08D4vug+jgXm4FKI/29bHZRbgzL7kk0M8vbXtWsnh2sT
kpDva94PQZ6sV3nAptX3TeIvsaRsq1BDc5xa8Ri5PtB38+meOcyvKp1xPRt9YkbK
7tgDu5Xrh0n46zlfgCzL6rpclIK/b3ocD4RqtDF622c79UdJ/GpiT4p/E6Gyajs4
J0LJvmmdXctELEDXW6FNak95EdUYnmt6AzXhoT+e7zfvXfGeB0kMd2hn8h76dRI1
EE7pnYiLHqcKON+cTc3u6ZFPl2Mc8LcLATN5zOA3f9O03M6/lS27y3K8zltk4Ita
7qo1MM1WPrT5NvLBT3aRQmkaCBIKwCX86eFqN8KsXYCB3mxzvCdmVzoZV8PEwUlU
kH4xoAkFPN57Lu13CCbuUZ9uuyWlrRsen+zH22H6jHwrF4q+px0/uKuyDRwNeNGa
iOEhvVi9zwVkV9djjDOs1ZH2jnvgKhA3IFRERQJTH1y/3LBcq9A4bp44R+vZ4QSE
td7AXo72Rw/VF2mK9prjgsTULn39rJGyd7k3+TcxTH5a4QeoHRGo8k/grLFpC9kQ
VQEC981UjlBqgEIr3KNI5i/rRPdHHh1V0ACGksi3x/Xt5+FaUWUSrjSy1QRKP4Q1
v84ALq9rTaAnUNbuH2bdIv2LNhuPeupYpiqlLoxTaGBKMk0oMYXtgeKKYqTGAHk8
WlOkhzG1jee/mH1dGKY4lOQvoynHstCpe4FQFU6hGBNesgSPwNB6fQVI50vLEZDA
PUOo1WxdRCMRvMbdhT5UOg8e9Kcwx1D9BLsnQagp2tjuk+A4W+TdqAacg2qYT6ns
tWgmn4Ttd8QIo64n0mQ++Iv7aGlPO01sKSJaPDLVkqziG+YdcLjfixDCGbpi9is7
W/hGAN7L6jLT2du8xGfD0rM7zHvZYgYUWvAbuBFciyVKyo0FMCL3Amk7ZY9/z9Z9
X0BOTfhuolLoOSAgmgumDYVv3Ooyo6cDC7PNSdV6f9iT5b67rr9rDUbvcK94rBHv
E4dUBJTcciI7Z1q2nW9aLI2NTpK+6u/ugVAXOH7UwCLfWIuom3WMqlPAOupAiI/I
wKzQhBOoUCQJi17Wtbo0SZbo1ROYwGBymY82J6VTRub6XgKAvcmX3ra83MoiQ2fw
nR468MkibY329aLSfdZVVGnevn1W8lT/z2Uj6NNDKNeGVoYTtx0s2Tl1139W+puV
O8qa8NyBOyF0aGB+nwGrutrrOCStjV55Rd//TSbiLhJIOHZoe3A+7dNHaoPa5GUQ
A4fhk50UW1ZQQqK1TvZS9AxG601T3KEOocAahO+kULHzgtH0KTEr1eAJHYcuedov
P8yuV9pKFs6gPhMCKZIk7oN1jgVCRE2UHmq5h6Rkcns9My8w3SiewKP+GU/HWfV3
5XzENAPDd6q9uPBZXA4/jUT4z192qt/m3b3r3hQmFsTVi5J/wvK8WsP942GsVj1Q
vxDz8F2Q5sjwoMsbsX9DGpsqmcOlGK6St+9IOcXO5PTlTpJkxbQqAQkfRbV5AVOC
MfuAivp8zDUytfW7KxmPhTx4XS+zO4r5etCna7ogPFa4xk2xxovx/bq6oh9T21v1
moB1L99RxWNsiNaazOmw1kAN+ASBOleFlmnkBtqH41EieXgzNZZ5NNhwi1q+9aws
vxJ9M4zjXeP8OsyMjCyMJmislNMlALVKgMrLAjMSi7MmrLH3UF8ew59zjyu2st4r
gr62skNKrcRGnAyAJdf8AGlG6xsUxSIot2Ry929APbCfAHIa+zTWnuIGJrYQAArM
SMau3yesT9xq9sUbdIDez4OqywxQHkESaRnWej5Dox8UB+Kx3n0DyGHC0YkKUKvM
JZncwzvIEd6Hn50v2LcFfzj0xQWO9kiFuvgszFpBDsb6Q3hY7Rq9QozgOyt8oylY
OJ0S0bCkQY9FsQi/ieyZ6b7K9hVp65gRvHOAB6qpWz7zQMKc3ZIYFfk9La9mWCiz
RWd0lBUTcxuiFT5A+mgJenY8maj3jAaS0Sgw8qsi47qqBtL68E8oJzON2V3RrnTb
h4rnjLHXTgL/9mmIcH449fWVyH3y1uJ5E+BQVRtJaH3uwz3Dl9Yr13RiX7x2sq3W
XwLJoeH9ydRYqY5+VocsVn3IX4sNcaX/mUFllTDiu2Le/JXfAp1pnlLJw9mMCd1J
lFAnD6oUtw+NrtvBoukXlbRD0asYuxcO/G7W41q39wbVBGoadlMwsxVzy4UcQAGZ
m4Fslp31WPAIRzejKn6jxca30l6rAE6kxgFZekelNO5eWv467OdwWD4L/IwTcS6x
d/z1HtU+7w/5cjqFNLgl/+JQJntc8jKLgvjBOBvKSdGCv8QMCbGthubpOQzjs6s0
BM8dwE7zqwEWZpYI/Av6NI194LYbC/5qK4yFDgPkLaWjYX+e+/ubAbnsiO/AaTRd
jXQRtL++dbWjfpINpqDIdsJIhSBFFxOdNR6H+7MOdFmEpg19OHEDCsNjiG8mcNoP
qrlWFjW2T1ZgZHvwowX2ysI38852wPWzAYWkMmulJOgxm9vFjw+4QRoB0J3uZCDc
38oArLTcBCxyrytwiMF7ya5mDqF9H2efNc0T/2pgcUBV/TCIX1yrGlb4GLWB8PgT
a+kDeDyrqB7p+x9qoD/pSh+WZVqc7Bbx8mfNp2/6Sg/0knDsDvHfzSIJblZkTLCq
rv11Kgps8Z70xmrx5BIrDGF09lnQW5JdwEOEw5K2MRSlab35yKiEyUW2BTbcXuZ+
T05GCjqhMmeXsARZWORyObw56hElSxc0f85V3BA6iEPjhr9o0b7mLJCJOQOUdrCZ
BYAcGqY347Ocn7EifMoIXE1EQQrTu1HBd5FQqgwEa4NjP4m8VrVshvWKA2bvjHXE
3OJmj0sjfpvzQF1mpxGK6m3gEboBLN7M/Q2eA2y2iq80yUetm0FQxJ0bBIBBG+l1
hoLLI476KDNkX5dAMqwBvrPF9+Ytuwpfg2dX3orOjhqHvTHBqf4uCTrEF8Vw7PAE
8K/QCpXnGDcEuphtGkMRbozHM0UzzROB47UW3PAMu9+KZ//rx6alwcAvEpBDo3Rz
n7pEBsJHhScCyv3EtULpgvx0hQto9gM8HC6W0TkthVo4ixZ6jfgyK1eMvVhGvHvB
icNVNB5qcUVHz+KL8KwsdPeLxUwUd++oIhJ439oI18uGBhQFL0Hvx2f4YMCTPR5K
/x8o+GmYGHAe/4uKPaIgFz5ZIYERZgMK2Mg7BI83tBHgIKUF7KYS9CSzlybPh3JL
muGQN4oD/BoB7zy8Q7J3Qph6qYaTnIrHM3cWuntDPQ3i/Ipc4D+Fe0VcGGtIFRwI
XrH1QU5E5cYKhd4SERqj+gbzJToLpjz4I3sB82n+PKt/nj/18w5jNUSiqm9gpjNb
lJ267VcTn7OwOFg7ijP3YUWXxAH5tSAxCsLzALJmWSuz3666M7cG2XXSCfDieJhN
0E6wrXFCiuyvYU3JPz3cxSLsgrGUP+N9SeVUZpESRN1hgaM7QsC6vi74KczCZOqn
5yAGS+k9JNb7slkzo5bPQunXBcSt6T2nyR8qsSedHAIlNXheA+SxRb0mzLaVcDXy
BcJ5EXswzEFzgm70KyWzVjWid1GdVk2NkvEqDSaZa0LJjKD0FcGAbPlpLvw/tEzK
O1MSUY0MPm2jQnhyJIRiEu61Y2ooatIWgdQA6WPtW4cliREAqFL3haP5UUmK/55p
58DnftqdkZ0nqiU+fuv4nEp4meAzDz3pnQQ+ZYftQqlphHqOY3GNqIapCyn5liPc
xdDOdPfCwwLNve1mzhjNAHHg6g31+oXFK/f5BXk2HUG5ewe6gEXs8TKsWok35tEC
aK/UAM4dka7Um5ALK3RAaEBfkGNUdxpfM5tgprUrrQiKHmug4KTQfhEez5bTCzzR
JXrNx6mpHVy7Yh9KBTYGTd7ti8ivr/7HW62pyvauHDGYa0SpG8zpKuAFM8IjVm2J
7BQ61y5tx47jQ8nRyG+iaXxI6T/RYxNPPO0acuHsiFCyX7PDwGr8FWGYpb2RRuyK
kiraG3+vJ0+ArrP54uFwXasnUPMw5B82CnK9vjQxXgTaBUdWCIti/zBJ7r9Jlrza
FGczwy7xNYVHUJG6hCHedThYbWH4+lzL6sQBZo3yTvi6JK5A+MYrhxPPxlHYyPob
dRWlP8N7birgV54G2jkfE1U6ZKaw108+xpKzIkuEq2LNG+XXHbKEnuZ+7KOTMKPM
gYuAWCT4z2gJDteQq4OqWF0BOA3NvPpplnk3x2IYzVKVL6Yg5P5I/adRW0jhENig
Hq710qHCapUtUvYwACO70ToMri/xgYDsfq7j16y22KJCKUK32H2rS0Y3D4pCCE2q
SkW/aIQ/3FnpBeS+AdTFqO4TD20BqKRfLVEFmDytKNxvfQ7nfmZba6pepdd+LhJQ
4rvKCqEqawaKK8FHqbuTFupslRIDYLr7n+fE0kaXhAbeu2BkF/kN7JcF1Ei1aDZR
p1NIXg3R+zUBVFf/j1HklcdRc7RIul4rcd4TGAZrWZgbT4++DWRu+mUsul1lY4Ya
RCrPCEIqHPtVhQOdgLbHzQP3J5yzVF0BEJwEZ1gvL2RVyn+hinesQF8DzIFI0Pua
44EfC8s9vLK6OqwhIke8SlfyGq3KvXtmjktMSK1nBtkKMZDfXKRjVrscL8GF/GMP
t7ZovYeWj2IIyTnSL6QqWDS0qbzUqY6s3zBnmXV0yIKOxtxcBDOARmC6AaviT+ws
NXisUHAIXMS9emXfYknfs8lL0BnoDAx9MTp94CoIoZZ0i/ye6RGUcELjXM19dgJX
Ly7EQCVyTC2coseNcfengwYkOgP5euAnviAf0niMgKOkMaK83O7U3s0XuoiCeHJz
vgDHF2Wmm8yurEE975LVJCKifotuSbQd4EBDvyag6qjMNqWLn7XhJ8e8NPaoKyXz
RPnt6pM+OwGC4h/3TabJIlb33l0i0DkBxNT+eGQOptibLpfMCgHTl+PM82QE/3JF
0Feb3cftKs8xULn5ZYxLrwU5/Csg7XJsKG5RDaCEZxLmku4jMk57rPuUD99a0ll0
UtaE6owsxD6KKDkRnDXDb0tAAklXkiFfjlrljxHg0XNdBvQf7hM/vAZIe25A5s3o
yA86rlFSOc/KQgvrCaNYbbRIiCMq1H0gEJ6C1kShCCXV/CuUwiWxiC7YBIQNO655
h3h4ySnzFh7CiYupYdnotE4joUHcwV4LKmlDdymk4qfL3iYuZ9zIBsx64XK5WkIU
0smkxzstx0NWrHo38g5uwVeFzg5OEFYqRtZ66hzFbUoxMCo4XP0ovU872+kReq0I
qKICiQjajKwYHABm16lRRdhudGIpzZTr33P8qmxtPuRilYp14sxY1DiKbURDHo0F
QDbhNJ7Yisz9fVukdyWBeTqqd4nI5CDWcTnQ0fXbeJa9VTS0SVg69w5zW3mGD2e6
ZGs39dvfS5cwPyeivKTkXaPPHSSyFBvpEc0MO1wMImerEzv0N7DMi7fsjSpwS+Qx
3jBwxYwN2WfTcJpLMAisGululGidl6uSdQiudQ9aYywlSngBJJ0aG5xRI0fNc3kc
yJy64CrM6aBt5exrjgrDpV0Y/UnDDujm00Nv+Y4dPpIHtGMPFCfqp2E8gA9C44DL
sXUNEYdIDhUb8Z4dRWkDKwyqWkj4WV+qhM8dcLN96N1PVJfHPUFWsihsqcAJAYfD
OWT4fUBGelmTynrX7OIZQWtsRkroFymCAZ2/U5zsQBBsjkgsMtYqaGezsO7b2mB1
D0r9ijV6Ag8KTPqXnXtRKlYwBHZG5huVbf9StvXEjFHIARyq9jb4AwNuZ6kX5QUw
OelOwHgmi0N9fFg2mqh1FibAHlRhDdI49g6I3kb8R8LBXNDKtOvG+oyHDVQCHCxC
ZY/ElAtQh8j3+Eg3vMv27FhcN5tXckgd0csVmBunSIPn90+Qb08toiEIInes9Elg
XzDiNofh+yusEB1vzx80wCwfPhcuqbXxd7OAoOQaxuRaGxvMHYGxxZAflJavBHGW
clt4iRQm6cFnZ1UN4tQPoCATv+Z3cIuYvmOXOvlZC+MaUhkrpTD5PnX7WFqFsSor
YCdpJ7zrktrvam7+6dNTuL9oZ2ERFuVRWeOgarANkBpNqjpKPYMm/ZNsZX7gH9rs
0LIc951/BqcFhfWWQRhiwNdtVKsRHt0BLscQAeKqatTk42IJeT3Wd09p5lViHImA
ip4RZJlX01yPR5knJPyeV6WKcwgoUMvcnAiicyIpe6FMKhcw3Yc/F9yALzXeLlm4
SmrCnasobu7ssbEltsLX9EnzXtKMKKujscNnAxuyahc6lLLgr2aReVJ34pZsRpup
H9n4KQoCYS573UulBS8/3wHcm8s20OSZNtNy9XQV3dhFJQRql5NCzIyDIZDZ7YC3
pwaAoVt+6cLI1AsOgVQzR2tCDo6F2aDourxui2A58E9rgu2Q6bcf8bAJQoZptNgl
83fYoAa4ZYqyEKBRYvEDk3CHBVDqIsb5Sb9yuBnjpMmWB3oJJWdA6eaH7QunswvA
BEMKgIY7RnBULNHGMCtIT56GgzUj4Nbt69OgeKWc+92yV0Vq6Hvy2zsvrdZLqvLA
ohHGAEMUOT4KJTPDMUaNBQ0xqfEG9qSiB00dk1CgIHVAHyfuijym+KecPhhM1euV
jcM6li1XIOUSvDCtzuHWR1uS6EXHASVSAhMdZYFFwiGKKcPZ2MJiKdJLnVjGQsto
ETxumMXK50U6r+zqNURoeTJB3dHUp+aux173UptGauABT0hD3goU4SyQQCIWhOsB
0sISQIFU7P1Du9kTiZUBBasPdX9b0ZCeT71xllROkpc3HfJPbJp4iHtoBGkW4auK
xpxu9htkSr3dgvPLbJtah54ty9QIUdKijFvQL8L43uhANnVlYQrYPpzcdTexWcPM
P5rwmrNn6zCOG+QpY+bA90N+7Rtxxm4zY9Ur34Ux+1zfY8cJBQCpRf4IP8JeLP7d
F0badOopU7rhD466IYcbOjZGrKBSkR/lar8FlQf0RrmJ+MSOI9M2hWkUuTBnMNvr
LdWPmNfeESywW60mnHte79OkplL1bCxlZyuyc8EUZ9rR2wuidsWAFgejTSZZLyq4
WYkzvSG5D+hMHwjXWrr22hvLp1PV/CSEkg7d3zzYtHsJcP9hZ0VO6SiuTeSKgwSc
kGlg5FNxtC4jz5IOe1yF507/+M5KCtdbcxP5XKW+A4q3DihHUyGEiR8R7/hwAT0v
fcnK3bHJOFxQykrBGSNQXFhvOu+B32ySaTaWKPYTcm8SAMMicdmZesEq/pItAQMC
cJmels3mADPR5kCX5+wWoCZQKxsx5sy8fVODxB4LV9wVGTPmeexrS7AhMjHz4kDM
RcBy9ACMespdN7inUyuZbBcOuemMDbwNJ2PJVoSoo0jWlj6wcs/F5EiD3t/JahVH
wPd+eUrQrKmQnqApZ7QN1UdUXUrlK8Vpuqu4LcpC5diNVpoEUB2jTboEsLdV1+U1
xdLtP5IvDfu90M5j6fo32IIDaux6qKAzi5v90COIO0WZSFmVBGH1sQm1KOOF4vdj
ULvIDEOgRv1BC5wL6cSGX+n7ZQjOM8HzBdRgFjapgktGyPFIiLjAjix60IDmJrz4
nnznKrBND4dos0Z6S558dQML+8QO1UPLlWa3EZQ6o2zv+jrZxUYMKLHE2GH64el2
Ahl6ycLM3QhQFxv3DZyCfGs0xkaycykVzURkkZd04ksf2Y84q0iXJL+mP8fQUVnP
OaGV7XFJh4S6SJ80rIJQjgtbTfeH6zgfBxnWrotBlfaOGXO/jbpajdPUJYHnZQtN
3UkHOBaa2aNVgO1W2ozQ8eEb486twwdsfaYYFdH8uM3iadswgniJrQsq/4lqzUKU
6sr+arsK8sVr0GlEeSEBbhhyErrGICbo2mRORPFUdyr9iLE3+QcLtMA4XTGkJRc1
weTOv+HRGwOQepKLXzvJBCqxyUNG2P+pAKD9EP0fBCfEAChMWxZojWr/gIxIixL+
IRfB1cOKJAOMQwsSdGv8ZOCfZIhuLykA0xfTG2nDT7xzhpI3dB7CaLHO1W7e1K+8
N8s7tuBQLTQ094ODFGBhwthqp4MwU79A6e7/BPqzh/JO5AYsOvNuTNzI1MrK0uN5
q5jvVGoPeG1fHNvfC6CQ4mWpADviRyY/lxcPzYRYgheXml6icBuvF9suDUF4jDQx
Sy1qG+6H3fACDFmQKp+3eEMKtJFy+E6IFAZE7j3CoMjQu+jppTyKGpsFgswT1sVF
3Ov+L66YXuc82ortEn+gK/gsvJu+XjgNjO1VV5L5sBUP78uU5Q5/QDK4dYSg7A94
Vi3Bqu1pMBJFwTu97uMl7a4/Td12WrCw3mNn16aKNFspeY+7/1jpR2bFvXDOPR4p
K6+pkgQr84Dfgv+SEN0qwQdYcyFW7pAD3JPRHhPOmK6yle3F7exptQ2VdN/aB4h2
fjPsZripK9w8pqTMETiHR7CniyxCi5kQ0+CMdtbLkEL5dC0G69Mmo4WvIaY4QlCl
faUkgwMEKullJk/AO9oJT+qeMRUH5TNZBYwoKWqMKb7Yhb6sdrRKD3hrXA+q/l8w
k8+riZk53t+h9PFLe8tIGuD7uESGYW/1KHJWlc7ViRN4ZlwjoD9ewBCoUKf5rQi2
UUTly87iFKEskAVffKfrggr+B8gMNTRzWWWyGMcLyJWLyAqsURAA3AG4/K36UAlE
5taFqvhZ9AoEU3iiS8jGyf/zLa3ODVKPMS+0jqDtsrn+sSaIpMlgtgwbLfa6fy1t
orgxXAITGkTd/utOHW/sCo4kf2VKsvivs+2Kmou4w3rIxjuffqLTXXm6r+1S5B1C
o1vPUxHtLnMsdNny5PvLuZ6P7AfQ5AGMdu7Ou2Va1NRX1m3r2YNjowe+L8D98m8j
STO6zOjXN26lW61MDVkm2clQ3Xv3w3NeSHOi3QmM0FTsZbazaBNmThMooi0cY6JJ
9mqYH9rekcwHFm7HDraj8LFVtXQ5fGdpSm3OIVNdQqiwQYJaygzFek8N8ZXxA7BZ
9QoFtozea16HfAZbS5NWox0EX9jc45WVRWmrNvw6n083Vw6Cbsws5DMYiD8TlzxK
4flQ9kxII8sLRGVaB/r6tSQvY/5Iyc0m/HejD68JUm6n4uNQNOZuk4Bowx/4N9r/
OOjksT1bHvrzvWeXpJKrUN5SSKh3lihUEIToOiSpDx/Uwm6ECFxdDo1ycAJvCNle
QnUTsQDS5j3X/oOaALtIgIkKg2gCzDhMXE+cSelYGg2RT32Jnkl+OMRy+ugkvzMK
2ufr9Bqfi/yvfwMTW/xjPrSeYJpPGVwvIqH9zwF/7gQ97tCwGbO0BgLNse0djyyB
nLE/dZE99WCE/No7y/0kaiKjQoq1wsejpO2l4Sldj21HqOAkmYBkMdctuc9ql/bR
tnwEIXl50oZCzbtHUileiUC3YICLmdJxJNX7CpVLja9n/YoDTFhiKiz8+fR/yKgh
5qsEZKMYrD9lBZoshJRN4Iv7YvVjH6VRoVnkZ48sowxGutloiJEs4EHsvXgl2Psv
fJDHvU5igxtXCtH3MLdCiP6LS5O0T0DlGZuhOSet3NZNLS2vEJAaMKOPCuv1PFD3
3+Gi+G/+FueCEupHtOjDHAmvJMILq2lruj8GO2kZ8mfF+PkQj+mawH5OOTZZ5ylJ
uAMMKWpTQF679XG9Kr38EPaDdNP5Ou6LD3MLJLjAK+lUahdFRmGL/rKvJv646DX2
HENdGjS/+i4aIacbN3luZwE0f+cCsYo+QZkRhCimaN82TgvTs38fBxufSMusEoXW
b6qqthU8Yt1rcSoAigRYA7tptdn3HhisTcx3m12cC11h/as5d+ZsCkw8SGqguHbA
SqURrcFtvtp06SNTWfMjEy+fZFZSoSa5+22pgCyC2LuHLqjlWDbUFtrkgO3fMXcS
8P5BG0FozpcFpajQJg2yd5MMn6/TEZe2lkRQhzZUGNHBwQ5tsn9IgEdqP6CQGK4t
AX3aK9NH9ose2DqQpFTbPupqp3kT0TuuUlkFfJ5cYANvPO8XqsT/Dpu07qFNbICp
/5sVmALS/4ZA2qx6blsQEA7U6ViadaE3Oflx5YNfNWibRbHtPHrHmMBta1D0kd5w
Rqn/eElX7bQTAoVFA2UGGlTpkXsBdZ4d6ca6TCuaM2CpyTElz9GnpcjKFDmo6b1+
/cB4ucfUyHDt7RnUv2Yff9zhwXk1Uq9aEuXd876JXkAw0risXJD2VS+BB6Gb6Tn7
8phU+X4CcVOxd2D7ur/oWPcr5bcniiOwg0yIk+PRp6MH4HsaxH6ama/3Vt7/1M0I
j+G7jNJjrMfwmhSBl3rNw7Q5fjYDSQ+LjUkqHP9R1Hv4OeQSvyyrOzSUzYYQAI66
4vCemtsRqbV59T1gzgX6Qm2bFgXXCxNeOGokjlLNJkm65rNODzQ3B0etb+bduKl9
gMu8wMn/u0FUQ2uNQGzst1pC3wgZg5mTSKV8k2q0ZBpKNqhNh9qrA5MxgX0liBcH
5vEtj5LfsuDT0bPQiBmEQQxoAdjqIxitf0PHTM5goSiFCgjXLqdCSU0qoELFABFg
JXZLHErVQtcqO40coWZeV4xdy10UkT+Q3tsGsfyuJDUXcNbRvS/0KXl1N5R9YCyC
ujqm7sdiUJcVRRWcoXk06GsTUpDlqLW3/YZeCMAoB0ds/xfnbdrXgea+QW2eBG4M
LsWR6RuuXaHJiat6oL/N54EupJc/vKtmxHKNboZl/FxoddjsszQegklb4hAaqWdR
xAlRWwY7MMavz+QHUCLH2nMVZYcYnWgi5/hq4O6bolYiDMq81vX2Os4OGeI9+Ixg
usA4ndvpvNkQJcJzB9x61vOJi1RXYnfA3TfNwtxz3jtxc/TZ3UC1bFu/GLB3Ahr1
ZXxokFNDaQbdJspWa/kefrMKbJ9KrXtc89D4qoPkD1RTF8+E8sHjaS1tmQ3hQWMV
o6WEPXsDfw+0IdQw1KDV0pMm2kQ2AGpf+hCnuO9vc9tgjHr6MB/gkUfUp0SyRof1
zJQTN6WDMd/ynykxditWnTvFf0kFLmMwclkmUs+6jCtKKJShp/vDKpJgb0XKSVHa
rAYzgWXMStKHhX9wDUzFNSxMYkk1sgA5dhBhh8yZxF26vidkp5Lcpg4yDYzB7xsI
XUO0anD1AM4t6mPkwjfisnu8VRP/hPYTYEmPv1UmMDx+f60HMPsqg0v7dwsWmcjg
6jiR83YX3ljD9FRrYryfsTPhkY8DcT+mnPUTXeBAR4kYbkbrIjTvtXDAejDJbT62
Ugb/ZCd45wAzA+H/z1NOg+aBEgg67tXs5jrjYlPzIqOL4x4v608KFPnhLQQAoON1
qSt4K0rAxFOY2QvkDg8MSSUzGJQwXFKFSDe9/vVhQRegnuncZrVi2BHMxASiLelh
MvluPPqHGkfDon0aWhMjWvxMFDfqq+zHfQ+E0PPX5F2yz8DLQk5oYaakmVFuzWjN
WElAS0JVtoUsXzxIxO6KfJUCmRkFUiwbGYS8vYYWzTFVD4VscposfCGgV4K+j26m
k8s0Lqtq1O9OMQ7uCfR2enW8pvkSdbPztQ3LU9BKgj5Yz2L9b9XybrEdS2lJxmZP
yqabEZtOVLAeMBzy7uAzPKRy1LAIMA54W5lYmx6Xdhn9TT0XoqfXh+ZZ0lMmJYGG
PiS4eT+Ut75HCLQLY0SnDQ7v5NQgDezx9dpnsjklwb3FO83k4s0iwFFrQlJv+sb2
Vno4iHp2l2M2wFmAmVB5tc8HIILeIm1aOpl6sZOFHvi5/wbHIzpbUGMBMwE61jUP
YimVUKsGjepmxXdxXSNHdthq5NTjGhGQ6/SSDAdIwCxUPOo4a/3LMl56Fi7Hp00t
fFEOqe6odn1SMOeWUf3+9abNwTqeqWGNZrPVHlii4/p8f8XjhlW8mgWlbzQc0EsK
DOo5rC2crUg8btZRqzQWxznpV5DRi/pEkyMabauVguDXl0Ldy9jRlLyFd69WyMvi
BeqvpNnO8IxdWqO4j/yUu+fXuMGBQe2nmIW3KO5YqMZHaYMGPeIgosalkf6f7/Dt
v7ncbVArVsc9Hv0JNt9xo50Kwun1oDAfxhXAegBRMUKFFKVuCTydZELZsrT/YeFb
Zs++qgEcqxtT9eKTrZMvK2xqS32AjLvT7h4KSoKJK+PgRJXpLXUGGjYaBegF9x1z
Ck/qg+rGonKPnp48t8ZxRBAQI7JC9OQLJLHVZOwd8kV7Ua2ADkoWIv8+ymytgBiS
MGXi5g/mVrc2LgW6B1CSA0nbfl2NfSB+C4DVwGy8T+qeCbc8C+Bni+WlBewAHuwm
s+xwCpEAeJ6f57Nl9yjv/pzsy6ggHytn5eu5nF7UqYVJt56i2PMU1ad+Cs60VWhH
PKXMcdj/eeqQ3zuELxpUN35Wft3gnWHIDJ6hkKyN8HMwTQ4nGcRJAcEKGuFKc4DU
0Qw8tgLhM/FL4zNRhiSliLz+iKm8RMVcchQT7mRUUec3vEpPAcQ0oCa4AC6Rg4OV
FsFGBzqakC5qyEGLaQUf9Rcj5IuXg7uSDMXgVMCVrrvzj+eGLIZz1QA23ibdQddb
SePBFGOZxBS+OmqiMDywzcEjzPDajIfY4W7Xh4jj+vwh9UgGtuOvCAMPMbAoxDvH
lVmx7bUIfGQMu1zPiIujsLlZ5QM4pAD5b0Y+YHTCjFpQNTVAGBXvycPWuvyLgMYd
H9jfTCBViIlOckY6IHifi8NVqCzNhHb9q1amfVTB3ZC8BjjgdPkFmLcQYuGCnbdU
XFI/pm5P91qCioUNsqCUXBImZ728nNptrCPRiY31D/URMlg2oaBsCqSQDUzv5uNU
V2EQpgfMq0lBPzv0js0hLm1b2jadk0tOhJ2nkM8METsSkpZcln11c1ZhR+zHySrQ
4FgD0NF0PVEx69RSeHuK2IDhh5RVWGzwDTyUKR7+bubDvhdVMbwSeuVF3qVBTvhi
PJiwdDUBiW9Zc19oMO3uHcDNNsuF8tv75cJXF/21cU3p9Z3dQF1xCH3WBajrs1o9
saaKNYctH0wLg9ohRU5iy9jeXg6sw96yPBEpPMMLsyKVG7YDMwyqeFDO2nEKd2pH
dxrC0sl9HoI2HexPGTTDS0VkzSZD1/RK+6Xsg/QilGV89ndg5qCOP3KIoqHKYoSm
pB2LLT8piqOOnuGKeKN485Yp33tzz3NYtYF9dxsp8jstsdm8HCkQT5UeYY/3e192
Z7N7qhxlRwj5lDlG3nexz1JS1kCZL468sbaOJQokSQS1TBteOEAGVcXcU/FqopL6
A2GgJrMskVtcfSB5FW+J+EghlMbrEYslaqLeTtZCdv1BjovWm0kkSZTP1ID+j2Fq
5gvBgdVYaLhYXsnR08bY2lgWAs74O5fvh6cFTmEAOQkGrNjOTfmgIcPCRrEjM2kl
VwBdbml7hoUJRZAP4xhjrEfNOfY4wayDM1W/0mCb831y3F8rOXxoOugarfDjbRQ2
NFeEBd18pyw388KBSEFb2mBU7AUX4jG+IKvonLoyGHrlDlWwgEXLwpKLtmKCXISs
1at/dkbugepClj+BPFTCMzpSDCt/yHk1OB/fcUCGBNU/v+vnG9esD8lMiyveYHZV
l4OcvRQII7WUYow2v+SsQfVtIrAUaURaNdpY764dVOcd4RCl+vAqyFU/fG1y/zrE
pAnUqbqZOkYqLBuFdVGBSlbFpB6OQ+tmPqMJbvPc6yk9zWFxfDYwcqqX+Aoi+xVP
qJKEPq7K6KY9ITrAlspFyZU6H8ry0unx/EuIQ6NTfg6y1/DST4iebdC8C2pVBUgX
23IOxcqYW5zWBzA/mOmSjByUxhhrOKEG9DqY9ZISHbjMIHxsGplkGm/J+Fu1oPit
ZDOpvVfrbO70DM3Vt7H7rVWC96EAANw/8oI6a7FUsgMeBdivwALkjcYCuWjPb1aF
mg5qllbZiEDveBJt8Ao+hjVptmqnBR3X2iP1F+g5QbhNqkCnYUF5HpV5JWFpyilF
SlQtl01kh8CjJeo07DKBsncmxLBGwY+saCMw7T/jbbuUgjQ0vrJwHVJzvV/Qqbtd
Le4KG8m6Nt9362R+Vgv/LU0cPAhYGJlZdxBt00hBWBbyc2sad/7zvOanIojjxGqQ
p0CzfKM1pXBFfv6dt+flghc+WU1B1MAFs8vB6sOKE+X4ydlEE3dyX8uGVRQpP2kj
KKCM0riq8rzJYH9bQ4bF18Pk5UgUN7NGcLaFcou75M5a1fEKd/5iTIbfT4D0y+uY
cmnkLlSUckyBcH1mPT6cOrWBlgY2Hf3OOaZFVWWQmXFLffpeMQzhpQ+29D089RWq
dm64fvn5+tBE54tcUzw+fYGtdlmxSnZkgIZ3kZ+Xgm2S2zPctgdIa3GbKjcZMkG+
ZJkq4ek4nsW6J+2H1qtkS0I7H+aQEQZoNVqyqgnIywt2hvs/mUXfOHxODJI6HB1n
wEV9o47oYzgIwQt/RswkrqBoy8/NiDhRpU+FBBJPOrQyaeH0GVTVbAGtQGaArTDf
2uvlNApaFFC3pXDJRYza4HJW9Q+FPgmHsdRrPLZWFEzBWm4bAUubRfxYCP4ALXf3
k4GFaJ/xvq9JhnQz77jib8Q6I9bzZZFG0IQm5Bsbs3PNjcMnb9DmTsElqofoixDI
EH0cXHvZoc2kGyiyyEAXPm7EhHHvndGCwOnXykWTvPXUQ87DtIALNcFxw1iyQm6O
qv9DwfsOFbax54OSVgc+8GVXBxNW1dwkJzpV1cNEFc0bmXqvwKWWdEkyYi4CJYRq
vmG0yO8bBSfgqf9GHYJmg3qLzPUkqmv4c2+W7Fjl1/XoLva72DgnQyEDMv+iTfKv
4S2SkEyOQomoLttaPmTJFY7r/HM82rV1txWHGZ0AscxeQqoxDns9oSQF6r9csgzg
Xdr8vREy54J9aKpQx/ShRQnGFi4vsH24v4xRKdpIIPjbM8iEccncsvfhD7yR52pk
jPi4t2uqQitPRrD3ruPFnnW3sGSPhS9mSWchY94IiCkg6LU+V3sc5C5MEsNkp9x7
rEdY5bmmg4Zu0v2L1F26HJJbEqxJ/vxX6F8hBEPwjY5O+LZwJk7jS/4dBeaAKksv
2adBiICp17J5RhOoZa/gYV/GlhSnY6bkvGVDojs8en7asGU8C/u/mo237vtEp09A
/liuk35SylmW+a9C1TQL5lOdiscxziL35vD8o1ouKY/PXknN+mhyfJK85mt+POlI
sd1LaRc01WBOMyYCvS8GaR3LhJrpX6b81lErG4EREq4prX696is0P71lmpyutmmP
itlTZWryg9+0xCOweTK+16qnoP1Pq6iqUEfuOu2YBSI47CHu7ubzjclURZW/RXue
WhYyXjYmSzn2QndwdKB0D8fRq+drgdJ7PYyMluGIbrrZ/pSKTMz3Y61qkNhxz58W
MSw3vQFEcRoUlmZuSz0uAnQfBX53/66Y5MaPTs6QLQkR+H5UvFF0Z5Zzs0zrxwHo
yRIKLMUDuKrg0XAn53Mmepf+bYL27LhjThrhV1Te4cziaUL1V5xjiJyNjcLxtUgK
OHXff35NlvrfR/Q8iDyDfCvxlXcze7prdDzy1CfK36LN7kfGtJ7DfHU46rLFsj+V
Nd+1DQDAyUvJzVifAUjXleUMv/12dwHphxrRWmvyhV3q/Lvd8V7apFcpbcAB4jFB
Q6m3iOn5xIkVNzDJBCIckwj02WJuex4IsmRN1rpQtNAbUgnV3DAerbpAfUJrvSiC
tol3IWc521DgqQM/O5Kz581U6XDHL3dXW1JCHBzaVzviAWcw45/HXxdncZr9D7W/
QSn89mn79hOnvERq0EPHSHu1VaHKGcgQforzxzc/0on7GR/ZyyEYpg2qvA02ODmW
wt7/PIVQmF8m1hD6mbIp6JtuZP1OXvQouE0/1iupE+3h+a2/Jt9wzQ+GBwOM6hsC
FMejJAZg0rrNkZQDjYweiE6FWUq2mFSJWKFCx8sh1/l1D7CwDwmw58ncqnlEZADa
7oFhoHgW9wjoLsPwCUQg5dd3PKZVUO6jK5doyqJIMYUTnMRYDKj+/5R+sv7PVTNI
RDj0WuCSr84YNveeazVRypGNFAops0/x2kNxTIOl2xeCUo5kJLiB/YHahJ4tyjuI
/y7NzB3EGZ4ycMXOqb3OPXzAnPxaNNhEWc2N1Bf3ZPwjIwl9BTsu3/lf5trx2+9H
tLfSidM7JkzCSUkdeVhk49GOQO15lgf5tdyxkJ8RVIR0b3Oq6B2zuQqANYnm5xZA
9zAiLIpVmef8LOI5+Mxq65W44BKD0mLnbL7cNe5PxD5oZ6wnpgvSAhsP2unDlTqz
9Oe0dtgHk0Px6Y4gTTfvXpYcaWjR86V0g2KSiyQ0DxgYgE2Go/+ATien0I9iHgNd
8IflC1xSOjo1nY4DXZNSvjsnh9BiJBBEJ8eZL8NjfZ1hUA2GdOyTIzR6d7tiwf4k
YBlurQ2Hxwgao4ukA7yhVxz2plZBDOfKVfN/m1wEaFHWMDtetqnmf8XIA8pMXI1H
zm9Z0ldK5JSu+wpsIpuIxzVCHrerHua3WTEEIdAPB3Fy7PDull2q6g7z/LdL5i/3
M5cFFj5SGT1bY/GR5wZirint5Chfe2fQRtzseNMpcfNHLaeNl7LQkZ9vdBnR5Fn1
/s6KbHGZ3iMNfkDZGMw/NHti+RFSB5JEG11UjzrLCAd7lB1ykhxW+ODFn3mkIzQN
rhruvtO1JOxhtY06mr7rhUkabFLaZGOQIhyAxZg5oY1aClSJbBY1wivLCbQDtW77
dHlQEF4D0OLrX6OoD9begkpfRRMmaMRlDHdEnEdAENBZ+DqkNW3LbUCBll/DHBWw
YC4DHUrIX/fu3hdjgKCzyVlVzze+V40Toj3LzwSh3xJ7XmIOPvCmneVwCJchsh4/
dZ5EZe+Nn8e5jtupmH7wQ1gBqcU88mePgkQ0FtIMFtR9JeBSzVl1CzcXeSoA1pxI
PSR12NTNpj6ijiqXVxBaasLX1F14qIRtybDnYfiIYjm19oB2SWAjvktbXArE5V2M
QjkNuE9S57FQiijEp3krfOCiNXebnIEQnLRaf97o6ZubPE80fzNlnWmSV9GUZoGk
ToxdGioUxByGEIf3SXrGbIyhmIWuyjAlQELHXAFKp89WDInJwk1f4lzpk16yw869
FkshMovKbAbEkKgS/Ke8+DNqV88Wdtg2sL/NFUG9CTR6R0JqIxMPMnaT304sTZ1D
YFcVG1gRnIHOp06MfbaeTcukiOPQehx1yme7YNMpe/8JPD2p/YYhnKtk/glYjjIJ
NiE3kBVl/obdhQtKM+LSXbzx7DcnKsgEV7QfHCIpAobz0Ck2JbmrnE6/m08EE5NV
ShDfOOGWYKI6PMXUWlLdekJEmmCmiR+pH7cRBlvYmw0zckVhSVfimgSpIhBYgYoF
zluur3AzunCi+Dn+min8rhj1HBJHRqFundE+W4eCAc2X4ZI39ptZ0/gy4EiK/4cL
3nhqKeBoMQbFA+hPrKvmvtM+pdM4zsyLykdsjCtzF1AXngPpS/BuTEKv7dmCfYJm
P65YpzehXAqL5g8Agwrsbcf6+U+BDryk28iwlvm2fsoATSJZYEmCxNszDcelfsrG
n7DoHd3JhWqVR+2NNxmRu7saz+HsjSzuwX7x9/JFQQ5B5BY6/NpHM9SZF9dhy+nr
W5xi8Bf59CESZxHu613vs4s/DsxxfVInN6cCTi45fAhjKYv60UQt42j2sdmEreR7
ofbqpFmgLgokKvXLShrV4m83tOJI79aYUM8vLbINHcWxSqr7ezvN+p8bBha72u8g
HCks1oi5RRYaJ6KPvxiGld7riL1AEhfJAdythSzA31NU5/E3q4YM6NE7sjWeTDPZ
MIk9H3B/kVKe4Fayl07rxYD3KgynWRkBVZm9EP3vSZSI6GQ37Som5G1ON4Gq84Zd
uC0SkQz5EDbJM7rN9F2l4V7bsSgjmv3oL14kqEkn8Vqg9nyks/UqHBMwgVF9t1Gs
UoI7httZ8I0JoDx4Vu6/Z53TnPC2eHVvj1Yb4bMugLxhEdNrE9sdRL0iL3JceOrh
FGgjCkYpRK/0w0j3pbHerEPGWHCXJOk5+HLKdIeAmweI21WhdY8YcijTtg1Ja+bp
RXLUQjnz2B1j1P4pnLnzdB/gBCCIetxHC1VZQcxEr0eWmpj4C4+KOcRqR4vLLqLJ
LXxy0+z8WEjKRWM998jFiGkV7DUKN8mBKOICoHIY77P8W1CLC/PZOdWwC4QrHBBQ
2BIe/Hdc9DUzeXrcVBwEK/d6hQ/e3LjRYb9BY6AhDhKwwycpnCS4PQ4uhyxaLCg6
CXaulj05jYnzps8qrc8tdpPOH2GIkYwABCOtNMIdyhNU1W8RhC5DnGSvK4qv33Pt
zg01zb+aMoimsb1csx/jZgJ6aoXPRIPONPr70V1xSJvU4Wp4qPrILL0LSuE/lFvh
2iUu81OX5f5KnquakHV4+/du4I3dO3rQehYEEl7atFe3qA6zYX0ECL2rYUe/lo7M
hqlkhKeD6NS/hzhGfuYTvEI+sv6rFawnqH2hWErSqM1XtwhtO5UnsEkyweOk7J13
sewbWTD4Ivza2q1P9MKAAUCOBmTtcQ3oVKIpjgb8hfI2P+CcQ4BqF2CnUSNy4GRE
LO6o3SHc04bl4rGUbp5HBvR27Php+rvaOvbvQfw4enpXd9cIpMoqveWtcvd0S2vY
7YIfBX88kl9RV6MMuluLqee1kxbNod2znSH3hIbw2JrRcc9vPJv/PzQswOBperkd
FawggxjUzwI2p5lwZfmXdT2bsiwSG1NTz1INwEgFIugNvZa+1gC6XyuS5VhRSuvq
qRIK2/DnjAxPTdBCWlfSSDk/QYWG/wNyk/NFXArL5HHgJh90UQtuOfjKbqvLb92J
spkpbuWntM9eMlw0jxs+2uL0mNSTUldin4qMqfj8JTrPODxbsr8hZwdRURg6Wr2B
kK0ZqcFc6p0CCv0fGodFdZ1xOI9u+J2bbI6jyaoMd2/Lw1EDHhZzVnq4OrvhOwxH
ihc3AoW/5Vs6xbsomUzafVUNtwZInKsDZQQxg2LJikhL2wQMXhqjpI7TYkng6RL+
EeSrSwsJu0LnuOvgq4+bq/6pAfTuWOQ9xUAaH8w5bK3hAj9GhJVL8UqoDR7Ql2DR
ckB/M5AHrKW3u3CYef7dzveQjv2hMjtYAWhRvnBHGEjthPIazslcBkp3kXxA+OU7
ail2DECrsOdkvKRr0FYEi0wmryC883wza82VzRGMsj/jyO4iIYyhGEWHbWZwqT01
x+hqU11rVxR8QFJ/q1uMOOyZeB/luFEWdC/M5jBNleY4aBAA4o8sud8LnjRjgdLu
JAD3bpDEYYrbDNCpMP3ybZ2lYKRJ91Vc7LxBbEtzC7ThbbeuuUSbbLVDMElW6oJx
WeK+yVZJrEbtGyFpo9m43xXRQQ2cYXc1304yoWv46n+W5tPwEYD1/6KNvGNtsXp4
Nk/5EOx5zUHNED/ZM/8bhtJyyCAsgwHI8dBbX0qaUrHLC4vpXBJt7J4mISXP7yM2
oyOLJiJP8K3QhReXpxzou+E0MuCpMClVUUbZshD1D3xckWE6a91/e502zgZHSDMx
mNYtdLyOd+DuMyVx3RW95q+v4Ex23lGYQi6a4VN9Jmse72kPU3npFYomOAptWw48
iWXcOjrfEib96OvGTq5bAGR7ouxE5dGbB92AA4iR6xlUe7ByCyFwpgGb7BQQRJyD
/vW4cC5aX70/30kFMAScAcygb8FVl7xxIGMhx0RnXqXlYwZtnT5OGWnLRAXdJa+A
FIFGUx6881LDIfya6fnUkDSDKBpCmnNoHW0LIzY+1Olyb5fwu3wfkDsuKs6mtfzH
UoAIs3ljsYZORKATjLS/OQ5k10nVgIWRBPi8CD2Y7e1Xr3u+Ch/oVnd1JkDoodGx
tFrpdY2eIFsiWhfLaEXfpEeOjc6DUlkkOkVRiLc4Z+ulLT+uOY0RjqDD51/KePGb
ECHSA0/hPFBLuwXkHCj0pwmKTk8Lpd1WenyczRHD1tzsys4ifQFeYjyFApAY91Nx
HMrNRMJwVEIzfWMVny4yYjzPQz4QiuYHpBZns9LILUaPLqd+wYYtH48qdhizS1UX
YLCYl1mUxriRqQd8rDpgcGj3vY6S05ZDh1X9gus9B2OAhLOzEoKUeEGzoGuXs2cc
65Klp4y5pWG6WvdfBPEsjR7xQRVi6gw/MZJJMtkqhf/JaPAnUsvNHAS7ATfeOQhT
YmM78hHLBhk6Ognz4a5CAbvzYu1jPT3VnJ4fzK8aJDCHnJh3ddC8TYjk/Hn7o50I
KqoQ5+b7F81Qsk3CKmbMF6WK9vaXBdY8iMV9BJE1VVUFh4zvbMoNxG1ikL92r6JY
P1eBXLxMDViWNhAte1cZyZXUWmO53WrNIl77FC/CxQin50DdUzqhHVFhrSubbWOD
7OOP2fdQXi6BEItK6EOSLld+foRDHuipq6laVxW+fXHiHfBRWZRwnGAPFSIMU/dK
bMbcgXf0hyGY1/3qqciYwHMohIbEDAZHbansfMbtM2EGw80Z7GN8N0P2B9n96JDG
DNP8VRs6E70i00PRzxO8o0wsQy1qnmwoHYcraG3Ss14oJev3GdcPnwCmTNKcbqsK
V1HA7NXZMo7Y/aUdPziwNMgYUunyeC6gdw1rw/uJPkic9ry2up3JWxUWErScpQY6
GGnUMjRth0keHFfUTJWpCEFuT6gXmVf00+6QqyeGe195nab50hNS3Z+lQ+f4kbzo
yB5ylTlW3AP2uurstfT4L7E3k2c2d6a+KezWRsmXtx1AETtwjenMv/fgkvmDsIaO
PHg8wp0Lyqnzr6caRhw9QBqRawo0wxUY75Ldfsrfao+C3EKDMryIyZeojRsJxlAT
+TEdV0Y7Q1uJmatvuMcDnXeR7E3I9lD1u91SiEUEr5KAkgRBxpxlnF5haFjW2mzb
Ea1Jw86XdtqkVL8LY81kyE2HpaJQdr9m2TT3x0vZn1ouHSJuZfQZHz5fjWDZImKg
j9nMUOe9ZVrOF0bwTRvvGniLSFCKvJAt/O9NEvabpKC0l6zf33kYLHPNPSCSmHvv
uCkru3xfO49EA+m8sLVuggyqnP3D8L9kklmLIVfaHkrhwdVqgIoN3P9XsPOCULX+
XOWHhC0C3RXaeTURI1GCwo/+4yW4zXjBUR2bgJC/k62Lq/NA9smM9ot1df4wshAB
VC/h3gcf7CrY1gC/fTxN7RsMCVBvcNp34PMR20QEikEvDl7x+vKEN0MT96NFLhLQ
AyfikL4FpQ/iq0JYKSwjCKE16W3tzeixMBLF7tbSXWqKs69u8ITEcOLgHoAosddi
dIf0uR6yB0UaF3vTm+gOldEFObE6KMGAOj55ZMyqTFLUmU0hpQzDFn8MJ1r3ACWR
4fl+co/eSTiUBKdWKotji+XIsCfPHqbA87o9cEukYqygPIqrzMU6Bwwn5k5sJ62J
mop+yQD4dUs/2w4skDOBREyxPz6Dk7O5EYfHw4Ux+ndBeU9RmD6nd6DYLnrDaP58
Nl5jFovmhwwuxHmEqaW8A4VQ1ft42H+GojqLHhvg/xRALCbvtS1ANR+7xeeG5bEy
csKIXQCIhWDXJShFLxZedwzzH32hrS3UDpWN97iL9in71AqThZmSIW41L+i456+5
CVFWZc9+dFAthG6s0hnQVagPC4V3EKinYbW4PSwvFcBG4A1ti4yLgzCkqu6CH5b7
kFpcdRl/M8L9An7fcUd2a74T1bNGCk+V1IDLHn9doudx/FA8qhnv3kq2Zy/RKkeF
NGFWnHWeZIIT/TkjzoFqJWueOR/PbtBIPMdEr0bmzGmgowWsDreoCQ0Q5Sp5hSCI
EVB0Z4pqn5b5SbHvfRCiMtPiF1xq3dqgtsdHzAiO5Wmm3uSlsL8KtancdgAUe2en
kQ90aFGsjRWu1OKb5BF6asT6kUk115dbI3mF/MEjl6IKXjXDXLBoa2V4XZTxgjqS
+B8xJBC0NXnTgKRTLjFNTzrKJSteBcIZk0y39Y9jMQr83YObGct+83CC5QD+SEIi
0aFQR5L8lgIHIQuK8kFqjazIn/2r3SXDGByT5FOXNLtLQZLxJL/piPK4A6eU6I57
X3drDlJn2GwZcdhUIvwrJ0II5Vmg7/cjskFiCroesCU+vtdiSOUzBRaLwkMjpWyo
WV51i2GrAhz8TTrKpYkTEvtD/uH0hXJkItxEY2ZdqvTDt7qtfOY2AERB3ICQUOR1
i04Bv9uHKc17Eo5+8Tcu8qTGcuIwydYkMT6EKORxrY7qIIzUOkAa067JWdXZ6yud
cMY7VURJUy6Z4Kiz7ZiOpyR2mljOdKN2khbo+LhxXLgZNaHA7ragdYpdihJzIgDf
L97uv5WzawOkTZe7jBEpvIfwGY29bxefiwy97EKvIS9nA21m2aLdU4XVtiwKYgND
GAYhbLk9/zzeYAEOz4Amgev6ohnp99GU3a2/Z24pu1iyqP4eWTpNHWIkV/Fx5aNa
F/JUl9zM9B9ffO8goKXMhVaOEsiTUGhHmDxbDSL4HEs7rqctvpWJs+/cV0G2fSOU
lcS0mFOvUl0geNe3LU6nMd+71kQ7P+tofzkYOy4g5jRoENoiAa32je0iHcPfuUog
Gj03SStRKdZ/uVjR5w6cQ87Zhm7752gJBpmQOUsZ5Waun9rVf1Apbr67Fj8NmGl/
deQcwj0iNP0/6dv+jxiDEKZGOb6NrZi3xMEIY7KixPBP4mpDwP0N2bZOpnLecl7F
DCpQBSl/uLYa+VILOa01B7+yD0kZ1lNOujdu9CKo3qSN/RTKCYiSai7BXu1GF9XD
vri8yl4SbYACd0hgbowFTSgWtE1n9VeoHO1XPPPrFUOu2XP1l0Xt7GxOPILT9kun
7vHbCEz6Ndap0G10vpQJs193KVyqe219s7WtmGfUv8dQUBPPBWoUkAcgP6SFnicW
Gk3zbfvcIvrTF8c/mtdmmrMb9VmZ3j19kr9+fxgvBuAIt0yHCiQ7fQgiEIUEeOt+
sTzR6zAnbF49T6hohgzxfzKSp4/7P0sfJ5D+yrGZpUYk6JldLMF9rr30w0hdxdSz
nnvGI19OIjXhYYHfX+hFUXf8LP9XSyaDy/SXz/VrJfZD9A0NADlYeXVFpl0K/Dag
K9hN2Jv5mVMu6AST4+hqaMS2V878Ap3u33508utK27+Vw4jPvKQZmSaM8zd/SINx
1r/JCzXk85C3aRn2sJYxVw0NH8QUwN3OdmH0Qx7ptJ4bq8uS9bMfeZpeBhhkLq3w
Z9us9DCJwh520OUaH6x/lccK7mxpsZtVprSSkS8tDLFHxINft9Is9pilv+0/j23P
5qOUR4Iv9xz0lEgFbufW+6ij1qKolmifC2mmqq9BZNaqFlDIrXmYC048MQftQxjP
IR9R9KxqRdVCIaJ4bPxZ/w7KAW6NYUwDF7dCeJdMRUCZYgjkAXhvD/ggSfN90aC/
4ZO3ic7y9NczymMtgv+hRV97mfWpKp9Wa0lP2S6rvPAksZ0S20kbKvURCbm03lo1
UaeAOKy0aZcQVGr/jxYbsXf5La30IINphdnjtqjJ2EgAesvpxGu51R8Oeg/0Llb4
1D61Zi/0vV39b2FOe4jgNBJd8X3HGn7l89dyMC2+75DJHefIIEq438TovozECLlY
L0cE2bE6iezxWzYvHaA/r85m35RdJ6F3YMQ6yIIQvpqKZ5m8XBv+VzAFFThll3kD
v06ZI4P+9/ibtKgaPCI0QoWtI/XBkDqdpg9TzIFJlqzTG8sCWvBCEcJq73LdRoSv
vAp+pNBsx5dXJoPjfFSz7oiYg4zPYZxzTw+2dS/022dwLS3wKpp4xiFx3NEHQL+R
7gpgQXTLwd4/RJhxbdhjIuOkTZA3mVg3Z+3EbQQZBB9djcydHFSZtLChPhAwbQmU
21qqzNjGLewznuuL9f3oooTrB+gLESEB6KrPPmpy4DJbOxXZsH+vLdY9salKVDbc
wbyb771PgWTl+k7zmHpcIHJE6sFn62cgxAHbg5A0y440rx/dGj+31XJkVFK8MdIu
gVXmHV3UYheZLxmAbDgHNMS4sxBSuuzo/1f+KM89GwMTtEEdSAXMIUS3InEhtxoJ
Jv0M15aFRrC5OXuU+/8la/tnOpYcLr/StGZYkohECgHqPq6/7OC+0J4VNySeoPZt
V+vq1kZG188spwWaDdQwD1pTggRKzb7IVPknVkT/3XquUY3X+SduVX1uTSD4r3eu
NlwhPJykkRp7LyZ8dGULIcw22xcNZCs/fWWCgmkOriN4nUdsI0LZwAeg2MmOqbtm
EOlz4Fu0xwQd94LhEC8HVvzv2WrRTELo7EVMtKZcKMdzO2DKBC8CJsPsVKl5GdQN
28j1QF/kgcFbXGUSCgWjJLxaaGhW1XJhn5jW5FBXex0F73apL9iJLuhe3QQ1T/dB
NfhcDy3aWdTmxK81jTvzXsnVcMSt1okWnI2hddrarUThgDUfns4guMkmp6IRKv4U
Md+vZmXWeiyvpvuomGIuQLArwMl9l6i7mXSs681gW3X1h30BKm979btoSHsB4+Dv
xhV/+KbTJxMLTV8+OnuS1TDzx3kZLQM1hOlCIYn2IKSg16CEN1RHj1oDbgYCBQ1k
zc4OoRABMcro23HUzhjaWff4AkB1xR8ZzjWiJU/dej5psui3Iwu2aDJVj1BWVDhG
QMX5XGfn7HyGga4v5BKxcKBNem+SDkwrYw8KgfsP+j3vBEu/bYMC28Q2OdM3h+1M
LI12PS+cVkF/jXPiihm6BIGcpwp1kOJ8Gvk8nlHdZEm4Wml3R3H/OUDgV5B01/gx
212GW9eHFwhWaxtQHXB450I1vrNXnflu6EiN2NYLOkdQ0z2T+Myic9/8rmZugoRV
ntRGsZxgddNWM3p5fGBWRC3uf2NO47lKIAY6lhmAnomytjoberDv28ULs1qNhO4s
sHO0G7s1ONolo+z9vi3wUQWVmGBcSfgUw0uA1DPDxaoHowCzEr/fZFpW20RLMOiv
A0AoHJlj68gP5t/sDLYC4VfTp1n+yph58x0GgCoqcIvRSDT9xWGZhifnvN8RFxg2
PcBoJTkFtTQPQxG8J5WxMvl90DTPJUi0baNAVcijh6Xt3XhLiHOEKBPwEfKgBUmL
zExyRz0ciURql7ZIacqRN9BlpTImroKoYGzNYd+7b+ooAHcguvjCBQKWBu41cHDF
AMif5fGYdhfVZ272nEf9wrFi3qs8jqphUPvTTLWpsnpAntPbpCV3DZmsr/fNdAnc
VJ5Jk5aJ3N4/4ASqX163geieyBb25fyI71j0farTGb2PwBJbRlMEdNgy//hkKBdk
mpZg/+I76do0nLP/QPYjy3N/0904/Nmo9A2HYDoN0cvJ+sRIvkya5mbM463+bsDa
B0fMeZ/FlP4jWXAp3e1uG2iBzynOrHVK3kPOXg/aXiCUbEb5E/2Zd1gaOtBT9fhf
2zOI4uEGVT1OYHuhBKoforNxWoCXQVHTbfPQw9oJWgAwhW/S3YHrsQeMukwJVgbP
2jC7AVftagg6MRWse0aKWYqvdQoXhys3TcLZAv+MsGUy68A6WkHRQRSFIbd5jqy7
h3g1ZlrKVaaCkR/8AB4CKOL6OpwtCwuo0iAr3T94cYt2+7TrRdtZqvH5NgCu+Lo5
lpg15YVmdwx2QKtn+kEJLrAmE7TP+BQimfRenJLXR+Rt9/BSUhcyxdaweRHiRwK7
1oc54b0e6GR/jzpTphVAsq+IZQ7J46Ud8SsXJcVuqy8Me4ruKY+tjTYup/0/TGPi
nOX8J1zVJbUJE676CnUbwucIN0X/UmHJtabhb6Qf0qcAhINzyiDG/GPZDsnu2C+c
0snzj0kAW/6hrMitI015RikhupWs4DntXLhVIB5FdkPZIZzqa+4z39Euk+qsKIvo
EGJWSJb6xNWXX7KAAoOxUeTl7cyE3LwjpBCKAgw+VCagQMx4mpPE56WXLdKh5Zce
6rGeXikRpHWSvjy+Q8nm1OQKMaJOmXGcvZw/aewc7qmKyBMobzkVc2L+mBFBvasx
WyRSBSY5LXI1xUBizWmRq1kYmHTxFhrDE4IrMxgeocNM8i7/cybpsk77zenKNHRu
dxYH1E+ZjpaaDOULIbEe/eRVG5l5n88XEybSP1H11gdKBUfWVKNahtiOn2VJS7zW
Ib4VdElW5cx65w1CNRHedxGGL/W6BUFE7GrIxcFwUte/2c4ibLg+U2Np2/50Ttn3
L3tYU/+F3anIPg+YgjTYz2r3bA2JwG4n5DYsQLc1VZ5VI+58mQSfiZxOusXR6+N1
zKD/Kmjm4PSB5QVhd3Ged9QF8k1c2xeInZgl1UlHp118ICtUYRPppyjOBVVKnIvb
0f+8kjvHmK+zXYWUHwuNgC6/viLO6+yo9XB3Ff0UmfQKmnAmvDdixX9XJUwkHj9P
7MmuB4ZatzqFaOgmR9WbyFpJILHOCbP5h8ndxgQIwqKC3JjZ9/oqvvssvCGK67ig
jW7xLMkcCXKtE+30Cl+gbLMNTt65WPyHTTFvAvKd8lid8BagR1hqOzCyH0b8q6UU
Zxzi107ajO77Lg+tZWrUrmN95YQa5OAKpuedZp2Dvg2NtBW2f4aSewy6zr+IZ/Up
ZOrXiqjojIxsBxrh+wpZgVIsK4JYHaynzp4MCjqpbtFRYcVQHvs7cdRzJuIxJ3ua
4KX4tTBwthSeAQ9pDM14T7CAxJPl8U94z9kNLpKWRrQrLZfQj39JTdxFTdcvyxMb
wHHVMHt3nHAijp42WL9CSUcDo79fuVO7eLt9D61P2hYUbf7EaxKbgPCegIEoVTIE
5RUUWdcOObNOjAbh4VuNoH9H0DcZFeKxfRfNWBfPtVsXAjG1GkJ2ZcaExEtVL7yC
B0adJiaGBcAgmLH4m30IKszFlTi8jUaAdcnPrkZVVIiMt7YYDwFEX0CLSr0AB7RL
wW0wPJvW12mMo36gpWnZmZp+r5y5sjvh/ct3HsSC7JWC6sHCJo64/tB3DEAbdmZp
rbSl4u1Zktlnmj6ffJ80jo0RLXEzwUH7S67UGKl2IKFY6hA9MSk2PyA5ufD3TQCk
ZHfK4bvNu79OpD5kbh/LIT0ff78x13SxdFnn9BgLkrBYcWj8bkjRhGTRNFH4Diw7
E/BQ4r2NXLq9BEQ5B4XGgiS4IUcRFBrJYtZCzSLgD0BZ9uS48z96m/Eas/Dt6CKL
H7QwlDvbX/ve0D0qwc3w3B3RhQnRF/AwmMYYVj0nQMp4F9TPHxrvPJq0Q0ynkmN4
XGc+Sq8UD0WCiSL+cd1LSkNl/P+MK4CE/A6oBwCIHPUdx07FeEHO94zJXqWnH3On
CA3tw4vuP85kHqZOZImO8HZqE7JgMJZHl2CccnzgLWFFWC8QBk5Ko6vJfIdl1Ex7
LDr0K4ztwFvLCrLZJU2H0IrwnJcEDAuvXHp3NpW0i2deZ7Y4yi+dCQ2XQofa3EeM
isg8zYnnQqpXQV9YwZd0lRL+v0gKvdOGin94ycIMYMJZDBfX1+c0uVrOcAFRhVlB
jpk58DBCsHjmZY5UN9K8IpUMvN4XCnB+fIt1KOrsQJVhi1EVTzu4Zl7DsNL9ndZ4
tJI3YY1GRYoB4AR5A6oBbG9ycGw2Im41/OnW6zHtsQp5WP8trlDbYow4k7EW7uJg
7SIOoYFOsAuZfmXq8I9Ap1GRpBWlP1hnE+vvjylAADocNv7WvF0v1Rt3XtYsLDhA
yGf3pKS/3+N3MNhLBr9NVEWmd28zniTnXrqHDSgHV4lNvREEFIMDybWxc88Zwmoc
pc3tlhihN25nVRMcL6KiFq4ctL+f7+NFwwRRP7gdFihKH9H1F2Nqn8MFzlUxaqbR
M9T3K6VwD1ZiL6+OD6MlD1ijrwty4mKSJBMcnjbWG3ixPOB5n30+axerfWz6of5g
hXfpjcXeZ+cwZeYZxu8xtxIuKuxpYOVdcztIXhsp/WHWjKkHG+brRw2tfX+cg8/b
3GjG3D39KUR7woVzyRlcE0egaesCHGTloNWIpzBBPCu+L5QLdTIn6/w4mNKPoiAg
w+IpRnkKWfUA5yVDNQ6+6WvC/nJ52fphAdMqnI5+4PAo2d5NG3UUNYbZQ5MjtbiF
qNh59uFCy4KMDDUU9bZYqMU9fwmGKbcrTh2UDieChrOIpd0TNXXnZs4V0tUM5kra
dL1s+mGZ3j+FsFmJ0LbagA4T5Y6g/Wt+pBkcJo7l89UcTVvy5FwOMfukz0q87K50
x3E/dSbX8xELv2fD5vKSDxG8cqDYf5t86bTV3ZZvCWIyq13DhFPyCnwdzMlC9pCy
yBXgZA3gfbNDS4cTci0ozZELXCuksMMB2FJFHb544kw16yPV4/tROsjXsKR4Rv65
AdqEUXDdEYc5oE9df52qofH+bR3q75Ppl6XKBhgiUnDttIg9btdfkxAA/h8xc1L9
I+8Cumjo005n3SIcVL0O8uYbfz0H+jB17e4O94NQhxnWoVbfW9HizVjQVGnNXEYx
CS0LdzEfKASueowa9Bh524XRc8nN9OPEc+L3CzlP+rUoAjeI43UQbvguLtpQbRc5
8srziVSpRNdzJPha8tmynPl77mu0EndqnD/G+/KugDKUW6TG6jfdWpAIVMb3uI+p
+rkJ6ZL2iSKRlPYSH3iN2r8Ni/PT9kZVxI+OWAjuKBe2YEPQGZaKD7jWHeEyzJfo
cPEN2Zr8qRgwOZWHp46SDbw/6J89rlrYokEjfKDNEZr2+03GeZZWPzvKrnvNDZFh
TW5TigN80qtXtTVS+LXOkYLPThJf8KjW8NsR2MG3LdFsE8Iub4QDScsZqG7CWOYC
eiCLI+Rfc8SOFReWDLlM6gPW6hbtMCdtnKUP1MgEmNLGtL+RW76p+N2UF+EtWlUT
VRPgPx30VGHkSA++dOPbHA7HNV2tZGHhwxLscYK8r47ztK/fwybx3m7xb0G7cNsP
H4DDcMXAPcqnh550abz6OvNvGe4F/2JCtD94uM3hc7R4SP/mN3HJkmco7I8w6zg1
NdsIe42bDzV7zQIx2l6U5USWBQwCVekX1gX51pI5yI6mn6lHTSdPJKvip5Won8qW
c/mbDqYAq/kDnj7F0hhOnM5DwgLaZwHqIc/yY2jjSjVJ6pntYtyvA0u0twpmyaIv
xU4uyaanGbyZE8w5yfGNk76obVoFLFXVfoq9VU1Q5YdJQKNNtczQKTEyF8Z27F7P
HHaDytue9Pmf8A4Wskcu5HShgjGIH4Jzfomy+as94x0nvmQDdCy6FrhTB1oFF75B
E33jIbPvnHVSjK+IHLCxIT8JuvIqS7clC/bsW4Gr8ArsF+ZLUThdl3ha0OPpyYb+
BUvF7Gl5qhXSJwBNK3z7zw9zIt1DtKZQl32IdcB/mnu58TSVcXCjC4FaXTvSY9TF
kwLRw9s7dNJLsIyf39do60rhR9FB8fSZDfHjuJ6+lzbbs/byt4JWXEy6IbYBqYvi
PiSN+f4aD80L4uCQiQbmSdHa8MBwBsB8uqafIxnCn4GzK21HyszCpjp1l9ftJIE6
6cM1dNAqotXflXl8yoLLUAecov7r7O2auPlVK4o/raGqwqhXedt1+goL3/PxW+YA
vCgT9UDT71b1n0LBG/qnuvth2zky+yfxTgzyCeroJQndyCeg4cbsJvKuGZKefH3v
Q1XoVVbpssv8seaFXqJVmxwXI3eH7aJP1LdKbxXiRTpsf/fUzfRMDR1qVmgVK5FA
5azAWeY1AbelXU32XBTCQl0kbDJIVs8oghr0IN5UGluTZDu2oY3aPVX3ju0Vn1Jf
CVI6baT6TfCSIv3zzXinvYZMiHfmkqQqW1inJz+C/5YAnUPhsyJawd3j9Crfs0GP
0yQE/Bw2NXG0mkh0Osa4hpwKMEn+7hbz7bly6t+I+A/8IZhtBAWvw8cA+mUMZCPI
gAdu5eul7kAQfb9pGTougyKK/b2Q9IiK2dxFNYA4cv82wl0AVnunvVIihq6N5ht3
DoIFMC6M/UTssLEkclMqU/SbRjeOpTz6lDGKz53S90p7Fv0uxycUabkEalpUz+7J
BuO8MVY1jNwabNsMKXwdnWCK2qzwqtnBSpbit4Ip5Hj8yOn6FnftwOOu+64jCujM
bRPQjYu9BWYrdCbHqM5tF4wrB+ukasClpWh8UFkeNbsKVRoHZCU7RhbhtZE6Slrt
faqSngxhcvnw8PWoVY7PZ61or7+pT9fUPzka9v9g/7C9TUcxzKqhDsLfv8Kc2oOr
nLBR7orPyb7rgLuOlPFiingfnMGxOvBoNXcBwJFp1WbRdxNhT0hx760f0gwoD6yc
K78A8pFs8Z6vdeqPR4EI4yrBKBThbdBKnbCQ6sikPPOAmccRJ44mVjYmbIvnV20E
ccQf7nhUNsJuP5beOKOwoRw8N5qqO2VlqU5yMXpMRowhZfZKkvHh0Peh8WmOGA1/
tyvsgfGl0KWJLFlj8XqEA4KcFsAY8TUT3rpXcuQn4YdwsD1qjmBimiM88J9IXDTw
2D30ufZLQVrJkmt3p1LDT4jqAvMjq+wXSKeDQYyWnohxwDI6OuKeVptUfybkJt+g
8NuDrOq/etFzBASir/nFkifh3bAplYpS5/H+rD0Nk/03eJ2oCUpm+XpDqPZVIucM
zoROKk5VyIlOKZX4yYK4O7Z4rqBOHREZAk1By/x3f5SPZCuEVEkDCaO9TCiZyPe3
6MFcoe6a0uw8ATxtc/GUiSUvhYeTF6fznz5dDkV62pBH482kG/qknp6d8bcDi+fJ
g5e2wJObbx3FmKFE0gTwocU8G2atmcIkw1V8XPbTa7RgA/fGXafuhKd9wEog4Rh1
hKSapWbPsxfF25wZO3RvTHDf0pfOS6GYHiclJnuIVTIJhewRDGSde/YaIEvfKlNc
NA2rvnsr2ZAlX0HQuH0LSAt7lOnb5w3TVtQqRm8IIlIQOqi4jH2yjJ1oqfe6oTbh
FwJsFCzFDRvPTWvORfmpkgLguxx58SxrWxJ4CZ5qDL953sCZ+7R3lO59FRY8+hl1
JsCfk6aN6saVRqwRWf0CPJ4e72K2lUOIHIvbKnApXwBReHhFwV9MBSdae9xF06KT
RgxQ7urJxg8Rv3jndnbBmJWJozUe4g3vtTBF2NKBs43dGkJ5E675t7fiKaJWs+Q2
coarQnGIxZITgWVHG0AGprExPDUPML4AVrdpnNEm8rhQG0UOTOfJAwUycpoWCfzV
AfCOTB6gRPMVvTDm1Fgjal/MbfhNF4OeXupaD6kUhfjTtgGbMp9/m251Y6CNIfen
2VkdRi2ce6ezSycnc0eEVTZ9vKz2ZnxKNf2+hOofuKW4Jfx+iP9lTgzRJXFn05cR
5dcPAHQDFzUVHVS+clSmBJixOqOGnNDvoVQH6dJON4f5YjB3GnivOJlLkUfVhdm8
/ZphiMiyI4cYkj+InTDtxmbQewUEKeAU3++cfsx0b7iyP1p+5Wk1wnFTMAnneHcl
EbRilgU8KwyvMJM8nVI1xVmA1v/6DJqOVggPuuAk2/C+9jC3vvEVW1OtQyHSaScW
NHo8Z89HDYD13wN919nWBo0Whhz/ausC64zo3TrTcjmdTbVYIOwekfOCSBILqUR6
xpN5RCPsCdaHRcR2G0/jh1JM1yN/KJF06b8cvcaX9tB/yrd1yO8jX8Koc6MAvogv
lZ/d3gamVWvNzB0Wo/9AwDlOXc2lnifITQf9tg/SFQt81MkNHmwRgTNTnpIjJ6RL
2xvC+HJoT0KlxoqyCmXPO5q+8TUwZXslC3S8Y+WokpnBxcIlYUFtEqmy0qqUtGuC
Jjoa+gMMbdeSkjW5L5WdKKewNU8/kr5SktnkjT1gSImLpi+h8pRPYKvXneZfR6+j
qIaNM0v8hBgnrQ1ksYH3fzHs/FL4MZK1Oo06roIoTwILxMqR6hK5hwJ3iCp8rops
VBlMQ8vqbJzjhI1JP60DLjiswwpFVFWnhLLTovquHwPT7ANSmpN1Y91jzvt8zyKv
OgRrz+FMoqUl7c5+Tyr7JwBYP2etEjwLHJImbRhi3TlCfdX0ffqiIHiE3GbVPUKI
ZlTjF+hfkHi6tAlN7tCPzVfCbsbMhktaIcbO6RmNYFO31XhBsYuW0a8ziP9uoPYs
+bt8zhECwYZKfhjN72n72NguZC4SNWjn1+V4q4sJZOrrOo1ohH8kAEcZvb7o0PSJ
MctzRlaibKMPIVyc2Fm0Wmfmd/CUgX+fsqkfBdu424ErP3H4kMGhzDk/qidvEu8J
/tstqBtYHTnAl9n5Zkhu+VOkQUIYYd/j8Sk+o2VzA3onRHasHZS2C066yBp1gO38
VQUfALf6qv62xk+EsO2n4rm2sh+E6DroYqjLBz8QMIIdusLw1uh5DQG61mHMDLCB
LZeu1oXl11AE2LVMCCr5qY+1ZlpyllwNvxVoryfqebe5A7qQotYZfXV7oIQXw+F7
ceHtclC+gwLrbGpEUI3syLSF3uIaqkFugwj/6lmlIEp8u+i1BbsDvkfW/HcYLw4d
kovdD/6pgsnoEbeh2VMo0YRCSpDT/M3Vc92F9PXF/SsgxjJfEFdPUYxUvIaHk4l0
GBNIc3ERljOmGS3bXNUxTZGa0cLZ/y8iiLAxuVhwedqEIm2cYZ8aGw5yK7fUDpBE
86WEobR+XSUqFpZn85CvRyTSdsZ96zf7/LHUde5xqudajoIPmAla2Q23URClm0Em
41cX9o4BiwogzbGphWGuq2rid53FsCOiGmitF/dH7r8aF7aLhA+wUs8TfFpxWTX+
/e3dXUecIoVENXFmW7jmO8sWsy9aOl9ibQeKScdUzigJUyrO7/2W67fSrFm48wDD
6rXG6NUZAWjiyWKoE2mniCco5CT8Q+tzD8XJCm7T/cTddZiD3DfkR/6ZmQ4ohN+u
Q/OqfjIW9JCp0D1BJ9GT799faZDDup4JRlfFjZL4YB5zvt3CRF5FAHBCfBtCwbzI
pk+Kfi38LmXkhUAZTgf9uICkjdVQ3F4ifq5kQyz8o3YTqQuZcg1VLiaahus1g45q
c0J6ntzjGzPJAUptbBnqTO7y4jiG90eGV0P9S9SkBmmYeULuRZWc62kISV4T18nG
8Hg6Rt+7kwT5kH3DXaT8SDyKYyAyweOTZLXTd1ahBC+2bxlHsI/LVXQLiTDSpfDk
1WiX4NnWDTSuXAj8dKvTpWxbola8mNOEHbw9fpjUPFPPeaBIS9k3TReS80Xxdz+e
Tp1CjZ7til86l9tefO/7niK5gsxICydhSHroOqVKFYlmPiWB+q2UJwp1/L8SSTQk
yUr/xqoFnw7D8yd4JZIFt0b3ZIlKgf6mRw34Yad3Zu9YwgG34wDXtHCt8+7dXiZe
hQEzNXd3Yb0pG5gywONxid1O2v8TrWKANy+htWl4b3SdVjPYU/qhSaCgb8051kuJ
63sma3lwHKFd5H9ecnqhEgOHwTx3+k+GUWNfY2WS3BfcGQLflU/z22ijeWvw7ihi
Jq+F6t/Fe6orrwWSmx3SrA83aNhaNt48+KCMFK64ZODKfSjznELonJUn74kvpg6H
wh2evS9xXiWIRCJ+9fkd8wibLsIKW3o0Wtnm56pPFtdEmvG0vh2+xDEV4CMZadJz
bM1CsdhrLuvfLiXPnzQDUboOe9uKXyXS9wup+lAr3wYwsiR0It/K0ebBzQzn88C2
kxyOBb9GC1UPjJXUk0zfDS4tsuOk3eZjH6Rd2SeuqqQZMbnhnvxeYc9ejafmCZgQ
RJjy+7AePA3zSPqwZOZOl0fTMDJajHB0zIpSVis+5QrlDE3Vzd7Mtq+inupViikf
1xnewYrFfYeHkI6mR5T9ICZ1C0vOy7EFR1DhxVcUtHzpkXGYpI5IDZFlYyQSr1uc
wur0EU/Ahn/+z1bxP7THLPMFpni1Lncq+4S9YpZsedCXbZwmtUIVgllqrrSkGp9m
PJQK+Flu0GWAkl0Sz13IpAPBSF1gARoeNJm8y7q24CKCFysMJqBr17rEhIknKNUN
PYi/uG3pvC0r4lA1+W08wVc5Gdo7butTRvLmV4kqCSSVww9lhEd//Q1wkBGgGRFe
k/6QKM/NiRFrwrCZHbMlCscRUh4+2cFjCxFZRH0ZZKNIOCz8WCa5kNlCoXU22I4e
H/8SmE5ejaP/grh1CcXpn+SEEyL7JD/5F7KBFLJiwscBr8Dc1GxY7RXttPa7Eidw
6WuFc019r1jTmzxVMZO8qZZh/oFPzydCN6OPWJVNU5h36UQ0VJda+OJ7lkVn6dna
9vgYC8ZhcxAgt0I4CgywBkES/MjTxUcMQdjddPJDNH+8mxZC5/qdIHOov/WEZtKW
p6p11Jy0aPVvWc2JK0smkF5XYgQtPrT7R+qt7zUYrMx8DEfG+TY0jrhV8THGE1Qg
w6tNhBk2R4I2VNxyMQAEgZXIEK3BL/CgGDpjHtsdniDepkUw6VzUAgCYuVc7Tpn5
4arEDFlKx8Jbb2Kk/QP2DAs2CmoDVSdqkZmX6HImVKwYnF129sL+Y9c5KBxyYgGx
xCMciWwNkBdAEmWvFdqrtICI9BhhEN99eqr7UjTxLm1teiPPUscTqiNWtoQNGqQs
EYSweBw2HxiLCwn44O8XRhyNX47kG5Euv+rygKWW/o6d87j9EsUcwKoBpG5wLpjO
juhphAkZODd3oAIvBUT0DWOoD/RqRH4C1mxoKRJNybJNW0MOt+T9t+Hw0wBGn/lb
kPfrK7x4wjV3ZQhI567y+iJm0zi11lI444JghAu5azu2CeDUZfGnts9kuO79i/XP
5jPccL4nuQ1m/ecD35ABiOjnE4kxfyuLzPT3P3yGG3jKk0rkrZYPzF40PzOHU0ph
RVuVRQFrxSC1rPD+Be79W6GmFYJP+xjI7RxHw4VS3bSjIR3UZwZ35h/MwWUYBJRc
ur6opTW4mjWkJVSstFKK4xWYnOcxE4WezsMU7XKoo/EenHLVnwyuqQv1pKrigHb2
M9PJNq3SyUuCqPhf1Hc74m6+/2dEQ4RmLTbqWws/anhsk+0DdktojH5eah4yOmPp
mzKqLsRIZCBoNEBA052+aErSfVv3Rt9/jjJXSiPZNh08txqZsbB5mEU9P49RryI+
tXX0OVo/m6fL6+4qQrTwNO+2tOzJDhHPHNrTYlHLcm4G5Bx5+ZaO99A4++ZLPV2/
DGj6ELNgvAw4nxfl7FNcy1HMAXUYpeuyVh584TgwGbUynHzrTqjJuB6M9UM+GFcf
yJ5oN66/K6uE7z9wqFKWt088Jgusub73rqIGCXCCl77qEluHfGEOixTxwSe0c0SH
7fc3AcnoIoa/V0/is7FeXrKUY4d4cALk5p4okNpkr9gU4ChZwL8v4PyZqUszNuj1
yubhMNZJ3fTF/ZjLAooSkd4cfe7Z626UzwUqg+70G8y76dBN/yLJn30JHxCkplUw
G20BiimEcv52TWnN4Qeq5Wl+pOXM1pZlzNRSAeizRLLUeQz0XLIOskwsWpOT5lUr
hg9kHRjq90ppAAS65g4F1/HeGU08mP8VRT0hneDhcjfCOdY4gIZL0SPF+U5Mxb/c
EFu6bPchq2g95oGgXkoNXR69ENrUy0V64V7ipTJM6DuH5qqUbYA5/uuGBhhbKH1E
QaK4lY3oiUfwETumSgkoF18CAYMmTTXwNMxSJib56yvnglwrKPCQf36dv6NCUPsz
t4q1sdV+UHU/ac0Y6i5WVwFJFCBM/23ngwdUqcXU4YeLr92qk1ctoXyHAZrVKth/
qCAKo5VoRc6cdRPNhwVKaFJLEFD0yjvCdS5Gi1jcd5BMUU/uWNaaZp6GHZgVvVlp
w1xYhP/V02j2S0E2k9C+z11j9PQpUuD+9Yd4trAhDIXtRWrRNrkDeCflTnZ+Ki1m
vcV/rVaKHAzAUEFySvfvCqgNGlgnxewvidcl/b5TCW3tYTSDD4m8yJTzBW/3NMpU
NMu52WXLsWA8P2hG+3T9xi3LWosyT17ccTjw4zvj9HWy4DuAIch/eo4C8RoJEJtY
TCvmLZLn65W5hKvAyPhzMqGSOzYz5Hm5M1OditZ+zfHWYKMly8/18F4nJIdv0woe
vGhT0EuWs3IFW+cdtGIXW4VFYokomXg+GPQcnKoFDDEHlbzFJXffMuu8SdN6sBZc
8puVmaNdUHUd/aM3Omhx889AUmg5LjCLQDqYu1DqB411OCJEt0d8GgIORsJtZa9X
dSMg48qqFY452lHfhnWvbfpUixO0+k/K9P3Axp7ZfePAuvKM8WfYQ8jXLZrx3Ri1
ZlZTah6h4RfLgv2lYMvHJAqmXhSq4alYGWDTrTpdiuOOqQCuai/EFdj5OE57fYOL
qSiGKSvP4YoBW7PbTl3IsuvoQqYIaEZgk2rkR9EIYnfNiqHhWE1+eo/iLqz6ZljA
b/Q/59HeNkwfGebqQDzdruwKvc4iVc/Zf7BCqCr3rp+VvFbaOadC7zyXyDSm5djY
ucl4m1quzKEql+JM++nueo62DlyqwXXOJxn+NI0ZPCI1IR7nryboPVjVdA+Tlevg
yWsM1Ix2V2lzDnxwqraD+iycCEHVkcPZBao5fGoE4BMq+zENvpTer2MY20bJ4ieV
sZXF/lp4lhYRA1ooqwvx1jCJSzDZ8VQZJUDwXm20luCFEswONVoTj0qT69CkEnFk
NOmZzw7UpmxJUZ5w8gz+9MH2mhs5A9B8U3qnqSK1+NU4bRj5EDsQ0bHcVHv3IH+k
K4KVvkm5c+ew/csZ44WE28WMn6oP08wvznZ7gpXY4VcXbQOnNZehaHqrbSj9bETg
2xDIjHCfgUSG9yw04Ii3gFpmJHjKlkxK2kLKtVIUOkOUnVLWlKQ4jnbUi2hGSenx
sxHYIaybdfoFStVBjE12PbApk/o/obO8nb9LW/mFa8tzEJ6wc0XYCwgLeo6zKIlB
FzYevs6nY6L4JwFKCJoyr2hZwt767XJNAA4x95hkR5hIL5VD4C3Pzzpv+rcY3OLs
HUDVYCjQCz1GMyv9SHGgpsG/WGs1TvJldThQhDZnphLfJLYZzSw/y3CtfnJjwkiy
Px3QMxYYefC7xZ40HvUsP7KHoGZw0x5nlrCiL/YuMeCcHM5+ylXGp/7rgoax7vCk
c0HmNCI0smg3WTdJbg563BKoMSl6GgGCaDYCi11yDaNiWUcakX4CMWUM0bBZAOF4
HWM5hgdmKDnwjrZWjIrvfqQBkXNfHOD0XZ5weRqF6odvwnxsmhh+OdvOATeNbKO5
hwrqwJA4CfvJyq0I+b7BG4XaKRA61JylUY0xZu78YlJWWYVDoNgXDay+/CJf4XMw
Zk+2Ex1mcmx/b90/XCgkNOsdMc+xisaPk3a9+JIvCpOm/SV6Gpac8CsQPN6rqh7s
i28elpb7Els2be6ay4qdMoWkhrHRPa/oU5ePA/60xOMjzoPMSQYtllHrhyYNv2P+
NNVaqzS6N9MruVtv7PqQ/zxPSturO9X+nYHl2+mHl99X4Klyp/93JLIpptCmSSZ0
v+xOHWEZafvA98oe/FKHUNglO3Fd7RQmINLG06CqyNsmwx/inhXMvT0VMJT7Lqpd
0zOJ/4CTLDNfMCRQ+raB1EfwjKaCspcqQEuAxKgjrh0+0VkuOpwm84ONcLvtJd4B
N8bgBYC1W996dUhAOXs9FvNgb/GPcRdicE+dIuUW15C5t+G2ze1WlhnPNFMZ0zos
b0cHzuwlH7zkGJ1QR5FrGwwTVS1U1VsEUMAYaAmwfDrMHKQbaRzpJav1EehdnB/s
N7R4LYUKlDw3GrRmTXGvZndqvBmzDuXeCtW8H1qSAoi7xslrOfTTtEdMH78SPnCB
+FiEIHTDIa287OCZj18/sF0CLuIRXapMuxZsaggSXkcOByfZgIL4qhYyK7YqNikA
VYfHDo1shRyeFcvtgSzxnASSw90NWFb5siBmgnrHxcRvImsxHU1Y54bH1Wqvj0FL
Hw7grHuuoUparjsGGtW/L27DCbPojSjFDLwpTcG67Eg79h6BeoPdodY1gAtMfEmp
cWnYh69iUjz6/B/cnTfRYtmaHLZ885uSeUIUdeazJBVsLZssRdYcWQNMq73A1mY6
3MinRw2jNPqQWK5u4aU020ZWPNvUo0ijWchIdjcJbOhIb8R4+KZOUPtHE/7L0ps3
eUk3AKyGf+nTXt5YElxFwFxLpyJJM2ZrxGwTHQNwrK/aL6YXphfS2TwP/5ccOa94
+1aNTx/TIJm2mDO3t5awyZk51iHaD5eMSK3gCxyzsipqJcytHJDMIpgfaR+9cW9E
BtdOrFD2fLF3gKn9O/5mJYMKSILHe4pTENEtRcfMCXZtgQ4f8GAqKNMsH33s/AhS
XHjkDYWf+EGTiAedwtlqlGojRPE7sIxurFaGAQjNQtxQOJiE6EfOrLiAbNpF4Q9k
Coletsdcdc4rjW+r4tGE204tzNxF480h6apNaRyTu/jfL7yFl48GCBPmFXzzlLjD
0Ap5fa62AFDQYr7oAzs0Cn/FCB871oE067wvKvjapUoGdrd2sELosJMlgphbAa2q
ww2KhF6b8rRyvPqeCF4nb0XHP15oQ9SNXo14V4fmv6j4RmmW7lFe8j7wb9+dTE7v
WWNxFcMcVAFrzCoDVrF+vtHguW9ghNz25D0XPQ4g1nljmTN1BoGttLFStAcJ9N/j
50Nhf4Chku6UWWdg3kO1VIz41a9JG3k6XNj1senGgW3yKfc6kG0aNy+4qhQ3gPuA
Tf0HjLPiofehZ+fr9TqY4vlYescnsxB893Q8HsQDKzdBiiq8Wqj4T3adbn1oOnnv
vEofA4XgtxvBtwiabP53DngVfcM2Nf7eRecX0GruUCcFippsKhw36bRQRWG/qsZn
6bgCElhAJwzSxnqh09dHgcEKg09n+5D2a2etjH/HUGwS3/Efds3foXUyQwOQAgQF
F8DpukKJwBA/ob5/dIpwGuS2yAryskllnJijGWMg+pCepTzUt5/PYq6rkmRIdusZ
Rv4HCaGsQevwIzHiwaRIuMLQaUkW9CZGwj1/rZJY+W+pdhnfAcK3BoeMmcdBqw8E
Wy+BU57V5zOUvIJNbjGoO26nWgCQbvIkK9WDA9JdUmkCZCa57ub9tDQSPRLg1VzS
u4F+nA0Y/SM2d7Mk2gPtiyppQZ2DaM/Rqw1wq0x5IvXPWrUDa+CmrnfWuCrr7p8J
LN6qK1XQ/GtPugxWQjbql5VfPDUr+f7JslXvJTZuOgARDkMPIbAXzKLPXx+2j/tK
xyahQ2YlNdAIAVspginFa4IA8hPavMz/YkKlJ3vlpNmrXsSPtdSsM4n7ncyxBVED
025tieDqlwpeRcXutkXNKb1IchQvhYS49Z0SdwT8axZdTcnJEf69t7Tm/VeP33Gl
hXss3jZ4UTvdeKZu/Ey2zX0QlaiiGVBSkkUHJVBaxPatB1vMhTn8CTWE9cepAPaz
Qkn1OfCEXQ9WBWnWUeRu514umUNZIVZO7LlAFDBhZCkQcuf+0SsLWZ/vztiXAHEO
lUlbKIJ00M4OJZxf1sO0D54ukt1W6aX3jxl32oZs0qEfd/f8YmROZbXLC9pK18i6
T6G2u4/ox3Z3wu/j/Ro0ho8gAOSrNYjDrTEDlbxj6hAQE4flPqSvuBvfXJlNzZb9
smO/tTckrp0+uipwJ/7vU4RB/AYg/N4iIs8rY3JrQ4u/tACSFs+b5vVXPswZkue5
JXOV4lCMtvVrpbO8+4CH/Hbd8DX7A9WkWDiSO3r67pIuoIkUamoQMOVapV1NHmVB
GPm+9WBjWtDQEBjXOSpjteP3bxesLqdWpRTLpiZKMLkKy9KquUXjG4MoEeQ8+qox
hWXI9Xj4pTUzqUJODd0HpIANIzHXng7LTyDvm9ivkpfAhojxCq7apcgovMT+9uZf
a4+YbUCSrch8JKdqt1VQgJFMGysSOC/tIK3434YqoJB0VawlBzj4Kky2B9OqBNDe
x9NlSCrtVRDf5Q+x3GgNKEbIIimNDF0Ov3HS6fAwWc2rtWZYPq1oQhZEO9QF1+6r
bEe9UqVO/RZXPAGZ6Xg1ta4KfqlwTcin9QtyL0ge0lNoZhMl9Ok575UT7Zzmga5e
Q7SIriszYBlotEsTZWJyEUcTKBv3e+GDE8PTyJB/c5Ah5aJAC4C+fIglHD5VCThV
wQN9AFL3CCsN9REV6D6LIFBg3cPU9yJTYqp29biFXRXO6OXHydtjEaE2iJUKBeeg
fYjJNgu719rdJq/4PfjxQPDgsZ/UFiDLoDgn1CZ2DPHRFwGJEYRW/VIbjsqlxdc0
EPU3JNbk3zfWtnxQi64gfziCNSJksKpUafG4O7tN6efzYqIiUFypNOTOUH1MdJGv
LzwBXzYuTvDRB45Avs1JRBUdkQcTMIa+ABQBSOCW6F2J0sm8ErGiWC82n0sH/kE1
vyyVFRzEAx0oUpQ473OK8H1ATz+LaNzUry5o95pJl5JiwYoFwLIGXItrz8a4/UwS
dVy1wqiNagOE3xWZtcjdI522OgFOSOeFnY/ew/J5Ekh8wRrsZ5B+/0AKoQWXF5Qx
Wl0mz83gcd2X5bUBkUSRfIR0bsWS/VpHwB8r0KWhBDr60wUfwpONl09SmN9+UKrt
s1oglJtvjO4VuwNieliwWFJG4Mz7IPghhgvu6NYVm5IXPwv6iGljN7sXsOHvoe+X
bat8jkYgYcD/heuP813syLGhJcgtm4MZvEI2Chsuhirhr5AxSncQHvBlLnqotuMi
1FzPLTI4sYSk7f1DDk3+Blx6n41OAByNEwdeJq3ASaiAdSyoTXvMUo+vXrTBkjj1
0x0lmfjIxXYllYFM4fV0Crvsy4jJ8OZLCyTYyr+ZZ9T37Yo8svga+S+U8q7wIVCB
nxS7eA1C0YlVLCHUQjQMfi7UkTQqWRkmcwfnJzudAqZCuFqA6pb6JR5uCHhf6KFj
fggcefogI+wsSGQIX0DLDMlODN1L9mLS9ba1/bYlM9jXUBRy51zKSKt4Aj5Pc5z+
OYIYFWowP03+HwKeni7BiSEhoIiK1i8SxvIyN/F9gTaGY9PNhj2ZOU85xseYT26P
Z6CcjPsM2+X0tr1gCIH4kbyIroE96ycbpfZeXfR0CbBmJQseit55VjygqHNK4UWX
USJ8pbyNgv6EfgmS4BWctqNa4f4Qd1ck+oKmhjzPIKFo/5FaCWm9CrTNQSZcCmRj
xHAWfUWqyrd/eIUXr8DT2cdXf2UmJYCud1NurJjUmeTV9z7sA9nMLtC6RSvFoAwK
rMXf840e97ZaJM3QzrLvt9tzILZL08x/2fwgQ1SZLE1xXJ5pr2cQWIn0B69W++KD
Y+/vT77KzUYE9qiIr8dNSIlQu4/l/dyOWMQy/PSIxE6UbRD/J/SkBAthphY1NuOB
qA+AYpPcl1Ru3qGvlcU1loyds5wZg8BSSTaxJ1KJg6fWT5rMszW7gIkijIabjZKW
eBPI76IARrMusjm0Iv9J3qCikwnSE5lspJIyyeCSWB+LxtlbvZZWZR5DZ+W8EesT
9CbFOUocYBpMdx0+hyix9EvXq3bdQpitHK5EL50eecv/cw/ntAsnqGU5Z45j8th4
uFpfPwLFMqzItteAbRQt2XhKV9maH+oQoJQmN56Mk9cTOJ8yeJRjT9nbnQSUUM0x
xN0Z0J7wbOy4Dq+QKaFd3IygPu/od2ZH8ICB2picUQ4Dz6nr33C4or3aefl03B0l
GQ5mwpUc6rj9dBX0T3uGS0WsDAjaBmiBe8HJudLbFK+6BeVTxxws7oW8O1Njk3Ba
o1SFl3Fy6p2qP0vCTyVezPnibmJ8HPVlxFtqQf70Mcs0YxPnwT7D4Kt/Jx0HJI94
Dv9Y7NHCd45fTBHOzwa9QlWDDc4JtxMtn2vZiVyeybiKlcvi0squv2mAXwViHTRR
tXH2Y1QzWJLv/bUZHE3spiy9JBsGI0cOBWsg4odqk2/sMuaqYiVmRw1VXhM7YxCN
8mBC5Lml0SkVVp9y6WjGTbiX00LA2WfMOMoTgR9AvvloYewu7Xf/0EaSJ48nL366
GE+9y8+PX3UgZzvZSYC4//5fsZesNJ0F/3vt/uORRLVy7CHszJuL+FI1oRc0MPV3
9V8IkQJOw0y5FcvSsBPCllFtbtABIrZSBwLvvZPqD2f1V1IGdd4cJ8n6vTSYKIex
v7c6jOII8HY/RHMOuIdbdB5VtUheiZqcRutlujV2dlGt0agNkCpO4m8BCtKU8zGL
9cp1cjRPXyOMSYKg5N5ZDHf9eofJXzrXBkgWuokPalHxfKORnYU7X3aJ2Rc9Hczx
Sbwg8h5AjGREQbwY7WagTdolwBYKZ1QRVcdsoJCSbUED6falxXprAtBBrdZtHjmq
H72Zu0lssSextF+sh+Jn+j3fCQbEszafDDW4KOuZP7rSVm2P/mb/kx8Jr2svw0kW
w2lLMwyF9QGhIY3kDn4lJiX9+4Fv7wnM9ZiCrfA/BVMiMVC0wPzfJRNTUUNZ8sk6
kf4wK0NY0vGf8QLIUq8wZ1VGKEucpvBZzRaD1e3NYvUa/Hhh85bUzJ+17Muf0pLG
CAYhUcb2zhaKWHdiePCSRaqCTPcMcBH7eybLB+uUFBuoJHnthGFSewSF5uT6T2of
sKS37pUHlwZsq33X6VEsovsKOqQb4Ol0rHQ6mjQ+bYrEYZpKOPP4IYlGYyKt6051
ccNJihZCmoEkHYjd2rpxDro2qMgQkNzPdqKJXNArJ2B+Fu70ssafi6teARxwx3mz
zu2+ijSNtLS0lawbTvxf8/3pHSPz47wlv7NYYZGB2LIuvCSeXcMory1hUln/+G/g
FYllQnlIRb66s714/Yrzv/nNuP7vHy8qbWlUoz9z07unSxqoSw5WLb83Zc5/wpyJ
9lT0ZY+2HRr2yVfbsvBSaqGHi8PO9MuDwRcIlcN66Z8KBt+o9E853ntgoeoEKvVg
63k65w2yrOaPoEfOnNpg2hM3TkJ9SwN6ijCcCZ/nAGaC53q8pEzgbG2QY3spAd+j
El/hhfvQ8ypmuhz+Nn/2O+HPGv5G1Ry4/l3gEoUiDYVX8WY25VJdYEt5G7mOfIZr
HzSwpb2w13KW593yhmMHVx+IB4r6RVC71u96mN0y5EGQjqo1fp6TR6+IjqvBQku7
8YmpO6FymcVHwbmhdQ0N/UhP48Gl1A9Iim0CZqn6ow5pj9Gdp3SiGGGVj4rkM/7b
yn9EXICZQiqJSDBXDB8nj1sov+10ikTzg7R4nqyHqtBAmhuLEGdwi/ZaHVl1nHDp
ezAbJcdYz9NbeZobXzBLpvHC6DmeGKaX55zC4C8QcqwvXGT9aYvTUR4CZEobCU51
RTB/31XVJMUEeM+UhkDbqYUNiSctY6Q1iuVFV9ZDL5iddNuYG634qjkrJAL/nxPa
SSOE0dpZVHFQNeycLi0+/zwflRUm8jdnOlWY+B9E9rBrBY1Me/4ysUwSOXo02UdE
NqwifCnqpBVNRXGRhZki38tNyicor9ibT5ORxBfbJvRsL+9oWLWXds6hVmRHu/p/
WfjUhdkM+sHctl+vvc4WLSspmAV3Iy7pjgLCc+2GMedVI9QyYfXZdgW/w5GyLYV+
F3dojXtgfxNxxOqfzIPRRussJVdTlDzPVSRVAlAM7sps9byQkz5MB2P74rppqC4r
Tg+UCbKw0R8Fha557DHbjYNdBxBzWMcOGMyS39wlCwGM6aVKTivVJlLSePC5Wi7m
Xxp4HrRGDrXDXAN03+B209oJuzqbHdZGxXYNGHY5fLTqImLki5Xp8SF2hMY4D9O0
iFEv3BlIunuN0UgUftDD1SK1bXDnd5NgQYKI0u4+GWbLcoT2NqzIEyMestbjYsRb
GJn2PdF67Ss/47U6XIbLUrSmn7yloUJYDT897kllCs/RtHaGCou9SmBnU823ChF6
zJM+cWvD8sfyg3gWInurD+rhWKVGOhx5IVruCDFUGqzXVBA8qUPziWwXGDNZykp/
GDKkTJC8sFFX/Ce3dLo+5VKuMjX/NkfdAOO5BtzvTuqKYT9XVcHF9ybg518zOQaQ
4XbAY7XlytlqaOrT0zkt7YhIQ7YfzH4DtkGT5SXo/74k95OG1oO2aBgn33YJkSCw
1xLk5DzlUoz5fTBXBR9xcoxkrISU3vjUBP05bQIq8gHQBzDyYaxyFizkYcwrAFG1
p6OOPMioPVSaObzKv03Y/TA1FPs+xIZRKLRZfxTAXHI15tknkzTPx9blNCvuUWiz
liABsBxcaPtA73aIYMsfVmdWoZNjzPp5hnK0WNzPnbhzRatjq10wk1wuhsI6xYB4
LSraWjAEAaXcmko/77GF+4zzAnmZbixZziCbGwuSqwJ+6G8+PWo/SRVp9iEnz4WG
4iEqBFd0NtK1RttNGgp8HzxvKal6smDaFkvHt1qSm4r6stSRF+dWT17nnqzTqWuf
24BqN+5jHMzVTYEJ2i8TZsL++PvGU2hIwQcm4oRUmlSjSDuiwtp/1mgEjYF8f0Ea
kZWZ+rUCevFq6yzwVVRzvQtYquugyW0Ppamds1r+vtlZ3/avqSgTpn62QUhuHi5N
jnHEBcxwUlqU7TukX4bZkr09jVecxaiKtlhLVo9El0hKsOTIl+npfM66gvX2vogy
09maW0O2fqjAV8bkK/fKF6+wjqBZ5J7YAG/Yv9yAQIByHYwebgiGhJGSEEkhKoit
WE6EwRBVgZJk6eDPMBO6FuKYXPIkO4ZKLNKQRHiDCYRbSDg6WIlgpFu+/aiZKcM+
uzL8S8ZvLwKcbGDidDGrTjRe3pvrpP0H50lJIAdtKQX7pft9Gmewkd+2SizGtZxE
NgWDyr9ZeBre5OM1Hf4oCOKa3r3wizof9gn2OYsLUtde3o4oBey6S+t04Krj/Ays
ubjepvWz9bzkPpRiUV5l8Q++WzzCVbskULaumxH6BZERJcaQeyJwLZiQeT18Mmqk
Iw7t73innHLcZqkxjoa22K9YSXbgzhri7UYVC9JNkG1cy1xj2sY5ZSyIJnOpFLXL
BFh2kuqIsG82d36hahB9ul96qxL2za+rexfRoyW8tuwHV0hLSRIT+DSpoQVsesEN
Az12r0Dsg099TMCUtGNXKNTtToRoisGsuPAjLA3lnCHFqUEPeNSDPpIokCQ8Y5kM
SxgKQVCCXME+XvA4UURngzDfCxLsf16XTnrljRKbn+a4SOJWSXZcift7EBIVqab+
0HG21ON1pxyFXxEmt78TkENrfDmb7ynwfN76DVIgZPDH3TNMoNNWl3sIk+XJOk6J
UfsbAzLDthv/yog5DdS+pUn8vtreKwrAM7togPLpqOY6Z+9wonmNkmtTXghS4nL0
jjEE8ukF4mn/fhY3/480RlLgbOgNaiLsegTlV3oMnCgO8M63kzTiBJL2HGJBrgkO
S4BLboySWUkb8nk3fGkP37X962VDqVOghYTZWwmhw+CNiYtRvJRsz/DxYOeaOJLN
4GbovkHzhDW3hgZyFDCAil66wHpt7h9x+elGjZFzHM0W5LdaP2pyWCGlLuf+mp2E
9Cbu3nqlj8NX6wLHf0sx1R8V2OQsqdnhAy+Z3mHGAIYRWZGTj2HOLzr5N/8nBDIV
Ua2w6WWCa1/2j7TgK6X9xzmmkq2UvPbt/NPCSkyZCUo8COuGGKjjpSd+iOiSH1cL
Oxg8PLwi4IoHXEIGKk5f5Q0A/6Ui/UuPLex0fS40sMTWpn44iVjE3xZZQ/76W88K
IIlLyoYGL/43dbI8C8TG7YJPucQeXfa6KAEYqby6RJmWkxLoQIgRqruewkBjI2tf
R5IhlERAklo/iMCzCL8Klk7Gv+oBVLc8UKYePDIG/53U7QOkZ2mBrKMbhwfriU9b
nxX2a/FdmGY2+Z/UeO/Yfu6T89e6kjoTRxhiR5jsY+tG+qhrZNEPv6Au13pwnCZx
EdPJJMXG7ChaFZi+D5NK1MKE8G/emym+4/ynkScpZTfiQxpbGjYq52jjmX6dJl77
4lReJakPl1OkbeJLd/oEdyuP97iC4gStJLOHeb61L4qBrUhTH3UXZ+sms9+6MwWG
CGnJ1ms41T49RMge2Y/5IQPpKGfSixCVmjQMQjZIvBWKWm+3+dGHpAU1QNTs8h4K
FE6/TnMnQ1KHzWjrBmY0w7ej0zD3kup4ym7kK1Q+rGEfQuAPF2mDiuPyTykrlvzW
VSGBmEc/c5Z5sByqlAg7Rpnn+lhu+R7wUTTnJ5c1k0xdF+8z1461BLne+jHBq4lK
dKMhkK7ixVgV4rUoBzDSSxQsxWgt0rRQTwhSkYexVLSa9wg+ttR2rn6BIht2amOb
wQj1J1D9MwGtNB5+udlPZpemKO2l8dk4SLIYdfpn0luo0s4GZ68GLEpS2fR/QXIO
dPXcobxpVVnJs/OJf4Z5whlCcdnoNn/KxPS2wLnyL95p3ixzwCFBpo2Hibf53h9V
CKz/6v9S+c3N6oMpYldCmQ4BdGQ6ZzrJoeLc+0tNeyHvsy5Rp6DU2e+bUUVxupb9
bjV4il1bJb5gPQiIW0gbugMUCDFwXpti0LRTyTpWh5FZnCPPSF0EC58vjv8Yfs6H
RJ1mHWKTDVSOh+95zfE9aeQxWWlalHPWPw6L+yCMKvU8tee0apAffWBpnbi7Nl8h
EVFCP/WSwmHO8kTYaDHrudj2kZ/6qcxzZAfmOqg1e5S8NNxl4AZetF2cvM4ZvRVY
Vju1ZeoKTVmWYtSisNNRRyg/AM4XzYtI6jn6EU0H2lk6NurWcpy+ndV2r/1+YJ3c
n/+Hc5qvz+g+DHOYiKJAnfjmaBexezWgsufuRYhjBVQWApBypocmd7UwcfLZDyBA
MDFp0mgqaEkPT5U0wTKyU+DtWY4GtWvV14ECSqFzSCWVWHCUFgSIgNFHiEuPsCcV
pwHFjoNjhq74GKoxzQpNlZ13eZJk9O8Yj3llIasQj2CBUbVyx60SI/NwhkW9ELqq
NREhEm5EebX0XCnFBdg4X0LO0lwhklxZUeNLSsITebOKdjpmAdGqmwzgs24j9e8x
okcd8WwUQeRjRnqyG6yBEWhHAGPiUPWtu8h4WYxrXv9Ollot4fiJW3e2CLIwicth
415MYibtoKM45dgE1JNONueoadDghtp9Fx31x4LVr8UlF5vFSg46yFcJ0KKRtnxn
TX9a998IP7Xg/Yo3upJKMJ+vRs4UEn18/TZS4uArv9wj3wU5VoW8jXAgwa/W+xhl
/WCdv2tFZ+qD1V39BXuazb3LHGqPonu19yWY8Ia2ex4EUKWDXUlVamD5ueS4j+oc
U6N3vxW6GinvZm33fiskvMZJ5/yRII5Kgvq63IDc7yumOz1HHE7J34ixE0VDi+QI
dm74x138IWDn3XaZ5ajvJnehqgMAw3acgPMYR7zkfB10CCogzlCSOGEetkIBDu2o
lo/4GnZWFPNaxoeFs1+a6hd6HYPuqzXgkix19qMobTtpR2yM+QgQUt6PvDjqR3jy
plFyGp4VkF6vcGErVLFjgMMerwLZB8CmthrR2pkxJ+aaKlzzoYJeUQjdmHigRbL9
RVYABzZNhBOkymkddQkMAL/jPiWkLMVLYm4b4b+kwuNoudTFtLeUzQ+vJ4D2aQuT
5igbV9aH+S/0F8H6z442Z0OmWE6HTM5ZykHnmWNRMpiP6nI3LFapUOUk3WH4QFih
yCmx0b1+jQS2z2YR0psoB2m6oSBQm2AY+2AuyTaN4AStK6JJ+Cv5D7b/sM2S8tnx
5aiFI5DbYnF0zwHtAlXUIIJHkAqKnZ7NSx2Eup52VqPJWjH2K0jiwUCX/cerb94T
pJrfj4yeudtg9p+F5SaJKRY/DI52iiR4/uP3Cn1+HZVF8KTkO49LuTqavxOHIQTN
cGZPjEssLglQLnCsA6lTcxvNW3/w3Val1q827R0tVKirbtMg6oxxbpDyOC6mHhbq
zQaZAzwFaI6t1g4Zi61/d1c4HZoR7PF07KEC8O2+RrNE5YGWL0L57Iz0kyuMUlaA
2GIKYSGl7vpJrUny2tt9QzkWUNtMGPuWo/CKaByI+m7XUn2p7iTNzyvp+2KEBCCC
2GrNMGCY/LSoPWtaQ6xhfXnHpK00Cn65LeWZi5nhBTeiv+/R6bTjD/srpAgwC7jq
EBBD0PrPnQ6us1G2+qdG5vHX7xWqnd5wuGsNCFwbYVNGvoVY8NasvttndTrPBMQj
fSjkvrjDDY7z4vuxzcoopD6nA8Rfs/EFb9IUsK490HuKCNNGW77/PU/nDlomDjHj
CaqY04yVQ9G3xgKprduaFTg7UDx97hSr1AWVWYO9Kpxtnfbj151j7k/R48aqSBJo
nmoKzMm2ksKocrDAZ2uQVhciXC+41u/D4F4JeGmsgJ0Al2yu1g9yUkTd8ZtPdMxP
ZdxD5LZwN4Ya1gcNlQpmCfHJFv03shPsLBx4t+WKbpqVR2OdSUIMsIeymTn2iKmO
CMSdX4S86tm8DpNsFtdpTX92gdXKrj6P31U8MvuFfRLuybfukVGLUA7fdhjEqK3W
DO1/7jg7aVuYYxT3bIORpAU32N8BPhKVohOErci+7K/C+K3lqxWsQNESQir61ohS
UyMJpyFlOX7YtBQaaWREUqVr237Arq324fWAcC9EqJN59Jeh5va2EHMlQO9g7KEA
IL8fSK/cEhT6UAWkhqc9JwpmjUnEW5ll3+i5Rgbns0kM13C+UpIvr94N98PO7zMW
qWJP3R9BUHG2oBdhLt3Wdne5ct0cDW42k0lNFkEj32LssKWlDE+8AMc9ZbWo+I2t
8U9HWXWY9jbPUSHalqw8f6z4aeeLDoiRWwojRxOBNHRvpW4xc/0B+qkMILPoXuYP
Jg24yp7BviGJHVuSYXXqPRKhqSVnRM2Krhr8TVmuDGzHtCOJRmKuN+ZAyP/mNMqi
+D1/rgYEzZKJPVxCxu3FkXwBabOX4pr8WRFbntp0krWG0t5KG3+lStudwh21kbCA
srfsw6UAPS6emeo413TuNcohendBhs5HakNg6HkTTgfPcFHES/R0s05mtbhjRWTj
+4ec92/X5UJ7J7Cvc0Qg2KGZvbj7mx2kfOlEZXhEqw6aTGRtzE9N7Kfr4jiTumWO
K9+J83p/xtevNFgpqKr4/OJCdttGZwIAUWQptlNosT93Mm1y1Cm3QVjsk4Tpme6J
vfF5vUyfz8c+mg5GYysJgkb9ZhNhF/r/0caj5znmGaCWjilgolJUfI5rSHU20mrz
6lPqP6qDusrfW7tlsKYVJ3aahV19bl77OsU247VKubFPZ72ccd4E44w/UaBf3ljh
x83bgK2XA3flDvMyZPG3f7p2SiAnmW9TqxNpOWq9hdw+tkYSlEEbl1r/jbwXGsvs
1mpoTFsZWYRpSReF7SxahUQluSktgX5BJzcbVYh1RDahXE8z4zNW30NjcyBts2SP
LMFH+/T+67H3LyJ4Fm9xvJl6bWy5Y94Td3yD1mmFu2dD6OO08Tvb2v4WAOplX1vU
1yBEKNsNSg8UYac9ucifp85VHrh4YodUdNQ5DOgDxpYl8FS7iQ8FWuF05m6Iz1wG
6ijz3v3fO2K4tzIS3Uat7DZAifIoE8FGS1jmIoWGxqMSk/QgJWkvqYa0gfhkDYtz
g6we7C/Vw8qEW1+0dw7kyLLAkXSjbyCeOwZrx86Y7rtGNgdTucSmsPpTHuYne5Mc
hzIDkp5pr8sRWdpSROWyZE1hRJ1X1w0F1m5FyWoGQ7CzHDSDFTZcwAM+8o0bM2Fw
Cazz57hbXqe5U1NBfHvGs6WNbQqIThSVS2h62nzDiYJdxlZ/j8hmvcwJhpb1aB+U
tA5hJ1zS0rL9/6yNqftZPviNcdU0GJ8I9P3gHSl3KU2K8CGviSsVdxH0I5VYRXLx
JPJERbNCeb+hPQ7XdKt9yfeW7X27X/tSWENmqprxt5i8nl8un1uYHApCZ7ozgn+Z
zja6y1n4iBfcJGU5mx0WHsgDTsBglUJ+Acgk6qs2AMQ5Kzy1MKcKcSpc7U3vG8yg
0xk9RJvSqSkPXH7od7c30l5v8R9RnVXo4mLvUmJ0d90i6miPBr6SSlr0lJDwVlPV
9HETO93ynn4xcPjlLRiHF+PAS7JiYX66ZZs/qU9wOVmleb3DN0ucsACUYuNbZjxr
dWrZPl7GuTCMsabFXi2n2REakvaEnawGgpUMDA3ER/bb3iNDJfBqpCOiSyCr+KJr
wp1yXOv5sDqk68xdiGUgFpdno11cyZLhu9KG7U4C1VnlnLfLE/TqCLdg6m7W+Fu7
NbdpadvdzGskQyzDXBEEuc3CDY8XbEwLWraRGAerfQY+ZXRYAZ4IrlyrF2VbLhco
c57kZINglSafE6jX4JeCnrhaf8IV41mGLXQLPrNiq3szqjieZEf2ynyFU8dU6V78
+voNIRHa2eoJow6kbEHjwDmZ1OMqp/GtNT3xC5piSJGlwizF1ocGIjrRa1797NvT
nM9yiyrf6C9luVx+AvdSF+wU7e3OvdS96tRW6ITKyaOIOOAKKe7s4RPpknNX2GVd
UeNf6wrQfl/PbNtWURgtKg7tPZ2XoPVFAxZh4YHjcTUgbEahyei7fKC9kq3htXyX
TaqbGAlIFJ8osWFTmX9X4kKRl4UmvjoWxh0e/y6z4OWbQ8cR4PJpi5s+B4Egud9g
j3C764BulVYm7re0ZOJ47MlsXdQFYzYrr6tD/FauwYThCLYv7UQwyq6KrhKqFtwR
EXKHRKGmJDSPGhgaaq8GgU3uurmZackdsTRX7QjWxSKGap2EIiWN57ENyW5nQFp4
OmD66M7jm7IAcgWLmw+C6jLZS+BB7JS+ClWwt3eqtvtfj28f9GdIfPSpHjuTQp5M
5ndVJzrLD9Wac1VFo6W3lD08XT02jF3BxGqbF2otnEVZ62Vvph9ON05eQfyF+e4j
dxCed+FclMy37qpYLN35Nn1RcIwdqEXaW8rKcsOYf8PxWEHgVZJCePvlBvox3MKc
SeLxTY5NQXkTxbi2lASbYOUq8zW3oqjGzqzB6VzS1gL3scX32pltmAYbLd2TE0Q5
rmN4YoNTTg1LNhKxSUzKWLSeYn3rng6o6fSM4M1Xs4Zr7NkrjXh+KoikM0Xp63Ja
6v7IuFLVrmmCJyqiD5JG8nNXKK1dEvBAnczY4sjGquDQSLVpMwOgIZzZPqsVbEYr
cKSfQ4hoAP5oIlaOd5bA6QzJHkqwA77iBy7CA7vOzrIhi/4VxEHznp4eEXHKukNd
CybrysO/kZIaJwDS3c1jxHtWyKz7ybA3D3EsZSTro3cWva8yJBEq352DQCk6eNhf
D+tnff9egI5qGgiM7cZdQUvoKmH2ANKviXSGB4BPvoD9byeQNUXe6a6R0Wc7Ucdk
EUrtU2d8bokMTHVXsbroWcpHs54+MI8Pf19JeeOGtGdBa+L3jMxHTBLygVrYC49p
p8yFIBkptc4chNcNliGKjBlo/8yY8Uq8rDfa9oDFcaX02GYAzh5tGVuwmKI2aH4+
cI4td3RRX18cylvAroDVNI1tNCunwJJ4nwz/yKFWB5ZWD6Wie1lJ3rEuUEXjrj8o
XH4bQzyuhC6vz94Yer4/Q4Gq7MHebdiDM3ORwHItHiKKuSJoYjjKhWhKXHOnNeMU
dKO9GyKsCveULLaJM1pzvrDR4iU1+4+zOa2Af0QrcIIV2ReVz8CKu9O3o2/ttHmA
PbEaVLRgfcIpfSFUGsmu5QXeJbffvVC9yaQtTKjHIdjf5FguqkdekK/voy5QgQr/
M+bIk2KIOQ01SAQ4jajD+kzqmcsx/hGO5wTBjk+QdWl0xpAmYbLg0/Q8LAdgMDYe
wMtc8lNPzZszwwp5K+qYgIekGnbKedEPPD+rfDpLb4yVFtVkQ/LclzQYUwjArtt2
D+VoQhu8/bX9C/tlAoAa6s1YrN5+L2TdV8lhzX0XQQ319tzIdvtyJI9NdUrkbMDx
5zrX9v8eMkYr5UN/tcw+GFsK7WFlWy+jix78k6rFCg41OW1lY6GmSdBrQeKMY1Zx
XiXaeWNJMZHaUwC6Kqs+icDB4fBafu02Nsshu91dChE26tehUP9o9fiIPGQd2ssA
t6dbYaVt9p+BBYCUh120cEJm2rNn3FFQD0x/btnn7xHwMyjm+drqP6BkGBtbOsNE
ltNdZB7dXd5HP9bja+pRLCKV+TpsBRfj3JIPtaWVIi0Jb4TgEXJ+kJC6IvuUqQ7B
WlsSHJ5E96ynxiPQnnj9oIuQ8UBIDGGm+h5LOUUhD6icI1WkI+FNzfdERHXN+7p5
0dxDy/tFO0JHiOQ7IAFgEJOF2/oKcl2zYamlfnk0DV/RAP4ISWo3YkLiV7GHA32e
Pc3nGusA/tQsNvHCymAuQL/LP1csoMGTYhM55dttDat3M74+dYL5tnrcytqzJa0+
QFhpbxZIXQ8+uvsuq54k3WhfLEWXfPxXacXvO14K1iG+9EM8lIgsF6e/7e8ol7zu
YBwPyY85CwNjbmoFkpt2x5wNss5kpOObd6b5ZZfSQl8FFCzrdsbNNaKa8F+hDIiS
R8zsJrwkrpglzNxZWLr5NBXBUX9Dl+iPpVke/S04+8z2umAckckfGfSyxbVnX7B8
3hM7K455/CqgetIbiqnwQxYmmUuEzityPpWliuIwvIoDbl34u/mez37LcEzh3iD8
E3C8WK/0CBlQsk441t8yqwrt0wecFb89PYSBlbSxkLSG0hGXrWX94BLOn3hfVf1q
dLRb8qZEstTFVC7P4RFOMm9/GdZmyUhv1XR5UzN/c7zfPGamKxpY4+MLf1YGl6XY
mmoQoY2AtZVkXngmKFWfyYbxYt2l/gI7rTW5HJzpfgZR97NgD6K6GfdGSaFkdy9c
DXQKHUUkU3vg/eX/50ePfOHaxgka/iDuojjMsBHVtUpu66K9XMNuSCyqAwcxAybe
7CUPdpsmuH4nSiLDHB+tR10Y2326/WOcxzMCB5alZt7b8jkf5HxUMkn6EJYgvQAf
/WyWfhQPSed9u28sp+bINQNkYrMFV3zlmlG514ht+avrtjwQOEEU7gSu8+Uyn2cL
Y//Zx2OriF1YVp2ih9lLudYVmOJqgLOPdPQg+XVpm/JNygXQjX8flDfqO0cNrfoW
zgYKQrWeCXAqiTCLFFM8BPuXtV4nTFeVP1A1L74b9g8JDwlN+XywII6bkTcI/6BM
LfXlAYRs4SW5ntOrontlhdf5UyylSjMsH8diCFw2RKzEyePaZ8fzDEvBFb2Q7+51
G9RkBYAy67p9xzAINtu0Ce699a8cEErcnZ9SPhF3GGo9NtQWD/3N3NzCiwWjvJn+
cbG2zY+F0FR//E3nJwju54RBYDclf5lERMvVRwEU9x2tOiw3Ozbol/Z5D1J6TV+U
J2Es3k2paAEkIAvX0tVtqpZ5YIwHoDZA50BG+S6Ez3JTY08belQaxAVOmkWeEqbO
PMou+yAorA8IE3RKyvEerZ/+wX9ymtmHb1dab4FhX6KNACDD4A8MViZSYyrDPc5W
AyPo9hpsaLt/HVAVfPYNnZc49YrSvRorvKP9S1nWCns7VU2ToBCocssV731yvYoC
/+RUdsBRSxBCIoIgb3aT2GT4Pad4afxM+p4uOAyiCFSPQ171l2MUuUDXTBwbiDAT
IY+SmJHzFXl1Gtm9C+rn5ycqgG/2Rtr3aaxDifgKS6E0DW62wBn6Fc43C0aib6sX
D1RQsan8pJFpMKtwxhmprvrwpC6vh0ibPEAb1RZLx7m8/cujKDGl4uFNmdNKMf4T
GavkjlTpnPNftXVQJoBBdvXtVLRXd2tpPyy7bAO4wKuh/N84Wz8wvsj24LRXso/F
raiTH6i2d6lhk4hLQ/b0kOFHV23jfEVBe6JX3PgXIuOz3OgxpCWGopQV+VPo3neM
q193ia371VfUEpLXobvIseZfOlM7bMXZFtEywCA45PiypOiIjiquFX2+oqWog5lZ
k/a6JQjGb8YekxEfe3k2J9GYMSeBmFblme2ZQOadM7qqxHfEw7ouSfCy5NZbecsf
Hxe8sbCcX8LkwfPW94cE41PlC5CECX+4NssYxH4WPK2zfPWoazAkpF9HxLB+O1xE
JeD6Z/AHJibjzdqbaCeEd6aMaK7s/A2C/akbrDbS3a+PaL1w+urQCNOGGNgNfxFN
Tok7dkNWVlJr4M17zA/AjsfqpDv3o/t2eCvXvFvbvochpJfBtJylfmJ7ul0znMAc
nf15u8SqmSp4GOJien3FW5FZIMX0Egu5mYkJFzZreOvK0EWqccsd5hP478MPzllA
VQWe7/n3MqTWUu233BNwIR8DEXJaSli09lZS+VSV1X8eZO99gtRDS/SnWIR1pq8e
QF4UyQHlgJaSoIIYXy0Ow+6m4iJmVejh9t0tT4Q0Tw0hSSyNIpVud5E/qd8thikG
bkJ5kXdkWy3ykekX1VOYCysYbJsIR/CxFq0+Yp2x7eajwK514rPT90ySS8AF3Wyz
TDxZ0ssRr1IyEQsL8zkiVP1dw59yD2Bd8iU5oQkgsfyPYnSVrKDy0vTX87XZT5LM
sPn4OhZHaiSbFt/IvDlGbg7ngBJDTpV9GJKMMrkIKH9Y9AxkE6w3+I4A7EgVyfpN
XtXe2ZVmrdkxhqZeuBv4WokAFsDPFrmVEdd0vHgTRSYNe29QInSHBS3bPljgehwa
AyLOSFrHw2HBvpGXjAaTEVKiBInt54v7r5weF1yz8HAAVuK2DTRXzh3WwDo+kVIK
zIKkj3bEdWCIE77TJL+KvTVSUP1le6d3aR6Oe7tjL2ToDE6YjC6Ax/hqL0IqIxM7
pJQWKLbuQJNz3wbbSaSfNpXfV/dNol1hEV37bYwWd6Cuj47CaVovWmlDl7aRFajY
9S72+wYD3QmKDX43y4XJXUuyp8cIpEHQmE180EdVv0vnjQ3dasSsMTcrtcOWYYgP
2mjcJrvjd0kmFftJZU5SUogpiO5HqaxHDu2WdiOCPVKwWz+fLznYe49oEODNchEP
p+koP77ln3QPtgWpVMoaxc/MI1YNRAWvNEJC9k4WyokaqvsCmrINh5tBgcx/vNYj
9FtYZTg50Fj6lEgYR5494hQV3zliLmNF9C+iiyUwZXbQQWeqcnYSNE5IBXJ6hBsV
FJbRi/vIau49GhJejeKipt+xnEFko1GJNhQaxT+D7l6dZpgi66X1y7VJjfdcxqx8
LON2USMQ/TtA8p4DGXZLUA0jqgqVpQJKlrtKhqVIIPkWufuyuB85J9ZvVGaIeTrA
IcQn4n0YHlnjhRzopjPo97cyt4far/ShrkPAcB6pl76ZbTkUDLgRTdFrInUIV343
KurrZcpWyO6fHqrEg/E+ZEylDVhKdZX9st6Y4YCoNMi3fqQvzgw0Y/a3xYRpje/g
Q5Yq8eQwH2BNNqQS8hLAG3sypZDo68pWVBpJkDqsUD5vS51jUQdgsePqSX1lwxcK
jjSDoiqJ00dJxxmfdZ782z4MtcDd4OXdrFHD9iyoUfYlw3h/Mug1LIbJqVf9Qt4q
CGiA3vxM6gr869nKHSVnp59N8JEk3/BCr9s7fGoHTszSo6YaeO5APCOtudR05ucs
sSq+2isQk61Qfa2Xc2RuHHoAZQitwmbN77CWOc7rdfaddaXmpvn3Vz4IO/T/tCvm
y9F+utnvpp8DiaqI937CVBd1v8n0RbFeC1Rc50blfP1C1dboLliMwrV+OWDlYoYP
mndn1sJ8t8yt3oRgXiULgFbiOW5UvANE5KUzjP3qTrbUcq+9CHGyma05PH1BBIpx
F4LRmKsTEaW9BgPNSxowjfMGLxS+yovsGa2u54Ok26cZxV4TDaniz1fYPvDUME7P
xrg0bT28EIikMGOb/fyzKrKPG6b+KryU/q7fvleAofjxoDNWA8/pV0DzB+8pebpq
IGwErE851HUk/EkS2jbVo9Byc25r2F7JleWXoIxVcSep/V7vVV9+fiR1hdFbYxl8
iv9z73NCyYo7FxZ5KeyO/A37EL71rtb+Ja+aJdqLX1mzmjF8JaM0grOBg01XFr4/
697yr9keZO4RxVv/P66rV1vsZH/MO56GGDBZzyAvKa50C4tRm23RxzwItoyrEytJ
SpfdXWAl4Fph0XF+4o31/0ltc6urFOezXMqH0dPJouSEoxaON6K3TgX/Kg7zuthI
DLQVL8teWDiOHpucSdzEZpoSOkE0mcEeZhqsiVqoIeba35TQ85crAeZOMcBKNTJN
86yvwjaZ1uGUI9BqqcDBJ8zPToHkNGWmB0asK54sgK4S/KxZBS9VTwau+c3E44sl
fuNK94ONfkd+wNubbcgnB01qd/pRBhPyNpLGdiWdrbHnyAebgzZiwV128SJ4MSaq
oFD8Q7cEnMeW3RAgzWG14WRr4UzkKNkfhB0q2ujOlW1FHbcnwnybJyA0JqJtGaiQ
wR2hRGR3xB0K0DGrkec/NlcyJ9Ocnwe2DG2i29TKOtQm8WLVJa2mTlQY839Ex65w
SbCjYpRinIYBGsu1j4XlLJfHSw/8ndsxuDPNCr+ayMwQrb+meiDzoNF1/nnBoCEA
gXsu5EZHqrsC7w7gEsT7q34b9Rnj1lqMXHcW/YvlaaA1rEVRPhCXE/AgZy3HEJoP
kbayccsvEUyol48zKMAXXwKdRMH9v9dcmbAtCmgvSZQqMwKwsTuozyuPTorWqLGj
m6GBvAwq0JR+Hrh270FD9Ko5//tBSOP9Mrn78AlM/61ZEu1P3soknQhujkRDSE+A
WIKTJWYtvW/oP+pbghGreGriG3WaRwe95iB2iJV95sqOIhY8srodTc/EG1Vv95RE
eh/HWBALdryELeFcisTdAgJBVlQ24TNhZNwvGXGq5WQiiS9qFikku0IAFlhHnZLq
pUDhLAfqMgDQP1XRWBqx5gpZFv77MEMkJyIvKWWMN7s5p3gWgxGnFUtvGXBr5f4k
xqoyDWHk1vAzWCfpxVROABOBZu3GIElldOmRmEdsHX1idhuZxOrVO4Esq6hcY1JO
/y4MgCZ2VWxQD06izh3NPsnoxdTf45g8C/BjFOlGJYSGZMFpJCzOmylTmDWQRG2+
KhFyyDrgTppPBovLgeljs/w57LVWlj7uNCRHfKVomb94s/mzvB0uxgkYoHfKuDDi
/YXiZ+76+bB0khm+Wwoe5ngFA6i9uImWMSJ5TkeIBGB3NRn5uMjZ///upoyFleTZ
JrR4lrFlXgUN1ks7hlF2GaDc3klgCqupmxqqXYlJoWbcVazcnj4lMbtu5dS/z8qI
63Oj3kugwgFpK2sfK+4HP9YFFtqMfunFk4aC9+ax3+XRlGDNXpCT0MsgYeWDzeDy
Aior3hVCCAdjOOPK17xrb5pY+TSlDE3iYnR8euVr36qXDL5pDfkRx6M9bQDnPlkS
DPMsYkv6RuPJF40k71Q0ZRIgsP2hzVS6xGG/9hV8SWJqVMPpYixo21HF++1cbkSC
dcRn7xTIRPIsEuZpgqdjbIp+ggc3xV93HX3ZBsm3NXTDNW2/7o7F8xvxofU+gFVN
uxH9B2AFGYgylYGPDz5wj05RYaB6xUxejBmQ1LuS8pZBxnalNY5nBwupOtuGIljN
syzaoU3oOvDqmhbJLGEuSi72vbgBzArR+GsQ5X3wNpi7xxLo40bkt0f9NzyvRM+S
o0awE1v5y8NcfxxLX5dq/ZpOZJscabpUpRgm8p6j0kGCUSpfQwQBc80/IbNdYlh8
5UwnqM0lrfgXMnWoWcsj8dVU9N5sW6j4FhDYC4kKw5X1XIi1XWm6MUGRZ6KQCPvu
fCQqHvXkcgoEOv82pIX/k4hv6iV5r/+q6IF3U5Bq17Q65wu6Is9EWYcGIFveiR4a
5P6tFoNOC4p1BvJW6B36LrDewPFYR7K9WcXs8XUOxZiDQ1h7TjtcCUStwGdg4cHJ
SabotIfAO5oWM+7vu8HmASQ76qBCR4HpMCj5kurf8Fm5ccWCrt0W9P7VarthsrcU
lpsp8DGJ+zBWla7tZrQ7g5kwTPhcJY1rl7QDFXotHoVUgLlINcPiVCpriJd0dNwL
bS4HUPzZrWDWDsfZhYEvxQRFn4Kbp0Azv6xICNIgJgUpl61YsvLrBDuqL0ZVy6CT
Nd/egfOnG1NWQEY+Hus9cLOoveK35wCuAx9L6C8668Eci4CX9g9RXXODDFBcGzgx
vtafSYOaIURTVi7gWK0DiyjZqEnwjn3ySNKZOvJLxirLZ+cfYUGCytEB0TVOrJzn
Y7aqEno1UfmISKkEhs21HUSiQMYm56xviDniJfqMYRzI6Jh496a80GXbBCLdTRJL
Pl7+gH13RMGAWXdVMr9yRd0y45nFICQS8wUaueSOBADOjY3CWl0niVjrLevwqOm6
D445W1+ZUNcMAoPw4bKVjVMbPFH9GprMle5Q5BRJoSfe1jBkOy3/dXExuCfISI1W
bCQWBft+IMtpVtu1TqjsV3obQ1CAKVS5S2bfN7UZHitJsr+Z57VDw/yoec4Prchf
3ZNxwxpQVI/UKi6H+rCcIRKzlqsIoLOqlCCZzb2lfEWwcE4I/UktlOSvo4EHB3Bj
Zn/x/wSRBX0XFdiBZRF/Ny09yosAN1w3HOdyzOe42qATz8f6HpDHErR33r/uuvHC
6DvJrTlqGwApq9lwAFmYDkM8yCwoqVpZwPr5tIiMwMOx6GH8nkkwqU6jcF5lhXCA
HdCZfENXs1FFV8hbqUG7aNf2pfxzAlM4s48tJMmi5VfypK+owvi4KOPukB8YJOVI
x1yqtj05jPaK0/8e/iEgmg6J30DxXX9//GS2wa3RixM5NwSGSuNxERZqFKIYOKf0
PpZTvNdCBtMACGyds0E3BlI22Kvi8LJMlTQ26PiU1h13vENV/Zyf7qBNAAxsDzZP
4r+3ghQ5JKmhzkPesbGBhPmn6TnSckpewFmCet/Y2/I0jQF4u7R7tJMoKtyoxZ3G
K1yONLwr4tlCHXmVA8Uxx8HNONPBVGyCmof/8tbKsBYcfNxv9jIQn068E64mc7Om
XWr8YY8PUvteo05Kvv9/kF80NDXO+t3dYsGR7gU/UKwSmO3QgmXUnMBQVZr7tzvA
B9sE+xntFTAoBgB/I4NrocnG93klmB0/nvfIfSnxXaxekXiuZkLz40cc4XjXfEXG
Un9HN2oE036AL+J4AkiroAUVnNDrBcu9Z6MDuTD19cpc7PLB0iKwbccz+mtsGrIt
p/kFbjR/ok5X1FkVxMHKQjvh6oU1dZ6RCWzCP9pa6R6Xjlz8P0IePHTOfg0laxmh
vkuuOp8yQrkBqQPXJeXDB0cBtQx9vnt/P1TT5C8EYyK9Vif/gYiHKDkEtVinAH34
HT5Ipc65uh+xcHN24IQqPwvnH4lcu9PmOW7hNib6ORKpZzr8g9FXz1ay5XotJAJN
M4we0Ckh7yu/vNdNqGhLctu5RZ4pC2PW/QgG8k8sjBOlQxFolz7k8xwOZ5//CU5q
KARVkD5lAMi2Xb5/qgi/TS2YdDwmk22ia99zAJFvXHpfNrXPlEfyDvs4SGgB2QZg
2JQq2o78vCxlovNONyGzNrVoWq5k1iKSkO340lLDrfzUqmIMas4LKfX70OXYfeY4
yspg3pmHxYa3+F6JCRTZEaf+0z9Hs8jT0AU4pPeM+40ftDDgfZ++td0JpyiSVmA1
AoLwPsWc0ImnB9CXJjdsl9GCMVCuzCR4zKH4UG5CNmK5aCOv6b+6UzcZJsg8r3A+
2d3WEbLpmMT7DJs36gcNdIBTZ03RffbVDUIBcZ/bPWHML4+JGUvWmEd1eHdD1SnR
G89MjAor9TlXiOAfw7yUXwsWdDhA0QXMpv9xgmXkUifnZ67entSwUYykSNFpwjTV
q0G4OW4BcFDjCuQZniut3Osm2wcAHDrfJmodcU3ofVZOVnHCzYhIAmfC8fkSpqB/
FyYXzLs1HWvteZ8J7MxMxnIpNY1bRJZU8jW8lLngnSSV7MvmYoTzrrjgOKedtZCl
Dj3ToDppsajRKI9/l2qYj8z7ir6ch3IzW5PkJIFehEgkzpCU9rxLiR3j1Vt1FNtE
leElw3sytRYtmIIUbq21HthF+tKX3smXw7fQ/lJTDfNae2AQfLDFY5aKuwDMV+NA
fRlE0QJ/AzkIwiJBjS4XltQOqGZqo7DHPPjnbUtySZT09BMEOwc/O/7QvdqlCH2f
8tKweBxj/JJQJ8muc9ixW2w7YkfR8Msrg7xOefcY7Wk+4AaA2d6OeAn6llelvh/P
aOXC6MdOXxOq9eDpYNO6LXWJ6H+11VYpZQNvgADsrEjfubblZStNszl6aqfjRCos
QclOaWkWsCmvElsmJVTCRMrqvPkIqNGHYOO2cDBSTGpSASRyCrQ+Cy3+Dn1d/jxL
sWuxzcuyuIu5pVtIDZme2CUYG5EH1MBtal1ShdTLskM38Rmscrp+38NrRphinp/r
dUqoN8CqL46pGAT7Wbgy2jHTyUmHQwbVOGO7fVZqqIXBrTQ6CAjUM/5VV+ikTBbY
PzSN/mXq3vBQVEjJg5GKrMMKgwO7gx9VvGanUtBPS2jxQZ4mksEbzKszMVz60dPk
R9NVraOZsNA+Eowvwqet3k+fQJ1LexHMNmY9qZnyr4C38eTYnzFjAdZazVcNyczN
zFFhc2QirHy7aHFTb0uijS/KJ8384LE6GdfipIr1Fgpv9LLmsNcpZRlBMjBkQVnA
jLCcCx3IMsYBVuw2mTjxVE/T880LBnKb46lBgdoV00lKijRPrwL76SVsZcqf0nuV
zHsnSZRdq3UJOy1jncLOVuL1bAHRYpUZdqWFOzuBMyPP2AO8cndeC4PVkgsYA5M8
BXo9EiOZlRoyg1LciJN8UZonjCPJIyzca5KHVtBc8z9l1BbNpGlhKecJ22YvLerc
nRNyMWfeow4zKSTgBNa7AZQR02RrOOfZ83l+0TAcm1zyU9OoKBIArARCpTV52OM4
UOEaLbzpZStA8oJOPJuEc1uSHnGefpMmbVI0zAGTcvyQ3120vGJcUmJWwnWlltqH
dQKE4eYgurWcxc9FHwbgtCNhf+/Y0/v3k4PBxz+JFOhdLWlQXh+vG64Zh4Z73G26
ZrGcSwRgfpUAvZqvSlBfnZEB7IR0DdobLKSnIrSsvMdJH1jppc2RDShtstf9a7wd
gddG4dwbkfB8vS82rbZ5klPFg0ReVIDS0C6N3tnv9V/tysGdwUvRmj5XiualYCTz
Ed6puPbUFvXh78Ct4gB+r1yRL/XSoiOexRWg6pTqZllHGMkFzihQR65IjiAXyFhz
hSdFGZIcwHoO90SuLOf+YcppWYprXwVr2IXkT9TtOrO/eG/McFM+WFjIgxthIa+Z
aGGATvVMAs1xJrAU9GDaX+fd14QaJGTrr0LO1VGbI0uzzsCMswmPHECsc4dPSeRM
HC4tFBeNJk4xMI0enKLV52sgl2mItCLknqW7wmNPp2ruZjizfmXky/tFw/+GC92Y
y4HZEfs4uUnNYr+3VveDUh2oQRABoq94Jy7l8CfygQL85oJULxV5aBfG/Tm8bp4v
+f8/F/ZU7eu1C6ucyI8PPJcgB8XsMlzlqC+i7mfpb8msOd/5ho4DFzggHOfDen2z
SqDesAK3nzCZ9Edmb0DctXo6RRHbJIw5YjHv89lRPeM15bbtRJVJXRpekAaSWObp
zBRLF/3vjed57JEclmzh4dgMGY0YYLn6Y8EhlMRrlfAtZtpEbG+wFCG0EVqfEOdo
eygFLVJWePSRBC807Tvm3mE4anJ1fHclScT4GlNcrq0W/29v+ulV5F/fQwQETITn
vSglxPg2IgT6sYZo+Dv2l5I+cQToHbE38qYAb4b3dok9tWyPej88aBoRaziOahSf
j/l/IMwsHTMfxVxWUGqIBIcYNGvxTzfe5a/mI2SYXlHFL0yC1Di6rj92MFI/OAln
iUnnsbVMWjhk+R0lwYJ7tdPtf/elH/i4AnAM1l/3l7NHyzaQteGrW5v7l5d6f9rw
oI5lFvGzo4gqQi/DoA4Y4gVPQst2dhCbJkfwgFAD8YOFAISWGd0s/XPs6/tkdHoG
k6uEIyJ4xZOVDyvFQKSDjpeE1jj3esK3D4wpGOX0uKIDbNKZdulqdSSouGwoAntH
uL2X4J+IKIe/9l4BxUTwIpdL92gQL/EHKAETvG0gDgN5gCo79PHBzNdPlkiNkL1j
3RO3nrjczYZ0+mwg1fPhlcbR18DT7aXJeVVsh5RWIVqwKKBrrVdAgTL/UmDBY1KX
yYr2W82Zakw814Q71vvAH3T7I7KGzqY5KPz7QMO/bO6PA8Y9aO/wKxGZgHgy/W8Y
w0retP5nnxHx47JWLmEEtNoe3lsvOWnr0al2vD/g1wpnCfc9tvyZHT1LWR0p57uB
xGUntlPUbIDhnTXAbOiN5doUZkho50N7WD27hF7+bSFXw95DOe1fBF6txg+sffzl
jvao8ZwSc58xXmtFsTZEMROJLpNNLAjl61uQeYqrQUMEczRlz1Uz1CUe17ybv++8
ldMQpT/61IaRkTqs4mcw7rhVtKpk9ysvK3Y/5z4kx9Bb7GomNq0nFp9YsiY8c2Cd
D6nmLZkEeDyGLV+mwZawtnQIEsZX9/nPua6vWUue41zctLN070rVM1JVl5gGAav5
BpNxJHaGNG997XkM6NGzYtbjBMBZvIBT9uqzFmR1BgDAswxz5T8BHo1gDu/OIdDS
sauTD3mm6TxX7rz+Aj2VMinp9fm5XabSCP10GAJg1mlt7HM7mXtwcSesZy76GbQ3
rP+fcdVqVt7APvcfKfiCJC912/tQfLODrs6RyuQ5sdFxxDtLjpitpoFYfIEk4Glg
biV+buh/Q7RZKVahrmqHl/hHa4S1+fKLlDITMHZVJerK0l7IwEFYhnXEZYyVz6hS
VMvoOKAXPmy8pTUPDsLJ1WjqFBMk0jISWK2Iv31pM/6SWpeXoz2vWXWz1W+wAlCx
bo2HEQEWyCypqDoXoZNxk8E81V9mHgUAK3NJUQIHc8FHcNf+helBCH6e1CJxEip3
kdlBxeE3lPh31fS0a72U+nMdSZOocnSh4+bMm6Xaqhn+6leITaiS/we6V3lHly38
wOkGfWk6jW8mzRNU0XXdyfMR6MF9lMSfK/XkkHEwwAtbjkqj5iIdQxoD9euh5cDd
wQncYnEAIpBta9x6oZqVt2Lj1GV/NOvUGhQ22N5AADXrMvFbwcDoh2PVJedAwQBI
O+kSB7yQTfrNJEfQJSmzo0DWtjpss5n3rAQP16RQJ/VhVz+TdXZ9cn8Ra8X7JItF
Cvf5Nvnf/hLa4uSow+h+vtyxFjU0hHRgL2ffAdE/pv/iVyNev15yOyfJjv6LWxci
n9TtzufGfZZBOQvmXk4zPnz+1ZPduHIZE4cG3i1XjCilWXKzA3jlVhJn7mZgvvbO
lDxO6hTQYf5h+0uu7Rzdx9VYy7c09fEdIlKFvWy401tL1KJDOcBYuE8w3K8ovjdJ
5uet7f5JJCqSKceiwro2hPTgjmyOzxXam56ftwyXzKXpO5DH6EaSjCV6IV/GNy+G
vMArWoRmoHpcJFQfct8cd/b46gzGMvJeafyb3A/bTdqWxqaNBJ64X8QC8uNJdrs9
zRHzk1sZsfG7R1IANts75ofOf8M7uqY3zqmegE9+KtNLF5L3cq/XVhtVTL09nZ94
1HR6oXvWdL0web+9ImlSqXrVfBKvC6IfdTWfbfB3xxHiivrj1XvRVe1g15kwU2He
GLwYMHlk733QhfgU7Lgi/qffBP+411qiVfZvlWjPJpkxnXKXaylXVnVUWbf1gNV4
1ET8400d6rt9ByyNEbr0x0Towp3zKiEWobUWymIxggYNN9lw1+w4/g6vP3+frenG
Z7sWS5LFHY7JE3BcRAYmfrto1F7z4GhtWsknOGWqw7tn6VWPtN3Cs4iqNRHX7j2k
hgPAgxwc1qL+RSZ/X9Z8PRZtSDyf8c6xPmrNm6Ker5Jewg0W610DqnOxQUdfzruq
Kccwq9tM/aheuMaptICX2eanGvVDo1l/XMS8bSSJzWnGYwCrX/xRl7P8zbEc8e/t
FoRGzdUYMFAf+o2U0r5ZmUGaN+aC01JcLysIIM7BzrIfBfUVTh4roeQZ2KUZUurn
Su7QGebPbRU+KzV9O9reH4OEwyxUUC8v+5KYd1t4RQN3fmiy/4rsUMHxXDm54O8A
1v5O5e+hzG17NEpi7UNxJQSlNWqh+vbX3WQobq9/KA6lsQ1hpMYZVheh2ULBzMLg
WJZhRBA8rcGTBgg3JU6dOpm/055gefpdS8AUKCpbxtf36MkhaI8FM6AdfaoOqo7S
633tBQ7vNQBKXZrMTlxF99YVE1II7mVoTOEdyaWjQNr+xmFDwNvwnJAzdn1lYF4/
rr+Knzh5LZ5U7dnivgcjndgrwr6RIUdiiitu5rI4o0Mjq4gVlJNR/mU/+WNUEqZ0
riDsSeeznz+UNPb0SSIU6kSpTKdDvhZpDhIsVfvWxX91zP9q9hD/9jnbwDHkx7YE
+Zj54f43raf49Ty6cVNWDeuz8EFtarZJnUtzOamXqVCROhfaNfWFhYyoB2X7g9I/
KgCNZOJOXkTqWPx9xpxYgbMoH3hrJ3Tu3F+znxBnXUD4IUYeNt8EuLVLqrvydtI6
1eqwNlXFtd2DSLWFnpkNMBl2qToR4ZCwpT5eiWrmGSCEQ/gORvAWwU4IRiaaW5Yy
chPF/r/cQCFfbbLr12n3m/OafanJjsCmMa9MOogEvyVXxoH2O6qrGJFy9SEC+G6R
puJy9Xc0tSYirFJ2ptrRAV7yb7MJ7Ca7tmxS0wg4HDhPJEPMlth1s+v6Rh6Z48ax
QQqwQuNomL467wPghTRW9bf5WBTwfzsNcLM5aq2X1D1w4VLqyvY47fCSlnU2y6dO
lYbUOSDBN1EJkMUNJQxTORU+ItlFaMHYI3RKJUYhyrVy8TzFFtafXsUFJxQGq4an
Azg3bRtqj2DCZ3uKCk7TpJFkJZX+hygDJuDpjmQZOPkFF5MPfKqyfI5a6cXYDpzb
P18O0P/1b0DgZP++ckJ5uMEYfCs9alpi3OGjL/7feGC6AJAKO1oXe/Sk2TfEQ/H9
f96sjTVD2NnUXvPEKZYMi/5UcYWKfZEhlhes3MlqaNCzjhdENyJaT76rlUfcokIi
IifTUEUka81V5pcB5mjd1wi1ink3yycNP7ZoWNLLdHc1zamVDR2dVB41qZ8fIBw3
KeiIcdCEhtAMu12ACSezezeHIo+xo6v3Lfx+ctCRctnpXOQD67XJmELrUR5Fb7ND
daVdPWijpcmud6E7PzzxJW0k83jXrNZ3kFscze2LHXhsuhlTM7qPb/4qNehIfKgT
2l+A8R3xqC/WJdGEOnOE/hGws33B5k1oOjAYFdwuiI2aU5sACW7Q1dXO1OXjhrak
7RBK2kwvWz79BNYaM8tZOj2nQaRpfbOtegrVydvltyi3u5NDJVrYjknHynrtlywg
5wF+5azeLzh+gXP9BFxBINXM5ID4C7s66tcLzxaFTH8N7eh6sc2m8ez+kGO9FVpE
z/ZbZMwrSvxca5lHEmJ+y2q7dnOkdDbIOtny5d8tzsGUGa4zb9zKoBymsNFeo58H
pa9Ac28Dom61kTgU4uoqsrwZqC88wrHUPrB1ptc3y1RX7Xpwg1dcUD6dNosencrP
ln545k6pWPFbSUULbHWAQ7W1qqyN6QxKFbhcIba5w3889EWEQONczrd0WtiF7CSK
8RaF/DZxUUb7mLQB+uNoEUny2gGY9D8w3Dg4akqF/d4blgpGaD4WE43o+LM/ATfx
K05McbQBqGSFQOLFirY89KlBtvK6zppl4FPVxmo98YdtOZBug79JlaRqimfwGDMD
VuLosiuL6StypMTjEcjHRKPrlBd27xHu7PJGeZq1n8rg8WwK7npSfi5nqFtdxHJi
C9JGII06OUvQjjHAWfKug2/ALhDYqjLCa48tNS2HnIuERr7krxOOPxfIfnDFLl77
k0CoH88aIJP0c/uDLNx9jSu1EeSgKUcA3wOE/ECF8xDBSgNwbMo2HNw46W+zYWgq
Z1K2k8JFHIRoHloEZOqAgWJ+6Lac7vQq6NEf1RGY/wGW5CQtSrO3xH16eABSqzmg
sJjZiyPcrFqJFIBsr6TKcJTaq62NEppfnKGKTfjFmme7ogwayfHF6NKFUAHsbuR5
fx3WsytlA3UkMchEPKhbweVIYQYaDEzoThXm8l0dATQpPI9DrnNkgodavy2WaYjl
8yTxwB/mpB/LOcZg5x3y0izEXN4nyC9WmghvRyvakw2pHfISpgufmgOAvG3AUfHI
2eVQGO5ZDw5pONgmrJAMNUGrfnyirdmCEN5uErrOz73hyL4bZCyZOtu+voHhq/MI
Id6nAFPKOCLh8I2ZIbwWePnMWJDWwhy2YXkWascTy42GZQgtWAgB7x/ht8mZawm0
yXQq4rBs1e8Tu3ZrnpvVUjHp6y3qCsbpofVXM09clLSVrhNluewgWkqfvZ1UjvPq
xWMIBAkRwqlCj+DV+1IgvLUR4nfMzdeKoBEyuQxTMaCwyjV1/exbf0QHotv9iQ0A
4El0FY9O6+3l+RYITUCXX7MkKQP+BR3yw03YaCGFMB4dRQbJ15469P0TxkBnlI0f
UbVcUEnRfamTmRnet6M6xyzQa3IA479u2JU2Z2+AddnkLXbG2wLHtsgPtjzjT00Z
1FbdehnZUMF1sz6i3lbmokF0I9gxN2rUbWqvMky5E+8c4lzwlwkqbxzdDEgy+RPA
Dy7tL8mVv7HKpi10B+T0zABTz2Ci+N1n46P5e4aZ6LphTa6H/5jqJ1K+qu0bkEXK
xj9hdPcEEWs+WEaRHN/N/wW/jMXy+zQAkdi5f5wQ7ZunjcYNA/dUoWcQD8JJjPCY
2IFuIkVvGt2dT62UQTKdIBDEVhxQeEWJDg2c7AoY4Z3kc5KvfQ19emYka2s0IRLX
pbMTLKnEvIh+1ynupaIb2M33VB6AY/IU08jgXw9wXgV5OFPDkjmD6XzAx2Lpm1Lp
PfXk+OlFaquoYdn7P0PMkPudUFUemNZJn2xdyTPg5CRqBvojY9h6KSTxqMhvkhp1
jv3mqz7d3JlT2qLFG9qmlkD+jzyxp4KUkoZruDBoFskXCfhRkSXa6VYoqzkoGxjC
PCBtBYeO2fs5HLb2r5r6YIpTXv+t9SSh/xAf4Ml+/U1uwpHLq4wTYua042hjzSg+
truxDWpbH2LATGsx4O7Gpvf441tI3j2SG905oKHdf1eyEYgcIJbL4dPUyDRGPSVJ
p1Yk2a7ojsGoTPLVqA0aKQ3jj4FsvOOLrddGvwN/JWzrC1RuHyMojUz6DOgABk9f
DVdd/7mf7aTiG2hMkbBZIHc2C4wfVFwEX1ZD70wtbsvBGnHWCS/0XfEuEe+QcTkO
9ahlcg2mt0uRSFDUz2Y184zPAG9Hc48KZFqiMCjz0qqUjk0l4SCg5VLU2HL2o0Ew
gFLepTGdaG9AsT/aXn+DVZw+TDeyOxoNIFews6qzQb4UW+TiPm9ncHDlrDD56JWl
5drkULKQJ3XzU+K4gt/hdRhp+m2LCwdNOHMpiHpMt/yo+4uIUXCmYw8kaDvdsI25
XKDGEsm8B0PCjhJoOBbkzhyILhogEaxo0eo+ZRLA3Rgry67z3qMoycavxrEx6d/V
vFt/1mIQRI9jh0Y1gt1L3Xp5F8kcKLRLPAou03O2a8rnC4kf5uLSU1etNUtDm4nT
8Hg6CRgcppGgmm82AA3mr85d0kU9sKC5/bE0opKapOz/89IGC0tHtuttz7JzEX1H
t5UCbUwYUwWJ9Y7SKNPhzPcT5FugVcIFOKhLJ1Vvwmugg+P8Sdx8a+7684/1T7pJ
mtKHuQmKsZ4KAwEVvgjGHxl8+5PseMLJ4glRiQGVfPJNULAXMgE539yIa0DMOfRX
xGU5ywDBeMQ43AtZ+uocwPHcWvBOxswcHMxRE/87QJ56uWBiW7Pucu80wJygEkSU
k4Ay0KJr0cn/MiecWtVzcjem/MvsV7QRFG9iWszlm1rQJHE6F0cMYtL1M6GBrfGu
U5mYc0U3nvhT6IxKSKjT/A1bj108LS9K4xQ0rn5eqbByW0O8mF4CC5qd5uphOd6v
+ShPZuSlTfBL709VqeU6i1Rx7cqB/vM1C47Pm88yceUtPN+v3WvMsHZk6/WiAh2h
4vaPhhti6flG5ij/AesSsmvXfkpFpyHkpVvKVTmjqPgDawz9BzyGR9UYLwy2q85F
iWTvra95VVX4BAfP01AsLht9ke/w0Jnjrt1tBnnaTu3BP0S4QyVRiDDgMRg15goW
UocENB7lRvDZp5JpdoWCFxBd7pyp8o9iWpHdhM3H0oc+ZTUdboFy2b8+ei1nTlqY
WhK+4IMpD8hJaq1rDOnasuF01fgKxPB1HKjKbFBeZpHWaYglGCVCq8GSKpcf36cr
zZxwASiQj7dLhTV48J/P6scE89qWY67Bd9Xar6k4nqGLyH+de/aWpzjJzgRtom2l
3aQZUwGehXJynBNNDfwup7yZL2gKk7kfR0QBEPpkMEFPxzNd1LtfFmIZ4s9TaVhh
/nBaw6CU2Jb/isc/beuuxgS96vLQpoi4Mxqi6B+BTa7g2Ika/3YwfHhJ5EcpgQ00
lWBLNrFLMysFt6cILUCOYlTUoLRZndiRI3vdr6fJv0GqqLWz+ScDrwgdK4Hm/60d
Q4DwLdgDfZllW3gsYJblBfohd9l+4pq5RKSf16vgwnixdjm//vNJb6DBYFannkgg
7NDIeGaHE8oqzmjFY5tRY9v6VyvGtV62H/hULs1fOV9PHpzJ6wOK/OhxC9sTzkNF
OTuVgLSyz16eRGiaKX4TUZiVKNMQl6TktZ2JVram8nQ1ZmDexXsIcCOCEwxW6rqD
vbKjRwsDS0B97mBVlgCu58HwxQekaCCptpXLXc5Yhjel38YOtDNM11ycf3YxA1k3
scemxvoQGFyqnhqpHgZvBKOefuggmZoBSc6gQpDooWKx0zbm2M82uGEg7x8RA8fG
jrXaKzdB4n04h0Cl806wSWyzOv9e9azMVxDNCckwuydjtekgDx4cOz+7uZ/RCdy2
A6ygHeFCsw21o818HFCmt2kOtjgJ9wUhNOoapEzhvhuhhYlsWFSx3RlquiUq6NnR
qEjUQW6smC593FwtZDFEDpwiw1zkxxVTN/DrmB37d0fLG9mgvTc48201vQnI2LxN
bxeuW7g3SPE05HjAY84DwLPBsENnlKh7R43TczyC+uuf7XmQmXvV09Om68CN08hj
AuJXHGuxWsqwY3AigM44N08V2lt7jX+Kk89fegA0RHMtl9KvFpTxoHENpTd6v0RC
fcdy5YJyiaOOOqp9jOcewK0eft48oydjLhA68EZTeVDNbML2RcfqEmPkQkesWanw
sZNUZV5HtARsFkynEPZVrVclwYFTXZXP1/dtEQBRtk++/ulQOvgv1PoeGZ7Hdpcp
zQ9e0CstygORW9lEhMT/e3UzFCFDAs+pGLV2ghAmmV9j5xrNm5ASZCkQ363nQV2G
fTpmAKwEaphXr7Hzumj7lGcKkeXOqLU+XseadkuBHl4U4APd0yHo0QoYRhUanupZ
CYdsiF25OhNdX0bvpZa3y+NqDOIPuzhvnWaGjWyGMOSF51ZxWVh2x1pf1gTv/dYr
jnKCEJjh3++ifIv6JGhoSh39xuJYJQ5C0HRsOtZewbkSaqJZgQ2sq5KzxKpp9Hyi
Ho0ZbnXJ2/ylYQd9cpF+1qMQwuJPTKJdEvhBQD8dRXrO+PdIxnQOZgEiZxlwNxne
WSRvzLJI3NzMmXCgmT4UL09s4Cjy+/t4NfkF1WISF5ewIjB3t9JweRvvxuKLradV
NFcwsyNHmHQOR/JAeuBiqgDD5gLHQBRGKeT2BQ2nUGymMPw8SMDMu15bGUqAGyTs
O6YgHwgZrhO3QTpLJoYu1Z+XaEwxChwZzE8f16TOsnd+5PpTxStXwYhUY6XyLlYI
Oj59JnM2Vc7pSo0Vp8BrC5322emlfId0liVJxNtInT2LdclIuh9y3xEVN5t56SR3
RBzSFPAhzbr+3h5JbhUXyIClx31CPMxmd0O2pyboiViGvLuSqhRTQOu6IPSHf6S6
XH4q8jceeOkxIzVLZVcepf/6TJMgGXNsY4kLHEXHqE7OGPwlRq13JkG/87Ofu6Mj
vXbKbIsNPmWYm2fLMsm+vtiHUartpEz6HmP7SKlGDbP1glF04i4eN5dgPRRNoY6M
Da7LN8DwC5RtjvZbmTrKzAsvqOoFtproNPR6Z+huDdbV2znWsYfMWiXF2G/vYpal
FvV3hpgzPVHVC2wxMc5DxedG0d7oy4RXg5SLcz/vG09iyNJYnVsRlYnEYcqg7LlV
PIxMOGEC0BYYUWcsKsFJb4mMDhtPc33h8UBE+0KLoSBY0L7H/ESAX4y6E88Hah43
SLzH4m0b2aWHpn5nLVZA/n7vV/BfV16kCtg26gsB0Uw1/SQRjZLLpeAebb6oqVTD
NNOGWMjtZBpVM1wKDYtPH2YbJKeNpE9MbKsUzfPDj5ai7HPcKTjJR+OEWUtJprrt
RbWaae8vc6L+11A1IDnnwQdkWnvTodntqmXjIZ6nY8n0sXsXMgBrEcmdfxL1Qwiv
ymfZx+o6ClXB5I/vaGe6e8lHruez2JuSWAAJSg9+3up0mjIAngMpUolT1wNQwhia
8Zf4j+Zcz/jxNoX061t3HSTREBhp5yx/qFTmlDs1sf3U18vZkxIwt6if8I/5b6Cl
/j66I6BRDGw7WG0bR1/vRtNEZcHHJKkglZCaVIwihmq9MwqsnbZ03076niEM/sxq
tYz6BXfqVWCcTKX7hHbfqafhjhBv2+YPJGpfOLwOKgf7kleNO9IE2blFAxDsjRbx
V2fPPYbINO8vBpTKxo48arn7JOhJ1C8inKdnqGOAl4FwjuG+BDalZRTiK8GVhtYt
Ce9g7Nx9ad1n2gN1yo9J7MWEwr0Vf9k/0OoTimlPpc2fk/VOlBen0ukfzeEomjmF
0w25SuO5WRdygwvywt9cKvRVOhs/e0i6BZDo/BRAiSPzxYF07vyKMGtIreSDHMkf
nwWzwjxlRNgd2G7wQCycC/Q/HhphNfT622GLJBJj+E+fAflI3Dk9oCZIMu0ZAEyb
PeHc+zKtaZ/OIYk+YKal63Ow2aEh9FZjWZH1JjITYjUqex6epJszFFgA73gyO0xc
iwTIIyZUAdMDCgU5GFIIzZ2qQCW9SzgOzMGtJ89fHhoHZRj7ffaVK7Jj/NZYFUZH
dHQcPM2YpVHGSQD/+QO+18Iaydgg/eUKHKu0xuVhWKg5tDBGwlMl5+NfmzpjkYxr
e/CMm3kBC2JwMHv/uCwk8Wr3sBDI1u8HTZNEFw+LuKk0r+zskAtfWj6A3o8i2LKU
3rPFVNm7O1YadTZiKUG9DhiGjMd5vWbMG9PCH5WQYnOOHxreuYObm/SNljYGU8aW
8dgpKmC+wOi5GxrlmAzub2jupMUuOUUN2T7HtWsYyYTzBVnoCaKpfIbB2Xb5R8/r
QQqdTBIdvXrpP9YEe44wihy6tsr3GqDAbpAZIUvHEe5bBBbx+tqYcE/B4e69cQcC
gviCHd7A/gKaW8DeAGJJKJxfofEOv7ybwYuHRvwIdidK1A0kNsflCv8pAP8QMmwA
cFdBBjpMzDJXjZktb4uMNL2SJGlspHGrgV8scLR818+vMn2zXcGGcY6VNBn95oT2
IQu2Qa1x/i/jgyll9m5O6uBcONhuUA5bfeMTTuE3eZjKSlGiB4niAxd+Js/blqUL
cQ7hm6Md1k2Own21d8NA8TjjmRQ0ZCk6FJ8eIS0iAUfFZgogMp//lwk7jY5yBPFj
nHjlAvYlbPkXRSAP7R6NHA8/QFFIcfuyvhzULOOUc6qXwDKf693z3TTHDquvm3G/
bS/p7rs+AM1vatrvxe/8OHzOPeDxNE0p8UZfeVQwaeo6zEuRQEUtD0eYFc6rzuVW
Qf/7on77q+4WcmLBISP0xSijDnXD8koZCOddDm3x3HSs18uUDCVqOKuzK7ro80T1
udmRUhViDyvfzj+pkfB7XhMSn7xQPExLWe4PJZ6SLJdxR3ivPA76Sqp3xaYgPAq8
ZOxIZQG70Jpa1TvuctA9q5SUMcLxEn2SeyYXtj/oz86C6RpOIjOFfUyw7GGPzR1h
4lrh8Jsw1bXH6YywaO2pptoNol3re1lq2ueh+TEDYGFTOadcHmKIEo5w+MqgMIHr
ocxXyg8TEfntByjrRdg0BMj7x87qhTSvglzLZBMvemCuV80DEwZJ3KfDcVcqjhZY
wH2f7xZWHvuVzSdDxYQux8wzpkgXS3TPv4Zt+TP8LJPJkMiaB3Aygi3Nk3uYZBf9
a74Lft0t9aJj1pav8sGQAAEm89TTwzJzMY02kqNYF9Muvh/iNeYQDfHuPa4vkQJ1
MQ0DqQWnbSx8C/XRGMsALjaN0XZtC0aTzFTIqj2axZtflBMDnZpGHZSgJWMRqKAw
TEFsWcC1tFx2eLg2ZoJ/w1r5ssFCBgIctmNAvtlmNdlIdetdaQ1812oSbqgI1fld
6SIxvjUuFgv0GNPrIqNolXezb3KzV14b3yeGjsn+MaAJXlUMNl62G6drXDal9LYh
9/toAgXd02XFbXj8VpO9Xj1V6LeshLgqBTb2xDon6CFhkIC2HIh5SgBr2rY6xO/s
VG3A36azSCeFX9YG/ogVSNkDZeVw35gUZLWDT4Z5b0JxUy0zKMJ3+3MsQk+Jl+Mw
Fe2xyq9r3kuU7uZ5lAW1KGTTGkNl8MJbkxtPASmFtYhZorLbeABJjN7ggEDKmqjj
qp8ZduOt566zfzA1hEV2Sf+Eo1Y9vzdpUxhQehEK5QxnhpDGP/g03hQcGb8ejRBS
psIWXp9dZNmQNQOc7RVAKmg9Vhfk0EYrLMNFhhgtl6abr6iN7Kb42C7r/c5RLw6z
g1V9OA6YlXQZjzz7B2RyeSZbpIpMMhKJiadyx0UkvcXOKLwDqdLuzynsjRMcezht
ygI+y1EcHUPz+IlUcmuLUwjeXp/+6SPOF7mG3qJr1YDD+d3LEYrU5+LRLoAWe49V
X4oXA5Ii3CuDjuQjA3mz3EIN4AdI7o5Iqn0/QUEbExXtlwjEtqMjWiCNtP0spuKR
0l4aSd8y2SrWHZYYyTow48/wukEgEOM/gSgEYlVi3C63sYkeA5gxUq4T84IhLc+J
FUxo7ucqYi99tb06BItg4Oj/KL26Lr0n3V91fBuczuPM83Myar32AYErhVeZmUj6
DuQvw5ud5nzklW33MVFqwqMPQkndHaby+fatzrGWcHPDQ8oBoVfXKzvubuBEySyI
+WLdw7930jiGTfIRORCHSE8bG8AIgo8zMzr/J1g43ir2pBEepeiuh9dLrn8rs1Ec
y3GS5UXN/gg+9eoX1tggaYcFBB7MLDNP6c1rQ35qdlpoU7hNPsziMR4uBI/BKvB1
BXy6fObQIoSjQ+vmGgdwf4g2ZbNR6rvtPWq3JHqE+GJ8MrlBDtCTd9gKslgbums5
ic9cwvtnf5RiU0mOc7bhO+WUkw4kWgnCQjpVF3vzrrYB2Fgla2iE3QAvU1XAFqFj
kNeEotewccVJ5aRolnIubuyULIbWpLqRDyyznvchmbFFCFT9akwefh6VfP+uLIFt
tTXOV1ss9c4WVxrvpyI23rgCQW+m4MH/DwKntIiAiL/GT+j+CioIg0WfsyfZeL+6
EVNqjB50G3salqDUHr1vjy86KgUm7Y9Env+bQNbN+nX7PF1nz2RzOWY1PeIIh23M
5WaHB4b+BI+gvQmp3O0uxd1seimZbqumqLHEZedw6uIXKCa1DeRg6M+rLXJZ+aaK
zvt87MfkJgp8nLRHPzRJZbL5BvSdsqO1CqNfsTNzK28GjiubjUzVtU8lfm5s2hi5
57PUgkXVjAj6tlQ4iqcmvNTOg1a2BtFb/G2Jl/IoYU3oi6L2TFwdeDwVMiyP29Jt
hJY8x9p26jeldyGxzl/qrcwbte4z/hq7/f0200K0a0IsQxH3x0NHP6evZaayTxt7
Ma2iq8VqvQhhhRUQwEOSCNDP8CxYVEOaOdp+H2tyA7AzCRsdYwIMztbDMzbW+iMx
S9QHMdGfX6sd1iJuo+iHAQ7s//+cROEWVSIWCKtjGX0zs9EuN/vG1OMy0mx5j3Eu
gfUqbnJa6ymQKTlF8rtK6SH8M/3S+1vK5z0Aw7Xf163xBTduD4z/KLClPsI+CNFZ
tqIDi43kjvl8S+w1JyUkZjyB6bZ8GRyL+NffImshuh95JX9KPj2/KGjALqJ1KsrI
jalBn+B2E2TNYjMPDMNaOAABbJFY9vE8eTvL6oMCgNDOfFxVYlIpomFmyvdrvsTd
91ZRNqM5ds3CY5y/H1ENFYDuX5fOw0584zAEyYm47eoiVQf/CIzugPY4MrnsrIe0
0woJ7j8LrGxH4mLonHdmzl/8z/N1ABjqUDDoM7tRiLSHOlBaf/E8mF/wEuVKeQfP
WARvKXeTc4nTLidAfxNP0juzZfyIJRiXN7ITrvahlh61bgPD8clzXTuGruYw6fII
b+iij/bHbndu5ulWvhPPVE1YSFXmTioh+oNwNZ047WORFM/8IVrJo4qEPOvzII+e
p9PCmnwIjLDmieZo2GVQSN16DBoEkrTpTRMaCCwWyUBwqI0f9PI/nXBXaQptnHh2
+v+eKhlhLmWQKxwVNziqg8Z1LbMGO23QbcfkebUc8HFs0G7ER4YW7ONOM+TNO+aO
v4bfsuOWpq/qi0IPG5AlGtO/+evHmy0/eD5aJjPxIxlaUwIa2Z7jIye9Qp9Itwir
AbrvqoXh5h6VXJ1mZUcDWbPI6DY6J4UsASBnZanuNRUYuP5Y4u8YDCxLJVENdHb0
9PX4AzBtnii3QYDBiRrnug/Zuhg8+LOL/UpdbBOPO+IRcbKFKd9CkOgwp4rlTh5M
DQFN8ZhjOjGJa4Fa10cXzLZyo/Mi6O2/8pVFeoEnH/xxdZ1U096kkOc07imI1EoT
YuZfuivoQV3+CZsjZ1tfbzjkuFXy0l06ACC7TEwS4qcVVpAhtg9Jxh+9iDrqgszA
+R8zBS0oahV4iX1pZ5/rs2JstV5xtNpWOoxgeh7+LvXdNGpyIB8raytU2FFQ6ufg
gPVdOiloZOYsaNzMjSJuA3i5tMnYTXdaV4pZ99kbDQxBXj1EqdtAokDJDmOCG+xz
fywqczeNKxY/TVBB3IlgdrL5d4ianZLt4HKgegbKP3RUgEy63OnSFp/gGhHGUBdZ
KtBzlCuKChv1icMRxfnLSjJYbSs+KWfiv0hBpDBzwvyAdUar9ECCJCPMBYPDSLup
BDZh5a7cSOq22olWr1h/o7sdzabAbH/hD66O0yTNYFvPkYzQV8NcaF+PBDVXugts
/NSeMY3Q+L/8FX8L3LrWOTyPZ1hwWLllPSv3uxAwuYC+AbCVS+6gwAJo/7Ih8dyQ
yrdu6R8eUdolxBM3sjc6DLd9tqpAjbHLEcqBHpsIBlfn2cZX2YD8hjWua/uuqy6X
4ps/b+XZo7RlCfAgWsASdwdLdcdBMHBOPdstwNLcDpztDM5+NW1s6YgwMBb8WGFI
Q9TeK7Qj2RlEInlys/SElbEBjy9NhdAnDlTR6UfHseouS/p57MSSU6brIzLLq8gG
Aqrywe1pIG6s+ou1yleTAVOhAukD2M7SjA03gTofvsmcaiS3PxSPrYm4Pr098oXG
xmOKQbQI7fdUVRurgDNsoTO8ws/1Vnw1PD5CzuKcAELDwnyO4R7AHD64ENFYJaWo
cUKxPDNW/BIdtIPEoBBTZeDvmVB/ROml988X5Y5PUHlsnDz0tVr8W1A2hkzPB8lv
U1IZZgtoIj6dU5q5KLBfRG8k4pZBH9uMXyrg/gEfyBJHT/sZyAEMwNgKxN72dvqN
ngvjx69mRvPu6Z24npfEPM5fsXT0vzG189CudKCxxF0UiD1TCptFDSbNDtN1KS6X
5fbtePUjkAIbsVfUGtZdalB1F+Z/06L8mSNBBsTJYrfKWRGcALDHeJVCS862NSSL
odaqhvg/qWkPDtaphXr4yUCsQlzmXTn45IgHkLF/2ONuZ4wTbkgHVMmgMkvHa9Dt
idLaL4Uy5EiPlTLRZ5JxEKGPIc/HmQC46XLYv0VsbUYxBcyfcrSej6I3bprE/wSz
Fxz9Anco2mMEKPdPpfhXGSocD927ARA2KFdH4SOExHvyIVTRwHoPmTLjU7skNvGp
lpSNVQ2yW2XmzO/EOmPBXAfQSHh0S4QYkAtrPdgHmrR2WjyqgSlpTS6UuwtjrOb0
EvBdauewf1TkmByxKeX+ETLnghzZctN1sPdSPUf8RgBO4zdrqYuXybpJgq8qbLu0
0Lbql1xIv4mArgvssL1M9xeX63Q5V8zhwujpzfu+wuMFZFbRDVvEOo0URU9vucYl
UGZ5L/D3teSKs/RY6zRR+mj8I928xsOfyYA+5pyIz5iCoAjeB4MHaYZdpC04jdXY
blFpCQ8DmrPHC0IFkavZD0w/UuoANVh5KZLbdmwYYUHYxTQKQjq3dDB/XDa06KW2
eY44XQq15PSHQ/0eQ8KRXvMSylcKncnvmtMKykXq3PaG5ZpWdYAHAgptKtmqndjM
t99J+ghjAiIkTMw6nsjpr1RdcGJ/h8me28PjreU+Dj6iZkHOMRLn6EnODnIC3816
isQdsAFk6xeaogOUB5H9SNDPhF95I1gkgmofEtGlvLNy9yQvJzPSCH56ySx7vAeg
eVuZ6n/dEA84KC4M+0wNKC0F6v8caKnr+c0FMujd9wSRMQykAeMJh3cDKpDY50Ov
PiLak++K6l7erqs1WRJxgJJ74H1XS5/m0H52yxXBoFp1wVipr7YEmnSvQWXgSa2o
wVo+gSLFjtMYzUeKZ3gkc4IGRnXyO/VaJbyJst9eSux3lpfhrSNRaYtZdlRaxSlG
wd/4+yiKnK6sQmInvmwEC2PTuXxNfhv+4kZnC4Y7abD59SvGQET9wr72bgT9JTQj
HfL8t6WsuOCoFL12TURXdD7NEUrY2gHnoGiIBoAiqbxS43DcLQYP6CNPj2dRB8pF
zhhU0lXEkO9+WAX6yNzE8/0AVhn+H+AIrtzuaQAqQd5UH6ATG8N8/G2iPO2gBujO
OGX9Kqix+x4SO7aKG8oAjdqJWaxjscKhaJy2NZsC9XR6sGak0dX443oJtZruzBWJ
zdeRKXcyU1U87SH5OCW0JyBdFdNWc72M3sadHFKF1mJLxSZIAtb6ODE66YC/yfmi
bwKLUizsLsYoS5C1voU1DVk+RL2gHGftBDaqCq+dTEbfxhMT92ia93t1vm3KmBQj
Bxd4E30Z53N4lrZdUDFqYvYISEBELvtrbXZ96Dwfd/JGSVCApV3XzJ6arMVzzPOh
mIp0fXYCjEeqcWcLnIslAhUFBxnIGKOHnzZWUj/OSUGF3dnQ0jRsUXtyyo25Pz6I
A7tgkdDMdnlWX3TXEwR47bdP8FRCfSar1kK5EQaIXuzQOV2nyVAXfPOArNvDQM+5
C56nXgkMsB7zKWWE91ltVx5yHiqZtNFdzAjfbVpPj9FSSlFjo2PUUSxfm0lpI/As
c9PCL3TED24hTunfUp+YpnlAfLtZS2sVUfV4B5cBbNBUkTyVQMk5R01pmGlhye7H
0E7OIxDfEiuQPZHV4zr438P0UIuATit5mBE6eAFV+Xe8vftR+9HzyIFyndlJRRgE
FH5jHzk0c7Z4ukm/bzezPEgw0nNxPh/5oGzvnD+fYWYCqf4hNRI0Akin9B5/qSz9
UeIJ1eoEO8Q5+fs1C3J4KVyxpGkVQ6SfGcTauJP5R+hQw84nPduTD/yKPm1zF0Ts
2scX8sUnXNMF0tWaaI9/F06yQlt6bmVO5En8r5pIS15YUwTvc/X5Mmn29WBHOF+d
ZvNMuOwCYYgHNSqJofdDo6KXFLExFzCP8dGrlXewuwV/+IaP29r3mfxh0ZA8bQ6P
+cyJZOyDkXaa9t/vnAOb5R3ntm8TipxCt9gxj5d7RH/n8YnisuwJHIeS47rmwPCQ
kXe7oa8IjKVahrcL+UQl6cK3LzjwRf8nO2c/b0sOgW5GThJUYrqYorgCurIHux7o
ZE1IFWS2uO9HTIHMbn6U0n4CETXpMmOtD3DqXH2MQe+XPPaSRWI0ShjtGhSQrC7c
+KImLYGPioLrGkla8RjfEqfMX0zVOcjPDR4pfj6vhnOfb7DMy0xwi+sAtgnAHvjV
jTFlC7CkX4RamytxtTsq9MDOkRa5TJZ4PmYyyjD/+kIIjt+A7qrjqf8CbS73+Qy1
vv9wHa/mLjqlQSsedyALvY6cnEUyzf4riau11H4IFZ2dEm4hBSHZTHgwspim7Owu
JxkJS+Y9RV0rhPmaPVuG7JM6KvxOcZa8BaWz0G1UakL6+qnBl/9WGlHtEf/0ubRw
1E132127ycW+FOPtPrLLRfyql6jUkR0dUTlLc8kzkPTdnu3dxvF0PJuwDc79g+9s
jZuRAMFuWvvws7d2O7ZLIUbK574SgEa1xG/+3MRrwUrxqDyQC4ev3r4S3Rs3CV9f
p/TDlaKXigCdY5JQmOoLLVw6MooD6szpYCwovrnGGIF4AEpc1pyNYabvojWcOCIh
3+in9+ioQQFSEa9uqj5HBlc3TMsZsygepuEiwWsb+PacLX4SScKzSAb8bb0Ln2Jf
aI+kcs8rUSYgz6Hu58rtqaloatqjXti1UwDEEVP2iUGP3Jm6HeMrtPH9rjlgKZOe
EJOe9cecdTeRPg5msylOxYXrPAYUz86vgfkdWMry2sQ02gIY7e1tGzjNSBw69c0F
ouHS4yDFaEJblQQ1lgyD46p9wIyZkAeUaf98WJwuaj5G/RhUg9ZQBY/Wup9p5vy8
gXkXNB5V2mo5ExScWNMr1aTwl9lvfuRAzo9RkaQcnoO4bAfAmdl66J2wtzj5x+zx
yMu49xns9rmth49j/XKyhQZnf9wRqAl+EhTPsLJXwcWrI8aRSzYU7Lup5XLTcTxx
hHWMzo2ZQFg/xCQfFGdQrLCZDoi5Df3VdLqCCdKlSa8bVnjos72godLqJoFNeCBk
DZatPCzS4JWni9ipy9eRxeouh9SMEbVObbc/GdtIDICw6ggk0nEotEMoeKMMxgiU
gyjgOCXZ2CEad7sQXZ+1Qico6YeMtqrfTTYwhnyzM6DFNponD+Jlm+1J0fRHtBYR
924MWlsmpp7Z0F6kFUMPczmUmv3A+yUAicFb8vKpNE2MxJo0zOUWUkofyGSNuY7x
cnCM2U4i1RWLM5DqUQ/VBAqDgCZTiqWk44l1cr8gqMfyPKLjh6qnpL7vPLup8OWN
EnEfhiN5KMewEPBbl9SmVLDSWf1QGaiTiBolSAYw1Q+JxYTDjh8gVM5B+rfzRzGX
d23/rde0iaXtU5J+BAd/Q+zMIsp19d0quVXSOLsCJBbycqvFfCyXf10FyDvHr0cL
lZiBbVjQaFUq2ToQR2lj1hqs8Uue4pMmxi9rcmwqH/s8240kjIvs2cIb7/b3qtp+
FSOPE1Ahw3SKvzKEOIcPal2fEXrhp+qAM86V+NNxQikEHNxJr6jQ8miMo4rkrFG4
sI0WR6Grb9BJ7srEz69G58nBB/VJMc2KDw85hFca+F9cusCrXbNEGjJYBK6tTdNV
bddzzdOYgBaz7PTCO4nI9kDmyq46vrzeTWeyO5C3XCW1MVQKgJq5aNtM38Oo8Ggj
d4M17PLz8vKXerUf6X6ov3ob/1hPH/+9XS1tvxkLcy7G9CI3AWbo0gzxj1iQb57/
gLGRKatdhea+/8SOfM25r20hw3iq/FPlr+ImhwQiyA5d41ap8+wXBX/Xt8FHbHAf
eKUcasB+qVA+uZ4TdblbfnJl7K4WcvJR3AAey56AcqXmyJoyEMsjsniIG8ys3+70
H6mGlWP0olYSfFoqorGD9gR8HWzDQ9XkMXQUi/yxyoZ92FaL7iJc4npL/U9IwMrS
BBx9eOnvBIeABubazMpZ4JYqlpHvW70lowZVt3T887e27e/9Ox90fleJAkI0bsp0
CH5bguy/LT56rJhyHyYzwT+BLDAxDad4v9O7GhV66WO1/OA2QFeI2/bFPupzO6E6
f0J+4CpAMgj7aySQPQHaT4HAid4LaskcrH9MyxCVm/OOftX5g0x0P04+DAcpt1sk
uODcyYBnoL6yzIFJrmZQ+fsm/t8HXHTuO9ALZ4hdmRhA9mIZ2ir1AADRKwx+VY/w
6ce/3mOMqbeGq9bdvFp6b55tGxT6kGhxVE4I3O0OjoGvAK73gNHa5RwnG3CywJf2
V1pltkwqnsMsJTqHiTpZZEJEdtxywSwRVHTUcD4zY7rLBYO4TSjUoprZ0I5tKG4U
g9wTENbkJLoG6tRNQ7VYudk5ijIePIa23mFtBwkxav9DcqHovrdXLY9v0Mr39Hdq
IEAp0nXFvgXIZxzRzXJEtaPbu6sFOW4sOuMn42olRf1rJSH1CKn/VkPI+JILDj21
0/rnfu6uFXABVrAPUXp7aoPxvDyQ2SViI1lS6cs4AHANtN7I3GX+v0s0XABD5kXK
Q0oP+00UK7weqSf7wQHcJCLHqubS0S1nddW+V1e1H8SZoZV8Uhj04VDSQgoaFJ67
BS7J83gOaZmmBqKtWRwfXYw7lOXuGbzhAIVDcclTfsLM2rlQ73eHSGL7ElbVLu++
P+I9a1N4NBRdIFC3M/v5C2EKisH954mldnNBDdIU5cTTWODC9PESNVTLPA/loZA2
hnUFnaK+OgwZzkbRFZs3xbf3W0pQs+ef76kxUqFB+3UDnihX2X3UlHvMIQMKuuWg
5K7WgMBd0+zxHtDpK6oAIxJ88Tqta68sajuhn/gXpottMuepV+tBhUY4YScBnlbA
vCr+dsRKGqz/G938loH1elWFw/qnzeqhhEfzSQPasa07oiTzxq5WoeZGhh5iNYFs
Vsxa/GhDxadycME9mY9o1go1hi9seXEWU0DoHgoRGtVHY2GBkGcbbr2uIua1QDdl
ULHVxtQLU2zXLBj62sIGC0apKSysGiih9tquFWHIuOZ4zrCrzoAWiQcTFq5KjWMC
sajgcw1/4YyQdpsGr9WtNCKdvUyFqj3uiepsv9DTPjlYfraiSaiaAwaXpcNV9HEO
U1wsGPXMgWWVerXZhpOt9nkjX9V4Q8YHulbeWCn0jMzhX5gNSOP3HOpThIEfswT/
BKfQj8kcL+dPYO9Or0O+MkgU3vjb6zvcQ7LXCGmms3MWoIOBb0hVOKC4eNSVtNNl
4AV7cHa1au1kaBiQgCzt26gH6OolWttkmKRat6sx58F6FrFMXt+6KqrrLSslK2kc
navwTo5YiAjk4xaBqNKvonxfc35rkp37wo/1JL5Ae85XgEDd9Sgapke/EyJH3Nfo
qCzDZV73y5LiW+lW4CeNWGAuniSqnOv5HhLg8yqTbZltddgTTq1p2JkKv30NPSlw
n4ZVnXXp71hQeiN4PZCtvMqrc85J+Qh+1WUvCEl+vrIUmwmRb4S5E1Cm48TX5LN9
OC3TJQQqH/PqjU3D7nsIv0EWpCEu9mmR2ioZl3Ui8vO+AxiHPwCDTWy5E+V0IeA6
i50f8FGHQBPEckBD2CtjSpVy39fC8/SZ7AIpeHlJR1sbLFe7KYlZ7dsQAa156sP9
iHM5YdJxCF/D68FyQHoTAUia0YRSh4DLjkrsicQEE/viLlzJJ384dDCQrbgfbfZp
XpNaZ2eNWArQCIhd/xI7Gtimvn06ogffaiK+gwUoTEe/Phqli1BWn2Uw9d4hJS95
xwoDT0zTkCS/I17NKGRr1JZbt5K2qtTtpqBMJxDDPvnHOktbKZUqmrhAV9wYVBM4
v/Enb7aBBgjX6/d/N0HdkL5TUmUq6rDB4L9/Rqj6LqRwDu/sFjHWEGu74UzKP7xV
ba8WqNiiiJAthq2ATuX0UmwKqtekzw/dnoelMOQ7cuCdc7rQtV4GrE6641pmZlmv
/X2Yu1nVKFrH29Sc9TYBrcAF8sqXlYFfw3acbpI6yclg3Ud+rdd1ma4R5Plml9g4
PMAQED1yWABDrEiSGRwMolpm/+RBK7wFX52SwcdXCon7gvVPx8Klo7tBzvcaCMmD
loi6L/E8k9Jn/PkLKWs6gZT3VOz9682mNVat+dYomJTFyaQ+smAjaRQNSOYqZtrj
AM2e/PA7nrHTQLmBto1yifS0DOidmhdFVi8cy6Wac593ip9nAWZufzkem8tGdGSe
HHLMgO+CmkVmJ7tTQClOtb9VWAQQ76gZ9kBY233NJyZ5VJdrgc3PGV0D0Rorleyf
S1D9h0Cx2o0oV3TDXbZ/RP8ayP938SbgfvvnDFev7ouvN4OkuDTsUvamVUb3HRbZ
QqjGGKfo7zlgDPgwN041ggR5uSqgLPGtjR2sQDve3Y/fZCGzn4Zs2k+FEIO38+9I
lMSH3hcbUe0HJ7eKDYCdOiUMhxgv/Rhk5crEmg6TVsKpRCggFwggEs2Q06xf1Ox2
PmED3Y/Qfn3hWiFkQDHAdDoLQGXbGBruCvIIR6GPvzVQxo5qjAXzUhjeTFQ9yj3U
Io4FtPc18jqj02QD8+KrRftYq8zu09YcdQnRdR+uYx9u4tGHdPp7eI3IskTNPnxJ
3GgS58k4xoIwl8tmhX01R92z0KyU41xPapetbR5IaL4rGQ9ySmT42zmVdayZtRA2
twANFWik68i0oOHtYevdHgc9MdeQPT3fYBzH+aw1UP+RbacTW9LKUosl5dZ81DMG
BX2ScAjmL2wJ7OLSkWR8PDWoclqrnjE4uXfxEteZeJmE7O519/pzeYrobM7XXhkR
wDz19QI0Uif20C0swXM0zQ1/ypJTa0y1EROx3C56LFID5USY1R8y9XVsKhB6d8xB
PoW/d0UFsyZZK5LugOmsHe/JVAIat+UqayOf0O+lZHMyLLuHBJWZLDZuYorCB4Hu
WrcajeMcP5D+mutT6PytD9B6Cl04HC6yIYjuEQS85M9A8sqfTUjx1DV3x+PkelXQ
+B+7u6+xO7CQ53mPCffsu0pVTGTK68C24VJ5UCorT4JS8sxSx0MVSYjAwWE6Uxoo
5TJQMCLwcQvtAhaexxWUfVET0pFvLP+i5+szloaBwAeqrQ4b190S6Koe8kW04f3t
ZxJAaC8pWLKf6bdPZU+ZG4217XAA862ccfoi6W0mL15AZo1Mzc+VsWxGyitHfLEL
nRnpCX32Juvz8tlzDgS5GwihSsFmlwwwZKXThUSqO6xAeWZwv/AKVavMT9BFaMPY
G6N/h2/zp4O+i1CzRNvydVdv1YnhLFOHRc5C3BWegZNKKDBBlThjcFHltXH/WUVz
1U2FXhRWNR8hQpadV8QlmCdXcPgW2J26MsMhaPjNE/x0ioqIyA2KBOblOMTMef6t
Sbefo9OIUv2n7ZcJtAV7vUHT6aWyOl2ZKd8derONj8kt+eeGSYZ0pQCs1xMXh4h1
wO6VQ3EiqetfiiTLUkOo2UV4fiIugrVgsMQtOnBxCF6awxRGZik7LdoA8JRORwvr
qDc0+N87iY5pWBItyBLIR9VNXNSWsNPcAe7wTDvO0saEc6tsU72LbmrEGLRpEcoL
BUApZWusd2AGQB8xmAVyo5etcsEq/L1ZlBuSeEh+0I9Ri9kioFJNgtg1wa6bPq4e
vUO/Z6KYWocqpTTMhEnV+Y3waGAeW2zuunRotDJ7Xacrf5/r3iMUHK+ePxMvBLfa
ks8NUz8L/sbvuX3zS87wgKRKdkLBHP/Jb/UXCE84FS9b7RIfz7sLk+8Qu49BdlyA
nJHznkgtTngR/eOIj5K1atRuKlEOKDRcpEOPeXjkheFgGMA773TX5DSc22vUq1G8
PRA4vLRgzioQghQs0TIjfqK6fBgQ1oGlIpgaBnq6QV83Tf1nWRz1GJnZdXSZAh2v
o72Sdv+I+UQctA4hsutS6mLEbgFUgwd+hW2ES9gTEqUh6XlmrAaSeTYHXzFsoEcB
14gaR7HgOiSvA4ijEMxcdrAFtSGq2Iv2LyR2dRDTiHu/vcKUzHalNJM2jLOgfC7A
IFjTJln2IvDy8zVMdi8bLqBukurl2FFw2l0BtZiAxIAtrRhHUIUSKXpIG3lkDhQE
HAtEm6l0RXA7CvMxnOrXSBpsJIgU2Z8oiqyY3l2Rc+7XSI/G7qQP6HQbdtGubVs5
sWCW0AK5kHYsPK6NXKcBTDtLU+qfUNqW/jrSogHEBoug1dhTLIM9izwwGur+Zfu7
Xcx34NKxbiGQj4Ms3+X4kKJ+KMKPLh44AvTwsXT3E+8WnFd1FHvgvYWH8FyQq2Fg
ZHF5zFF1/BBzTeRajdyYqV4rNbx/gNQCRe16M/w3YhfrHuJRgi5PgTD/x8boOJBU
OvPqF7Es9PR3+EsAliPpUpwcgTkPfP0O9XKpw6E1rPGl//MGRQF5hkf5WjXM6sF1
j/pMe6agI/d2fU5F90iOX2oRuhVJiypRnaSd6j3KzuZsRo3s9gkio3ugQklU2xIA
dBi3mxwpP2ClpGfMxMGvXVeBr6XemjFZSc0t7OZ/WTlmpqbrLnkkm3DxmXRvotSh
0P6f49ofdw5yLQlX4x2kSfl4fjqnOTSQGdaH0msP1KoqteL160e/Vy09NLivjhHg
ZSlBwJcQL7bCG0rdcjvBiq3rtghf89WFl35zt7yz4kc38gvEUGfkLjkM9bgKks7Y
4Ye0sZtk7UsLe49jnXeTHRVlXFwkWIcsU6xtlMoHS7PpsSp+ebh64TDWofRgFlw4
cyvTNZTtnRowAF48N0ljr269FFY6DdPp0trD1TMK4CEOuqJxOgGpFLk0kPX+w4Ms
/ucEJK0BwRsaOTe6WLOiRLCQFeE592s+iSmb7awhlz/YtjxNbNTr2rzCTdhkvTlt
iqIvllV51CI2+2nrvQZxGPnDaniWtrlik99Ux7IczvRc3yBKOme+vNUvLOv86Dsk
nZvUsK20OxmvwOa3fPdqDzy5HfT3FE18VxvMZV7h5rIkET1Pq3fe7YoonXe82P+a
Aa0EeR5jwWeWyJeul4TXjxBb69zykZGRgIfdMF2bPtIn4ZegOq3n8R7D3QtL1Frv
AmL6zlOa81rrAYSUIy+jPOuWrIvBq1j6OUby1oNs/bqztaVLSNpqzh9SBfDOCDc/
ljUOXpc/YbcPnE1Su6ft/TaY8uJJV3Z+nnDr06HHLzWmy9J/D5XGCbNeP0oIAkOH
RfA0WCs/o/hhRSMfmqghCIDeJW5RpNHhmZxbf/gWS++IZGsAIR0HsqE3fS7pPwZ4
Ghfw/7BIa1vUsb0sY6UB2ZAPPEYV+ffmQTd/mB8jfOLzrC47Qj1OB7bf+9SUyWMR
4qGIj2Fa/91p1DTQuGC/M8Bn29wEr1fTVE+zIbKhUq5s+bLBesD4trWsuJHYxdmc
Y+tWD6v7s3JCuEKGzjMkXJzZ+KiqJa59dss7gy6WLlEXjxJfLanCCLL/GIyHA/S+
I1scUCIdhd/FA/1Z46U4uWU2JR7Nw4oFXpHkUbNsrWz7r5zogZzkSA78b3Ff/SV6
5EbLYLV1T95E1Q+bZxF4CJYUOF4Z8AZQw8jzxxri+Co7OaxAmQ5frgylJCRhYUHk
xunUiKtMlkKDrpAUPFTuMxsKiclGQUwCttviChZjrWeO4+mX+8NPdcqP1NexFOIE
gxkrTR0oA3KVm12P3ES+/z/ENv66WbtTeYbQn1AZd82AwD7Rc3mTv++ZpyyXyIhb
Jvi7DIHwAqWoJc1eK1+/LZp/2bcOBNbSCyRTBmSa26MrHdN1Al9J3t/Bzcbc7nvT
7aEWLyvycVQmXDFE0o03s2H1kH2lJQ0hm7/+MJxlB1M1YmGrDF7Kr1QETWp1twTT
CRFVFaZb4XxvusQH2zMsrd8xl9fKdYdpMios3SbfQX1gccrH23JFznNa9fdHrr26
rQxuAv8+G9zQXfUX8mis6yoyn+jy5gjz5GcrX+sth9BoGUvpjQOQB31D7RwZSE/5
ZVYuYPfufP2twzgaGya/xt47duKfBN+RsndeEfbtyYgrwMg1gRUBkpWO+qBugUio
pdUc46zKnLHT5GMk746JfJM1MtFJxz6bZTZyoKAcPEa2Tc/GM2dRVAqJs6Vzv9Lz
DB5szvOLmzS1gZt0RB+1NsS/iLIZPKxpXriXfM1acJ1qAwHFxzkizPDDHFUDXS7t
JR2wkyWDu550y3NgKILNBT5q/TctglldSBmKzEm6mtuHXMgHOrY5Lu5VU/pbPEgb
MZiF+okYD1lM74G1C5LvqIa9sbdt9yxV8IRjFcq2SeT9cAXG2OuBb2xx0SdPO8aC
V86CrCQ3bk2wbqgCzO8oYB7moI5xep8v/ed3RuaGpy3AAiljqp9yJ4xOvsnSTlLb
W1najPKyO7dQPCykgJhyWvtidN/wQznVgzfNXGyCtLyUcs4xFhxknxOYs8GsiJ9D
HF/mvqUa5jw5pxwdRpOpUGo0Wg7gba1iFw/kaHRjDew++JStMGlVV8laclW2h9ka
3JNLpCvgTbCZOl9GjuPea65xSmUYEvkvzGX7APYiOLYRzn9SM7CUj1TkmoQ/up38
7ZXcDY0CuFld8PWbRYo7bUc9LrKNBpSYXstNHbgEf9f4OwfrspBn4zKCiK+PPqcC
m7s1VTYeL4/whFhXQBp4Em78m94TzFsDGiJk+EJK8kBDD4GYcA38AxmsUBRTnQBq
8PkBV0nfxUEpRMfU+fbawR6ytDWAwbDa5nz7d2+cpnx70D3LNyqXBKxE1Xw0VUxj
DaE7lVEf276WmY4dk4aL+pNC2k3croeJYnZUqNTAHXyppWp2OnTC/kNY8fbEkzwu
f5DjgcvyJC1HYBcNolvWltP7qtT3ivSMBFv87d334nvcJLTz72h41PpeCGsXzcUq
ML/nqZ7KX6X/04HcPqmbwmHvlY0rpETGWydEOJLNtX9xgzDiaI1n7petFj7feU9E
UO3XCixalT5LrJrIbZMlHWqi5j1anjbGCj8KQQo4kiBqi8GvoIRr8tLgdZ9dzXAP
4i9LQy+g3TpsgeO4voD+BYeUkDk2pau0fjcp2EWdDxnymKYEUCtKkqfIRtp9cROZ
uNSZ2SXIu+alHgABWCPFbVS9Jp98cN5F0yABas+fPUDvMJDqp5+zFsorAW43j47m
8BVZiTrQk6fX4P5o642zGDHAqdA9ysVfJHTNslV5+409z4bF1xaknpidlPkAAHrI
RhIQtHlvkm379W1AVU0LkNRiYg9zvN37+voEhXzo14KNBrFeBmre15hBclO18/F9
v19LN6uQ+OBap5q/h19n+XHc/Bxs/TUHbk6S68oYbeye2zISSKCumu2I+BJxk3sH
axLAhZmZG+reiKY3FA9q6y0YRrCuNPuJf+wS6+B6MK53tVPp1ANLwnrT62hy3JbM
ifSwRCq7wdmZidNwjzruCNizPExb3262Bezx48SietnT2BMQ+Sy3KGGEuuZ03NYD
EdXBTknO0XdJ5MNOMXdneiOmQJjvZNRkhtc1mF9QNCig6z07TD7JRh+71S4DkeHw
wXC/ddGuM0Be00CofTBJbORylAqJd++gXkf2tK7B6s0F3dxdNQ19KSWi36s5kho2
MT9qYzs9F9IRQQVaTtZ0JlWw9vvVdwVmSoKN/KPHfj4f8Q67aTZdmTPt3GUoc+xU
g4LPE8zTVuPoBLGuyBqwjiOs7C9NhgT9lBpTS1MF7nwy/7H0PMbUGsDl5d/FiCsj
E6F+eDFbaYTgqu9RzqPXdxqsXtTkDYhoam1qlRtkjzW93pOpPm1s1hwCH5joY799
UmgLHsCP9eLAHQLd7kuUcQlldLjXi62inUj+TeHY7vVVVReAS/mpWX6NUSZa49pd
xUibJQevrTysOurkNcIp4UwZVwWvZN8DePmO+gbtGyMixgEgGVj2KYB4j0gVqxdQ
fUYHwKFfwLMuWdbUEC2djqiQrrWXAV5gA8H/wNdMkqI6GrHu76T9GzU3No47RGbP
9g3zHNRl17yeMn/aFhoIqwPflTjjIakQb7mtxI4R6lzOMe/3WZy3cQoTtp2XmmG5
9O5amxO8E72lF4NpdxhJjAd0LQAbtyhevZcc0neTwDjqWmL8LCp+ewm9Szjae1Me
6nKE3WNlFEelynHg428Nlo1rcUzLqqoHSXvdeM0XuJxJDOw3XfK2gwqqiOTemxGV
Wv/A6zNZrTk4JYqKnLPDRPhLf9C68jZ9wxcFxq8sJgTZ4RPquZpMItdcIMpv1Jo2
kJu5fCrKtfpHpjP/iwrSgj1jxefhB9Y4zX4dT+vIQAgNeQGy4lU+QxAEPLbKgSCV
zqBkw65z5WpqgmVagsFRnsqprc4ycLH65PPccXZoNBrnFl9nruER8iP5hz6hcTHn
btvqsNxZaxJP8nLRpHaqtQj4FEUy5DQhF30Xj0uX7iyudSPCRkoGGiAjLWrbk0DD
oavDxnF5g9OpbbXXEgrBzOmTPEEQC82ImLROMAxvMYtsdRZYxepNDocv3AO+uicN
MRQUouytzfrpgAlma3VHCcO9I46euEX0b2T37QT8pkIK6E84iB7ggQNNtdfiEMyt
0gp6DA1RCyU2OJceJ0CP0YWFcdAkNyhhZKCm0Z6VcylAsjvqocaEAaBGhytgtDzZ
Tp5T+IUiwd9KcFAqNAgYLIazb5qr+nIYB8axppVlo+luRy30TB/zV9hrCU1otiwh
X+NPv/pVnVbBI3IXqMiktS2FcBT1pqJYlXfMV0o/v08A+np5XCQzLK+czGAaSylA
qnADCVwFrL/Wb5w9zVuIu8HeXu791gosqzU6YYACfyFR70G0AFkyWupyqS/FiHL2
ncj5f5MqmFNClzKsa8j9qERJZU+4qC+hrIsqj7jwfHS154rL0pXja7Egp2PKaV+h
JTOPkBFZT9ZPQ+h9U1XBHgVdQz0Pwn1jgbbnqB1yl6qDkUphVQjLd+pcDdoNSSzy
/p/mPK+qikHr8yjVl51NifETAfyskmCK/wcFTme7D2eDyKU9oerHp5bX05JFCnYu
9a9MqJQ5Zk9/vQLaZIJ1/4WK5f3M2lni/aDkZLG1720aiVZQOtivfVaBMZOdLzeU
geIhT51B8Q2ZZxRIXBo67zHOl8xOFr9nV1JcxoI+xKBjf5JGuMReLWojj3hM7LYE
gzbGnMs/ThDuBpaph7Y9alkfsEtbDOcKRgAJyruxcvXqJ4CRIuhrZeZEHWChr6+/
HXRXt/1BVOKp24nzixEnm5NkZEg1HChi5lZA7QrPxpsw5OODhZQpoQRbFv0ImeNV
k20oPY+UCNE0gH5ILfBmFB3K6RptQiQyskI1wOJKT7xM/kuA/6ZdoywBn1xiqxLu
WxJu7vlpcAfGZwOK4JPxbbOTBO2nWStf1jzmSO9erbVUbdJc43y4aesS50MvNMp/
RicXXivIW+LHpTou9mTYUns7UE6IWLLT3rCB6Me9V/jXSjIxG2sB20zkmSFWCF4p
sYpEt25lFcIe5QBUT8jUJcXHktTu1nkN7bdZKS4X073pA3SV03HesXEN+TVr+Kou
kMNPcHtypKDqfLP7lMkVH4eIaRclG8IMlyr9FoPQUH649itT1FbqsR+cXJu3WOlk
HBiHld/WG2NpkaygMBIZGy+bCI1z/Q9k/hBCb7VxKP6inTpdsaGNqqmatRPQQk0i
LgFHE3dTRMt09vuTUXz3w6iXO6CMQomk7kmskhGZi7hxswr7QIRD4Hnz1htc6+0l
v0a86nsIootfOsGfa9PrwUcSHytEVAzBcnql1rAVHxvbOC7l9nHSLAiRmFkwZBxf
TjM9KnUzcdJmyHRMFRQ2cAVLdglREaybjJG/o8pyUQtu2NRQZriu3N3uXfkJrm+Z
37Slu0ed3TXrIVqAgyO3qxmT1rdKy4zqkhwvu46HnPhmZk4cHBiUHvpOnVC10G5V
qa9HoRTu1MnBqkC5V9QgCj6m7UvUwjoKToPvqhz/kP4AWSI1MGtdzuuIpUrLK9Xf
Yw6G6gdBRTcmo998XhPioIJSbgxqGXvPP5jPr6jWeCjd15sRWAIqC6m7bm8q2lnC
ZwsgDzTikdOk18aXVp7E+Mowa9t7isacD26JWUtcTEss0uvwHco+U4CByzIpxROC
N21QgEhrcDsES4Kt69Hr2RXz6ZAOWnbsR1T8SyJkSwcquyIdRft1RL8NhVOUBj3w
RYpC2tQBMEfsTf6kbu74Z89EweIvptmn+GMfuRofetLLNuyPw1dXxUFw5gorRyXY
O/8KYx50+WX0aDsagsIeFTemo6olqEAmkjk/3L1/jyRpeyPzfRi9fnchOvvrRG8y
Oi5BE5clAxO3BXOiL74d/R8KF1dwMVv7I61tAbDwv4Ny9Icfy5pYSGT+TAY6bRIN
kpWhax6uAj8ODn+uJktCrlWhRJ5/cP/pjtEhVL/mnBxsS2MaiEE8xUcCVbQZdQcz
M3llGNal/XqMApH0MulJslUew23z2z8EuE4ImULYsAyodBDdQ+kb7fGle62wyXEK
PS81IhCCEjZ2NlLi851SjBo8WM8DBAmJWBbaiMIDsZ6BB+KO/Sx2z+/RLtw3xqi1
8nCNEaweu0iNXVg8BsUxxPBneBBX67ROkIQHcKg0VmStqYxiI3Ep/XiaxVQyHbKC
BVvVj0XAYWU9dm761+4WuwDhIH6bdPh3yiU4/erPeib5uLEYb9c8XHnoumTm4c4m
fzqD55oR818MO5zO1TZaD2faDgXO9cdt7zD4uq1n77fXX1tAN7F1j+fwj/rScg39
wEJFrGbjYo+B+cftAWuLZvoNL95Vbef1AxY07uQ6P9c1B4dfwv4Dz3/ViXGUULM6
7J3l03K9zEpGdgbPhErXWg5xeUO+jV9jeliNhz5wzGtDHyXFynpLr0UM4QqifyL8
hflNMjXr9lv1JDxGN4Rf5tsLXj/OrkWYbu9oJt3ioU6m6FSt2AYgPt7w2hbav2mK
CTiQB0AO6ZXLGnLCGxh3NYldIY1ok0usf/ZVrGx5wUpt8qdiOrQmE09+bzKRmhUJ
upG0En5k0Cm4U2p3Umj7aHBv4pQXUZ6bE+W4qjEisJ7nA+YOScM61f7lxliUsY6Y
6J+aGUEBLYLsn1EibIgWLGyfzBhPr4mCt0BnyuU5FmVZawr1VSzQ4rcPHx18E/kP
4ki+SuWkHP1kGAfHbFss25U3GZWk3CNa3WYg3SdWWMLQ0QdMaEEWzPNEU2PFDmY8
5va/D1+n6OgqAbq+RGjR5yoUhHr5HwqtKWDknFNGwUNKZICv260sVm1OnQ4X7KZ7
I4BsD/ym//M9/93VTh/plktdwvPoFAgeqzhj1uNHJI4vr6BjK9IcVteJ5NtasfMM
tEvGi68hHayCNC51/zX31//Oe3WI5MkbrdB3ZwFi5LppDNQzfyUAxSzNEJbXlWAc
ri3HUFuVkx8cjI0LZ9/7C8ykMcjFVlmzSnAXN3/ZQf8ou5JSvh4ci0ApajIOwLAa
Eo1CY4dEWaZMXX4YW08e+M68Cbkb5Nno/OtESQxE5oJRFSxbvqXGkXJQWrBcoxP3
W3U/szjrBOgFPvHI7066lFXaQxS6Cm/+8cSS9J24fOFai7F9F34xi0/3VboyqcHW
YcFfwgD61b9sukuE3hwHjmO6sAHiZrYOdn2wjoT9aWTAZuyPPA2cR4l+pFJ9tWRr
XDnXC12BxYZMyEh3JTg5CTid33Wy4AQ8RQAZA/vKms4dJgHY1aQ+Bynd913yqGtw
JWrnYsZZ7hlastAMqrsOAh+V09LYE4n16OkWoO5Mxif13TA2b98nL2PL1P8LRWlv
KVCeZGwJZdvnsu9gPbGl7NbbZhWXE+7kgHk3HRpw6cZwVMWU8Iy+VAA6mZuhpYpM
bM9rj6uczZ0qOaAcg6c40Vc9VYwOIyHjKHZNFK5bXA+I7Fl00ex3QRoogoeCakAF
mFyEuUa8QZkwn6oRa699G4gNHaDYasbM4KdPzPDdmeVnL9G5D84iGennc5ADMhJ8
fV/6aRu8y7b1C4K9uRtizyK/G+Fm13rLT/5j1/Z3ews9Zw2SMvMOgbHH9zltMpMg
RDgs13JnOUdHkrwZlQpSJNljM2tlkjUFAg2LiS6pyFaEF/XuNOpmFdVt5G+tRam0
Qls7FSKLcmNI9HQcdu5YO0PvE36m+XWUZkXFSLmXKNfeECD19QGI6fq23QX7bEWf
Z/W+7oFlMpsZtfgOx8l1imQaQ7+58UvFO/7tPKX4RdmPAX2irNJ05fXsC8WOHPjx
4HwecZFZR5TRLxdqck9CES3JkayHXKhE1dZ+AD6ZwKz5V8ZSg05IrN4StFWn6fpT
l56aRMY3weNLgom4UtY2iuC1wNkXGnFzQwApgL1etzeHBQq+Wuzp9D2jytzNoS8Q
kDPbDdvlkH3f58YPR1rsq99uNuODi3+572oiMUh96rFM/g1jj5vac4znf/pb80xv
BoZHR+vidoAr/oFbHb+o1rrITaq3TDQ2TTrqlhkTSH4ig9jI9Wx46+DOKkbwoqBx
5cd/c0n96JJjXvvGbYdvOG1DrElJSfvHaq1APXP3NF6X8nM90pWQwwdVUpgXRB3W
nLAfOFHG23ltcWeyQkuFxbK1Gk63lN18vPsmuPzn7XHFNtslIOzBXCQhNeC103UL
NgDBsOGD1NYDQd4jv7dsr8Ot9YuTW9FklGShBXCm6VLAd4c41Z83vnCM+ecwZqst
8GFnVtsszERjxPTQUDzGcndT+JfeMgfStr7kzvGje52BKZVsN1bbV7/gP9e99/Lc
UwAjJm3O6zwe4o9HXp9yxCUBQ66OQKlIR6Dg2mGTCpZhMaTaD0r11BixzGLO2Lrt
65rOYn4VnH5yVYsOV8KsaeO8OE6vvqCh3PNlr2FCvJZpGqDOP0YHkG9QQpodaHnC
Q+k9UZTby7HTD57A4CXC5bhZ6k+CL7Ne9CcbFFOkbO45k3VRCglj3tp61rbkMlpz
zcjDLz069AEblxsov4fHft1UEeoZDVsljhjhecD7oDuIxjyGKChY3XuURzxpf4TL
7NfPwliX+YtUNV1SrsYWMzuJvXx0DyyyG57wewC9us4I2MHTf7fINYu9oA9O7L9v
jPgHZ18qfsxeicLYi21ULlxbLPirt2IooNRdX/waiu4ygC3/eso/Zo92ybr0Rtf5
D7EbInIeN+vyf3xOzWeoam2msc5ez+Fd0CHCrc7cB+rT0F5aXikcZs57tP5sE98x
NvhPn8uN3ellhDZIA6k31ZSOn2boH3baBgrgMVmDkmSG/b/SZMT2xvjoPv6nCeqW
yVbWHNZGxQh/y+Tq4o/0r7iYDOdLAWk3myhz+PTTVGJvoFLAcJTORLkdbBcBFFyJ
NELcTYa5JqqZrnYEPnOcTV80vsDuF2sFQ8vPPDC0CvETcOZIRIh2uw/BZkAwTwyn
KGUSAyxqZQXQ5jR6LEMgeL9JzDk7Iz3y09f96v/0bb7LR66v+6YsQR6qnvKAFwwE
5bag2HJV/5ubuD/1vBCwwsmFdprkEdfEPk7C+QjYKdhq+x2+3BjTRIkU94RnBD+B
2fQuX8dbDdpKiVH2e2uFe6fJMtAdEs4FMoPf0+N5D1UyomWKauaFdVDjS/20CBcB
SRP4dzoKTh8Yh2h/1GjhvIxgxhFlgKzw9r6wOX9hSDDbrZmBLr+uYSZVwdowriJR
hsWZQo9wQ6sAn60EU3wYN6Dt0QzIlN08Ez9+KVseHkHEST4/H9kcwF9jmoLa8sR8
zRbwTyhLVhUBDe9qLBvlfaGdnLdOqEqRz3i83sRYot1A1SK8cOW2zKfBQ0OxFcFJ
DQxUBhkz/XLVuaqotwabjZzxS0jhS29om0N5a63nrQpAhCVL2BWwzL8VkH02URpF
QzL+HoTHJnFFvMMt6ryJ6CbN54oh+8rl5JfREbbb6O7PVQBzrlMWVULnei+OCcb5
T6pxPqcQ2A3PT+LEaAeBOEMNjiHqZ+BrpyFbqW72IJDV3H5J+jJYqHWUHx1TJ1sb
yNXngyXQI90XZhFMQfiTjw1fIrGjr4l/UyYPzLv0Q+qr3UpZh9QI/QPbDM3Ao0j0
Aq5rvYZduyNPePpcAAJnkIreCNX/d1q+9zH1Z9gGg13L9592X1DH0e4arInhGLIO
DB+ahuCQFnczpK+1kx/9UwIyVlTMdqoL2MfDFDkDrjxurESEW4HHRcnGtW/J35Gk
eKicSKVVeu5+5blpsm5WGR61CdnaGXZSbI6dEyPvqLrr9/0eQIs3uhEbI9TQbn0h
WXWENbQcWvH+jq4BQd1sm4JooiFUZlErQCnjlMH2zBZ3cmH52r+zF/aezpA/hPG6
vm6+/Ln7/HCse5EKK/QcJh9ozfk1fXf+MhV6DuSCbA7li0SO4klmMWtHckA+ttA/
ajzkSPZARVqqusTd2KEnY6YkSMNBbewJVLqBsjTH2Mwh60DzcNSakXPNfJtxGkbN
MYncbf4vRFB3gy+rHTcAYPOPPwUXnyiFVbTzpZ/GEIWQWHJJykfC4o0b4ULO8qni
VdZwoLjqtYMMGvblCwU9EE0eonGfHnErQU96qmL69MITTwYSxUTt0s5fYfe8z0Ga
IKalJjHPzyRGfylseNgGLO2XRJGVqxiKJkOVCzPPe918dGau07oiZHmaYM+kVAqR
TRbFoJys4c9OdGFmwZglRj0UNFNlEFCKWVYd+x8v9jurJzyEY7bsq1hmqbjyZ04J
VEh/U6JEC/oE+t8Zb3+JWeCGpHIlESjz/8KD/yWqENmt0GDqs3IRjDopFzEyvXIc
Ul0ZVNKaaPKGuL5Hs6G9JWjuYWM+XG0CEHnn1a0LNc/3xglY2o6Hn06SYq2mcWYa
53RRq7PMggVclzofrjUDHjEIymSzE0KqOcNWLSIKHXt7gtmnOE64L0eLPkNQ4Rgb
SXItlzgAS0ykIezizBWJC24pD6RATTYHDpYxVD6iDSXu5CXzfbR1woOjELFuy4fd
AZw6O+RK5o9bg9iIeWVn+/1ymuZdTT0lCXEAJ1acyQNGKRO0GmGdg0Afista5e4I
exzFqj4SoXF+rq1RRD+eHCHSbGINAhHmR39JQk770rJN2+S/P+Xpwg9AO+kn0p2H
WV/kk6X1q4J5VA2HHGiY5TSsSYizx8GU+0+q+Le385VDwkJh7L0Z34BMy66GEMBL
pckkftQOOAS6w+2Qkky/CIr25wb+7uYPxNkd4GbzaPEX4+plgS40Ouy+CvZjv6P1
Il5JO2NKDkKN+SyISTfVNd1A1WNT8G4mOhVut+Sdhw1O621rPNiLw9yxBR4Si5dC
4/wY5rS3Bmbum9YjNiAwk4vsPY67PgIYpSux7uWaCFZg81lOOb8yLPgeHxMTmhSz
kKBpltTqEnYd2AJcWaLyqTdwFVXXw2/aZ5SZ83R4+I9PDbXJT+Jcowx6UgaCdtko
RpwcMvWITWWJteuoRxMfNh6gToVVkpvdRvcYhnMMazk/uRViWdFoVjocrrLebUmX
ycYx5zUfUoZiw9rc+wf2NTFuPp/XyWSCj+j1fIB6btBCkapQKBfxxlmWoaSD13GK
UvuAkmhYGUd+/PJR0nxXYlP+0WnABRkhCtqLJtlMjca17biQhr/IcbwRocxDD4zE
QsAOsBUUOSFjHODx246LlpWrHL4PBjEe71GCApmbmsjbhWYmyVSTzd3DR8brZol6
FxRJsedA/w7YkhJqgK0MqfGzMcKWKO/Mfsmld4KZRIb/BXU1rQLKdhZWvRIQsR2C
/fRnq4V+8IAFkNuH5WDeRfQcSWlgA6rSb6ApAyPudvw/DS0nU0OI6D1NitqUTyvm
HzP3ubUNuFkGCN5BtoDP635UGZFHigiAiJ8q6v3Qf/eskxbJohcpC94eFYtNkuMD
7/6FEJmPLfIpc3BBAWGymNDmuaUaUwrLn7mWq2ovABOJ8abI2zbLYifdjwSrTzvC
cu0k0xY3sZ9Az8Wv8UxykhjWhAMjIMaZrSP+A669wJNkQrBAukF9nHQGp644njvB
JN9tshGftpYdVl1CFL4MPjv6NEk4gf7AFV5YJxOOPSygFh3QuzlT3OchcPQwiFA+
CAd0gfPT2sc8s6vKpxG3PqlQ2QjMCHrJmbCkfKIxWm5phUx1B6v++HbQXxY29fvc
VNEMeCYORadsymdWPmAaiJeB4YKw3qeKOIBUX12bCGQhUYqz1ANIlnlx+0qiajWT
WzJbYb8Zou/ZM5oqOrRO0uPWmJtT4GugWJgGstet19LtaiIN1pPmK3JZ5scfPo54
OVeICIsFsX10vLPqfvE06d22LrU1UPYxOE3LdVd44V1d5NR7bKIqnAz5O7/FNK1v
0Wqj+U+MM1zAnGXvkwK5RDsS2PG1wgABhIfP9YcDNN1X0Fl+uvbM4ILCBcjhDJDJ
/6UJUXQKXBMPPP14L9/pARPHU8K64aOjtA4kCe5g7aw1z2pTnGBaFy3yIDGEW6y9
/E9eupXgTI8Q8o433lhJMddDDP5wURJJ+Sx93nJDVoT9zlyeMey/iYkaYyHzX/wt
upRs0bKyO8WZEb4Q7BIbdvK2tfUHdmSohaCsuCt5ATYczYFpyu+dRRL9f0xSti/O
nvHMC2uicSnwcgAagI3q0ZyZeown95ePFqYNOsFbCugBy9YyQXKZhfF1bA8b0/8r
vuOdqMi0fJ9UYgdac3aMC4JhlwUaa8H4h6NdnBszlk6qdR6PuAhA7OQB+6gBzWRT
K/KCY308BMfQHM18t359HGB67iWXFRd9bUFxAg/RXA3I9LfDDlRiIxvE9lfOvFA9
rwEKeu28b1y6arZJ++PUOeDkzjREatSZ5zO1kl1+7Hy/qF9sjPccZPVn5lZ8Oelr
KpO/h8BVXUageqi8gHKRze6HxXhcNrPAI43L43UPLXGKsMXc//U8V8lbcI4CkTnq
iEqROK5ADyozWAZJcW26WBpOify6SHCEM1CI6u8DWLKgkMVhAoeqgCVRa/tz4Uih
lA2u9NN1ElHH0gA15cwMVb+mn4HsiRHDjhMToC0u6PN3QAYGGrElx3j0rncz+zIE
I6UrrqJZKP9UifZHb2GaM7wD1V8EOHLEvfwiezH01121fks9U/NYe6hLOv5A8dmt
+znsmDMae+cnWSfiHi1M8PXZyV00SptdB+BgYcwDJn3cWO+CfTOL39gHEunIw23k
SCwWdaKCaT/UIHVQ1GIA3vzDax+ZpNr7xt7jR5ufoB8z1axRA1B/d9Ah+FxgMcMs
0R1gaBwwo61v9jxnXjwzKXyYKZNG76cDlyrCR7fmIkjEGVM55ICOlacA5u1utMp4
sC/yb9yBnY0Z26OVMUAAQr63ktFv+nwqSzhURNk6u9nLibjDv8GWzu2Kerpy3iIY
yZIaesV8vG0iyhP6zOrJap+cvBLSGOgyiUEvmsXKTXm03nCM/s0Ur77lsrCUtWl8
LRWzPa7zkXzhZUjAXXv2EvGwm1Tut60/A0KSfcm3XsLcI2w+QnihY82HEJX4GxAG
rQEWyWstzH+ibvk2wfGp4c3KbYdd8+HSkPfv5HVTYf0C5xcI6/RnW0e12X+ej9IG
m47qhEqEElBp9Urg3UoVZkNSL9eNHrcoHlsWZ66nq7c0PIRrFShY2T3oMHbTAYkx
0dkKUQ3jU9zKv4lb8io9cA8a52sbvPbz7Rn9HNndF2Bh6qyNOdiK9XJkXkOFS7fR
GN7v5L5GBAnvOVSFAv7EBIbo5PxuhjsJ8PnZ08198VZFb1FrGBgY+dDbXRoN9tAk
Rizwpz6Br1q5zV5Xyr0t6cx6a+awa8c9IUc7gWFG9lK39fpR09oxLv5fIuwJG3Fm
uFqdjdspWy/2UQZ713w1w/aZhtvlR1DmZT280UM11iT6m8g5SECPiqAPMGIn5ca/
HIuvikuMsOsYEClWRW77fbS4tbr8muCNTuP/hWZZYhnVSYmsaj2BiPb40GURFyvz
z9fcGk1fv0LSJXUrHa41pv/EDsxcvAUJkb5IZ1SNAAoXb+jcsY9F84PlrwcAzUWC
WDO2Oijn7in6jorGn1cac5RAGagp7xdrffNcmSZ2/kVWCjmJEpEGamZ+pE9p6+7J
tYoa8V4mLIa4f0CmRKZrtqjjSBlGBF8WjEzEJhOjJDZZRiAnrbvMcfbwmOYTnPMH
N1X9yVr1YUetpHwvPaFylKqxoKGI2p+xCDqPWyE4IQYitoH26rucMlIadonQX0UW
0FPsQ1uaIm7DgXXLAbLbfUQehvnnRwTRsAKoKBlNQtorC5X9bDzum6JfoH4JOwuT
+wt9VWLm/2u9BhHD6wOooutGTGV7M63b3MpVWYaRDuN9zqXH5eW01NaLBMx8Kh5E
vqun3m7PdDcQcGhFiKhz5Ytx6za/YgvC+bqWnA2+3QyJAC28xCcY639zYlSdPeaQ
fzOZBuAKvLImUlXW//hIfe4k2HsJFCN4KWY6n7hbUTp/3JWnatJJFY5UU5vO+wie
JQuSSKpFo8/4npau3VkRj0vQN1195WctOFLeBmAGVEG2BTwXRPxqBxbgn9F8JSCa
z3ocVCEeqnOAmIPPHS3WtfsjDC6yFF9Lmwvo1oDlTed/2q9xL03Y4RAbRfNuvXmo
PQj4hiL0Y9h4PY+SYJ+qDILykjk+1rgv6c2djNZ6JsD5vSWbi/XwNYzY9UdXbi15
3Kb3GlY8slNc1hotuT4JtkOMf71y3MzBKfgWuHN92Dens19jOgzWHt7u4GND4KrH
h2B883SoMZMyZ1VYLcxNMGVfotNJuaOno32FBN2TDjaPA4lEjTCImoJdqWMgmIPm
j3zwhhlgiuOfoSE61El+AFYLx35/cpYu3Ds6QiG3c6jZ5eqAILp6Hbz5adfDCVyQ
5OOyrG6U9y/k9tTRiXtYaWu6HzBrbE4dKKSYzVWZtqD6AsZi8i/vUs6AhPVZuaFD
A5qm7PXFN8TyBKGwx73T9bweclJODlM9ynj/XGVcJHkwRKhEeZwNDS3QoPmONry2
o4qKVJH5a9009RnLK79MjtGgy3gf7YG3mrf9j7HEFZWmUc2EL4pngNvBNWzqwQ0t
/tDOCoW2aR/iygvJ2ElZ1CZnhmkAOCE9MuS2GLNXuaSnKI39T2eQmjCEZ/kkRke/
K7SVFxVUZjnShDgR0ybg4Meo/I1khDCFJNKUvyHDXBikV3W/rQ+MNCs/9Xisba1m
EH+yLgw7vNP3eROrucO1VEjC/+wJVzv0+A8/48zYs261UMXlqWQmZ5+YIi7PHzSF
9IuckD8I0yg+Nw//09wNiYaxSruZ8UPP5f9ygiHFKrAn1U1TdzA7ukeIIObqidFw
Fm/3DJ5pG8xmFE2exJnKsl5EzTMxu7XnBrmreSF4jEIgUnRV9eVt9mecJ5fCQN6U
tycD+o94YWRbfunFDKdqbbLzqJte5bQ/0CpFO9YFjj2MPNXJ1n4PGTV6s0So3efo
CwUjEx+tyYEMIerCsNsPa4IQIRYRP21Tt8l2Ub4lIOHgSXk95zFmrmp6p57gVltj
RTnnbPFpoN1nMLSd2epFZHr/2DSj6J7q7rVGRI39gOJgNSeoVN6whg2eZnfEzO20
Qstc2D8B+Org1BcmpyLg3USDjNWr9LkhPrqixVGzVbCs8ygyGCIk0K2Umh1fnpxp
9EucFsj+0Jprrt+GVC6TXrDXckdbjSD8rBZm1afZcDuaQdEJ1HhLK2NkXm71GibU
kc3a9aa9zfLL5hSLfhgThipX290EmebOw0b06Rj4K6++Upcb8MCR679L9aC1gOC0
QYe2yTIhtu/NX2Ixd/R0CJTg0xO0pVL6malFoegvU+L8beQuOA+1GBaCS4T37wwF
NxDP+yYuruGLHkV9kZgEUvOxf4LQbl6W4BJvijOO8gXGRFbcKmUhmxCtgDesMPoi
du59NK63rCE+zZxpArd1mbdEvYqrnJeDJ7d37awOgPL968t8bNx79IQeS7O3pocp
rDRFdoe8xu4uQSMxdfw/JRnSiRxqbaYczS/Wbuu2wamFKvA/mId6dqgXZsyNxQS0
mGnQk7W1JgjAtrY2SnT1CAN6gMGae718VJQN2I4YhPLXk6rLPyYPb9v9XSBABzNX
gsWhVb88drwTNFZFrrtq9NIJq2JBR3L9hFR7fd6fCbSwaxrWMNTFSQf1PJ/nZXGF
0ffntdtwu+LfDYRayWq9EuZL+42SWBoBYAhor9HX0+tczhMu8V8VIjLkSZk+hoj1
WlffnCjoS+NG5uYbfWYdHxMIxSTdTEb1msxuADEkPLOhpbSylexP0OVzmCHWXsqy
6+++LTMvUpH/GPLxnT6T1nyUzju+OQ6D+0aPilxt+gtIVvkrwnSjCRN/uqCQPJ4y
76RjErmvIGBwcWAO9Yqc3D1BHsBFiACJIfrLGVLAxBY2HmQqb0D+1qDgzGl7Dtqp
m+lfx5MJBgSo2x/s3/my3jj9y74YJLCMmcIkPwclDjfvNdKnNCbcLHdnQixsl9Ck
1Y00kZ2u/iIo0NAhz3d85aly3ffycm/yy2q/EZgY5Cww/H2frRaz8/eS9dvEbemQ
Hji53tvOR4ch6MDVdn7EDI/3gP4JiN8TbplQKAjlbgExdLzjfDr6B9fRSJqg6CMc
hjHr43jUQaNj9b8tdmWvx3itPdwdVtJoiuo1mPZMxYC32NNJloBTrzJ3swGbxs0/
mOMSt6MuRcIJX0yn4H+9gTMQKw95N/Ups4o3DgvAmoSt79ePUneoLU6M7jco6mPh
CI6LWymTSIFeCPo+dyC1odi0eB7F8ep54ronGrYyBATcUgOBUTx2M6i0PqizljxC
o74WeM3ClPbphqavjRSDUCzunzwgS5LGZH7Dar8nDDlPDmxwA/Xcj7KA3ZgVGAXu
NB3wVK2p+PE7CvXqqJqiDG4q67Ilv5ZOa+jmZBwTjFQBR9M/8FAoz2sxguoIyoyb
P0xv68c3L6QfXQlQb1M7qGy1mmbBiDbmNSjq3H0NWjJ3Pmh255bg/9Cn602fRhcY
0BY8M1qWV0Kcs1CgGaVP968EJXyrMfDHWjYaaM1xqoyTnzh++43DwLHRdOr2WhYM
e2/N1jcFoiL68XmrB2VVBxnuWalVPklfuPHvOkBDLpVw0YEz2hW/8A62wotWmcG/
7qAAKZSWknMDiHI0gHT4GCEeiD+FFVpk2rmyiPgyW1OcIYq0DeqrhyHRIS9ZMtiA
DfcSRhcs6i0vqN38rnAGPgtNnFkICPXUPWmEwiM/NAxI0aA09KG6oVN+httQniLh
qklnL7r9LXxLgc46GElCAEUdx8C79/PVdeWERmfys4reftS/2BtxkFhgxD0fILA1
BxbGPdIf7A27b+0Ydz5+4CABZ6jop9cLWOe+C43Rp3YJaxp7qlEoV2PRy5qQBrQB
H+drkSCjAcg7nQkFJ96cBes2VfEBUeAWAQ8GibkcemfWcozP0GURcuwyfGV84yqj
NnNtFOZaCEDZ75jBSloAuRu78QdLZ6Mqu6/UcJ4UNafIqDDda6cET18sctOrXHXR
pqSNWDfdFFF90qfvmBQVpgpT8XNLEg9RoLgXY89ZKqYFZermZaUuLQrndP1PjJtG
/a67PxTjkVEmQyo7GwaAfRynItPHWBMd/MVd/d8IPYwf15qXHckfoJMVT5rAfPJI
t/QWw1WIkzbeRTQ7r5JTgWYrT5T37JgchwkMq3bT1o7yoSZBztcZzYTbm4izAC++
PbN6atZCrNWP0f5fKLlWHvHNNxD7MmiPmd2UPw3KdQ4CE76+KETwvM+Co/tIIlkl
vVrt95YoSElBV54GXXz7KCST65oMoclyBcvSuyrsuWMefL4o2+lbHyLahKZLHd+9
ZSUlHIbEs4PmSPFjdyTBegOk/nq+ABsz6P0/d9YRgnOqSpSgkl5i88gReYxnb6kL
jgiRM7643QamVibGEPIccUaQgTKgSr8NyS9az0TGJ3ueNJuLPECurn6ILzaXH6OA
yVJ4P3bmheGXHSVaxLZQw3uFh7EvcrXqfQPpMndFlnXT6E8telBhlaUc9oqrCULH
Mjhx7zaqnnFOkUOyttdNvDaibGnFMt0FVlbyyi89lfQJQhvy7evImwLZPkgfVkT9
+zxTHnk3gwht3pRm57Zq/7JgsKFIxe4E9K8RtF6IhFsms0NOD27J9dHMitUWLrsV
s+Gx2DYZoW9GWtqLzYV/h3tQ9VX17HxfEcJ6FaENKY13Ky1JnfQIH0GE/0LtLO0M
B5XqMPgbnYOwTHiJlZXF+5P2+3s+exrtpoeTfyze0JQRyo6fbsIiF4mPPCOhylOU
OlLsDLmdD4qllNtDBrNCGwJTPQFqzP5ZkHB0xgKjrO83sSIEGfJtn8VtXFl4zbap
aFFC1yg7O6R5FnqHaO4DVgU3n6xFv97GWwSLAE11//MAC+p18ZPo4fd96VqK/CM3
Lwo2dDVcAJyHoskMnAg3BIjtwkSHQBgucu8JiP9mpW5sZFhfTYmGj/l3zJukTSif
A7GI0w07mGjYPYD2DHJOLkqkrBhA4FeSVTvw3FDIRzxpldl/kjJiQQz47NTZS6cS
Jdq5vOidGMjeb+GoeER+HyS0HCnSDrPQbqbNSriU5Gm8LZNvO76eYbYgC+z8+flO
ekmtNrcDaBUCWBqmQ1qgvHxWD2bY4UK/4qCoxkdFDUKHy+TnVAB9Ap7+jZVYvVNF
A9jlDd2sUlpZlftinZk4ruU0tcng/rTdEEEyKh9gSpDwUwYB9dsCjLWe0p9vGgs2
mpjQq/441mIKsY5gMjPB1scVaCtbkQfYG+JuK5k7gP42tT0414X3SuJdIa0Zv0DT
5DfArb0mu9x6bq9FTTrBCGte1aPo+U7+V+NjF5kpDi6uq3N50yPdbJXrq+7RfrI0
c0mxW/ue3/EAmzYKKFw9Tz4LrtUuq1s6JQnuCey+ruokr+jJNarhy0GS2w9YZLm/
oNQSG400sJDVJDOCrIcIx4vxXNS8/8t3UazlEGoarHPAx2J69zHp/Dwdi+NNKKAN
ihP/+r/+lGsUB7FZAJIwMkCrRQZhftlD3MRcFI5XSFIcB3DZ9S2jtDqTH3K5U0o4
NfU59B2a9ckMz0eB6HMzfr00n9IBPYf34FUm1Lw/88z7ppzwW0+439zraQDpJxvV
wggOtnlJ8MYJm9p26tuYo9BXcwlxIWD9BJAteG/tF7Q2HIyeYGLzdfS1Jh7om3VW
aZGKz1tJgxK9GpVFrIPgshv+Qda/mmgPaTzH0FvgW+2eZQ80pkyywdil83go8cH3
4lrPR3rmh3l2Jz7kAFdQBGcjbLD2whVjY95WEoqpDSFFBDE9AKRNqteALX8sKNPg
M0fIZnKj54UfZw7e7fCXv6Papr8JnlUcRqc09+jaInW9fNcll8K0IYeI+nuMad/T
n6o7xW/zhG/EHafJgvyQhGRBQF9k7ppPXo4rlZAdYj/TbKCwxdubPvLz7olcYjOb
j8y34PSa9EQ/Q7NX5Gvr0pLatxqeZTDvbRgSCHs+u/3yXsCLXFFS/O7QLOOpiwHb
cejBRjCtYTzFDAhkXi9CHvMbC70AOZC97+YKVBJXcZGTaJxb0Nd3uWUGkT1P5KtY
VE87d/luzAagFohmnCuVrLwm1pBDcC685gJn6XDI+FysNwrNNiBKL8dJO01ibWLa
tixE3ozyigObbaQybeQglzyLMwLWuIT8oS1TmppXXrPAGwlU1hRfp6fQRlZdoJAu
7cck6ZuOL8MeQ8M9CpQ+mvu/t3lUFLq++5c55nDVciMfmp2jDEp2LF1BmQITA7Yp
hvg5b7gkXF/MPCoyKfFVyUgDbXK9EQlH7PseY1n6dDQSDSiQ8X6WZpCXjxrsh9mv
P+fxVJ4pmBcvEG3D/VHED1xK3yudQbqgbOgCDMW1PumYwmxJPevozFar8YVAp5YP
6D9qfCq+lJFlRuyqPflCmoL4klS8jDzXbzj6bUgRGuSj7UH8n8XCl+KHSc5Ut3Pk
Zr+SqRC7dJ9MxBG9rK0GEYjhMYOjY0dX/G+CCISuLOlgRK0R6AF/DVI9lUkNBm0T
0SXii1ZC3bjJn+pxwLh9c2jSio2NeDb6M8AZKFr1vJppvGJvht+slbbQXp2+PZzn
XjCdOdRwPeqbJpuKE30sCWQk3X88v/YS3cT4ZDBloo3yEAS8GcatkaFFwBlA7/PY
t5rWGjDH/vS65N5qRZy0jwkYDiM4hI2tbhB4nB7s0HU7BznIDlEpcWSZZ6IK6nqF
2CsE1a4OOHTo1DVopO5neebQd+QunRgUkYMwGz5UpMHrxJ4mNVyA/1bnHVVYvLBe
4rLuTf5PPmTMvY2aaPxQC0DHPrBAmdAMDjQHCmsk1Q2GeQg9qd4qTLzd8pwY7R4l
6NdspsY0VF90k3ZcaE2mV0xz6B/57zpgn7LgQXIyJ0xZv6w94wCxSxwlkcchb2CL
sBpWQXvWyr5sl9XUvbqLO4kYJ5UZMHnLuwW/CbtzYs8DXE65fiGic8IB7Pi7gBBx
0dG221BTIoAUUcJlKHGM/IFDSq30jYOuqQSAk6xJzTXT0grgbpJx4y9TLok//BKG
B5UsEmsWihSfzdIx9933lz9zirjun6b7x3hlFg71JVvlst7thMoKAHjCXqQARCsB
p1pmEz/fYzvh5zrn8WR9F9oSoBciz8iiCorNWUWn+CKULFB6o/M7oUgbhz1VnPg1
hsn7sPw/nkhLCe2a8DXQMci+Ymddb4Al2XQ0sOMQdIcySKrXcKXFPlvIorG9Kfwd
g4vSeb39Wg0XYviRg5YIxp/iaXrnkRZ+fjFIEyUNihYa2QofdLmeWcUcBT/Ks6Lq
nYTvd6Cau8ZEG35ULWtVGNxuocn9T8XtFicQoFB7d0AKWXuZiCeyuGH4xiC310Ho
g57cx48ARlY750IWAKNTAQlrYwtCTGteTIv3XZqrrT77bPIsIhNsBsig8nA4Vk/O
E3Pk1/xKFYzNZHqmDVRoY4ExZyE93e80MYhsJ/5qiPLbZu4STJ9jvylDSJhHMSfw
+yqwrWTi+8s6b3qnjU7FtQTDd6eAueXwtDUa1kOZwVUD+Lr9WYvwWeqe3u5vBed6
FjLGxrTgTlPdqOWMLFS1WEhwp8HZEI5b+hgNli5sCYOA8VO/It10/tB5TufcRdUc
eOjCBmPp9LNuj51s1Dg6BA5r45hFZa9tUlls1FkQpSOjeqOWxnjaMnnjmPilQzfK
M1G6Vs3TJMhL+oNLwMrCa8btvIVeSwr2LZV1NzIAJOyzF5+sI/bYcPTs4ukb5zc+
5crYe+0JANQy2nxzrVNPTWbGJiYQBudhCM32rvjPLCZfHgjzcHbTzYATO4sw8J/Q
U/Um77gZORo1F4qvFHis6mxa0GWmn/2e6I8WOP8G/lxdhJ+bSlfmU+hIa7nI7aXS
BC2ujsD26hiZO0YPSfEdpj+E/l2QgxiEri6bkU9Is5B8GrZxHUKQoN7EMX8X9683
/Kdp/v86B2cK0x5IadOJiiJ9Otqq+tJUiGk6hMI4hNaKR98CUGVlIriI1KrGrOKg
BWGgWM5gaNIE6pdAnrtmVBlKoS0eaGmTEfl8uKmkgcyg9OWIL5kMpHlKW/Yht4z6
XO9Rh9saxVUtni6jxxaInUMf/C1ZOHl2rb7uPId7o3eZtLHoU4g6vDopqQbu0vqb
I8zWnHCO1P1E7bAbQmeBSmzprDit/ktm07fbld8tMVNPqbmBemeR9lNFc+UvJ4PT
66Ca+O64tjzcCjvC0I+WMS4McPe6DvIJYT8tgyuG4QwNcRtFnRphJwZc7Skp72am
jgKsLtGOfnzkC+JMlrcW55A34kYUMQoHgmt7BRgA3MNXLwS4EHZ9AfjEsOMSGuzj
HnbNOchMVhfqMbCBNjuVBnEdXkYzOdTEWww+Ok6QSie1zdTdO0xVyL14LOdZH9fH
TFKxGfaNYliuWMKSq52RYuyTR7i8whI8PQd3e6NIvcYyRDT9DBaIu/T8Xw+S2I78
q+CgJGlSPg5NFPK0jWCFj+CwVBF1czXKDy/wEJmefgefSr7rmqBPa+8FNWl8Btex
B1l6UxY455PRqawuQ3EMoZ/htepaNPLXCGQIXddTqeWQ0Ew9PLVwdsIDTgdRxH2W
eaq9ME82YjPEP15uCgUBmsh2tdsOkZdlh8wf6Ruqgi7Rn5aXH5EwKfm4fmp/NU08
zRzV4lniAVil9EzC/59SxtMcsPGGRIj4rNyhYRzFPzA/GKtwsjirPpXTZDrQl5ip
cl8B6Ywq3Uwpi1CnnaQqeq1ggDs8PpZS+bq7qqwscoeYIsVdRmvNFvmVxpOaykaB
qpf0gj014/tvv1K4PItpx44/9CpfGhUCFEfJQkoewB5AW3R80duV74cGdfNR4Lq+
E5qensRB3STJNpjamT9KROMJuMerTnakbdxefFIWfdRMEDF/LYZXN+cxoYBOqNcw
DFlfaZbrk/htwadaTwC6r+zf+BLVAjGj65uxium+HnICouzy4iUQu/WP8O2Dgpv3
pD71vrzVoYk9LAPdqomXA2EL+2wlTI6i2C+RNiRwabC6KhYshwKPLQXznzhK4dBB
igGZ7rlseblll/lZcyvv6NlhKshW1cFhjoz/670pLD5myf0ohoCeQi5jay/OodGv
yylLnR9AyyUFT1lzDHoVLdV9bxhMLa6178lEbOyM/9I8QbXurkFdsfaazbv49DIh
XSDzCZVA6A/YUebo93bwb4NKuaWEcC3zasjiov8XVrsG3cJFezqCPnzCkN4J4geQ
/5NdC+ckMXr4KfDqdCHXr4wrjh7+GH9xszts6RUK8V2fk6H/6AJceDeIlGsLaL4w
W5OpfnEC+pU+LPM6O9zQ6QvzRKUsPcs5n2cdXiITdrsf/MFlrz7OrHQfHM9HDASD
f29W3R8/6N17TNgtw8QOUthegMZXKP3n5phDL2NPUlBVjhlxHQdJqOrKE3vKM2i2
eXUroSd6JWb+Wg6qDlqDlEj/fyVM8xlX1eqbNwcxq+SwcsN3iMui+tKyKt/CsPx2
2rQd6AJcjdTVftdc+fF1glAcIYo9InLRHe5IszjPYOpY7nfhAtTBqcma4eWyXb5O
FueZ1Ck57Bgy1hWE5uQBeJaHrscGaEmSOSWo+k5BUrWPZY5+ztkPpE0nC3MlrP8v
WN5rLhmiXPd1OvBXT7xc75MYwIf1sJBYWJZ0BB6WGhsv+WzklPEVMhFS82l6toZr
uI7ORqzmGaXfgXgQ7MVs7JJORkYItOa7OT/pg5bBPgPe4TWpZ8UmtVg0ptck8Kvw
6znLFeFYP+Qu1LhRgV7ihuQgf7gkNFz+S4Ibh7wPVTq8HbOPoNvytGeoKXMSvBqH
WyeyKrtMlZzo1C2LQRVd5bo7a15rd8dy76fOUs+UiKuwMLLRbyr5/H0eHuT4B+Io
ou3k/szGvkeF6tj9/9Jl2vdz6/9sz44JD82skYF8YN/Xru1sbpl0BPSqeoMVP4zF
dBD/xdQp/ZhPU9dFIN3So16nTdzUHnKRP7OduWTJgjUYRBqyyYBPZEHFuGkAjmzc
TdLufBAfE7S1mnMWVuWaoEnX59MTy72ZP+dlg58z/JvlmTV3G9/+kPftzK3UgSE4
rmK1SMe/d4Sfe4TWWYna2FueC1OL5IUVRSzsR9QJ1jeYyXUPRLIuW5WCSzz4mR7l
KEwzHV3S5ni3yJpArBW5/edkHX6T1LqbzutWCGPSQtc/YXBO32Pxd1iYv+7s2TzU
WJofq2jsxC1vuvKruFIu1imQzkjKZUWsHT8oIg3TAS9YeS+iZ8j0TkxvIFGl9wJ3
8LN2yz2RHk7nf0WI8onKnHC5SU4p8lskd+lUd9VwjakTrzeIxdztxjLG63xSgDA8
t08sl0m65HG2sy5eYqVyRt5Q1MF5IbJF/OSJXpwkTQ3M3fiJj+MYkqX3QAk+eZfF
qGyzuLSgfGWMqt8Zb2QtQYSQ7WBiqzAA/geih5hDNi9Nu70swjJ/svct8k2+WcfF
k0OU/HuwK1aHF7lldRRKMyV4YsE/0lq62NThUNIS3ksfmKWPxI7P5Dw6qBkO/KBi
fdVkWxvHGGO0h9VGJ+HNg2psWse2mp6bikDpYzmeJpdJdxtzQBHwHxfoN0/uMf4K
pZjy+p6D4ZuFIUb+XeiVsMN0/+ZxjazV2jdaNUSC4EpKDiXsaJ6yJilcsr+AIEP+
mc6qRfMlIFvDN04ThcMWh49uHrRFImuMi4N4BbILt0zd+lpSRnsyQzu+GnZbvTEt
jwVrEpjJx+qs790Ik7TiUMqJ2IlFeAyBBaS+mvJWV4k10xTQXFfi7D2tvqXlsBFS
TTlb5gnGJJpC23AD3wQLiwu6KLY4Kq7SRysvqzpv1RHyo0dTG/hsyCOEc/2bffcM
CqvZhB8IDLUyHqRlU3s0LNLRezup3lJp2hQoZZMAcI+Utz2I0b07vlUbkfONazLq
LG++0b7JnIWC8XivD5MA9tnh5Mc2ed9ZpRfobVRB+bAyln4CUspxet02jChVZDx5
uU3a86s9dk0kppUWymBo074hybKSHuV79aGqNG/0PK6u+MBE9qmaWPYda7vZgrFK
jc2TS1mxakF+D7F6nHTJj3Zvp2uykeIGNexA8y1xYcN3RNXTjQ9yh6qPPuNT78xf
YPksqwRvUZMty1kucnodDERy94eGKkqNwZYvVEB2NXU/izdF7+tqRjHPJ5vXwjdz
+V+01eVLb9nFxwPBaUF12vBQFrGkaV33IuEnLptCCdSIS3vX97Nn+xDWRRHIwqKM
P/hOXoXa7tn4JVjHByOW87wRAkcak79Bc1sq3PHms8j2CKRR3ryLJxEVZHuB+z+v
pFYWYDBAlXfK5Tm+xrIaWrV7IZ1m5ggBhrcSVPvOGzwNtLfPfct6QgUki4f64TBg
slcIAmji3pYpFM4dnXpgWvM88B3RkHEZJfV4v0EZsIZFXIKAJkdGbtuRsOca5bcr
s0ZD13lBd8xgW+uDHSV5RwgAch9F76q0sDurCtLLMK2nsw4T9In4B+GOUJrVobeF
1koa758XrDlKZllDDGFWM0Vt5QN/nxOM5GEOou/nLba0I2c9G/N6C2SgK0Z4Dd4c
uIzlffpwM6OwG6qzQi7aq01cbxsgOWUD9xCXpwMVIqbADKi+mjo9KIOop6DwU2U1
nKeIgEh1o3X9DwL95RUmjaAaw6pY9+VCc6/zRRU1zQzHI5Lhlxx5JcyEgpWvN3/2
r+rXxZSNipD2T9S/yNPgWT8nZlZ7bmw+v0dCHufRLmn23hTckhN7D9ROmmi2CCmx
Q1Wok7o0QTsgl8EWkpkaSE/rU1hyG5DndMkboL1nECQAYyE8zeKQM2DfPGQ2moA4
wZWmR14OlZCkTARTLUUud/tsY6Zs3xvn6EcYbXHKpkb/vXPwpHIlnXFQLQPFJXf1
l8aYaZdKgiWg51Bfs3rRzIcYmvgb26/nZ3FdRif8lMNZESQFpmvMjsOUEHWEGp6y
GMQQZxc+4IUBOJQAqt+RXh2exjmBZRqFpv2u8oQ+ZoYQzGyRKmsRoX+RKWb8z/ge
JIqNYrHBn72FD6bS79+jXWZF8PEAyE9bi17L84LEBvpJ5cdiJhkygYQW7PkZSHVJ
z6PQ/p/f0ulpW4nQ5E8oqJZEpODkk8eDlYV4Awy1i4Q90myv5PZxJnrrbcSa+tLW
ro5+coH1H1yGrPc+QtEqsZ0ZF+3EI2TxZKHJjJlBusT/56lgb6Ea3Wsk+8SKsPnb
ljHEMGFMpOs9VGUXyR1wzsKFWq4Cl60NBkS6AaxAxVg1ZvnM99RpWzV/7Oecs/Eo
gyU1Kj7bRr+MmmJqQX+qPkJwuXTA5bzyl7SbfcneKEhP24+Gs7TH6At4Y/OmcB+k
LdSdSnzjGOsWJJFP7LgwlhxeeQNSMknoDK1jabz2PcM2wGSpy9EzuSeUBCNoW7Fp
eiK2+gx3VMk7wkxP4y2J37SaqROeTVqwIQS3HM1uRmJnjB7eXdkuzX4GUgAqVXxn
d3AtfCjjtZBfVx1RcDwfTXbmTuFgUXByQUvf/tyZ7aS2b78ssVnHQ7L5KL6vy9De
uojqvS9gc5hskn8rcRxjhzhTZ3X1s/vyIgMR86uFZnD9Xv9fVmB6Bn2nxFF8S5Tl
tKz9BvOeYckUGR4+4kqYfaNNVIpGaZTLAZQd1tnBbPgiPnOZHPGbBHUm+j9IBVvW
wfk97u6X0wrcnvJihSgezqOo0GRbrl+hdqvRu5t6nZAjcZ1X0vvMHyg3UC6UaozP
p4iepgT9ynpn+eP37kBM3nFMRyrM8d6y0DaetTufHrInQKcrKqrFwrW178OXaz7g
jIbLSfycBlfIna7Gk2Lw76waoDBLJuNTPRheB0zLRUGLId04Bzce2HG+mf8I4HB5
xWeoifo/T1EsSYPVZKWu3NcAXueqg7sZmh02xiwkV2DBCZjzzLwH1VqAwOAPdVie
hAGxM723Vz1d77j8mnICIe9mjxKox0L8xVTZBriTIsFrvXJIMUdejzVzx8R5Qfvp
CEgXOjXR3OX8exkbu2rIkkwzwu9kkqznkzSBXiSU5OqG7ITUXCd1ol4QYzXaNeZQ
652kmLs842EZPkCMu8ZA9+3vjR5iEVZxqhFJsEfEsKi0MKjvdPfnsL/D2ECN0GJM
3wxrw4imXHqcPmgQ6Ui8c7V98pk4ztT8XNvjnDWlq1UsBCbKMm1D+o3xdia8LCtZ
rcGZopUyzD9cywQdWdtw07Y7L5BctBAz019b0VOr2AYYbXJ0diWrp0TpE+1xGOle
2dzx3VLbkfsTxiXeeOLmeELJJx/R8R2pKsVTeGwIMWPm5m2Sm9YOcJ5ChvXd+RX5
aXytTdkKXqN5ZgJcP2eSNyJ7LSRzd3dMvm3dJeAYcBDle5ivncgKDKQTTKOK1u7W
OnvnzloAAyt1P2fXrYG4GcW8vFtmt2/pzxtN5J3gVDXO2xbx08eRLO7JGt4DmBJ5
yq1x3hBWjprQ70nqhzwMgwKu/GAklwQ3CmeldNLB33rADjgX4CZmsr1a+bulMBRq
eKKGEYNqNuiOwrD9NyusOx74A6GKyD+LlzpYf9inNzc4vkXPW/JIDYscmjdV5srb
9q5Ev4HNxplNtd63hzKpFcnGv5tuUO58Qq6D/VCtUCsQN6OClgY5Qv9eHKX4V98b
sp2Jk4dU1CPqSQp0LqIk2lCrfj2Qbo40uixWtLZkofLDp4d6d5QF7G45iALkcvdm
wedJDt8m5HQ5epll+gLlQxd+IxoPagbAKQLRn7j8X7AqubU4ln/EDosyjLrfWmZG
2QG2PYCZuzms7vQwqYgsBLDAbOvh6roWDq2ju1HP0XJ+GBiATYRVQhB2TF68d5Fb
e9a01kDz3T0I2fe+6iBngbblpjWPrVv6cobPOeQQMdkBWHKIFsUK+FdCl8yJrdPD
z/LdjZpiBNXyNRJvX+fU8/BO20Ipqqm7ccAZZDgt0nzScZQLLDtweOYsXdsqywQ6
T2Jkbq9t4R8UzOJeg9EqESKOyUjguBP1I/7yNAltJ5Jb5ehiNdi0h2U4iCcMA8qh
l4DV0byoU1LX4V8AnZ1D1JFKYfJwVRlg7CHLn9pU8QXhcmHFUjrwRSPOnPFPBvP9
daTtGwYFZ3yJQClpfvrczQq1OABuuQsUuZNHCvW+M517ymiClTr0IOElKrx2RTb5
aejuC2NhVt6i0Fdf2XTP+xWzIgTFD+kiah4tjgcVqkVtkJPuQXRRmSpa8F6hP6FW
C9KwuilSHFmqJD5KFR6Wfy0BLGV3AjgxP/QR7i5F5zzVBorvMsVIKoKDMe5F0zd3
4yzwXfB2RECk8Fki64Fg5R8dCod9MqUYzGs7BK4gz5j22KL+DX7eFyuz49PXCGaf
+HmA2WmocJMineM2Bly1da5WT/DILjRsBqYiesmrwGLbocPhlXBHWfb/x1g1x3wD
Im6OATmGuUsk0Z6hwwwh2yG9z8PIqeZrRqagiQnIj6AJZhrnC5zjzORCLWjCyaXp
IPfltF52WXCvRbwNb6ohgFCl9/wKTyd+uk24vHf2ZKMjGJEq03ibk7LfDHJJKk//
b9y2vKk3AKebu22BEY1V3JVaNnlV3iW/u0aoj+vIPswZ9U0FpuFz0FsmgnDDUpul
yZSzXWXabKrJdJbm9hFo/Vxm9Vvd8MB8+qLd3HzWiOlgY9/lxypxSUpg5W3O3GS4
q4nnpwLiqsPpqbc5sgWZSPGrLpKvpj5sy3hL3FJpXn1BsF+FsP5N9q26+qVsDncS
qDw2tQjhaTUCb0OLLEDg+WE0bi8IXmckvxlLytzMrWIQGvf2CWwIcYo/EsS03IJQ
/peNe1FEOnl/kyyzk3iuChZaYZRfhEM4uZm0a9K/wJoNizOq3aJ/guECCYVQZPqH
KzboUGyUx+uphaaILkqAgmmkXGLDhiT8Ptgb/1iWpu1gtQJi1zZzffU+OxyZ79TU
8nrlEc1AmRnVXP9jm59g0pQ4nCod1yBvQhj4v41Lm+yMIeQolRg2mpun3KdNm9T9
gm1UDsl9hanX8IBQh/N/i9+pQCDX7QlqfxZqOW2xD6zTW6EP9WpZPayOlD83zHuj
4r1tbAqIiRKa5J0aIi6DiLbhwrmc0oOypwoOVs8sqqjYfM8L/hbDyNF+YvIjarm5
fzyjZ0nX5IPFVA1K2EQBX3s6Bp992W+hA/Qk3yXDtqvdNnikGXDg7Sg0SitWcwyQ
G2heZmtrAEnOLvNJ/XuB6utCuGQf2KoXOeOrdffh4g2FWHd5l6c+3mbfAA6QCoIb
WSKFRuylY+JWG3t6zLg0NV8AHit50gFVGeN11FHXOBUCuPsQDjl0MCSBwWuHzcUw
PmGJvQFgfN2gWDI3/m4bDtoMQvIJ0Lf/4+Hl+h5Z1AYhucywaZofUeIDWUvkKKWN
Z0f+2vx932fkO8qndceNwzXzdmHLObcJJp8sL2ROaBrX3v2XkcHVXqVk17jDh7+3
aEONKFnuonGq8ESDAwVWZ3+bfF9Ancpc2uAA66xKQkEUWfOqAi7foTZzavShMYU2
8EOrHTNN3MnIabr//O3XY+vXVCUXReDYM1S1LXqjUM+i5unn+Tg9PdGz/Eqkp2/+
967q4vfjFr7iZrjzU0umLM+ZBYQ9TdBmeMTQpVn0l9mojdX/7C/eylSSkZWEdWzj
aNEYJo15hBLezzkp015ROTBVCYtc84FFds7QZr1vKhM2WaUZq44lcmUTAm3bb+Rf
U9XZLQVopMlGbs9LI1IvrlM07OKZWSvOuNsh8DXnCEt6zUlPG8VCmyQtZxMXjKic
LXa0N+ELUjjiJqaeM6xxdoPLAosNtD0N7vvdG+T0OxRrdM94/QEWXUUUc91s/VK5
hejYjv8pEqKDu1OnD9qsaLDfX4o5iGnH4X2k6GZ0IsGxVMFd0dBU1g8PA1i9OVSs
A2duy/ojEC+WZa6wUR+OOD3KftZupx6h++G0FAWtKLnaVG4JIYupNdPRTlJqqRPU
F20O+aj6daoiib1I3KcHD4w/VZLPfjU2RaAc3nf66L7qYd91rtiYdpkce0oTnIyf
pIUqTu6XhJN+2dNW79PYzA3M6rQMgBRDVcm/8VTExFqoK0oTQX+ItAn+wkTQ6N1R
ZH1f3W335uaejxPe2MdlFSzcN/t9abA9GB4gdC1vhLzH7IAafAlUKAOjtjnbIUba
N3Eg2VF8tN2YZBMUtWnF5Ucw3IgfCmlflfqwBpWuPRKpM3jdc83QkifKWhDIbab2
4xB6lp4lDj6flwPCXjLpSwUh6ptim8xBDCln1utALOXqycomXWYmoYdy9VBqKVaM
g/zY4VLOma0nb01Im3iOLtxvJ2v3rsmeOAEYaTQyJIjWP29J1ylMHxQPgalEOSpC
LXE4zB/njGTCLzr8pkYmFB+llx0712Qu8hiadXCf5FqRlsg0eeTZoKgjSmG3egO2
4Hvp1ASN2xZMwiKSyX+w2ApFSuAcBzGnPJABwt4XCZreoprUePA1cm9baOkwKw43
ryeBzMUthpW1OG+PCkQZpmNga+2nCltcwY5iHaNLKM7LYlBPk7VhnQR09/P9Z8KU
iT2UcIUzcPWPqRWC3T92doWCZ6W7azkxZxtLzmWMEMkrICtpFtg/CEkvi3Xh45wJ
bCf68zWYrKKgLRmqROl7PODNo4krAtucuxFYJ2+itnSS4eeEV4bP3CnGtfWf/ZpA
yakr1AcB2Lsc4LO30pE5NLIqrnjBnhNaFrpPk3ILGlkYfatdxs6y+Vz+zyVZqy/C
iJz1790xLmepgVaZzlF3lYwvrO9vqm/RNC5koPBUxhP6zuR3EdvgiCh9gIMcf+sm
Q8a6VmcToAoAVEJClYpSz36OI7yuD1bqpQW8qSanQJFmhGIsmPt7RJIcz09SjpFe
Ga8/NJxQa7K2hheazvRnL+Fi7yB2dgdke6SO+ilK8Ex9USaX6jIdEfbiSEl5wgMT
CVBETXfqkYgcJMFKYguWxdV7WgNqXGdIWcam7nMQWSMFdIJvJ0Fk2gHxbcZpprYd
D1638JLofGkWMJk3cO+l/ML7FglKA0+CcXt0T90tgienXhSGeEW2F/JHE8eqfOzJ
WDXkSJKm+MO0EHgnuCQyZtc6BHxgYLu9CQ1WkvF3dACLNKnv/yIds74g0xw6v63c
dKtdOERNIMn0Tsf5hIzcEXKEe5/CaDZUEeF+TJA+UWsilSTQSlSbcDe5TlH1Vvx9
YbV8PkkhAoEdrF2TCZVP2i/g/iT7nttv30P/qtGR3e7WJZUkDdkrtTVpQ8FqDFnP
cHAto8bZx4G/pVmoesoC+GPEd72O2nXOXjc6bUTNeqmJncoFtl/ng1xJCqxQdGEW
FMCFlgGbc/kiDWHLv1dkgy7hTJ9AjUrRu4GXyLyJ1vZbybu5lG2kqOCsi9eI6ssm
gCaYZOV4T3ia8dQz/JlA3cs3kwuRyidDOoR5pCYLLSOEAIY3p5gr5VwfZZAG+MT9
Hze1+iunsuDLzlexoMrNw201/ECVCAxrZHSckf8w/687Ev1Z7o855Q5YEXeegp8O
IDV5kXo6hm37VkYCaR07vYbd4KiMBFxkali1sMEPBjpsEmZ13sMRL6wW5VvQHvS7
8pI06Al6hQA+QiOXrYs7oGeyfnQ0P3Wv4CisinXnrB7SC0vPXCqikLCWCVPFhsoe
RlrBmMW3CFyOYTChVxEk9aDMbiCLyU2FHFx0uI8iXIaBKfm1rPDb2hIL/hXaEZlE
avP+8whYT4T6xuPTWr4XIFAHXwLpSjh7qtX+TRbBhVea1nng8IP/8jFZSj+AFlFI
xEZgl404kFdWl6+a0vCYqDUIJ6gjKr5LkgoedhNBuHS9ysUxcFD6lSb3yqG7jEJy
FKfaamOJQ0/RspOEwX1RbWBkPIlb7yPdHH68oDS2k6hGz+luHPkvlAipFwpi6BgY
vao/5l0C1PfigKq6KHFeOPEf79U8yOmpVItF4iZZwWZWw93DqTVNyQ5BcpuGTAbI
dYu8oPGsU639ytFVsgN2aniz3SudiBGTfx9v7HzPMl7m9LeXO3j5gvjLjnc/hMlF
ftoIcIMj13aeeJuQTWhX/dbE+z4fD2xQ5iJmgJ88s+Od5IM2Ka58yWXv6T1xlj3y
KOOcnkAfNbfge+JQQadPWVJhUuDLciqsrfa12+YE04BKQu0C+hqUpV0J898G9JiE
xK0DH4tGOiDSbiIbtsNe2ZjToPhvquPBh4UXp0lk9McT7hUjkpVcD7Dn42TODRIi
jfTBB9HDZISg+bbVYQN97gbCHjMpr1I77QhQWr/k3SAoTEl735wb/YYXr4tVd77K
Mc+UMuqeQ3CTqhSoxPiwtJ8yIgI321zTnLgGh6mtiPZOCOkpT1SeU9IRbCQt1yPl
8hn7P/y3mJL4FJxg4QFxKn8BHl6HHfuvIvtnYqtH1V0C62BV37dIj2jHPcr2k7eF
AHYOCPdg70kiM0liiF4FeUCYEvdS/rc8hDCI7dp1d440BsiEQHOrw5R4SwYWstdv
Re2Sg0oZoq9K9g73GrjhA2DPW6twpXkmBIpuRweN5fehvLn8QxUybX7YEACIYYrN
JSB94oEIlwnbBe5gG5ZZZ/otR1N+6D8cxd8olreeizP0Y4QWVylHDBOjmjgevBxh
C+dkAlNIBK8WzdSYmE2XTWxfwMeSSJ+42+QRCaGCksGVQ2Zoiw35wfhsZfby5zJU
mgCP85ogSrRJ+kmjb8HI5NfvrosD+UoySvsiFFW4DNu5i4Tf6HlkvaYsl/K/Xt+1
IYPaYwFSMqKmbWz29+ie0CpIZV3ERwDUg4/8Ip+HDUwoUzdrhCgWtQNu/iEemTZw
+eZ0vCaawljaL9pTioSSzkl09yoKgXl7wiJwH2YodSFLWm3PGv+xDNn7j3f8FEWF
Tyza88AR6pF2ZVRHQkJJLOzpQS8KphIySDhtO+4oqbsHAqhPdWBKZ8Kpk9e/WiGS
wpKluBRIjeU2kRQKQtn0qRMKnTFpFMeHnmQ8StlOpqGdCsW916jYouzE+3wrX8WO
kBXzOHH2PYZmBbczP5NF1obe435O9rj8iizPPyHEVmPj8dbFOICyEJiJcOdGgcOp
Br8i840VcfB1ERZtzwiVnifBbPRhnDRysk9Jf6H9Q1zB59bLP+0p8LsRBgH8C5v8
WFAdm3Uwc3KefW3xX9/q9U+LhzqZbrqrF8fGaM3+xWaMtMsWQD809XdJCvmDZt2x
IaBluX4CuNQwXDXus4PPt+Z7kd6rv0v3ra4CJK/MR4rp2EiEtdsGiFI8Rd26Gtz0
4B4DpMQao+WEBJAL1+ky7beAeaCc27Dn17jmNLGhI6L1BOc4AKxpa+X4XHEOrJMS
k1jad8UjIpb+vV6VA/I2E6HaZwU9cAtA1UBihcKocqAlMdGCPiHmdF9CbeYOyMy/
IFuwy5o6LD8J7/d3PnXYJW8/VJwyKwctMZJfG/foaWO7gQWlYJdklIBEWuwBC5Sl
Ed5TVwscM8yPQnZRLffg2E4gRV4y033Tpy2kG8Wmu9wYwWIAXawIxU6R4iVVjXEh
gzpMLU1YzgGouaI8OMlsHKF1CE+nQneJyTu5FRswXUBkYWZjD9lAQBVWYg0qq+wW
8QSST+ultUuHKZx1cGPgVMctBJe8VAuiNRJ/lqK8A7MQ/UJncmhmTD5lRYSdVB6D
FVcdc0DnDFM3TCj9I3d3MuU5CMemIcpqz8wdwRrCaPv1LbhorbbqibMZ1gEdl+31
+NZpc3EGTG/hP5xW5Uj/dXbyH4Mb+7QsMiRt2lRpmYqNJWE+ecSSUGm9slliW1vM
DsojLCresGMSmeuylnhpnQB0rMipghXIz5u62rQuFKOqIT/loJhhnmpEzOf3dMVL
RqzMvO/BrrqaimNF2XWCDsV8SVZNJhFNUTwwnhTKEPPvpVk6w7mR0eKfh7rRWUal
MyUQfVUb9IAKJfncXj2at6sCg4+EzZbgdt+4C55A0WUkhEV0nz3vSd+caxc9qPw7
i7js3EvKHh9XT/0S96CY23I4CG3AjDv9X9XMJFkRHdEjULdLlrzJSAz9DD6cyE9t
y6k706m6QDJO800ajg3LTZ+OITxN6yMJiRVmihFwQKNLXKKyIrxi5X8f1RYS0SKR
vkQDZryeJpJxYkjOIdZBV6U0WwSJIwF1W0KcRGsEjAmxNnF7fqeCet0NsK8VUiEE
viopuKXv3FY2THipVLPtd5TANX8gy4do4TamYnJc8siIQaBAVSUWaN3A1odeFtWH
O2BnoJTsFPD9taexnO9TBJnICH6Dp4lb+Vn0Sr6notytVDhC/7qJ/L5DdmXm4xX2
YG0iQKrJVxoSAOmWF7wEY0knXJH0AzDTM1eCmEbnQhDj6mTRPymq4K0XliGPvxJO
OLtqcOBT4VBqBmKoyGjRCgoCJg8HhqeJ+l3rEX+USPTYm1MtM943U3l/m4DgXWlX
i1yhRw+I5Xcw70SjPyloMNMByfrRcufFwpBwMfR4iLAE/ng3HTIAQj3i5DcmP8Zc
+yWFqktgo3+FvsaxIQ4W3+xPpQH0aZK/o/7rxxD2BlHFKfBWHW8k4orotWGB41sh
4dF9kBQNFP01KerL389MfkzYGoAfPZ7qk7N7znj0EViWQO88HA8J+4Smm4yAQBST
4HJMal9mdK/7PaRFbhBGHLItvC15ZSbY+T3WLoj1DBAByqyHxN6F+afQCF59qepN
ZzuaPxIqWdiTIF1Qu+W+vNrO+MprFyFoqkwgeLypWTGG+6xw0xq4B73Tgb/LLGH2
sSQggVd0smOEMNZ9mmYQgdwMU6JXColVx2DoVSGqRh5rbmLkP9VjPfQ1saLn3s33
dr4Zfb2ioMHiFYS7rLhwKZ6+9zxBt2GWHB15Ox+ZPAMvwCOH8HKJAdqnXjmdCCJ5
IRMn7kTc1x0gI4K23bSRYzUloZ91EhjQEOZePasQRZrazRZXC8VE/0BVjCPD9LFe
clDTCoGx7cnXKngdFvL2Ja9pKX8QOl1EVeQmhJj4EXeDkaVoURsLKPuQki6c41rx
GlamzzfwwHtHcs5D2klm9cSsRXx+SPs7aKvoaJUh6HKghPmpTX1hvRQLYJywFSLF
OER9SScIdrbQjxSvhnJQG+CNG5FLZgAv0MbLsTdxWXroEOgr3HqMxOVQopPNxjt4
dWUqFim6C12Xf4J/JWSVCGsdzZcMIrX0UbWuggPCNvuaiBjCOrGLWTyClBjmC7BM
iIdQdtYsVvoL8WshFhfHBUn3KANSwgoJi0PUrwz7FN3YTIUumsrdRSgbkOASnXw0
3yAAX2s8Gdq8ONIHBCt1NRm654wM5dygs1WGhhKe8bRhlgOlpluez4DvWcfWKz+S
12Rc1bJxpDnNEBY/Nud2xaFJc/GbRCyYZpam2pxVP0AWIX+Jtc85fXRTKIs2DOMy
r3uvQchCnmaK3UvbMVsKHpJDDYJr1dg3XNwXqxXjnNdf9pFllANf/ItphXnOe8lm
wOluVvOdVP4kGmI6fpIQJTiKwia8QPhaoAtrX/rcZU917HqF50lJXaMXLCDOjoRm
0SYAoQ6lWViA0KjpzaF8lWmCtiSXQk+AwNUIZPFv55wtA5OqMmUAG2+qSpZgdrkw
KCYkhTzGzkOkC+ryTXtZh0Vvn52+GPPN0JRF4HYL2eTf2S6g36T6D3+RVjMqhies
5bvJX71ACrd/g5Ps+N0zITmgcNndBViI7uOIdfUxh9ZUbt36XPKez7Dxa0seAxbz
zzGvx1QXR4/q88YvQ55Wr5RvetQMLikYKP0ESn/gPzUaVsTxzGq0NobbnrA6spSh
JCMqzeCWRaaXjesTimMZpxpzF/OW+48MTAhLlQykfawOvExirz3C1mBRao1GhBjF
vZVA05UorLti/lv25CxlEBejkvUPhxbh9RtDUAjHUy5VjZ3PIpAXZJ5uZVx9KQXZ
ZvLwdZ4lxa1ibd2fc74phP4W+YhlhFjhDNULuBDaruLEtApcI5cKlyiShtsVfCsR
47x3/Qev87FPiWuFT+mVrGq9b/m8OXJtWwMuchLfr3k0Dey+ShN07C4Oz1NYvLUh
fZbZ3hg5ToSsW2fgSe4AM7tddk6IAh9+HkXsfpq8WlbiX8YYaNWVxD9+0lkHh7zQ
NNauwCC0hbOCgg/1UaSmdK17Ep7sUTjPAXx5DW8jwMNRRNGPZjXOPPCMiw1fuobu
E1K/5O70HtmqMleWtiRj3b+I1db55ZVRlg4QuV4eD+KItvl9bdR9MYSviY/88KJs
mdkRBhC5j9B+gBLHrESTmk6oYOIiURC+Jd5w+9idv4cdKjYqX98K2I3Lp2bZevor
iK8YeS4slV8G+2NWzdA22JLwMd8V/8Ey/4WBUBx8M4PL8aV9/PrYrzMO8zIb9aEG
XeQmTVOmC3kj/PkzYwPlx9Xmwc47MSXtWxGU30yl6IPmCS9Qk8UCjtyF6QfxbPrs
KtRitSs3vN2IH0f0FuNegaLu9jmeJFj60hr+G87K7R6t3ORjqoopG3iDk5V4/9JJ
UUNS4jovmw1BOi5k6ktOQDNbQ46a/eq2dd509O0Y4iGtd7B3k6yewYFTOtHQZ6U/
oqydUZpIBJ6IXfhp7JNZkUHoRX2piV0PtLgU/05uEHVOXdtoSsAJGiN3EZ/M/Rb5
DZua1eoN2kcN81X5UrEL126BKqqCVD4WENfAg3JTOMGVSxAsVhdLrYffGURhHTye
vaXnLywPGTBI9Uj51CgCEh05Pm7vlrIelUzv3qpnaz70EfelNpl9aUhurgbNH95Y
Vw3x+xuiisHZmB2xkNT9kBfAInOBW9c1Lp044Um8CXY7vXFFrW2oaP+/6v7Dsg9o
+d4wj16pLI/Gjev9+25hB/2FYju61saeABvrYIclsLGiz/YgB2QdN/W4AFl+xlmv
LGqOuGYWsWFpVVeM7n/F4TdF64OcgqMIMBMdFxlJ3DxmzhfDnX62RSsKd7otBeST
qzKdK/I49Q6eFSbjxBPGXpHlQLT/W6w26v+FuSeSnAI5ncgjrfaujb7o2bhVg8qw
D5Wv7mnMmEFxCdDkKFogl8Z9SM0sngr1Pmyms4OTxyfLjgXIoCafNfcXGXl7WAWk
CZgQs3wdxIDaTdD7lwDfzOP6Qs9qdN0uqSJmoImfXmS2Fh7drF+GU+wwjJDb5mA4
49/QH/bxawiHrIy3iNa/xGj7Zf0vkd+wTghYrU7aRMtLa8GXu4ipD5UiLglTDnv8
kYcNiJlKGiAntOQDiL+lS3WDk7MSpq/4TI6XMCzIjA14FHWaHJABLfbnTXaqYxWh
uRUCpyIVFb8oeZ7TmzaB7W+QRaxZG1/KwFkSlHPeeoyfgJFfBCrBOnvJFTkWcQs8
OSj9pKRUXx9K4g7TCbmaSgy+C2Krap9JuX3lgsZpMbbu48jblSZJo8gAr0I1jN5M
h5F2CaZGgCJ+tgSIIEXgBDWMWeJFTCsK8WmEq+R2Te6gxALDKPj8PWp3Hr8ja+Q0
Ook1uLyC1B7YFVkj49WylFJqG9PhCRVsDUnGUL3OMgurszprh+jwgnynHOlVfUn0
Pfwz+3+FRfxLpSYzZZz2zskPEtPFgqBd+SRvg7YAfGI/nPy8/4pyjTx7hbL/4oVU
fa3gp+egPB6r8Yu4IPYtgfESzxHFxGrISJvdEs3+rSHcNzK9e8pEj5OdqVvxuNyQ
cz+CDkcCY0eXLonlrAjKrOmAFnGYHrZzrzo0rAilX2NsTYYyIKy/ISPGtYBq2j5V
KBkhc8KG/yempIJHtJIhpOq99JqTW0MbTf/nmmgSkSwMPfSjFjrArBXQgUxB+7iT
T23VBr+s/53hDVYaEaM1H1+IESSzJOEmjEkwu+IRCVRRQ+MAaO0z3Pmzs67lelLF
E8vwM4vM8g5L/NVd4GEj8GvvShAPRq7Sga0nf4pDXqA1MT4UwtIPyIvk0MpwpnL2
07/D9VRBfieGeO0i8fAgdb/woCDxVQoB+F4bAqXqujYQfVRLH1uJMI3wqjLc9NDx
OK/nJVF1nBnXdXxKDLjdbA3TIMtRY3vyLTBZ9mNow3Jw8kOZ1Em/oAQdVJor/Kjt
smwQXmkB563sd7/8I/mW+5qTYf3AuXZHyaakbB1PaJJxmA2RMNJgNHiMTyVb0Blh
RXq0PrU8fuD1dkbm2YA2r3JdhiUhjcolTn/BCRkMIeA14GoEGQA6LOezuVYlx9zP
tVw3MMKFChetc+TZClkU7RlHopGhLVrUdaVJ1twz+U8hEpIEeTWCEbJ2i5ADTyk5
71YFalYOJ84qP8iZtXsSgAtRv3C4jErbKBfVHZAVH8YjV1mhp1U5zWDYluRQBT9r
riYJhML4rD5dVzwu/xczo/6l8IGkTLYUvaOnG4d6Qja9DR8AndkzR1ibyAeDYe4o
OdC++HJFaPEezfbM3uWtPYmtkHWS0ZOZJaGARkne1S0twbQPYLA+wlwZuTOtIGbW
oN1Z6e81fNQwP8m1gL3mlCbsCv1B56mEq153+cm4u9mCbXP5/JgFPnMsJgmYjBHS
dXgdiaNijA7WE3pah0p6FcGPoRpUHm7hu7Aj+wtUqFVPkoPQ/J/JVhk1gn2w2+zd
z1ZmuogSZjF7Zomo1uTIyYbZqRoToll3iKzls3k7vAnbGnEFgbRHX1t/xvkPKNhT
P0PF/6vRY8YcUE9gCzM4+H9rQ/GpPGvGz9rNs9kUwojZF3jMs2QRq7eqFlUFFZwR
BSe47nEp/bttuLpSlWDrGd1UTj/N0/VgyOH8zTGYU1oxXX5GHopmhz907RovBk5z
O8Nf/UNxJ6pz6l5uVxYnN+hSiicxsuIO6yk6it1FAURliLqE3Uqr+kuaaxHj0mTn
GMWAPy1kJKXXXNfg/VMwXOcq47UEK1toqHU+9tv8oaMSeYNDI89WKYq488m41YzO
KV50ZTenNl98Y3nvh8OIjPl5o0OYCmSrLj4TjI3Volh+DlpydcRsgDrtX/Fg7gZQ
W/TSwe+vFDrwDiHRGfkb6qzz3MaAsKP34kLHWwSYHfZYbfpfqJ2leZOaZC0d7c5V
3iGq9pW3zac4Bw5qMYiPC2F8ilw0Fg45G+nR0tv3jDsgBZ46UKARSvsujgUNkg6H
tSx6cRZfBgt7Gx0niP2IwVw3gKbEUZ+2ZFR/jr3pK+x5PkS/HqhsCq0kSMCetgy/
VfoEGei+RP3Of4IzMGt+HT2Rgw72mMcV0TzY6TMjsHJ0bkO0mu4WcjkBlLwx0Gs1
t9CXg0/z5qQY5y0GHJMmvfumCVB8pMrR64zM5ozAzCry6b95jv9/p0dpcmbCS0/k
sgCd40hnMRNMVPKvZowPNpS8tGTVOTzrxehJPRtkJ5f7d9iDrBVSO1vqogrv/VlS
4VXUdeNxrzGDJu1113QX1vuzJ5hOGMvbL65T/ihxMEcgMomldMTaUHbACdU6g5y1
qoEfx3LeoPXn7a+m6gUIGtyHvO1yxIU6dMO0GC6tFAI+LdJgRv3iRmIVpPx757b2
9doLhLk7BF9tzSdh+rtVVV/PZEecqZLD+S68SwkP4IVc0hyeY1K8aCkaUyIf9X1q
D31BtyjFi4WUX1mlTYJM+Fl7BHkHSfHBpIf0mdq4CD73bRgLdZP2LOJcR3+X4IN+
b2JGSqogHGGRpOnxhdUDmRcREgRTL7mdkmxzYsNQwXB3BWrE2E4WhVkyLxrS+MiX
sB4hsQ5jcbTfGa71Abbj9u9zY1lPXWUIKCoQfI/TH2Ai5u9fCnMmF+PMrVQtscaN
WnjSWstyoCSnnbdKd6gAAccjLNIBe7bhBIp8S0tShypwD50zB1Cr/xFiJLOYph38
C6n6wXlsu7aazy15rSjGgTk4r+XjoupF298/HJ0a8IhS1nEmx0bMz2194W21vZ0D
JJXPuYgzebQXk3EQjH3QRYzvboJXlasseHG9qBIGDc1drTcl8HmN0yaaZkxclIGc
jfQsheHuN3BSCi4FgUwT4S0Db7RAFR/U+EQq8GRT7Aty9Wzm4OYC2ivcILKjbyUw
ZtvMvDO07ID4D/o52G+egCHIfPgQFjEquEAG4TVtqSeZWp9wFgZkgYNEc22YXfxY
l7l0JxJjYaEQJlTF27L3GYX1aOw4d7qpiY2jHBSSw2MeCGXzIgxXC6YlP5yYcSM+
vrLVlfXqLh77losNCwY9ebKbnZmx1pbUAD+6b/6xkgJFzndqJYegQIWTnbCIOr/e
n/Gv7MY7PBQXN+PO+jLTu0abVy9WJuW6rQiir62qeHJAXtmNlddZrAw3uwMoKrFk
GuTTXJ8nTCZgmMeI1HD3Bmh/L2aellxCnNFhELsNisNa13jD4BYTvGDSVDCKMieD
RJ9yqen/8eB0pe+muuVhyfRl4Kcmbh+kl7o9+rOVSSp1Vv1T7vnhSc7Jfa0m5QNL
unVJEGbUDskB6NvTQLHcYAa4Lw8cNnB9el7K6HwLLDOeXHBm5mz3PpJjlDJtwfTb
BgzFSHXJgb1RI4pMrOQyogAq81XoONNx7n9ko2lBGBRSNm4qYO27dtgXv7zHebPh
llF5c2p+a8NK0US1hxtHsHKZgtgDGzL5IMRadW5fdaCAnjTSl1dR/gTHM9VQYR/5
qPPlef2qEctYAcud3/0hogq0Uv+6s98wr77taDtaB2dET7Reol/Ti+2AQscNm74r
Uj/zuHDfd3bFgb/aNvHGfFyq5vrUA5H+6XREfEuBCgEQ7VlMNn5IbwlRMwT8JAjx
IV3jCbqaFLrubWtXYyM0CRU0k8UjXZgqUNXriuDigE0wA2NOii0Xq+prEOFG9eNE
MtLYK+GfxWmkcBiu4+wvoJQ/2mZ5PwIc4IhJP7onfR8EReZ9j4ba8FE/cirP/JBT
s2uW7SSyGGfJm9EBNq+UPEqYIRAM0ejFQTXee++FJs3rtjbnqG9/V804YE2zC8Zn
hlBfX35JosKQiUzDtDLHf8SW444OjS2DqOCT+o2cHGXhAent+pGTAzdMy8fsGae+
cZdU6sOsZxTQpx8Ypw2KLjTYaF4CuPUj9jlqgKCp1ppM2nxJJI+P4OzmvBqg8mZC
bXeZkexJJNf9t0XNvyCAkbaRE2dKv92bWlVe5atSLhFF9lp43zs6W0e/1YaQTTd/
ZNwbnJ9mWlrr3sMzaU8VUNjV+Nhqx4Ee/WNtk4vAwByKXX2wjGpt/gv1sTOCfGMh
dhWJ+eQ2Yh/pNcss9/3nWDJ6ITjyaVCvVpEZlFQMnDhfIzQhlU/ctVykkNMwYaEm
DH515llucPjQEJgH0kXVq4xuxpGOWGrIgiQ01/qpLt59EjGNoWakg5e2fm2uXd3r
2BlO9OxZZSI9k26kW8FIfF8QvAErtKoJdFhrtaqOXDQ+haD/lvN14onJp2Kq6uvh
6eD7xYpGaDjlAVnTVC57GnpFNagf8/5MQhTVLbnvODu/KGocHoP7l51Xj8C6Dpq6
A3ABVBeohaP2sX9I5EC5puULOi7x87TBWPew02BnAcr/nvWFxtZkR5U/+R4jgWIY
ITL2WE8sJBH7GtRWuQklQgLtnywTFqPHBtlmOFrpbtcyU/o6dHvFt2JVsqA0uUDq
i5Afx7rYDyxkqKXIdsPvB5H0s2WdzqHoG16Oqe0ln2vyZTVqFcxwNvr8r+n9Ciia
R1aprGfTz5xAMltG2v714fr0PMHZG/WFuqrKuWbac7SF1nf9NsUOhT1aHVRN4k1V
RBZoUcxVZpE1hLusv2JstZ1RCHht6jX8MYz6RR7O4JgIMJG9yZjC7Kv9E2n99LUw
nVk24w5+Ti6E59UlKm6LAnyElpP/r2WzCg1JN84rSvxJVSAYcT1oWvkCAqs0AlO8
X22Oyb9qf0d7ThFhqY04LFoieAXRE8vB3KaKPwk5g0r9AxdCUduZTz4trHOtyC05
Q0UNGL66mEn1rYCYiP7zeAorjg1CKXdQJ5Si94c9a/wsWfnlJgvxK2xvaK/7FCTd
IyT8PtuCR+WCBjglxSfLFeWBWAyCqAFRFLq16iFD/2RAruyIvTu2fSVC+kSmFIOD
v0rjxaU28z96y/SWJCS0y9xGE1VVpiQUH45Dqio1ibyksxCcS5c8YO9Q93uvIB6y
9N8wrFepM8S9S7Sm8honkJnFSAv6rIJnhmPOqGIBLKyN9V+uO787AxdbtGtVACzq
cQ95PTFcMs7XZC83CzJXHWgEIWkyDkWXafXv0JWJhrdrYyCDHD+Mg4dEuhAC82AK
jILLPc+qEhCfxaTMYR3eWQc90JEEqivXvFvRx4o8YD2RZeCASdno4h6WNucEzHPA
lUsEDVn4P7PPdBdkZtltcFfAvGxnsl3m/YR39l6pFm3+y5ZjbpQBprm93DKS6vpc
pldvVOaWkR1dXMjwNEdOHgNesIYE8mxPJ49OMdNMaQj9I28TuJUfnJkTMshLk7Et
XL5EWrUzOkKtY7IP+9drpbidT0hFyRUUy/s6v5KwK4YEfQbR5jmK43b0y832/XBN
U4a6sssWbn8IVq4p2qgA1gL7whG7hRlmcCyrLuBNgM+uTqZsL3sq+c6dvpqbBLvI
cmPC2m8aFPPxHuFz7P3GdOy2Y++2c3sqZW1jnpBCKR0YArxVvXntmQRzc6i29BMe
kwSa9an3CWWCNojoWUx6IohXUDyGCAsQAbZ4ImE6VTCMB2QfUxTelNU1muqOOwb0
m5dcfS/hRsclkhSdblIzI8WmUA0yR0HeaE3SliCUaacZDjVz77e9LL8IW1sDDQFg
3UTIaw0/ay1Eqho4dBpN/JEnLh9NMeismY0AlqkCKsVXwRAqVGPbRLr2bxGQmz1J
bvnA9nVcrQ/i1IP4i2N2d3H5OVgoL6b7tDvUos527ughzI4cTITbj+xQYIVXOtap
zGLU4DY8O+nZHKlNPlf6/A+h7iieWxsX2nmdq53XpWsO+nRXDSjUSQBLfBsYozms
jON/WaemKVMzDSj08wuxs/sJ0Uh4KdcHG86piuG+bDAVaFq7wFw1IJx2I/BfVMsT
44YLx/DFQwSlh1v1z1ATeeCEhNnvwR27ldDTxshIauPu65oyZI60ay/GopyogWQz
cq0ICW1OmwZu9MF1ovxrvOAOp5EijJ+3mba4T3y3hJdzOIzdiEeSvMnjeJjCqMF3
FkA7jUOOfE+/g4kh7ir1ujKRuO0kGGrJ5aWNkAbj4g8HfwZoKFCoS9oAFllX0Uyu
Nqbm6Q49Sk+jLoiYyQdE2HV/Yw2kTXMRpzwyOnA31f/CcVBXKJJ537GMoRIWJBTf
UZdCeaFedBDNnxyc6b0OQOZn8DeSFY803ptA0YzLtP055UHi0Aa2hLf45IvX5rTW
VqUTGC7khub7VM5XD9ct1dW8d0NbKE6urcn44ynEujEen0SrzTMiqjonw//631u/
hsYnxu0ClnRRRiOR8853kZH+ult0OvcbU2ePWRzOcGb/MI5boE+cshtOnrfgB12T
Nuq40yK81L/XDgbdcLTvVrHuHJ+Ev8a8VbB8ji4p7UKZDOvBhIX3d2Z4kiz2HOMh
LumdZL9koamt7hUCSJAx7JLp0G8alHl9qxhsV001xt+ncCFGrNzf5S0QmiYhvQzz
Bq3QI1MNNJTYwjo1IDt3NEcJKFaas9MaCS3K2vQy6luFSUdRIKQb3C3AYsuxSHEq
rNMfDgfPqMk9/8zqf6h/2Ov0UETrq2+eAPesaxrUc/la1no92947l2bqX8vWAQ/S
bsVta/WxJQAvHUv/+grDNQ7N/fW0CiBI9ZgKtQWeD3efsKdKIjwe8arIIl4UN5Fc
P+rMpBmgCL5K4WGoiHVC/G+1w9GcxJe/C46qChjOMZ+Z43amkxdEQYgy6RQygHl/
+Oz47KG4UXWt1II+nGtxtYJqq7sypRFHOC7LYbYyEMybw348huyr+hiisfcSrXxe
WyYUv5Kn7pGnWiYgSndGUyyHPHTXGrB6Y9y7hKeks/6EvB4bLll9B0O7NZWoZqVJ
T+teijR6blXctfBBq8tUp2HenmET7tA7TZ+E03iBy/VMtNqhCb8QXRIBFFrEyD3o
I+5gxSVl5AaU/PS8953q3g1eJHyFS1ZcypRWsJF/8mwizJqIrwKKQI0+cWqlG/W6
GdwYV63+yM7+WIAOqSVZmNS9gBFKG/rBYaa/VW3DuyJ9sCwtyuimov+snDfwGtVu
yu4BHdVFWcELHGi+8yJPLxKme7htkQ2ET4OxK2r4F0fqGkbPsUdBKlFWKRV7ox73
XTbajjoyc5q3+jMwmqUh4RviqS8xyeFcA/jjnYPB+Yf/aK5QLOyhqa7yR8spdheA
3L62g51wrsuIhO79fH+ffIVeHRDkKlkwjKBDxGURk3arbqz22IEBNmIl56FLAK8T
EzTy2fVNuH4Nr3uqn1+dcKW3pkV0BgLMlQ9RO3Hzme+c9qr03P67kWhHvVzWEp6R
+pOiShdW63DAtX3wveBFAtIQrsjWLvi0VQjRH6qoXRUDj+f4EWwZL+F7SR/aW2Bs
EAMNF7lSYfUkav5GSmmIA8YRWzNzOAqOp6RFQSv8SlF7Zamjsj7LW2JXk7t043Bm
ebkj18gTfpZtl8aOtKrO5lZpgytVOL+h1yZ/O95JOTXub4jIApD/z6LD91kNXYFd
XHw3WYF0lwTHB7Qjb5T0i3JAugWguOZAbcbewolzNTu/Uz52eOmT3NZOFmA/kigX
DqvS3JkkNsynLgzfO4IYGo14IiGj7BdknsvcLgqMGOd9kWi+PARMg5FkNpdD2Xmz
TgqGpssAq7HFmfxCkU8T1gHubZbGirmB1hIzN0nqHxV/y6sGD7HhFzuXkabyt5C5
Z0wPOplEaxDmgIp4P8eJjsqHHv4SZ5IsWBdgzyxk7qWH87GTIfWtVE+d2tMunucc
xRU94+9Giu0CKdrxErGTwJtsb0tFLw3PpZxu92bUEU7pVZ0ZgDipPUGfnpUYQj6t
XhKEx84WtTdcGHY0NI1pklM7gWRNPNoniX9yv7zYLv5tGGPATF2rYZuAvmPig/Ep
3uQ7bZnF0CG7LK1CzqOKY+h7Lx0rduUfPMp1ZkVgZxkFI9Kd9n9JiwwANUZTGa1u
b2pOzYr3yQWg8YPM3BiIZfUTD8O3rmnfWCyirqykOXf7iMSmoATOcc9YNUZd22YV
Mv5lde4gfFwrvnFv8SqgI5KALgoRfVJr9+0xj/LFYP5MWmqZ2mNjfXpCpYU7ES9c
nnKTErOCI2KtGcNUdudhYGpEH1FmUAcHTLA4lvVtoO8uBWyR/hnafPGSKM2Hz0e9
CSFQojU2Y6KfH1BP5Hd3sje3cJG6rCjAOySShWZyiCVKHBP/uUdo8m8+IgdHOkwE
l52olJP/gVmNHx1FevdPLInRoHDlEvN/6Loz4t/nl/6OruhX2TV3QDavKyM7eAGZ
A1K1eL0Hd4gk8wQbAVG5HHFsK2RBF4a+kEex8qyoI0AABPW656RzPQEhvq71UMv1
rPEMvMuMfbzXKsBjM0CoxQDB3fQi37YsMezscMtJLRQnBZxexBmnkDjhVBkRc8rh
sMU2VTIKAEf55sIZI42xKGxlQ4CQGH3J1nj2cIQ0ochMHJ+tmZC252WdigrfN/bC
+8K7oWPfg5j/7xmAUyC41083H2LaVWBCiKATJsfTD36Qhgo5f2ux2f+SyoaLcM0X
UpTEzfMchOpGGeDDVAEMr2axoyQEr7ie51voRobNY477R4G+IbovVOU9CA4amOp/
Ts2qqPQmH5k113G1O4xcNPBsUmAynCZvYcJ+CeBG8qg7E2QpFBfgzEUKcx4JpV+s
9donNmKrq+WoJn7QSQCb+LfBx1phedD4hkG1oxwCqOrvYF7EoBPKKflBNZj6Pi3b
RJbUMyXfvSZvohMjL9lGQqx3U49sMIMaRlv+TgPo6hWXl/6L4CVubYmLJYLrfC9H
cqrZhhMqBgS+A5MmLPhRFuZFCgB+VuxiSZbz+VIsBy2/4MxnumzQToriCgWJOqrp
RbibvBGig6ytg9DLCsTAXP6AXEfPGgP1yYUaH4pMqT98T/tQuEO7CVey7VxfeRBB
2an0XvQ85vTZa0BUZQqxoapyX/CszDjj2PSgDY8dCIQOS+8B5rW6YHsbQe50oT5s
KhiYgsKVsx5+AcrKktAg77x9WarYqhK+frY6shjqjKEuUsvPC0j1IgHuMsd34pOx
DQa4u4zKe71ccTorNY27/WkgxfMws+ncVlq+lPUppTz2LEHX/lnJlasP+W8ylEZ8
wuqstfnaX0MHpC2c2PVJBOObLPgCzm8XP9m0Hvzp5K5JwpbVnZcFV8Yob4WqSwUZ
6aoQQqEGZHq3B0eyqzqjiraEgK9V6eDzQ2FLX7+RMLAwf0d672ggHtblHzfsRmqE
SXcbW0/u5Ke+6yw/P2yd+fLrskPl8slmoQKmtuoKILwtwCzyTQtmpTIm7MpuscaS
FV4MxRNsSdZ0gpEJmQ7GQEr4ptShOdeM9z+7BkExtDFnrEc1e2KqjogN1vd0miK5
aOdDx72uyGYTP+RcPNowSsOiLC9pQ6j755rUA/Jys6My2ruKxx7GOysfA/5EhlUr
ZtczHTZwD/tglORtxcXFTx4isrlX0fXYB0x+sQM6wY/hgwk/C0o8XVry3sJM1+BX
2JSKUNnoLL7FYwT6KI+1P2ez55UoOSavCK9DCjB4qx72NyalowYx7u74h3uYtZqi
5pAR15Z29tq0SzBA9u8leXVe2izSfy6My+tbBptVnr3W4QNdx6AtqJDQCkITF6dn
g1A5MbzT3K9PlEELCPyiocu2SaNbGpaiECKAF8kri7Cxjs/Q+srunKYT6m91H73+
c1yN1JrSfGpHMSWGpi9v2ajrARo2LLceyLklM9O+pvZ+Bq5f9KrHSXy0/KzkY8a9
sRg9aceFJTYqDheX6VD42tXXLCuDKR/1D/3T+bfy6c00Xs+7WyiMlIDWXwUlI3Jx
V8q6VemFuGBULr3vbtBippvrrP6C4PXMrnmT0GnaqkQg2A1e3wsAKzk2HsNTurCF
yEI4wnKqZHwkaxvKiYOAKbMhEivsgKpi49DuDwsAQYl534hdyl1npv0bQLplAA0J
5JwLqHygqoLkN6+pYrmukLzwLeSeMsTDl19vVtahPVcr97HNNW+hFDRML16DdaBo
54k6jFF4tTqvGyxhGW4nJV2iEgsiiwrLUlzz0jZdMsGJcl+0tg5KsWvNzQ+p+FZe
CBtSCOg3kHbvNQthwNcLC0d2sCYq4Ojj7IwQUyZdqYVJgp7Vv+MDNDYvaKnP2nK0
7QEVOWxTPS28H2+iIsfaw9IVwyK9p5xlFPFF9mAJu1bGFnG1w7qYX3zdzU1lEhR5
2FH5FBIlMU7vLx5dijITXF6f3JynaSiTb1lLeuukHm0bk2Y1o5iT6jJ2SMhO+2d1
yz6sMy2+A+LagQndlvSxbx2RrP25v3evFeviQXyNwMoR6oOK1fYA6MEd5Ht2vPe/
bljPkJ/BWqZAJP6zhy5w5CpG/K1lCYwAhBiDt9r1l8uSTG0+NoxmDyhfSxcDbEEN
FqIMY45KOp1dCbDqW2E2rW2GREmoBvZ63dzX4FmkKO7OtKISNn9NhyYNAglgX7E3
Yj5ZKXsv3KgaHm+tmbJ6hgibl50efpgJC9QBhNbUyQVku5glL3jnssTbs+SKqtM/
LeL5xLTRcvvwXPdO6AZLx5bMtzgAIjTrruZCW5tpq10Hmws1aPJW3NYNtsbBE9Hn
7fPaKtulI8vSRM+hafbB1Rsvxa4dxp2+jHSafNa4igNQWEubSrZ9N3lJ5f+WkarD
CNuAZqqhrhI+PTSc4a34UQogFFzJEC4faqyDVoeh5OzK1znSoIZsrAqfP4BXD+AI
Fp4aL5BrQFbTK7G/q2pkKSGufJJ685Ij4bh7S8VoOQq9JCjiGTPkylWrS3V2I/WF
w/uSr1/fntXgeIo/KiXezVlAF0B1KTdF3Y8eY3MkYIpc/gEy8YkaOk4ZgqMZ/jbR
Wi1Whz42lYWxUdplldF+EHf2FdFfqOVDu7PT/4A0LspmWEP7XMCtYpyv8vLLsjHd
GOZ1DhLB3tLA4ew5HbGKRtEQaUuoa9Ih971VNiARvILw9yc2cmrm32RwEm2RTINI
krnww+qlWrN7RR8iekjwEXnSCyLAAT4RyJcf5Ww7qXcMtolG+Kf3K0BVOYG/PkMF
dwwiwCCSHCnve5rh7ESGUoPxRctCWPWxa8xlhQiYM5VUT2y6GkgKZTd19o6qTFtQ
aNJ2a4l/P48qvXKRxIkbMcEnJnfNdgrvZKdbWyvGe0Lv+7KlEZHebUcVE8rf1hcy
KqiBYcNdVrbai4SyS3660281mmY3oMWKSXTP2DH1ktHVN+lVIgmogtbktoi9kTtA
UhM3a9Gyxzhg7aDpAuKrstjx27kRZXjlLzphSNM2tVtfbVs4Fqy2gbIBGKVW1B9U
u88CdVm6DcpeF8+656WHIunZgkoJlthAo8tnJ7KvqIxwdP5uH6B4Qo+O88q8CvM/
wjNn0FZmLzn3v5rXi7gNH6bvbicSYz1NmIYvxXMORN2Rz4qUmXRVDIBt9XjsXEMY
oVR1nvhd+X5rvA4xq1Evhd9L621kZvDWz/EM0sqjWF2zKFy9pjPp0AsaIU21VpXs
wePhNZUVp56vs8h9l6hd72zZ5oUHcTLbQOQJ1Efmw0afM+l+0ri/+8vAgHvEDblj
GNYb3iPx6t0roNDwLGrXIrO0bk6TU1tpRZaWHJSp+opiI9G8AJvU7JV93n97Qt8d
5ASDc0T8gG6uo9GJByB+M/O1cjSaL0tYZWN+Sr3zJL9ln+0pl4KmU/Gr/d5Xt7UW
au+xAlePx25dAxil0VzzTJhItXRlN/plYhk2EkHOrKKLetoEm1NP5EiZ7810Wq7W
cUa+PptXTjRGi8sgDkgqFfGSvmwc/+yY4WnXWSDKd6Jq1rp4rM2xqcY7K8vaNIkI
Dp5bKc3jcLrsywosg0lA3gRjDTUyhC6Ft7uQiGYaxzNSm8BU7bP01lnDEpNutmqm
sC70auLOnPvquLkfRZGLX4e5ykyWCorkpxu7xFejep9JiKZi6CITnLR/y80+e6Jf
2je+15CEfA9Udv55QuVookmV/iN+aRyYd4dOqMw8Fm9xKHI5vYsfzdhCvzoWH+aU
mo8sIil8qUDrQjES/yTiuej+y/CKvXn3vEXFSleTbU6jVXcMeasLj/3u0orQUA0b
xGOxfrkqEg6ikY7PaPACj1u3AzwOQ6JcYPG4imhthCtnnStYDcORmY0eY90KswCU
oTpfdSvwK6owaiRrtZLMZB0koT6h+N3Wh0qCXoRrYp0ZpjFob7rTE5SiPK+HLI1o
1coWWuj3hYAIsqfoj2IGkhRhjFRci87fZUZE0GrQOGeLjB6gR86X4Wmu92as+H/M
XqAuh1o7hgGwqBsWp0OFefH18ZFIuoaF+1FO0/hpygOJcuFELXeVLQslCACo7/FM
Q4FnnOFcvW8uHkW0wo0Y3XKPV/emDYMIfTRfnzDTBu5miIvML2RD/YgkSyatFcAS
H5QVk/sVn06SRAzP6c3UgpoxbGOnMzoPYMiLOZleq8FDmHz7WDZxieUoxC+/ahAD
XH1OCMqe7moB7hT/6ZBkQXbF0lYfOfHbH2JQymmWPBGaEEGJpm1oV/f74yd9vWcO
fW4KHJXlF5Mj/+ry6vxCC2qLJfGXDwc/RUSDkBh3ZLV7TSwIGsjjEIhKI9Ge4kqd
8Z8vaOkst0U4sgvxR3P1xvNtiPpNsnZRgfzkZ8BWSNGrS/VRdixU+IiG1nzXbCJg
2f7ZPdLPAEaQV7q+FsjYnDU4a2OBP6VAPVKQnVGvjkgdrvAvceS9ALSjm6D1YPQU
QuCCMxFeDKrU7AK92lGQdDVMJA14VcX154UvrNpLES+ncnCZnOCvEFgTsnAYjgnl
kJMSs3fGbc8UOJGtRvOwH8Q3GqOacJzD6eh0hWpOHKs1ePDm5yKd6gs5aHdMoZnT
uBhnOyYdDtAhrDKOiyeiSG4icfQYE1QXV/RVZABlZc3OtQCGmSRg8HVw9MiiSCK4
Pon3xfqEgplfR2tWMXGMjhZzAqOM6ughZFU8xmL9pqwAV26ZB+69Ukq1GRGZWpmH
XCvfkMWyqDGifUNVYsCgsfsgUlr/cD3aSGFS6SvclS8p+Ef3JvBBaMA4xk6m0pm/
PSC1pCBh4YtzQTyKyjjnuQCIZrV9CY4PmB9ea5rWDWVWIVJhmD8yRcil7ddBh13R
KDL5h48tNKSF1XwIpQD2fo0VTqNWO6hDhm6kYzCPwyagbP8mrwfzXeIrO6WYv/g7
MB3BxnGHavyFrGbh9Abg529htnLMoTAUxODMHHPdsm6c0Z5g2P3EJnxxG7j6SZ86
5e6VgwK+jZb9fEFALCOUrIpPdxYk/tV0EHictZPv4HINYjaStUDu2BJEl+qsL45y
A44om6ekRd2ClLsWa+pB/Y3h/+rW2oRs3YviapBimM0XGnYcvUUIAS/KF6FPsHlE
bss+k9qVK7NnED9czsGWwoQ8Wq4QhBc4fPWuHaMB5sE6Twd25oVOgZK8S60hXREm
xlndOhaaFTJgIoAn32hto1aSiP83wBnxwpQdVh+LJkGaV1R1qvSacjJ3nfDJFYQ/
5kbiX45Sl4nsNKr948D9yzk8p6Jbr1HUMB7aVFRdwZ6vDhwaAnN874oSc0NFaJXJ
EziqqCdHa5knmcXtaBU7ngByu5doUHopkv60I9QJjXewuo4CHOq3n4lCsRAn0owt
v4YsPE7vY17WOMP+pm792iuZfKK5roLk30y0zaglXPiBE0ELl3cWHgcCsg8r3D1g
xVPVgRHwsIU+c1cd2L2l/qpcXaTcfQEIenM8dTg4m4vX5ug2xKd/mQHFKGUtGM4n
7VQlDuOMgsY22C8IQv6+8MNat3lthjHIMqvsFUHog/66bbprInW5Xnrbtv6yS782
QUmJc+/9WG9lnYQt49a9lS4KmVwQplD3o00W5RwUDnufRViYgGMN0DugMrZnZcvn
ofNWR7d5Op9MQWllpmzw3jsfy1axcYLzjszZqsy2AO/lNC5EfjXBhGmvxqO453Fb
DrokFToQOn1K7fARJchRvV7UZ0kFwg5lrOfAnDsopxKb9ui3ik2U9y4uf8rA3oOz
3PZ/6f7ffo9aoGYZqKbGJeWFR+nrPkDPY9bzEhn0GNMZmYRjYdxZ+P6F5Ry/MGx7
+G17bMJL73ayzMwvtw+AGs7BwdbHGP9LleIdGbpow9ZLUVWqSX+hWsITJXdktl9G
2174sbZMQY/5uhKn22StOSVUHCBx3FM/oitMv1tm/Ue6fOSnHGZULTd0uaCDHbQ1
qPhekd7L+1a8TYUQph05gX+1d3fdcuMJKJ3m5UBUYSj34Sb1u06WidlMxKB4i9Ro
f1kO4vIwayDF/wcc2mbu759hf2yMq4WkIaEqluQ7Mew+oeBa+c9ds2FPTv/PywDy
sSFBCwHEA2zC/p22iCtKxtF+rYueOu0wibiejeLy29Jz6UDVHKAgMqXAFcLnRcGE
Fzvr0wMwgXuSzGrHGXyWiGVzHwjoaIcfj8yYMfw34BMWHGaTKolqyxl61HgehiIs
tXzBg0YYDFJU2NGdwQmm+EEMjsAzTwa/zmENNIcDrImsaMzJCcPqrHUDoT8BRM3G
OfpDOFNeuVRgnnjg7ecp00dguNrD9IE2m3smuMnoIemtXS/JDDLvsGKBdx5DhD2f
r99LlNWRQoMUy9wRW4QtxSpHREOnyScRv6Rx1TFtEzD927hO/ElMEyC0lkF9QFw3
VLnG/+qtDUX97/r23KncnoZzagF71N9bHzwItDRgAMQcR1NDYBi4Joa5OH/mXalC
DWeeiXzlTKI/7Ylf8+ZaOxILLYi/JEYYxDCcqje1XL0FUOJJOK0eshaNQQxlNaV2
rSqRNIr8IAYDTUNbbTqsgsbCXcZGsn3+kFbFmyVk5m1yKob3ewtcm1MUC03tHdAg
5M8JP5pEqAsBbTFboltTxBfoakCmlAsFjc/fvMuvOXdX1YFx2kUOrDb/8wFRgPF2
qbjLQ3Ox0l+E4VCJMs/EJ6uTllNb8zvDRRZTPe6mqG1o0V5rxepemfc3dsY4Wu6S
4i4GilJgR/ncOYgWsDHCXmDJPwyre41Q8y1VKpe4expGHDTVOrs0pjLObRpHJ1tj
xTeYBGJjhT3HyA4CeTvk1jsRKDHIXAvjapBgkxctwd5aWuhoxrAaJBisFY8Go2Pf
qx/idGNRLUDf+3MH5OBa/Zlf3Bdlimp5ba3L0ZviKevVyut01IcWpNfI+IlruNRv
KaNPka6+5XY29K22MCcFeoTTkcSmfW5XqXW2R/7RuzeEWN8aDHoc8k+HGPt4Twmy
sJnHp63QX4nGmYGo7cugoW2gtgc0ZmR1sdLZYsMMpsljrGmImsrf/zi5Mn7XlwCE
KFP4/mcztFV0V9FzsFMtCv7apqNZsPIOigJvrbbpvV+U3dmJ6wXMqR4+RNYg5Hyk
VpbKyfDmwIdjkjkN68818PPtThcykOWYWw0yj3y30tZJjV/OpX+ualvxlKFFQbqI
zdWz7Q5gtBn8Ktq8b26VAHWhKsFCi3umL8vJN/njcXoAUBIzuSo0IxH7pgK7y6WI
2sWJcXL1VWyTavlJwvzIpT7xSnl/7bpxHBqMGRaG7ZJZqssI/bcI1QSz5vVSLHmE
Ps/Dzn/H8Vn0JaxqEX9El96i+ZIxqszRLUWYCXj0JVH8sg81MkZEULYGnR76lEdz
8ojG/lZNGskKLgDpaB2kebcwoHkDWjYQ4lTXFeYpxZCo2TltgOPz+H2YuR532l9F
KwjfCpkgLPZFwYWriiDhch/c/TYDA+FFUAUop/Y5dz4gaS4C4jGHwYttozNtMUss
DOa7KLEwLFD+omk4HZ2Y33R30ibIRs+8FZGNea4TCwgtMf7QUsdl63Gjybrbmeo5
sC03JyabgazYBUjGmQuPD5EF3hlcCOx6681637xr5ZJN9izt60ep42AYTNsuj9nE
ghY8wJUYSQ+Q/eb64wgQlQSETcZjkP64hlfAMiM5lD2xjbnaTGE+XpWR5yp/JhW6
MPQdaiUDdkyGPODVC9bL9KVThGrGR3MQ0HbInTTZaNZNI70dFVoypl60TmzaLuc6
1nh58pA+cWh8QHplwTWB69oddc9UuJ3MNZoXUBPFKCl6KbeC4Ntfw0L77dkUxATj
sCCp7JU4yqqgO7kaF9asxDt9K/fOuqkOv1/XI1CF3r3ujbF5tchfq1o6h94BCRdh
UZWdWl86aHfGRWy5qWL1duQETybOcXDgg51bH12sLTNMD74eD3LXxWp/AmdKEcMe
w+Tt1ruojlDbXN1PHViIhBnzPk6nkBPAOKfcgH/Cs8lhAFdN+60jCTxj4eMZSPKh
WuVR+XPbWj0nmQlbqj5jrrKetUcz0cZrjY9ItNZclu5yM4dn8KEglAWVc+3r5Na+
QYXkw09v4qtrrunaphI1v8p6JMg+AvRQgVcRuCQM+0JW3qL/mXpmD5K+4ydu+KIc
6AAh/j/Uka/GuonXgP7y/IrCGqWpKhaRKwqIf6VmqW4sRCEWNAsXePDY4iCNDsUm
CeW0FJQIASnUEZK7u9q/4+nmMMmtafYtIqUcPSXo2J5/ab0v02DtkLbV1QAcb6e/
K2h95HUP9be0LCBgdw204Na4yw7s18wKKVgxsQnFra1Poac1Eep/caOV3keqkrJU
8WcVLdh9TGhN93ITC9mfPV7ejA7HKBhBInUmvhD2cFSfw/XokIK3sWZRkEHjTCot
O+FvfGYPw4nP6YVL5hclJ+Uv01/cZynvfpiDXT4C+sJq8TXLmJ8H1jgKwaYIR0VK
TpKUNyHRYrhzFvT6uThQdy5d7LdoV8p3dIIu2E2WBsMoZ4O2kjoCVm26HgJHUmBw
wu3b2aES3bzOqBpjI0QTLJM9jWGY4UDGFVZUpAy131GY6HM1ThB6BZT55u5H1ZpP
aKWP61/rOiB9jYVOEsRUo3ULHRlkpVeiDw6MoOpO2EknnHjka2IiFVmOl9QXAhdq
jmdr0hmPSwZpTCPPcOh/V5+mt1keATHRoj9vqbkk1H3rlDfu4OwzUyRa6ObF/n1Y
2nmJ66eG1VyXZJByfEpx2C+xHXYpkKM2/B28KJCziAAMAs7vbbJMUT8gI4JcLH/A
8f+cVdFuyJQbzFPiprkLtlH9hGnJaIptsdneceISqsPZLoQ6hqnu1YWPNu359pAH
xbx0720O8OnYTJrQCAeQ0wZ460w2f+9FtZduJcrjFq3YFazzzVUISLZ8IwbLeBkx
OvFVUvn3d3/77MCp3O/YU17tqlXWqkjF5CI+lYSodzlA2Bq8dXwfXpwQA8dVU/Zr
toUJzW1FLIQJU8VReQAHRTrbYuZbF49yNyPvxeAN1lKdxPLYew4ZMpo+pqkSFTjp
Yp4k2FZX1Zr+PAa6A/9FvGtS4ukhmzt0Dox9gWaNEMWnmAIqPOG3+e+CtvZw85AK
eL3tDSI6nbPkOLkvKpTMSd89Nh20sEk0Qxre6j6dCAmWyT9a/1xTp2jqNcZCiIa6
OL8wM4KBsVsmcz7KeF4mwme1t/4QRcc+C1nHIrkAtX1UeR1FxUFXCItmyhM0ZBoA
6H/fsqo4QMBbOYT7D4cqqgBbu376aruwl/plq5o8I4Xf9OtFwNPahw2S1mh2GPZ8
7sLQ42sygyfHl6f/BoUmsKT4L9ZrlgH/ElXxtqe6cl8fMAXSp86iMqyy6qBGXbeE
zBG84vZLy86hqMrSNyjrASya51Ttq89VQfVaNN/iJxL3b0D7R85H8wP64xy68hvw
qNDqstPr+bEQOyZj0e8qYAe2V96heEsWxjrOexyhpIvCFdv/Pn8oSUZTBQj34tVY
QntC65dHw0cVvyHJcO307CGkYCgtZxSpW3/Ai59Xe8bbiBlAkhGFF2Hlx3EDKDhY
Jjam8bMDEbHXiIRVRbBirYKUS/FxZcZ7Oq7zHAsBDsiDpUpPTRg5Fehpvtzn2UJb
TzYHWS0hfmEufJUAPFqDQahMUQ1dVZNNlWD3URIe/0XnPAsKTLP2MCUO2j23KWjc
Mw4VImlFgRX2SitfzZ+QGULWod5RNww+726VpjmMEIrrmUejFBjOUg7Ay99ZVxn7
5aSt6rmb0d6SNY2pXFl6jCHAchPIQ9Oj1OdNuSzqAXoSaVvJ/c3NUtZgZYvoLQEt
UOynYsPVYVIlYT71YU1io8UjTFlbufDVyzfxReRnEhEqvZs4+qSZfnF++viZGAC6
wg5Q5oELsrub3/DOIq1So8v+KLcPbFGwgV4sjLBhz7TinsGcLfH3FrN7NI7Ge+WU
2WBeKCEIZNAi/rpQvNxl6nE+Ru+ksAibP2Mwrw6P5BdAnQyqdqpp4JMwBDC0zHcr
yMhvo8DfN6elKFr4c9+vsKz+otjMZv8ez7kS0hkwwrn9SRKlPNKSnKPlEpOn7R+K
KTksZ4JzrTpLs/twQ9hL50eV+6Av5J/48DT5yFQoaCPRVT7snnqbnBWkzb3hcnMF
zNDsEIABvqwTSbBRjQN8SW8RskK4Mp3CiWcwdXpUjpofKrorFkfNFPfDSDj6wG79
iK0IhoGUiKna0mASqGTJqiGQUBwarXpLQp6x9ST/h7RkGW7CZeO9oDtCxt7eNSll
BfS7LvqE/aigZO6ibpvT/mrpiDKxjqQ3DoQN9/4+g1f6/WhtP8G6i3CMCIk6bKjS
n7xdBGkmRW9kh9IG3vndngMK7zYs0MXsfCaYB+mKAF4Zl/cHCbqYBKgq37trE6eI
sGgZ9o6en7me1mdBfVrjCbun2oSJVVD/wqo1dC+rksPQbESf3ilm+exJdIL9aqZ7
DTygsnWOP4MmT78i7TtNSGZnhixx5M5HkjDCPqsH2BlU/jHOY7kj1tPjCBrtgXNH
tjTpEiAv5ZmSs4jCFCIdFgBpI35fSocb8KFnMXApK7KX2QVqL3HsCL/HZ39qZuiL
4ZiJfYHwNnzUXh+XC7nIXWpDtKMIuxjeyv0ox1i1bX7rkfFYpLobpirIqnxlAhxy
VpfBFQZ/sGNgLnG+eAygOKLs7gd4RkyElGcQ1VIYiYxNWig5fBSfjVJ5wDZvvHtT
//06HZJqDPEivWkVMpEANG6lF9Qax4GedwwHvLYWqfXmRVZzZLyM519dgY9bCJsc
OSrUNLgwl1rHm/k8xceui7T2v1Mtqt+V9IFjb/CW9SCu2g/sB7jssFacDMEq5DOj
ahi6i7p1XTk67F6E3yx8zJ77hlJrgEdNUmbJkjtXUbijCvEAa4bMbLZcRiPGL+TC
NYA5ojNJ80Eh+VsyKkin5Ixw26H2c6OCkYBxJ6RSTT6JjKXsMJwPDSnhj5IpOSOp
S92+UPsnHCzTJIb34+shyePnYo84LXrfHleINBtZW2uUwCYBUHeIx5oEJI/zoDzV
PqtBBevepVN/3fkDVtVdKKAE82QUsVIFGeIh9lYOPp3QqxpSOxlwAfN2OXj2xymp
t+9pgkumo/NTjKCLtvjT/RJevtgTsP9czRimYC4KXDREHSLVrsI+tJkvwCXGW4LB
SsXd0CfIJCHd8Tco4oCgZTBsQb0jCcAEkykpoZGANUDelSu1qGZR3nVWpGlSqRDk
MFtYQpmeEQ8tzDqT6BfX6Um4d5LKvAhpIQhIP6EiBcdl62YvCexigQCos9KOWcPw
rIw93c0UUVYCVdq+ssB7tMCGWIML0IVYm6Ee1YdLgEeJMglmJ9fcH0rSWoPUA+aP
gyU/Nt9f7ZzwG/UPhOAlT8sDZzRWotTSLwFwixboszzSs63qwRtGNfy6J4XPKN4n
o5uUkMSO5YdCvhVpPxtRNmpCVSfrKaP+8zYLTZiukAVU9b+PM0uIKXiJCiPMWB9q
KFVczPOe9dyLQBPrxO51VCWEKjRE6/I4rpzStYKEYeu07Z1AI+nOv8nf5OilnezQ
ZY0S1ijFZv7fMj7ZMheoohjZi3+pbEupkyoGROWS09pNk6jifHwVAtJ1esDqvV2r
Hbb7Ef5s5Z2b22dw3XY9P41Mhe1glko79IDwhwvwzcyQjixmwRwj4qcrr8htFgVu
vgPAupELBHgHU3g/Qp2vDVBJnxWOyu8i4lvMNuD4u7sn1aGibG4z9xWeUAVwHRL5
u2+BtXSz7y/HJ6Zl/J2YIt/tKpJOV3V0e+svd1zCNGZScFEju+hPsan/4pumoFwR
wVzNfdipGCsVsYFroGQDH5Gf/Bfi6b6M0dxWmhLUt8IXxPIdmd3Qho5m+xuQSlu6
r/VMseAKkVjFFuXr+hp/DP/aq6TM7/qnkgwfPFOZmcp79e/2DAqZmEP5+/he0ZZM
ADJpLXBJJgTlZ5tTUvk+z76rKvao4N0ShYSbg10fnlcA6f1d/k+M1T4L/hSx/FIh
kh0sv5iEIMvV37D3jsXbMcPKhVGVOnr9XSwcT9BG/S+XqB55w7tExrbEGMsQqzXm
+EEdQI+WjlGhJQEdZkGruzxy6y9vbzJO94SOq6A5S1EziQaXu6e3GczrMLag1uij
srf6sxIMbRbQ0b438CtcZTggNfCg5D45pDYpkixWJty8h2LChIxgtELraSE76sNO
Z2CDV8BbOcpkRODr6wodcVyLCBT+x1kcMcMjo1bCtOIQXPTs4kUKC0hrnRVaxOeZ
x1+F3u0JQoNGtWBzrmh0VOdZOn7y8EqKUQMdpAw1c52+sx8Jz4zBcjhXuKGIoZjF
yxjP7tBPjdwT7edNRtNUBWIhlRB0R/ADr+agLQyqv0OJdfodDdCDx+ccmpmGtp3l
2T9NkpC2Z/kX0cEYchcPeP4GJHsUTqHTNK+agJyXmYAbKODRfIz3aEXfndpEgUHY
noGJcaTYzrgm3woSqXz/Yh66GpO+GgUui5m7Qz0J3F/tRoCg56K1f1ZRzbK9mQH6
ZrhkWOhUolYZsz6k6o0r7egSeaaXyWlXam+jrImi8HB1r4HtsQyBEOr88jrK4UJ3
ULNFdCSGhi5AMUNhjTY7AA1p9vbIazeBQT+leYchwAFQrFcUk6Z0hXdmUbeL/hmd
HiUgHuB2AVQ9GMsKvNW25ZRdhzoEuxOC7T4AWiDVKJq2HwTD+8TcrZ9CDe824OZZ
R3UWCHQcirU9hjX0foHrg1jmB2MTldsgYiCAYFcrq9dAUwE2H+xYQN8lXEG5+fkX
weO/nfU5aDF8PEB9Ggo1idMiCfWGpj3y5OlyPuEN2SuUytnJXP/oAfWxOaZM0C3u
XzAm08iXFuAa1p+zeQ7KfX7DX7uwUCvnMRn4Q+n3+fn5YAak9oYFddlUs1s8rIlk
VYYBPxhg7DYI/limHlzMDBjE3AcAkdPjwE5rb4FWOchkyNiIx/1LEc5l91Ts9bMj
rTob5Z040FrJRPXjsFau0+APufXSQAHPrnxANm+7OPabtM3QRNE4KcTCmKe/ueIB
AaOG3jVvwmEioTCtM3EVxuIz5LtJ2PZmOlw2gwz1N399R5tP8rQPiU2VgGC2T10R
+/yPiHEowyrsAle4lzuMQZ6nSFLxxvPRw3NzwQ3Zkga++PvgEJ1Sl34PpNUbBtoU
GiFgf6Oz2wuXnSAUW4NZEYIYbvK6/lcWry/CAXyKwCxfCtBo3MIU0MR8ScsgF/ig
FQjoLzeQqIxd+IYv7RWmJ7ywL13GPvOEMIykhvWYjFQ7wYhQlWDZrqMEN5M1FUyv
aJ7ZHCFNDYIoaeR9BAa/QtIy0OCFfFPUdsu7kQVaGDhteN9hA09Gg4ioS/xki7bf
25HACGAF96uSRwRUJ/7z/QZ6FYeFtVJUkJ8HPgH3Y9jX3YZFPpTYTjqt4B+itVm6
Me6qwTfRoWY447CV3t6+S6NI6jvxFqZya5b0bcuosV43MmLLwdTEyC2aWEZUrkko
w65FfFOW6Rgy2jWoT7iSb7QMPdyB6Xyrgefd4fmT7v4oaa4Yck59FLuIRLKagJIQ
jAnwRwOI2GlXaS8qAJxIwh6jvXnPCKv6EGWeRPWnjcqajwE0mvQZbsyYdqcZ/sfT
WlvO3WaX6jspsSKzDqD67icF0Mn2zk2RehHte4I+3xUbmPMw36YCteXInUGLScma
sDr91jJLl+LZJxpDq4gl96id+ba474ubHD3VRjaGR2/p2Yooa9YQmKmCtlLCMFUD
OcYDNZ7dPH0MKdARTVmOmnePyYA7MiicXb5ZgXySnhRQcwf2FHhVpRWatkrKT4Hj
+DUPSPtxkQJtef6L7Y6yhuTEVOnJXQ2BrCF3HWYSuBWhZiGBjnsgIqaSz2JAGYt6
kg56ouSteRx75QxDwEz8bv/EyLXPn8Z43q2LTQDqSTb6F6yqKUPh5tgslIsQDc0m
2Cc9ggQTUQvm9pn+BrTBnxdby3iweKRXKNB7UAJkHNwAK5jAvTquZVu38Am38EI2
HSh5hFF+NkGmlE2m6sYE2xhKj1XEGmapqBemoqAtvqX/KCqZIIJWFG1t1WkFMOM8
pwvSgu3KQzscG/NpG/iro9XwgdXI/Fr5yQFL9IUI0XvQy0EWRIOfmuXrigqZUfoJ
kXpfIdql+m+XJUNIM0mISgsnZfVZTpBAM4cD3DvCrZ2cv6R9KllxEBlhPRiChs7o
ygnTYRN9WG7RxO6eORxpwiwxWt1cf4tALphrh3Pn+YR85cma9JxJde52cTSmVfB5
LuWJSdBYnMu2ygnVY+eZDc5CRgweg5MdDNIGw9e+lIwsmQrr2oTyKeMhwLp5B0oz
B1h9G8kZCwokP6D6On7AuMly7JBkU5tWYzawFtiHMlNxY/Lg1RGbmUY0+YBuAq3Q
Uwr1jmx+5Cb+oSs9qC70I39BJFMigIyLrlU6T5Skj8Bj3Fxewu6eCiVEa4DNi6u1
P5ypRNSpYHCx2gH8mEVbzH9HLnWcQhXH6LiM5COgMX3wxtUdIbmkVp4uL9Ca1NcO
vlWPe0knWb0+fvv31yfhijjcwbqcZ5lRCpUkCviKt1oAZHC47o8VwZ73uTL/GoZD
3M01bE9npXvyRmYMvYtCsNQKBiU6kOrZ+hy7R2vPJtC4ygdTkgJa9A4X9WOYmIml
Tj0q0j3RBCNPKvohYdUftvooYC4xpWX4IAHA11vZanCJEZkqj/6vNclfxVYsvsFO
5UECYn3NqeItVbnLOWKVqAkvl4h6ESGuIugTU+cWgo5DivSST0MeV8dMpJers/8z
Op4RZiZ28MR68R5gV9JPynNYYaez+ic4ckB7SddGWej78DWJNkJgTezDV9vivaBs
riUGiN8CeHooBYyfFQDnZuUpFQj/ASFZzY3kUVL5MVexD30/wu/7Vr9+QAnuaVXe
5RHCzN/dpD9wzHWdZJIISydgj5buD2DTUaAu7dBRIiWQLJkaK1AnlHi90Z6VGBD5
67fxMqYLLP1EXu/ynq8K568PHdDmikAhEAOOUZhVEr1ynsqAkj5fqMuUOxIlFkdG
E7ukxCUs2MWo8wpezBoigvDaox17rrLqcO6H1vldHxK3RinQrztJQm3JYyiN6fvo
X9hL4Fy3Oqvs7ccWyl/dHsGsgnbWrxThznfSFT3Z619f9iliyXHEz2pc06kqLv49
qQUwyV40S78x+hawoCMJzoeJZHektL4UiGVKVEQfraJ+n/hsJRrRfPPGI6aCfGT1
KhPWs1MxgukLNbb7jM2in6PEXq8XQieAcH2ESWYua6pvOm2l3EDodaPlHonaVnFu
vgt1b0fAp/svXzYGZ9Ecw91v64AC18GMo1M4h/TKu14bBYMStt6AF+E3x7Gz6BZn
QZppH7U3j1wmMDjP2q3NZK4bB1PA2h4uYKUtwJB9HNDDGwKoX7UGJpTjy58iDNjf
C5OyEIi3vMErnFRvydiZINtr0kEpYMo9Bk+NyL79tFIXrq+3MqkqKgi/YTgdsAZ7
lAVIhmVDvQCs73pMnTnk7B4Jl+c2s18s9nGh5KhpI/DB5JsrXafZ3C4KNixDWpKn
e4aZY/Z5VfaWVoVMcu7IzvWK767jr61Tuj4ev/cgAIgoVki2OgaIl5fwcJMXYvDB
7Z9ArRhIUkEd/9hSmaXXxmlnHRRBKtMZwQ1BzZe1DrBMML6/E+NprefIKTjrh9MX
HcpRq59PsdF/wM4c93EUaw7B08zwLHSc0L0P9ummL6ypcL6cVxSuHXKKcgcmEeEv
WMDOgkNWCS8RXlGxEYVdYnjVE2mS5qYpvMsLhxZ43gneBnrOC2cFNbEOoUa1+wMV
Y8PmwhMF4JWcXw8RNeGUPwy7UncVhGpdf8iY8eRgDcmrc766jGXCs0zIWjr0RgUJ
S2FPjk/KBW3sUh6L3nupGJz0rw1MndWjXuny+dxns+T+X7Kbb5V6HnWkfSw7UA05
g/EvkfQFjK3aHBeUUk2heylY9n0VuXReC6AqgvjommMRtz4zQM+OYE98ci7A9Zbg
lODOn6aamgxsf3sFY2k0Jdd0ju7aDYKkUoDBGSc+PAkv4TMTgLFiP6WsR+tW/HPu
5dmES5S13navhVNavut1n68wi10+wgEVuQK2MSatkrzgtMwDDbhuwojpbYWIMdiL
h6v5rnegDoEtONjBAaSikufMyABPqI13zftSixKb6q9olkq4+ZgAs0xtSHTGqAQV
XCY2NEd5gAU6R9lHRXMs1RXOQ6/Iojc3aaz7rIy6AyPssIKAKqTlhjESNxuvI+uJ
YvIQj1bsoTrBy8+x+h12eIAOKXhQ4hkWptLmP8pdWdzL+hKdQqArP1sZlhl6eDSz
CS3tEcQsLWe/m9VUc65cR13V6JMj4LfLa5uT3y46Y8wzJ03cOKxsYT1PKKbqUuwa
hQlWfhUy7I79OhQYwdpCiRcmNFkaqPlzP6Iz06zFN7c4qEq2s83e10kaK/oKPDcQ
pcYHOfIbmJB3A6EmTcSWE13tx9NI/H8rKvcRWosVps6IIuIgJk1GKQRjsoxpqeDb
9v7LzKCwcnc44bpPSBKODW5c8MauNBZt/pePmht8imeqAkb8nkiNg0qOFmSE9gPP
WCEQXTfhUjRN8TSAZNJbOax5yu1CtRaAZoONkao34D3LIVRergCYQkPWkV1w1GNC
9gVymKWDyhhnjiqyHRFjQbeuITk3nEe2EbP50fXoIB61nvgUurctqNuUpmLbxS1n
gsUdf4BJXo/7/8SzKzy5hSgmjuUNPBE25QIq/0YrPG5Egu+QSMuKZrJxYGuBfIb0
srbUT1lzI50bAZRjdRb8/SjrL1YJxDIIdx6d2QqldXLNYJDPBcwK/SGuJX9TbV/8
ehbITidvvOxuDimToBV0NS0TGKbAKgodgLEHwmL+U4PFYHz9w1xIf+8acRvHc8MN
jAFGbkpHjk/KxmNOHMMVoH2IDWkZSVUfk7PyUTPrLnRUgOHg4rAAXUrub6sDFh84
3XAvcAnCqYqI8A0ChzVhn9ahGT14dfPbsdzCcv+II9MaIh9nRzt07Y6Hzmn5K6MH
AjfTc0xqyTFAbVipEJJSlsYuZ4OoaLYbuBYSpAiJvs1DtJBpZtzWu2QEEXf+z4ZX
ftBBQZ56Df6SXBFm/Yl/vfYjooi+chEwzRMlTqGmu53nVMu0SlOnpFB/8osePT/+
5VrAY7GgfnsESocV6546Ou9emTPRQAPZsRvZUNoRhjAep5P8mV0H5xypQtqI/pcr
cVgNQG3jtU/FECtGDBFZGyrK2SAKmeJhdZh77dZNCWbKL9c15xc97bFPT4u8viq3
Jqbc0ww6+COZR3YLUZmRGdINvA4oAlx8HBtY+bnjLCA94LBSxuiTDYEeaoj3s3fw
qAJlY10Zy9fAvb0DwNbkJUXqycO9piWUuiGsu9i0nOyV0RLcayO1F60uRWO8LwgH
qX5+Ls+sRFSZmSqnLKj/QBJoT/OnJ8rEqZkKf6FtVWU7PBAUoOCjTn1qdyMIVU63
n6G1TLIrizyB21ewq5XQexjLH38U0yg3WnkqTy+Ad6JCaq/CTGg2fgVxATRx+XEP
ovmmOqVpbcChcf8LkaNQNC2ozDzOpClY52AoeizSqjxzOTw+7eTbt5Lae8bafshE
VNIoJt3B6RAZ65fWL1Bwfm8y/W67Y/B9HZgBMhXY87TJkCf89QcYLgZXZ55/jhIb
lxry/g8aFoLCx+8vX72tM1e7yFylIlCY1eQ87TsFRohjqye0MQp7ym8yAVgX/uBM
Eysj44lJWPdVnXvH1C33xV12idXAFXxLvdMEPsTKJ9RH5mc0vkeFdPEHWaW1Ajbj
uLYGuXS1ZXC8CKsZTqpfTLWjO6VN73mYFf4vviHuxZbv7zP1hxZl04Tc6c/5BDax
gkl4a+HqrjygoaH02w2FzjW6vGAbD5jrKyizMTaR6WdYR71F6vYjitmnIfuqs5ie
QH6Pd410Vm9RdOc2wVf4pDsaX9EZLY5MoRa2FNaeeyv3J7rgmrxmS9XyvBSeptQC
UNJ66Q9N0rsm/S9OPAw2lp7yZ466u3N+q1o7SdOTYEdGkLANgMHPy2v5UVQHRMpd
ffC0akqkpvvPU4f85cysF4zeOBgu5WvRLYDsM++O+TGRr06CoHS1DS1+m2QpIxN1
LJjmvmV93rlhenMWtM8uA2LQBdlblaExQkKtNWeuj6uvumOlW9aHYenAg5TfnjnW
700XaYJCNhtCx65yE+n0df3C/NsM1RYdX7F6rUqsZc06rS6I0LI0S0E+0pkoUYUs
3jN5NnknCcT0t2ZVLTwwbFkTN6o2X8T/mSUaB8ikX2jK6ebBnW89eZZ4rSI4Kb7L
CrU7AiqXuG4fMbcFG726sIl7qFT61yWjTIJs6p1bQQE8nPwCagEzEBRekvCK4vIr
ZwMXVMThOni4gr7QMy4AGHTA3tQ8w15sXyP6wm4uAj7qNKB4IBI4DRCdQ38ZvqGg
Y7NlJ2P+HEd+VR7p/qgQBfosfPbYMBpw4uPF3K+fIe2zrLfDQ6HySXvbl4nwDdJu
J3H7sZ22vavzZ6Q33fJRLOUHO6QPA78+0fKuTt3v9p3Z3ibx257ogoQrAbL1P3zc
M/CZk5VMcuJ9i96Nz3zKpObEoO/qHdFFK4Go2hT8n2sp2+NzK0cGGi6tNhvmpu+s
aF4b1ncN6JaeKy59SAFIA5LKZyVbHRsJ1YDld5O/nOym5r7w+CHHXXoDE37WeeIz
dMlV9dNRrCZ6KA9iiq7T8MyREIEJSM5O1p9LafpFZ2w3nCCKmB5NYaekr3THLTOf
T2dSo6WKdAJmGyZHk2Ts3Jv0Dg96l9G9IMqG56q5tPOLmEr6GTZ8VAjjbjHRH1Bv
fVhjw+hzkF9e7u2RvHrXkP1gyvGdO/nW6lu5KUbhWHIuPnSSU0lkoLNnhs1yTOTp
zTDt5Efy+seR8d5OsI1jjkixADAKpr38C6FE+8H4aEiGKZKbKhXFEm3meo6kqg34
QiFfZE4f5JeIBmVdmo3ruAw4q7FO8Pcr+OIA9NaQVet1bOsZrAgqDPCluGWQdF+r
b2x7mqLFQ3PRMvkYpJpmkY8UByBa3PAtKm+pPU+OaKzVBHxjsNZaLNKLAARX98Kr
/pj8gCYcI229KAONVZoIeXBrqKgzNHzmfAqLhtu/z4nTdfYOg3wWpYxz68JGv0fN
F5aHy7RG+p1PX7jXw5TgvvLcdoKf3fjMWC9U+OoJ90pBV29TRJ4t0pQCwiRtHMft
Vj/wiYa2iPH2bmc04R7SwCAFelJpQ/SSsiWanZkI3N0GjUZvSkOr5nLExjmPEYPT
9IO9TdaGCXnhoZNBwTfrTHbzeXlqLR55n/LaXRyvid5BD7pJvBcoK9uXJvWbbaZq
WmsVFDf/mlwjEt3FqRaOo2yrMc0I0ZdQJYj1iWlv7Ab0+kcLumAN66t9OHQDA7/5
VtaNk/GInTJ10u3ZHtkOf9QuiQfsoK+sU2os3G0LzAymdlnFhkP892+huQoFDXad
LFo7uzeCNyGVdW1SW+ht+MKHmWrayBd+MzCIoal9GO8xdqbrk0tqe3NFmKHQt99d
HTgRw+B7+QEP0AZ/1K+EkM+6KkbRrwybMQu7OhruB//2p/s0RNjp6lpqpBPy5NOH
Pd7YuMFASSxCeL/TXGKJpPfz6fgKCm2jEWbyBIQNuWU0Ax1/tBnJScnanuABpD1g
HD/bnqIMu0BdsC5Gillmronve6pMVr/hwkcw6+96NIEWwZmgfwISXYGkt2QaFfOB
w04aWH00f4IhYmf52NFbDhxFsvNrHDBACA47Y2o/+zqteYp2ENnSokM+FCxL9ty8
BCwZfPk4g6yiYsP1FR/WV/3YUzAZazMahsA9CNq7joRK7gmBlPd0BpX1EBoxflve
uqCI/j/jWGMcH5aMd/KEV6D4DZEkQAQGjpFaIzgzVZBm6TorfFaJ69WjvTET/pk6
px7pUq03pPs2JNnI1q0nbk18n7EifRFLzh07HGryjb7LWCptM/qaKQsbzwBZ7/Sr
36DQIB0LW/1cADSFs/dozk6C4jPEfQStClwRMJAp/36Jb2XjPSlVWHOz+JD248Cn
4lzDzw46cIyIU9WJHxcFUfYoB8sP5QMG08ghR7Rz9tI3BpeW2HqZi8wnS+ZA13Yo
Y14GoxoioHiCk+sOQYxOHxYfs18fuL2+CYYVZ0ZhBlFcyLCTNV35M+MWOvtLAyMK
qVKid6BEN6SONUAaAoMh9KDSxPty4c5ai8LIPwumPrU0NUJncckdTygjoZvS2EWw
8cw2ox8J8rN8mK8wf47Hh2bqIH3sGyV5OHFeJS4C8MModRSO3rCu5n6SJfMMFp2i
wQ9UnZ6UB9BpOfet3odUm8CF4z0HC+64VReY46O0350ibGMPV2e2AIb50BSyDici
z2K+NF0bWHFL9zkPQseXweiZXdL/yMCGqlckMyjeusR3PZ0EsqDNdVMbTF/zVE0y
EDFFKjgCIpLbGl/YedlVZytRNMJ5adjCmEL2Mm1VYkwCBUWr3EM42cgGAgP0k+F4
tFykAZpLpIgvv4Zkt0r7ILBNUk0BaW284hMLgkO8ebH0fT1Fc0zdKFRwTG+tASEA
m2NanokuakfneGC7jOhfA5doc3Rs6pmAvCzhQ2pcgRKoPt2pVFweSzi32rhLDsvM
lxn5c3Og86LK6OOB9J2A79nChjtallMmJe3LV7yA5B4QkOOl4z/i7QPkn4JwgmYY
+YjFL1x4/ewkqb2xrkfan/QtPOZxulowIpDqayiDTM7umWdKERnaXyXJBfWmlrsR
LlijGzhaFJLc621JUUwv0ylnZwoavHmn+ETCbLjxqbnILsdtW+mrmc1Snk3/g6PJ
4q/L9QVcYUsjlj45w2L5or4v2zEaFbyhFS2H39WmfVnem13lfHVu0rioBvrQtvNW
/WALidmKVk3kyCn5XykqBrEvIRNtZFG3rqv9dYavi1O41yEYsdCJRBO0ONzv3L6D
mceIlAui5pBY84OlIzH/vq7KokcO8d6dYr9jFVAbVKwoSt77jTXJUA6UGhLXddna
lqs8uxZosfynOjpZChBbkZhzboGGkJQS07CbiZAvkFNQnMLCsX+9Rl9bp2OV9vDa
Hzc8R2nq40GaXIP1NXMyMnJ79oy+0bXTYwYiu3ofBy/LabwQ5wX/nao0MuJNQIca
jQ8WmyUL7i2pvizisZrMkJjRCJPJXqOnSmZhn0HspU8ZgaF+d1MZXTwOXsSW1bOS
b9+LBOgvp5agYlLmJNA6zuIu+89M4xFRkafM2mtBQs8WYIBTvLBXkJJs0iJmPpZz
1cr14xqa60qGgza+/5liaGxeeMuLWhjuzEh0vhpZgsxqUW/R6ONpvFLGkxjtrsT0
QxP1SvCv2eBCHPv5lxgaJ6RQolZPPC+s5eE+dtTtp2AaA+AL7XvE9dnHCHwhSs7k
qgYH7gzAIz0sd8LJIyv5ZMG173ZdArVVPtlodaMBNmTS9jfSq7oNbjGlx6r5sVNk
GofoVkNvuKPndkShwNVIh9BsEQfuJJg3bMXs/ell94qAIKB91aCVbgz9xbukPJYN
Sr/Qg1fPOVYBVCiAzNNyltOSySzIligYOCaQ+x6W3pPxj8JFulcOxco/HPpwbfkh
V6iowX6Gd5/3oYVb0OIr9+O/vq6hvTQcpWQvfvJgQy69k/uSd43tuC90NgakAjxt
Ae4peJoqbzwLSL9VjOq8taM/434Ldk5vhAqnUyCqQQsw7mJyXz5lfAnv6ZMq0AJD
W7pZwuX/nOv18n/q9cayGLVOX4a9LQS68Rs5zZS+TMSihEibI++YCNU+kpzS1/tg
C3JARf4Wq3yOdOmLC+qwEm573lJPZxzq1uuCf1qdx1RJ/sTuWSK/Azh07h3BoSS5
GSUfNE9uR+4h1EmiFWsrN4OWiPuBhfCwno7XnIUa2hpDYgk9jj3cP2pXKvQB8sBy
/dyOt3smudnpq84twoBGWyFchBc0wn/oCVtEayfkODJgBcmg6xHbojkvZB3+PdT+
Pqdg/dOn2WndnfodOCKaSwiE4qimpKh60zDJredKjGfc3QKbw/BOuo967DLloHC6
Cotpe6V1bA0l56SyOmCbKEDHCwnrXk/YcI6vYLqykI/qCwRBMhdnBIdL11F5r9g6
0B0TIP6eP8cuNAOqEbotj3knkkZ/QufQwt/Q4NyBPnhJgLJd2xkBeX99IHk4Pzn+
PguPt1hmpECgqdV7NI5JfczCumuReaYVPcS0EodffvrDnAMH0Su2600SCFPk8K+W
NVjvCD1NAPdTjrlF1QGdMcfjE2KiVhpzmqzq6KCqk0cMeEawUOQlJ37P3jDE5lEu
rQiMD0/IVqUgNNHs6f7wl1IFRPzUQd5Bysoifm3qHUXAhamDZXzzQpH6U/5JKAlF
QYNOTRv60kiddOabmWH0euQKKli1IF7edFPL1EYbg6abH+0SdT3u8oRy8aRrsbf8
OAbyoNDVIMya7VzO2MjregyU59PHtz0Mu0sd9kBVfdCQZB7oF0wqz5wp8FoLbZ5J
xeRTf/eUtyR6aFjrvlrbrtLFkQH59qhmNPIQaN+gjICFZA4HhHt7Xgb7y1/ZauCc
N8biezah81AD4asZrufeBaKMuTOJJd23CJX2Wu5a9aDg73a5DPVUVYvlYwKowTbQ
4K0azpJLnPUI0Tuy3zkcsEMEPmzu1JSy0clgBKkqjK1qdA1dYVYM+4D4+IF4dEb5
Wh7Mmg8toIaVIENhbrtyfbcoEFvLrflVPfqBNVzw7cGbkBFGJiTPiNz0wrl4pjpX
dW7GwKWmVB/fc+fQyDHKYVZ1XmNnMURb/bAeKcxL3bmpuSzFKpPOUGVjqOdv4PCm
QWInK4jiT5V8IaK6e/Hp09dfQSQ3EMUNQ8H6alouGxf6EXsA7AJbpL1h4RbKTeVo
77cngyxCcemZTY/IUBshts2Qn2QSStlLI4wXLbD8fs4oHRjWPH3vTKug3QwwG2N9
fP4OSWrY3dYfjteSBLB8kaEPLj9zuKWXy6di6UeGn41pz+KtyPNehon+aEdZ4USH
Ht+Q/zbkf6Us7ud7DPpgQJ99PrdWFpGnWj/YnWplPQ69hFoYlPFi+3KOWVp9tB36
pz6sNAg1IZ/4/mtOVCDLHlgfLzfW21dDgh7rt661uDtxHTicnmtjJWK3cZNJ3IlK
uSmCXEfD6MwGoCUnG2+6Vmz+w/0KI+FHo4c1YmuEoi4iWcmX0IX0gjnhi/9fdELX
vuiH3juZCXYrsMKs0gBL7eW1aaLp836SkG+XbUQL2NWv5Qr+JZ71R1J2x1EzV7qf
7ciYTxQ9wx9rPNnPqYYFwCHw/CdKlXcssVurv/CNCJvST29hT4ujtdZEU7Q+p67/
xFRYgHXv7TArxH1ZuYW8uafHc0DltG5rIAPew0E+QPTHHeeml8TUTsQogpeCC3YZ
LPIWq7ZXr/DaIyOagrBONjfRKJEtxv1HJ7ByekWFsSarTxa0ck7i7Ppj85QqpxRD
eSij3Q+wnWeAwXIAsvdvRjuRzCD4iR4NJyFzm014yXo5OBKUBRcVAqIchflcATMq
aziqukZYZ1bc1eaQ4ilPf9OAswEb/JMsaiC1WKhn8bnqldV/GxbTbDJez7QhHhth
Lx0j1xUqwgmB+q2Q2qRAMhbYmBitx+rR+kR4iKNvhk1ErawcYcVr9gUfaVSOc+ir
piEw0Za+S6zfdmapR14THeulmamBCTv9A09b9YVBRAiN+xNYF6ZHu/tI8PywR23W
ZcZEMelteYDJEC+MMPD7N76/Kt0Ec689m6ahcWBqE4Cg200sfv6eGYfi1QGXo4mE
x7ea0/6OGxahdvsZuimDldiwHrwHbdTQoHQLnggC8omepLyjng6QI7d28FURh92+
bxTHeL8SuZ8Utpy9NN35iIeQuUOhd4bNbfwI0T8hdyGXv6NG8olIp6dJd7lVgr3F
yPvTmvz4Fk6v2RV9gfDhoC5JCosYnCBp+1kqWSpaP+ahwDr9Y/wuBHt0k9lDpUn2
vqu2lIAOaZU8bXJ0JsTXysKrRzbb+EdY3b1vVcU8XFrpcz0ggsYPAjlnqR9hXIdm
1oGgceIB5s0xLqMv+ydBkDdZFmytnitLIPioRY1qS0C15Pf4z6Kx8nfQ5WQwl7ZT
0l+S2qHqTw1t2degOGiC8X3JwuhcmxpUz1wPsKsMk8ISW3v1iaET/xsrxjAdU6us
g+bCJATBxKyU5BlADCpjpuebqmnnlYtyD09ul7EevBic5Z31RmSNNFm/ctrCpI1+
8fO4rfh5qFEEfFRgbjWSdbSg6unddVmMxyG91ySO1VlOUXuKurbQozWdMYIn2vmv
6BmqhuplWfRva4bahksCtTUNsinrdEdgLa66TEmRQ/XZ0thb80ElkTMkugOO1DJ5
1eZK6QQTBM+PmnKpVpmUSBLgIa9oBPD/YrLxVw06tnZyDEtfVrER2AH/azG+Bytm
3NU0AgB0PsZJNdebbkjnQCS1JPApe8//IyhUjFrePxaYNA7OjjhPC9fAHS/eivkT
RNox8CUtnj4b/bzk3saBn6BRkkwhcjtolH8uwai61Dr/jGDNDEm/X1WJ+4+eK6D8
Fv2U/P0xBM5UPpkMkSKaJ4XXU/buCT3v7bCWLqq9djh+M9hWovgR4/wCh1psiVXk
gWQ/dVs0Hy8woWa3RJcYvM30Li8YEpszJCcoRKLuor09kvzEL1kj1OJcLIwJl1JZ
Tj6hSMk90kKLFV5QVUPAkNXCql48JsfagDipD/kJc/R3xutkoerv1O0ZhTeKJ4H5
HPhqa0Wukt+rQzrJ4svUqLO2BvfQtY3ZoeR1c0m4irBcALrTVACfeAaH+tQbjyb+
VAQsONUWcWXhuULFdCDkYnQOjAFGoAGheTvJvmn/kHN7T/3Addl+aIYxkRvbpg/a
yLepeXsxxKyRCs8nFQc5La+4Bz/3R8LnSuwz4Exw2FadIO02tqC1YyZFQQU0U+zf
vXoZFLUTZ8Q/bCvOMu9FR6Wtgvj62M7jg9mzWCjlY23z/S/BZi+ywGjTyJcfvSjX
NdYXMKR2UvV6NUyX4dWMSAcJ7uNX3WBcAXMvr83Rl/f6tzH4lNuRdg6E/57Hvsfm
ZWSVamMkFwPI0R1Q9WkO14DE59/W6vI5rCXzLz5ewbFLIKyhgbOuBZPZm5ot5o/C
SSCnR1K7C+0GFzPj337LmBFrm83Zfw4idlWJPR47IPw4dHGmvISzhzOecLxagVRw
Dpc2Ptb7cEIL0bNIWFQhdtsz9SZk6NhARyIskoSZZfYGf2yOnpRxVHJaUL4c1icV
tbRq+Mp7bo1+SiPGRTUpYs1jWLsDTKeVjOgRfbcZBOcqN6kiHnROdqvPxcgHCegU
ir4zd3ub9S/6RbjJFBmybDiVGfhKQfJys64Ir2vleJuEc3t2b8y4jDoqx1ohRNz0
HHRKWvlHsycbbu47nDkBSFkx+txW/NmAfAPRU7abywiuNfgubH8d/d57J3yVvOry
JNWCK507Xdzmf78GvN8qI2EtoqcK+BzqX0tD8jUdpgJrxrxvQf3YU/9eENaAxhzz
d7Y6d43ECbUZDcT5qM4+MpBjCfxUYr/iKJ2EtO8sA8M+AoJiEw1ysGUOIQbd1q/3
707WrhOcHvLW9DhTMmBrdRViDlGHAodtCD5No7wW7QquJEFeQYitcivptyxMH8cM
UfLMuCjJqBgEa5iNQIetngHeoHdmBqbP0QAALChtdzrqpI1Ht5KHszWfFVQHMAsz
A4zlRw1Chl4XGkEuvy97ztzbtOKlj9aHdC/yfe+eg+vI1UQnOHq06IMn77HB/vJf
se6lmRdtH9mbnmufgmXs3OmxK0z2WhMEOd363nySPIokmk5yaq57t1GYC5JpiwjD
HdfUZUUQaUyOqvDP9WRnvp7soSXjjhXQe7SNM9/+glrkknT7gsKvGhprPJeO3ZXd
mwGGRcKC73pFXZkVonHRqT22sJ97932g88TNdrtrRcz5EMQwKgCkQ2DHDkK2//PY
F20YdeCRWXtbNbi4mmVsaq43vYUW+7aCs/giL8S/N2hUnm0Q1zJY7kzPej6075Li
8/ZuxgR2SFjfa6wOhKFALxIwMLOoOfyNMasf3ivGbaF9HAkW/HkHFA4qadQgxjEm
MOjw8erZSUgqfIoNu0YHHTPDEh62aKXeDJeuDzCnU1W2WmpGE83CFFgxKM9SLa9m
0jTA4BXixt+CkplXSXxHRLFHIvPLWQy+viQN5u4Ref8ky3MJlW8KKrwcf5wHP+Bw
kvwvDzHkovLUPF2NwLAYkGxIiQicldM0qly/Vgyr7UFpc/jG2a5BpYR9y+ZEd0vH
mQRTJ/qypuyCrQ99IXc4QqPvafwd0NW79YftYavr3AFcspEPg9GQe68bMAId+pWM
6YjLU+Jgcinx+KntVqRcyUyJk5zoC9ZArOTAiSVRwIGldKgcp0kRX+6TD07Sf7nj
JGwQKxatm4Wf77K8VyKksoL2NiyCf2K/8LbM1p4XepsupNAiEnhzx0F3WmpnMiXY
qpcaVzUOIRaitGuxYB+ckmKsk6K7jSETY2qb0Wn0RCeX92g1E8cATVBhY91kJBx6
9+Frjojp03Hk+77DAPRayVZ9OGHm+pE1A3j3Jp8wZ2nUHkbbtGqpWA8DIsAGCjES
86zlY/OyJpEE3tRpUEvA79urrWvTyW90Y3RZxpE1p3VXH7goj2BVjwqsJtEiAJFA
xMLIuJT6nft7T8/3Ty9deYA6Jrh1Pa9+xUIn8x5gI4JuuJzwbuzFHVkLtqOd6DW0
BL5RNTCaDmpXruOChpmQE729MoE631fcQbporw92gYD9Z1XQVysYbnHkPsBy2tWZ
faDjviXdDAC3bKju67hsE3Q6rdI6d5FwWDz8GWjsLylqjIorb5azx5KqOPHNzEZc
R1+00kUIzz1f7M8y02nzc4XpOC01j0GFFBKDSsDZp1+P+GLKA93v2Cb2jDl71/8Y
4Y6by514kgtLpqZU48ssD/l7kgtp5YKITFKIT3aAXKwK4pZigoVhoMZyZpOd2juC
CAH6WORjiGrqOTdXSPRZV1Dzq9uEmMiRaDDIsrR6oUkZiaYR4doqpe3ck03nWQFr
muTwt/SWzM6I6X4S4CDzwjlbO7sbmmQDAkJQjMunagmtRw7dKFTNdi5VIEjBdhnK
TMEqRTkeevqWvNF3+hT0je8WlF3bjLVAe7WtwDJJlcErc6YxXMq9poYMQvDCztdj
DmGTJ+C9NDMMWtZEFvxuYzI/OhAoc+vtBeIRqeuMeAJ4zHgPJougYUFs6YD1z/wy
P9iGamdBidYbzc19UAs4RHuuwEhhqhTdjVynubw8K2lekarIWkzaA82Q5y68Fq0M
DEyyv2digGAA+rMUuTkVua1dXUPskBX70k3Ab0HRbjpRUQt4uakR8pax8JAEuv0Y
8ny0u3r/gjGdEB4NfkcWgi98K/sFe84OLECt2DZEr1nko1YUh/q2+wPulqVdQ/Y6
GS7KTkfZoa1sFexObFEzWu1TE9LAdMgsGwYdf6/bpRn37+rZHVEGRj2hP1awbalL
LXA8ynL/bEji2m8c4Xx9EpsbZLICr4436J7MCJPtzF5okrgZedg2YEDoxlwPKxjd
PdMAoifjb4Fq6MiDjCaSuAynSR8HRulPUdZQmcWM3qnCrslkv+yC+gMHpAHlr6gy
IJ1XAN93+/Fp6aPJAj2eH7sxUNz9lasdD/5ozdDgn30KjE8GPcQBXm6/NSk4Ny8a
PsVxkrfg9jBhZ77fFKuOSou6o2vPaC5oJK0H6v9+nnRu4foCfDbs0KIy457Tp/lr
j4qg2U1O1HQHTnuN+mGnkqw55DVbgs5SSNqv7p2jANF/lDSluQbBwzQ6bj28MQ6S
9nawU9dAV82vdWjApXeqc3eLOSjAjHf4IPo60Pw0qmDo81+tO7VxSaElnHxFdB3e
FcAr1gCVWCpdgI9gpPSfyi8zFAElwO5SEAkEbIp39wa6jGQDXJkQLYeTaYAlUzIX
Vc+Oh6Ug/kZlgjGzaQBqkkS/ugWR7WfuqAbyRONDMJf40YGzI+W/JQ09Vb6hq/Z8
Zru1YUTAlvlVixCnD4azWJp3k/Z9h6/OiUzHXo3O1DfsxwQOcZnOpbIiIxaQ+Ju7
71fr2C5Lj9gZcU/hohq6uOabJi6va/hLxxkTtwCIrlrvXr3xFkwSSBBJ+3B4+CZX
fFGb8X3ofAGusjvwz6+amvMjeu7PWiQAe1rFjG5lTvxfOXQT+UISJaRwzh6Rtlni
9IlffS0tFrvquPg1fScFjlRYub5IVCd3GAsq9LUhmSV0ffEx64DUFSWu+IHIKEns
7/H0Np190oFxW/Q82hoxA5dwg3xN5ZYUJkqVUrJjLdZjStY4ayXn1pAAH80P0yqZ
z8XR2W6/7ajaTYN7eFqZ905laiG8Zp9Dd66B2lym7g3iCS2Gl6TliCb7Vp/Ln4IJ
NayQn9BxHa7Ot1zwkttGb6UR0tnbQh3vvlvVM73sKlj14PWZCgEL2ZYmyGSHxnXs
enVNT/sT5wCi/PO4N1Ra/iXSp2vtWyNE8ehW3SF8pep7o0/2uYPpwHj9Q4qdO0S3
s0jG+VASJrDp4wdHd7RwNDDHWz2D6TIuF8GdN9GjYqbUFeqfHmeeBCjHUfNFbGR6
Fiz7yKXgENW78NjSVtlB+FOFJ8sPr1K3AOpTexrGEkWhlXrFdyKwKpb/EGfzUhod
H8+L9WiQyqBntTtnSMge9HglVx2uA6JqsuAnasAiYMFuys/AXxrSqjYLgzFsPdwA
ZamNfPexwlODiP/jpbdD2gizUfmtDeMWiliSwFzQ5XoVO1ASb8CSngwmgm604AlL
hNQYaS1KMFxlkT3Vk35JVquQYgPdeUSVqjpDq5FE0oVNbf0CkXFFIV06XtGbgT3V
obJ0xGLGP4KmrgFKv87LLRwQ23EjoYCTYbTVhzpTRk1aleFDoipAchflMFd72jkT
9K89+TnyVnHRvW4kHIzaQL405kjmVUnjMRXeq93bmg56L3FcCVuvxk2ULp6F0EK1
zRiNFQfWmlhpbTWo1h1vtPJVgAWaYTgFPo8Sp8Qv+9X1aOH7t/k/Id1Ly/ZOFvsf
JtK9z2E3P2UAH+xtya/DWTUzPDFjtRTF3VKlpduQgjr3EAINoep6VfNatQg1x3Za
sffjJlLJ3pjCyyKjeb1Xb+0du12IedGkh/f2qI0WY3wAn6C8lyENQqSizORbJIk7
KGFRBPCRKFoXIicUpswQhuMlIgJvJt2ZS4wtY9IUUPqUOnOPQlhqJxdnRVzog/zr
ikQ58VSwkOp3ef2YHDpFF5hvQIih+Le/5MPr82ozrdje2HqoqACLTiszAHP9UpLf
s9NCcFGXOr+Mc1KSWTG1a0fk5UZ8gNVbKdnU4y5C/LlZuLunttEAQyr4u9NIn2p/
eWHJuPBSE7Dvvs2/p+cPrbZ3z/jn+LpYvwfnG8Ljbxl/LR+9orr1n3GQZNf/z7h2
R7LuYctEKgys736eOw/GP9zGEi5A+j4jIBnL6MIxhx2MRD8Fh/dDlJTjvz+dFLM0
FqwXSezzwkevyizP/IeRVex7OPS5/TKyO7W/WqDJZanaWIn1J6VjyFW33sfISP2D
APGRZB3hz2F/qXfv5vp+h54DVSgL20GYegQ1avVzxUt+b4aXliLGP139nFhD0BoO
RWbWkxESIxM+VGeafeKIrQ+bHNNC8DcRDP8z7goqPjFC+6Ot17ju3GPRFyiFP+ud
UmskKNn3hek7XDhy5+nnX9zi9+6o0q5LcNNeTYFw6h2NnwZgr45AX1en9CptGQXe
OfwtM7tolIZWm7LH/TZ7LCn1IelGk0GaHOPGaKhFjzEwkAktle8qWI+fC7xgJO+B
gR9aLXRuvZqD6053nHZog8rnr8WGd4mvtl10uyinikgdLDBiQelMYJjhnWB7lDr6
91G7qiediLf/ED8SSAcrDOfe8XZvXlmtyffi/LC+MMcW0nX8bCqMuarWMBjOdMnA
BZiibPLHVUdTmFx9+tuenyjUoxcw+KZVSA8SPrmeh/lsyvzN9PghnvZXJAbvbKmY
sB3MkLXJ94KpVHfESNCEyyogY6tyxVdsWKBqp+XmAq5QtChorKTh6JDE8R836qpO
vQ/sSbREcFhYWDdOL9IFKN2zK2qnYdXD/rqgzFeWgy9kWkOdbb17N6hlgvBIn+Il
Ns3la4jZnpahSKNS9T+6DeqbHXloTc5fwtGWw+Qz8uo1gK33mJS3Ip2K17B3qmFF
SkvwPGnaaz4j2qzbJIa54+48YU3hLZu76NLIFtjkcfPZP8thY+Z2O8lSgy8l546R
vmNJySm+mfR9qoZkldvucte1CWNKSMsP8TE5wMSZ4ODnAvNLkKIJ3fXg+0J9SFVu
wF6MHnxnEka1ZfrBum88TsQEi26qw4rDzol59Osgl4h6VlA2AeTIXoN9E6IruoGJ
g+6y4OLqazdrTLZ+yiCMm0vFmrc8WGlGF3ql/qyaywZf2zdoO355lmlBnPGJ3Tm1
H/Paq62qdnROWP0IGYwbZPkJEQ2J1rzNmjL1kVEuEWp99jajoGG1GeZxKWo3TFpN
sGQapQiui6vi9VCbxRC/erltDVAXib+aGNQQGvhz/crCtnX38Uny4k7SCU5qc73o
eDjlCeDBBjoUalha4Mgf8Dbxt6PaRQNcKyDN5twhaHYnViTbscZBERgLEw62CTmt
5AATrMA6tDLAQbW0JxOjfSVECNfwVub7+sbimuPanDXuN3FPKqMGC4SUcZYIbMjm
in5uq6nXfwJQCUvm1JiK6ZMuOnjQ1u2qyPpkeOKxB/qB09ApIC0JrDCNNBEtKn3i
8SK7CUXnPLbaMfw4Q4+kyGqlX+aH210xRIjFsGdNDVFYXO00Wi3XHR/XpPuaAqV0
085Mx650aMd9L49bQzylEfmTaKIKUQTQ+m2Rv2CgccO+xWMrd5R3vX3OcVseuHky
tZ9nZt4w5dN6bVPHQx+BvsPMirCdMxHzpjB7AZ7xaj6o9yVxvIzlJb2F16g7FfGs
JKfpqs/EtH6oWfqvJa6qM8WBFoCP34ID6go1oiB4aA8AEuUPM+o+CEpUgou4I7Vh
CWb/ScxE7ss2ZqCTLiNDDnKEi+v1kFe/8dQEUbLYqdZRiwcmzc07IWiCvbJSTzhA
jCW7Ns9Vtd8LiV7jeIXxR2Rz8GOBDAQZRCbVSCKq6TXgzPcjyYa3bZnYHVwFNu80
BwWQfClDjPn4XdCU2ux0LpwreiByXmBTcd7wahHpsLp3Z//09lxRxBrIkPz9rcgT
TZAiEhGfkBHx9rVaSHjHbAFd222YeAJNXsgttcVH6MBuGOSCNB8NGLFUY5NjezFb
HaYPYrcaISHM8IQDVNrrIF2x7rMUKlDPhS4vOQK+9dAk3rzdtGY+ZAcdea0WIHVe
/lwP6DiJtiXL6HJPkBBF0DH3SO1Se7Xj9vxgOcld9czC1msQpvonp9G9Qrs58aus
8Ujb6Hz96oE+L9yGtLr9OnEdM66FWHF6OzIKGPf+xnIyUGvS5qEZaGFh9paLCrrW
PDnUq7WgVyyZvfdrDYi0x8yqtAAF48f3XTYhp5UGEWgd29SLpwgPRhzqs4WeY4Co
2xEVPAWYbQdZRC6RxHcv3hUhcmzYb7gAwvUXP9+4ivE3E4FTyzq0+HW35p/HA3Ve
1RlgGtkIhoeE9/WEgIvkJHZNzgqR1FfC/RAstOA71g0NwE7pruWk4sd24JXiL9wJ
v+FHRXP0hBOEiymV/Pto1f5K7nWpHzCx6lFclVKWV3F+qrYKSfS0uIVSgLMvs/rS
EGX90KEWx/7zTDM9gGuhphCRJ4LKta9jWZIGfgXG3CeQoT9hG+JZATzc87XeqV8J
jFYYNZgOvuvV9MYzHywdt8z8hxUGsaFARAl6wmMX9eyLSY5xW7BgMmVTSh4XJaNa
cWcLqQ71nR9lvN4OKpFvRIcGtXGonWczsn/QU2w7TXuPKxdwYLAqqzIFChk7lolG
pltF/8r9uWCggUIf2Fr2p+t9KwYzv3DWw4EDquRwDDO/J8BnzP0Ej7VW5RXk5hqb
LL2ZBr6qRKVBgJ7ynlLR/HgdWfHKPEHpn5FQylXQx6I5cuIMA+x94OzX3kDYRwDF
06VBkZUTVT3UkG6SkcHObMJfY87voJLJ2Gxw/GVfnj8UG5YZej6DcFlBcFMChnCt
xHBgm3QlrIiAISem6t53CeYz9vmSt8upHgxAPsW+r6xu1XCoJg+dtkj8jxpLIPY7
bdlOYmiU71MfEhGN/cI9V0oGSoQzYmwoBmYXnHoUi8Jmx0wwK4D1tlm4Qv/bSlmj
GEzgcDj79Ekfvme9dipaN0FyyIgL5EQeVUH7jLoAAVnWylVvsZBdMuuTwToo429C
yn6THOAd/KWi/41xjXmqh2o/6V7xm+wxYLo+6/5iLpqJuOdQnC7Muki/jAGrnfcZ
5FFQ24YoG76oy86dsJNDqMPq2G9NS3gOmMuVlFpilZcnDTOV/ANRvlzrGnm59CoP
TFokoGdxJxNKPbSDbgF8UEw5nKL5qOXY2r2bsgNtqZbqhK/rC/sXxyf7sbWjnWHy
ANNs9/mYTtSfEWf7A/+Ju+PFiKozQlpl1DxpzY13JujT/URITDvwe/vE9LXkTNJL
A98U4vzBWWs2vGL4lY/uI4Mq0+i3pBLD+N7sw7sCd4yAbpQzl5aRXuuPaIY+Csli
j/V2djY9uLeBcJ28zyUX0u9XG22IEf3B3aGgvijHj+TISRrFlgxmAoIfPBQtZvgZ
EOnTBmrM7lnpDoT7XH8urNeWz8+UGtFXDYfCRYqIe9ikxFRjyfXTfIdopclscw6R
LGuKC07SEC/TsZtbdimiU1q53y5sU/ICvyFfCGsCXhWriH3aUUvgDgSV4P6Dpqr0
2ABQ0XDgZwc5SQskcxhetpF2Vo61xFkX5OQp/u2OtH7HbXX9LQqlDdLn/bf2dUJd
Jjn/KvALUhH+ZiEVazsT8GtgFZelares3J6/JS5YI9qPCylMFgynBsVa7AKFWKZv
jFiG/+7IhXa6ft98rDPxNuFD/gNOhJZR4wzeQHbualbqbL8HACATvsups5m46xCY
X3XmBzwDPhjxfL6EMJyzlz11BtXyE5FH8TtBoPOe/ORUh51LkSuAm9tFndKuoEqg
/QNWUUvjqbQPJ5oyTXk27eqK73RqpZ/zowStfSxVa37tbR+UHpNpSd8MIJJ4Z/Iq
KDNXQhJt1lXYuFwFyQhTd6PQfIqvKqwfpWgij7J8s+IvW93X6ChflNz/Em/GeWav
OLlXAvSNa7SWg8mEW9T3TgdM3PbI65UmRm3CYSUBMSbPQT4TbHGpqCcKykj96haw
PFUFxV+MTVY3lkGH1VpMOYOpdNenEW2PJY20/NFlB/g1H6ypvTAp8KYaJ7e76SwQ
WVkoadA2SClcoJnA5XTnEd3XVFcJc7nWC+sYGnmhcNr4c6SNK73tqIqHIFAImh3W
JDs+u9Tfkgt0hJ6rQGdvJNC4ZC59iB56QSdatYfArjAZpoGaD5qsrLSd6x3q/bQi
4FY5UnCTJ7yViaGlSg2+aOm9Gh2K0+Zz/QZROB3ySHXxIMWS+REndrPQ0fhHsPQ0
OHWs06/hWA/yuqhP+aqH4yNvVTv5XsYhWgIf2XePGOOZWwSSIoXIspw/lDObL9g8
UJt+bi6KQRojrG13qmc7cCJLE8si5nafoCYNMepLLPqFx0mb+7EkzwY/CYR+Vz4q
Xf+dGRTvyr0eznVc5BZAYH18GobaMbZS+hZSI9Y1FtEwfuq85k2oHLmEAg1mJN0h
HCunngB9vr5xb7Cxp4nWMWIN8kR5SuD9VwDgtBhG6cJ6i7xUEcmzH4Ol3S4Ft/Zk
1lPS4nzatr1MG2ai4ZNgurZZi56Fj7IMPmqQVzrA7xsJjM5THNGhVhmhJIUop4n9
O/m5qlqQs2D0D0x++FSOrOSxVZ7SlAh+qmwOm78gZt7iM4xqjXMfhS9GrpeLOx5e
CZIh9gf/vtNOWpwVlNuZ3d9qsMo1UKSTh9Nyvfu4hUtfABW4rQhPMuWYGeUZmADu
3c8g5vKPrJCQ0dj18V103L5QuLjqGCPC7siawN5vAmPrir1g1BdeKTTN9m+SfSFH
UF/Je0NYuHX9lDbo0m2bNmhvEGSuBa+61QtXK7HlM6HC9Y+VHCtl2hlCgd6l6QHQ
C9gMdQ+WYMhxNCDFlgXMjCMOqnT5t153SgAaWle4B8w0oRRm5n1GboHmsmNq2z+n
opaXi2Qxx7G5iotqg3MdrTmQUzMq7l9NDmu329dLAqQ8/zrqcmNV6GSFPjaFJr2b
PMeUBE/5zKAwHlzVdoKCwssvqEH9ovXO/7MYgME8vT5Nxq636q03fc1AHH1c6SAi
voaGw2sG99Hrv755q7C3xUnJq3x8qropF1AutaaWrQN1ubqi29d0lxZVXNcs6PaC
FDfPvEi4rFWBa9OzDpBQfQsy8OfjEvGKQH/wM4fnC2SBZPhQ5Wqvoia7G0zAf0RS
pLmREaxvMDmsqQ1zs50XSrkt/oBxDMRhW5WbiEUeMyF3VooKxkBuv/LV0rJdArG3
5xW2Yc8gakNmAtUWpaUdUD0IpxoZIPOeBE2T1deK0dNm5GsRasjnWkI0IStW3Ysj
AS+SNupZK4SwUnxcYIvM4FPOyA2jvFj7UMshb13q5SpmsjCe03xpzagpUtYxeiip
N/6IWyXqbPnanLuVhhtAbUTUS1bZIAnhJ1Z6uLAYA9NXTkPfzKjnxS/uYIrBjerq
jn3d8YwWO3MOTqt5qx2kbby2HmnhLLYxon/I4ZGrS5rGPaaqUO3fslJnu9XU1tyK
ea97lgN2r0ffYNoh5AZkBYGxgy7keY7+UOvLR+UUU4hmKdwK6GYLKV+s5VNH+7kr
rLOqpCETRbFACkDbBXX8Z/sxSHpSLCgqPONgLVLWcQdvYio+RZzNWqCn59BS7uJL
9X5InoOsz6eWNqs9CHO/EfBs8/EGhlHKSx6KiwWrBeS2cN3IqjlE3qLBXNRQ/TBS
MoN3BkgZvQl6N01Es1AEwIsL0OYf68nwYx2dpgQN6mnoYgPQ3rylYwRJDv/X6Tze
t6hdefOd1ia/uFg/BOGsSXLp8j3vGS7SiEvnFH87/QKNBTENevfWn9HriBgAyEvz
5ID51+V/aCiejQAvDyDhIcVXfnBPcz0em7w/fx7DVN5ARUg2d6MLKnDuyXxCrX0l
PgL/v2F/oVmUZyWLgHHJzX20pUC7J5iXH72Frl5yIXtnGsFr2z3X/1PNASy3jC2Y
SvHE3ZW8wmpSRzIKv5nyG+Nga0EWtbDhKDa/Qu412mg3KlKGquvFgk5hht0GMwhO
xfphW6fZ/Qg14ggopXb9qlqq1wmy5JRoXC5ERmO6YMQanELQSJh2ftOZQTas59Em
1hylhv2Cn5f2ngOiKxJLQCkMkubk4bCGVy8BQ+hLIRvfYNY6T+SYXSq9ZLgsJ1do
fkoB2UIH+TTYAXbTeNEVN/r/PKA6sj1Khi43N0xxeYQqlQfWASt8fey+UV+19HQk
bKQAC3H9bhDQuG6C+P4b63QXW4aepjavYoI2c6BIhmXxDNRnkio8uMjctfxsOFnO
M8rhdYvEFxWt1V70giCDcQhuvOS8FdJJ5sj3Pd9UB/FSqaXkZEJMDF1CzvI38viY
05hs0hUo9RYJPoYWHJIdwltuqQcj25a3UPYlb1hFOV3S1p0LtvaFD14mm2HavoVX
GuUYZcxwArX5k3J7v9g3/+dE7ZLt4FZy66JpnDKqtD6XuS3Pc+yE2llc24tpNmF7
OY7MDssPfdWwpM5eqa1QLdSCzlWQKZypRvoCKdYlttUH639aQd0pQgWhahFW5204
qUJTKqnBplK3fmX5VRLL2nWDUDed9nlQes4ER05etJTd1riublBjcZ7bvfCy5XLJ
titoFQOdWm1soS8UHXERqZnSXg1062Mw+9tFtrkYgiJJoE2bDirZvNZXwH65h5kJ
x1ILPcrnI9fy6o4RE+XmtUEEhu63eOUUTG/m/wVhb6iWqkn8+uqPa/mnQ6N29vEG
yMF5k+9kau5fT1voqAYn6NAQ+G+PMPNZCCM47bgLxGZdyDMSG3vJITlpGl5Xj7E/
DCQycpQSrkysskgsYS+qopfxI/970R4AvrxsbJ94782k3oa/x5AbqxrrW2dB5YD+
hVlo+kdjj/7QwChKIfZpyoi9sJzSfs6gxYqzSTqgzzrBW5DcIwMEeYvx8SNOVgvv
YUylOGeNK+YR/rVcP/Krytjpeo07a2Kz8RXqIyx2uhJEBnUScqeNQtF75/wYWzNd
0YF+yEmGhiQP/ms430rBTLR0nquxqW1QH4TMwUSYsHM/Eez9dPd7avyAWpdkj5IN
dKrZx28qVGWrsdu5KsjUlr1e7fZXxHlI7WBUqwMoWGqmxKSUr7124d5GKpfhyyb+
lr4Uy004iI4oPrpv8y3E8gf0vBSywMx6oHWNuSNUFIdXS/xnRRuhK8MiK4giQwFr
Tk9rEAmsoeTPbAVCXtMOyrd1BvuU2eyiGhSCK3cX+aZg4hQ7AdHVW8pEqcpyxKuZ
mDrDNNN+RZLaK2hhc8CE9wlTRw9DvN+2d5tBSPGDOC37wLtdMUCDr58iY2bnuMPA
9FrpM+UeOa0IUGagBZiZr/J9h+pjTGrSQbEjuAhBGNiJ8X7Xa6eBK6AJUV/WFb2y
gZZCFs3injXy/nKkcQt965HIw9sRtay/ZcbvE0k4ysdWnD3PouAcKQattoh7CBh1
Edq7VpYb8u8/dqKR7ajOM0VYIdLkPSJo4U6YhSDjU6CfInLyn9XhjNbIPVwhN7AH
VJGFR2IUWnUBEXRmiJUWq+dnixklWlf7xhN7uIJPjZtrYCc4NXHyEXKk66G/GHKC
LZ1ILTYexGKavgIGY5TRcrdDUcM946MbovISBr5gH4Pp2lGwVRNeYZVdl/UZEtNM
1AuXiCUYQgAcSkBJRgEUS+gcTOUD8S8akAl1VBDnb6Z6aJc1lOL9ucIxMoawNdEO
dJjbOeKasunqieRWURLc3PO8CBO3QaS1soz53rJysOsBvdbDGKPrD5iLFqm6CX4r
JMEZ+fG6qOi9mBRfEOYeUCrqQeVGYIU2yc/b3+rnrvqH2Skf70e+hCZq1sm8fxrO
IOAnraKWckyWXNq4XocFuBxLEaKISaa58ADGX0aNAVN0Z+GrLKK+7JOSGnPSjYb9
oW3pYzKugy31KhMgzLZmt7sYwrcYpudf10qc7ZtLXjDsU4+KY8klsrKCI2UG4CHd
jxqb8diYh/6fJ1nmUOVgt57wgrksVP9so2u37Ho+HZhcs2G/nKuhvvBuB4zTmLx3
vR0QQSrX/0ryXkGjgZeuhUG294zbfRfxKPnzQa3KX8vTdGQb5Q+oUGPrSS/dt7Sr
c3mtnCXnYRFUz3Jh3ihbOCCRdiSlb9LYilSSOMaR2+jLD7Gog+QUY08m8pfKGU7J
HFQIkNzoxoTzIFZYYWpG2OI3FAu3loRgV5VArMCK1f9fZ+Av9q7wLsTB7uYBckMG
tu9BilAkrsXcqKxE3eDHLhU5UPgeYN8Sg3xPiNafC+9PacF5QwUQd4a9Gqa9KYAz
rh+Du0DfLijhe0oTUy3+ovj5KryzTtbRbyx5OZVv6ZXUgL+FbXQ2Pun6of/XYmB/
G5MlcvLq49JczfWkLil23RUIXJDUXKR9t+sEfa049V6q1bsiHz4jPl0JMkhIgGF6
Z+ncLvqmwZ4ZqcdHPVxl/DJ0Pn8sZmnsq819q5G7QxlkQk0qfPTetwbu2FWeUq2a
ucLGt9GgmGGQahI22g1UWcOIs7rWXzZSE+Txn+Yn6c4mFp2LoKZxxqeHi96Q8Ga7
0nxcCV5GGCTQYfKCFpUsCW6gEGzIqS/qtQ/KxS7SQEb3fov62k3tYcJp6+gX1mbe
52BfnOX7N6qLdCpEC50dqb9pzQF19//nq8pRKrcOxGxg1NouOY6/7DRhzDzBIdQk
nR/YPVuI7+qDyZii1mWuTLE7HV9cY55jnGsS8EB19PMlkrAPeVdHXV5CMr7dAAs6
8Hn5aQZlSGRat2LWzeNQFWbZ6SOH+g3/w5H01JbjkJK1SAoAvApj1XcxX0Ficktz
yu21mp54YHFyn2lXFtSwnqymLJCEA8B/C0pnz54mgNgPnSC7yamj9zuwbs/ADxVm
x7/DMcvDU/ES3koMzFkAagMC37K6XMxQtjC3xIN2hYfHsQl65RsEYRmO0CAf0Cfj
q38T/ismwaD11Faf22A98k/t3315ZmMVWBKD0mSsfjW1Lub5Oeq5KsYBtGSuT23e
tTXPrFd+JnVtSUQPzc4VFHvsd32+zP9iNBps5CGBevZQrjgMugj1Ao7/QjDeVC2C
LDoHzCaD53NRfs7xM9qMBoFHJfx20LTS3S0XPjUPSS0H9Io7RXW/hMj7qC5Af8PL
hKRQuw1SDiGi4PW71UNWC35lFvZWDNklgRHMFlob4V60A1ER6c8ZY+b5FVjT5qdP
he6MOxCbOjhJC+2V2UdedUG4VpgvEF+hmUYJanthxRWDdRiGqUIBhDRJDK3NQs1r
vV4l+bacOTJWp9actCP+zo3Og1fcPDcCct1/J9vCZDNVLzU16qh+5tChDiIgdAxg
U3HHFyFwpZhVthhYHZmUl+pnZpg+4Z+LC/3DyChGuMAvZd2QgHotWzzjgC5t5aaz
shPEXXA5PsSSxmjRYiS3XBQEQgI74cfLWp7WqWYU+gzweHP6gGA28yMnzSnQCiCu
3O1j5xk+ISZ1c2hWistGz+Ye6G+2wOqh5SBUcconY9ZU8HZ5jc2up4WBlQGHTkbd
LhsXozW+kuVqUib+kYMz5+Ug0RBzmrRWj6XJkk/+LLwAjH6O7v7bxi8RT6RbEhYI
VPHbLmfAT4K1WlBlrttU+/+cxxWJ/8+vNrR4rcsPt+sCov+kM6nkvY9YBUW2a21h
T3caLZv/lI1/euv2qG7uNXUtxhKahhUXNpeZqwBRpyQU8M7r3dseW32SmLsZ22Ok
kWf+I0OJh8HTw4CZ4dOKnBN5h0VCcYKKIm7LWYjyn8Ly6eMgjoRkah8oKeZTx0fo
ifhuH9v6h8RCw/j5vJAZIMQSKNkEHzENCXNefPvz9bpwwRFQCqe2tlgDW9A4SL87
+gey2hGlJRFN49O4WcztzlWXZa0xoY1kI4cSgMy/VFDxRCX5lNySnt+3Ogpp5htn
VtCT5o23nDaIA97cg7hefoAtovcsS0uoZ3NwI/ilLkIBsZLBZNk0HrZ162aNV+fW
OdLeeZLJZOwsGhfar6/I6/+M6fdWMGSYpzYhVMez3bPRwsRIQ5DrVURB42kMZffX
sYt15HGegk37yeW1cwNnmQLpAd1YoJ6As++UGtP9jtmIDadpOVNAehh8b8QPMnfg
jRAmPF4tSV7w98q2a1JNdceAb5rQNNiOPopJeWoUtBgflTM23GWvvrIZgksRY+ok
6X6mVyybzvd/YH//Vov47gs9eNwwnLaBAVS/gcVn+C+B4koXuNfhmmH+eqQwEekz
1h7nHZCpAm4tvrgboBmPhwZE2h6gCLlSaLUXTJrfJ+MhHOGuzlVsjao4e/n8Kd0f
iZGcQijy5So79lTQ8ZoQi5e9nwNTgYMOb91hitOhIlsXvwFHBaDfrEs24BotnEdG
GisRq3GooOAJR3G0TcfQeAUVGwb2BeXeTlXzuX4Oc9KaJu8XDbf5e4iqX3cKpPnJ
BJ/WjQdoOvm87JW65KmvmsjL6fIAJzDAdT17GsPfbhBSLG+eLbW6Ey/4Wf5/ZFDT
jKoCz7pZnN9oLwBTE9n9XiQ/R/Iepk3IKC90CHktI/lJ/IL0lQzWhpSd8ukrB5Er
I0/QaEWAZft1i0UL1BO6D5EIUu/0nwLDiDIoXKTM2j9k2ICKKCrYkSq9C0+JHc2v
VeDcSMuPBBb5RTbw1fpJWfII16n3LRofsmdXDA4fkOmupQpql8PPFnhep0wWVK/1
FFTRIjvmvnpA+FCF3axWnsRFKVk0iSFxfxz2VE21XEoRPcJdv5/m4bXgGG4mBSvv
+hWuOvNFgfT66alTA17MdLu2d2Kvi2/QS8J6D5ohih8uTsBBkt6XSY7UKdLO/Fxt
If9qqzB5puoQHE+t/e7NSZjxfngmQZ50R19DC431yCkxnZPlVGUQtFmEBtBHh4c4
nqoXEvEU1UAhxwP0iw/yXWRPU3X86TlL4CbwZ1e9lU5RhJgmCTsITLVvR0GzmEEk
dxb9vlupsXlYTjIyo1EVVWbp2DNON7moJUph92GeICk1m2SM18ucPR7HVAwyj8i9
mBzqjRHUNWbOnDOEkieBzXdvvhrjncUMcTHQM1wvZYOdg4G2svB4BU5eUmWRANS0
nMtMZ+WrHw3lztRcUncfVN6Yt59c7RgB3VAfO68pVNyeMj+gPHgj9RJbOe1iOHhK
0H/0SBMzYVS5z2JxEZvjLkIg7kDqCPlNBPUdxW0+RSSuG1ol2eUeM3z7Pbtu3puL
cMMapdOkedsjglubmlyqHY4ydWtfe+z/wGpCyBpMShUv6hJq3TtQWY0v5ZCZBwCK
pITpRSUXMD3pZ2k4dKcZKFH0mgUYLJQdGlmFyPdt/N8LIjZh7Ew4/GnjLOcIkRt8
oVumR3475ESwPxAnEtqm2uU37tSkPqI3AQz+cMFeKyiWRXargkwTJN1VN9PqEhK9
57n7+8a/n6geQABN7fnfXa+L6rpsX3Lih9bhdOdGB7s5cAT8Ga9JP3ABufhx4XbW
FUMceWyXOq5cJgc6GwPpPNblP90KBo6Xe9cloUe+j8MJ/UI2pUhVWikkVgpZO0rj
2Gy7Us3wCnw5JnSQsFUWlG3zZ0wWVpIGsNx0TAxxJCHGrTxiw5Z8AoLsEmNIpm4g
/3Za1gWlBtQFxl5tweQgk66g7rDG/bDrT3Bw1DK8Ean/J7rvZgFDjIEMow/86QIw
h+hoHaHz0X3FBqFrSfxvo///DDNQOH5SeHlN8Y2hCf7ltok+yslw3LXYl/QFGcV2
CB3R1h9NtWbA0hHC2YT5qiTHDG1Kz1v620cawMu/a4a516XPOXxJu9k4ZrhLrDu7
xOEoU35Sc2RzgKsgmTEimI1LeZepTUsxZ5fLceypzDwpunGYOava0njvqemvIUwT
fNZdLEqrQqhta3YZqGBRv8nYbFyOCJbCw38FrkSPwjuyHJTsjCovtxbSF8dnbSfo
/YD8hA4PILgCgZchPZjFz09Y0TtkuJk3Yo7BHGQliyPKG4sNds7pxeQbtICr8mww
x0eM5u+k5/BzcCqtZEMbxtOv75ip3a++LcT+giCcMw4LF8z2KfPqpGZ7jp6XtPnh
YYIZNLEqbV23gkMK/fI5JxXiD6nzE7BBiKxpnIEJwGjiTPg6F1np/kyAGNQowwVP
lqyUcQfpJBJs37MtbM4RLOOWOc1h//8M1iGv6QWf27v9iFdwCfMHq9Z/V8oX6Khk
P/K3KxyEYPpDU5+wP+AIY27RGDqNmmNuv+yvnIyOLl9dPifo8VDOkcMd9oTTudDX
t2eStHYEkR1mjKsJQW+OqOkOTyboIFwQEIlmVEmmDVz9UAAQYwePr6OhGRch9wFB
g88ek0PUczJDDnqLw4VguuXtOTjWv2MZPgB2HlBhu7z4pqRnvYlBIEy3uZX5DAXf
jfuNhTnedgi0T11eU9NDkfJP/OAbDs9r8rQl/AAS+jX69cIiUvsyDKqIifC1H6Uk
ITJ0pGQsc9ERAvDJhGHdp7ZaxkMnEV6XqwUq6dG4aDwKmanQX7T3ouNY/8WkYJHQ
k7hAqTgDCizm6r8nZCFCeStfBJWqH3K3YKPun6hLEUNMryyXb+5tmcm3p9HXnFhV
aaYcbpCEWrgWCCBzSOBWZvpxdvdeEjuEynuZlB0p1lYb8VHgEOZD/8xe5ISs4iij
b2AV+IaZr81Nfx4f8sR8tqoiZbLnwHCFRVAs5vsTzPQczYcF79PgToUjKvTlurxp
RZaypUvTneqA69yuM8Bl+lNVfA+H8RDe1N3nC4AN9BCh5adhg7Rm1fS738O1t2Ya
QR2M24bt+hCljbBDF3NTJv2g/9RaIG0AUPcUTRE5zVu0q6bIxRW7XDWjjaubFo6B
c5NrhY9EaP1xjWHhlBAivK56bzRVhUktZlKhiqJzdehxx1zVDdCtnT7gb631qP6f
TeSuflvwxMlsxVruwsaX6H+RCPD7hiJyFBS9v2yYIardCZ7hmGa/e0XFOI+gG9IX
m6nl38h6seKwAfBdVOOHBOiS7ALTbB5Wr2YIA9h1bBFJp4m1IgOfJYquRLB++RTM
2XK5mwK/KArwC0OLQRnf2o0mVIE0KIDVOZKUJCQyNyQXtvQS9v7EQVVWwCWSrtu2
1f2OLo6v6zGQ1gHBv7khuSyU4a2Kj365VCBRxg7wOLjDBmfYlFxRvDwrG6DKA+Pb
+TSbsQevs3pP/JvuSUvk7E6RdV5SSROMgIy8nwCsid3Sp+MnUexjqfY3ddQMcN5S
iRbtfzXmqL6kAXcuScNZ7QBaJSGEAiUmCak7SpKFTx344LGb1w8QxT3rJ3IKzcvG
6G48n5U6QoQUKdOLuHIhveLmNRVNFxAtq+vrfBbqq88v/R+SP8Wd7ObSinIyxade
bg8jrvSvXm8yDzABBeWX2idwHhBaVszv4sPDfEZlDcEfcsLxN0V+iNtmMwguAt6G
xg9u6Xx4OI+lNf6W1GRitnZf2Q2wfgkj6zLDauDRc5smwSye5pfev7GXY8HAZqtN
7GdmG07j87yWSElud9Ingl53oFygr+jTySTPSyA4wFfTBO5NRDOIVNEzqTqqWF4L
9qfARdczu0pOyBGixfodkgkD/98OtoPVATDgjooMgzvuiyoelh5z3vqJ9aAlIvUy
6Gh8JvnwnImF4Q7338w9hL853vhaKhOo6ODcr+216TnCykWxlc94l0zv9zalDnuC
eP12XRGR7EfBgwcGMjOwSDzDFXxE4aZ9IAu2HuJzYKxndRaBUk8BkiKT+/AUw1xs
fxVs45etBAXpkaUHmd7ySBkJI1MDpxDJ3M1eDzUrq4IyuL3kv2gogjZNQnnwTMPQ
MZtB7aAtQbiQNXrU9Xq5AgicLqSJNs90CjZ9BPQpRm1toWnxXapPuT8EEAj6Qtut
vOT3FXVot6hSb5zv3ubLZAAtztZRXwZR76FK2o/NBFpibxDVf6Frlacau5Qrqlan
xz9eH84bFLFLnyHVgbLlHWMGNwrXQlzNvngtJ/X6pJxVTL1uc6gkkb5sl8VsLAyd
ATWFZEifkuy09mh02emmE8fZKRVNFas019+N0sySMUIWoqTL89mj8GTXUYWirNyI
FNzU2p3XEXADjj40x1q9Djo65ZBPpPjdc1yeNgIpfnwyabG9eeGOBTKm4Q1rDy9k
ufTOY0HFGI7Ye3plXDYupRJR+BMy0Cgd6GPjxal4sFfaNFGwuC1E/fvwHeYQljCH
Whd3lJ5MODSrMy1mV067QtpJrd0a5fJzoUt9AR+vfI507o1zDJD1YHvuD9X3QCmJ
kY8FWx8knLMPssrumu6YxZNvltVeFqHFrTFar/yTHCZJj1ttJkB28RGPxwzFgRDz
8mSIeH2jByCr3jV37CLfHf+OQqTh173DXXFBMc2X6C5SExhcHuTIuvn80xkLeety
CbzHQPA+PIa69ia0ucy+ohuVL9il2LRon8C4uNOfS/eigBArHC2yaoynuk1XCyL2
0tpdmJ2zqVjr2obtAYAoiYtn+N9lklTcWtxFLffSLrgv9M0JnTqQBecQ087u3LqK
PCEzAbpfc+Q6JOgHQwHcPipRDZwbJAnEbdnXmScpk8XVGqQsMGfH8QwHb+tbW0eB
PqnkGRBPyUxywybSDfMBHAeeHe6r8XPIrjjD8zlK1CfiL/LW3ma3TiJ/Ib73uYl3
QOZezWgCe/C4PL/hkSQvZF3K0KgJkxcfLPWQD+9sS4KK/DLGprM3f6a2gUGaiS5/
3rmHv5rL43oRVFi2dTTowepbsVZBU9cXCH4rnRMF/L/YOeOBZiTBuMhQvbBE1btv
8MV4oiV9G+t+Cl9qgaNMXb6+J9fc6ZW6m/dWXup9EK2ka47Yia7Ch5gAsibAA55+
Yow7p0Su5hG1Jw9CHg6JLqR/fZg9Nb6TqrYCufUgjZViHmJLkxuozp4HNluuXyUc
DLPEh/ZjstnDj+fgH7io6mDF3XVCU7+Hul2T36hdOTaKPP3oUr7ANCmBgAYvyuD2
lbJLqSHuKRJKJkB0dDVGAEyPcMRYBfG3ROlP0WoO5F0u2fSeSrvTs3GB0W0GWrvp
uxSY9sMuCmnhim7sj4ZtiYrisitX/31NUPVRRuMc1u2gEOGBZfTgBphYb49CjMuC
xzQ1T41+gZl2vHsiUcDRAxACp7vgEVAeRB6VbNjvNoSJtBPMeB/toGkajF1XR+X6
7lEi8oyOM/WnBxZF2ini2yPA7OF4w7K1qgGb4B8lpXd5cK6gkAxLTlXwN40YChPi
qisMnh1BvSkFEKvJnhVgYNPMYGtzyfMwKcNYpYQbEldM0AylZ0I7RMdCkJRFfYfp
sATAq2M/2VEPuTLbxLkfN2j2ZhWPQrVYOTy+oHgCKNn6ba1+BE1c2Pd0PM1wNnGK
Nx60hD/ZEPR1w0h7pgQHLrFSrxP/edCW+3M9+V8u9GUdTrAF9Vniuo9SZ4/4vptx
jm+RgZNXuRkuQNe/vCw6FFSyWFgqlqZwuG8t3LIgdYdwni0WP82m6PhXvAILlO14
2+x2gHUtcF2tA+DO6+wlcN1aTJmhG4RcGPFdj5ATW41utrl7m/NgubDmf+p3Hz+X
hcrFZjiqOdTsooo1V2lSBd4RNKvltgJi15ztJgXg67CvDQ6E3rCxO0WUKdfAC4wB
+Y1Oq6IOIEoNAQvzdb73I6yaGMsf2eUcfQOwiRuuSCPITQvhZ7ab8inXuRPhS+c4
bvgDCKJq8sziyqwtzrWx5p/FX6lht22838bpZj/G0bjQb7801nwbG8/qYBGh1mBG
HMugsmOaMgiDKe8R6IZcs4AmqFexvAG+VmMbFBFIUAgtqBBUcecrjYhMfEcbe/iV
cQnhDjCNzPHXQaMDRMibpUKgdeubgdKKMcMI/PnhfZhzARQfIZO9MYaq7oIvvYmL
NcpPfu1t8jT2In/9dxGCPP0pRZ3EEJ6XFsOwQY3cah+XA5/6YZufv0he/zNZE5az
X/+0lTjE2m2gFBXiDfsClDbMGPerMuPl84T6xD/oFkaUehLcWHkD6+t0iCI618HM
YzgB9/LxLmf76anqRMOwFytlgKrIzfusriJsyysE/0M/mq388tPJtEYcOHND5a3y
iSIRlwgY6HLujAqwwQ8l/a3OGGV3EuUf2xJ9LIt+uAstDEpDhMsMLoVvwe9YX6FJ
qryN1tgv6Jf8Fu+nGylJVsQYYT7fAkc7Rt8h8MyITbU4Ext9qeZURX+Bjdz9xd5w
hsxp/cSLxrrIEIxKo0u/wFR+E6K9DpAmtMI1Oe8px5J6QnSu95bLukDmPQGob1Jt
QK9nYireAPW7Xq5d9Kl/65IuEnJ4YhH9p4iJN1VSr/+Qo1NGKN801686VOszplR1
rygjXGVsUrSpFjUFAROo7vnjFdck9OURywUl1O/bkP4DDpQCoKvnFukcyAT0HlYp
fKJuSmVi2x9Ct6pBR430w1W+Qd7p0BWWwGD1wKBKM6CaetA1NtgHkzlIv+Bqx9XS
khQknPYex669hFIKmbv5wKbtfCSjrUs0lNnTBypARzoKMUaCRW1Mg4QpmU8ID/Pi
jERRf5xvAtvI9xdmpcuA/TgW/1gx0OhBgXvwLBm1EOLExe8/wXJZg1KOx9WlmZEw
8IhB6fv0l6TMdZj0CrIDEyqRqhB+1nd1lqHIbb//AaFjBQIYaudw7eAK+IRx/H1z
/XjMANH6g//xTOS2d9sdkEeSg7lMFz55Jlb7SraxbSZdqdsyb3Jk9MNZzNcyDIZk
+QMuu8E4L6vkbpI1S8QtkAa7lDkPoXzBiVWwH3vjE6F2gn8drOdNWiO2/IXlEAoX
6jBPVx20CFTogshMnj5+ZP+YXFqRoHjKV8s2vhXOQXbgb+5N5tj7CJKOw7FHUCUn
HsTu90GdZsTo5SgyfsIYIz+Tm4cyhre6g0HHndsxTMO8DLBum3w+6OHiY9GH4mWr
EYVg312bVogpTG+ynYpyB8h/YgoLrrYTcJ7sBkAn7Rnz4nTq8RSQbYj6Vy/01083
LdlIR/su1K8XPU2MBWmNrk7KCxCSoDTobh3B5Wc+JEIaovnQOhWxLF0RHwzoWn69
dl8SwN7RQnkF0GF0BhOHav9EPittT5s5oNkQ4cngGVXLu+SayZULNSj2tNPqf5HH
PMjjrXTS5GJs+5urSx6RKISvbOuPSSZHuZFPhqKgZmpSQNzQaJuDBM6AZBTj6Zns
vtYjntkxlD02Une+keH0nWwpTz9CV1s3TGuO20fvBYyCzmU4HzF05nLuTBCSRY1Y
8gjI2VIL+XrN+y4cSrVqlVvNfe4Dex/g309hz2xKElMzv3ZypgzlQY08SMkT6/eb
KHnzYWh9uaewJbzKW+a8ClfxwiFLoeBeM/aecskCCnkHtuXr9UYuAe/mn7hOOzVE
G12MN6/AXMkZuwaIOlAFULAT2GEVqLpvPvEQ2Pv8jICR4hUb+MJqTsrCJ3w+rVkE
tD2Bo8QE9SYniLH5SlwlpFA4huYiwrAqGZkvknvggC6Y4vdERaqgEIMG76w8IlXm
xApY13jpFnimYoKOlntZHxw2wjGvvXAmmdD0Xwqe5qBEShfOrYFAGqD9+fd6+HlY
nul2DtHAOQYRao0k+lY1Hvul9S98PRFpR/S9lIOuZ9JX+UmhBZWQpE4mVTVyfkhA
tb1K5R746LormeEZFjoarRbNRcStXN5Jkat6fGBLqxvMDWKZuC/8iRsI1c1GjMFN
CuysVwzUThkgV501qjy7cJZZf4XnnsfaEF2C2PHlqZVmlAkkskxYiQunOn4AzChO
zDDwcgjKMCcYd4bM17BM8vhUMIsaqFqPA1eg7mxW2fcBNmXcGkABZbO/4viunC/w
PQP/Bdn/b+tbPQRgclqIAFJiwDV0wPiR2U/XAJy1qU5/CUYGr8CIglPcERuibvab
c3W5trqlw1ZLFqVCeQ5c2X5P6Hmj/eNiAuD+1evT2HS7lpEA91e+yCNmeqqBiq/a
Do0f2jbT6e4ItrPwo16+VUriKzN4djfm+FnCKtjsFOUZonJ3FUKKLgf4z5M64ePs
rNNGNG8lV1KfuFkDXNhLdp47b8SIbTtM0E+GgLUBnLp5QiweOtVIJJHQ3v46NCGD
o1/zXDYXm8XF5vvJ59KNY2zTSYAgZKg5q+uz4lOYjUyYt0W+31OsmoT3343NRKrE
R0cFZMCx9ONqsj1drCxzW1IN6TO39BsyaA46PtQsHGHcth7dTxaz4yfNYuYrpHUp
0mMLiUy9LAjLG/K4H+ZP4EWhaiQuLThHqxu8ocj6S6qVexHM/FE/Iy9PDsHLjywk
E6v9/9FQ1/wPWQ39gxQXeuX0c/LY19INR8r71Jip6J7pa6m4/oZCGistuya8cVlm
WY5W4ybP74QKZ/VmoaLsNEDTL0apRqwW4cjZwKxd1U1FaXEVs75Mgk3Pjg6Zt/ZX
eXexV9Ce/9mKqZGS57FoyX1AL4U8LtggEnvtFaEL/6r0+d1tFE/0YZSDYLivixmK
NLAMJDdxm7CTUQKBPxuZgFcTFZZ+tyOvmXlenOPmxV6QMtZ2lCzGnjHcITTjwDbK
1ce2d2MNlLt1Z+TR4hv5RFa6qQZpyQk0+0Uqi0r4aLOr6ds9IzKcDU1IBUJzJSvW
whxzJyrWKDz4K+it0QhaI/l7oGhhzSkMWE/vEJCwOw0ssL3s9J884lGe1VhPHZ1x
Bz+qEUBXK8/SEzdm7ia9wFwuekZgzctO7zxMSiCQZH+UF9Pxc7EecmTuzghxzK9y
xjqZ+pFx9X4BPWvgL3I/UfxXK/4KbxAFuWAYjJRQ1Kr5RaVfyS0uSRNzEXr1eEhx
v/WLAZJDhJe/ofuUPyCTrm/wFpfYbo32a0X2MIcef4rxb9eGkmSl+Ygr6/z4CidA
8YdEnBKsDESjLiLzjfullm8D9zR9Vk3COGhIZoycsj9zO2Ip4ircQRsSAF+QORxv
3hVTRfUSgqYaFdbtA7QSqSeYfAydkni93gN0IWcz8mt0qeIF+vjzVs07LKjX/o2I
klhOxprJ0LdEgA8LnHhYfe5EJzZt0sqvw7Rrvj1xqhoJMjjUSpmj/mCt8UtrxFbu
0v6GOU7UBfvy0RCLTYhZUtxmAzuJJXsrGdToC7BvR1SDMVZwtAeqiMywC0YfxNnH
p/GAZxaa881EStgefTOMHHylYaO1sMEp7a/GMvVE7FeGyO1FWC9H3Djht2xxF1Lg
tYgkNUO2pRQpAL4NpN4f3rcqOLi0LjnE2xlLMlAUBBlyYW1Psvz2Y1kBHtFEa1v7
DYjzCO/+yP4VzS3L+8Wk48H+MvaY555tecB6/2wQKUwt2MkW8cIw4n9FMj9MUX5d
y8QOfy8ovzy7PB1OQRtPFG95KsDBLAHA3qDu04hmjmPQIpBBZjaqDdo/1yi0qOVB
rgv2egiSVBJsBM+5lmzIXI28N/G10SUxZDQYKpnW0z7lvw4k5SmDQJyVMHatPY6h
O/yW0qeEW8mi8nngey5iPws0HOWEdKJ5hhJ8D8sQao6QDmSZKOIDOYerbtgud0uU
g+txlaYU+HVMbwItS5pkXfPTJHQyzbZZyqrR9RIcmQdgoJjS/642fYK7T5LTq3sI
LaMGMrGN0wR89pJME0XlTvLiYY8phX9hMnAjMLCukQ41pwd1l+a9gCp4cE9ZbUpv
YVkba4+gNezao3eHJmQFee4YRroG9JXtW7av948iZl4oCass85fdMEQMeFp2GC7Z
Kz67OSlATk/M+0u6DE0aGCVTFZBGBOGIw1p5viVqFt2mFFMm3HTM7JYUb23K8UdE
BBr/0WmlNAStGejWpPpu5qmYwy+oHv4qguNhrZNjZMZ8j588Wos2m9y4xNELwY1i
ooNUFn8PeQYG8aQmpgNIFwtPvTkLYMLZZSZ0eiww0OxIo1A1sA12rYtRwg+u2SuD
yP+Hof+cbl6/tzJBIIeZ/nbULPuEuY4Y/mgzK8+b1bLOR4CuCwdOCRKIcwgS4fQs
Ob5yX9iBWLMMCIf8QWLsy1veicc4mCQDblnSMlGc/zQR8kofyeKThXzvL+gDXZvD
emnAtkZIy/6TgbAdbq1wm6GmaJFVeOyW0SXohm6dgFpHH2dKmNxRasJBlJJzwWXr
lGIJSqah78awB6eEVLCPysVu8bFVVKgkyAvAS3+8Gkdl0prRAE9czxucq6kM2Dmi
tgocGGd7d7BMYCwERI49Nro5uEa9Wz/EH6NVYZaCUtz0vwktl+zOuL8kIwxty/o2
8q2MLdDoV5VSEZfK8Jwht2Oog1OtFmtG+r4MOkS0829jUER9CL59ukRGV/mYKeJz
oORfvsTRSZaZ2ocdWqQwdiq7KBxYLuku8gR2X+2caAVd33uJDBPSqzipPDmWlcZl
J9AtzUsK2ivgUlom63qdaUJ1FExUYWvodhttJxIspAXp1UJsyRDWYcU7F/IZNNfW
fIR3Io74m6+fT4P2tUmHINzbCuVZoJjRnUTaE/NkN3w99Pympu9ttEaFsgP1n6S6
tlPEJTgUQ/0OR1RAcagC3grMv3RbXCFU1Xu+tn2/DJ3ZswoyEy0cjJ72aW6Iip/g
wl5d1MUEqqhQFaCVdSUwZ3cMHOgjn070r9rB0sZhh50WSAXn7ffwn8pBVVUcQDGZ
Z90+lzHD4PU3ovoCzwuxv9JivW+N3Liso8zz0NL4dV73Nti4xjfMbhsyM4uiydTK
vSQj1X05QDkc/1I+vBl7wKfCutpGCCpaFtZOhxYkb6ezZ1z2/z5Pk7S4uKkrc+kI
En1YH7yl6sBUNsMkg5NSbZV0Tc4zaKrxwltQXLArHhMVv46I7TIOQKg5o9jspWOO
xzW+EjkuBa6kcjbs0B5MldudrMH8GvBkgQsNcJImN/XjtAVaXBeJl32ueQBXTiGI
Y3KRwKg+SDkQ9WFl4amtM8HMnGAlj5IjuOep4EjiImV8bkoEsyHQsQJgAOXkLx98
1Du5lGE5loXgwwRTTvmvAOThNL9fbxzNdhTjcp9J8hvz4YzbQ0oh6f+jzOZQpaMP
vWr2EgUpbnvFC4hDhw7SwNRN7/PoQ//8UEC+h2oWTscsc5/iBD5Oz94CZW40p28L
6c3g1oxqtLL1kXio9q+j4E9uPiBaFxwmrgTdzjhuqTo3dpOrz08dlD1vgiMREgbT
bEwJ49kmuqLlabhEPEI8R8uW/f+jmCPNj8nEOjjIaaKcghNPdLawfpvaTPBaQwcA
Um/45mxNBnpywUdE6R/FUf/zlCtWwl+qyy0+CszdzzVuRjmRSqB9Ylu52zRJKc0j
Wr7kC/m4WuXtTP1XXbkbqEdVPsbpFbxm8C9nHnsOUMru20ftsbyrUDbwbRvz9WqZ
wo/Or7pfRKD9Xeh/VE5qN1hGIGzaAYe9mhm78CHVHrkTjuqoAY0fqhYqq7qmSiXf
m8gDKqlc2Y0rtw4XKtUcDOt4hNCVqXr1cgS+0L8FMplWZgjB/RkOwkwZNtb+13TW
N2RLWgwR/WrthEv8dyZF4htnK6ZBJQOOaXEVIn1bcDf3XzA/TZbpcaRdsOmZzAWh
63gSy6Yp15t5+CsqdV1Z+fHVZorRBqacQ1ZIQdjRxu+mjW6+aSuY6pGLePn0WFlf
oV98+npP2T1j2X8T2VC2omjeCzU3UbNNMOx0DWZ1tFw0DYgWQ0bdb6we1U83ndZ2
4x5T8W/ZofDtp4qaONiCAWncaGzOSunRwPBqfdSBpPVP1y4cT74J9il/VpLw5bGu
tqpk/57fF3jHBQEJ7iRPgX+/gizb4x4MT/WOGIE/UdutczSN9J8o/htniEe/foIZ
CLA3M4CJgN8J1v7rySmVACvFlDx8fyVLge//eaXAEJVzt98mF9yCX3ne9GN+Saa3
0u1wES54AsM17ODT0hxVuW6Q1uIaxJHZQeDShB/xVUmrYpVFw/kmxfIzEI7iU3jv
o5kNSLGvLNn8YN+2G0HS5lc2V5PfrmyUbDZOACW3jWoO2smPoojGR6PWabEFDa3h
vL5QkgMWfqTuESw+yTveYHLrk1o0E3dlmWwKKfRI1MLHTOPi3IL7O2fbq29ayQHo
EXCCVs86o44Q6lJb7Hcu2aWrXX9thHhcKhVXQxCYO4+qmjAFc89ITUKGolGozmsc
RibRxefGF/wrc1koJpsoArxGk3StoqhYVWsWHRD9sC3Hf8OMKwiyLA8Uwn9kZRFq
uFJW/D1dK3Pq9zOiRRI2+bidO4gLx4gxopNwowaKWF1uvCzNehHi3x7VrZLyHXpx
LZ/P1QYYlANWKoGiyuf93zNIF8RvLGd+LhdWE41c4VrYTZTAgbIAzWcv3SYFpbmq
sMbYRD+5Loj/O624j6EBeG0Sn4aMpJHzJgHRbGjFK+/k0KtHfLzJSlUf88BKfk0g
7D94AjjGDenqjtZhTnYTvWdFRTdIBUyQjax8XR9xauJGAJN5DOShhoFAyu5STmpO
ZSkXosFOwzcHJmtuY80Tj43StFYVXV/AsLPSCGHS4RsSebN/xQW50R/HGlbyzOPT
1LQAW/eQmJLMPd8QXssT0qcyjgbP+Vu2tiVO8ZIdjqUSZLAgWATHWJz+p9eKOHC5
TiqQzcL5yqC0WtWHDDrw+YmCLUsm/jpsjLGAKj788eJfCcSpQ446Fd0EYH2QdskK
e04Pk25C9pde1zw7bslG7Ri0hU4PbswacBQXt9XlKc8rRE6kYMx3r+jpOP8XweQB
sbN0kgqOQ+ORyhaTRCVSjnlURkxbh8JuIPT3lC5yLCUhMNEv1/KdkBdl2NYi2HqM
kHpjYswBUGJ9x+DUxyguFwL/mhACZmYfqHz0YpuU77Z7MedmAH1XY2xUrczNZmHh
C4JHyXT7hRBgofczmeKqktL60BO7QKtA6rnWUv2m16O6PHqAUbKGmIFllRaG8Wko
QB47+f1JMw078n5LHrXp7IOXFkIJzJPIovRLeF6Fderx03EtIcUdZKR7j4XGjzbn
KLblZWFiyI46IGqEpcTlLEhsiFj52Ue/yUijtyriSXH1ESa78qS0TkTtF4aQnlWu
fdtMJFWyr8r53Ohb7ldoy3Wlvc+3Pw6G61ASIXeCUe4o3jr+473r+lBZuFoHuhmi
Q8z1Sf8xhyODINC9KGD/YtCG2G7yZ4gLc56SbHu3yVLhy9UTv17Irs0PD+9545zd
bkzAt0olxlP+BCr9tARzHQ5QISECfzwRqBJFfjWCVgh3Omnv3x68j+UHHBeh5bdA
vxM2WgwpgPSc3gsJRkVKxVrD3CNLA2Qho9SbpMTI2gNxVJ/AyCaJce7waFpuyJCl
4EP3MQlsRfJWaYTCX4QWjoEqs14Q4D3oFrEaSDtt+hvlahdRx5Dajt9sNwqj2Nm9
aVlQsYnMq64eCR98/a6F9FYVw4ZnZj1Y8kr8iw0BgMRBvWlXT11ue3vTBz0XINZ9
/f5kG4D399CEO92ofwFLHUYod5NxL4ailMLc6kTqCgWsn/O6YSAs+UeKcu+sVAev
vojO8EmUgwkS3meRUYX0u8sJ++LROZQ0mPRSnDW9YxBkmJx+2npGssRhMjq4vtAt
I/DvJ+o3/S9Q1LYqBcLKMBHLF36XLmz++xNmcpW/Zl7IBNzqgnW4fIFeUfGE2wE2
5Gk90wpo1tgYqdcgMytQ6BTeKQd6V7ATJrJ5VzrYcOmAZ5xDgLCRSXK15fZXHl5g
hUeeHupmRxtMwC24t6IDnJCTZKRCVPduRa/5kBobjPclgVhznalouni8qMqE/2RU
DQ5u7u8stORJePlSJRxbmbp36EJz46eNa7qwjDcyeHsDvVBHvy2mB103t3IA00M6
OgtzsxwC8sooM3CURpSA9cdeU6RIS8iIxd2ytw+OgvDkQHfV9OhKcqtdZsO+a1Kl
c/ZhSSH8hxEYtaYHcrSXVNy9O/ofctxloWBOfBWPz4Da8uv45DZ3h9gB7AcvR2hq
t828PbFzMg8W0aA6AL+dsnbiT0cEVw5PWl/HB6U4shssQRbYMnIASm+QNgxrQU25
yNX7PIBsreBKwwjYZayqrxXa29RJ0wadOSw1bJkTbzqWIHfyxk8qxqlKPaYaJknb
A7u8H9StvWLcnbfHo4vgWLIA5aTMZkXHe2WdiBmvx0VurA6o2cTc6NbppHJacgFZ
6v52vnVk9mVQ+VlHKc/pJHzWuFG74iyj9A7ZUMvz4TEviScZsaRX3s1nA0TidJ3O
kzHIIJa0dXNe5FF+RtMXUf9H2t8YpH8DgrNV4EZtrfXnzMZHAlUvr/f5DWBAsrbG
upQBgr+4F900uzGVIiPI5bNnGffQKWFeIMl0dlSjxzdqMz8Rfzi7NYb2jpGrpzvz
8+KyE+qUen6nzuDmJgXFGV4Xh7I1epmT63C5kwJZZdypvnz7yOp7rFwKJwBo45Rl
jKIqLma44Cc63uW2JCO+mEXrcFqDz/7tCs9UMzNxr9qLxC44sKqtjQiWcVIAur91
tte6VnonhFl9LE5Lorp9jb3tGSBu+8mnQM8+nDuxM+wGGabRTWPaG0FvUkwX3wPg
Iw0SQMXRjlaApP+KaeNs+Zp5k0KnAgYNhl5SlNGCiIM6PPBY6GQTC9Fu5FgpVR5k
MbrGJ8hL5xfq+M+woEkFh9rQg4VFeuwcGXJrTdRR0p10Kpf06V+fmKVuPsPsf8pG
hd73ALTtKVqnCYHzYma3oPgNBouR7h4SKo9ts3HvlqntPyBg5+7imKLRyDCRlUgP
NeNRTCK3ePLLVfJfiFshpKvFtNUy7BB0LyVLuKMpl06+mIARXIunv6jO2HHSKQcS
OkVWpLCNyWVesJ/VTOV4X5Pjuov0TjoOenpWJ37UluriTXJLbqPYj4/Gqwkh2n3f
IBG20PzFBN1Nzlvz/+0lflgWUDW8BjpNDTSakIm6dnlwoXaRZPvk48s+Zx/YhQHz
HhQsUkYeB8e27Tz2TQkiDqyYeGe7qrtC6AI7iaY5k57hm0VieVaR8vmzwO5ejs88
dkVCzwJB7J98AH/FkAxR2vTXq/V8U3iD/btnycIRCZk7mw3jG3YSUkYxeudcmQkF
bWZ0gBnmOCrx//tMrFQnAH6JeeUfROSPTF+JMB8hH+cniXzTLmR6yo3lV5tO6ej/
YPt4ocDj7KSJS9ItsZmLzAJTDBMXsq96F26hyvZZzc1S1VN4yC0oSTk57wninCMW
skv0pT/yaGtju45jqG2vtT29BLx4qCyMdMqhW3NbjAdPAk8O2IplXkm0CpTF3ccT
1BqtnZMpaZnBDGqGAR7HAtK6G/IdNZssncohBmncuFD4TZ8/0GXb88dEmbeZJCCf
EfszOTt7HVgEIfH8GTy/c3B+CBIfqSqnH7c9zmBQdtvmCQcz1OxMYK8w6bS/p10/
16+HrMgiuvYaKkhKZdHU1OS78gLzknX1wtzAvYMLRfjtlNoyt+G7z5Onta7GmSyx
iwChiIefVmAdoumtGg2RhZWWKrqWtMbadNCj5rd1LYdcV0UXxaR9qNV9mrui+gLF
MmH0sjEutRswe9gVLTQ5B8ucKnVe1jJYtwUeunnDMDs5N8HIJCONPPmTQeeMp1pW
myRQ7ssxmMM98C4aK/X7G/xfYKb+9IYrwHC3CK5N2Gy7EVoQ9dB93MOtv0QrbCwy
JAk4x+Q6QpejeW2amvcD83pRHj/6oFDCWisBH21dwjyEs8fh787FHkvHj9qrDDL6
f4Gz2VfW1I1H3hMtNY89oxWJEpEpN/2QYs92YkpBLyuGSLEVeq6EMyBm31iNHRjw
IOcxGR6nIqJU56I1PxGKNCpL47BMBCfS0ZR0nC6rCM/PgHyig5wo/8VVLWD8rq+8
98+lm3XwkvN7E5E5lBFEXWCT5KeZhzpKGzfw1qpynrYj4umbe6FHPLpfaEnGfdfe
6TAtc5eKgEACLzXzqhCVO035RuwFQ8h8139eNj/P10u4Xza6dRHs47c1OLgZZhPB
NUlmYybmH8lqznekfhewpHFT+SuWIOHjKRWfb8i9m7vRXf+HWr6pkuvIKeQhE4L7
zJGp4KNUX+NM6VOw74iOk4O5OU+XCUz8EreYI3a25YVpPw3g+xf1wstZdU2QugMe
h3qGc288HRMzf7WYm2T0M+DzXuXU7yfCcp0+wZAJO838D/EpRLWX3IYwkZ5UDhhx
7ET/UUmcklIUnO5ogYVYzn9kBSXFrmrsPxYB5kUoimM4HXq2H4kd/qPbkZnOHIiV
mecggK6wLSNEZtDVZ2l7df/jd2jerK5r2ukTkyPxFBcytPrhe6ZGAjxIe5xybEDe
BthkQ0VNTFTIU9+RoOLDeEwJ8rVXLALjDFHm8KwESViZxwaZlMJhKO60UNrHJUIs
lO5wsyAn9417ngpXaWqApMh4wLsKp1Oy+q4XnnO4D5jw5nt7GC4Q5SWKzKqBMEKB
ICKVoniWFOUqM1g4s305M+dmnhYU0heq4JulHTpO77cmsix87OP70uQzZU74Ofc+
lIIiMoh0QGY5q4QhOkKeecAZ3e6H8eGjjLBveoU0eTOtQF/WW+W2YcpJGwJ3kvki
EGz7EIQ+/SkNj0Zo2XZChTyDnYSWbXznYp7zCVdHEjkl0+4HCmwh1KdcoEDQELq4
Z8h7Z4fseNhHBoQxY3JSdwLQ+KUqQ6blakZHbXGcH9DQxZ15Yt7Rh8kEHaea1qpw
nGCuTTzC/ciKJsO+8vR4GZMtsmRcJfTWc3xNpE2WNcjA3kVo1h8Y+iVJlzmMQU8S
MRX1RbN9GHujiCF/UcxtFIlZlBP2GGVuQYSRU2oZBLohTy36BL4MvBGjshkdY2pT
lElbIUrLY8aDkcHlazmQ11CyJ8Vez3GCzbulMfYJR6ge2PNoOIfxY736HpLTgP2a
ci96mTnNIokYPMkWjLihMMrKA1bJV98lqFuPjaIoCJ2frsblTQhhUugzaf+28YML
TTRod/3oElfzobAo9Ox7QEeOovHfACqVTvC6dAXuEiufeZJs30tKmuPMmXpyf7b5
VQFC8bSLKYJGVtAIrEscZ8UvBX/eUuVM4eDJv/kLNz+u0o+YAcAwVYFrp+B+p9E3
Xlkw9xPdCV1WvFOxvqRa2LxrWYXF267xFG0RBs2LIr0tPvDpIe1XWGtWdyXDK6U0
O7Ag4ZKWvOj3f/stQ5dmTlM0eR2mCyVaXhuPJi1YHLct6izZBCql5pMnlQegv2g4
7tLcFaDhr6j9smrZdNQUB7/kOzdbE8beyNYrXWjSe2WJ7h6mYRhbGiMMmRgnfm12
Is0BBe60bW57UzPAuzFqCSBnEfy2w+rYs0EOjQHz/DUyST0xhRiqGf9t6sK6f/9h
opOJ9RMaGCRX+atOF62wA39r8CKPJhG/O0v53a3GUzeEsv1hKsMdPCC+QldxBmI5
8reixGtcpVEf0ePa0y0iN4GWiD7nAQxV1nM4FIB9BHaQ+oZ+iq4uQ7enl+Z+IsTQ
cP6heRtyk48tfPAR28vW9CoS12ZpYf5kP45G4ER/0inqKMB5JEfxTa3TtvQ6syS6
fktD4506QnSsiHLek3ODAsnMVKkrhkO4PGMt2CfhqhwTIcBcMBNYrT7twr6GfT6e
kt4I5A82jwZeQRPm1C/h/baksOwZZpJeEJiYtho2KPcTqUtI5qW2GcY51l1PhkOZ
Suv3mCk32PigFnD4zZM9Lp4P3zsP3DU/nQkMENsroJJvarYxvdltFtE4f3CzWrhM
FNahQdqmucK6GMu3AANz7IStlswpZAlfVW/1gN0DgcvqLa+CC8iOw8lM9iLCTiN3
lh4X+fAmL90rcGEwMYqW4AXTye0ltTvEjA1/4jXSUDhb5FyKiF8k4BQcGcMJPydt
14lLRNAWH3RWSosEHUgCrvZbafIZe/lDdyc5re+9EblHkixEFlq3gPhckVU6ydIz
ZAZTD7WLUWmFxausWkBKkx2q7Q9PWALNBPjb6dh2F18iaaIICjbE7vY+8HTNXGLW
BgUbokuAnCzIM5hIaqLeblEFw1ySCLx1K2t6FBtKfcuyQj1875RNbWTbh2nEMfHN
hnzRXlGw8SeAijXRMF8BqaCaUGpayQTivKITUcsUj2Ox0xJLGgwYXt4GhEqMBFcM
Vfx9RTRs5TKQYf/boqZJdUGWgIc/KzQxLSFR2qg0m8yIHTpp6ptHwprVyTjaLHRL
CmRc1193F9b+wM9MNcPLUbwWqRz/7wzc513iOtRGJYNkalDB71oN8eXP6JQms/m6
iv4BHAmfrA9X2dCjrAMYCK9IaooA+0V0OCP8GwrXfi22Vqqx5L4oSl8iwy8AItPj
Ncv3lJeyc/QxYZ31/npvn8tDbFaBJjriG9EUUoXKwbTCcklPu2Fgb1KDR8B9lK2J
C4t9qW6HtwdA59msxVTHguIrPJOt+l6HPumdE+49knrl2znK8wzFNeG4qrtY2pPW
1cnYnWDvwmumpsydDfDFz3CmOuZFFmN10I3EPT5QNzudUYVUl9IJV9J05pQboncv
2EKyz0LKGIXCgLLQhLO4Uvs9GnK2KTWY19ArPTeNKP51TMfIsAaBpKhTN9ZHxiib
L0wVVdVyh0oJEW5WqQW6CyOv+eTYvQEwjHRqUI/hhB/0giMXXLh+/xHNwmJJTh0B
fkq7GwyG4/WlkDxR2JU1clk6IgIescPrW31QYDv6Clp4a+8Yu5GRGyl7LOCTh7Qs
5EzO7GEnviJjyOl7S5NVqg/dzkjMLEwsLewm6/ZKQwtigQ85sfq99KW8jnyGIGkJ
3EMU6kjXe0bwpqfcj855aeJwzoB8X39Im884UHWMm+lu8XxjZs/5WdAj2ehkQLYo
GP8p8CRX/tWDfww5RlcyFZcqE1ceD5pqMpEgzbpNm6adlslPeF/N5Pj8Q/7IFyRc
fdqJd1cZN50/18pixgAZ2qlSIbKOkzd3iyRx24hHpBleu8RBpPwuHK9T57XEJPxV
d2v6V3CeWApGZ1I1n3jwVdetuRe/y3mtUJIENO1ybZ93xqLDMrmXgZmPDB246UaT
y4XQkVnveU5VwhdsZSGvfUBcygn3eopxHPB+TkKZjOzQ8QLguOb2B1t9iTZ/BQmG
OD9L5KjESf/PM3GlUMLNXcwSloQ8XEUc9R5k2w+YZT751ec8N+FInyJ2eUgcfIJt
t2zSGYJM90qqko9LA7VURUIatbuKkKyCC3xPP+N8TIqKxL1X/CizWoHaqkGVah1E
IlQaxrM4PH48dXmtrCYGpEHpQzHxWmyylRYlY9bJWTMu1D5FsjNhCHsL87ADb5E7
10HyxYwsfSl2EiMTIcl47eMTLGFDFEhR6nZ7xzMYksRh4LOLbzzsaCGzVHGrw8Fm
Vk14cvwIv6GiGPMQ4BvaHol6a8NtFNuWauiLRm1aULYVjfp5FC64ogMjknWy3BIl
6krYQ9BcC/pX+kbZ8XwHDyUJFMbrnrPrpfxFo15ocUfC6Fl0wgZsXmySXjwAOpRz
ZhS1V5UWqyISAOPedE4DUH8JV8t3YAd4kKJjxHjbw4ZjHe4Gpq8FiTYJDQ7eU5pI
AtvebnThiBgH4yuSrJjCKty0EK6N744rFNdB4IiGFaSZOUX3zg3SONpU+Spt6wfY
yIftoBzO/DBbVWVRXk6ZK0X64MAXFHaSCaR1lqPVLVIqMXjD6+Gf5djWLIYZ/RoB
+5iJwAabF+nQnSAUKKSwB8GYIkS+ODGi/I9TopG/oknpEG9v93F1iulutdWpnyiu
LQxuvXF+x9D+Tp/gOhnlAI06MqSbv4YRuOGIJhRkjS6F919KMSGfCe/gVbeCHSwJ
cL0xq17lPjkpjjKrH3Jq3xD9077TjopwMDggrU5a4c8b20y+hzryiJYCil2khxzb
YZJ7UxIMlzutWwploOYLaJ70nfoNETJfvPOhUhZtXvKF2/JdlAYOJX97SlPTXtqG
P63DRtsMvRDRkgmTxyEgb+XV6qjn36R4sP/vHkCz/X38KRUMgLQBP+Haj/WNcaYW
0mWK8TUQfadwiXTuPNJNwU/0lhJSRd4brTz5oTxHm+56sODrTOePCa4u/oHgcfpU
DNSugFg0IiSSy8f8JFoqOgZJmcmydlhd/IbIEhdnLEQ0vmVQerztqe1uG5Y4D21T
KBUNMFyaZOGHIC4Gwgj2YZq+A/mfyVS8Us9BaV+3H0yRqnLlyQhXSscFsluuXvXn
yf52arAqbbEQ9I9IbFxU1W+qtRffPanU4o6UPgZX6bQZooed11GK6IYdSWMgklu4
KM6DJN8XAeyxB0u6C4sErUDkoKcPRCWFP0d6TFGlct+hbBX3e/xYNWR3F/4Jefsu
5Ckul9+Eu5//T6W4Pd7Xa+HXpqHfXSQfL3lzpVsUSz2K62dBd6iyF8WnMrgtLY2b
L/QI4TPwnqpGD2wwSnRMo39o0MDcGj2G55R4WKL1a0X20qfI38TN9SUXAdgxTyul
MRm+YoQXZ2OOA9zv30BQph0k4OwHAyGDHctnOFzaqYu6B5C6hFN89SM8t8nX1iDt
xerUxYAfXoqoPa/QlLXAz4DbZ4SchbLUldwstxq8ZvENQfZTOQkqvcAIHOxlzUKa
oZb9zbJJi+HTKRbOu179vyB034bgY2/XXDxC9Tav/M4BYZxY9ULeLQyYlHinwbCI
vdyXH8K71yO5bN1ED1l/7t+OXEQXj3kniYHsisNFSzKxBeXjkrWvQ4O6rjAhZOg7
qnNS5mmDivr3mGbss5XQElmAImgD+YWBqC7oPuva0n4+veErQPUU13/MH9bjmJpR
5gZKxoEdVF06nNJHvwmeG1DoiqluJvaVqVPyKz/vGioaWjEH/NtlyQTohJlpeg4q
KJnknTnMSh5AagxjEJ7llkJ9XRpQccsMT+rxSa7A82qlRlXdl+sIfLQa/a/AVHOy
275vRer2+ndo7Ru6mIjKYdbh3bNTb4WBQkUAYFaFuNck/Zo6aLuyzCZRp1Qz2uR1
/ZFP8tJnrcz3l2FQSFDyiRrZM5naGcse64IETvFLRH4zfatvbXs0NHlHrKJrVvpE
elD1xYhh5qXFJnoi3c7XGj41BiYVAMpJLfeJRuBH/W4utkA/fbRm4Do8dQ1Nb6ds
6BbilCaspHMP8Znzgg8jYx9lW3xnZWAKfVvKuwnWnFukliY3+FfilBXRdkOujzQo
phPCqIviWNYP21r71XXce8PtrnLcpHI0ZRCBdZ7FwYsqeh8VRPEX3nXCXpGHm0Wz
i7Ew4QzkTms3E8xoi2rwAV+I7+/5PWIzOOu5x21NLZAnkmDMvobhZt2dzKCd7aK8
2zgcAXtkL6ImaY0caQVTLk7L/C6wicbHro+1tKbvbYHj1imeQ0v7XEPTtbmm4TVi
znmda7jBXT3bMdTVX7/qnPRpNpG9pFudBbJXA4+TSGb3o/tr6pKHNnqaqlLYt9UI
E/h/f07tu0r5FLUZ0t7dnpuauNzDFIqR1dTRLk3pUKzfh/WJKHAdmyaGUgyTjq+G
/vb9cVvKNOkQrzG1Wgcc7vm8YGYB7CaBwMMc2mX63pWNhKwujx7Ua9dHP3tO7g4x
OLoZ0AeqP0yex7YrX+kdLXuM5DrbAOk39UTY5u6k1VS68oPIIqlRmi1gv0OR1CPt
/DjekG4gc8jt/jSbdXlBeU5vtYJYvGeGEMs3NkDNyCgv9z+HMyEcYWHlMOmamAIM
mVxG1KnetLdY6fVQV1GToQ7Yjh8A714RdwTdc2BOy302+oEP8tn7cp865JEA2ye6
XGoERHxrrsvZp5PYaJC10WCU1A9MCdQEjNft7zZZDDGyDouEOt+gjeHKf/DM22cd
DeErQMrnrv0bB1hu1AoVb+yX273P/8G17Hs4D9D7pZpqFQTTRki2IuSKX7W4vbAz
CnzSGVChp/5FQafbyTvbYqUA2Y3vs5lyl2ZLd07xFqXQH3utygkMq8haLrujz4aV
n46SwdAIXRNLWGABYl8Ed0mGsVThsxUBJq+reNFCoGMINWVQagmxYkMu148Ma2Jj
jttjeAv6HqNrgbVH+DhyzZWy2/K0EwSbA3FHvBCLY5azcuxfpffzGRAW9K2tbVW8
OAN+prquLiP0I3Ht9x8AFSXvRfXcewblGQNdTtDNq8kljR+jgKU5rMBTJlAHXoIR
eewnxnc7Qyu8olstk3IqybKdwoXpvAzc/yGjLYi5s3TsqiL+McsRyjOTlR+Q6TJe
HQn8JkzF7rPS0nJKfdTIs31NvQEhwECTClP6gYJLYFmsSwGGxqPQSB3SJ3zlUPnQ
sDJOstAYyTdRQGqGHN44h2uZx/YYKVae3ezFy3uUUdQJb5btvXJ7TKfzd1Fa/ujF
KaSeojOdrFfa7uwteTbAHq7D0TNk3ONhLdMAXnDhkxugAUkX8k7BCfHiT6JEAsxO
WXdPRiA+TtStWwrV3zMMQty+7p1/jhawq/ZKpl2qFYzwgJ6sW7LJltdxhMIox4UP
xbVV+fvfpetUMDKDzXYkxWUyRAGpnynUETTFzWMvkaCMCX/jyDK5j7KMwdoA64x2
gj5z+6b6pV0e/xOdVgfKLBtDuCjIKd/RhdbWNw017dY7TeX/u1bCXL1J7fcPywuO
5Wi5mGUen5QPaVJb+FlXxNcNuxYo/UskbwTcqSNiaSMATWCSax+9yrS/8WXhf/rF
84gOMnoN7twlUgk3+l5HyzVt12TRCMMr/qY71Gx23kEceTSUJ06yZ4sENuT67XIa
Ur0VwewPqn5THBHsfa88M6i0mGgCbortI70BM3fD6dki22iXVLzCB6BYPHQdzXgy
0x1NZDPPYwoCYVRbCCcr/M81TAl8HqxNiy57JGS3l4iB1riFLwO7BZXMDgudsYVV
ebwhP8sQ7PefKDtxTESAr0wkhWG77s4+5XTFNk6UiMNkkZcRTHROwSh6XcSF/h8f
bBQy/g8NuZtcWFv5AGE9ppfUnwSQM6XXHx2vNQJR5+K3cEceVXUYvny25QDDHysA
8HA84Czc0uB1m0wxswIF/T0xQA89CoB9H+4/wDo5jVrr5V0mRPz/Zc1Mvdx9BG+H
8NgtuKNhKpJX0lwJ7gznnYCIWtXoBRAsbuhxTB5VXDuUs+9E6mptYjVAOynRem48
ZX43i6j87/gEPBFeJY7VFpLDgaslEymtw3SQDxuQcPIvmzyvKXR3naDK7VVAd23o
FP36LYelswd2SZCsHTXOwyFtAZmZI/oUNNnEvK8jFjLB7V5CWsTtDFl7ZZvipdvn
2AzWiSfWjecI9iVUvEVmEzKQ2BuyjqSwBUGVVA7AKFykIDhW+vevp71j4nkDOers
SRY40r2WN73tijnA5T+kbaSYRK+awkvK6Gytbl/AzRu+HJ64pUjD6fUdIYlrz8E+
y2RgRudOIl9AEAf1J6QEYMJfeUUs9sRC866gGT0XoI+eP1s4Xmbzt8DYKQpbcMIW
oWy9DHT9WhUzQ+p3nBSTHeTnAXM/sinEwmlGeLpXoWMd9h1FldoG/XSp97IV6OwK
X8MW+9hhF6H8vF54aDRxuGRPcyO+kVDWrdiM0MAfCZmt4fDdmodiwaoOyifHjTqG
kiUsZRjRTQpgSQ9vIvQ0CxSGdUPwCkEKn/OZ05YL3cLbWyi5qiS0SpOTsJ8kNM5K
tkGi4AKyPD/dltBspW4bgDpWkFM4rh7OD/CzZLvhphgl2qDcy7Ga7aZ04j++JP0G
JXM6rdBCuchUahuZWPmzlfa1NfOIPbnabmaDA3DMWoZRGDKbcEzDEaOAmzmwhJMz
xB5YLrkgAI42SdJweb+pBtY340ZVricKE/C8bnJFi3OzN521FVKkQRqt5DHchAPS
31hz0oJOvaMxmrqLX7S9Pea2nZFRa74cU1Ouvpgg5iJ7bZnN3n3QG+PkPwkJxI06
5DK+BimkCbLU8ekNmiroC/hBejh+MVatOg5opMLks2wZtCzJdhZL84WT8CSDRghU
V3pSgscYKBf69lrB9ujsijiw7vq78N8HXhzvJsJ21HQb7xV2Rhehxl8fbxO0h69S
w16fiVzVCSGuEQ0r1U1DSBSj7QO5Mt8qKJb6rzrAz0AEcVxzrxvRlOwDNshQ9wLl
fY3iy0daX6CzA/ApbtGTBave0NRg305NaSjwS61lvB7X7xjqAXrgS4pKQOwliQ8N
nhV/TyyiTHHdJ3EW+yaJe8afhJxk82icFx3twK2qeYvCRK+/R39Uzt8TrZfPFbYt
u1efiGFp7H63gGPziPeJ6asDcjdXOzxChl0UzfQlU1fx2BphI/ga3dWQ9MBZrOjY
5LGtBMFArK6dG3z6eCoWEz7Zwuhy/IdvuYvQPLfsZDHgJ7Uy2lwJJ794uHyhVcx1
8G931YTcPTKvlDh5e9L1GjNHkEtukY2IAxJg5rM/YI5PBm1plvYcf0/IzUt2T+0W
hONGQEOmPy0mRYOBfav7JXmDM5lP4HonocoqzY6Nqw7aKwMV7EbVaTxDdQW6kTFg
o0m0IdB51Q6SBC9WF9ab9BEqks+aejdSE9JVuTWYRp3U0y4+k3ICXG8Hdw/lgIVD
eYV3GWxkdqt63eDWqmkTNfgxdDrc79V+WTAj7CmwXl8vfQA4c1P3uffKhZLaXwUY
CT7eYTU1ky1Wo/iUN8FrgexwYk6bbGsII2Hli8xWJ8r150Raw0Pz2KDBPXMfMnj0
5VHNhp8BHFQoJub0SSMbDkbAWCnWnwkpLEFVmoAh7HbnBcx49rEou4f54pEit5mw
eshDynxQRkhGGzIx0XfKhsWFA921FpWQC2wX0wz4jCwqq2Sb4ugdxly47o88rhEC
ww0RG28LZ4Ab7UPnTDuujnd/0r4wB5B/XkKTrSJpsBi6SWWnmrQUIC/eI345y4Ny
z3FaHFzOVDrAusd1N3VQD2/mhkSavS2zS9vGE8XG1xugO0q7O2Yj90KtTBpN7t+Z
VtPHPzXdq0XitS7S5pSNIWhL6GJZJX8Wm23u3XvsLnRLJz5wpiU+YJiX5VViXxuZ
x4VwO6Pf7Ynveud241g7zCInGlLw7FPivv26ynOvd2iAe74dBAW/qOoITcvFbZNH
oFx8wUA3oFe/4yv7AyUfJ/scbATGMarejqlE90jbZZQDTYs7/E8fn10OLveWLE38
tDDJZtqhFFZKLgva7lUpxl9JHKqM/XSJ0l7NXMAz8h5RaHzk0clK57t8oIju8cNY
plfoE33kIXdXkPZAqbiGNWAtPxo8Fz9C7+TKgSA9ukqcUyT0+u9xa0s09NNq5TM+
u2/Bmj+u/0OxuwLfXTYaMD3ClZcTik+IvWLCFf7E/dXfzL7443TLAztZ9T5T+EH+
HFND8R8BgjAPBVQx6PQkWg93ZGXnllRL2kF3bLJeqocRE+JuG32GbXLvLAvF8n15
XWsmg3ZptKPadNxqa4oCoqmuItPykaam0Y0QqndyJ/DFKtDxpEv+NmtHbR/XPakg
52QvlkMGony+zJxacP0NQUE1ivQ4cax7OSRKrWIeQbdBKi6Kt1xHNpf/0vucmqlP
BKj8zNbcQUCNhBoo/GSSSlTPiJ5aoOIp8MCG+IHAfvi41pAduSBAKPfiHZRrZJLX
FIEbcBmNAAcsegm6SH82To973KML0DcsO7yflI8Ki6Oc3Gs3gEMhcw5FErMTGZQL
EGqJUaFcsQoCNFIEbzQrbNaEEcex8GBZlP9uOJTqCyMwbS+MmqDVKMwB6gCJGeBy
F7ZDObVEfzKgsqfZmpPOe3yQMIa38F+92yh46iP8rQBy82crSPCyJiygEiNsRIgp
G4SWs7WQ2eKzX+I4OshCgcIB0P11KYwyPrhdaT+i76leQCWLWdKLBmvKqcOtXpQW
gweXBDkhSQc8XO/o4oZ3HDmKc14YsWQdbg+obEFHgfMoR6PuULli/vSzd/zMcLFc
TX/dTm9WtiBBl6NJMCXp3IsKlbwKdMWF7pQiJIPtP2rK7zDrQ9xNlsHAV//qpZep
lPUsWSjE8x5NAgTyJT015HoYipbPy759rsJpKfpBjwqwC8wdMDgkRlJS4mdj9gV3
CqX/YMgLwyJjTEud0HuohYq02UbNLTYX9Dco/orTa00jdcsdKbesRTvnC7fHJLn/
dyjlvkTUeCrprJMi8tId7NqUd+tw4LudmrsR+c7j8yDW087jBJ/MsnFCOynEQTsp
Zx9+EiBYTziDpQKP4T2bjmATvhiFZgBDiFA6uVysPZmLBuLO5CtVcqmFdPQWOCaw
HNFx3vA9LK640hjLB0iPedJpQOhdRFV7vsdkIkOTbYP3AQNlpmZkVJ3ZMFBIi4GK
fBvCmaC7/+x6cjRapjQ87OCZi5VD76srQgJjVP8t7b9NNACukZWlAU/LK1ptgUwn
gkPQi6PhSIUl+c9jRxZ4lETRFegoe3WIlLKu+32ZYYeinkd8TFAVRj0zctIJM1Dz
weRiMppRyM7LGw7xewNujCUNbabMiI3mfUYfYtlz7hMlT+hKHU8pJPqqbRwImEXf
NqZTt5rVYAq2n8gax8yEVBo3Kl8fUknoHVcW/JaYriuGQS0b+Z+Bs45sEfRXVnHe
zP9wfZQzLRte4ztfqO1iHNzETQblqr7ZfJUUNmCHZHa3aC8p1BVJUn71cWjI13EC
h2yJy+x6DNxNs9bbLSYDRel5tGp+tAE3USKh5GiJQvmWYQglCyxpDnAO+JdUfTHz
ZsGy9fpbqGdcyi+dpdEJg2p8EIqjAmoz8Dzt1sF8I78+NFlMB8vnoPJDTGD/+eVu
kk50iNWkkZl6hc+S3SrwLs99CZZy1gwvkZslWYAIPGGIoabLB/41Rhz5wX1caOxE
SnTFsfjOpGdSPNXYQChFPfBne4zJRnG8wpc1zhzZw4eUn2YlfKGa6BGhqsQkP/t/
9JBxMbiY9hoz7FTzH2dvKq60BJRqWEKuzzw6PmMTvUI+NskmNb4WtjpUN8E+Mlwl
WcHAlIATZOgiCgwCwkI+E+ah9jP998qYwel9DJtMVP4Q9TCNKrX3V5mqpCgnwr1O
ZPCik16QJeY2BcAIAw0IXGRLCzGYE3hk+sa5Q7KJK9rrvQYlUJkDvWVu4EGQiu3Z
74DyiIutQP1mvxuEgn9UNqd9y8uSrFqhq5ZrnuLd8An3zb3eXVMFyOM5JndOQXc0
P3OoHx+Xss9E3dSnM5m0aUnQlJH1Iqsqoa5Yz5p06S3f/YzwRF2AZOcFspWXf2kK
w1cxXp+R7aLXw4EOLcyzhahQ0+UGWlmQoyGuzZPcYDh/BooVuUAQ5tGDuY0VjHQ0
7Ky+Dm4bydOj76BOsS8hOlEFFqIZHmQp1rFGj/+54MOYGiCmixPJIMbWSqohnGzt
zmZY8RPf5ZFSu+h9aK6q+63ZgpLn+dElWXsgCHmnZQrQSwqZYpVm2MbiE1Vxj6gy
BSmG/SqiKL4IQQVG59eGOHU2FwonlNGs6gMil0V9ue2YRqrH2iVlrAAXm0epNMPi
WKwo55vyDCXpejwvOG/pVtDTyCnGJgIdbBGjj7pMJeR7TaYjWKxqj0sEMSHlhg3o
Ur1XecMwrf1Z+rguoMpa7IXtpOEikelpTlWTx858TaNlLh5u3ZnuYUjepZi5SRsX
zKRCfpSh+Yb4ncPYadOO1eyqj0yMu7tVZMlHR91mnoFB/uQvz0Cu+ftRATCub9sr
0AQf2VLu1YuNbljFpHdy5+aidtY5u7Y5DJPFpL5vUpK1xRLLC2T3jFSWclHE3iin
FsvdTBCPfFkDR2z0BA45zfueJawhxjtWspO0I7TQPZIfpydQVHpRqiXuezl+vrQ0
z00THY+iOS7z1C4U5ZVYJRAOcCAtyGQEAXvmkIdYIO/phLZHTjim9F1jzEcJD2HK
09cQasNU7MqSzaRbJL0NgRrkkTtqf+dlNQ6wVUFFUQCJwJN09JTGu8aRuq/MgU5C
EdS088VJVX/0te+0P6SY++uwHpNZ8PTLGVwpn4e8TVj1P6vuDz1GO1sgserT5DWF
XLlr4CpSHWWYIiTpIN7/0lDdq1pjW1tbT/t9ziQntDM/Auaw2DPGal+K1tghd8O6
uYYYP0ErDaUtToj+nFggukPYe9EhrvSfLQINTO+Wp9WzHckA971ms4oifLfPYX8F
ymjdG3YS+okq/cAzPJ+V9qnwy7L6gcyRvHr1Yajb3UwdLYClD+t5kXpX8eKZxwJm
1u0xrgZDSjVOGTahx6gF9eyUmZCp8J1DDMQs9Bt6XNjGaz+lNkCY1RUe4dAKxyN/
OcOGpGuUYKpHDM+EJJCyTufbMp6sVfOMyRyyedGm6GHhhzzjffgT+w9Zcf9Bzsc/
BTVuVyvPZGGvHRsHlzrpXLH9Oo3ICP7/eADL7NilDOcu/sZ/C+4a/T8UPAAaGEsf
vY9tz2rENxtKpX3u6Qef6m/Ap8tWjm6e3gPEqWDhMaD5DtiSjxWMRiw3UdoFf9jD
sFiJD44EyNzJcF2nwS0ZqJW6IlBq9aa59lajvUFRt1IDumOYz3uu4g1zm8Y+mXxB
PIREjXKbSeHMFr2dSYmuP8eBMHGtdzA2meQsSOpGNO5zPEV/S0mDLvYJmnWcUQjn
u77j6jaBE6yKrqFlrNESiXG14CfGdYmPYUHMMnOyr/1t63kG4LK+HHP/QEdF7EtZ
GlBZdsg72NPBKjbXtanYoKCkMbqOOe0VWD/xWZBu4hgJo/f5tr5O1V9aLH4ZYUuD
wW9+HBJfGQWMzAjgGBoGAXP6mTOu5XrEujji6PNuVhaFRCFqNbt/eUle00FahZ1o
h3q6MSwfHxpBiU7cmwMkH5LdwR4Yyc5tQ+6sTe/3F5kjviO1e3+VYrDJuiKpBwN2
UvkNgV7YQtBDVOh9vH8NVT11zTk4y4+4mnk6WGQEBKWwVy3ii/dn257wJnRMMpb+
KCTCCGYrFgYqcse+qMPJ/uQsrKNHw0fFcUkgjZlqYX/T9OwZrwCXkTF97j+JDSuu
xVnHCdF64vnPGsw4ElgWCjbEB1w4cwy0cIyemyd+I5CFyGMPj2ciwcYdcRz8QZV6
h+aUdGTmRUIyDNkUVsOjKbFnL6NltrvDCZ2btDU46VJd7jh+O0R09ReDWkyZfGkI
g68voO0TLeXUT29+TkMc16OD59f6KPRJxpDf7jbgM6ntg8DEF+bVbJKIWQc5Ep3S
SQ/MqZ+eXgcCdm9nh1a1IYW/vrGToVNQLtaPJh1ECcta97Mqqot17/y51nMQfLpg
PWj5GNRYUbsUy01Mwca68O7f74jlcsvjj7T2sMFV2TG4cvfs7vfxPD6Dv/aDkanz
9K3kPvQ1Wx0CKIaUx4OHd6ydSAXuYxQ9gpFfXNuLJwdLrDSOzQxMPkR3c/fluMXo
q5FO99YW3AE0WzzMQFAm46i4B5Opa3DrKk4TMxLG8fKwcmbpMlGwvZe0061B0kwo
fQOag9lUfMqPiRNUwUS9gMGNNmao3ytONVSjuOR8ZJ0c3wmMfNEDiv5wmndsPpqO
NinsCt3YNVtNa4RJYNV3w0peZxHSFmEhf3AVjsPpnXOJDLCfjoCD2kb2RlMefQpj
3r51hacHYMKNgLd5xsC+Gn/Psb3eZL85QFG5NiY3Uyte+Xryg/pdAOhxIkuZe/gA
KXcouy5Su5KKQDaLgS3gPWoRPAdZEoYEw2VBCjoqZF1VV0usCms2u9ZQOlfzHO7t
wwJTfmwYLnwtqZKA2ewf2EFTy7A2XxFJYtXJ2X9vnjVFJfeXq9lpq9kxTqwcb1H6
r3L343f6m7S0jbwJZRohnjT7syX8aIBWjcJ2mUc0jI6rKDCTm1cOCEZycbdg2vOb
0Zik2Ju0bhUjN7CqEpqzX/DVPpF/yYO914NlEHVhvGnSSZbMXkcsGneBYskGT3qo
xQmT9ADCGpis64a+ikO0RhZRmBI08bku9Ne3+SFszT3UW1x23UOMbyIT0nzzpayy
RLXKEr/E0G4/HHGfxZfJxqZ+ucWh78Qg7/4fIKNLaZ1RTYh6HhkYwDW3+lvSlyUF
YEmolyMFBtP0TPJiToFGcwUtgPCr1B8FO+Caw0kHRMaK5PGSJW/qeDDZcD74rjPH
EZgiZWhcU3Xzh9dkuN4Mf6K4JXBIjHIfO0UCl/jrYgLSQUfs/T8g0zQvEQoNHhfq
b1gI65TX6oHBYLF+IisA8B/7EACDhJ1YNL5ESG7LCxbAb2DIb0MYEpb6bS8uUwbK
3eXOVtmIQwu1skxENj/cpNsCNeEgkrSFjx2RK1uPXJx8nOxBpU047ITVTTOh0sQi
UOdLQDLaGfqZd8Q+7mZLzNyzIn4IFYjGxIxrO72jEHrw7E3Dt8ygGeHeXZFoKOrG
Eq/OqP0Bhroju4/2VZpkIYUNY3zkD4PR8+fnRkeNQoCdOYeBxDVEaPM3MmCYoEqF
ya5LtDfEdSKyAJuEnjAJc+xA3d9x/doGUmlMOzJz2GQoCnJQiH2pMFHJ435tec8A
ir3Fb2SoZZDQdUYNns9CVrrUgmRNvqOTWKz4VL5ryXesTfnQa18KVTJrujp8Cu3z
g7nCgztrtzeg2NGJUwmI8SbIZvwmIIkFX9nfXkplBsnPxHozqgYWHLtPYt+xkXdG
FQZmU6vRUeLR3uFHm8XAJSy5dc4K/NE4iqX05+BwK2yehazRvE0OdSh256/+OQjm
06CYcnPi9vzoIdiBNLjuXuFezbGliu4pCXMWsIfHuEVQOk3qkOt6br+n7eKaJnAp
VU0q4oYgAowN0OVquApNngX9191q8aQ9ODVIHWR9TuZEE19lpq3wNt7bzlQOh4zY
2OEr8SyB23W6pEUDLjYM87sI6X5aD5pJnmlJcfZ0WnJoby5k3eDiQhzrJcj6SkZ3
stpo/Y4Kolgdr1NLwmMK+qL2vPwoCEtqpvGu7Kb1aKfWrfRwMnF52e4zMbkvgZ+b
UjhTjRtyiP4a8iFSZU9AIn+XoEE3mJL+9xG4Iv/0zib3SIkDmltF+zHzRj5wwatU
6blQpgmTwIxLmq7jNK1eYSavQEmYG69MPlqum/xCedoSAJqgsgKEMcmhbTROtM+s
Ou2GM9vIKX+18hkHrL0+4hXsiQ75XMObw7N3aIaerSSZogtcTDtfGvCcg/S+7cyU
VqwWF04+WiidPaiGllN+OvGFnz9W/kfZdHIImDTI8FEfQWJGyuSH64NFx63ChjtG
Oy5jOoqFv0AOG7fZ93VYgw9d+B8tiuooR2SVK5GLgx9j/tYw4hZ/3f1vmfPsj1eN
uRiyjMuIvte76+LQXFx54/s4tBcR44a4CjJbbdJ6fW7ffxAZW8GebXYXJZNxfC+K
631R6BU8hzuoyZIdPuO1QDvLYGOFFhvq3EabTDPqXyYaZT/rxdyvRnHx3Xv4mhCy
MXdJaMhjQ7XiwQB0fKdsXlTgfR6ifWPvpFuy426WVCcSRiJdJVpY4PtB6GS/uxN/
Sjq+B2dvSG9+L9xT4WQprf42FgFSz4POmxAlQL/NETqrpv4zKyapovpnr5/wvTaw
PUmMyq5epG8PtYHW51VwATC/1G9ES0ehc2uc8P8jQWq4Xjvp7eVW+HugIMegHU2j
1lOOcJbWHIc4YjYIE0dU48ld4rIudVcZpOsE0tatm6bq/3sSQHPitqnC03V3o3XI
k3K/XSJklUJVQ6H3tOjqHEyvdeECzUip9/Ii4HnKaAr4RoIsO54XU3LRT2BRwmXy
yL4gmr/QBh8cry67WObYcg0lA/fTO562VKSX6embHIJi+HljkFyJg93l2KRF/hi3
zlJa8DLOfvsQj740v6UoSi9JQF+GCzOegkekWpGuw18nYZHqzZDlwDI5X+OaQKN4
F/60HhMKrYRQD3i1WJ3R15OXlDM2+6jT3ckXpYJbKkwTLsHG+49T4Ea/06ApacrT
AI01bY59vxLSjPYsDE3MW/qpVZRlqU5KVO9njYcsi3643q2nZmG0XUooz81Nh/mB
S6zmJkPDmgIk3ydVxR8mUIg66EQIPvjnr33ZUqG9ATo2X/7rE/TGe+2zIQe0KHs9
okZbchioA4Gn1NAPrKrd028kE4hTjpfYJq2nuHZq9/dUze80JDRiCaJQwkEvJy62
ImI0ET08vnYmqGi/iYy2wApyRJ/kpDpSfPqGd78+s5Khs3NwdthO7ce2lt4Aaq+j
SH6SgUJ0yj11QrS3Obd+TmBJC6rGpu7a6qLMDVB6CxTb3MyrnKpAMTFvHcBwDE+S
J2mk5h6C7r0j+sMe3108SFZ6Cn0N8Q9cEKAwXS0lNXhnuZYnH0qM8udXywr7HdqX
Z+nn7dDwmi7oGFm5yY7qqwrCS8yYJDQ2kOUxsJN3EkD+1A2BWCOZZLmB2Q7XaT5c
Wkzgn9/DUwkNm9ogFkLF00uAtx5hbLeIk+lVO5CvtXGWMhKkknufZQbLJYnhnSTI
2FUQyCCNb+D1pS+KQ62Nm8G+9+qDZFIGAmROnaAH9RWt7DB8E9892kBf/ia18a2m
hPFhmjgjr36zpVWDVBD14hUq4+f7TvXIcGBjUPTS/YJ17ORUnFV4PSeOUR4TVn/i
P+7cG7+aIvo20WJBpLc2PKpx37xanPnnkmXwj1IXLdHb8sZYnvtnVRgldZw05CJH
bBihpduUaiG8HTHCzFLpqnbFZ3z7k6Nz+A2Wp6WatDUKlr5sqLuo0U9Zj9TBYHri
Ty/erJX7F5bHXzOki68h0S+Zl3WToonUBZsViRvJBirlHCfOVpAFSbFK9C5g48G2
7tmbYPfX9mz4MnoLErifkkCqZ2ytVK6bP+gLUCOCDFvSSt8kqnK03OL3Z4F6ePu9
8+mrodw93VpCNQIKkbMZGlTFvfwxDRGLpWeoWoY/AVBtPBhi6fR26uyUWAwOCIfk
PUzkZ/d4dhanr8jHR95oJgmXEwvQXlV5KqHqrrNrn4aqgtNNU+5tJIukT3miBFgC
d/o0yOvG7un+P6vvAEboxL7JWpZfhKcDSKQ3HyamGyrxKooMbFi3+YlpHtQENLmb
ZVRrqk8Jgk5TWvgYaKuANb0f1hIYitdS31hmiVXjeqxKC0lqrSKbEzEK0x1QZzK3
JlsZSGLHzrfwUo5mVaOJ8v42+eIKy+Lj36TgBxEhDooQRGYUL1joenaDPrwMFWnw
q7WO5TGbahvaWRfrJE9sCDO0zziML+3rlkwZy8h53L3d4oDNGrzMIf1gipzkApl/
E5JIREBIP5Ri5QZxftqAa3JdIqJTRlAuI77lPB6eYEWMiSwvargm86hCkCNe3BN3
fIjETpLQ93+Q4F0F4JqyeYUbl5bxYhyKwWiz5W9JebTsu+v3TInH1zcqmE0An7we
0vqD09bALmhJCzLg5/jL+IwALjv4z0qzF5fap2O/ITsi3ICHM9h+dscjiZ7vASNI
TfpYe5qrSFwHQpPyKLFAkgqKB/VhBSgW18sUW2xU+lEdqAa4e4u7ptg+Pat0nRbC
GDFmhfaKE38rfoEsI0MgFadfnxubNa7cCcDboAG7lOwj+Kln9sF5Rkehi1/488RY
PDbaYqvyZfaKXaaMHFxF1pB6NHyIimUO0FC1yGTxvo7v+SHrFYfBLWB0686Z88dE
PHlTIDS/2RM9gdu6RzlhA6ly3mMz1ekdg+ii0b42dznDt4WHL8mDN2m/5i4x6Ybl
4Gm7zZ4InW51+5Lvaf451sHJEIy5qnmsWeS/1S+zP3RNwm8CVSEvUQls9Dn5rl/h
0cXc54sIyFjHd34XtfCUYguE2NaTWHgL3autlbaoQJgM1NCvwiX2ciytKbU0/1j9
HesfHpkScMljT4VGbLysujsSNwV8riLXTGY+lJImcuIalZXN1lCLNCkV8u4kpyjL
yUfjPnh+ivkAZltHkHOgsb4XPiDl0XOEVRb3/1+5l660l0SMpFrrsjXz/BBQbUAf
xk+ykntdeSANNP1zfM6a6ru07xk6juulQr+I+fLRrDyJghNtfxbvtcBQl8TgXqWU
EoVr9cBMK0AZ+/EsCSBKKHTffMBnIRpODNrBSH0gr93Avl9UkIQNGYOLbVFGQZJJ
S60Bhh3LlCLhxarswp1C7saYoS5TWp7msr2TV38RNuOd+0cga3K8TpH4TPCduzDb
rHgGUU+VuBwpQYwmp8RM8OmS+STZR1RLraynl0HrcRydj51QB+d+N4cHBK3o2aXD
V2nk0Uc0Cxn57zo7h88UFCcsXcmf4/u5nTMSNp2Au7QbRYXq+inre/JSImBy/xiQ
mVhIMna+rVcvNtalXO0I5zA/YLwVUfPAh6d97OQVbR1oaxRSvEN5/umU1Xwb+zQd
Gqprl6HKED94HuPY4j4e91nk4fv6Gb+vklfUgH+zAdotBBzD9hoYnx9HhdXUT1uu
7FOMUcK9lpUbyXeFakHRZYIW5JUFP63Aka+U6w5kTwLuipCIhT1FNyUBlX9a2ybn
j+B8xkrFk2tmGzepVWORSrAdgzUXJGbqy0JLZ3VpU61Ka4ivRbvRl38GmgX25321
85Oq6oXP3kM8JLQUIY65KL5p5s98ecJIuuCxDri2+b46/A2L9CWQYG9nrKMAMq2/
uuC+yWpmZm7GFuT7IyUspdg/q3skJBXeg8MUci7QZOworrq4dh+T8mw8I3ku2jmP
eqoSwDv8LFwclB7gU4LT2I4+p7xOQ5FROxt8TzQ5qlmmqBRwXPCOvePCri8Tkf2Q
Qgm2pVf0UqRLwTRM54ExuRr+kEPPJv1QKyfKk9VCMkCUJFaBwQclpxy8JnY7Ltr9
OW59btRKoaFhXumtTsLUduqHUdU3cY6aHPsRp9HWMfRH9zo8asB9MRSJEWsSONW/
Ly5Sx8qn1zcFGFfcLiw5+S6RcLe6sVcOuKAxfb3IJlRBh3qntFTvLR1YZstys2Ih
3WBBcTWTY6fWJRbR/sty6WCsLjoLVYSE5N1BH8AM/2IRw5NmVvEGky/rcoAa3v7S
8koGkV+zNj1c+oljurKptbplj8IvkVKkOv+99mJWRE350rugqq74+Zg1S3bw8yWq
AlnOYfZdFYR1jhdJ0tF5FoTHRflr961AUSpAQIXAau+AT6zEUlFJUGvX4dI+eF5k
qw8BTz0qX6MAxj0x7P29eVIA9nrh+uhCxj0I6qeOcr/DenOkDUkPFx3RAFvbgjiX
rzpwWGIka8N4u9CVzbC5nZM0pslTkt1npUds5kdnjGRhUKQLUP+czmDs6XSJs8bN
+0eluMAdIlUjmBNTfHCzaZomj50+qVI9vAG7qxKwd4lDGrC4kc9IsCB8OBtIA4Pt
8mqRLlPu3D7LIrnISxDMtFgliMEc3I/seV4Nlb7t2q+yHM/xWbITwhFJadfLZz6/
qxsehSi588ap2f7oKBPtgAXp4eehfxXGVrjzttF0iNSZT963L5jl/SR4ifae22V3
dTH1NDTfq0y5jrCcrpOxM/p3ArgGW02Q6j2G11/BQgZ1hOMi6Lv6FjZkNkrbSsOX
wpORTQus9QoGkaO+9Zog49Y1tIz7YkX9WKoxt8RYkDBWzh/ly3/Ulu9VNKAb/u2q
OmFZLfXKHAf7WJhkPbrWMemwMtes93y4dNky5bQG1U4szELlL1Iw0am8E1UH1W7l
sUnS0tnbVScylwTv515chX58M6ZM+7npTwKSaanE3K+i4xSqqUOB2DrsIEHSk0Ja
QQR0r8YeRfXy9nD0E5jtuoflhbdOiVuGCv0hjvIpw3lkajDz+NAERzqjnoqs3zC2
i9uSO6xxIYrMlQw7KqmN2PYcJ4klBkEO1W0FNfSKtOO4eiPAet8u5OjUVp9T/59P
ZBPKaGhPiz3P9zWwCZ2p4pkgd24ST/oqEmjiljzFocOJ1UrOW3j8VBuZ92xHI+gC
KNU5VkCZQoRWQFdLlVFlhzU05g16B/35iUg/HxPUGgzNMtffobmuTkhAH7dcFCGq
+9F5yLUvXv5621ygMM1M7Dqi6wFqNKoYIg8IJS2OQDFSUek/Ea6aNfWT2F7sR7pz
qPB6A26UZEhP0EB8OZY3U0tucZmfEyww3Wn5uuzd5fB2lRdiyLRQbNGsaU8fvV+s
uL3YN3KKGoSzNG6iN3ejht8bNy4DCUnsfHYBgkemO8c9ZeniFybfJQ8kVJjYDYcK
eFqK3/xfMrs+2zU6j0k5bcWzj7xjc/9GL+I9jTSE7zRRkFl5Zh0mM2jKjslyZppn
wgkMfSU4GUcOgkviPASr1ZYq51KnAcHW0/JNYiVakUM55LCCeYNLM5Zb5NKy9iiL
fxoEnlV1iBQMoBjJDw3+7Z3fB5BoUmx+YolVICGzcunz6mogmI1TgplyxTlWJOI+
RAqcmbBqwg4hXXKKELo4dKw1TMhYOINPLJDrl66mOeA32AtsqYbNKRsEKcyjhmY4
6Eh8MBYrcldT0bC4jGOmaCfNd7heClwlp7+YAdZGCg9BQu4ZRlvN7brm6eI3gB5J
QJkr7atmjCtIVgwCT9NYdS40xxd0YZF31NJcJ0wyvza8Nbkuyo7hQBUBgqxd6Tom
96CTCFtfuAJ8e7TrU1TTcl1RxEDOSnO54MfPxiqJwFjCboZUvfZN7E91ZrTH92c6
1VqBDtNh/va3WJhVUPtaeBWrANCieEx8GyXfMrdL0PYxrh2hX5W2X6FWsKcMx1HX
359zIzvqFfLIa+fFkNReQmn0RheDQa8taUm4zYwRs3kRXWEVeIahzt4+UMzRRqPL
+zj0N7TJzYFmDXU0SXRitMKy8JK6ikhhO189jBCE00V5RFZyWRlVt8wusDF7zOpx
OpoxUv/fTKrWS3FkqAv08OJu2BXDjn5exGz1VHjjU7i7Ud/QUpMXcCwdanLIseJj
9ooUdZYxKCCUeS8/u4wgokrAheNKcg4Bd+VBD94FW/beEAnk/m3E4vymIln868/i
stvWvo1gvDlcaDZLloM/O3KODCAdx3CyXxak/8O6jGgisp0a1YzEftJ5aK5otqMT
vE1EGniXfEPvu9psT0uHBvG8ybx+7URmAOp/EFLNYUvRWXlAARO59+SkkTVXcHRw
ak81dCcATzGLYI91Ge+zuSsDsz+bqM7kqYCTF+d+OmJxk7B24i27LqEAK5HMpZ+v
Ki7GnwelXaCQPM5lwuHx+frK/RGnf559D5NQF708vuhlvq3XGQtE9++Zc4psqq5Q
AtGQe+Y8w9WKP7NhJzy1gEKa+gmQnCQyLudunj6UlyIyMycP332EqI1rXrKpIDXR
28qcBaauanS3SnVOmu6oa4iPMSQtIfDzimU0ajdwubnsQcg8z6p/PuT05Uji1JiR
xIT03aofN2JHgRDjUDFqSW35K0NpcaqTNh4sx49O/2lLMwU1sJynQ8ZfO+LwBvxX
uOEVbEVNkmFQsAPySIzQP+jV5uOVNmnw15FceT5wqX6pdHW2XgY8hCXbxny5+gj8
rZglYppXUn6V0Ba/atW7iOqE5OEjuDJGzdlWYNOWBls1axtkFDPKKHHbBiYOdcna
6EhFH28z9t6ekMllQrEFlDCYVEVzZ89F0MPon+rPLSnGGsrKA5c9PH9p8kEou/wk
H+C26EGgAKwutAgrOvkl9Yc7NtvIQ6jsfrsj2apEm1i6XN9fauGsSLvLr+SANW3+
NzKiYGpRR/bGN9G+lOUg2ofzB63UqMg7y2kWrEO9pIz/GR6x7FB563pVzeMIAxZ/
oiX8w0UFCUVYO+J4UKZPKnojQ7gGsXmhmhHLX7zYfK+RqygAtEwI+fXXvIWHHb2p
lrtad8El4MieH7EJRWRUddTQvaAuAG/2G4Nww4cmbQY8TNQ2I1CNMAcPeKqBZ6TZ
mxWb7B/Im2rxIvOcPGAVM/Ehze2HLHBtID8LLKZcBZ3eufqPKqzsbL5zHNT58spP
EuDoRLFd/t0RE0HhJ74DdwZ320ViRe8oNp8DfR4By4q7XrEVfg/Mm3fmVl8HAIiq
Rel5Dwr7vozbdA6ZJi2owb/dofkYHbouBENgFgri0xJnXd44pEwps6yIcFCl3RWS
R9UvFngN+refaXVmTcnwMrFLoACT0fI724OeBo0QYYLSD/ghca2PwJu2gcC1DMFP
24e13ZxdgNHiYCHyZvobArI98s4jf5DNHy1zvMyBD2BfkmiS8LQR1qWgGvvVjuL6
OhTgDt+rkp4t6nd5GNEnZdig1kNRCU5JR3PmetFlzluR3Nrx52HQpfkDs+s2x3Un
4Msax3mcHIxCxi/gFTnDIo7YW6HFFHq0kCJbn+rDi5sPRjTS5Duh2AOE6yHW/hj9
Fw5knJqkmlXyF/9c3EnWOgceLrN05qkycmYxsjufaXIEHFnlA4FA+iNTDYqDwYUL
B5eRfDLMc6YgWRSXXBnZWlH82c1U0itU4oMy5ZzfLdmsvtkRSgeBpnya8BvfmVc6
Kc/7uYErG9+tqKAEPKjAa4IYZmvFpAODf7h6jPhn7MGo4kC0+HJFc+j4EqnNncAj
Ht54KwN0tJVB4pUjxSH+Z6HrPAJr47FJLm8r+TPiUZsHfJBS5XL6ZL8jSzGrXIUy
HGqsvYyxbpdEXXhptrYsnceTjW321J7PLGVj5fikcWd7j2u8InyeA1qmkHE5eP9i
MxjGnp2FF4WofnpaqRC4KSppWRcVINR7vHseuP2WdfVMVwhnRePNhik/T+abIDEK
Ag2pnerQN3Q+zvcszErnZ5+UnSFUARnowJy2mH11zRYckCdOB7J6pjVtI47jDtfd
tEcj3kcNYkrj6zqeEr1ZVWbIO36Rvxt4a5a6wym1yrLzTafzZOjV/cTdTul+tRI4
VAblfjjNk8MAmGrCYojZqnIGFc8y6sGeSD+d2TAqBDvOOviQT7dOm1/nKQtzuLHB
0E9P94mLNUTC/SMLRo+R/aYWc97nGOsIDLq+T/qBawx19q/OhE6ZTe2exIdw3P+y
hVt2eVqFYFARvPJXVzHaRaVZNCOFPYnLMXj9OHXM1sY+pod6bgCMlFLDpjIDtqII
AQ/2DYy4/hNB/49RqnigzmJkv4aC/ZbrCU6BTGcu7nXWWO11drpZszePt2vsBxsb
QyE2A314n9vvel/XP8pVmvPuGnaP8B/UaiHzHwVoj17OkULoiXrofieWNf6z9HaS
721b9wmVr2oXy4E6hXJjN/l7c43ADuRnVuheJ7nXAQdpTR04nmaLK5VsqGqL0DH6
rJzePIhvDDscx70JU9kn+TBB46VGl4KHSNTLb7MrzcdWH3bqneCDmPO/kLhhYZBO
Td4u2XbgIRSJCtSD5dVKHWhcXo1RAwg5YlbayZoAnYMAXKx/gUE630O+S/n9bl5C
UskGVMQPwp2PVnuXacoWRtcaNhH+e526oHtAJYXxVQFfHz4nspt88ioHrxlPYafd
Fs+HZrAcnzQbQRs6670MscICyxwtKbLvzOIINawkNyBaMOiAG3amY5FWvvtvPegO
D5o9J/9RIZCrrIIRPqZ3ngdeuXe/MtxtKb2aQXZEyxx5gbkd9SSUfuYWqbLfLfqc
6unk/lsasLllaY44tlM9JoHwLXyIglYccmkBgBdB+u7X5a3bUQVZ05YwrCgS3W3y
2zYwi9cTVzNgJq7wU9mHZhl7AXywnLVbSrPNDRHyK11zXfIFb63tlXd2Xi+NWJR+
xgUVbLEyujz47GhXrDi3UUY0Zxmff2sxwCUqB1W96MLBHWEB60HuwvXyjDJQSHiV
KBiTBEUjAsLCVRuPulYYmNU/cF+/UXFJMlXBjkblUTxQevdSmEjaPj0JSWeHYQwD
5M8gQg+WEKPJqO/CaovYbRLKIBHoH9FeVRyFMordB4DrX26jf6O2Z1yfOlhgBvO6
7WkraQJIOE8+xIwrLoBicP19AbH2+XT4Gcu+lAcfQizLXGDqEVpnDIYGnEx8gHMx
QnttC39bDnCVX059xBmOx8WoDzW3JRK1Jx67aoJNW2FD6QTMNAuD9ZsHqPqxXFAr
AMCIvY5M4gjoFhVt0MnFH21iFq8T6BzKvmJfCbUwVYUl3EZoo7+8HuaoF94WKC1z
dFN4km1OOH/a4P5VpPJt7HGQQtKZrUl3OgVZpBEaJeaLvBS/+IzG7tXXhoI2BqRM
s6JqBYIDhmBMgQyMT/zDm5HJk+Njql/uLeu1GeInDBqf7Be01voG6KJECTJVLq7G
I2aW2y7F4UMQHH8pLcJO0uad8lgEVlpQUPtnSTYOgRlAVUYhFsrO1PRVp7dA9qLe
2ngTxVS+eGaTP0QuAlIfgcXmv5Kar0nFJ5XSpXQFORAnM4vB7PmogPCRQwcWDDf5
G83HePNDNDQDHfbgX0wiZwyZ1AoBRx3WI32aFOoE94UdUmWhLZOUaqN2wwDTpLW7
2KdH+fPBp6rgoLK9kyFlgAxTiSNoDTk7ExQDRh1Zh4s2NCgYjrzHcmOSpfHgVpYu
IQVe+bip4u+xhxkolED+WZwQ5+aa7X9RzPB3xwmbijawuvH2XUHG9LaUpQCE6U5S
v27Cfb/9wez9OunFZOnjWnxOafy2PhvvZaG+c1yC36C4axfEGDajDw6yuSIgXUCu
yfkXMPocTFePNLkjtr9gAghTh0Zma18qC6At8GBI33eXmUJeuiygb9ZrfqwHnLlz
8ok35oWYZhsRPit1WWNAokuK395oDt29uGmLDJBlXM219U0TrWqsvosTzgPbRtpc
VrPI/rzKhiOwa+hVEdTqOy2Bywgoxw9VkQnfMR08Tie1HPPGVDKlsA/I3bwrEvV4
zYDoTxTr1yW9bp/qonLHs6ZSk2OeN4KD3rh9w6k28ilg/ts/PPsj/7gYibsKBFQU
SyyeEUYxLOxnAhRQyaxQJsyVJ/WtTCmdP88OiRRxMXhJj8ROTt+uUTCoZO/naHra
yiLHhHAVd6uFxaHVkvwrzhLxxFH8aZoU5WnD5ryjvPpAskjjuYO6GJ8TgDEfbrso
fBmtySvP1Ajoc9Qs+Qp6AGxrMX1ISXmdaxT75c4zz18taYqyk+ZQDWiif/eumLlJ
y8xiV0sfyIV+i1Lt3a6eUij9WQQjWIrdK60AKG7NZybyF41YvO8iGMfChQZoa3P5
DSmcJbFKXlNWU2PourkYbfPyibdHTNz94lpC9771kvXPKjlFNNt8Oh8PT5QLZtBz
pjKUb4SChMFWa+XVvUhiEzUmPuvOpjY3hMt5dKmaem8z3+nSOCqXShFyCfKTjj0T
VziOZOPSujZmcDWLfHUMGeR4b3gQvKx74BVvAJyq6w/xIW3K3YPHP1+W6QcKa3Jv
FlTM8jL3/e/YGupMQllyEFjR2kmCbFTnfhSoGonaF2TDKPKDo7f/Xaf5bsOTlVAN
u7FUjdlL64iWTqWlbQtR3NdBTUeFu4t16ey1nPdIsIF1t0GYSi72Z6WHE/Ty963R
+P/fcnPqWdLNOpMaP76Cp3tdmliQQLRxZL2CQZREHlGdkloOvDcghuylbg9X9bcp
IB4YbzMWV1Oya5BNyMby45SQWCEjB+uqm5xeJgPGESHLJFwEeJBdKRM5Q6l3RP6X
57NccJFS0Q9nMZGAzVZgUQTCqGC+SkAG3Bj4eyKN/KboOdVPZyvFIHyVf8YJ7P86
ZABsZ5VUKV/5IM2SLY2RqjKKwQhLPPHJQTpMl2sSfVioBgXam4vk3I2bbi2te0bK
pSj9RbdXc7gKKZcSykqRAdNCYGNWtmSdFaA5TaO9WxjH7p3kOUW8ian0TAx3OHnW
x8eG8719t3KawDHFTLzwkyABT9eyka02EkvbZ5WPZg/Ia0x4Rfkmndly1nnwTmub
OyPlpjTjb876c9QyAiM/vo9dHNCae1USuubIoBGpKt3if62bYV/r78EGpDU91yIS
2gpmwUZFAccIDyovyrnQuT9kIkgpfyLuJbBOMbwiMQUmWJ+6rdi2WpJoT7CQN2xH
P0TIux23FlYQR4xqDgCV0JSWVZ9Ibq5xLMwJYYM1OxbtDyFvK1cK/CHAmiRCp27z
KaqeO4dOS9gfvKaO3ySDTcCspnXajQb3ePst9YP41l8pXPsY56mz2xlgwdBqGXwm
JwyXUsvw5siNQ7I7QVnmsMZtdmTUODtSzjepczwNFz+2pZbA/cFLkCVONLxxewqc
bKEt5hKIWHGFZRroa27Fk4Ieobpiof7SrRAgO5904m9BUiYSMqOZkcJWjzn1tzM4
rFFSYAifoTcSFY6N78eicUc1Z5N1X+t6t62puq+8V+xm5ZSGLcCscKVt/u2yxaxZ
v/goI9oKxaEF28l0KsIofBdjXOO9D+Vw2WAsHyise+rFJ0/CXcI41susOxJLN+EX
lqYRCfai7hBNSRMqeLZBv4gSbaA63s23fWhk3iI05BA0jx92VNjSZKgO66h4rgNo
RqmqiZiHoM+t1kjOmJZb7+/L57VSN65NeLckzugDPLvP/ZAchGzL6YMYmIlMtR27
v0yDKvu9YZpapzWFrHeigWLnjE6ZjCFbjsKYECwDotCJIskWSE6GfUPS2ER224MB
ILMZ28Ybhu+Xoa12epAnmfY5+hXsSCUN/2TghK+nEHWBXcunK0Av360peGXGRcwp
v5/dqRPqK8w+8z6R8Hkx23bHSA6n1feW4xGnnSDtE/9waEVB340piUpcIEr+3uSo
oy0wz8caxRjqF+G+TXOJOWxwEwNEi6Lah+JRZTd2ncUYNwch7sFbF3+x5GVhyD/x
jcneneEkYEq6Utk1i6CKQX8WncBbLnhHC4rtyYmibSeNCkqwe7008/LP3/BKHs5n
eDFzdZtdDSB5bd9SP4nQqc6GuJDPs2198W5InufzfOYLsXw7nDp1P8/pZVYjbu7B
6FhW9bfTtMZW1S1+/wKPwGXXzQCwdSbyIqpDJlCCq8dPk4TAkRGftKOLxFiZErSv
oqeRYTr4ljUCSGIeiheCT/Bn6pnwa6J1UJ6zEUpJYdQjHBi8R6gvKvKwBXvs6y/T
Cbzzv40/rpQZIuKLxNI6hH4nMtjtU0hFTR8LhUfMNivNAW8zQymQj5O57Nx0eU3G
JRoRbT28RFk4iRRGNrENVSWySalmVgq+tOgww/8MAzgD+VGgGzQmqlWyn+MUC2RA
5eISF4ZC8sqtTr9S30PVNY0e35eoLFU15YxNE44hZY51nHX20EXYmxvSqzlMCgq1
wXRGcxsmTo9e2mT/HARpSao0pX2Gh3j3HYhPY9wR+eeNY82CZ7KH9V+61I0CxuL9
A1k+TYPZoJods8dtpMJE6a+IVRK3fCs7q1V+mjtrLzubHWyY1EPhRVeRxIeOkPs5
MKueIGnxwAVnw6LYeLn8KiTa0BQx7H1vSGuCf0Qe0M1014roeazNOubLiARWUTJ+
EvX4dZFWh7z0dV5tZHJ+UHEFmPNZm0dVx6RUxW/ZoxjJHt+6sJog98C+w4WPapfo
b0IZKJW6bO1I2py2hwG9X9WZS0T6AQk3UBP09O3JBUsSeSTEKfelLDhIWSRheBgr
cVOZmSZphbLdZjj+MDrM5qd8RA4urizuVDlImRHFPXJT7WtfTeAjYimvtuvJvswy
IYVDUikKCNHcWgCQz191EMG0u/5r1+mvVtlVxGP1D8WMz9I7ci4aLOgzjGPgA0h8
EiUm9lYnP41rWxOfgesnmbl8XknmP+ja6qYnBhpR2V3gemSL+5HMzW7SeZ4kBbbS
G//WsdvoFaHc0DtGI12XRv+dq1dFq23HgSvuBtl/uxIP8nEVvs0w626escdmsmLf
3LMer6zPeYYiJvq9/IjGCWmF4iilZFQRGZm85V/qo9PCEwJqYJzgr88+X3nrI9mE
bbcmCSjFYR+gGDJqZIPROS8YpEZFFGArzH1L7cyvmrCFMn6Ccv92yL78RNIUAJOu
0z17wMsBrvHC1udkY+WiUN2qcktq0w8aA6EbEjP7WJIi/Rq2TBtchdLn5NNjUQNe
M5oOiYb7wRW4jAoS8aGHuiQauCIJrYIWi6/7gaP7oK9g5ibjXPe6+aq3TPHANGJc
H5nvUCbQwIWVGOO+QiB9WnIsxyj1Xz2xf2eEf+c2NjybM5cS8zDQx5kcm63sDc8k
ES5LHdeHxQ8Is7Vyd7ohrweYnJq7bBGua5+TzGMrIvtSITD0h15ypVsbvLF9Ubef
su4P3X5pElEMD91dzPFZiv3LGrqIMLV98FfL4q4j4lEroG+dxf2XyJNMrLsUlsns
bOoG2CMW9fkkib0nvW2TftUEvV1B0+46IaiTpIBAg1PRT12FazU5h0acTCyr+4rd
8cGTzn+obnFmU1E9VAS/3zUPaU2FMY7G5hOMgVuNtUeelHIN8z7n2Zian5zxvtIu
M06x3lUO7NEL/LSKitNk/L3GoQeJHuSYqF3UJAVLrjUAtYDuf8uIkHqc3LAQzt/Z
gMOni56zr6HXbqsJHtMEaQgrXoKX7cltTxDJydhtMCXmipbE1wIJINZJL+cU0XqG
rjUcMj3rGQMezriFqCvbpqdSm3VvHBRILhoc9Hk0tp2EJUZI+Man3ebc+IhWuGiS
6wmvcFJrlk8Y/MAfmDR2D8KfA0a8HlwkwuG9/8REH2jPM2V6zZwS2T/17QPm2BAT
YSX415dJ3a47sXFJZwyk4tGD8w1kCZ6V4WS8WuNxDP6Ge5z5heUkXlUe7i+9LzkV
0xp8JGcjbsEQtghJEMRwa2LUUgMK1r6/RTCMOKYR/Je38IphH53ouh7b8wHnsfGW
7AODXK9Fy+R8zhJF7BKaZSrCYoMP/l7checM+TXerspFvR8H0BLWR8IprkK37taB
gXwXkT+aLxmxMqKykfJZOGb/vcoyGfljuu2CLgBa/GFY+qtRsOGYdHtYoSBoDOGL
D8FtoMKCDF+ENY4AnfDE/5m2wtCoysHzQgI2QIOMm/FLCWSVnxyed0vMIrQMKpv7
wmwb8SWjP1kxi0EriL53WkTiyjEEnfCzEXbLCfTifdcIiib0MhimpzHC/3z2Jf2a
7ngrgnllqvBbPZoWp5yl6OziyuaKjcFBD2acrNnfddHM52VS0LKV8Hr0Fn1di/EW
pnMNK56B1nEmkd7YOxOK0ljum1VJwk3N4Ao+q2CCaYYlC4eQ8z5yxPe21+sOSazz
TOuGw7n0uR3+b+vLRKjtCEKpTiAiyp33LaNfkuWykOEsoKynehDpoVQsysu4eWKw
uqshpXa+ysdQ+4+mByr1+T7qPpo2R6Xi9TFRchpY3h0gQh836a1WjzBzTqWu2kg/
JitHTqC6p8/ZAzgYKOPMlBuCg9dkGvUY1PntI2mXuCvQJsHhmq4pbTt+7I1FZ0du
gcS1fQ/GlbJCGnEdqZ63k3pMyaSNFiSSNC47SjsoAmdy1DI8V5R2WfaLZksJk8gE
0ntHvaFeIDyO3mgDxz6xHWvn/c/u6Ns87lSRKBgZfRJFPLkQelXFhwAfOUTnKsLT
o6qHklFAouU1qw4daCpYzadGTStAjcBpnB6KVbhnx4//Obr1dTaEMZCn0hSyKKy+
KNbbRYLZYLs6UUktJjWN+xk/npM0rjV/MA555WAKkkYXVDkNnmFbPdyRwNq3MFuc
vb2KN1jC+yxVZAk6ul9hD6vB4E8h9/Wh7r/LUN0WkdSxiZqIzwAXl2seZz4mSUIl
qmOEcKQqu0QcBff1jZ1ZwjPGko5AdeEUWKJtJR+wLCmwDVvMlx7WYFPX68sUF5Dw
qrPt0h5iYuSAny5QrqQEYce0iD35ILXlyQJT2PsqXChtJhYXDkUk2i3TJmhi9ixT
7n+oR7khWmIGXgD4YCfSKmbSnNt+nDHSSC6Gss2Wa3amtAG4doQ76Y2Ieb28FxCs
Awn4jG8OsHBrilpt4VSUXvqpZv+cZuv7c9CfnUUznKJTHeGeolUq1SwX4NXioq7K
ovkxyf+3Op8Q+qLT6Y8YGsuQHa6rXK561zzAyBbxcm108cihOYuMrQQE7sg7xFIx
FrymXEH4WPKpL/MksTCtjsIl72oK/m63b9qFgN9uEFU9wgDzpSs3UFH8k00QO7xd
a7ylpz09DJpkI/0PI52QOBkNY1nnUefznJ7c54uPkE2biSt5Bjb1eSeGbVAJ9YDM
YX3D8+JAbLigYE7JxCsO1cP7TDO0wUaXcnmwCbR+EBiHXLJ2gpwd5gk8Aot0EloI
Mf63zUDbuGfCHPYopZxI4CF3jCN5Dgsg+qYY0p3hLY5I7SNokrQZZX7K2TN+I036
NfzUWFYEhlB279ICK9szJHWuvwD7om6Xf+7+1EN1CUP/G3mPvb8nBC17FT+IP8s3
fWaoK75uHrS/vHTg6qtFgl/Cs2z0vZSy66Ic2g+Wv3UEu5ISMbks4qUsbGZeNWvr
WOtbApWWTRFr1MBa4PGAr9j6GfaeL3BwEhyTf/OPDf8WVJMx3dL+2ItbANzgLyek
GvM+sItdrJPIFFkZ8zYquagsDjU77djnO9D0wffcBpZPsZM+JPryIn9DHmsBL7XX
3aXhIcXD71XmIF4IGTJpuk8y+Y/v0DhAXPSBS20s+Iy74wRnKrhhzq2GlzvkiEEg
ZfxyuGCJUr6xh899tU6kO3GPnPVFYqKBIoSi2+T1quPARG8x7dEZKtQ7517zjfeR
9ATp+1aPrvK9Sor9hhKih19EXzj50wQsxAIH9sJOBo9fvVlhfg7EB97YdpwTqUlO
rWdGsLqD6rJud4cD71renfGyF/3csS4WRp40EzB8JB7lisC3DbtH2M2XqABwdGEs
fIgtpQxZWYnKQDfYl95EWdQGZ2eHBeP9Luhy7em91FKmeAJpIWuYBAU3jpoGxWHG
6s8k9P7MF5cp4sOtxLl+/QZ808IJ9+8AOIY3hGAYJKsJTwc2r5GKr98qzbr/MRWG
FJfF5oGaphrcGDVndVNLjtgw7F0IQiVCZa135MLG1Sh/lJF/IMqi+TCmq4BeoOHS
yXwLD5ZDZee70nXA2QZcDwEm0RPbLcTxbiiMUmFg6BkniB09Wzq9iSW4JNt7cu+i
qn/z4zLDy8qCy1BWCK29nJ1eYpXMYD7/jSIzfGu0awPSQ6T0ZCvDS+nVZoOvzt6J
zFzfFOjesF9IJ0KeAf11LTRD9LUe7Kc5jWUy9C/SoORIdw/qHbU3cvdBSMvIdFOg
k2lXEeT6LDfoF8Yl+Y1HDdNlnZCg6nkdumOk2YxXrCxv+IFTeHP9YIoZJU+cUhkT
XbxS4pbpoTig82Rv369PLkSYYydoz0WmeFwug++td+6bkySO9i4/eEeVfzK9L81x
zdAo9+W2AoZX7ttYtCo2WrPB2dYng7ByQETlvImFNiybRW9Z1px8x/kwQ2T2weQF
j+4iqJMJ8sLK70HBs+1l7uQpMs3vumMU0ZhA0LOy5Sws1OcntlC6xOX4pThc3f+i
TywhBaHi4qouj1xl9dnM9Xw3UzxLWJ5us02lTe+QgBQO+5KoJ7R/gjdeep0gVDeQ
UOHnqttvxMONBhLTIvS70rDXWPQsvT2lU46OkvYouIhx8K5zi5F71MId3WJ2rj/4
pL2uPlHtnwYSLqHy9Bj5AwcUIAHtxzqjh8ZyHMXmhC/rN2nO/DimVNM+HpJgwBPA
Lyf90pKIg/SMu//dzrShoP0v6AGaXJhXBry5YUrLrtjAZdJBdVVNTYR3ikGlJP//
LPFpXKtMFzJzBGfczj+QzrNDjKsSpGsReZ4Uf8cF/wRISZr1CkqKhdqo8d/QibVj
09CKUub8MXD3GlvycmViLQdY71mhBqW7WdGu7DpueKP3ZvA0Ui0dHmVOkB2aeeyV
xtOWPpTbc3VOFpdO3whQzZIaLQERXc4T9lwH5M3Wq+rgz3OiqLhBahhubzWCo023
A3HXChx9yDiir7U4SdexVeBfudxVSc20JwkKW3oVHItahFbBHq7rGa3jFx+4kHce
rPSWxtEh2fpe1xq7yJVNcFObmzpTDNfsD1+5z8c8otcFZxkmsDT3JbqRs5REMQBg
mbXD5LPoVxo5sGLs3DOYxlt1cSxBVeY5ahalDCVT0Z6gbLhZKbO9oman5iE+VAkW
Y9ErcO89QzQ3r7+/AV7VG9VfFqrf5CS2WGP2YoE+Q6d4dGxOUX+ZG5rl754Jbewn
h/EdhB2VGab6dJiq4mk2U/DzNE1UXG2TX3EFM304uQGoYypuoaG5RhROGYynnSyw
+r879pIlrQ+Ldni4NvbGcQUx/Ija7rbVapNBqxZtwZC+DdH6zrSKzFTnfpt5NS65
RLwZ01pyGynL3o88yAKo5Ui6E1IFSVn9ugWFFuGqApDA0UUIi+ia8QTUjB4FYdKY
RVbHPhKbavFxbiT98GgB4kfjrkr0mwQqrnxtlSOYhp9QI40ddoQ+w6B6BNQOZUFD
JT+82kEz/WSPeuuTdqHPBgKXYkZTiB10nrKNbo5SfCZihqK0mBlSKlNns1m1T5XC
C0Wuo56/j7o2UGQv6DLI4J0OLcleIccJQyAU0CmPp6cs6E2W4VKxasUvUy3qmXv0
gdpQivOFpxyA/UZBUqSx/oit+5q0J1cT+wzlMeOajDPlT7KovRO0FVrZ9ItOJ15F
xfTvGw6zthCdNeSgHDHivwW/D+OtG7IaIfxuwLOsGvTouYnbMfVfwlxAgvSw2nyc
rCrYhxaPFASYpH40VZfuYjbk9YAGFwTaqMbRW1eV1JAx4zQHJPRzAzWqi5wlK684
8M3+oUdZ0CM2+5i4a8tJILit0lc2z3s5EyToVaWTglS71Zc5cy/J0DTIbSEICro6
qBtJRdS5NGI7LiqzRbpNsZVL9kYshTtbmfRXxCsfg2sATbTjbanC5D6X10yNRdCo
qhD5GjURxo9ZlGZTzRLoqD9wPQ2XmSfiRcwwXZDfQfLf/EJgIZXsST1CNz0Q20oK
paNIbmJag1IURNTFjbg3leoKKi0DoW7gCcHllMQr6hr5uUFZihI7kBsMc4cf/XUT
JG7FzD0U+weqnbNaKcjPaox9wdxwpo/C12tMAN4dYls2DPTxzTCB5kJaZ2yZmSqu
cyGgur0C2xBsDNmGHJx/hboL55oLUclR+qZ+ykMrFaH1dkcs2vJrDXtJcbzY9gpi
dMpowp+PGcNI7vnUr+4ecXzHkcQqCV+WJK9Mt3QmQ8XWZM7gVsFXXcBivUpyxNM3
g6RjzkjxC9aAjUZczZBp5eQTAhdWo5kzsd2w7WZ+VgANgq8comOJENF3K07aiXxX
YH6gzsMAi4QA0iQSyBNocyoufG8vyKXbRzTqhpTBzQ4vyc1SYB+5sSFkbjZMkRPj
3wbx0YawDq5cIdYI25WY0LllwP9n3H45hQuPDBKUJWOinph6MVq+QeChnZDzIXiP
EeEfg8KgNpYX4F9WPC9FNaoXqGmdWEeGyxdlet6OT5hdLkXi5RlSBj7D+Q6dJNdE
OyjwH8eacZYCL9qWKGQeapw/KykAziSbDvrESp9VRU3EIZqeeGJ14KwDQ72S0CF1
4QPO6E7+ikKvBV6kMQ/xFwOxeNZ/XyvXK4wUQymK5P2bpNOZPgBC0EooWENsDfdb
2V7B3F1zhnp4eed+U9AeY2ofLcP+j4QHRbtr8SnQzhigDTnzvaWkxeoo9HV87qYd
CMk2J88uMS+5xRFhTHkUuqjPrkLANE/OUdOcSTHAMfNwWzt4lqpLsTmUY03lAs1I
ubCYp/qoMsgP0PWgaSD5g/PdoOIznmlLrSI8usy2HIkz14gjX8d3Oh54lKNcITAE
7dsA3w+JF4A8V20CzgKr0axoUVNCij2k/TI0rE+VF7UBAIdvA4HUOLgFuN/vMS+N
G/TvxLRyWB9mgdbXaCnp9Rvr8uki6AnWeuTa2NSEwpsavJzrQXDgR4KoPqkolPIC
FP8qBJMYA1CaFgM6DY4aSjuYxYv2CqXcTj4LlKw0rDUZFyNZ3IgJ/O26vn9cYaV1
zGQuiXjmc6rAIHpy+cHYChfsqZ2MK8yPsyoO8hl4sIOo1skinER7gD/cFwOtjO3Q
M2K74i4vp7ecBaiT5eML27940sdNdZDUPxf6zN46fQLCFA6lNQ42UKGiu/+IOFol
x/KDlPNUQew+PhYpLKqCXjHXIJVa0fK/MT2QDSvKHO8xgZywBtxYaXtIAeNhph7B
lK0jDrF1FoZT4/b3fQG4IrDs64e1SlKsw8+CJAObgi2XBg1vsZFTapSdXM9O0JT5
RGVCpNWMqwVUJCxrb9bQ3J96SSQpjpbcUvWj3alIwqsrNyGy31qKPTrP1e4cdCUl
LsMLt6WrpzXQPus3QSUmImxVFSH+2pnAq95bao0ofMGILOtyuyrg8Rw7QM6RH5KB
IrO2c9jnbXB9S5DVM6Edgv4OjT17frzDoEmps6dGnMiqhXCDKJv08g/heoNGlK3m
/QOdcJtJVrBh+U179rHXiaOkPfTv1VsYiGq4eFPc5Tv4QvZm1Kuc9D2j0GXI3b6z
P8fRnuYLOtqsBGlO6+lMQBeMnDzw9z8BN/ty1217Jqowgszp0m5+mGZ5Mi0iFSOD
t8kwyJNdjIs6go+Iq6wp6BPNuAGNkYXDaxSpb56IkabxHXHMjzsv7nLUuLxYDvlz
V3J5NlCgfZA8l1gx3SlnOfPfyu4S3YETpmzJ30YvFudY/EO+OOVipdIR3aLlNKpy
LM1g5apmeGu071CMS/g2hv5OUSasIzGqo7uuFm0F1cIUynkTkPbRl6wN0MxmwyNt
DJDTq+HZXaUENv6IgZDDDvDk/WxzC452HMuQE/gdePDUeczFg6/i3KpinLG4oJqF
4Lb6HW/nZaVUDSTV9PAM3gnVQ5zKLKIOImZViyiKH35hG65zclx8pPilWHw20B0T
nxfFawFPqYN539xJ10JkVh+IDz7sW2ESWCSykJWRoxqO8sxKTvNr+pte7++gzw4l
NOEdb2r5nCBMtr91DuV0ShY81zajjI4YdKgJThac/XYLJg9uNHIqkrw8hQ+eQcBR
QJPS18G3eKQAIfk1dUtm2FhijOYkcAntN88xSkL4Hm0aaJFhlzC/Vif7NZKG2oWE
a35RRcszcc82dl9YcjhhvmlvhBmmItJhKIvrIElrV/mACsK6vdwZlkVoy+39F/Sv
rjAhh0K/4hJTKRsWukkExI+4+x6B1u4KCjW3PGQhdo8bX9SHwMy92q6zE4OdXtQE
cu73avpJVmcoND7TLrjpjvA7V5Bw1ogay//mtv86b0yI7kX8msUuQSAx3lU6oore
gZNXNYA0gseSLr6OhRUYA6Hy8Hp8cEPKE3rMUZcE+4SwNidLaodyCHdlTUYFjA+t
7fZsLoAZYIkJqjdk795SYA+VPi2QOoiLjwADp8OuGTMWNvlNRykSZc6/GXnMOOzH
UO6/vMqcMK4Ow4N493SwSpnIgwfIlu1/Yb6WQG3QoHDBz7FdgwDEANBGkTox+9Bl
odJeId7kxTvwTP7tt1wcdCccJwtxaBcp5Bi7y7QW0PdvmaU5I15Vd8CljfqbdE+b
qGsLFzkBuz3ls3hMKSOYqgINwfBs0yAcFao602fcqjAK4Y6/mBXtmxyo0LU4EGlo
PUUWvQMW2SxmmuhdAAKtt19ukUQ0djzIto9B66SItxEKuveS5uFh6b+fPoIB79IZ
V5XcAkIU1nwQ0VhS1hjMSWlQK9o1RVxaGMT1qXOoZWgrD8gf3QipgWSLnp/WHbo8
hIZJZ91y+yBe7J6VI0AL1vaxbVR3RN0YublcnfpNAS7vAnlcYyh2n31ARThIDclQ
NDMol6t5v87U85dU3AiSkfU7dS6pU1mDg7roY7mS00O7KebvAKCTn1u+GHdfgbFT
F9Ea39VhzcdMQQ3O+FhoQOfQgDmmf+EfEHpwbwP7TmAuIAMBfcnHwnA1k2Y33lQU
+p9+qoDyKrPGDp6RCkVRnuqrRqwKcjVSaLzeF/qZ4oyW6wpiQPazw9Mr3pgEd/lu
fe1r9EpWwft3hv+QfctfrlYuuxod4LMVDSxZbCSAkAj68YYVUTEmbZGZayRmmK7U
tzuSgHVEkvHWhwVGtx1WJZ8EBpyTy69XYyuR/Y2Kp3T+cweDT5iSDgmcxbvrcRLk
iJ1qJuOz2OW/x5I1wdwc6MOdw8EjjpP5xB3uXXPfER953bY8gWqBIQwt0EbK13Nf
lGbeRK9plt+eZq9aUawJ8DZXMbjZbo4jGgbrTKE0y3ofMu3rS+OZ9lPCZIt9pLpd
nBwUEB65x8PZbHrMbftoMG8joMWkeq0g2ONVq8yyK9XzYK0HjfENb32E4WWOz2zs
jepdcEN+yPzv9MZNtnVjsYDwi6IVLgN1mydLroZuWSyW+9Cw7E4kD7LBnM6NIPPD
Ev6KCb+g62a8IBxvOk9RwPPz3Tq/Ya4s/Ux0VqjaFwpKQFXvKEFm2+ng4ooz5x1w
R+XtQ5wAFYdkq6aa9aWFXEvQl7Qs+kABp7TxtWy6pdzX9t85EzsZe/eJtqSU0wLJ
AuGnppMdRT7N9hGQU4PejTdcLwMWYIKrxF80IAErk28aKSOtFgTTjYCn/Q369SoX
ZFP6/BIfxfgpYvFfmsPIiZORYZrKsfs7WdwV4N1Qejy7mEMJpYTfwuKl5/wnGMZi
oazHz9vAuEh/8yO4TFZ8/NV1zpAVBTfsfI4LgOtkdMU7IPxZqF6+uJMWB5Rt1FC+
yDTM47LwCJ5rlULNj/Mi2g4hQVL+SkkQfGpjfTI0BknF9iZlYQxS82QfpXiu72gD
pPJ7LSlV6NlfiAqmF75SRfIM0sg7Rn2nXXK1JqxV3H2qlFCyaVm/tsXLFvmJb2Dj
o8wmiUlEwaaLVqU7TJKgWmH9dn/luG+zD/PHR6DpGVPIA148PZlJTZT0BVAfCQcs
LiCOLux62955Z/CPTTUlznFbZMnwcRVSbYHRZ9wgs93g6+5botmZ3FzbJ6X73FbK
A+mW0bltyi4jDYTDHe2/Wq3oyu1de1yVjsrNtXnjUeIPEaKqyV3rA7wTtYn8YpNX
hqRcc0bUEBFrj7QIG/DIIfJFLFWnHvESG/29fzP3pcO1W3TvA2hUdqJtyWHQwbTI
GofWxz4v1TqslSKP10G6Q/E6+eMiY9VkvdifxthxdnJVtCyv4YYSgClDBHlJNWZZ
dNFDRsZ4JGWvb4Xj8N6uz2A+waJBkRimceN4A8GvLm9wkpnPJd+Y9wcaCZmwaj7A
N6tB8lE7imvgXGxiYAK8yBnHUbw03c+hq2fzpW+oa27ExgraQusGRtAqdF24+Slx
e+P02U4RnkKuZZZ298AiJngjvWVU/0HoF4UCWTWCRQKpP+oli5+SgAAD84Hj6vPL
FtoLVBrUDbXLoWcE6wBW6zVSngcdt2pLWz5BdJmPRrBWwBNzBE5acYc8QgY6zCAu
v2MoSJeOEDJZCzhep3zA/2pP3hNHMk1sUsqlwXD0cLZ0h4b3N/3+B4OjJkpBddDk
39jiR+QaGh3wYFIE2+jyhXquOR4g4UNw7NfhrxQzKbN5fbAiD2xbt7Gyobety+w9
tGZvHhbGKe5Ja/HEeCerR1PoidGLeVS1oZXERp5PRZpMmCtVBeV+vAQCnISnlCC+
tPTvvHdj5PqmaHkgjNUTF9yO75FJnePRr6mAPuxsw/ohOnXHSuvHAhMacp5lVEHC
Bh+nfCJ20utHuAtDTGzISY2Hecpv+3yA/ZfX2XsS11qILe+424QFuE8X6TUJgHN0
LcPAwdgY7Lox1gLyhmu9U072ABNU2DNr+RWmPGPDmm1FzqkVRf4n0ds1Urahd+BV
CE4pMLpiGJgDqZkYhMhEd4pHXBaSi7GKkU7F/H86kkSLxvz5jCrJ++9wZ/ec/a0o
c7pHHlNebwbRELUFwC6MrnH9hK5XzuOksj2HSt4T21npoFoa3FZykAbY7y81jYJo
eck3Y//kH7MIYKMcHtyqeQXMPVkINqHH1erEva4e7yMxcRu4uLCKPvEXqGkUiB98
i4+k1rDCRldDuI0MRPupP8FZfUnapMKmPxbhbS09SzEXAoAAc95uFN8mM03B0l0U
zqZo6/ZvtXqect6bDGWSnEPXIvBeQAr538IzJHa0FXnkz7uGEicqfZy+5mzfX4zm
7b5GQzu4M82TrIpDu/nlq5dTAJH6ZIVugtQviv0LTAGoGODelcCNJkjxynvYArP5
e82SJa0ZZvk8BWDSnMTNvdApeTmSLbfMl5m3SwhLg3MwCnqUPy3vXEA2+iDwdLhO
yfCc3PvoabBCVKBHeWP0quh7cGcqyi+ixZHyf8lpYj6jkcPk7eMtrOhZ1VKiVpBQ
JHv3UuXaDVLXGx4kOs9SMDbYzmZl6X7dHrHnAazaH8ENaTS7jBuSeja9KcmEFf8m
qrvcEjA0rXg8X82Hh5CPHZT91tEeQjwUuF0hvLNfWGzDHGLttE5k7UP70RUW8YfC
VbG/Kh9KyQ3v2njPmDIx2ByI9u+8NeIfpY/wimRBsxf6CeYSb+AOOzYBJ6noh+zy
VKFQVDYScIKg+2rBFebl35hvY22I3EA1GvHvZ7iciGvB9+J5hdH1Z0aUsarHkgOV
ckur2IFMF04TnNT+yZzin7Aj0uXK4rNYvCVN6ybMX2jFo1pM5bztgmUaV7Z0DCIw
KwGBqsERhPBCCIXNEPyJufCTPGYHIdT8iYsjN3U5dySJUqgJP2HRP2jDffljnqPG
TJIRfIIm6DE4a8vnnYgfIFubWv7K2FuYXG+uT3j+nvmT6pr7e73PmuS+dUdWvyxQ
a3nRHr6sZTsQJ9xdK+FlGzqqmipOzUk+gQCE2iUv6eVXratNaemRqViWbq9Hmymn
nqEGQr5f+QPkGD0scLwJUQLAG81iCTUTo22O7mMyul37y8EQnWrV39nLqwLZGhO0
pPu6vAyZu7mW+zHgzwcKPiHDxkj91QVZmlhN2DArrDm5UkXz322mDWgV44MOUmhC
p8AMP6AaK73TEw5g5YdfJkzOoE5lwqffpc7T04NGggY0wMGgygliO6lKHsPOoj+K
KdBgX/HoWDM/p7h/W5C4YoIZhxC5ti8AbBxcH9Eup14dmSYVzsldE8sifwBXuzTG
wkItz7Ve7cWM6FMTylqhNdrY5YKQoL0dg1uWMyYS28b3SFgjMI+9V9HL1vrKXqi4
DW1oYTVEbw/r9UhR5TNH1zgDxIpyW2pIFzHRoOQgWfuXvIMN7JP2p57Dd7hmJG2j
nzbEN99Lw6IhapV2TsAaxVW9MhmRoxSS75ZKogwzvF6R2HwQM1b7wNm6VpNc2gct
Mez4ZWiBVFudtH1sLVxeyO3ec9v58h+U/qEuI+Ilr+9xMxOwWAxjfpFVf4UdZI/W
JIgKsOQaak1gB1HH6THhKzveXCjl9qnvhGoQ9yxtDN1fnuYm588xNc6q9uTXpzvl
eSG1o1iGiZumbcqLjRA3D6JaAdiVgiLVv8ary/ln0XfYt33415LneYMUTrdynXuJ
IHdXdNuVQk3vfE78gRNfOfLCsvtQQlpyjss5iQiCUIeRcqeqewqQ1AJVX9wQPiEq
wV9Q77x+RmE7TYoXb4gFcpEbQx3R3d1k7UQxZVEEzbHczrnJPlklNBU/K/4gck9p
B7Dz0Z+XEw/TcH1Kj56RLlnZQVhcDTg4TfLCJ0CD20HyyvbixMjuldxOPR3fgyoQ
+V1xSvJ/IQw83AJV6/2I0fRyscBBSNm7eY+mwPsxyyzOFKpDHpeayjUAquMf1smO
CVgz0ulsXORj7PDRnYqux+stb4gw22oDsfyzaO+dSE6XYHs2EcOTSBq6QnuF6pRw
VBtUQEZhJ1tj5X6XHoks5eFqnderQBKR8HoS6eY58Z4nmXFGc7cEvY6KbgbDCU/D
y7R73vmBYMGO7dX4x9J+BufNKP2yzrzaE+bz0aPpiHXxRIc/0geRGMn+zz5gemT9
SaJsUY21Wb9fS4Kp7uX+qRZhM2y2DxA+jQIrJGHcLHg/jDDGt/fhYKBbJJB+SpBL
66P1tOpC2dHGjFauwqs8HquuTDARRVfmc3i35ZFtg31jQ1MfK/78amqrxA5lfcIX
YGGQjEkgvsv9t7MVnhAE/Zd17Sj9OCWbhy+1oGOc1xn8j8zg75ZveBtj4c9iZWbP
sSfyXBzYUJ49BkAdfkrbtsKKfQpFpbLWeSM7zTLW9hTEh6WjJD8HbCR9s1I4OwKU
9HHXiqp0JJxOfmLkI/8XeI3HqSF4GXxi+ove+Q+5ywdmjCHoxe9lKRyG8emy/TYg
Ji11Q1VqEe/AbbWk2drR7meozzyiyfokcWiqMYMl7M5f/+fTDp42b0JenC+zZFI/
5g/DHRvHP6ZOLRJ/Dxs61pER9x8+JWZbT6ACZeW6f5hy4DoZJVqFwsCNyTcH98Z3
2/JBrjVQQvwAK7MrZLfvn7Wyj+QHVGp3H7k2H688HobmfamZG04LOQYv9o0h/fYP
gqawk9R9Tz+oM5Vj15GVFILn+WCUj3PdInp3gRvL9J3pitpYSXYAmUXt0rS2BCbf
UDf/hUFdByGwzhw8Q8bUDdSOKZ/wIC4PGzBls5LM03wY48BxRtbfherKogHlaInL
k0N1/BdUBZJBKdPR4FRpgPSj0mxx8lqDlCwv+D/oGM4FCsf4Ubw1A5othpBiqVES
jKTgcssK78FBdNmHbnOEf3UUU1iRdDfGM3/wGo0BqeGa2ETr5dVR8jt/C6/gIyqF
P+WccjfgvPHOyf0Z5bwLt1NQ52bFj2C0WEO46qVGvmFYMiSdIHOm7K7HldTtA4Um
iDiM3xQ30ViKiQ5GCCIEHmkaz3dy0exH+LGjTNAyoAfHOBmC399JyCebOagbfNgH
GK9TkPFwwcVb0sKWkNvpLZK08JCrGcdjn/AzGjaTAvBp9ZkoN5OxWytrltHBw4Px
vGxK+1aB8o6yo0YbaQruOaHc8DuBWtK4hiB2Ni/KVOwXKfJyLKTwTOr6b6qpibI1
dz8xGXzzLeMPu9G2M6lmpkiyN9yUSZG1LYo87OPS3CDYGzPtGn0HOJstaN78DnJx
J4Ms55ZHbYsEV5NLad4sRDZzuiKvaIT1VvmzokEjTkO9zuFZrBqFwMYe/hy+SG3m
aKLWktq0HnLVodHbrY8JoqyRtu1IUXw5//v2zjuMP0xNKZJyM3Z/iJx9tmUk20b1
8kZYU2Fmvpv+1HdmIKvvfmZE5mAzEoWBSe86uilvSTiBdnSEMYR0c/WpnneGR46z
OV2MGDb7FzKBrPn7jSrr8Z8YGYHRSwGxndb9nC1MlSEWGEZ2BfsTQMOtSa3zCX/x
Jv9UMPI+pBwwpnnQoqlWbHU5SNeMSfF7vSLmWMVc+J73KhivBeLBrpF4q76hGk++
ws/CBp508bKaF3PKXFEu8gof9Ui4BpcuxpeaxTYYIVHZ/UTwCI5Rdu4P4isCxEzf
YbPtw2pxCusvd1lvXt3c0pLbIjR4HKjqwfPlpGvKT2cV5bmZeDXoBHcUMbt2dcnn
5hkheD0LVZv4qxGkjUWZJ1FaxQdKnaeam18qPCQtFyBMoEdgjn9C0cAqoyGdEZUY
HjxMDdXVxFqzPHlN2rMa2OJEccHeHjd7ZwrKuQcsxVUCZQhW+A0PbmTkdV3q/Ju4
95svi9D9w6LG9ht4H3f/3SOf4VGP71pRbGclDCOXH3RerTrBtJNnAtwxlNSIoqU+
dbPU4c96XWqJNt9J2UrAVaI1kiObQR/PqwtStD031Ogrgw50PHuZzSq6HUqlZsGb
wGFl4c9kvxEFQse36Q5Ej63DvyEuT30CBwPdUmy+/JLG2ycDqSgPUJ+YHUFbzc/N
IVUFea5InGYEWjpHOHFYY5yCop/t2RMWJ1TmDmgBErA1P6kgv318sRNib7hR7ewp
qDzkbarrlHY1WTU1UeOLhppzQYk/b8WkQfXd4DKDF4seE6Sr8n2XlQZk2FCsvCPt
QEgMff72eS/YD8j0gu1aSjHcXRSUsjOQasUMQzzsRl8qVROVqGN4rYZ+8pSt2iS1
J7+SOWfE9Gw0SgF7Cal7YU8L1evmvs3m1n5sorSTc7Or81nj4mTD83MH57MLCCXt
HndaMHjih+/Qx+WHY0nksdbIIEbbAKEn6IwnpywBB73JXpu66GGYJit143G4LkQ2
q6/lfucOKJq1XI8cxB6kUeGOYB0b02fpmIAYytVC/AQjLXByPZbEJOY55M8+Xdw+
zQRrpy5zaeeQyTxH1RnM74oK+MwIU3bTDTXuW/CvdwDep4Y08Ciuz85qoYP2ynPF
2Sz06kvwViurxbhbNj92O9QURkQpvruKRQQQYCSALt7T8eYaFduuPWKvcTM11O0E
/C9im2c9V+YrQI8CwsdNlCJ14bGjAuHm+KfyPnM+cUzLYxle5Dbkwdz80yeYv+iS
cm/Hdpc8D0DguVKaLOt8OFOvwOC+QwRbACqmhT8FStxk5umNMp/d/dTKC0dP9cNR
/+frfL3m/Ah3otz67Q9FQC3shDeETxOwmZbaPl2ZkOJcZnh2eEVhFwVP9zdPMTtF
erHSGIfVCgett01efczsJxNovhSZaAm/7GJbXBgPSg72onRM6UqW7hjg+q/Qxtnq
ny8Je36DDZ8A9+JsZxylA4hB+Zopm5WVOzhdGz9MOx8zUxny1F//rkmfKRgr/YN/
24PWH2+xOenHMkn9TJ7bbAa3I1Ul/t1dnOSv+r8QYt1IGqIxkxgUhkIz879xZRbj
sog6632EX45/mK4zMTZaHf0xN5Wl42y8jY2U+8GO5GfisiaPxdATe7lD21TNqQEx
CD4ZTh/Yfv4kH9fZyZCD5B3nDM9GjyIYL3dH8qMX8RrPvT4wydvk1z8KXW1jjAeP
vTa1mDWGarOjN+fUhjP+xV/qba9gWDGYvZWXIdhse4IRW3eMamgTipM7FEYIu4sx
KvGqFlPRhyvorPZrA3sODSMqIhrIsc3vV6FaJXtqUCcHSA1o2xR6ySTQbC4NE1iB
uDfvt8t9LUPcNuibP4MdaPucU5dvLjfu9LPBYTZGij/WCjsjjg7m7+HSx2dQbJaq
ZHF9Sieu54wWssdZCrO8SA2eRycDEMX9RbqIt0THdDXHDYPVjhz8BURtMSakLw2W
X9i2xJk2M5GJwyrLs8baVf1biKNBkeRZVC+RaOW/JB37QJWfUy317nsmSbkmaD2E
vM4bmeGIYjeGFZlXD4wX2VKIws7E4tQDXpSIqyIr4cLZzOgQE5KhuW4M/s8XHr3Y
KZbyddNSC03xAhbctmF8x4OFoYJTvvh3sMTj/Cu+e+lr8d4y/EO8UcGHSgLAWJiR
l7eWGXNHqRoNxLtj7hu9kFRLX+Doj/O2ZrgKHxTE6wn9sFiQ8nvqmb1vtLAhD9F9
0I33gidAMNbCzerKmbbFflNA0G4Ka6tHO5PVhTmKNL4VW45WsYQMRrR/J6cyWnhC
noWEAM/seoJ/xFUSJXkzPahTB1ZOu2NsOluYvCR5x9E0Z/pYteidUYXSqb62e1f8
9RGQSvAEwf5LBPqbzMLD4Ogn+/TvhjHCs6f4mX6x0RZgd+xDmUR54/MmPzuONpNW
9oOrUBZARHFoC2DQP+RIq2oSGGvEfV4PUDoWFmuRynUeDIcH7rQ2OwINDkKDCREs
f0VuuMSx0vRqKRUPm9eHiT1jw/3jO6gc/4VIdriSicH4cujWxLR0jm2UmnvvBc15
jYtqQ0FF6I2hqH8aW2rPMlZfWtZ4VNfg9tMZodoXW5TgROFPdjFZpOUsTmGAIjWY
4fuq8c3iEW0bnd8Xn+0ZXXSL2aRvzWtYqGgYgG4mmU1ns8/E/0m8+6+y4Hzhkiwf
DgxayrnpXBGr9g66/HCP8TMa4oBZw4sK8gpR4nsVEupo+ap2iSZ9bNHiiAKNUCrd
Zwg20CA8G/xpTdYbQbArmd5JFjbGIJrz9WC+Tl4qc/5H9ODCUDLF9Z4BTVoYSxH8
0p8wHuBcI2u6nkqh+TyMBBHVSiuZF1SWDmXHNTPJHV1eSgLeR/HuYFslIkvdhKmq
0ZhgRrE7YCuWl/cm3cPT8Oh52GrwmiN1+VhfsxIfWQjq8zQyYQUiQ7yVqkR1QKir
8e5Fw01E52GoYOK2GgLNnLd0vrnWcuNCOdMe6EvIYveP7aO9NmxHQrQRCmKR2ksq
fXjrxH156OWlT1HdIT8xxPlq1vAltebFrF2wp6a8BEwahipy5qYQsH30cU1gA68z
vR+lRT4AcyWzpeFM/UY1CW5rI9ygyFskK/CHsOQ0DA7uBO4lWjovZuNzr0HH23nY
r6iyP4hjFYPw+ipA8dSK9yPezFFmlrvnlhWf+ZTTdA5Rsq1uYrYzxgegs8qXauRW
4NVFaVE7GfeLt3PD0WveG22Fi8f37UKAnu3uK6WsQHCYqOeQyUvYD9kVJmfmae3k
gBN9tg8ysltPIYMBuc+KmyyzsWRnRkTxR6+bBUAeZYg4ECO8GyKqCgayExWFPPIl
boMipbnT50+qeH90MUZd065Zl+nA7A8auv7PqnA32kVFuC6pHEjMfypiuPIq/wfn
clexakvWgW0/jYgJAKW3pCpvfSGVWk+jNs3AgAYAl27OK7K3tIS+OU5Cdhmpjpy0
M5XZgRod5EW7aHDajwmiHDspe1xfWn1o/dq01/Bat7pgVwtdMwp1B68PizYchXpD
lSu6VguPLKKSxoAnbqKXSyVbuv7zQRvi5FegMD/TLsXgcOXq7/MSVhVl8cjk8nGE
Hw5G7zbx0WnQ6BMuLPZSPWScicp9r3ozcr9YjqCnlrgvumAFS3bmJrW9O/Bkpc1L
IMCFpkxX113uRPktRy6JlBV7DgWHuYp/wwJk+uKS52HRUr6PJcl5Zn8jB2P4R8UU
LhHSa0GO1urL0IvnuzM0ehCIdHHr9kSGpYskfdstHfyXTtidezFUkjOetgxTo6i7
LDgPUNYmCzibjZHLRB6fwo+L3gPbj2tjn7yu9u7bpEoBAfXPJW01fi9nGaIt7lS4
aIsIC9baJVv1Vshdq3LhfPk2/HRnnb9ko2Bw9SNJMaNC6yPsb8MQjvzIwdZoESDw
82idrFlwb4ybvz5XqoRBvUy67lm8vPIHXKInFT63TkTmWRVkrpUzWedDJHHTgBlB
dkJynfvLZC2316z7oNCFoSdCddoLGbeTvhyTZqYoCD+0DAEbfVg0CYhOhlfKdZT0
k3lnMouKGp2y3CdFrga6BHkwsEAPRpej1Jz+IBkyp9YjCW+QpKBeRh2SlX2ZXlm6
RkvArwoa+gtOkz11VMIkqwfE1Gaw+2jljqhl3PfZtWAURvVghlxKS1j1iyNvUlga
x9SNjQohSFrrSZwMb0/qVql7XB+7KAgsGJKGWkAQ5Un96KgToYO81RXDNt+3ui2E
QD7rlZKqxgKI5PlWfuMrEwI8BVuJfls/jRb62pAe0x/r8zghAKjmqhIJRc4DDT+n
6HzdrasePO6yI4dBFbQwoO7BDaT0f+Vyj5LnYKBB56KMjDV3MeFM8v72Hd/M0Vsa
FvLxlDipVPN2bDUszI79QrQ5a997eCeJn4N0b3qwb7bm98vYgt527vbN0jR469Vf
swZRmVHEYmMl8U4Vwk/8BmDqS2WUYf4DvpeDiyOJ4u/vxsmvJvl5v0VlTGM5ngps
Hh8/xji+yQrj5A3fzmKyyI7pkpjGxcDSLB+R002bwRKuAxh2rLmoiQgpiE84uJ7o
woqhbrPAiZQlY26/ZiJnU2LLWZl9xk5KqWSe6bXNzJxR3buSsKS9aNyhjm5XopPZ
d1VYKyJaPDgYE/JYoHVhOg2iPBPfyzpRnLaNxyBQ8Ozv8A8bg57QV5k2dsa249+T
krnFVBrS5E3Z99wd1S807pCz0grkfm9+fz294ShHHD5iioQS40IdJd+6WaJ6xngZ
kofyXOo+2TCFuQYpGENRU4Sd2iQVzj6mQpNJYV5ZqNaPHZvYYe9dlHw/UDfnsEJJ
LV/YYULDvPkNBE+zQWcDphyst8jbSWZAqQaVyzRYQzcc4jCKWnodVKCixtn6Wd9w
0jJSdT0ERWOCLFbmm8S7M9Ocg9dK/kJpQyid83GGzQRgIZ08nPl/1CYEJPqX9ihZ
2Y25vKXYHQsVJTj5fkUo0eAfTZK5pgUXB4Pux5G+JGBkjwUydelSftEnMEZjLt2z
b7uqhbXpVQLnzYYV/zdzaYUwYQAb5N4zzlCsvE1hhC1anzmDIhqUZmCPlmXbRnu6
yd8Ei0spDZB5OfDeIjJPmzWuoAa89dDhIaH1uUeHjueEGKw6UndEAkhhI70LfIg6
yhkqzAZ0yQaGUiL3i0u/zdFqRnRbVM2OXHZnn54+BNcuk0DzQQMn/IMadU1wvFPP
VbpFZwmkbIrJubvDaWaMx6opehkL/UQk/kyDPA7Y6XTykde7E42hTY8Djek2J+5T
U40aJgFXOMEJaFiVLKZSSvPV6cyNnzUB5piRIE8p7CeZ0Emr19Cb3OPql42EvLVj
Nx4PNgQQLwROP9GsCtU8t0xMnoUF/6KTF7C8rzJVm2+RRZ7FNb25dR69YUtlE/Gm
QIS9bxjB25xiRkR5EU2cJQy9qLPvEZEG6FHn6voj31mJcA2z4pD9qbI1aKtG467F
3MfZI+S40JMQqZKgOvwU8xz0jhE06OlU3jQJ5ZxWgyscvhdyPsJEUzx9VH2D4bl6
ibbL1ujN8/C2UbGQJ2XrEN3iSgLAT0Ivirgl4wXhsP0GhrSgwLwCy00KZIw+DI+I
zQCZCIes93e71M6QC2qF/v/DqmihohjUOkHXh62l7fDqVAXqlbDKE6y8T5Unm1MX
LtH74Bisbhz77lG+OZIP9b3EmXe1xVCdgN3XurkYNuZF9HgZqy+J9Bq3CHSxtkMh
n3hy7srhda0HTpYveWM8hv8FunngrEIBj5v6lmpI+ziXYhpBg72OWG21DC/3pgfO
3O11vRKCi710+i09q/+14v6mG+p+rgNXqW0Wtty3NHtIvW7x88Umku/E1aCTKT72
2W1I5FcnS93UOhJUO9c4RngWTYT+ow7DqhH6bkwazArhgzm/RbDCctcOBsmkt6HA
vw2UjCA+VtIFQCkU12uthW1Bq9IZ3JAeOjG/g5dvYm1ZBwPJYsFMYwHIWd1Gmmjq
NqMpTjVPuWFEH3HfEpJ0DmBk/QRLj1njT/x9OETdnt/CmCdlknfUx3Vhw+sGDtRb
+GGOCI7WMN1h3Wm5lzAKhIRJ3CtVEkbqSgk82tOdR25qC7EHtFLZmWsvgvvdvbKT
/odFentOacuQ209o++zrs/BoaX+eUBixRmC85en20s9czcrfse9aNVMh5CmdheSa
AaLY2RlFRgw1wTioRPwN6IXGTb2bB52zpCZhUw2w7b+S3rMqXq+EIWzeCNK7Klz0
mG5axB/HlPKiQpzq+UMFtxJJB2oa4ACp98DXE7qgcWOeCFsBSRD2yqJc32xEiqje
2kTxQpodGyr1Co9d1jXw6vOG/EkFFK2jjOrgBeRZHP2ix+imWx6Endj4AYDF8l96
WeIZDYuJU+AqBDUd5Tt/KIHegRQ+wJEUmJFjRE42uyJfPWMph1ggQtXDc+2MrnBW
aBFnbTJZIxuMeSbQV8q22segc+pXub2Z+6x6YXRxvR0ZjJ7npsbSOqLL7fax5v1l
IuPKMPbeffoHMXnv9/zXbE0y5K7HC2IBOMKgLaprXyhBnHTOpO+833wLBOHaGLQN
9Z6LbDhVwp1pAF2huLntJHi/3U3QAqOj847uC8A0VuZZw7bvNxpjl2o+zfXp+Lpb
EZRkh7GPtN+ztfaL+kU1FivQ5NRsyVK12WmcsNQ5iO97Qov9tMpViFG7KQkQh729
YHuJ7LGnBoUrUoxXjjnz3aCTmcQwZxDvaxt2YYmIRU1AQpkywt5CfT3e1T8/48sB
r5uVX045KebPvR7HMpLOmpBvWo1/aT5ujNZfMtzdj/lSORFsZgE4/gFSX5YWCC2i
6mIzpOr6rYW2Bf08FBdo0Bm1tpxGKdVbk5Arkmdfy2UIMq4xWCYy86tsX2csK8qe
+HbNeM3KWS+nSHLrvPN5L7neacRzwmZc6aLiMO0to/d2sCk4utCz2c/+wxdWY9DX
s2bWtFsJqrlWjD/1L/gG6FqQuxbW0euwrUx0Rz4ryVj683I2CGptRD+fEimTIWJl
B/nQWTT7n63A5857ydYnNfNILTwJElhwjZrKKAZYrH0WFynW+SZHAlPOoRyEFXXz
LDPgj11C3mAXsuFgA795I7SlKhS4pDRRWUBQ2sskFK6cceKSEyAYwCW9aOk1oa56
UDAeAe3D+DGQRaV9XucrSlGPuSiqF9bkC8hT3/k33F6ynQhGzIwMgoEtXycR3NYB
2SJ8gxf5smy31vxmsBsj6r9k5RiK/gbbkzG83cF+rbNqy66wmEEr5Zooa/nM0Cld
PjPkvAmrPZnjt60J0um6duwLgX76ky6TG7nYZoOqP3Aoce1M5ZlYP0YIadKnYy+l
233ASXnhc874Eff8E/RULdXzA7WX3md7lOA7m2mRGNokYIu7PPkb9oWNP8ZDc/9e
YWr5OIe6rlUQjnFz/JLBHK/i+JQrXa0YudcZhYv2eu3G22tjxZnvY13usHO8zl7i
QMJn7Qyi0CQqwGTSUslexHWB+B45pgGoGzFAGOKw9DbmM3XSW1eYTOP4MVPE1vZ+
WukUHpJcDmILxSds8P3GKVlDm/RmDAthT20wK9h8OFQfGKAXK+ZahRLsEEZXaiX0
mU9YbONQtNqRANRm8X+f3FS7iCuJgfnr/aQlE+MMpkukBsPeqq51Uy8Z47Tja3j/
jDghOKuVako9ojJmr1BF8/de9rULiIU7pSjGJyB+y+5YLNHq4ZZj56TbtyWyvb+6
vb6RRjrdKjPrcO+ji/pbLtFiZoEwbYHAkVdTbCVi9I7IrDY8Kx99Nb2pBhnSd3xQ
mlApsCK6kuVi02npwEC909lfcy5fa5DSHqlNCUKwdKsQh0ssl0DOq0LFdg6Rgn+l
9nfVcVnIrSR9zZ7MIFP32PpEC8I+AnhYhrt5l/pgxI2PDP97vLOV7ZnqHXub0Drd
+AjoTM5Nec6OTehPDuoY69N5EGKDHM7v4m8cPp0M3iKqA9sJrBRYAKAFDdezJgfQ
/AV5nOrdH13itpEq2PD7C3sXVMCIlV7bgRwskrJWlCetyg/zB+rD5TzGIYRNJiIB
B0+dxcgKsNDjPT3zXV91vw7wB4GKXaWi1UnAEj08SHYPOEtMaFayrxAgj0NT+Ed1
BhLf+pC5J1ldm48C2ZBPFNZ6qHyG6sOa8oaQp56/sZ+aVEAAggYROyXrEXtD/37e
RJjdaHvZczscCEA+F2kYStsoPtiKJoexkYipxe3ToyL8zgqP2/PwxqcF5ITH6v3x
1FUZrS7+OFZP+F9UsyvU4h+TmtoQYa8auVE/ENkvZeX6V0/I+GwsnK5lHMq8eKiX
p8GdYiM3ylNTtsZlbXFlZKWzsQ57wiRPEeMeQv5Wj23tTd4K32e/m1yZ1BHa7bFr
PiIf0jmRhWSKAiXmRxJGCo257c4WymgEj/O8NTQ5icxraPfvLN7iWtJ/bIGcAN3Z
TDAAC6rutUuJ5VYsOw+0h6QDd/FvF0z8Z5bLaltojB+77GP5IP3pbI61nIVAh50M
W0IHrzt6fdoORwAkGOJhH9SN9Ce6aj0ppXnwllHpp9SQk1eNsc5O+ry7eek8evjg
BmIZDg4wT7JXQvt+rAZG2uFf6VBfu6HRNBpkC+6Lfvh720LxK71BSkStOKbeeNOq
K5rs/cjpjt6kxApE1DxBAc5F3nJjtZyq3+UySGFip4rJyotHsmyc5iYT1/nlcyBE
wh8G+v83SxGpHmpw8x3H6wv8T7u9TsSjlXr32xTmoCLPBEdLAvt0krLbrrLG1f6n
kV4sUYN0GH87tKbxCLDurQ4pzf4MVTo9CSBFDaqGyYwbjgJ+RRLA6F356hML+oLQ
OevGoG5nHLxqav98v5xH+iBa+XXqyprTJkkGQsfZXBx8dIdu5SGg2dtFtQWVZ/OC
yC435AGVjTIempIDBLaAIIVSv55LElwSnq5MnJEWP44OI6I/1KMANXgdSXoeNBNx
+DvDcF8HHyTCr/ufk5OIOJCfaaRqO1cFy/ywt6lQuVgn4Pz+j/YuQhBOamhvFn3g
nDMw/VNUx7O2oZVWZJHi9+o39/j+Et3RmjAtFvqorzNgW4XAnKIUmLAD79OUxEOI
nBDE8/XPuLl728GAO9DZUz1izxR869zPK09M69VJOZGs8MJVjUEmVUvNMwhFFu3G
Y8c/6RmMkcz4OnxbyEMR+lwv2YXYYGVX3xj2VNEpYGT7OlqjrUXQFJ6jQ7A0Ql6N
MVpWZrVVMnn7NVe2KN31Mp4XmVB7OVdEG4LOybo6zlTlIRiX7iT0h270L7Wd2zAE
MOF2x+toeEGyfdsRMAqZGD+UbYK3dOZDHK7lLb4j6ZuBWj2z25ZqeJWahaSSZ6cS
l8Z702gGmPC4xZAGYmn0rCTAoMOuTsNX9v8LRIWmGtomeI+lo+SHKh3QwX1cPWbj
r1690hjq70++TZuP1EAOhfNLMXlnEbEazdY4lEzpYxv1RpHC/Y+kA2sIwPTTPDh/
jL3jXTJeeE7IBKLbRC48yOeGo6tCywlvWKCI4y+FKKotsAqami1yOKtfobqp7Uyl
Lz/6HdRnY1NxGeZPvki7rjqMUlLC6EkU/WF69Mri4w0yAyzgjIo/h4lpnWGGqBFo
RLcZyl++A9zXGyEX5uucNRbweyCSUyEjczt6l7fwid7crdVSYxMTZAV1HC04yp9X
LEsaRKi0pYOk3izT+IcTLn3a9+Rc3juXC/UxaKj/7YUP9ergri1Yq+Su1aUAgDA/
fk64UrgIubyDpyqw0uUQeAmCw1fq/nDCvLxBXCZZLsR5xX9EmwMaD1QS5HZ2dwU9
/5ba21JIKiWf7O+o4Ev8qr03PKV3jqwSWNk/NlBHRIXgciQRNt8sjz1H4lCuGLlQ
V5WAQAtMDi6UaqvC2OE7cv/Wl/CMU8Bkt/VdA+mfT+94f378dbvgKdgsuSnZc5ow
LCq8R+jXkx6CZpEGqASRaOi2uvKFDikEFn6CJjGpSqHJgPTBkgZaa+aeHrXHhW0B
0J2rPrOvGnR/sNLlggSJD32gMie7qYgz/XZqrAkRC9hH8tLJ4PkQuTTt0nlniPk4
Cfs/KSVnB7t7G7Q6mtNPhQpN3vJ4osbjXLhh3NmZnusEBhjLGcxIsBPWmXgaIRzu
UfoQXliWGHMz6euay83SVQOdnIIMlA0lthWXJMoJgUSpcvx5kMKlHUrOM6G+OXzR
MfvHNnvFmGdJNg35p6zQqlASADW3B+sje2d6DfumDBWcn6eXwxC2xnm+DC7evL58
lr3h3KT3gUoDciiUL21Ge3b0WROJHLQg9GnrGEtF9liUT/pf2qrQ7/A7Im+cTy/R
ow9LrSj/189A7ujeFvx3pVYMXShIikfb7Jqxpg2GZS+mrNqxPspLDZj56r15x5jb
6XULmQ86TGSP2+NSwq/kJejYl7CzgdOx7TeYhff6AaAsArZhlJ3kN1H6B+eJrqMe
LmeuWtE4VNSW5vmV1migSj64CsvvhhXrnxNRDbguxz/kYqJ68sMNXVdvnGDgt5Lw
a450hunn4eQnRmXhHELxOHuotutIowSkn9gHQjgnwDVbIh6TTyVTVSpRYX3ZqcVq
uFiN5Mfk2mjBCnbjnA5ZBmlBk70TGs/1gHCvSOOKu1q1oZvpj0SuJwuQMBDNwoRC
dNyf/lqRKqcWLwH4blGrAly3FZHD9z0HlFsvU048IqupGvG5r9g9SGeQlVdjW/y5
notKOdqETHnReubhtgqLQAIKzeSiKFbLENDS65PEJtYK1OpuuEyPIyEHKYDwbyni
nBPnRhJy4zvxTnaJRSE0gzjRvUv7945fLbGezFpTNr/aunF6hgLLPWw367cBkLB4
2nWs9bzXNIzsOhlQbss2wdIaGP1ptwHtosAEb4VXLLf+N3sXWDRm1GWYLL9VhrfP
jP3Xa6b6r5PmeTI+g5XqN9TNmOggHFBWe1CbZ8yyGbhTsX9VcbFdpmYgbVOw48XR
+9lPZlfHprV7n3S+JmtGv2B/IYP+cN5p1/R+86EDVbRXrZ4fU94mOL8mV0QzJVKY
HiId4uY95IkBIBKry36gpDgM7h53dXY4KyAYbLZPN3QkQ0UMr9unMqsEhIl3Fpda
RFvCUh5GqXoq3rTkT0Av8GKm1QhFtI0WUcJhJTzx2JTnb7hJpgkdBuevYNopqT/z
jhMUD4r+EVKgZ68j8C2nvnkV4LTiYvh/wtRPDzs8Bir88ahyOSylO66yeHGWza6r
sB/F4DexzwgvbMmQXSbBl0SFuEcaZYU2LGjJfMwVWIGSqaO1spBWzmN6MaCTLgit
ycqWBmp9KfCzyyb66umh8iItQJzIaV+gsAmu7sr0Z7n/BVCrjqJz6MOHgB5K24A+
SsEOc0fpXEx+9MRnZiSlN3OLiLo3uPQ9MHxcNzDxmnxypgZNctTgnFmbMs6+N5y7
V/aj+cHJ8vNmElJIXJlBCbM5FmJUQeGDjqq6rUGivOtWeYXoaLd9Ozi8G2yte5AY
YTfp1LCSaW/r4sGOEcfGolxywZIKTQnVePFWQdMLV7jYUI+UGG04m5pNPI4bnSXt
tLCKYXpX6T1T4PLkmGhwdNkeNm8jPwgM3rR84Cy+7IcXxaDhKzkyoyh/oqAM3fAt
JvtnxFPNlre3l1HVOwa3VQGSZHYO5U0R0OTxIMzYvhUKgDw/exhvshJqUNcYR1p+
IroFCRtNPwsziveX1cTqirLBs70ZfG1zSWOcRTvF50DU2WoEmbRWgBRgejf+PJV4
Wy/TgnFlxaYZ23l2Z6CDVyviTh2FesPmsR6eiveMWzSXM6merMQgwgsucl/klMM0
aj7RFZRpQiEDKWY3gsw3+9paL07JD8ZqrRUaeXB/ZuPXa7Spq5RKrsUC6Ab8AjVP
PtuiQ5B/YLTSsd7KnQ3jBmlOv/pIU4H89cbCU1zC7nSVXO/XpzuMtOUx3ADRbIYP
pDZXAB7FvQ5qEuYnWsUbbgAJpuKu3pxk4uMjFCFJwhcIj8LP2qWa626qhvsgQ13j
f/rL1iwO2RtC6qReBtQXMt9+8XahFP0L3kUkLbtfJPyGx65KjVx5zNQ8nFfKIleV
pfsib3z/PZF3FtH2wbavF29vmwZUnYUSzxrx0jsKTeFPhlNJVF+BlXM6KzshK2NW
phSdn8mO/NsBLT7iNDmzUIQM4JfwknkZwn3LQkKMT83enFWX1N3tSq1GNMKAw9CO
7kHLQDVNyZWcN181si8Jj+61oEOJqfkBb5A/KkVthnKxaqg97sZhwOHReMtGCJaH
vGQ1bEa2MYm0995MIAm/XF2B1DbbUE57mkwXGj52GYMVFUsgvyaNCl7rcwkgAB3p
O0cYHezStk+FerP69Gwg/RV0PlI+UOEFPlMQGvEPhgwT6XLMcL6a7ga6JUsE1U3U
qXdjTBs3RwGcSqQLF0Zn/0PUst9CXKz5y8QVvpGHfBX2lnJxkEi/rU42NYmQZZuf
uhfJnrYZOpjfdxcwxjEiSVsv9Lfw/naEueUYKTY0RRqP50sSi2kNoD8iBwK/Rm4v
y+rQGHPvmbe2i85yWpVw3bppPaEdOoAxfdL9KKE17WRvW/PrQBDG2ORCEKzvznJx
6VkoAY81p5F/hW9GExtBn9YUfQo4qdVnOh31920dGaeyyqLFBKmdRkQT6mnzIwqA
2whjwFb+RhyhhhUm0vfaGaB4ueXrNwQq52Aqa73h01JOuKHnBlaG3W7ehtWki6Vy
87qD8WEPevYMbOHa/GDAsYuMNkx0SP8dBYwmEy/z94GZH18tNeVp3V7FkbFcwRxT
BtG6xtaMy5oUbQIi7ju4o7RCPBsPGpHkmbN4KqB/szxroqhfObhsddQy4uM0ZBpr
50jI2WV72zEqYePNyRsLYMvs+nRLGUFBJ8Owklpse8hr1mc0rhQSlwgGVrYUiFDY
X49v+Orn8Yh1h9H+4vgjOI1qy+HCLhxvyZ6XyL0l0mqPxzxllWqW4l45LJKgrreJ
6IcSyjrn8KxADvB/vm4XIM+7oe+cw76v9f/L9UBI1u0B5Z9b5+eNXz9QmZRgZoDH
cFYpxvWDMuB7pDhmrthTUF3+8ens9Dhwp+cjr2Hg0MUbueHmMKJ5aORnNgJBiqU3
Kt3zs4hRWv328qZX9DcL2D55AG/fs42J6ypwPK15d0pt+Pi5mOHRwOoZ9vUOIza+
jOC6hgExqXYsUfKMJgPaRlgOLFVGyVwffoIFUqpLqYl2GNBCUwEiktCeanENnakt
g2s9auuKeC2bY08IBxt/x9PAsPhAqV0G7gi5Qp1AqyjSUZ//+Y7rvT7gVijaZcUQ
iWil3akLTqcgl17A5OE5Yn8Fn46V75yg7pygqfJqWEU8+qC6kQ6dgv4iSGI1f8Eu
kh4XR2F9xBXCQMIYaIGZdXXLCe3rYin506znLvWkZOefQpmCatrSZmqlxIjjzDeP
a0uCpglrnywioarqIDhPLK1fZWYwGjDFI/4evi9lfgME8vySYwI/6UbbCm1PlrLt
GhI1BS6+Knw0WoZEvIlBXCDQdbq0OiEBhwJARwijRgbF4GHwbYTbFDDmOlGANtP3
kL1zEz0OVii5X5NG1hrQKEJ/cC/mIr14yHvTPQNEGiZk8acM3rQCeNwTtTayYrsN
+JMJxUKnd66FFlZ5IlB8bjM2f+p2dFRH7cRojvawYCwtmMxGZxU3CB2PzLpP4zEd
aobCj0jBi10Qk6LIg9A+D1+IVySBcO1fmGddlE0Ygf5eepEndf+BlcA59YRxTI4v
wCPERTuPt/mDKmy42w7MTa0TJZVe/jrTo2K5O38KxTU86j7dVG7sWX+fnLXzAfyZ
N+/cjhtETA6Mj+PhJBYlYtu6ltxOGDEObWThsU819fkYeH6I04iH6oXg/UG94QFb
5R3LXV/YXTLcd34Vu3Imix13I24c6/cfE1rj+3AfQbqSFBY11qFZxkF8dw97mmZs
aNgleolhQ/iydq+mjiLQCxQlcBFZv5wKCiYRw2x629myTHg6ZoaOMXZqaLmY3ANn
M6GfCDde8KHn0p66TJkKTVhpgjNixj2t4faF3GYVgIsCXpbMSjf8jvSCn+Q9V1vH
yOmn5VnlQ5RCKow1xnKecF/eImWBGasGYKIBI4/F48woxFKSnwMxX9UVHvK9pkBG
sUBXc/eWhp9a8qMK5bto7PL6AFPKcfobeupWch9iTvtJHXHMRLdMIBLqmK9/DoVL
XWyv5AlloGS8sY5GcppLdN+sFwy6gDE97fRRtRbWkBsWLec19agdvGqZEmo5cJGz
GtmEn951fEb4qZW2COhnTmSpdDBG30YtK5sdwfI8l1NpAMnwkOP3H/O0K/GbID0G
gYlbbE6A0j+x1/pALqYnTtjxDq+ycCmgvqz+fc8+6FHlM1P6v0yLzmb/O8Tf6Kou
4h4nWRShBxw5J7YtmD0cF9rKzB09WeIHI/eewx6vAa7Pwcvnr/Vbq3mZrZzE4hWs
Q+J+MZEd3TQ64smiI1wVdGfDDQR1tYT5dDKvoID+00k5Tl6O7ffma3uu7oiabfOu
Pj4T13t+WXBYMgvvfWKfSGlc5GSJBK81iBfjiLDjzX+hVt9iQRYhvpA5g2qXFn9J
8pJjxDJuEECXlF1rqhFY+L0JHiHCJ/OVBuz1CHeCDXxfTHOhMoVveoEpbKQfwbMs
ltIyaYILAohx/c8XJGHfW6G6VvRsYd2B+Cq4FXf/dBUlZXX9rkwBP0BNG1ZIg7qN
LKbspEhtX+yxYgNihYFwC+IHTyGXl4T/heF9NQ6GYCO5FePwT0aDOkbTNMpip2wK
kYr90M2iGkjH3kP+7+pWsZsgKgufyIgWcKrM0UpNPhs6FW6CO+GWFrJUxfSAKokF
stwzC52p6Qqg2gN8UqMDshyRT+92uBRLjTr9uplGOw8p1U/voS6fAmDGkKEZaWzM
Ah20nqFCj3PHMgzW1nwgtOjHunLcw3w2lDVD4yuH9aBicn4FzqCtJA5Ahln9jX05
i+I+/Gijt8dEWBRD40/PcgIHjdNBlZdnVmBv3tL41unABdSi6lKPuv2SQ6VPHGSu
/rT+Qytj6tPQ1YtbLe5eBOlNA6bSPqFbe5Q+yI0LuGM8Byg92UcClRJGPzkMgGYM
+dLk3H3+asFeKSzsKfwjYbZBlFopDL6712n9V2OG3u8BhAb35NLESmTTIY3oi1IH
GyQ8p8RUzhMCunFasoCwXPNil2ELPJpXp97l99LBw+q1ysZwbK8n+cu8ZF1PNAH1
M4VhJhz52sMPBh0vyc7Ugx8guU49xOCtRbrqCjxsrBvRV85jtWtv4eIGmuSX7jiV
RK88VcGp4gB8aRXdlKU2VJVQVCjtgMC2mA027xez7Ty4ffCZtbAfA0yHWpHVclDR
NCrccULjUhrETXYLjKaqXEHnl0U91P3pW/9erplvSe3to3FUGENE5WSdi1QkIw/J
qQaaXQppsNth9CROeDgG2Zhy7gQzxn4tW42ymkaHS5DGzxQ8V/4/H6jH2v8c9cdY
Q7qcUSbjml3OC5pk5mMpfFzKzmbVQesJqAta2v6DgpRLUz/czWztDL23oXw1pkTq
UcjDMvO0aW75RVeADCLx2xTmlS6O7r81kh93/zkx3FuPSPSAeOX9ZPzaRn9O4Lt0
lJEeGKvlgYfPt5oO7bRZ+8N1zK4r/M2zOena8kKI4MyJW2cSp5ORuTO7hL1yhqMV
Lpt1yijQusUGXW3Ps+20a+eptzvWqnvZoRTpWymW6CBV3rM3+ht0X8SnPBKk9ju3
MjZEh6wG1DdgPudZcLeC48po+EpJVXnEXV3czCtPeEZAbYMPJdKgyW0uxsBPRkDO
V2au3DKr7BNi+KFGBKwFl4bs+fX/GnEoJlDvbM5TDTIvAT++2/FINJIfb/isTBkh
YtOWA4JEWv7v/oDlJ/lszbHsYkSF8vfQ0JrE+e9uBzdLvI6Z20uM0KNUTIECOThq
Yw/gce2l4VM8fmT8T3rSFKkr7zvudHnusJPSzW5B6QIJO141Ud9v3pG+7zY4Hm+j
OYMi1IzjQ0kPumDuflLbe/Zq1oGbgguIl7jxkjXzMmaRHX+IZQ0I0mQPMH0hJtg+
1QXI/fyglsPdMUJlVBvluLC93Rq2qJi7ts9lXGPgogdf2K5s38PI1JS0pCuU7LCL
6vhtjRdYbX1tYVUPxViMxQTHJrHjnkpeVhsWW0z7+pNowS1RmGZ5rHtq0KGqLg3a
Bz76wKFlyienmwwZiUHLXKVw+Ijiesp5uIlynJZfkHFzkRLRNDpdUx1DaXYBzrMJ
OhLkWxhTmqOjMtI0zwLsB9E3f5yzChvt4nXqp6VxvoURyd/wYkAQKdQbtd6iGiH8
uHdJUnmFyR4N+mf2NcsOVx4XIwtl5GDrCm19dlgecyrT7hfdW6Zd4QQte0d4CpD5
3HlZ4JmEqoY82UOuZmyPHtovQMc6CX+4bElKipMrkTzxHvcx+gKt1UCqPZehjXF0
pYYibOns+fbgfRi00hjFp+sSHkvTunEFotW6+HNB/dMi+5DbDhrLxyk6wVS2HTPF
GpCF+NorNPIHnpG0dALZFaSnm/VHbXbScqnoDsJKv7Vh/q4DJ5twVAwY9tYPoVif
UPSO/6DJSqXZhw8D0ghfzzMNiwJu7slv3OTb/8UKC49q8Ht4knqgFwrx+QWUS3dv
tM0VAb5uHxIy2Do/ZEh5NRfFZzqR/P/hoIC5NVsWuq8YCZM9ds8sE+KE/WgHwB3U
ivMaj3YWYFJIrVu2+UBFRogBNCutXI1+Q8SnMGoXj892Fhx35r6FvxPcsUA8FVFV
guFOa7KAfLGhwMZ2HEDUO5R6dQgOtEoC3EWuuueBpMDHgcWIWZDjnAfwI/wrjK/S
JbCuMLcso7lnpI7qSm8zqeFzOnLv9TIksDTj/AGAy5CC6WvNgRnxaZ6mbxd901F5
/wUpIp+acjisFOJ1v+dN90mxOnhTH2SDHCNpDqo/RZEdNJu8H2rolpaVDh254lko
jG7C1drc7IpmsHRZWE56BDeQaCpkVgBSV2yZQZiSuIIuV5Q5tv+hNGTN2c6FiX6/
KU0F75LWp3S9Nb0eVrDjoLIa3RAhDaIjjCck3FNnsXQJtJbIottzixRWrS56ZzKy
cQ67inVok9pET5iOBKrDm/24kIOidG6pBHFTpJOp+PCjSipw1XtiutyARt8YBfDh
bcM2NyvnEVUVvx/2+gVHf/uqvnQVtt3wyCPI9vGmURCbLa6RPN/eEjUyGxbNnAcC
iASYoDrQyOxlp6AF3wxyaGPwbOHwD1EEh6NsL3kg+shv14INvO7jwfm/WzHPdEfH
2cpA6rkGImu3uaIceMSN04Cbu+q18t1OCyjK/gm/6eJcjor/J1Z3RJ13eJPCi+IX
1lKq6EGCoQ9Zbhv5pmebRB3jRzwfwxWzDG3fOVuqrZfKrTVqqO3akychGHXseKyL
1j7ZbiP8GNn3T0hOhgVBznqlYLZUpf6Y8Kfom/vg+RIOrfp8n1PhatYwBA6N+nw9
iH+Ir9CNKi90qJ4emkPUCFP+L0zS3CtvMfdMzbqyICteCpUZ2zWgDxE0ihoSvMF4
MjxbWo22PLMeIUXJ1vGPYn0TYdzR0hlWOqZWv6wmS2WtFCLkWv56wGxOIEUORpgc
E1JJvC5jCSf+SiR8puCLh+ajWvYwNZdRb82AKpzBGn6rOHR3rIDDbJgNbP2rhNlT
Wn2jIJdYwoTnv/RyWH9PfbTJJ50xAwAUhDee4I93ROV5QuM64ISQ1tBdHGbRJfsj
sRC+suBQgXUbAF6Ax0kr/CKehaRoqjGFh5qKPZVPYFx53l0Up1PkFe3C+ufZVlWo
pft/TyrhUw7Tjs18xg2KL2AOlGInW19odo1Wm/c9yJqqJ0DFzhq5HhyWFYiXq3Xm
cuoOLZnX5tHBj8si26ujva1jhoqYXcu/Dh63soXkqiWJU8dI+CC+kDrYM1otTO15
LZpsO9s56LtfFDw7klofAy3DDlfovkr6Q5n3+S8511uc/R0omzJDg0AvAlHy3JsM
Vat760ZfJAmwgdxkXg0ygIlZnXCKdssln6KlC/PEOqOVSSvqgsiNRacncgY9GiaJ
Je5maM9SN/1XRtMp3ucU6obWdU0Zny8N6yPZH338TKSO0tVCSzNc9Ux6tGKQ2f1I
id9dfKQAq++1FK/PA2i9wQGoKEscsXj27szNPc0gEqbuQ3ibZqBylJ55B+XtUMkU
HP+oA1R7x+9buTLsOeNGVhrH2cc5QmyER0YAM2KXhuL8IXpQz/ZAT44jVWunqbX4
qW6VKKapCUIJbsFwOr1zcxC2pRT6nnfjZEug+1SYgGRkqHNENoBURqcUXX55RH7U
2LrWtOkGaFgadOoDBs3uM6kAl6nNRvqukhfD+uTItSEeZB+IBjQunLmzhRW1ZIG4
W8K098JE+Q1XieYiOholR+5TomX7Cj7BTKIcULx7hKenKdATsPya1JZTosLk0cjz
KQYJNjAtkoO1wsXy9yVcG1xJr7xR+FyROs0TCeMFSd36V4wZgQi9bSB5BPk1jDay
BbnPOof8F3RDhtdG2uJXUnG2igTihXOWmNR3G/Ofmj7figu1O2hZ1sJevT6a1wca
LWO2Fv4sXMLzMrwyEPcPQODRz8ZoeYlANkEkuGcNdNJkGt7d7yb5X0wBK81klPWn
49SJXUKmVUIQhS9EIfebUwLwrq7bimXr86jxnUycAz8nof+BAj/Y0bZ58vGzu9DV
rQyWvJ1F1uZOPUtfQaSpVicq4GRBlQVMqkYOPpL5GQzeoTU9l7BUCsqOl56uIpcu
MlvgxyoEBtDKFz49C4rLyw13ehvtAvSFF4uGnP2+btjLQ/EecEVD8SQDRDFt9YHi
SaCMukBM8pCXUg/DVN+B4/hmNYyQ08R5qpPo8zu88txIFgcn7/gYp8O472gdXkfW
FIULFc8YQFc9cFhcQpalVCM+0h1edhFt49MCMJTDF05eOhpFn8MN2HzsNykG7LRp
Yd3r93SRQtcAuEE+0TM3e4ib/il6nZ849YelDsuMbq+aJq6SLvi5UfHvxJ5j9dLl
aDnllK5X6rJuSUA8x+xRzCFM+q+yrxU0zZnfEPfO7wdcCWh87FYNlEJGuQZ5tmbD
oK+jbvlKPLGlY1mKUyK3/Mnuuzz3K7sEoB/eoEsNiTjSWnuzCjf55TRb3WLohICV
DTrL6WUFHEzYtDbPFUygnlDKwEI55AQmDER8mvVx/+g9uC5+o/wFJzfW1Aygrj3S
fS9Bsv9Tf8YAU0Q9cL2qPLfULVw1FujxI+H3CYOlMkDM74ia1R69AUXrV8UefSWY
BS957hsxSgkWqmli7AqsMMaDZVAyEQtizCDVW8kIUFONPsecPOV26RKfgwn0jeKu
RHj99zwVMaNcGUIkEB45eYj84PEfx41P9y9f4Kbjmp8flBr48SURcK8F4lXDmGDx
+Ic8s2eN+K3Ka5gvDHcL8H8ff0QOtXCW7ATPb9eBoDcXOBjwKHpu12QaVw+Z3AFt
nODZhcfF3J3xvZPAb+8kbJIW7LQdU52iJ0cKec+dLj5go7eUjf2Ut7D/7zbqpIV+
FZ/+7lEtvwU34m6A7lDzF84bgeeHmIwM+wlox5iJbyys/SIa+a7fUtPw8GjwQ42A
MkU0wuSAyWGur42zT52BdQZsW+OerGa68jwFGxbDnXgwpfSVylorOKIyHOS5l6JC
5dZ9soThMWPQv9SnKh6ZA0V9oLXZ/X82IUIIBA3Jr0T5VXqVkTkBKKqzozf4WF+H
omJbj5bFmmc/ASV0YNmX/przXMziw+/qFPP7Ar/6xCDgaooLN9KoX0/JQ7ELJKNd
gob0XKTAbjl5cCwngAY9SB6oXUFYMDz3n181l3Xr3HSOaiFUmedy1Rd/wbzhrrVG
wfwlkVuw+4GPLz+9I1tQR7t0Q6NXbnDfwBwpNVDhc8A+2M/k1Rn7G9k/U0tuC2H2
T8kBZ7FEfEeaxXvVTQBQYWBIdR2DpGYT9ae9sb5lWeIkhFABamhNnQLUBQn7wwHn
/v7/xTuIkiKCkzutWQzauPOfcxvNuNe1UR/7IWbnx987z3TFyp12PQNHdewdr6r2
6pKC+zhz2aYwfvHx+L4xGugPI+jS0Dd01cx6R/b03burUmNOggdK/RzeOY0x4NSH
ocVpghag1ozvrcHiNpK3OKnbDc7o4ZlfkSfMzoVKcsZ/+xw+xsMI3s7AcZHi5Wpt
vDLOSFXpXnwnZpDF8sfxC4pUxQcSAXI6p3zQOb4M3VW6qQQWPjt/xIjXadnF9/65
l5k2x6U/ZO/pGw9DKw6WK7E+MlJ+atKaDqwt7VZDTQNhLmS7pRpVdFKVUaZPrrQv
BXHDm6vbaELKizSCbcZXanLpX5LJTO9KLzGzsTSaBcckyDUHcnjlhmpgH7o8U9En
c2NNcv1KDQ0LExgpHreh/q1dYNtYgZBgmCSwRqc5bZebBwnJAZ1ychfULhsGNXOD
GaEPi5XB4Bw2+4zLEL+LtpINGSUeP7NYzU3wlyT0Nk1UeB+PnTzJkUjfYpoGdzG1
37v8GtMpjjXQBNiu39Et9LUCdif8e90vRhkd+mhjW+D9TBeUj2Jbb04iTjhjlewU
tJSubNe3yGu1a8BB2LVWD9oNmsAru2QMvhsOnVE33xh/NoaznngZ89FOGRNSZZLy
wDBuZewB0mueH3ssXIbb9LuhXIkjs+6309+PnPcN2/oA34VKFfEIcMG/Ywcj9ZGO
Ci8sMHp7GLMPZg55Stx+QvvC9tYdllzGqKBF4YclCGQlItBADywaVNFwn52wNz35
ITSBeofTiyXZYXxLySqdY2482V1kYWol7RXVXswCdFS6r/iYDiR7tYeE1ALvJqjK
LTdEnXZCdpLIulhxh7SiaaUpKWuNB5ZP3EcsFsMj0MfzlBLYLolMxC6fRJLOFxSW
iO2zog9PK4qHhJKgoZ5v9sSqMXUZM8+XOd5Zo1oU6GytZnpMcrXy5zZsCOGxiZGa
PUQdyxZmdBnNC25zCrFvRUTkhaxKhbljG5AoXuY1nYKBqdv0jIA8zuVMolQVqYWa
2KuEfdyATfJQ1fh51yNgTCbfpN72GNu0WCKo4+PaGC5lh/23sSYN7f6E07Elhs2R
C7T5HImNd9gtoK/u6s2e+7zneQRY3FSGBYfW2/yk9MOb2OmRSdDJGjgPlUhgK9Kg
5DPVSImGPoxXd0uP2M1Ad5oRgjATOm8AEOxSU1/YI5SauIkx6j2VvOzL/wZHHmtJ
tCtRT9dQnQp+t1t8PKRo24QzEUCYtr7IbI+mSCM6/OPEE/5pSpuIIYC3S4wxvIza
dNnpyPs8sWFcw2gDFfN+V7pgXzRgEb5tMucTsBJydnDB/ZU3unon3NGozuifvJPK
F9fvRSEPhvakfAEYOE1PeM1gTnrTO162ntMEW/N/nnEAY4LM9uxKFPJoROSA/LgK
z8kv7l0AOME5OaVKhc644yhlc9f5Aq2K9Zj7CLccWR7k1vebmXmOIDPrFajH1MrN
k59GtuELvJDbTYpIlOqbXNcBfsE/KA8TmLhMlSGP3Gv5wpRYeg/bfAj9K3OJTvZn
mmOBo4CgLTNQchrEw+tcu9UQwBNRSwpQ+20CbwWefL6pApq/xv+NSAeHiuH6vrBD
G6pQY3iHO+b4GhMtrT3bZ9CdGweiYEuO1lHYynuLOwEAodpwdx34rb9OLw35lK1m
5ejMWnQUqrEITJuujIdOsIojb3jioZVCTwV2Y4IsU7F7rjrrrzEeaT2xSml4XS5/
6NrrcUUbxAPescM5zyZU2IxsbdHljVXRRQQV24hjLpZ7MdUzNJ+JXDDGSUA3Pfjv
jwdzf7PJIm/sa9/EbXpAfvlcEefzqPID0cBwmlpcv+j88xxQcPC5RylBCo67B1hf
eH1ytYYFLW1QCbpOTbJ2X2CpAYpt6ZOBLVIKXijsk9XeFNcHIrmY7yc52PaAsU2R
oIsmLpURVEoU9WfA6yCxaMoinrUUiOsELxFFA7bebUERtcPK2Kguekq4jMwr+CV9
FZxf2Bnk9QQjgMIbzm7kiaaIhFCLGDQn4LkwY7EcguIVXo+02ShShs1c6EO7bBxA
XQ/nduLY5DRxmnENAdu/9TpFnOVdd74XtmCHpm2a/3YhdddZAdwkH1krov9wMSgO
Z/O7TQgoi/D/oecCGJLz+TSoqvJfOzL3jZPPsP3uPonZFhcnHBD7kJym5+7/U2Gf
aJpbANSmL7Gp7AAUBKILHNE/oyl1DDnDqJNYGL8jrCVxL/3jXsa4a+1Y3Z4I0iip
npYYpfCZgku0xPVZhZdHmfiGbeQZIt8bUYnqEnoYqrnZ+RNILUI6BNU4Ib7q30Mp
CV6sdXENJEESzFd3LsEMoTBIBvXNO/PXRSkkVegLpdnfMIOUVeEydsGoJZdNdh0a
tnVheEPgasxa/1wbP2EKH04r7w7+M2Ev1maAEYM9utwc8f08w894UBL86fAneqSp
4pQU4LWTpDYKvHgOaLYBP3xuviQHDpzRrRefVr5a3GtIWUae5aCUzjw6+ZG4YFJa
PUJyl7Pxq9kFVMt2NRyOz5vLJ6wBDWaqK2wGSVxeH4IPs0bwya/G4ITK2MwZjPdE
o5oaQsFX6e21MfQg8WwGix0ESOY8dKDdqSHWn2nMLb1mSldUX6KlxqLEB2Xi1oVk
J8w950JPQ80Kf9evULR8YEB4QhtM9jDXDh1yxvhh10PrtO/LGhoKVOtZlovMGMSK
O06BJEogCLt9rMakHez/HvBmqmg8VnaNIoGpArRH5MCeBtCzJghmPDF4lQqdCQ5v
1A1fWFK2JTTBxQZiBTyFh//uJ2/jrcx0EbJA9b8xZBquHg9yUU/zR+ajB58cfhj/
f2kq+N8FzJ2vDKidNh26cwVdRSK6wZ6AkKCJZ2A6zWrn48ePFuBKZfoqjE0fRDMV
gyzSNS5S3DMCx3VOPmBIx1KNVcdlsvekiMNvnXPPO9LwObOQxDtCOFluu70SXRXD
0zhnJxn3Fjp4hvFXbM+CFomhOEO6jtvZn8nyaFt5FE+SynI1V7ei2dvvPug5vUa5
2Pmp3DKh4Q33cPXmPqRyDnVwV+GZ32smJ89uyv/PSdaWNS5A/a8gqGy4N7/vY7Zi
DF1FNQur9Tyfvzd2WIYgrpt5RP1x7HGm++xuV0d+Zm1hInbVymHpyyT46JFv9nDr
eLQOfxeR6kcLmTCnHrRMgDjIPtVEpQjTB8Sp9LxJNGY/ws/5r2vNCVUNLGibY7yT
ZZGfFVtKkXFFs/qJ7hloVBnkaHeKIGIDzcgHL8p1QUSzs3xsP3PJyF4iHzrSYHS4
rmYkJjibTSn/iDRyuinncpwLo0zjyHR5neTZLSiit22VHd196kWP94kOIi7MhOaJ
OsJU98+t86eXnA9C5aOUx87Q7q3ASdeOLUCOjvEvW2Arg/AAB5ntkOLv+ucm7VIS
53m/KmbD8TJmfnT6wK1o17nfLhUG++9iTjjeQtLop31LQ0aO9gyjlyJScZ86nswO
XdraNxrZKKgjrsMN4wS9RdgFsCCBRtLlyFOZstVFUzyJJFnXtwVgVJAv1PUzRTr9
oShdzyFZutWOmyMuPEip5ntk4DB0b1WYq+B4Rdx3pDbwLfUM2lVy0+Ni8YqBFO7y
ws3ReU2BeSaFLbnTSI9ujq4IX0juuEP1Ts7QetLmvF42HOT8TC5yiPcnMG77cw4O
HpNGfGRmLaLSvC8n4BQr7kBc8QyjFgU8dB1mgiLtJsd/hzqX1+FmePEv0b7tGt9l
L3saeErgOXKdU+ocikWvEqdn2XNn3p8e6hvo0avMvuDQ3qbn8yxHIWQGMPRVL064
bxSe+5/mfZxz5oiPYn4sYUom+6BFUQ0ZJiNHyyL1wdC9My5JlIq7QK6gVaH0BKfa
qunsEGi8WzZHzxLJEHGzFFJ+F+ZyQ7eB7a6B8EEkrFXsP2gZBKmSnsmv0gqIzWF3
rdQEzFsMonv8JIkoQKZyo1jbSTqaswAYqXyXLggjq1/k0e8Ia2cqdQVzeSL3KD/4
TK+7JP8rFSwrJP6/nepMoKz5J3n3/idlabn+sYZDQPOAzlA61qQrete+TbYr/w4b
JZuJ1VWbnTcb04+LO4V4ttWmOvnYLtml6bINRFDccVad5X4Wz8d/sIuGkJvjP6gO
bKyepa0zkcn3FEH52V8nKv5k5Q9KqTm+R/T9ICHqCiqjSSAoTn3IwGnRhzIZvknZ
Sad1g3Aqw6v1uag7ful0HSxuuSyt+AW+VkLrEeK/hP/2VqTf4IihgVJom1DmnnPf
p6+nA9cu3FiGMUagC1dIJsNinOvP0kULdzNQ+K3AEqHPiONAewiqhY1kpx4ht12b
llchmf4r1S1nUX1+Zibbr1+TVpL0j7N17Q67H9Km3WM/eoLtnfPoM8ZDg5tWWsBt
DCoLwOqUxUgmuQYyhSSVycNLu8/5qrTGFldQN794hLuPSAL99evHUoq7xDdkkWfX
hTjp1lgzxH9LAXn5oOM4/bHfh6cT6fJlmjStZGrFZDC5ABzRiPEGFryDBT3WOm4u
TkGtnSo4E3QVboIzGU5HVPoT3OilOXxNUC42TPjJlSGHJd/xKnSMmwJui95fYQJc
Va4MbW/RjJKYYWD3jcy5zvIXu43yjIou5pznaFMCRXo/r0/INdQM14AwQPGs9+Qd
aIh1Yb4zPhbv44TnSPpvnOKVbwxsmMHSxbEbMBEtf9nHjzHt7xBtaafPdIlNWQPJ
5N8tujMISt5GrXyRQtFKIMB1AnEivNsFtGz8sdjUCg/CUmbxJgvzqKCPCOmGEjLE
yBQBWOjhfQkxThfa3ouu+UtBZyKOrfvxlBWBarZyzOclXMgS4jrLfBwlF7uKptBC
MKj1UdSRM19Mz9NFhADZogcXiLFBc4umluogLv273IWrsKaAQTmOGRV8PttZIG8o
Skln0U7fLdflMoFCZGDw/V3BvyrMd+hnNH5mhBMZfmgtlryljC49efNAA8m+V5B1
O6EC155jiHmmjKwnE9X24pbfYqvyGDRuVUp+u8TBwSfUd4MlGxXUnhWjRrQqTy3j
NYcRuqGxw0ZNfmdq5yj8g5R87WhTpB/9PNE096oNlXZW6kcTcql+To0BEao+nssQ
goo/V39AdcRoBSjmKhgScmTGWGwTmPz7pTJgc8JGnGQr8eQiyEcaw6ijtolmMvFl
4ARyismBJJFXtRagrUeNxKJ6ej+d4kx4x18fzmBTPoR16I721J2lL93mEZ09B9yC
3TtC00JCpCNKYIVpAZsRKR9LwxcMxS0IjbJ7UNu3hwqU9FavDKEvHkLC9rgw3nXM
tT1LJcv5Gjh8IV0nq4Mj2ruqscqsQDJMXtnCwh6A9i/BoIP+Nn0F6DxZLcb199M2
GLUs3NgqSkGGAScyQ/Dv1Ztd3OntIxLR2A3BTbxLMW3Pifs+d5rkyKfMd85sNApJ
jgfcRfZFRyT26yI2aF73YLE3ZJWqtVtXHUEihcSpSE66VeJj6ePKZdcezQXVK6S1
1sFgS59OGk9tapVdajCtr/0PJGLQLCraGFXJt5+G0LRG+DNs8MtgYO1ujzJdfMBi
vW/GTdE9y+feWR9FXBjcaoBjFhuxHJLh9wI+0dG1cbuycYDCC2jqOKofRVY8dFDG
rYMFxo4Jf332heLEfVfkKr1hLchY7cA9vy0VpeVG9U/tgTjwOqQ/QQJqp9QRMlDR
6EB3PSUNglJQ0hjc4iRrAWI4YHp+PDP0vyHBJPo0E6oRztKPC1nWoNm02mzETaPA
cKq77K16wuevSkMficS9s03WyJMYoBnoV0UPAFU42mAO/1OtX9E0wFrqEDSubVCQ
cQ9Z94yLhY1L/eHnAlIgOAcyMqpDA1xvCfmK4y2jeZlP5BNeZ1DdC0eRhgOEqY7F
yzZMioOUfh4YZbSGscfDylQxEGUlM71MyQd3CwG+NORm6wKZZ9o+iVy+cjExXUxh
ow5lFNOTAjJX7zZEX+1UWCFHCXnxQBfp7GwDDgZS2JZRmGWyKXNveO0Ff7sMUrlY
/hv7LMlwbZwws23vux8GeBjO5ulfIUZiiBlssNuP7s3AOOfZQsGpePTBFSDMvn46
sAkR1h/9Ov9j7gXzhqa1JGWg9uXX05ztPZtw+7Qgp7AcyLTAoeXphbeDrRCthRWL
C6DJgOyt0p9ep4om/ci3MU+o8A8FJWK/XNVBb2wVw5yEtF9WaUc0xgOCv8fmbB8f
vzdFVGl7lU7Ih0buvS5WigEz84pK9NAwogJrx9KNyxM4J6B3pav6hqii9ETcWoqq
UDoEOqd4ZYs17wYif2/pG06f9mzWaiUGzt3rAOvTBK+tAqUmfo8KOy2a2q3QCE/3
ZPVWQDGzobyEPdD8xp/yyyrQqQkPZ5XCpM7pvSvPLzwLnddhaurNkinkXjfdxOO9
oy+JCGdGgpN0TWrMnCQu8pDByEky6PEyt71eNJUjqdZSRepb0ueL+7VcYnie+4+v
pT0NXBPKy1CgCQWSf6GOyVLGSp/bcmWAmcZSycLGoHSGbaRqD9jzOCiDJlL23n7N
SzLENlWbLKjix3sal2aLH9+5OgQe/2OFMZfj8seMVxW+gGyE5AebZQq/HyiVFK1p
ic6gNxtRYUSysPfZaR9y9RA0zm//Up4RV/Jqkmi92TChFDYAYvzEebeHBfjCPrKL
4ZHvLpEpI05QmVx6aJFwNu4NBEIlXKIMivkughhzZEF04xrAfKMghHI6c1/DcQDD
Z4aKYsB/sD0NmGNrbissThvEKzZQfLT3T0rR4WzpiHM+rnW+IEJnBsyf7SypfOtk
Pn2jmIEV5etAvC37PRoYq2IrwTwU6QHzVA4h+zxIK+CPRWNjF1DCrNFr6XczED0T
NhU01NYMQ5xiKV0Sm51jRjC53dVKnrE+5Eb0k/zz8uHxnBnAPw6glk2nBUQPIGYl
oiGeXfqqso5QDCNlTnCZniR+vdUCRnHVj5BWlslsr024tmfnJNQ3VGOKCbyfe8Xe
KX5cdpoq9jqWIkL8cvBki7u5ZUuDQR58c9dQdoYAUcGQ5WV+g/hP9CARGo5qzHZB
9fHfVVO9yxmMhoqKUhCRCXNEXx166sHa3rWHX/fVSHIm0Bibs0F4x3ph7M6xhYh8
VfuE3s4yZLBnhfPjMWGtt1SiwP/PAR2NJwQWBsv2unFq4/6MsJkz3sdcZ4/cQAI6
ukuk78M03Hs31IA3xCiNPHzUPZIE7ZAMa/Yn/W1UOTlJuhe5QeATww+7o/jUUXFM
ams/mIpd68QRyQVWvNQ/Jq1h/NvQzZMY1UWBL/YCTSDwSy65OUjuQTEiHH5yYppx
86JUltGHtdTm12XQnAltDk7hDZNR5dvmDlOenUnvZcqsqmbUbbY+bpMjmyQEkKdj
EV5/EXlcCQBtaRZYOJgQT1WI5xyJ82523B0gn8RscsntrkgcTED19If2NRhzq6n1
lzlV6NnQbm4Qp41cyHS6Q5epzTovDhi8kLvCUecheEtIbX+XVhz0QMyjifBrVTBe
AoqmK26MyxBokEVgBcGEAteHDdNXaY1GVYj93zN3y4RdMwM9obsXDXjMWc9uhVkY
VRREe09XV4haM60H5coCMxpzRuRrnR3pFXgR08n3gqFyiR7ejZzruWDFPkn8lkBW
sg70J+3MLuO63Wa/6L3RLB+iQ5gIaDB65STjk2IWXHjboMjEzcjIWpImikOdk54v
LFJiKvHCZ3ylEGT2e7P0leJ8DYbbK9XG0SOSwk5ntzhTuTm4dAD7T2ev+j/0V7Ef
Ofjy9WYPLi8ACkCvnbhCzwyJMa5irQ0A/UwAjSJTJfY8aNJU3Et00PcGvHrIQe9A
/kwM0QQJR9n+EjlRMg1B9X7fGGGC/w3LPwVLfDZUtR5X/3ZSdSgQfp5fwaPwrzk4
1/2wl9Pk7ha4kSl2w4us/0vkzO4s1RjngVPmPqEgA9d3R1q9K1wwIqgjpHH7q57q
nBsqgRDUKtJKAmS1N+nhLyGaTGCyW3FSU8JsKbNUN8kG3P2B3o85CA++Od8HbgTQ
0OJVbvpEOZ4imm83uiW5m179wewWLYwIDNsa0xbngI7WXY7PYMBH8SwFucpcYhwK
j0slsgUcDU1WE2fAUJVsFSJfXdTGBapAkOFjtURGx+Jep6J0q5boBGXuy6IMA6kL
PbhCUS2zWMTn6JqjV2fFT2F9r8tDBsVVtPfTz4yHn/OTY/btLQsqhvhfre+SQ97M
XQqnw4UQyMIsjOGT9v1xW+5kTVP+O011ChDV3rYiDeX0uJaxbwIgLIFfplz2TUVD
Y360X5nEMJboGroG8gCsHqomlIp2QkwdYs9nLML3U1iGxkWQVk0/6ij1+EWF5CVw
wgTbts655X0oZkkk3HzdobJsn0YwXMUXmNVf2Lu2K2n+dCfD7ozKO3O4Pl/yhyry
hAVt5bfLEsJRfEOjPGInXqZzbBc6jYKg/te9GWRSMyM9s6GObj1ze7+5U89i3pqj
IljRQTlZazHlWFcq2FxNBDNhCpbDzzTNJFtcVJrokRVaRxXXekRmYh/fD6EXEvmB
1L9O/h2Fbn8J4RBoTT1EzO3ra1Re20K+uM3Su8RxnkgBCRds1eHOhBvi3xFQWnJ+
R3DbqXMA40CHPnq5nPCmw55wYAyAcqnOlfcmEKluQT11+09e4FuLhTDEwN03srRJ
JKBvpxNFBzi4G/15+bk9obY3zvp5L3NSyrDWr8QDf9WmWlpdOOuA0f4n7qb1279P
a2fRjmaJWr0zJrYrOXYfT1v/D0pGzYMjurXtsPUoHRu7LcHz+z6GccDyUq1L9/S/
IyRZl/HdvpoBgI2fA74cW7WZHdnlTwwWDJPDERStvXxG9Lcqa/z8i/3yXSUP0MDD
Gvbh6p5fJ3Ojma3Pv5CPDGqOWtLBceRXLQnMIG5LHpIG22P1H0Dzwk+pzj53pAzW
8Q3A0e+gJn2H9M+5nSArOnFJbBecdsVsX6865ju+adEaH7DztGv5nToRj/b4zho9
5RuPsp6url8bnacgQ8Mw1JFDDtgNlEE0Ne7SKEUtuazKDtaAriM7N4G58xvG4skK
olEEz+81d/bzr0U9LnrwZOwaAmzlrel8jJ6JwLzy1FGEmT2fondGqPV5H1BQ8wVl
RVZ2voGF9d5ba/2QrKyxstku5BAXXAnEmqhatEVVVcYiFLdlT7mXr7LqWHHDPq51
26weK1wKuUjiNrD8FYlcOXndaq2bvGwHW8RyYQ2//OillU9PMHT19/avlUzn5iL6
7LoFJ6b0+W38xHjZ6QpbIf9FhjaEASg3OZttYI2JvFcNoBmYmZJsPkLtzwna3dWh
QBejJ4TU97R0CttRAFbH+AdveVjeGabf4fDQxc6StIScRMIvP8kR/R8zvHxxsFNb
t1OYYDKYjivxmnD28ks8qh6EyoqsIj6HDifrEvMY6DDj/IxAXSEj35PDH4D5GYbd
sAL4Xf315DbJkReCDIG6d5/7xBkN6gGpmr3RWQx/4VnHWz+qdxsKWogF7xnyoWpw
MPjKd0gzm6b39YGtzQFLdnZefjCpQ21B4lVcLQNadiX6fdqWWEdolMOYzULaXxE1
PEO1ijeXDD+ozaaeKPo1dh7KhvC4HSdqPxYdD3HhbQC/7oiWLgGFeElasDAZo0vE
l3XkADNJtBI2j2ozsDH3lJP74X0FRS9YHV+GHP5mYi2ZxtyxZt2jpgox7RUNIAdB
ocnKQlTYNi8IU+PuzbYCBW9SkE1I17IgRKXrnTfo5k7HyA66IeNgDJQWqdfRVRaS
uDC/thvCAQWBTtTwPYMlFE8cv1UkU12Ag8UgogEwsjjk+Gk7iOGVcpB+wQ2ELG2x
7M2f0IU8+f35eB0/afzHjTCBXatYsyqRQ3wjdu+QPz0eKAEDk3XPnlWX9tbF2CYC
WJEkfFAep8uREJjGm2bAsnycjnSqUR7g8w9c24Qm6SeGDlVvGzmOrLZBuHt9pSQ0
xHbygX+hELY+9jRdGWUpMVJ4ARgB5zEbSCfWKG8cOeR3cs6YLBn5i/q4WJq2EZJK
Tt576PJgKSgs7j3NDD60nyTyIpvB4k7AA5wD2dvaJXvJs64vFrzUhG4zBEbsR6ZT
7+veN/eXXs6kLgO3BvtxZWFQwq0ZfeXWJckC2nxA7TaDz035aK5qOwHQk0elz3jW
Ax94nX71vIHmJhfJQgKBi6CxR8EJYVlQiG06oZfDNum58La8xFpeceNp0Wljt02z
R0FlAOwdPLNL40WJBzohloOXplT4CYZFfDp88xeku3EiRXHXT725+E1Kkpq1wbU+
nQYKb8NMM9cKK5OtJwQge0Drz/fjfzu7SH3/iFWUnapR8/4cNnmFWqqRn7l6echD
8WLa2K8n3s5iqG22szfjjVToSFN+hJmbYnWI1FQXlwHjntTtizc7LA+qmw8XtcNN
EJeTp7Orhua4r0xbNa8NPeAnaxy8AW8PzP6gnXBrGSfwuoLoh/FX3r9UbVdliAW4
Q2t+0xKu2BbnJrXT6P/jNE4JiBO0pJsXkJw8gFWRpVmlO7g5YMipEbTSi7Ct9zbm
x6zfrq48yHyXLRpgdiEyefEGI2Xid8qBNzM8iu25+JYXY/S6C0Ikbx0EZlEbvlT4
4TGACkZhvcoqymON865Mo5wIq/9aPTCEQNmU2zCzp/QygsGlVQ03NncVAJzJCTyT
ccLwX7t4TEbeDfFBYlpLePa7S5l3v6vncMUID6puLRo5RSFzTZv7ofuc9cZ1c24A
nTJfg5O2hvwJTh1r7GtyTAiylfQ/w2LuVfqYxQXyGzGzRNZxR/tEK6T3HGs4DUr+
0LUDmZvpinQqZKfAgF9ugaZgBXELeudq/8ZPUj7HlaLek0NEjv3alKXEbmWxlTrV
XCBcAPgdyxLRrboZRL0kJSE5IjQITImUYBqKOvzlG0Vv74kY1SOJJ3J4R6zD45b5
14cSy/dEH5flud01YaSMNXR6a6BFhfJLZbE5p79a35txxLakRYXXMvWlr7qO59UN
DpU5GsMAwVz3GmyYEkBRk2jW61oo1/WbAEdVGYMY9mRXXxXUiw/JruYt09d4eE0C
B7YGkn2AOKFcH/PncUuyuK7QMAiJ2QG7F1E//hxIb5VxigkkOo/7OUrzQhFOsCj1
A+qJu/CQGq7xc3LnccRJWmUZA2ezgF+FJWVfv6TMUCYF4q5Y2yrgIQ0ZXFn6y3pu
fP62pMffygVjfbMD4cN2OvPe5kCU40RMmDGpNR936InJfXghrDTO6km96e2MhEWF
hVe0+AYc4/riJivac+PJIxQ8SUpWY2jOnzLJ7Nn0Kg0mNgn/qpOoXuGQNX35zR48
hlxfLfLRIADBvXI2XDDDnb8V6a0+mGKlpgExJXaa4In9bT1Mdmp010mnWazH6SSF
DCQTDsydckLEiSvoMawUMt+0Kzp/GPkZWreRrQ0bAigGCJNVe+UU6q+lx93pMNsc
0NlS63/umuaBgMkJtEfFPInVuKp2NtBIVMY4s24tdE/CotjIq0POqIS8NjL+bXDB
8TdRKL3JEXUIMaMAksf5RuY3PLRHz9dw2by2yQDGik1+LrTy4Bj8z4nWIiHHKelq
f+ssQ5ED2C3eK+s4WCt9mf3b9+kQIwn1QhTnDSNL30Wx6gsUSDrAfV+pONTwBSa6
DSkAgfIf/WnBgByQ9DxBK1PN9ZtoS89IOuGcXS+AlSbbi5wHdvAaZs+5648ZZMH1
9uSZNTz/ySqr2jxoH7QheX2mpLAOYWtW3wpRDm1DyHK+JVvk2fbU85qqaf/U1yhC
R2qFXz7G5JKaWYrw1MCXC6SqYGgakXx149Q64vaJeFyw7YDJ87E9INEF3QGkxgTC
fYjVO+sVQeeHElwoHSTr0GuTEVT2Bv2UI4T9OnGHtQAhDCiQxPrUlnYfIUVw7mlr
EVktnAO4OWMhRmOLxGlW3c+W7Ce3uTI+hoAmpGJC/SbPOmkRegLQ38o+w7R+ocMY
0UNKBzRjBegbXoHrwmUBNv7blmw4/LWKrmqeKg1pHPQUiYygouaCRzqNcXyjF0vS
GBLEstcui6JymaOIu4xXNjy+qk94KlaDRuMueY7iwFAcmN6OVxu4w0SNLxum6DjU
lEkkyv+iMkVugpeKLOx1feYrc//VkzPSbkSJBKY76tEpzvBpjubMrGXVT6CPt3TH
pmb9Buwmzu9psNa97yO6gzGhAkuDdgvjzIF+hZeaD0tLanve7Tk8g/DqR8njaj5o
O3rnc8TnDRdX/L2GVh122sG2pLpDCmFb+xxn3ksjxQ/zV1iV0YS1FGD4VT+8U33S
PxeyqhrA8ZIhZzX7bhELKMOOiQGh+eSxjxVy9dETFwcD6OUkh50BI2ZAI3k9gxMz
hJGh4poxUbj2gXFwV7o8nV0hNWC/7irs5HrwaZrCtliKLeLjx7G+s+EihmuG+hFN
yYZFaxH1qoQYMhLQexxnxZY6IadLkhQSF/YNrX9cN82JvfyO1oUZlNRR4Wy9E/jL
W0uhCf6hMalgkQIS6fpNRxpxq2/3Qlp2LavGZu214iHKEx2zwVubqMz+OxfASzwR
V/2Z5K5szyD5IFOws3o8gXPjoXULwZAYwRwMq0jURiBajaxayGHRnFQHpE0XXSBV
ExbgQPw6UomZn2JXQQ/XANFl3mOF3XwussYLVMKQ2DLjPol5Q/sbbWnu7GfMCOeL
Nd+op+D6RObg4IiqzR10hb+ZGtC827+O3ZT3qgtbKQAQbRj4d/PJxvAoIouc9szt
iAqugqhauwCrmZb9VSOWaX9Ukq3J6mi7kEruowzkQzEy+sCEKu26MZzCtC3cvKz+
mG1M8399oSKwNvqVQs0yKyhpUBm3UjUxeDUpChBJN0pCo3fMPQMS192le9aQHOG+
HFsORdK+MpSrBdMHv5qI5vJXa7bPSWeQOlnK8Nk8SKY3M4V/xQPu0k5tHndJSska
g0yVIwEUO/KU8C1XC5PHmBxYmyPPgfphf2amsH7EmhDZYwa89mRXXUQc3gcfarB/
eG5nnH8ydbJYPq/t0+LXKkK2RrM5ZQGGgTaDjR0aPJGw/XsLqG7nimdbZiFNf9Ai
7l6QrS3JN0Lx+Zb7YwDIjzm2BOFnxM7xAVO0hOei+2lvNpcliMSoAzEreR9B97c5
6+bOMgYJuYKevHCm9S8qAJ8KZzzUL3IGCWTRLZQBGXz9sPyU+JpDWOvFgtG98bl+
J/E9OD6pPifpjdR0zYz8XPCyDMtuY+S4se2nDfRSIeCY79XsULRfW5yplyESsfWJ
F32vzYGNRl3Xt61ak8OQoXdlc/2VwTQmgUWXAamKnf0MTt0SMmHXTkxrZJK7Rh7y
YZQ0Joa8SW8md7OxGjxA4mUqx/9QPkf2vpnoxpR6xnHx5Fqf6ONJ4d24D7mXtjrO
sy4DodAcN0S0EZO2qbOuUZOrNgWzsqE25hRidyN/7G22J+QgKBaMdN0hSxOGTmwR
03vTWcxUgLc2fEzEsq3mUYhPPMM0rwaE9IsrsrDmD0bg9B5z3X5S+PeihPE51g0H
ftP2H8QjQuLKMeQE1DdY850EvWZslfaHKHGfZ6OUrvMOi+N2kTXxriTY9jqR8iDj
3bIO5qY+1WR9WcHbo8m6NMec3hdIjET1l4WWIiKu0mh1QEQUMWJN8sa+iVoq5fma
Qo+He9BzYYEfRVFdy0eUKjo9YYPkqbsc3Bop8xANht+YsJgHkmsGjPm54Qa+tCAx
jDfcmZq9t7Zkk5SRVPhUUJqG/S2l/Ofn9wBZsZpA0pTyuWqtWlRu2lpEOoaark4p
nmY0OFBkAVuwgd4LKjK4Yx9xAaoyO8as3DUX+7N3TLL0xiaseFQeIT9CAB0VnG0o
Fz9wgUmf/FwwJUgsf08fyi3Is5ZvHodwBiCDs3KKZrHeKig0KJSpB36741GgLshr
Wqgm4Xy+ezITYT0lqe+slOK99s3hYaW3W/C9i860lN2PWCvX0+4IeQncLh0pwmYJ
VptoNAWOffJpIoJD5MPiljW1DEWmgPE9UQ8t8C21g7gA8LMvaZm7SCK/FRnx4lOj
gVMlt0n2F4/wyXjmF21Qkubbp7I1iCfFmsnCsVYhndBjrG3jBRhPMyCrFqvbUndh
8tmLWuEWRa59lWoFiKt0JPsJBr4VrUnXKJrY0wMq73vu29N8j0IavsKFe3tKXGwn
f15lqXCfVnnnnmcDjLXasCpDF268MHT3atFzCiyfrE7OpLBjpvBrEIikHBG+8ogu
w4rxs8SPIJIUmDplio6sK+OPpag56o0AZ9CQZuRaKJWjI+az38UhiPAY3lE+n/Ce
tmXAz0vJWV9S8GthI7T39ZBNgcjyhc3mIvdYGXt/fNfOcTgfYmGN89Qfu/oSW3Ii
3HD+PlQ0qXkmaTYk0n+QMv4OvzTPKGuqWpBhU/e2zNcFN/XLbrmW8YlP9vB3HyK7
9aJnXv634uIg3HLB4qlCQhdLDkJBdKAOsDkTgUJ1DIOudH3U0uOI5+slWEwThNeZ
dxk9rvOJAPkkOwPZHRkvQD789mIk91Oj2YwaPBWCcPhS0+ugDZzR8pBQpopSwh4j
79pidJgPrgcYP2miyPHop+Iriu/NVBcv7LItZS24DkY35dSmIfWAOvT2IAG8XQeB
z4VeiuiMj1iLuuYf2tDdonYHB8i+DT7vqHc1KDdr4qxIOZFqieGuK9plJ8YRYnZH
Z+8DBd0dXZqLruV+1uL1+oGEtaPRTXWJtRMsFNFvELFEbd6A3HsaOq3f3rFJxxis
6qTonNdUgE44NCdx+ExqV8oXc7wuVOJPy7JFDgMrsTfIM7ldaYAymyams1B9ZbkD
gRWZYRO6LtT8eCOLw/PEk32LquSBtZA5Hq0kFj8/DSdkhtjB5XgbL35qmF9aPHSd
CXYGw0ipuCBlQ/TwNfTy6iOB5ibTz6E5c/tFVMErBEgGZIdLA3P9flhqu2pJd0cP
km1/pnDTLSwFF1WtPwX0ml/aE3GvEhiZf5ichw7K6A2CC72NCKW45Xw54AUi64f1
jd3Hcj6fYvHNYKXyfFowArN1zxYmd1Vwg8oG/GRKI5NUcDP1LZup7HmE8DIEw3Gj
h9fNqEn6BRt4BEd7hTEJyX4SSvuhKmjS33DmoSFGX8n5bE2sU0mNxUfMf1PcW6lT
wVQcjDWm4rQLQUziZ7gIbDrP04SAUZET1F0L/OSNAIaVWgfR4UHakVizo5wbZMQU
IfBiesLr/OktqTLesdvxy6nQbo2LRRH1hLziwnlFudfe4N9Lxy0y5kDNM5ZNSaOr
vw2ahYiWywSS2iS2dO/LNpULLDTBCiVUkoyMSlmdPwNSf2cSNKaSAvib9I3O96wn
Yhib40uH4G+5IGPpJTwaD13Rp4WtXMHZzGzMWHFhx1TZuaag0TgoOmcPd3eSbXiJ
zFdLs5JIlIRebPciI1s1gePuX+wl2V0/0p1FATkktPfILX8/QovRIbHihyRmFEgT
eK+dHHh42c2nysjK5cqztEKQBF27B3g/15+O4/MMTKl7Ch62//AmQkOePzy44OTI
JVKI1YsDUQaLoan4u2jrEZ72s8ARj/JInWuULqfsnKPQy6v4YGwFmre7FLCO+sDT
DBgO7mqLsT+4Zk3HNYkSkZ9HdQwfSJGaaNS3lgTaL/lugOKFFrGSER4Jq2uTJO8K
vnhhWV4+Given3ZVLE4QW/FJFJUr3Bp/XrQW8f4RtaIQH/kC7MeBnQfwzD5/F3Ew
siAASFBHDXyVMqriV1j+xdZ9OYx4qrQr58eLNeL0yffX/tbJ0ZSUDTiTHDrqeGQO
DWTbSFhv7M5dlx1dHhVgOSohPlGpzVwPRcm6XN/R+1lkucIi6/ruwAkZpea4le0i
vaHzcinWAHLRUkV3XtOy1dRpYcdyxIcApj6FbiMNRWWqbxxzPRNqHpEmsa/+9dPY
uAncNMaydqgVwM3q4muDspwE3MY/FkXJ6A8JHmbRqAbuOHOQCyXHK4KDF8BBMpym
l0/u3CstdUxZ9G6wgMtevMUGZlyeu/qdiguLtxmnUl32Vy2nBBXu+YgYq5VzhJo3
qePyjCBTJvqIDWmmJxGGAfdoU8E6Dwh4Oeo1c2rQfk9C0HcuIY9/6Mq4sEFFfbvq
9srRcsTfvakxYYG0GowBGzJqf9CXG/H6FmRi52/E3lAVjC0tWez1FqJIQ/L5mAYi
i5laV+oc1WQEm8oxzaex9i2ww53xP1+HjgRYAQAniv5w/Aqq5WSRoIF8ujqNoqSy
jfbuE/W4Mh357lQ1wLlFwZ00yMpopIFNnuCnlHTm8V4cCmDgI6zZK2830Y9sXFn1
IfXG3gyeDjB7ir6Hfv0bjcXT9TCQqopSHFye6VezVYDqZ+79pqvtNZvbS0QZYgpd
D+ujYzGBhsmbz+zz4Bour//k7hr6RedkiSqKYdxowuW2nN34+FiVs5PJC1cGURDP
4pJoPSkG845e+CTTzo4yQi+wtNS5al55FwAUVIC4TkegfzDUhvLi2g3PNG3vpM3d
iFkoAo5hQfU0VwkvzdU65IjCYosG9w6ZQaKkwCd8B/CJ32ryE3yGTzRcnO1co3fk
1qk2YtxqI2Npgp8aBeQgjcYYPupYzzOI+kC/EH4nnyqWgBicLjX53ImAGOdvLc8j
ACAeGNKRa/LgOxAjo4kB/ooLDhke4njVOitemihPm6GSZnGe61YWlwxUK/xUtMVw
NU6nuZyVy3V9TwRqTQK7bmXeFdXq+O8iMO6i2XenYax3iJXPY3dwv281DP535ks4
OA+ivzhDtC9ZHyfft/r6sWD604bLeuqJgV+69wTsHRA6ieXXOm9upibq6O5Jn4rJ
sBeRdvMecWHxK0pFRYAJaci6eL0FbZI0RJcBlSdFECPL3gP3pPB4GE0LRiYqbqFS
8DztbX/jPY/sk8RLMlUtfzECLG6u6WfXne7sKxiTVOokNGgvCe5WUtOD3+yPR0nq
FfBO1jVE0HU00/wpJKS1E/VM6w1qD13LPVXgJ/hLhtdap4lWtNaaMCTM2sD9IuQV
kRnv3gzuDIfc4SxbBEe5E0DeGIZkg0YOHvNv9y3MbBkn5sYAWtvAkCj9UsDqnmcZ
HMZTy7nY88yJ61xZHuvFUWVHhMbKOIgjGycmo5SGtPjfKk5vj791GKERBlzcW9ul
td/CzSlJITB0uPmPdez3J5le5kJK8qhLqNVJW0IbMSlGQ5fV80LEv3/L1jhQFW8Z
+iz/9ox5BfQl8m9xB8IMMhYBi9u9lnwit5HaEvviVSnVMwgZrt4wDcnexrl814yu
Kutb2raZlDmowHoDjC5GX/vfk0RrC5Kailizb3FYp+4eua+CAKhlvrRx01GitrCj
DFDUbia54u0JIMUtpB1kbZXzURwZNrz03ittQzGRUbcNc5C4s7ycdXd9843TA5Ib
e85szbv0wGnCvoWkSChf+qILr5Rc+sRZ96Bk9o6Ehio+QHGy2EU6p/852mY5PTW4
eNzZ4xo4qTwCnnWskvlp2fyZFKa8uLN2ksn/5xTQcjnGPAhf8lfggUZz1GRwo7DA
nORuZ0ggHM+jzQCp8N8PJOazBdqMshAiFsLePSGme6uwnAF0UFSRlAR/BH08fb9x
aJHHeK7++PLQgnDtYHzB/+FCkP4L/0VdqaVfESY5pt+1O9XWXNa+w7Z18ShSpdeb
e8welbtOpi4nJD/Op7JiJOp315PfvkXw5P5xwQTD7ZCi83Yg77lQ4xSKMENXvi9H
bOAPYWjhADoYW5HnR91sXkZ1oSmdBDgArQSRLGX5p6gF8Wg2XnHmuN2NW+pJy/2d
Xv+qwPJC+lzI5SCAo08sdKcX1z30ScHruveWy3jOCkCBJTFJHNhLJRkdIjvCxsjt
0KcjD0lCIl/vzIqOREatGyg4tJuWx+b1puxbRTaAj83ReQJSkCuPJe/mvvk9Zx/D
s4Tvz2l1bDz+cQR/f1x7Q3uNQmWGgU6XlqYsamEcTuxr1/ikcx44jAvPnwpykbL+
VTA6dO8B1PMCUT7z+1F1b2iOP+XWu1LS5Xh9jrrmuoeCIc5mF1vPfHybIYO+4h4i
QR7cuUrUQTqCuKOXCK6dm/Xm4E0cavWNmwN5ow8UEvj0moGk0bnFTLgKpFVdtmrP
VkutTpBhxKufpEeUT0rngBod+AtHUoZE3D+Bnd3VKDrPw43jNens/hlUit4Q7dJU
9Fn1btwL71zCQDKqclrCuwD25iKSck7N5YnmMzIpPQdvowcj7wNnddoF6ys/Qsyq
UUYgreiKe19zq/f7XGLs1JlfKcMc3grWrL0SGltQ70myuBQBwkpK7sgA9HsqlSxE
ft3aw74QsSv0/k4JFdiFeoEiUZOUvAk7l+HGHCOXDRoBK6lifHoJug5dGzOijzx/
oaAT2ABcWe9jwOrtlU9rk1ndUyefEGawW0QjM4dw8TM5ZffutnMM7o7JlJxtqe5O
46Od7zSz0RuMCiH5jhNFkxX+sQUmGHUacW2M4KCOlloAuCuuHt7qfNl216CpG3+9
0GUVtVcEBPqMhe+t5Edw0sy8Of/XPClR0hlW9W7MtBVY81Fl5dSJsUq2XwZ2Nw2c
0IxxlObRWtAquuy/X+J0mFZLAaRqEwPlhpSWph+2Be3Auot063Pqkvv+FVi7m1+h
B6z8ektFD6no+Pr9eaG2Fu4RSQymZUJSGnBwi/Cuu0rjt4nFSjyqbZN9LaIy3aot
Rb7jZwAB8byWu8+JbFFwZX/42FlQl9K3qkwiS26OuzpaFgFiq81/Pe2gRhCPj6Hy
uj8jeyHJmk11bujluZIjXNc8goX4Nyfb/TOpP/aA+sW4IM/FHZNmKT5JK4gYGjRL
MK3SCMgpEyvaJ0JrdquuMIM8QrhUHbmw3zS/or1kzrSQ+RQoztRCFaadWR3I70Fy
1JEOc+PLHDgi3K6LnUGXlvkOyRFiax99VNBjkSr95ddky2R2iIydXIg51sztQKVM
LNdXJY6bRWugBjFXEHZxyqZ5wwCF1tKFhbHZjvstw8/+Pd6N5Cz5b4H200p874jT
JH5ajXc6zDgmVzEee1yGt+gsTwOpkgspmlAE8BwDvq9ucQBZBiobRoGormEvbzzX
nAqKKu0dKvZWhIGkbkQL7qK7208wlz/hlnl2DdYOHr6KO4egZkmBE2p2VVdTPJjA
lkuEcscR1tz8UPPpqQ6C5DdCllHQvJQXcpMVEIldp2IJyDEyfv0LZXjmBZyNHog8
vyP+M2q92m6P31Q3l7KouidrxhSJgn2/THwcsjgI05aXpFiHQJeIc2vq1tJhpzGU
GchaiwaxG64RgNmVLVA5/jorRdbYGNVpF4I1MBroHL92fE5dJQUI8i67EQcWHfCO
p9pWjdV/OaXk4SvrpdecpUl3ARALfGBoNI2coAC7r/5acs1J2U/guLLi283xG4Bt
Y8NCjjifknOlkGoIeXlCLSlsrsYHPxQkrzFV5PIqKhyIo7J/koV01eCy4Nyv9Paj
G5vyRSWGK5kqrnBOFXqTAhqvLHc92g0M+RYmA+xG4UsIogosvbsirXywBsjhO1D8
Xq1hYsGkoRRRtg2s7LOQCjyTmitw0jFCzz0r94+tElNlQrGpa0XgAJHywK9mDDue
WBHnpjXw4uUn73LIfYX0JAyFy9GdzkTNES4HyZ7O+Ec4rTRu/WJRgp6t6pbezHqm
pKgsnLnCr7CswUelQxBww5J9ySR8PYanfGFHxZgPszX6TrB1TpVBJhcKAUAE/1th
iaWQHb1L67weAi82fkz0fA8EKluqExNdlwgLA9yH0orLXamEhKFqp9gr6ETwlMI3
1Ab8HmV6PlnRRDP1afNVH2ct03riIjchRz+p34gOxj4tNIcIj921mOd7VEQYmMcJ
RHfccpyYPdIBKbSOEqbcqoa7XfZ0XLeGhvTcTAG81oiX63B/GbbENKax7QDks0yF
i3nYCKKtI4UMxwq/3YMAZLqPcNqqFfv7CFxPGz21hg+MChMtfXp2TTHbuRS/z/hr
uWI1EuadHjBLV4JUDRbmP15Ww78Xp7AYnnNJlmArj9yojGHadQAVexSlzi4hDs15
/+3FyefnFpeA/Ck0xNlO104L7bMv3PG1THrBTjQqY3m871D1qaN9NYdiLe0HWRJj
z26uR1pgYJEyb40QbtkOHgvyENFti+JE//bJZinfDMFiXBLvIWclStxk8NrY76G+
1eEDqIgB11ObRDvtJEol3T452I6kXxzkBRqyAf1iSRQu4Mi9OydyucXeJQJo6Y8h
rEa6IvWktg2JKxMkQ11+oE2MqVpLa/nkKMC2o7s7NRQN6FywbdVSubVX0CKswuq6
RTXT/yRAtjedoLKqS+ZmvbKsTgJeZs90iLuMX6EWKzIN/FLp1uLiB75Zr/SDNKVm
8l5U5t/cErbFDXBnYN+8HLd0RKveMW3i39RqyKmJ7DQ2rO02xRWxjgAifzuQuaTE
mlAX07hdLgFQsBFLrwEAGRR8ccYyvFHVSAmgHOZ9oewnSz0x9MyURl+kphWVxGzp
rKoA1f5FlHfFO1Akdh1dfO8EPL527Yze5spZO1nH+5gEaD4Fg7c1E+LT5pKpqUhZ
bZ9q/Q4E/WaJZQY+tQX29/ZD5sAitUcnsOwZLoiENSSmfKU18mHDzfRDTFlQDgHJ
434T6f0wnHngHadjnxxWRsugA5cELVfKbeXA6mTvPNDB+quTkZaCvaXNprWVSak+
57OQONJXt8HwxwkXGEOVTr2AkWiQ6MI/LfisKN5xPWeLlI+YFXTkLhMJw2Htxouy
8vhdZOJW3OiZ4+MXPOhLjxgdkbBGrVu01A1i31+OZ11tPDT8dzGyU05jQLEZd6td
zvjeb1eMf70p6fipQj5kiZtux0Bzhqdp18kGyErKeXi/DB6BEXIHD6HyEce6oqG3
yO33rwppajsDfsgQxkzm7nWxuqAdyG8KDEZW29nhaMDEyuE6zg+raXDEU5ixKWI9
mUszO9Wr3M/okwcX2QiH5C6J2yqisbZJlN2zXivrPMD8Vq6MjEiOAN/Ka3ThY4Wl
j/fHAHyRuGqS6LqbwF3/6MVTopFQwrZQfmf9FdHTwjuGZqRN+Q/P7lh6hny8WB6J
SAzeiIPLBFK1thOLXPXdFKHOjoyzPH58BZb5RswHlqUtiOkrOAAbUABnRynSfOif
tsczYzZ0sbt/1WfxTEPtv/PK/IdhGc+peaswPjDZykKVn0aQaljkEK8ffZIEmAcB
vxHzRxsV9JMbhFcYU52Nj04gBzuxqLBYG+Eu2WKoXcQXqcHZMCHpoUng4Gg6APrn
aXCtNZjaKYCfnBrmRL6tUKx3B5NfiMCdpkuAVf/HCNKNzcxWdnAYqQThpBxe1lbk
037q3tcJR/HEaUpbp8NLO3YgOtFGgzj0OfzOSd+XyjqxZ978myje2APVTFX5CIY5
95BwaLwVQiChr5uWlk0eVN1TrClQU9ZADzuuR1T6IXI8pV0V7y76cTTxqDe8Vzo8
Bh97oNeAFst6ArJ3m/r3E9okeD+BNPUmLM4IUnzapckR9kdIrARXPV81gyUm9s0A
rBFwRkLtjDv9NMzJQM561uT16v084Ys94MU4pnRcY7IIlSDqg+qmetRVDUeQN0qA
Sukp1j3D0fJtPOMAeiBjkkrNDsFCM0nRRvoetASyfA6HRS/DnDDwT+IVV28rxy2Y
oLw1veVAF0BLfoi58IJF/8yBsE1td/GTCOxEDopWyN/+w//OsFmhuF10w7F1Lpy2
BYdfjMv/SLnFbSgj3biGjQ1duaR3ARk5Fld/qv5W5h8xD1nbpa5LuKDOjv5Stnpn
tly0YVD+xnc9AelBZN4mW1U//CKxASjv626G+e6lhCLDsp49DEMFAUATtxz/6WY8
Tvt91GSawjxChbLLMFByh0JmODFlfFosSvOUwhHLQ5p8M05vGjMk+P70JMe7Ks0F
WggZ7m8XxYBBLZ+47hjAT8VwAI82YQyou7UcqwonxWE+mujCVsHX4nHFVkuzEyM4
TfIj9nfc3xCKp8Q9i2yDmyIUVTQemt471LKFFjq50Riq7nkzq56664mc3+Tr/hwO
jvgv+mSOd/9Bu2CFI7UWJrKN+i70mpE7OknNLm4e4zotQmZ9a5w79EcF5g5ZzIpk
FsaSIZr8UYdzZOod4tvm4+wcUM/LfIyx1siyjkwX4S30ZndDkrDqDgT1rn4iVE2N
Qh3Pd5Bl1BpAhpn8FQYhSzf9OVW5U/5v8cwmfHmhIXUo6IfH9RS+GswPN2Nuzbtr
vQX1+pU+6NaVN61ie4+4SMauMrphwyxZWBqVybqbOkG3KqS4SQZ2o5cZxIFRNFCw
y8v+QIAzro8dY56j0MVUl+DHrLUzxseLmRxbmSH10PEM5d9kgyOCoUdkymNJapGq
u+WJcUzU2yj4uG3L/PZ7zyHEudMYhMQMsi7mYhjVhbPI8evymG6PhXhUdAC1C77a
xuXg6RKr0bSIbzvNpyeMmKvdKIlVbVtxHZIPDGCa+hpm/jen48GsM1OMac5ge8lA
iTzT0W/kWl2OXo/YWN6ZCSsVkJ1rSSLs7Clws0mMMxFuuB67plZnX1DTVh4L/wqu
SThUxuwq60U4K8ueztU6Gx1R5vFLbkdvnxKQL9KybhpVsIS6mBFcryhsghjGZnGK
5oSmCEAaQ87RMq7Trks/33MSpsszt7j+EDXqg/6lUjSCeS5wsYUq8LWrUOY6mNuO
EItnTCW6DQfwOP25vOATsWTN9WOTM6f156VXaxHEC+We0Ql4wrvSrKRaTfsDgs//
4YpV4o9js6MB2JnKOxvC+1cRbns4LHYntAfP95ItFqEieugt1trlYDvqB5km57DV
YT+FEVJ7uniX2+ARkHQDzXr3PUgOsMI9p1xZ6aTll5K3hojyXZhYj8pPOk/FRjGS
egCGgghMsDU6oUsFoqzceeOtbRGZ7QD2kzuxTGmR0UJbKy6+Z4hIGpCBNn1Tijfj
7m6hZY/o+84wdryz3LSIG9XDBeM7clDv+mnqtVlIgjGzkVRDPlvBEU/JEp40Ij2Z
E2d30bvMMlPaJ9eNjGy2sgbl4cDLgWZg7njTYMYD8U1/9ccaSrkf8jPYNTcw0rpV
YIOj3nO/83kAkxRsCdo417RbIQCSvwkG0eOUZbZltUfFnLOjx79Bom7KIJn9J5o4
fLgt/ktNBg8Bk+q5zripPYXE+KAddLgg77aD9qBjPOV0+91O9b8dlta/Bf1wmGds
9bj2d14ZnHX7d7nEoal0Yk7iq6nmKTYvLk82Crn7Wj4BNQGfxThvqfahSMz0kZJE
+l4AUCLPeR0A3EmRNkIiN1HHThlZWeyvGI5kbRKlj4CC0scj3xs1wpnHS0RM0S56
I1YobUlK97JOEawSkJ2vRKvr+L3XZoP9pAOiVEyKj4NwgBKIlH4qaBR45rjJsh5+
Z47CpENAPkeODk893F4mm7T/tC0ZN2ZEa4ULJ6yCkZwYu9UDe6kfSDAqF3yMu00V
kotAokE4kbYvq8SHWsH/9/b49Wclj5Aa2PUQrjGhho7mdPi0pGgoUaGAMG9ApsQf
hOtWtpxQmJR0gC6jtgj/lZQOMC53blw5szXsAf18KkOgn7PgR5TqPxr69dFn7kE/
UiFy5njm4k3pkb/qeWpx8kIjyRS0RBOJI0UXKbvHx65LN86xy4IhoI2Dw1xJnNKs
KeTRk+KsPwWnqsUa//5aCX0q0ldFmtB/Wxl+vsJkC3Ln6hfvnnji6Bj392C+p2qd
coLw+FcLRPeF/H4l4Ts28Xfq/bwAGuA6TIULmqKi2mgdsH5o7Y4YVpIVTntf2ZZE
mDpdAOGjtnHpolTKTlO21U7A58jlUJc297fMTDYJQ8nZgXn7d3F5VoJoqD4CGBV+
nLCEmi9vyzOtetg2xWxi7yGyhJt3vJdxrWRYeYCftruJjqY/CJX5+/ifiv+NrSCb
ewnVS5afc3qG7lv+fjRhTTLO8FjLF3uHHOpMO+g8XZTXDs8YyU9LYoxdf0anVIYn
WXMJGWCm4I1304G461YdDYvuRdnixKIj54IikwJSNHazEHz0nkMkAMo5N6HlmtHB
c6wBca5uCwgbU7jAK/S5TTbOCuigFFwj5AoFlJ1RQFCw1GbcJD15AKIQBtP9i9n2
No98c4PPV8sPcp0yA3I0FHpm9ERuTSaeSXukF3ZvzGlB6WPgjWHdDmlUEGWxkHgY
YjYuJXxCfhpAUJPQRAg4OwQfkIguXGlsPLYlMqeiHuaEsRiPMIO/fQzfhFupYR/1
PCtUtBTtFTOJmujglr9HehGmQ6dAxcwaCnayg/79eLqMqvc/Z06GcPCasz4PDOEL
HhKncU3I1I2JwCLIW4nUeo/R4rONRj5b0kpE9f0pPgNB89yKMQlg3W97PR/CGKiz
T7w30ZEZCVW3214Tgfhx0JHi/xpfvrUfsqZElD7Krwsr89b6qhv6EoqAeNnsu92k
67UST3Qgox16y38hAWUBXJBKr+/BPdQ3RYJOwGTah75QOj1QAbu+3TCYKgHsP/np
/natrOGrBN2NFMhnkzVHj5bAx/+4krTmyF6aNWdPif0g7LbVLytzp2zgyoHIDyfl
fhPFmALxYfikvojNChBoFsjmPtpxYJyo4bKCX89/Q0y6aTo7aOBIqvV+Pfx3EXP9
SwINXLjMuzlyYSZNQw+c4Qhy6u2mT41JeEtfRCIXb2jH0nL2pJPjducMpAdAv9vh
VDDuKYVeDQE6p3QoueAwDKMqJoyiPepL/q5MwUW/BCalnvQukbYKA39OixgDdkYy
SYyP3q7wRw5SHi+IUPyVzkMcNUK0YHHXfshfubU0jsrbHcyQsYHTOEXJHrfThTZn
fdZTGorPQgOP8fgcbzzL5Fq+roSorLP6LpPWYicOcQgFeLmqSBtFoTN/L/bJjYdh
N9/8URjnk9q7pBdO4UdCa36I4+M1xWFwff3Rewp1kE7gWAV2ghpArhwi/E+tXJYh
vrBFcEdNhOP3V5YzM4NAWYq3YZemaPyKMXbMrXAS42WrTxoi50EQ/sH5TkyIfsrz
I/wZujE3/WgmEL8GypKAn2RlqxcHB1m56LQ0pfVI7M4l2Kdv9XkstUZy7nDDJmwA
TmYaxMNaqit83tLyDgW9zVwNv0yl7lie64uPK6BcwnFKJvNXSnKoaqknpNZNiwzA
cYDhWliIOqVa9VL6qFzDlg0C362vSwAx5qW/wLHrFJn+eLozhsKu9/SXkIYc/y6c
FcP/mGxXQPIgmLY2fsNMZeZahQpUX14O8e16DgjCfCv1Ret+7QBv+Hspz4R0pdMs
cTe7RblpvARXcE3HX206EzVXjefNRyNWKY7LCI6uZJ0K71ASfuq/m5syrOyVvT4c
ORfK4hji4RoKjdeVIWQZ4GByHnYycyXHnJbowRjImrc93beCCpC+fWfi8ILhFh3o
guqqKcEPMwt7fvLkBRF/fZ+YuTocJqMoOyw1YRwcSGN59Itl85XVF5MIiU9Ud+RK
Zn1hdWRpui3odDh1XeR72HoimjhokNvxUEvCNQwOUyx18Zq7OajhqooVBBH/KtDz
TmXzS5P38XKEVInstCtuj3AcMHv/rtOhpeuA2NsifrfoxB7eIQDlAoB54LLzwNBC
p9hLWRDY3P1m/xT3BfnAlnvw8DJbEMHTg1SKMX8H3Uk0xydGuFIRQ1lEQSk5Woy/
PpkPFaUA9XLcq0EFvTFbsxVGk9YXum22+ikKyEV57QLeIoMUpVlp1WMXlViLL9kZ
jLFbpkL/Y3+D0WCGXdI+WxR/M9abyt0KiJeFQoETdqX4N05qBx2rqTcNM2eFyvN6
aAvLZkOTQh+P8QokBjT2w47YhQXxs+ltIgaT203AyyMwG6Mt9BNMLT8gH4kXXn4L
XnAmKouCBRRsj+r8R2TXaxQHQtFFxWfyvIEqcwuYMd5XaPFQAcxus5rz/3FoWAef
3+bRDx/68NF02dR221xdIqc7eQynyyFssoF8YjAqye0nmcRMFhtm+k0OUxH3T5C1
8arPAMLisX5vjQsaZIEfUAEWdKpAqKkgWEUxbju3cuJdFCAk4eeSrxTr+4heA372
Oml+21KGeZaf8ylHGl9Lnc+VxZc9cGt5OtEKKmwEXNFe2XPfuNeJDMJ3X1PtQRzq
D9B6P+rFzFSENhEcPDWFHGvqzO26FIOClpLQYpCYg/6wbPEQVLvEL7vf3Nd/03f0
LJM6PUT4OVZDjn0xO8WnIkXX2gHr2mwFB8XnIkIhTDExVgnrOTFvaC0GN+nBrE5f
a7HtXdVF90TiPP7/RaXXs+cdsjQtLbxtCCS7cKKl7bSS2nQP1lCThMQhBFjb11Mn
6ZrYonLmHyfrEbnhQMCG69XelyDr45LBy3PXZOVpBFPyP5HVg4z6CrSJt2EvoUKX
26urSE/h+Ebv/0qs43/ja2i3PpUihylftm3ah6Tg8z8jZJHYdWY9m2NaF2o10U3C
iSqqWn+Ii0yyOTHcsx8iDOOeIqpCGmAHdMmWMhRkGF2LP05owSt4U2XhHKHBVdGz
tIg9QnSQWnh+K1t6lEoYas32uuVLtpELQ+2/MK+rBJ8gvecVZkNDpBs9udg4Dh13
eEwP9eCNDYArBN4fnyPYV8xaSqQomuAxt94EcO8A12QOgGsaXIzr+pMVt4khXqmr
hw8rMhDhnox3OEShk8r7L92aaFzRkAZA9aVjTRSXqSF85PtT4+ZvSHhIS2hH1E/h
OTLMj+rW4Nk1KHH081tlEJ1BSXncnlxeAYt/cKdUZfroASjI/3XQ0wAV1Jz41/Co
q9II7jaH44OdrJ6zKZkYQggB+nBN7lwLtwe3plrDQLhid0XaNRGVkMsqhwxtjSP8
zVP9Anm76uaZMeDu63JrTrkewYUJzs0aU8BimUu+9lHVYJHy541IuKWSNLAGMqH4
nbw8WBktk6yQel8klZscyYNbXa1lB+1ZrrJ+NjbvvpNNjuQJ6rw00wTRxCmTm8Y0
mSTPq6mZSUdNidO25PKAxW8OnmRkn7ol+hlTiMqDRiU6QNt7ZWGx30QhkwmQnVQy
V+fqbYyNewYdfLT4nHCdZ2LD8q+B6x5aHHmroswkm9CBDRgj42Z+9ei0UMDqm6YI
bN/GScqtuJYJKXQPtVXSpCyZhML65NsJkzqGL+E11Cu9dV+jVqoOzj6sR6utnY4M
sM/xegoZBjlfjgB4UyXkXvEEWFzQfkz5iOiYZluseTWH3fofaxRmbPYZTj3QxBdv
Hw0eCMIrMvx3Io1KWsglCOvAinS9x+S4eTGZY4oyhY/L+lDHKNrSRxviyHyxleat
GrMtQYSTKLqZNMZzqqA9Z5vB2OVS59idpwA4EW4tRV8rn5x7wkGP+OO1tNk09IhQ
GG2+6AMUAEHTlIM1+wPlSMf5MnRhZQgo/greZkkxESmvF4N8Jce2DO85wVLJBmi6
9o2RZ6tdzf1Q4pne1D3aa6eH6LvrT1LhUxMKVnOD2ZrDFsNSdch5lsxKq1iTqvNE
xBfr2gc30t/8S2aRldVQVkIGwUXyuAI1whu0C3A9C4bjw20TUQkC1bIoJasPpjuP
O/63692yR4INtXS7SO2SXNPM3Nb8k6dzyVyJZ9Tat5FxQVr2OfvdPEnlh0cihUCv
Menbrx8P6HZWluuFoJlvmbpG+btOyEv9KXbGoO7hDQZN2/cf6WTa0Md8ga6nCmU7
/C54m2GRviZFud47BFbpnEmZtioD1jIlyfP19tiqpjNhPA18g0M8S2U4OYGuSLYB
MjHHOocNMzVLM2b9SYI2A/9YCM8o1/49NKgosH0HaSfTtk9ZWPhp7+XKYq7pdow0
OD03R6Xn8mtl0mz9A9kSvt9F3NVLpTMYuWxS22tWEo1dhoOGrmtTnFBU1t/pK1Zw
1Oa1B0eb0UJK2hKVSz60tlAjD1rz4/p+bo/mmfO2o69pirTGZNLmh+iXfUCrGddN
3gZOoZelrdRFl9IsqWaA7rDISp6RbeCTRpv7113bGC5NmR2r2XBIMrw89OFGpvBw
5pCsY7nAlkSZnnS/8ahAegBojaUsOeBxTYm1wUzaB/17u3dWLQvbG7RjSVHxXBlD
eXZmthtD7lUrshNniPSqeWensQEjRjIJOLF3pneIxVn2TRMyKd6ObWKtboXZbU3N
WSlzaKgBi+LP9CKMAks2M5mfgBCTdLM6T5Df5m9JuxMOCzbzNYp6RK36zY70246o
t9vsDkHtEoesPoyFzx2xasgwEa+UYHtyaetZqBK+uTlO1g3pzXGjTMdwZQTFwIvc
vx9w1u6Aw0wRZOMYRWsJzEPnXtdINe2Ob9IFSqqPAG70Ajabtdh6z/cUwQqp93iR
fQBZVtsHMIt7641AWlCHlaY4IQYK0fkc14kjMExSnMDitJ4qubA96F6TJbN/hXho
aH6qqwsNDmtCNsqsQTDhLwwcAVdCtujeilhmPAqMgJWH1SAciX5K88fl6VJ0Au0t
b9ugkelOrGD1HPFOcjXfAuuv4I8+BypAI9Sj3SfdCctjEjp3vGketTMB9Qf01Xdl
dFmWAUlxAuAzgwCDsQpuI89hiYWp/S5Q0x8YHhNZXOj2ZlyiUEesPzy17Abyz/LV
s00ZBR2XokgSj8Dla+a1Fmd2E7I0CpXdVa2LbkM0GG5tSfIMp54ClCqFMZQjnP61
kKOSvcHFSAlS9hdHh2oER9Z9HiV7+LgH9hdFqgKBJuR+HBMrLDg50mJQra8DzULP
1ikHlSk0V/wYjxq7fYhX3PGurDkuuWVc+dYGJkT1gwxURyPCNgmMzZBK/kqd25qc
lGPKTKE5c2nt/vxos85sqWtoq/u1eeEv/OLAUPAX8Ib0IcWgPdfJDHeKbPNfnpYz
Ynad429K9h0p7YQ8qKtY33A5sM7AZdY3GhNHZajyvipmMNfZs3Ox0B9jpGNKggXT
o3YPqRmM0TaQL7KAuTyLbbxGPKBicg695iFo0ZMTEvKxGihMGBKng8kjF51vFT3U
PRJOHEpRap5UPoQMI23Ztp8I02Hh2pRAfKj6zaPSUaNJIJoxZ/vvct3BdZ7cqMuA
CD7QnKEyjOEurGDqQj3nvywebIPu2A37L2C3XVUcx/BwpJZdNyUiO23rTdgdUk0Q
RTAZkLLaZyx68AtsLKyC2avBvw7SaBz/qQsfI97ZBQPzY03cc9pCOIX8ujO8POPu
/yi/EePikRnWFNO2qOsbt2/dC7d7FTeRBwVvykxta6TbSUdVjZh0kaqtY2y0kHz/
HsbUTdAmokbQiBCR6EiYDqLWn2rrK6dbiyVwRw0j57BMNrRNR2bzGO6zmDl5oaXR
kfu06tLT7LC32cmHrmhBa/SaqsKWCuzT9Yafb0akounZS/0banc7tHHYzaWxFsE7
SgAvWNA6gIfoYLy5gjq9sgMuYhjenM9GU2Elet6dRDdXVhnO9jVaph4ABoD0iqQg
pN6PjhyoNvmv+0dxWBF6nJrxf2G2FAVUWfhGBou6gSl5xzhI6+TdMJ+awSfpnaHQ
XFwYv7dsZnkHwSxEQTJcuODOGBmtFjL11401k2b6AEb8Kq5dMUsgGDkW9BK2ExGB
JfhVxdolbBeUYquDY0SBecgZ7iXMPcG36mMqM21JlL3eigSKqHNN9hZurDEZEYQ4
wL/R76TFs7sjCwhLd7bc3xbh2M2l4oUa4xQF857+gvjL3+3ZbQ8JNjqt1D7YD0eT
xwwsuyWHH3SzDQcFdWVD6kARhRdMcQFxTInB/gH1HrxU1bLq81rcZeos00qr8TIv
vCxpBUw8bGAkCYrK7uTmJSkg8kC10CXDFDOL0hZMa55IweieUlI3MENyW534AfNB
spxFEhuA3SJn/i5Eip20MS/UYtzRe6Ruc+yghxIE+CRpSWixiCgLtAiZkghBU3za
0dkIo2KOLnZVZscHypdi5f2M+dPgIDWQBZYnDuNDq77lAA+RILUh2kIAeJ932Kx6
bf+VC7X7KrYyuZMvhOU8uCKvQrSDkkWSq8JoyN2kM4apOGTO1LPTMExjaBrtzF1O
xQhBBXxwTp/j/bVColOLtzw+jdKEU1qIcmrBZ/Ec72NgpmKwXpx81reX4FdyXlX9
2diYyAbY3PUhsrA4OhnHDN7vjXT0w1bTKct4fEQjONnNq61fzxRtPE4rOZvT/H6t
3A3BndHQ6ZQKG7yCzhl/4rw+rUle5DmGL99dam78Z063vF7w1PG2Hy9Vx9oxU5/S
A1C8UTvs7KQQ/wLgKEW41gKots4zNDBYYbpmEnv+mavnbEaLW22MnDLAvzhm8CPq
u3cxd831+Ixobv2f/AO8RfZ25Uu+ML5bxO/HkzwdIawrIztnXYVWYcN+dFHwNqPm
ijbecgIeZkR+iEKdDtFaPhtSklgSCGZQCzwtlJxFzdkhe4unhlQ75toh2moCxGaT
l2/MEMnL/59y4Ol/07KVY/HLLHk63pH9dQYY7iypt1XWivtLeVYGiknmTk0kfsr+
3I6Ka8J70hHs+o3g+Ah4uQnt1mQQMIC0tlJoVo2x9ndmFt9KI0EXT9ZFnDG30ZO8
+7+AheUWnUWd1HB9NMvfq0Fay7XIg3EiJjIkRDFGw0I90FvBQ4AaEwohEsRmSVVC
PZF4ojerjrm/gklGh8g2ZFMtgKrSQScDwAW2jhXM5CGOZp9TfQiKklVeONz3jejj
L+zrIEEEJ09/SFnGQNaipazrRd5nGSoWype4BktVmbXlQU8hUv36tMpD1MRhPwm4
r0MdO562CVwlSk+pLK03R2uRtLO+pHxn604iXVtyGX6ynZHdZbjaGlKYFa/oBvs0
ZV5D8vJ8kXCFwK2Iz3l9yBIlXq+oaoqw5jKNXHh1BkpPV2U9m7yEd3wew2vkU7oa
IZUUQgvmpId/RiPr8JterNEXq1H1d/9mSpQNLr8RnmVnAFqEafYIhilDCx6ea2rm
DqvAt4O6+2ksmrTDBdzgocSEMb8pjauF1Wl39yONjd/FVl8ZtyRRJl4tcTRJEk0e
2to5fnQ0kjP9QzEDBjgb1HoTHbqke9JoUs9crCNoV3AzjzlOK0EAE7niXvAUzDfT
FMMvJ80JCMKaH6J5GUCKAgb0lIl32g/qTxCV5vXI45DeUZeXOZbYfmrDPVv69YWi
hTPE37xwUmBzhERjD879cHq34NgkCimDeZcutXI9nBxDH9TeGg+gp2d98YW42DTt
2r9yTD0SEsLhi2R1hRuTSppIhsIbFdqqIV82Hz3X1ZS5UOy/0IeXBQ52q1z3sRS+
BpJ+Ar3doakIoBvTAL4wJLWVWld8dAmExsPyTUsY7M9HotpqbqVF7Kyw5jGWUNDX
i6mepWWf47dRIqtVSeklQ0qzxydea1UEObXtPBOss7RHS/E2GlHeFqtMpAOqQdMt
GIU3t00Ylm3J7SAC4WuwE1+eaIoGaJInuY/Tswszcfqz9zxgcKAdEuwEYHyuXTdi
4Mee15j8crRY5EVNFAiFCPUWbcvHOaX3DGjQ8jE8rkByPXW3M0gYQXmyi16wwM3b
/mIt/t0Yi3um6nYdx1CC8JDSRBd8v4oQ2O6s9QAWvJ4LvtqMrxI0iBOWCNxA0ve2
CkKxh6HDtqvgDnfYg3pu39ucHhbbrx4ibh5xokEmhlGfO7ALdh/OzeyLhV5XwJa3
foJuEwGVmtHMJtqwR3skNFJ+ft/IIEExs9M5BUTEyDUEw8jrf5hOps+SGmAk3mqp
m/Bcj8OvKhiuNqPLul6fP1b40rWm8Za8/nfKN+rzsogpszLpzDTYKokmAR4hM3+a
xX2sH6tbhkP3/kwJbjPUWnVHDDH0YJhqEPETygKBvw9+dok0E022iacnBuetyPL5
TR8DhiDQiWtvvZH/6EWM+M48pROytDRJo0uZFvIG4fSmBPFHoFEMyymGs2O5fDgf
0tPdsqanF6y6z5ZyKUO1C0anAm7YyuBmip6BRKat7KimUXf1IuSuzYJcaBk2+xE8
lFUfGLl6BA06QDLlQ+jVvNtDiMNmVRmSpkHigMC8WXTTCVfYpLZzjP5ObIMELesJ
6CUaPCM+gJRVoBIXlDLQhaS7q3Ce68fwdtX8ThQSdkflglA3PYuHf3EQ/pPvhiAs
tJx5Duw6QctqAYbstwTI0eqrL7cy0FSF2H/xsJITBs1JsJnk58wKu4xDjljA3eZm
8iN4XMQvsPmj/IioCyv2iPdSu2Ain1PGxshLodtaTBrcB4grO4GDQdt7JpUxKhMa
/vb6o5bO9nWNTm0AUt3/Wbi0eFSDaJlM+9qHyBIIbBxO26ZZa0qfPueR/RcBdlJq
vcZSnUkcv5rNNmvui4KUctglow8h22oW76eKyoiGCvWR5C3e4mWVkCaqQ76dkX3s
I5bTohl2bKlZb9YqO20hmFITLCJos7lslszFiN0XfI+ios1FpARAYmFvSs80qNl3
peOMpDrK4tI+SGqNDk6oSdeYF3EguUGPN1uL6gZaKhUXXJIP3+V+oyKEJ6TH1X3O
pYWHa0qlBEu4tF34hUFZsXr2e1lubxp3kRg+nk8oPG0isQH7L1WBegxl5O+MdJa+
FAMu4cn72ASLjkHtQhG05TYtguXk2a0gx7cqVBglpbyaqPtFDcPpJ/zcpRMZFlM2
twj31l09XkYQGZRskBNoyzCW0mub1ZciHnrponrVqUmXPpJ5BI+QXL2gEg+abC2A
smGGMwI3UBedLblgocd9jYrt47w832nhvKKpFh0BGRkWKV2wwkLCmLHL3W1bJCtv
NrzHi/Mc/rSV7rBnvn07ZE+7fNkwHOj/ZRWK1bT0xE5/XxTVYxl46oLC4WDDhCwk
M9PxXnRoYdVfjKgvzH9umS8WDHSIWaEab5IkDEOO4UyOSGYx4Na17/p5T3YVucFS
fAwODy1tLKrB07RgRm9T4RFY5tVMCpXUq7V3yNUiITYg9mSrkzlTTPTv8mo1bxD1
h6GIytBXQBbsPS4MPSOsZKXaPnW/dofGJVRgC6EkjhaRVbmKvTzJboMRORP4ZYSz
OhfQKSES3ZY/s8tWgsOfXS6ksJr2FFHZkIG/PctQ3AbOWT5n4qtfcQma2qTJc4IF
e3YOfTxqavzgyacu8eI7Fq31ZzNINtD4nuo7tjnMx/0A2Fkm6lWbh9qeSzyENAE+
8IeKB/Bh3r8xI8pXSIDcPq5HwHppIhaHrq79dgNvD6bIkRJfYS1pZWOr429JbuOr
Gzcp8OkVhMN2S9iV/Z3SfIlc6vZRjnYME1T19sFCCdKFrWmWiy7pH2hrs1vSEzaU
T4J7lU5gYF3WGFdR4LLCpNWKgeWW5yx5UjYUL+3QRy1qVxy3SNLFwy75ky+/AptR
U0rZI2ZT4Vzx9K1YXwwSWoabk0zcHWMGCVQQeB7XLVQDOpCeqOyAdW3AQD3dZLky
Pw5+y7pfQczufpwG0YoHjY+Gbr5dTXaH7iaOrTdnqAj5N7rAMupTCRVY7wtYcw9p
qNEx4udKdX3j7N5G9iQnAbEMbI5tZZ8qmfzQOAbw6NiY5w/U0cVN1/2MCT3DRJps
9UQrj8IY9UU0cGMOq6ZUce/nRgoExl7sUChO66fhgJEh0SjHi9BKDah7aud4wUE+
cEAtiqnKodUXMKkpZSJyiy5hWV2LUKWLXySXiG60h3YCaZtDWSoypowi/OrMCIse
ItzTbU8RI8Iq50jHnNQIqqXG0h93gXJijp9kawDkOokYBPXVsWx9o8eWwrldaVl6
BCvcbRVAvHsXny67DTyfIZY0LjGIRKqIKkXzNXTlx5ubFyJ7E7NYqoDcHyyN27FK
pVtIDodyNH4tOKn1Iag6N0yq8R8s/rzHqCAgtLBJKZVZ0J38+2SH9U0acNSJkMs0
lXh7VP9zp3/YoxzfYcSNQi5xE08/OzxtsaTcAx8WSTRmd8+6wFSH6uLLbxS0wmld
zOrITo2btElFK9+BaTJrCupe5/YELu8Ec5vAQpocZbUaB2PbJBY9w24W/+uAp4uA
qB9ZSp2kjmuOhcqjnO1+ghuKJCTx9Ghi6iSL4DGcPgp25Yx3Lgbk2O7rv+5fcx3/
uRnbGE8e2GMVoUY9EbUelIFDQfo9kWcf4WiBg6SY19CNN87qAbuFZ+AcR0rDWtQt
SU8MpY2Mpjx+nN9IiEXz7KpX8eKJgLkNmpdcIWGGk9a5OICyQTUk42FFXYULcIK/
FSQyJL3DBOihIz/ja1378DLu3FDajKqzMQgeJT8TFbQQI2Q64OWTi67UfVsTNDXR
gYPWbpFm/7AZKLNceEG5NlEBwueS0PXAxlXEzoOfR66KYdouNu+/5/z4c6dHHXMp
W8XFjNmvXZVyv0vcXvQBQcO2R6e6xrdDBPleWE/LQbE9GChvtohbTTkJMNQXVyZB
diy7QImT41f1tFPSOI7CbRcq8lKNyT4xz9zJj3YBLg8KEJdkjwYfCsNKtihnwZSL
SNVadl5yIKatwjU9hHfb2lzMkB3BpM3O9MH07L16zv20wtkdShHO2Fu/FOknp2vX
X+cEUpVvvQh95p8Zi9nD/K16XSuuLnjgITNRI4vYgXMJlSvHrgHYRRtjvDFfogX6
nPaxP1rJ0+aILa+TkLw5S0O3ARytYNYrQWg7q11iCa7d/7XI0aL3bgVXXIiRSmRG
YzpgLKwtUA5dRVgjX+BnuWiTUIc5hrDYiSqmNDNmhhKS4ZgQ2cAFlSopXPi9nJVA
v3+aWKQROj/oF12ZPeMzRmpffgLOl8uvoW3xi8wOkb8RHUsyQ7YhR7KmqDmscPMJ
J91uqm40x7GvQoDQqwgyl1OFFM6bNrZDdIvZ09zbe/URWNFCntj5rIn5Xcvlpus/
MUmQmbApb9TSz/4NOaoBoKcuqORgKjrpin8HPw/v230ORH8vNjyNFxTSLSazYRcT
bG5peLf6TVRnjM8u8M3/LJFZ5cIshYp22Y7GB64uqEIuKp03lw9txJk5oJoWqQ8P
BwMWXM1GlMzJMfif/p9qBO8fNwLKxp8v6EJWxYSyLbXz1ymumh37JnOmUMRFiosL
Cbx5LiG7OGXhS5rQOZSjKpOR6ZJ2/YEJDowRxbAc7xw+rQfVBcVWM0ETRbL2Mb2t
l08Tr2UA7s8CJGTvu2SiZKfOmp7zZ1ETtit4eLCIZa48+KZwBumuf8+S8DWSz+JF
wEgpYXNcc6KEbPIORn6sA+GerZKX3go9lA5EoUCfwVrrl3PqFIG7kV4oALLvWBi9
qp+J1BdZApstNVCSI28wyEx8WsxIdpheRf5BV8cl15/4fyiPm1gOHhXcO/rl1NOi
19U7stJw0YgSN5E66au/Ekgi4H94b6wYovwejTt4KK/AfegL0uK9+IrNegbaiqsK
p0zkcJQCTweRUfpOl/XM/t+9coYZrHv69QXSnFsohSXrBtm4OE3evK62SiDP7nge
nvsIHdPyj+/bP5HHGxCGp8brMWcjooMID5fZSsH+PDO/MXtYQuJkxytXgCbgIGzM
9L8kLqD9U9+kOVN7TBciGfuQBuUIU/hh7f5U2mM5WEziO0MkPEXCFi8Pu6YTWMHN
i8zyc/Rqd8E7Tw6O7qlSIxT9Aj2jbVmApzb9wgK04Qo97waa0XHQSChminIz3rAD
wto0G7thKmIVP2/WE8wLoI53fLRrQxyUgXcVRYgOziX1wmu3L9l8SCynj6RK0Y6e
oEaQ77TQOcSI8zQcKAnoz1VUjOxOmePQDeWif1BO9emPDU0cFaGeBR2y5rmvuuDT
/IMROyUgMImQgUuRUEvhin+4zvPTLVndy1MjGpwjKTuNoXVnqx87mx61mvA1otRa
FMX+J+zumgP9p5ddzDBXf/JLFVNFGyRD/lswqfS3tlCG4TIH3o5FIS0MmxEbK+C9
mFHoPBss7IZm4ZwLHc9tuDxxNMZAc1l9UT/EvdxXVcqfF3PChuSD8FyiY4EePH3y
GN0n2b/njxDEgfg5YAcr78J0yGnBixtrzIoZKuSK3jPq1slgya9MOPAbjULnP0eE
RApMfN2f8HNAeJkN5/CGvVaWsre7fAViS0xi+P++By5YCxvI8EsAMEx+H0po9Zb6
owmzUrsQrAyXpERcBzlGqc3sgQESd8iNR3QdM4lH4QJnsg7hunYZ/DIJci++odpX
cAD+qLMy+PLd5/39r/l3OHhaMcrDKoDhV2iI31AGGWh47TGYpZP+vG1WVkySylSb
p/uGcXUbvEDRdeFxg3/+Dj2qm3doAX7ISwORnKHpYikePZ1SfOmlRYJ59Q2JHpMR
lVt32qeiP9YN0Q8gZMs3Iy4jwFH+mZ3uxUcEzoFwMlEbx4EiutWUtFfGTpsU9luK
p+0Lw4q7LVTHZ+JTPmY4R8Y93T8IPc8w85QZ37/HgMbqphHUG1lRQI3dROX3JDps
XvP6WUbuN8gFVDb08iQQKS/1Y0Vmxdm8oe2zeXvoc59mHua5aHOf+ZVHcE5ewlMe
c7lzpQtd0xhjMoEMpRgLf9afKPFHbJosdYCLCcp0cEUN3hwYwuxxWO2j4RLQe45J
LLtXIsEcXUq/y8dHHJnkfmfNNN2CiraKopoaaO//tc6XO5pQ1Hs6zVS87lI9epK+
Dc+l1BskPJXLe6ydbyMJ+ZhZ+8AaR9EdIkjYHC5T+Z4/3NFDBrBVa+66gkNdkmoc
5ocDe7s32IU28QpfMHB6dL8ORDPmUHtsGojCJyFgNbiKkrtzwI3eQU9NWRaOXFwG
ach3j9Qb+ZfE2erIzd+YOCRWxuT3CIigzxZSL9xGXd5tfWU/nchbzmuB1pdOYhSC
iptvh/dET4PpqIv/GjXAQ8+hp+KaLNmnTO8Dxj7vKx3rw/66VYuhTyANvxjdKNGW
ijNkLEfc2mHiuwbF1Zg1nC6nkcRAQNIvDAvceO7yrd748yRc5kYvA1idXf5fhpuf
Jqkn/84JJCFV6/Vda5QR8puugYuDP7otJCzdsN2UYyOW18p1VjJGD/usxJiFSEz9
HXoLo956OBJQ+5fC2A2Fz1pWkk3Y0UDMRVka9JaPEG7kkJGUkKtKSv/i0gStzlcW
N7jxRgDBPTHOLz4RAVRPNp5MSbLcWCoixH2HyvXacMeKqIc15FdVpkuQ6DNycnzH
suhc70JihyqvDGrinyWXPQ1NDUQLBAkVDYOWOtUB6jCfwWehnRNm2VGhNh2ZuyTA
BCCrbsyOTahU43qTJcICufxRSfvWEKzYAY4VlDG2p4CFpq6Xlpr7+AwloFs4tyVS
7ONrVlMpK7LOZuxWXu8UBUjBTz9ofsi7AQvfsi9ESpFlsYR+H0XUabnEt8coaHqG
yOHT1fTlQgvlHGChmMj7vBngh6zfOc2QRsL3L5Hwg+8sP2vAwp1Iofr9ZqRWiWWJ
d8Zm2NV1Uow+ZQeLfxSOHMELVkRzAufK/Jt7UGsWtOZNe7x7sFwecQMdmt/v0aDH
eW0Q09UVVBauwTX6L6/I6dnLQEcMyNZFWawLDIxf8nWuQ54887ElNRDAxusgUGwB
8+N9ZaXzEb5Xb/KWoBosnRZ3WVtVPnLPQ804eKUH0Cg2O+cziK51yqmhzET7KanN
wpJQH9enfBCjZopseDVNKt91443037FWSkuxVENh/fZbvuhlSGZ3buU/T4e36xNw
7QDkO5QENfcmPeAQGanOsCRsacCpigocDW846VfCLRHcZA1SG94yBnhBbWv7Obw+
AT05YZwTBdKXkJhlfdOM9mXMeeDIq628u0erHStA79RvrgH+zAVeLqsX2YDl4fxu
n8nABQj3lx2xVW+fCKL6J7/6A2dkvu6dLWWrrVSIEQUcprgB68qXmac6ItDxIwzh
pwV0kNHFDXArIewceKNQaisYyWjGw6GTgxP7xtZOcCTFWWnYJbnwCcM5stUtLjCc
dixmAs3ypWUzSiHmp6+PalSnkCDIIsXmJ9juPXFUg2OM0TlR/qFUVJPcY2n5+XAc
hr/oaK36952+DRRDTG9v6p7SHBqrA2md7vsnFw7rOoxj0nVnmiH6Izx1XwrcvPPy
pDdq8SW1zcJO+yb42nEwvk23DOTKoQyJBKrPXCL7zOkBnpz9Exov3w7v5GJyoegd
0KODidsFQ6CE4ldYT7fuJZDgA+I0S510aTU1UB2CkA5OHiufwgznqYvqrHpcijCY
YiVLFs4LkOFFX9N7bubx2/gI9ftCkqCBZ2409dXBKfvRrYF4qqaESDoakp4Hc1iC
dk3QichNCvZqIbJVnQWjOWBlzuFALVmxmaL2fHI42Z7bMlt6Lc+gF/o2BLTZXWfY
K5VN8T2G9+5+vpUng2PHhJnyEWGNGGENkE8KeXa1zvHVBy5EV8SQ0PhDkRKb7ghb
BeCmvjqkOCpMGrs+S/TOzEEqT+kxhcOnufUytFt9jWM2rzWIHLVFcuFhp3AWrwVa
kl2bYxoIigJkPS52xK35v3FcHLmrDhX+EthZnZ5fgoPnTcHwPWG/OgkMwyYbR7nA
sl47kZR9GR4wI0Q6EzngUyZ+MlKyDVtV/zfGWT33IO8siETuuUeCAbBBo0ib8xoA
5rya1aPsA1jlBDGbW/w1TmzUPBnbudAOp3tmzjrKsd2eZsaDpDMxLZpEsisS4iQ1
87WBq3gyIaptn+FUTwiWfjuFPGmooL0Oa91/lQqYdWU9KtOKsV6a9cTyPrXz8sYt
9bHEeuLQhp6GYhAB8hlPVJXTq9+bixG5hkzhCHFMNpo7Pbw2mk+0woFZaQAea2X+
1+1vWAeaWYYZ87aOtymxgpg73+xKXAwZFqaseLPpN1i7TNnX/PDPd+QqCwysjuJh
7h0SoBKBapcfzQOaac9kstTkunEixpGn5wl9GpZtC/OOTfjeIMt+7eg5izcWd3+m
jZGYKXHdofLvdgoOCq5nMjI+/OY13dXAfiJRawWAuhGqO7jizZ70zz1ZpYn1xVDa
J5Vn2EIhRWfyb0qCM60vhOH50DtUbW8K4a9iC0NqGtB2tFMnmLCkuxZjT1oBC61J
qkdzA1su5nBD8l/v/YUfcotuaoy0nfMPc4iP+Pi1MAAHnzviNJx5IuBYV4izmeq7
27TU3lhGqkQWbYGTFm6S+vF5YEk82Lu9Y51+w1yZQDWr/XygZk+BxdQV4blyRwUg
Cp/cebfIMg4PEuivfzzd6WxTwkiRSBCNmf+v2iaawWTO/s7IwDuT8qQRXR6lgVE2
4N54XEcH3i75hkY3Yg9uBCvNmumrvGAUefbllPNB3wt07hEbU5/IExmkWs/bSx0g
avNJ6L6yELZGXaLiHEt+vf411PPwC+MjVEazi/EIt3Ye7YWMx7uIeQ9fZ1q0ezuX
NZEUWUr+TqtVaBjXiNdG7UHL30rBfmfQ/fAwQuqkxH5xXDGnRb/Cs6iN/61aevKB
F3FEa1WArW54QvOuyybTpE3caUyoK7A7l+5dYW3UDeE12wP5jGlQprs/QlN05txt
qJewbD3YkAKJrRJNeSnrMLN1RU34OsVDZrLLY9NeRXPu4f2mR8wI/LjWei2cYJEb
Da1RS2svdcqarJEWigF+5zD9J5cG513sFQFf3wllNTZi03axoLLuekKErqja/4g5
TjbjATyIaw1TZNESyS9+vh9SGu7tgkgAhcgtLOcjsBSdNnqCfIEL7bqNZQTFPj1z
IgEcxP0e1rZjd1rlldezWJf00v686RDej89NrxJGEspbrLxlnu9gm/sUN+15li9E
yqkgHm1AoMvwSn2VxojZfa78sOKgYjRpTR23AKTm7kEARplVzQd1slLR2V2YlV8M
lMtyqLc7fmi2pyEYeu5/JDugFSLa5D4jA3Ey4oHXmqXmkW7ev6bAfW/TMUyX49zj
9nSSvoWepwu/LyDQGvmtTQy7AgPju6/GXZaB/62wIxlQKa4ugp813jjR8BHc9xRJ
KGlHp00mDNbQARb7hvIrYslH+s7mXJ05rdmP8CPe4U2AthPQmFOmMc8vMZpIUvYU
RrWdf27/vETfwGpTxgNmNdHJbIirXOFdfnrrtlZgXdtqPoeIS8NIcRU6O9zT7sWj
UgkcFWW3J4wrEzKnd44kVIgSaNwEb4u1ESm4rSd5YRl1uVU7bU1JEzr84s+yAQxV
fhTbzt5SnylAurW93dJfBBKXWf5mOQt42lfBxnCnCafl0GZtweTwrBceW1zYHiaI
jX/NSIjJP9jlYBhC/jHntosvuenHNtggORfJIUwJZIHorhDzgHSzdTZn3By3jBby
d8HVxMJYBCPaQJH5gVYfLRUP8xX+3NpZ1ZmtHtnNKpEjUS9RnIHOTMyLMPYAiTgH
CodvLBXeAkaJxf8VqbE7qkmY03tfGdwDamT1n/8RKAWMsAiyA31PDg9W7lTjk2QH
0PLAOUe2IeM4RcOCDREEui13NTVw+5GyLSZQaeo8ufcIqRJ68ATsaQSbifvtkWp/
XQIkmaDbQ3KzLq9F9vQ+IV1s7XxQov108O7j5DULXcgzIC3f2lyNAwYQagBOLiyj
BmvEax7rxK9OE91YMiymsn+3dyBozRtVdoH/d7E/WR6Cp3wg0fx3JRTwCBxjdmEF
p6N+7XnxzYd7FcPE52zHQ978zGC+w24BYASLdHKEyA6Lb8c4g3kEzbtojEiSpUq+
466VEBnv8bQkFLvBMKS/8RbiTaKdpk70JmkN54KefxKSKMvgLCcVgDTWoeUeRWtQ
h33sPx0PV096yLjF2GZxPXCiSP93LyTli8kzw0YG1Rsqn744qRPFC66XJCmnz+F0
9zSb8qIFVN8JkluJ2Z2Fs2BI+xbVgBD6cQLm7i0sAUdB4cxtZREDZO6vPFeBrDsF
N/rOqAwU4LjqQm9fiSM6XW9d6QVIVAZzBdHgW2yeyk8DIWy2tA2BGni18Q3l+AN0
4BtKGGLdEJPYyI/z4ZBX9dVoU9kYWi36jThIr26ApovVascXvJNBpBXbN/0H+u2N
fiyF0bxMk3Eg6TKDqJGBa6FeLH7K2HZWfabk8hVC9VrboS4q1UaJvVfYdERkbMNL
WVocwdxsSWzNV6febcc2zo95S5vkScDWdcppf1GNfqe/fqQaOxqWIWhsihOrN1pf
Lhw950d8h8Z2vTLQ9Oo2ABX7eVK8d3POYHyEImIUVoxEYxHGXph1I5x7GqBAMbHD
nVkbQdi5Aeg01QMtu6IzDvnE6rz/CHHcu8JeK7wndKv5DN/GnbIiRUOWiLs6Pi4J
DMkw1Idi5GRs2HPw1zCGw6tk5CYA24nu9wcFPsnVeSUB2dD/12KwjQfJEfQyEO3a
HJhzBsAnTo29GS96hWW8r8GIIxLjqSOwy1XXs+gvbW9RrsZYJGQrUrsZL5OrOL2d
ZqsvN5ybe6SivqYL4zCKcziurK0IoV5HBhe+hcO9rAtqhLQvl5ZV7y+RWxT2g0Id
2E0Ifxvejlt9E6v4Pp9TA2s7xxaMlqTquzLcnDWt/lJHDJ18q9nOkeCQcDxS1sAs
IBvyDjwmYvOe0AKzMQdI7+GIw+KQipA3Ietbw8jxgnHpXgMx6IYxKWMDEuUs8M7l
1BTrk6+OfuHd3cudXyp30G5JZZMowdTe09wo+38s8SyGXUFCMkPpOtoE9Go2J6c2
l9xUvZWyMzEKvPQ4wCsEEdnQcPLJ/RbbLET7pj385vsIy2b59C9pEVL1GGK0kir7
vBP3S4gxldtMfiSj/r2BGdtQFfHpk5W3ftfOCBvhk/dgeseAG352Z0emhaqFM+mH
Q4z+7QBh0kegyXLmldQkwpCXrQ5QFT6cEbBY19FwFWWn2Ahz+d7VX/Br2+uh0Ido
8X0LsoXpxv+fYycqYAKd03NgJY38lbfUCfAyBthPa/XpE9B9CcMuLx3OFGxzS9FL
aXjB2d/LxIBdAsfilScs6x728Mvtn9G4fiPwzyh6arICBqSbFSwjmtKwYXY9Yhsv
N9OQIHmjjHPpSmzf4x2ae+jCtVrTcW7Tmf9Eg/dMQ0Z4we26YCwJpHjgzzMdgepI
ijt2ZUcDG1W0BtwHYW30O5ZosITxmzwUzK8OY89K9gy3fszhVw7AncCQ9jDCsFa9
UlLGOAs3Wo/IIWNnTArKF8WC5FaQjJt1bogagqlHZTZlssjd9QaVjslUMJ9Wp/o3
XCv05cfyvZ36Z1WJZ8ybIizR0Rnu8MJfFSJW1KZlw3j0O/75038UAzBdAWDNJHur
bAwC+h+VvRJCPmWBf5M9RWVJGOunT6kYELTjDKgPH0tFEUmmJdyO03IkcjzWdwem
FcycPXOk6E68V5AOoD6UAR5760P6AonQ0jJpUFEuZyonE1nBOiwT1cq+wtjWIwPR
0EfnndawKd5PgDBZA67jysUx2zHWHKsTea0w1RvgZhq1v6a+CMVu2zdy76hvfPsk
0LWz/4/tAEHq8ABeeH+3l3YAMV4uNaLF6vbnszEqs5ttkVbcRM2VFLwu0l1mCIBN
PWK4MeXHQ3ePtyxdO5d0uWTcsAszd4ndGTU/SRLEYd9vALvR2xIeXht4vSLXqQjt
2e11/uiuUtfl4jXxTta+KrOSWR5gl2/VKPdoaMc/8N82Cz8gMIwY/dAP5pfv+Mh7
IbitxGZ7rMchYUZR1/liTxcZYt744kM7Fg7U7GHeeIdACxDEtuB2I26B5aNWXwBN
spcXj/JJaeasDCbrvSQl/LBgyI0IU0ql3wsBvMkjVR7iZ25/UOcpGt+a/oznbMIx
wzW6KCW8Ueo9cQyK4KLPd3O9gpce0u0wCbCBKtJeCrJm2yu4yMSRa2N8wVn67HKu
llPuk9k+5MtHmU4Wtrbq5ZI31yFuhbkARC6Z3s7dXwDjX+kStIOlTpwXERKsZ+pD
w4HQxirBAv/HLyS6nk1K1c/pUrey5/IwnLeA1cR0Fnh4ytxE+M2ywuK/h3fz9md3
emqighg8/ifGN0f2XxM1csJe5HMzZ4NaggpY42ADccrp840Eu0zTU0+tyXMDz8vV
WZMND3LoBA/mEi/qc0F5YAITzB5m0/TKYoN9Fq0epaiFFqnLoNSdyiZo8Eti3WJ5
OJi/3De98m1YUeM2+VVCrb8YBM5IEU5DNTWoDNsr6qBtqmUnkHZXgjlP1cuimSMw
G/6TprdhjvDGclcpKBUG8sIiygGtZZ9lfwpCggiHhOdUy95panIhI7rAuOaaqsty
dc/GuFiwQX4+ifYvo3vIPFo86/XRcRONc1xJimxo8AeN2cLxpVxEhVyhzY4NCa++
KcyuxF+S7xMCPbcQgOj0ktqphI2wTSowU5qQqdRdl45rAbsR8acErA94zxzKBr38
mqOZGgtZpx3J4K7KSywTcdza3Qiuz/255lLryPp5v7KhTYhysdDq4MCx+NLbFssU
PLNPMzZsHNvjKYq9lVh2D8k48kgAvTWR3pS1FXOTDRqZKSjfd2uceB8SCgc/xHCZ
9FP86B82ZX9UanU1M8cJkYF/nhV/rwc738VL1EE+DeCbWiRdfT5KA3sDINVmz/xp
jjpH9CVHZo1O7hDoym5E6CnDVGf0xd+tSAdbmz+cZUWuISs3ypCx5D2QvxiULxHm
XQEW8Z10zjNV0YyS+O2jwKHnPPIO1ORH3EcNPLjYVxye+l/YDUzmAlfBk5m7NKDD
u2cK+Yu5DYDVg7O1RVkGlL/yfkTTyCi4KihEW5q41cTvlr4alCWL4AKnTqPryain
9+1emDCFrpagjmeMu7gKXx8mhayRFeXAF8jWjCaOcSiZc+oyFgjSfup73WgtAeZj
jHQ4dB6IsSwPeq2fXLNRoBhMp8SoH3W3iYZDsQ04UIyH84QBml1IEUbQkQCNo9Sl
9KdpZ4R+fLq4OVDKoijy0w0n6vPdiCqBVhQVs5lN8k8qWOi6xya/jbAWP909yCeB
cd35Lo4i9v0Mn+4G6Ke17hfoXW1f9xt5XaRhdskz9zPiNLeSz7WiZ5bBbPwjIVRK
411wlqvWpxx0OzrOCu6Y58vmfft2RbD9S3Xelvf2lwiEX7o970TwT3yqCujpg2bu
GE+gjNPPqrCmngjymtOynlBKc7V2tuefeYe+kStmcPn6Kxg+Hyn1ulUXnIVQyf24
1YE7f/8MvLKc0/YrqjscMV9wA3hafGsgXzHL9zIFfklpqJJkI7Wb4LpOcR91RqEz
5HyuRV6PfDQRrXWDc8UUehVITew19Kz0lzF1HYWbKrdMyrj9U6LQEzhffzJ7LrAr
U1TaVAqBl2KHoAtEHqUt58fTtadsYbxw4UkojFNOvhJybWKl2UC3zmYDAg4T7pTm
vnKRgLw/Gw7vBuwdwlnl/moG58g/AW5BJiREcIQDpAlJGa6pnZQGPwBwrlIfATsk
2c4pijHdiJma46YZiQVKKDXPDhdd5R+29DmYIDd8C1ngkXfOsIozTOQqInD2N1sR
8kbS6x1Cjf/ayApVuGsq3fuXspi1O4Fb27MJJjy4PBWqxCbx8KjYrCE1rQnJFE2B
u0/R1BKPulOpl8j9IBGwgRncVMUK0mn+H/KASMhim+b3AKk77vwG7GaxTHTepLUv
sha0TFHEtMgWQ8hNoHye1NyqUYh9341idXpYTFhfNZysVT/DBeFWN0AdHwyocG8B
mdHDiuxbk7MdzpDFZCa1xXavBcAGGOWSaA8uyVaeZWQQDoTXstY+cg+D+xaUOsAV
JUrenwoXy1Qo7A0q6vNAh5LY/rtz7DdaXORGNtEskux2rM9XnKdXGldI4y/4+epD
PtNJ8Ol/5DKSi7wFbCnqkt3hb4VIg4pm6lHqUDOVS9dp/gpyAajUY8ILakY4UVNn
557wlPsAqIIXcPRrq4gEqHeAq49QiuOx6PuKzPWL8L3XjdIdnvW3sT52C2huGeJ2
s6wQOHuV0PpRTuldPrNjeoSi8cQruuPiAMGE7s5bzMe8+Mx5MjHcMLyT26C3j0ME
g7BtE1XRNzABLhoUKNQrxBRPIDPkH/juxp13+c6BFKOW/WLQ75q0Ojov5zPMsnOa
QLSPmolVzC5XsZ2HpuA7GEf+4ailvnmcXo9/GTuwS32JdiihuMEm9zRalp1BbdbN
S9ZYfgAi+1BgmuL5TXNrPSV2H7+eepBWNB8uyfB8G5zof01OCOcBXE0qTp4LJKS+
UgCDvWtTfPGyJNR/529k/onefR0MCIFpul64sNIea8PMn41djKh30fQSuZXSwihr
BgHw9WI6XpnnPLwqV5jWRfbhx/zCS2W6ELxplZVqUoo/4ICzYi8DF2nnlLpw6BXV
4lww+iEp+W1YfkQvanP8ANhEJoY/pZ2dM1wCAfQP6GzDm5UtGYKKD623qH3tQ1HD
KyNJ6+jmkuDqtrGid/XJO9dq6jwCIl7zC+grpbXEnTvJq8XxYDaaqcqdZz/JdzPC
WLxehRr9pCczAr2H0ciM3+cvID7zJXtGYXZq+76Od/Lg1X9A+NJ4M8m2w9bEiP3I
1CQxtIRkqlJZmaAIQYGk95AdsIBwL0Ns4WK5ZTN0NgA+YxlkV8S8a97OX/QthKxx
tqrRvc5ZqftOS6DCx7iVgN3dE/CVG+LMiOc73gJSxpyg6u7TzPatCdUZPYIZBDxY
Pl/wwAVbzIxrtXH4oeZPZfhwlDMYREGzjsUpFLmYjg/Lk9TNPV++fau4cYW1pC5b
SWsgZ7RCSNiVO2UKad7jI7t+UIybbNU+56865gVyvYMdS21g/fOWhSPdAIMybkmg
2h13rYOShydrP60SemTm1idzbKd3H3xbZatPhX7ytideqnw3XD6NFLTvQYz16E/A
4v57ZG6CobPwMC+HcSmsOFtN8JnPlGLb7YHOx1yShRgju7mspCfrvdczYfNU5irH
wRdQfizQJwB7RCcc31nHlArteTfoGYN1rQLZdbT56ae48lduMb+vYboGR+FBTAuA
AUEgHhPVLrDO8V3kU3RAdWPlyiz4w3dstHEXoh3boqLmRR9o+0ymM11QxYYf0dC2
UEmbT/EU4/6FQLeJBt3yx3oBgLNlkG4YTmb0jfe7uoXxye40PmxfoPmSiay2Anj/
4ypojG0WWTS7X3oghtEK6+KPHwav4t6Yk8E0v5B7VDDLhXGqMMDnz2vyhR8ZK3qc
oT0QrYbUntDTaEDUhVkvOIxUv16IUAWDS/HhFPWkzbxpnJf1F+tUHC5RaiC8KpGE
DowZNeJ9aNNBk69cx9HrTMUbt7f+BBjzvce9AZvTpFeRuQ1bvhdDJKkHukhon+a/
HKaQ5/fLrABMWsj+n45EbDLMBg5GFbrRRz7mVZA5dgyrEukzt/prqClra2IWl5W/
bE3ZpcxFja3jtBpfz/KGJx035fOxmZ6iaiLNzmKk1CdobwEUob/8JOMXfPzpNPNi
OQ8QczhEZt/woXxQYR2dSXGb+IYECJyVBIKwAv9k2ooN9758x14bvlpYheaxTv5V
E8as3PRkL5OgqFh2FmQ3vTlqzdDyd1Ln3OIY9vRuzd2IyI0ZPpHewFbT5XKB3+B5
EODZtXZCAnq+Kl+xx7THC/leUbChsFXt64uZh2q94d01hDCBzoyvQapQlJ2yQhR3
YZDMh6YuAnl1GjN/ECHZpTA+oM3uZkDyq9qff9VnZNAJMIwlm9/DrHalWBaXKjCu
DwtArKIMK6bKsEIP0rOzHSr9HmVggCVnfPnBJUReiITLidDihkDG4q6r4v3ewrSz
ZMGS4+ceBjFCeR0kHW/kUqy3nv/MJF7d38VTGa5k3YPPixekfhCI4mlP1dK/7NY0
rDecb2XJ4NmEp1TO+dCPW7R38fN/BXEI2T0qhjy0/uZ/Hn1NJF3LQG7B1JpcKrFc
x0xj/9a7YOeAS9mLv3PM+0FxEMKBC2NsFq+AJ2Y8nE2LhZCMFoSaoCnqnu0NLKZR
i95V8lvSVIL0B/xW6+bs87by2FLuYuBtJ5EpMjbBuCkVzCBscr6uzcJMVj+lEadG
4JaRuE4sURNoMh0g++IsuLKeznwfAlW2KFEpj9PhpjRCX8Ol8qE+Tq+CSxGZNjfO
zN9bGzNBxHsit+MoOc/xBlClbIxIkb4yIVImlVKU3MdIfn2+nbzN0C9+hcnji2jR
1/+8Krp9yjqte2m8LQugmnzwf2lCs6XHc+szHlnRpx8WzQnWj0RdyCGtZxJUItYd
A1IG6tWYpTW6vlfZjYyg65cBYI+taL33e1w/lYN56rxpNWbGHd6XRghaFjPkTDnP
HvTtE4DL1aPZb3TIeYdVntvMhmKrx5tJVcKynL4XGUi2H8c48RPGikKFF+PoKBEF
qQFlJRUysupXl4YB+dJf2ARQv2C30c0BDuYph4vSmoSPRf7Wwn0NEkEWI+iF8886
shOY0qYYiRdf53kSSUXWKNnEC1YyI6XZl5vY4tu9V67/mgYU8FI7Bl6EnW8DUFrr
QMHWfuccrJIYdz60rGQLnoZBKWCWLYqjihU7LoWTOD42kJPqtzVGTl5CA+F00t18
MuxD45zmuD5VIEKLyDpI64+vu2yF8od/G4bup0U1QKAyJmIqkx0oz0HBpY9PxRdi
bSXyskAH/g7/FXJn+rDPTUNowHynJOszS1yy8Y26c666Wh/hbyiq81s+B8893IFt
LQ9f5M/fZ5MMqORGzqjEx/56KZ4eBiR+deldmZR48aVWDu2O614LLRRKLafL5ReE
W4kcHhYcnR/x5orVkQG/mApbSYFYwB9mkRBSHMONTevsBPEuO5wW06Vg/ADVHGBp
RtvabS4+m4IE7O+ModHB2TjaKJS8ONsB+xoxgx8qqd9B9EZbBwiYRs2WDF9wnAxB
AbT8lQwK6hf4xNwqcn+GHCpGWJF5ELwfV8pbPZVta2Z4eTlrTq/+0Ne9GpM7f6YQ
pEOW8KfJ4GAfZsoJRAgrRSoNPBXkMxayRgCdJ3QlCr+5E46foldgFrvauXRkEFzv
BnIxFoy/TcLaWj3fkR07ISIXblYFXmxP62gg5PnodU1Jkbwmu8lYvTCkG7yszsYR
MmbExI7n+yAQmH/3ZhHX+6hWNg/UH2MvZUh0UbOLmxGzJh6EVLZUmIPWyPb87U0A
I77wLB/Vlknb+oE9gJ2djKNxuB5R3ZxdpLYqZckTmmbROElSzDP/cr9fq7G4Y+kV
NVCFOq01URH9Euszb35tomKtS2w2QLwOjCP5yTOaTBrNdvvaQcRZkY8vgfNTOV2P
u9LzNs2IFmoojFHESPaOVnnS3K07idcA+8q5Qqy6R2u4o+8BtvQibIDAP4Xfmesc
kM9C45OJxF2SNVD9kHh51QMM+z6wNnAjPh6PMIo9GRiCBEpSJewHbiChanjRzrhE
eApYpZOm5qWa6rHQwzGzPvXZ8UHlAkzVfdrTds4RJJb2NU3YuhLJHVWHTwmGDPio
kB8H7SsZYUMz5ys+Tio7f06aCyxMw8HX5oMS7ezB828h9ygkazyhPCXE7juURaNK
QiTnUHZ8n/Pn5BYc/P+Xaei6HSOy5AXouZYHbPYeYHEMPZvRTddi4+6jSowhmJzh
Fpd3txi7mephoZpXaJTlOILz9lmjwVMtor9WDV0dr/Y+QDKs4l/CgmrzigquC4/u
fD+kxVNOmypOm5wYXCjgdTEbIWeFGobQnokJ7N1ev+vFZuIn5arlLrwF7llOm+zm
k6DwhYwQRDcKDVtP9Da+OpnBenV4BDelAyI5vRdXJTtUraASjmdHt3XBJxTQhjJa
pTJJkzLqt798Yx+aDDuK2agdYntr6UaQn9ukQ1Y5EX86lYqE51Qw41pta/LuZWfX
rwacLyvxAG9AwkPW6K4fhEFoGCEgwSWBRmhDVCB1CZ8ROQQc1dbdQ5RwJvANzM1p
ElAfcU1Nb/ArJDHCBQkArnPPMwvZJ6BOYwSCzWctWRWUhfHIWtvWuGChkJd0P4qo
PefPi2vZgrnclMZYIDGD5DyRXg//nEDeIdlwdF4fnLLap+wLQ3HophPaWJQc+7OY
1MJCK16Qx3QXFqmsbeo5jzbb3Tlfe4wohuZPrseCjGyXME2QLoVHm8NZZcaSfsKY
28hyXtRmRGSwhdyDakgVUpiO9ulk2fOAQccZtmJlyL+54qy2HMJuLFRkIqeGUYvC
ZKcm+g7vHRmxFwBTJ/W6fcm7KuVbH5QXE6rerUMYN04Q0KQR4DI/dU7hkshxWvGD
lTF24U4arAUXy0p1YKkDb2kMYZG86yV+YC+cf7qDcI0YxKmjqPL/ei/BQywsgZO/
2remCBuX5Hc2NdbyHo4x48SIN3xiOB44/bfrVPNlA6pmYVVN/CGYW+rA+FES455R
JEwjGI/8PeJ3fdj2Vgq4FSyWSX0eLzQuiEu96EBXCs1Hscl0H7uZmhcprxdZ01Dm
RWRP/y4inRYPcisPAcRXpaQKD7zf2d6/myy0AkmHXPUaqbrcwTTQd3D/Ki63X2ZL
FSDPRA6rQPzjRF3+MKcnY7v5DY1B7E+ivCQd/amsAato5lqPKD0vpNgEUf/KArPB
6/BMAkoAqB9upreKW3UaJVr1iH8j/Y1nqCP+ykBUVWA05m8R4gsOxUrEkRfuClez
rMnumFROzUUkgL/fZ3X6hPZ72B2WBY9oBefE2M1Wq4qoF5HQzIk8fuCO0h8ieGfG
XU4Dd6f7XstFJVZwsgzKJgrkW0955E7fvYs4h3K+YjrcD4C1XPd9lGIhRN/74cIk
Gl5UtiXYLIWe4cNLgKR22dWArLnHcx2EtNDl8XzYEPjzSQ7S/sQz8aoL2fYljNUo
mzMuiEkD5NEjR9EJ31MnNlt3MjUYJt2P4kknJ9OndNksGhQ8nZlfANX/xO8C3Fby
f872lVSv0NF/RD/8zgIAGNrcJ5EkpMgxJNjJQlFPuGUfIJJKAROlpqAcHjBK+/3T
3uJmwbUmWbnx3yRyijkKJ8RGCn9Mu0eF7tkIXehRafuvitUPZJDP7Ip2EjWcx3qZ
nLcJ9HeJqMHKdNehosyGZa7cPaPJ80vKp5T79mhz/ZBiONzn0AsPyimqEgwUGfQK
QS59CDy97CgckekyABlsu4VL+PEDmvuttx2VINMGyifj/26ZlNCGdaDtHhRDBVAm
1CiL7srNiP1mEqv9+vq4HW5EtF4ISU57afP6dqAF45uPMD8/g7fEqtJw3knX+fKl
AcX9AfRtcfHNevxaB/CxrqvDr+8G9vbEFTsl5WwlH2K7TNEyWNUdFoEjRTxmnZ2T
t//Q0dnDAgKTvtXmOgXLbADuNLVasaDomrmi58ETEcADBigNUj6prdVRPvdRuJmO
19pFsPOhTQT1ejP/ZioWTVgBA6z1rCGSdD9KfrAbumYgGROgSYsuG8hs5hH56Be1
uY6pilyWcb7fyN7q3APbl6AT6BntI4X75cNpV1aVXjrRoDz1ftb1qcswQW+f9ixy
2e/59s5dZXyIfwl2700tOiRVHXdgNb8d4OKVPQyP3hvISQLHjUlHGV811QsQzuxi
/cevucBRN7HTYI15tRXrQiiCrcQeh681sAl8mWWAQJLfOCIT4c8+Lgeg2RTPwpRu
Juuvhkw5Kdw7gJL/lztHJokK763U++RhLt13CyhxX9kjYXpzmupxpyfPJUK+K/HI
z6fA9Gly0Vs2kuH9mq5CXjoQ705wt0EIZ4EpuUsWz5A7wgYlL/RVxerdGapm6LtA
mm+LN6qXAO2SSb4lv5PbTjHfinv98j/aefyShPRToF3cBPuxfrSfEylh0DbklrlK
H8EeTTjoHGqG/Es6DACBP3cME5BDtI50dBdbeSzT1MznbXsyODy6KLMBi0U9dXsY
dCDams5jN0I6IMccCRgULvyDH1EXRle0EfihVFifv3wekbexmIxY12jbIZcgb07u
PZ93A87dJZjKJ4RsIMu4pC6LmiGDjiDgTJzylFTnV0+11r0x92QqWaaV0iJZrPIT
sLDwpVrC2JrGUprfM9qWsShHP368X6I1SMQTN2NTZRy6V65YZfPrlxVzjLaPlxch
xKIuullMbv7rPytA8pa77sg2x+n5xPUSLX90kcP41vOj3QkJ7pBxi2lvuJr57+dY
2zzD3qDN0bGJyop8gGvQRL9YyVyUbIpmpyklcoZeNftZV2YXPx4Dap5l7XT8Jk5d
F3NhWtHueekFWxNKawtZ/6i2iOWKiYAQkRgCEiID3v/8UYkadef6Bho525VE6UYL
xUtKDYt5kQZD5/EbK/2OsDGZo491UCjH680Jg5cTgFaiSqoWdkUUafZjAQmABuIc
DSRskSr7PJPAFyeXOikSX+azqQSpr45Qh0UTcPOGbRioBA8cel4PytJ/lhhAovOn
4UcxT2um9nD5s7z0In4uprZPFqvVYK3bS2LSdQ7k/dnywDdlYf+wnVAkVXpuxZ6y
ylfeuHIQ0NJqHSkgH0xMglpSUd9sNYVGiWT0Mnj1SdS9P2wRN8o6dGmAkguM7+h6
ca5sQ2HpYpxBGwRVUOym38s3DJAjYyV10HrRfVn1ASFHxVtmTj2LpSJsh4HKlml+
VBex+HpetYuSYl8MSFVW45f4qgZSq6m43IKWKxKZB/NdT52ElXpvUhiXgSLdvPDW
4GaR5HjfYOMZ7iQmKmJmzw96V56wfYD6vI5PE2vBPCNHJQ2qbiCWjSoOpW7XJntE
7U95EPv1lt9tRDDlUb2OePSx+1fZA/4eOxevRhSe6ZRDRwQLuRPxzFg9Da7trl9g
3+P+bbpyTgMD/fKA8w2OuCeaqVyYBKzB4oKzJaggFLufecFrF6lw9fwJjSdQI7co
sjV8YSxweAj3WX+VmmCFyb+mVXMrw81swfMQljBSe6KTKZS8QmBdKxy5BAc//xEj
JT50xRgatTzHhtTXNQjq35ue3y49/zroC4m48rrf8vMVD0+y6LY+OBLKwGk7HiA5
rh1RLZZ9XFSxI39qEesmHH8Tz/tGh0m6AvPsi3vMK1exsF5WLO53xeXW+s9GSVIY
euo91UiOVR5vdhzI90TalekenVCKfcaPF+8CX5iEEpLNTqYSmqQ2qBC2Y3VcsdZk
H/ksKxQ2IQUXMbZwWpoJFZa90EYRPKpjVOxo/h2/FUzWsvITEoOA/Xz7XLasL66/
9zddrtnmAsAOABagaNNrD9e96I80QvQYleFcTWVGlIurkSnhKO3cbSFb05kaFHPk
Y+5PmKZ+FcwxmG5lGsFtNqNFx401F8MaXfWA1qkKZBf/6LI4q/+HPuim+XIOgWH2
C9YA/oEk4u3Cg/qqxHShbzokzDtnay/87PcmV9n5jgyWPCqP5q623doRR1f3ApOP
guuV0tmU1rTTC1A4fKFI5omvtYPOq1/uTL1Le7L9FTaGQtj8LDXXHeFNxHUt7qyA
05zTqL4a/WwfjNJP6P3lS2wyzH7qrmi/0jcq26yjCWjLLyot8vfyFeCY0LRh3ikp
/of9T+Ueht3PYAf8UbZSiFXIzAhY7QYohJ5aDcoNSU/Q2yCQExGtunmPcqpfAIVC
XU8spNTun29afYGnaxoT12MeaFt0dJ9GQydMfryoxw/EoGhFbwBNJMZV6hxZhQ22
VLSp8LDZ8LBHCOJrIpWQCcNTouyj/+O6yDMAvia/m0OQWFfDqmEi9wnzVHvszTVx
SEwb+YY9Y0oLCOFfcVhCePNmo8Kk53zT+PPyt83DKa6MKrt/c5pI3PCZTwymNv1u
AyY94fPtaLLpLDDoEkCa4P86dgyvdejWNEv5cbfseUsWt2jz3EGA3IVCzK0Fm8WD
wgeU80pcSb0BCNUDkElP3cYoqKjxKy9Ycc/493LXPfbK4AiORNwuoxws55JhyaB4
Pmno+74tYpTfchWObZO4ZOPPwJjh8YaGLmZq41KFLL/1b+GwqiDORKz/QbeEx+9K
pTKOx6dPfWg5p8B/ziVnZu1mVLYzoi5PJytLOhBUjQWfEuHl2T23xJXrjsjfww86
JpjeXy8M0MAVZSayRzqxzx6yzhiS8BL2ULBMrXLURIABZkAnQX1GXypG83q2sKZ4
ob4xmans6qEROWNeZ0kJvliOmP+0IY0qPFWuBnfuZvmDjhi0xNQU2XhB7hYaih3j
vy7zm3wcFbS2krPhTDda4TS2Law3+uxfHCZE6JE/6lBwJsiyPE8rfHDYL5FWTHb5
0QHEqBWaeivKcccN/7Te+doNkMsiWrj/Knuu0ObP4eRF2GjJPmZXPAFhjjf/Roln
x482JwMlF9GPD1z97ak1shvTVi5TVZ2z/EQkeyiCAal3TYEw3mR2YTfbBRP7L0jT
8Hr7I4bSH1Luf/ZYhrI34ICyi4AXifqsoVjFwcNNOAOUBKeY7h63gPs7jK6kdAnp
3ShCkj24xSg2JXTY8iN5W/FCnBRlCEccMqpQLoIeJFWBVGP4qZ0OgP1rZfKVBOwH
W1X0L2BeH4oSPvOmJxXR9LJgjhCnfejtgQILzRHP1I4wT7xh+C/Jvd8mM/Wnt/lx
WwihfBbbbOdFQ6wnrtVSt6picPQMO9F/CV6po7KDpyjfbXEj0cskQK8hcBJuPXfy
/1cfVGtAiBUMHAdartiRJ1SHKmrAkRVLC+yJqZvi9MdxjYtG/1GWNWODSg8lSBx4
6LNPgzETYVZfJZT21V+FaWuI7k6UE4XNiv7sfKHANPCuXNe5yGkSccTo+6ZM7ZU4
QUdvdb+dM8sAKOIk0HnPsNhhNr5HuQRH1hu06qtMkPp6xN9XzDCmPe34B+8cbPqk
5GR2CRRnQWjifVygCtzvQMC9jCze7h9QAAFxdL8mj63uZ27JFRG07V7hgZlcMzdK
LJee3ev0LL8NBJanmuWtJVH4jI5Un6ENTmF5+hh+trQqFzBeqb0QaFeySQ9+Br3k
GQAFlAGzapmkAOqmI2cGXkU4DduAPGc+i/yJTTC03Nq2WRfudMLSeBoWqeuSbVyS
3U+zHf3seD3au32LKPX20zfqZSuxe6/XWJiB6/RBtI7xItnyn7q3kfkNRNX22V59
U2oOMHIUxYCXMj8iylek3Wj+6UxGlmd4XF9HtWJq0PxAoG+p1l9D5K/yyT8Zg8Ev
nK+3igkEort+jkwEKbkEuJ3/PNwBRWMCIS5U8ysZwhkBaE0MCxpM2ND4Pyl4i2yH
uYnzSTbm5OKdj1jXTjsf7A+hPM6Wv5oLPFcxxmQhQakHBPpIxDEasnqwOfrE8Twl
1Ao4iW3piAijLbwtcpS6fSzmLgCwDh+0VqB43wYdZzY3SVuh0TZqOATc7FPJ2m6o
F1SYE2WLon4IQ/mLCXm9Ae3cytDKq7ls2hskBuv5oXT6bKUb5nw01nd4B2TCrFUo
H9tg7wDmtu+HpJH+RHroaiyFGgZ6QGH2GzyiVlidMX6S06JrwcTUr2MO9B20swIb
2oxv6XSA2u/3l3S1kqvx53zpext6pOvWV/MgwCVuB4j3gTbSNhZI97q/XwPv8oF6
hGtn35rI6TjQ+PNr6tULBV50aY5yZWch+WptcIaDhGZ09ZCDrC5oyUeUIR7SOhtl
ZbCq8r1qhsLi+miiTFBpTxRKl46SVizXfcPw6gsKjreXk8liOTZCQNmtlMMr3oe+
pRUnvZi0K0gpgXCxCrCS/MQrGuLldXDnvKIWN063+wyozSwx99OwJa8hJ2T1Qluc
rR5kn+rZ+0hm1cTdx95u7fCvF3D7SbXgYIckjuW1YEQRTIbGB2vPl16G9ZNCumDI
3XvQYUZrHfngh1AsNVkjbmBrY6+91hBgo+TVNoIhyCQI29h3yRSzixlOA0YQb5Nr
U98m4G0LB1htbH8OaOYcSdEK7AshKOOWCOc/NYk2H0wTPhrb83Cl1sapg87QGZ6u
jvAUUSL+702ls/RJN57Vx8qfE8YwJ8XAZB0n57yqvKJNCJdeEiYOH0ot1yMl1lTh
eASD/o459fRpYnk+KWKOhZkp89Y2vXXlEmuZYVC2SLHStXldKlbwAtDP8zJ5/yfX
t8ywmGGx9q6VvsT46dLxVRst//Vhk0z1jNIapN/exkpe/tptB1w2nPE7gC6GzMLl
eS0OPGh+dmuJVgWAAqHPlx7MqopEb+Ni2TqAnV/eT/dA15duUla01nTTtniR/csK
F2DZRtme68x6MBsRHIZsmjuRF0ep37bBMKZ8fdFZtKwR5IjVlDqBADXSTe1DWifi
+X3jb5FtL/mb5B8f8gO919mCgi2rPcSiEAJAUp57NOmFbMqKQdnMSl49SlltILkM
tCaQOy8WGKU64/EgdbsnpY6fxCDoVQMisXi77fyghEf5YKe0fVJB4ZNZtO19a/7o
IliX7+Bpg6z785eKGcJ10zg/oSwRetsFecyWynogpiGI7n52C+JVRagOZWvuygYA
cx7dJBGuvhdk9yZfIXMNU6y+VR260seEyvA5hWPatidr/NiwEiQL9TD2eH+nZgNW
ACgV1o2naZQh1JhYOKVQlV3HM1Wtp3v4LsoGK02QEwsIBPyAytEfMXJKqaQ4XNbC
ShPSLLWnfOycLZjbWEvpuap2p3KnPaCU2DikCP1m3VqlSfyjR5Tb/J2m+s71eo4h
0YgyXJaVtlr9BC3acWaRiTC5T6GglWhWEDNofHbLkWeeXfZKU12UaWcrBsYnEmrD
zq7tH67J9wv0W1atuXPz2PVC3QRYfUUxiduGPfjr1Mg018YeqLaG2/y4hsZ/JRo9
Quzy2syR9dy0Pwwoa7FEp70QSuGUF/yeZtwX/gFKJu9iOCvkA4GIYxx+yiSnyu2k
lFH5ICV7QEaCCrTX9PUfwwmf+pfgP7p4N0D9m/xaFSdkmnPhFSxAILqPf1nf2MVB
BJ5KqxBR6m5pXX2Yu4oQ3TKIRR+sVpbP1RpLWzic7QXRJ9d2EskVIBQUrNW2jx/5
euu5/zlsybl+B/hYE9N85k4stcSvtUNKgIrA8qRutryHkLiNkYq3Z9WDEYpiptlm
WSbtTkViByOb45+PWh22A5XJGMthGE94oJ9kzPsJx0CHzADtmlSoRRqLseuefXR0
ASLbPcun5gTvijjrEXGUYfTfvbS4aIO4Wv2r9S5A0+lcieDVM1bwcl6sKrdG/u4L
YapXuqbDuWzIEvlr4712x3170/0nN/AsFuwXAzWrCkI/hSsqxxNwDgXVIDHlsswv
xTfeRMAL+GpY8f/rcddm0rI8agUGpfeJnllLUEhTP7Ce8qZapsd8w86sefKcLjp+
+1+ocJ1eYXFsgaBXy5abAvr0Z1Q7iPoxHRZJ5e+ICE7Pm5Vro/ft4fepsaV/vcmn
hU7gyolJWl65yh+oHxNP45MJWoD71jzrEMzirKqQWdP6PM9FOds5SASLjw9LyqZZ
Usm8Ljepd+Wie3BIHQbRU9lHEGnSWfFkzr13dKIGJBfK2H5Vjd7ClonAfclTTE1s
vIltj3EOGfLXdiGPfDY3SGcltRYzsgTZvFBUEjb4QV309YxSiQHUBkxy9xgMpcFq
GpSh2WAmZAsAY7upeekPDyAK3NgPmS8Pa/tOD/DQPy9pBLbVkRwRbIA/7GwbbSS/
jtS3/zGrhZUsFemz/tEc7zd4jFZ87rYiG9yQw+PjWhKG3+o9/GaQvfXQfXnOq9za
zBkwciBoR3+5nEc50VO78x6WVzmu+hQw3f+L/vFs19V21wC9XPPs5hDAlZ7GwlW4
uIvjQFQcOkuO/o52xuK6dRX1fljOshpbUxea30ktAJkocMo8QLP7JnFG5pEswMWC
xlUpoX2fz5+n0XYIxXwRnHeAHkCLsrTfs2rgAhK3jlqM90z0T+RcoJ0qrB06k21/
PV3cQr79KWnvNm1iT11WtGNmQhzrOJW/2PTAuthb72dXSUE/t6HQUmHZNhq/bffQ
ytt/esmm0J+3WHbZn1LygkY7XPZjCD7x/uui1au9L6gu0SdCwRaFZnp64OH3N21u
ww/MULdyx3ukwfCbWrCAsOOzqKoD9PQYwfblS1yIW/JH3tkldRCmNaVTFDO9jXpJ
wjj4c270pnEBG8M2a3LbVLi4yHt5kNv3xtQ0uZUlO5Olrd2XyCxqC+nVlhsTZIaU
SD06WgLkp9qyvSIQuWT1Bw511IN+TKELy0WdrCCjC03MWvcoNGyWOjz3uuRDsyw8
Bn+b9BojJ3283QYCHqhqsraENRDAU8rQXV+myB70VSoph/cKREBURnOIRNrlQbPZ
VkCWxhgYtgZDYGeKLBGGxnqcdF9LNKOcQO84Kfi9ezf/+LNdfw/uNjU8ZJHrr1l1
visu0fasu+gu4+JOC8ykth2LhwvgHsTmPBbdkb5cwdA3IbECXpD8tClhx/vE/Wrd
mBbpcTJnKKSouFHnFTO8E2AvTMfJ3/vj2EvW4vhDDeilfJngRxn6aNjqG7m/olyJ
qN8orA/dS0YyoYFz13zM2dc/WIfVhhMhn9XYnS+G3Co/0Bj3YPSjsKnvJuZLb1nB
wTDhWmvwtaeEo3o6ilS7+w9B95cwQ0QMfLLS+fRQ4AM6MJd4lPoov8Etb+1XldiK
bydElVAsmIZMYsVKSDJ8YNLsjy3oyNvcXmgw52oJ62Ynj+79ueLqbf6DCqW8wYCx
qkXTuaYlPrLBaDwU++tu008QzFUgEvik9UUwDVtbjFIRdF8y2muVDqvNyqlByWzj
dQqXBckzq4g+6qc76rF1dFl0ADOif4QAaC6Tz0bPX49kQBez2RaR+pgJKNC2XKIK
LUPak5KrXSh3vpXbV+e5qGoln1yTAyJ+AbTSx1Vmo/xF4bKD4KnonFhuICTDsyFI
sCm+pdi+bJ3UnsFVfp5u2TsfVKgDkAIC2f0ZvSBzt3z3+qbIsQVblkkg8Zbghodf
qR60lnNRgQUtAoNbp+cbXebk/UJOGEWrr1Gt3bTozAklsFkJHBvlWi5eEPQenjq5
pKEVkp5k7dBMbeYOoD2xkoavgWNa/qAhpQGJtTuWqR5vffLvG7O9W0MyH5r3xR7q
rUSz1ghIuZM06Klgxx5TQvThZbiRWkpS8s1NmnygV/8Xnz72iA/tVZpJnAAcWWQd
/JmkreIUJHFTYjrotbqBoAo/ZMRdlhbuqhiL+21r8zB2wCAmUa+QbGuzZXKb4uhv
8h4i1WEF5wpdX77Hamju0fe9iwyQFSe83lsxVeK2k14BgAmyjXF1l2PbahONvYC+
LPW390wRVhAh10L1D0R2xc/tsfjDbteY+Z3Ueuu+oFk75RjuMtyxjGp1YC9lDzit
FK8Hu92VdRAwK7Krryu9oo4nYvl9w1/1KW2hw64t4pEFEurnZvoR2hfeHklr/m80
U4/Um/nA89Bu09H8ukyEIZj0gOjuf2/t1IgSeV/A4T7nbnozwcpJJ1nyl5NiaivK
waIXSyLp5Zzm4kgSPxR/rWPRCICa3/jwRKucz9WYKTTipFSb+2Pe+Dqk0DaUcf/a
O8euYxIQKF3EgaRlSOwVCgFVTdIJG3SwuyfB8sb3jHwHFmmShyawvsjls2kc5q3g
jtTAZWtiwbPDJLLG6UH+Kt+/S1ciMolkhqHkyrsuB/wGrFVR2lN55VCyADyX97dp
7FkXvPMhMIKbE0YDsHXpgmv3ifzGbapLnH/8P/Yo2P56YFP3L/Rjdinb2PIRwvog
suSQLkq2BgEStSVgV1pCCAJq2EM4Cpi8cvnWFCU5Bblo5pX9Vv+RMegATl0Wnqas
RTXcpiABKMLQdiKFjGQ9YCRztEyGQzM7QOPfMBDdSR0zoIK7MpZuOOTShpUs91bD
qmVXavumyQo6vKWZuEu6j+aKuab3YDtuUYG8bxIYbaNKvUCMCaThPnaAwhWyhqKp
cR72/yOadCvTdDB/sDUk0/cUMcglb2SKg0jcA2GGn+/RJcWRRodr63E+QixjFS+b
m6xNeM9t+nFuzqw/wzkULPbsaQbZFTX7s/icwTgyWEqJIyQMuz68OfyK6cVTbXbb
IPjW4PN0iW6Pe18UcFiyMsWGuaUoA7u/3rY3/gVVoz1QWHPvdJMDc0CTdZXCsnlK
A/IIjkYMUQTccQnIQwmbdWRjELKmUPJQoVq33+sMAkDZ/pM1q66vi1+f4lizPe1K
HaEPHmCp5ez3FfgCOxE0zlVPDGUox2TybbBzR9Iw2bEuoiJe4x9KMjtDTNT4bJjy
wZRhNhQ7GNGUj5D5A2CjGrmhxD9UYd4Frs7SQGFJ1PeZ1YyO/YhlUcTbxvQqaqE6
BUXf+0bQ5i0jd1CzUCQy+p2zgkEOBpa9aW5kFxeGLVNQn0prgZwBoQS61sjBvZwR
Mj9PQ2Zg3ZWD2E9v12/+EFxF1Nn250JAgRaYLZZmr9F3ai+ntEDnmVSVvMbMZTOf
wnsEJuFdZ6/Efe8NC8XVJ7v1IUO3YmMYOy6wZOAZcZggtJkfI7QF3I3rAS+oiT42
PB4yjkJNDLE4LOfw6kTb7bdY1l3gEAzEsq86xi0t7XfH1nVhE4HzXWZ7TA05Hyzb
Em+IZU7dQXhO8rrcbhi5We8DLyGXkjrZgrG5lECd5aIBMv9HOu7QiNwNBwANOA6W
O2yWQx5nSptBqMRMeq8wPZQ5BljBRl4Y/4Yt90U+/Ya22QeY3Y7ike8hwtZgAGbv
jJusGmTcgXzoCp0s7xaULcAcTZI7JeJ8KkLsDvo9jx77EzEaCMIzP4qq4PeLi88T
QuQAvNx8AyPoQvJWdh8IDbcnGO1KeDD6p9BWFN9BCyXE1TUCnEJ7q27sGmxqEQ0+
cYLnaf8rMBZe6UgJqr4bsVoULklDaJL9Tl0sJSuue4QVtPkTIRylvT9KHGnGzIvE
29KOMwaLDtz/vKx+pH+zKnVRTWflBgugzefy+iUJ4QJDIikHNFKHqYKTFPvm9HNz
q+rubqn9sS/tEAFTyMCQnYl1FGsmI9FxrWKiWsLwPD4zjJJUSgPvnFx493enYGQu
JMyrQVxfQXXLtNXrWMUXf/wbgi/tC4uqlxeQsix0zmY8av4Tr/N1i8T6B3fRdrrw
C+LOoP8tF/Q280IaLRG/8L6yYZHjJCKV6gJujX4GfUZtnIsLkdW+iO/XEwzb8XZY
yseBE02dRtRVBHCL8LOYMgg8qGpD/13d1wM9J7hjEVxMD9un53VdCpmwJIs16sn2
+CYkiGOCj5B3jLajYPq2zU0fjXxjPdB9dCuh68U3geZaO02fRsjuoJVXdKu0zK7Q
L3UMBXMUgIWbUuyflaFXR6XxeQPTbq0PYoXbrNFeAU7dmv3n0Td6O5DlhQRRqCZZ
vGQLS722IAcUdnZGB5UrApbEe9iiExjIkhcKvyBAi+4bX55aVnKDvyE4E5rfV8RY
lEY2YfWTQgBMZTEvL1XAB+k7IpxcHB4PazVJm7fckfSLGypA8SEt+mpfcs3Efznf
6UN/cUg0vZnmnPds+GGCMhO6+qoAzP368/T0SMigAyynVyxu+GTVerX8CI5bS6L4
ZQjtN6ZhExVcb70XSZkGU9dlVOqslJFJZpmoBWo7PKmbJLpEd18Y+igRtcnnK/z3
IUG9e8XR3SDOczUWGxkcgC2KQydxCx1C88/arOQmoguzKLAYxPsaLQvFtJbSoDCH
SToSkeA6J0qx/Hd0XzPI9zSGoYRFLRjpMDrlkPqh5HphPTg5YrSkBGs2IgiyW56U
aksy6TpVvXzaIvHCtK8w/ObGXN1zogVjKmK3/3yPp98YyEFVFRt6kpfH3ZppSa0T
8dJB/Db2o5woQ2g4stXP1B+Ev4FxQtvRjCZEZF7VTeFn/rSGrl0IeAZRbVSJAXdS
sMkiAaGTu+1+ranKY3LjU7AZIdfwvIaOGa/GGRLn021wwdVYx8v23s2ZsSSQSiY3
OFZYUwKhlOZUiCfZXgRCpaCEycgVc7uBplv5Rn3O7cFcLQwB7i+2x+qjN+h9rI1q
8ldv7IRuQ1Se6XjDApITkER9BNvyzvjpXCjX+VTCsuJdDU7kD4LC0J2eKpbf/9X7
UCpJaGpPuAB0PEwPIlpVkr8gTavlBVU7iGhXbkTjaE6LzVzqtGotV2PtsTo96nMU
nOR6I1fnga/lIubfIwobI0Kv08R+PydfHXcXlC3kE7Lzs/UG4+8no307XVBIjgSw
gz6zfNqwX1+Pd7/338GTg6/5u6SxwFNngLJA1tOf9LKM4ohOw8b5P4H198laN6W5
2bY3ECIKjtQ+/TX9UKCsC2T+pZIMofnl0Q5PuR5ZUvl/trhkCE1SQoAlb7Pbwhs0
Y9JISsb8uMozWzQowjYVHxI6gK08C/U0j7JbjNkUQoXlsNsDDxBQq9H2RLP8EtlY
C0EF/UK2sdts6HJ+VUPxoccZOsU3s1snkFdYQnvdzXeUmUkJ8dkCKY9sS9uHk8FV
uncNncsIx19tbYZhS7in0LViiYI238D56xR9MMtMs030PAIMdtx1u+Y1Wmfu6xqE
URMn4BmC/Hkd8on4rIkP9jRxI7CC3Z16Kt97AwO/1D6+xcnzh0eCvwe7e9xkO4fJ
RId8JX2VJzLoZDEa5YeR53xToT/sWGMPj34I8KYNBP+T8AjrvbJIIPgFWMoJ2Flg
fV2Pf6/QcvOZx5V8i8mepQA1NkkZwQvKXrw3jGnvVMnb0Llkb1fuUg3O7nsHxDBJ
Emd8f70l7NixeKrzycuqLBAUk9IaERiYNd07OdavU/d1oT80bZBbjz/bwT4WtOFU
x1FKZvCZbgQnC0IQD8Pjme78NmLoK4WY7vFPdla8suThKAthFAoe2oUN54MRNfNE
Tktgos86XoNX7ZxHeMDp3DWXqADLhh+zh6ViRK0ZfLP7ninYHQ9x+4Vn7INev0jC
02qB/EsJOCYNNXbh16u88RFXva0Z9sC6p0zM4wqbgo5Tu1GsYecge6uDuObrkB8E
T8kQAGBrAqqPShiSI6Xom4c63JJfgXCcR1xVuwiA7x8vrrwpd8XNhjBASzm04GIj
Pxt4uP6uTT3MEZp/Vif6NJAlne+YjM7XLqOOG7eCqzaVnIP7iIvn80Da7ULHXnEN
CSEXj+pqxM3m7vYvAwFvXVeIMa60tCKnvOkE969Dzhrcg7C0hoCnwR26W9e1Kc1l
94XgtEgyfKDzJyD8L9krlOp3dm3CxYK9LH0P301+75RSyPOVoFYwOHBNuqqwpn26
shPWr2tziW4pK5XD7oG7kD/eHZUn69k7Ic4k8d21/iDSoULWbYwOCYwPhK3zSt1Z
EtsikAabY5JL9gKPbGFb1ltWxF1tiNxDt9BMCjNbuUykMvncGav9NxCOettVSeZc
7QvXcG0N8ZNXtE9HO1ELLaB+Ira1/MBaa/bydgBTaBG+9jns+s6gwFhnAs2WDAwa
II5ioZzUUvOI5xSXW6Ip0jbVMlD7FXv5dXfZFjXxHzsDpTaWL3CdxfSwiPataTKI
yXG2IJ6WdFK5rPhU3NepDjIYbnPaJoNxslRnGrPGm+k/+ZNo52VF+9rhhGTJham0
6FXnM3JDx9XnBdkLkuAQyyA+3kekWgJq4hH+edsu73Q1IpYIbaLW3vT9DvWxeamk
P9ma4eCdcXucmnzYHTKaPezIXDSs039Qkt3zuHbylRmQDx6/7rZY7Yz6WCvhRSCG
vNwAoEy4us4NtogXOC4RD/J7nnOf2bNJW29vj82xOFGuR8ycQHxO39pHq0q+R+r1
ah0kH0ej2rNzm4qVdlGBjB5smWszaorth6x3wzKvLDQosG8NKeRys8f9yIizhSS+
hXGpxjQMb3shJzvAbX0pFnTfOhzTUwxoarQJ/D4q9/nfypVfLYI41dN/U4a8FwXD
rGJbK87sfMUoR+uWkivg6kFjA0NK91dL1osnZ8fzRAyALrRUWmKQS6x/M7FnVA/q
c4srZAQMR+/XX+l97x7QX6Dlgg1cbVr3tbQ3KnaQTmRbarWcGKrkWU5lKuSk3ba8
Jq69I1DqAT/9ce2UC6PeZD0Ly9BudMNHY/LqpOY73Y25dVzgzPpmIw6HJpt1lIA6
wlePZXvtuySTg1DthQl6/b8Uc3PY5hastCP9x7af04vxHQkMz6WEs8Ulp7qWpzMz
aMnjAsFsE1krT1OwyiU2PzEwRexiOyyRMYBmVk9bl/kFAsAkH3cbh8lsSSXNmzvT
+zYlR5vi1EoNF9xJ7zE8CVIrMpeBURsDJZOzImWAj1yw8vhLm6/G6x0eyHixyKgu
5UT4348IXV8TdFysjWKSFugRJ0CakQm76FxSrj3gmX3MZQBOQwezmSmaNtEOvGNe
EiTxUf12i90VuQnMGvOc/P0zoiO87qXmGKAjH6uN7dZdJE/zIVTZ0jcvnnVObBHk
okhC3hzU5c/H0Y5BPlTujNdkmdV1s2bO+M2jWpL5F365Pmmq7HGGfuyBTcz/Kgf8
9RMG0qJOQ4a2/BGF0vJSzbNrYlxvhmglxM831RXYBjUMjmF2Bx13wGWq6WlRi2mA
b8hVH4HV/J/lgO9cqt64ka17YmQdZYRKzHvvsHJedzqwUvGdkx4pWtvOA3XF9GUq
oZKrUB5GIvcKXSI2YyPmPTsqHvbjaW1M85l/g3SDhuErIODpSUNW2SQThPzVbSY1
x7anBTyJ925jO39Yfb1UFQ/DZCwK6EoSByQsJtVMBmyiGr3R9LYZXTs2f2g7DFqp
X8Hw6xH5lPaU4nTrJvcUkW70lBa755qBW7eh4E8DtDVKmJ+1JHOkwuZY+USpUQhK
R+k1BLcFo3Qu09d8uYftwhLSlnTI+kH7GZdalKQrzq8CbPTYmTGiOkGtbTSmE1ak
3BY6xJIWrM1XWO4kjryA5Ni5B5sCVvxVjJ9PCgHn3mk2qZa+q/SV9vdNIBxyGMUA
QSefUe091wl6VWBajO+dorgppHcnZIoWIHtPGIASVwzSk7LK0h5g7wl1QCT71HW2
Gh6XScPPrUdwUQjtbBclfJZJXxWs2NYMznOThVGAV95WivszwN0wwPJLEGlP4NWH
nrOspVhtU8LX3pDb014uR7CY0va/aujuAPbbgRyX2+NVnZo6op1UeDsUYi3klTdk
cFQG3RY3seeUz9Hr5fX7L7ONy5MT1FbhcahsmWqFBj6gAq5WjVvFOyCpU/mEj9E9
+xcm351igavf7pWa9nElDeVGzkml8S+e1VAkteQZkbf4F0IbxFVGtCVwJ2Cup8oR
d/bMWWsQMVe0poyPIF1nZEmHnEPLC2/XJpbBxW7a6qXl9GznB8oBsKshUkcLnn/s
ykFI2Z8+PWoZgm9kjtQaVJ8kwBoWmH3Xe565HQ/r+r4HkDJ8LCVw1G4+Af9atTJc
tZVRcuYukJPke4FKcHEHyllOK5/iFB0g9MneWMaUefzhy+8jDxeUCoQF4I0IJLHb
YKFyJ2lCvYRadYs2beJ4iy3Nv0gIGMOaeBjEm9vuYA2JdAMOLBXO3STLhOcaRCK9
vBULhOZRccrX7ZCIwVCAEqL4z1pXX2HICA+0+2IlKwQN5IXVdf2mzDRcj2QxakG3
bmtdO0f+c+w4W5OyL32MtPwGpbRhUUeKMI8yD2TLTNclQA2ne44yQcusYuJv8/io
xd6CTZCGM10rrdSrMolK/vGOHD1KyhTDDRtYLh/LSJ01ES/QGNbcCXSJaD9z6pmi
NDLGuwa87aoTjE86UlyN7PlwZ8eF1RfOpq7UpbDKfSnWbNYYFMRakVS2TKqW0s29
yyFbz2q1lHqaTYZqAxNU6tX6eKaHvbOMbEwDBTDorBBkyonXZYq+WqvqSKMMjZHU
m/tpkpBCopOZZWjg1gnlLNnqHYZtDn8UbxIXPWQtrwv5sVpSeA5y7oT0sGpg5IGB
kOIL5DNjJ/nLuzZbpkOEWmg7TuAA1SPcJMaGbSbz900ejmRxTduWWKWG4VbeGwh9
Rcl5PDerNHBMUT8mwhFZQvMtO/9eM5ngB+S+Swnp0+U4ciy+O8Q3cKwROQSR03t/
h1w7MDWbC6dRyvSAQLoKHbKwvoUu9F4rh04N/u21AncyXYlZtDuOTQFQJc/OipxG
CknDdbNAXYCSOrm2LDCtVoYCkesiB7EaPqlW7k5sJQvmO2dWEO/LPTLz44A18vmi
K2RYLjUNHayP5Uje8wfq0kNJzyhJW7UyLZ4TgEUguTbtrwgyEWeSHhTNSshKwbN9
qjFoqKXiB261koYke8f5zcuh4e7u4Zc/5kElIWsVllkpsKfSeqTS1zwK+CreghFa
DOXEPaEwyZTJlpYDc9bQ7S0zxjGIWgMKg4IyzSZ+sMKOYg4V/CAv7BiHc56M+gzw
Bvg2pHVHq5DF99rDjRNbcP9n3Siog9o5boI67iaCQp58WoFL5okwkH6lMIxZ9x1w
dWx+EDYWdLCObdTPX/XNHVMej1K4kL2tVV2sfUlnyhJavi1gwoGbnjCPF3U2OmUJ
iN7j4ItnhLZXCgK85tU6WPx1bH3maLZsbwmiSK3rY5fvY+Kfw+c5zmNPpWvlPkvv
JdT2d6nPysnsMqr6adhiR4SDJVapCddvtx651WsnuiLQiQFN7Xkd0LzxDPK5Gi59
8SoHXJJybuy8o34LC5BK1glOsnN47vqm6uQj0RjkxdYujcfq1l6Al+HMkOTDXYvQ
ygOjDv1DBEIceYU08aQlfWYwFEEGd7UauhCdx4SASZ1GhWZH7uu7rZLISmnPBbqi
GQhTH9j6KlKRH8WiWVFV3mWaY33N+xQQH1/zUZTGEVz5pxjjTg5ZYnbg+H295MUj
Zip10WYDV0roDTajLJPiLzBSWbZ6RiCslGmqytVQX91IoptKQhXRHLxEaOZEUHvT
ja5O5k74RFHjpGbF6zBBzXOnHMu4agnf5oDzfyBfYxqII7a/rMDuhwjCAQz8dyi1
C/a8+imA1XltqODKCFiGhYeXG5aZ3VKAA/B4Q/wHfL8oxhIn8dpXL6pL9edgrP1n
4Iyk4NDRueagKLXCGsEQt4eg5+obXnskC2J8rLUZANfhmsGZ5cGLURETjlPR3NNT
Rw8hXzvpu+zuef5hkH0rCVPCPoEYc3F+dUfzFU5Lg35vfWr/mHejhUdM3mdKh4pp
Da8JVLFih3hUEhQj0iZd4EhbeQ78Nbc0qnamik1UVsDmVJ2LZ6SPTKOHBuCwsj/J
TLRPI0Kj9iOkLoB9wFdXrrmMfQ4lUJ8CXLHO74fGH87bjOzVtdYK3OSiPw8AmI2Q
0xGH0bTVWYGnJbMHAQNtVIZHQG+PpQlm78WY8jqp0UsQODDFb7L4ldRZpV1MdpC9
HgXYrldAnqkc0CCGR3T5BCJZ4wYqqO72kriNvCZm8ImZ1SRttkrSQwtdAv3YutSN
9WWUE3sWuDsBLdBnmAezdZ1M9rzqk5l3YA3R4eep4k4R3NixBeDk3VGwDbDGFOlD
XvrSyoZMuwZoKz+8PpFS5VVM3+JFbAJMBZWre/dDTVlhywFuOmDWryLv+YZhj21S
IdYIukesf7WJtoykNBkuuh1ejGHS3FWpsrPx9kqF/KmFUUpTn6La1Fyw6ypbyQh5
cQfcr1es+fcBpUi9wAgSC82CVwoH0TZ/+e/NW41G50wP/2Z4hRCZ0OF2GIttOjsY
RR03CurKsawtnQOALPf04OCISqp3v8pjq0PCNMFeC/XVarTcYHu1ymsp3INPWS04
6I1+mdsuiivoZi+yGseixpkkPMD/DQfoy7qcKraFC5TS1y8SCfxqtTOukyozExIL
JnHVid3jtRDh6Yq7CX+Z3/hV16eyFFkx1dJ/0Ze+iYv/VShdMrD/LGRlXJQ+EhTm
FeGcU3hsX3JA+ljRHmvqMFRVZa9d9KOvYGh6OnvRfUoULWAphX/0O6AzVJeIgCn7
VhaukXbO2r1RDK0giEuB3bnNFs5E5nL186497qlaYkrOoyVRFJiNOdjGTW8Azzxm
tJsFbxGktQgLKAoflBovUpynXYrUrT8EuFrfg7QbtPG6rSk1DwniZpus29ObddzG
ERmLQ4unyv3wtnbSIra2ckCK5QudIv43h0ECuu16B0lSnOB/n2MaFp5EgSL/7Ddw
waluqjRpqnMrDkxTYaWt9XYlEGhJvrdA0CY49TSbOdMIWeiDVoUt2IdxvH9oxcf4
J/eatg9PQBVFphco5jNb470zwE3dZF4WN6rQUUzkJZvplyaAVFMLDENgtUNUSQ5d
lwg9Om+BI6a7p48phHRw21n+5U1sW3sDuIoM/GHcL2qPy9X0zoch+veuOhQsqQ4M
6mXECtBBQqopo1/gpoOOfrIU5W5WgPGxJJPBWKaAb2K5JNRZb4s+Bb5ILTdVFPko
6CY9MG6tEPuSj1ksavUmQnWTkdhS2wFQDW9mAqbsBpdAwOrFkuBm9ieY68heI3Vy
NxB1xltk9MGzH8Fjrkkk56t9GEMAXh2df0c4C4dUdGmbHByTLuBz820ASDmfGnk4
PHKsM0m+h4x42iWZ2Dfp4ctVc+5tVNXh7NA9wSp68WKqidnZgEzmjQXsl5cPIZJY
j6/+xAUCHU6CxN5mWNjBv6e4PPSphh6CmSiMtoJHxOJSy8d4BEKxdfMIjrYXyjZS
+tbJvVdEc+ySDWKp9GL7U9UfKsa8R6Dqi4P+tTZu3UI+Q4XeOCor/VymzG2OpT2S
PM0kBiRQgNC+NEPY5C3eI4ePJGQoIZU6qMMZ12IiGO0rbRHWbGDIZ0lZSc6G/T0U
p6Zuq/bCCIbXlllvHqjatM2zUKNJSkHyJiCK2OfjjX7F7ZyGlgbqbp8S6tIHg9OO
Ywg5wb9hNj0uaXjof9TIcqps05kXjmyY8mTZLb29c0nBLtAs9B6e23/FWIBl2TCj
kymtJgBPfIT8SwFDsu5Sol82DlaP45biW0GiCMFpLIIC3g53/edvk166IZW3TE8Y
yACNGIKPb2KbR/FgeqTrCaw7B+KXSaS+dJX7V7d5Up7TBK/iOZD9xh3xRHWm5nwO
DleVqm8qm9X+vnly1BYzyQBoamIMJ5OAxRJETYkUB7pfh9pXU5XshW3U1Gg/sG95
33Y/XMdifOa7J5DHMp7DsOA5Qgh+lEUAlFl+r5igC96ITVTl/SkBkYXNXTSiR9FT
NRwo36GeCXP99L4zMlqcu1Acr6kN9o8dJp8RsPSwL5J38Jg5Y3TqDGT7QP22F8j2
ltf5Tcl+g5MuSatdb/gJSGaW2kxjbVmEDKMOJCJNWvfiefQ7yrMwR0802stDvMUv
4w4Atbs1f89Ctv5o/ZayBeluIQZVPz5LIzHyn4ZCu/7L8zo4kw5BmIuXIy7pstir
7cR88ow6PO7EYYNFjm3K8GYGqp83d6F012RN3P80G8Bw3B5XtBkNvIq85wt1TF+v
4LwVQtteRwcxIDdvHbzkBLSF9oO8g7S3UNUO1udKe7r4aO7eeQWo67ZmbsqlNmRi
xKzcJkWqVR8TCbBB5TbIk/Z/wLCGkAAunWi5r48eXTO/QzvVazST7ZVjDPPax4x/
W2+ac6gn8h7D+lrswEz5V/qAeLYiYTO/IQbP9JpaMRAufyjc12+qxVP0wuSoBEQf
HY22NiTTd4cljm+9VZ++J8ZIq+SHfw1wV1yx4t/vaOERGPB7Pgxqzcitvz7pMwUF
ewdOT6F1tR0YKWmlzfDMVOWyywoMcxAxkhRkdi2hFeNyyeg35d87HMjKYlsgFr4h
9zFpqwQr5Oypx3glh5jpyZiRQsUJ6j/h3Tgkfh4JhuVLqgYttQr9W23Fyr4nEjQq
kPKlzcTt1v9vdiVFdCn8xAomHf/WS+PzZ8BwkEIU5KFvPEQPrRVlCI5PnINOmhRp
UjwoPbQ5/Hx/kSCP6adVsPuLZEMfutgZQYU7LRiOcUrxuhWQcPED6g2lg19rfM4+
2bVxI3Rcr/5njofyJeD+fFihxgMAry0tcfob1FHhqvaovf1lA7tvmAXNqTgIc8JN
tw+QxvQJfUEQG3wY3Gwe1Avmmsde9qcHR/vzs60CqSww8DIDnMTOSJ+ShfcBwC9P
AtRu5SJxgjQaCKsIqo5pXMeIcQbR9YPzAWE/o5ee3HBzyv09k9e6mAPuXdMm+RpM
PJ9H9y7IB7rbBjjIhlHE6nAZawXw2Jn9lzG+RaZ+aNgNode2mO99nWKebvZtlDeb
OxuKBqDw7n6XrKHE3Y17Va6amoG0JjAcZPlAyvgRfRzkNW4l2F+empmX/0JYyM9H
uGLH0XYidrzupAZO/JQCK39te3yojYpRIWqK9wGa5HnEfQUB2+RG3ML7KjhstmcK
i8et7QeEX2wCtZe6ICn7PrgDP0KyP14or8LauIDcIH2fdTFSsAYmnJdVNAICeCpG
QjElxfWb1wp4e8VffrtdD8hazWBzS/xDfGQyfC2jQmCVMrLhZF2nG4TxJ2k9qb6K
+3gEEN0CBI2LbutlwObq03pX9mbRHcoMzeDeCWtpxM+iMnLpr5UHPa3cfBGREnnb
sRp7zCimspi2bz97M1UO+xDwr7akIGjRNN3O14MEnqVczZvjADhWHG7VBWGEfA0k
MFRlVRki9vYawLKE3YZlF3r1YnclxsWsXLr35V8Niiv7cdHILgpFDE6KRBYYHPdW
L8mSh/Z7xjO5c4hpnI+k72bHJ5SdOkM8vtRAGL//bTtatZHRgQwqQ2qUAswvSO36
1LY1ULa1i3YEffhvs88NQ1wRpgoolhnpLAYAMA73UZ49gF4p920tAf1kIOYq2CUA
hkIbxy3xy1bWd7rWfe77QrvxdfGOvydH4EjR1icwUGJumAi7lIC/EnfdovAg7DtG
IGGPnJOaIyQdT/WhorzdjCf9hufmF4onjUhVHsQiqQaSu1yTm21sRW4ejynRYi17
XLYnYbA82SmBistEkW4tK+mz9umdQaWj601AFlQBynehtZLB/s7dVhaXIakfhoMk
BIct69i51rn+r792C3Ef19XSGb9we4ObIw9EolJc3vq9r9QuUCuNZTFpMqw9Tkys
oK4/+SZCoCh1Sm+G/tresaRGp90BbB8naMx7FZMIufXd2hCrUDjRopNlHPDVmwp7
v60OHN5OxxQFY9aMcQm2bMLA65y9xnaanpG/sWi1D1MyFgUtG30YiHAi8A9dMtQj
4dw7rzo+0zQ9TjS3/pclibTbgaRszcebFTgSBPvM3jpgLwcWxo6YcrKSHPx51rHo
1Fps7RbsyfMt+SDUjJrLVD9kFROeVZB8P9g5XgcrA6I7Ty+fgAdtx5yLn22wFicc
CMYKn36dNYcf3JIsqcqLacI1OwquDY6wm3lHYPndvRi5LR9oze2YCx6y3K+a54Bj
+nNksLhp1lI4m+NHiDov96nKsF2kzlSgnCEzDuY8OU3Qo/rrX6hHW4sPbn4+y1Wq
s7x+Ffq6bL4DAybxOTotCbwwek23exWHGX9zUgxYBwMMZ+BzRerwjXZv7bHHFQRJ
aUHQJXAOWQ/dcxHHMiHGiEJ6MX3bh7hjA1TCiddvClQsYvxOeOXhb4agIeP/UjU6
pY6Huz5aNdFBNEndXLMekHRexoLb1YCnZgMKsoULCYx8fWlfol6ZLOkEcxaWn4tV
3I4wgLHfEIS1NCLSGCGJnNAuf4DfBFLGc1T56YrcDEj1PuRB4uY1LrZJkQUCknFz
86VOT+OUbbKrd0oM/XILGjHu76NxaA73mP4d8PWsccnOyqDxQ84S2ALQWzqFIXZX
20hrLL3bF/HVKhnlq1oEwTbZ4Fc9pnIdldV5Hw61x7VgG4VTVZ+hVhUkzNiDhNGP
dzdb7TYheqaQFGqUNWAUpJeTnzzLlmz9XQqSRzZ8xWivuNpr7tRn1eTwWtpbaNBY
VBOIIrTm3hoPk9UffkMkR6qpcUBaNEooXXC7WrSQthLkWp4RxyN41JoJ+yMHFDqq
ZbkLoXwOKgDMoB1O+tP9S51DnrmK6QpRgpCcTOkTEXYmS2/oRXBt8vnN9NpoC4b6
1BVuYG/XShrrWE40tQwwZR0JDYq/lqV4JJrlkrUxIIdGkvx7oqPcP/doR3ZhspuY
uRxznimdAvY9pk71YIwPWfdyZeVkRbJ2pGWMHDL0My85khxT0U5GehQoHSphjQDo
W1ld6WtWJtj89ctf3xUM0vH99fh85fZQggtT9fDd7ceV+OhmIB+7CxrT8T7vuu3D
1JuYOBoxsj3Dk4q6JAVjaDbvBCmJejaMZovXkcCZrFstknUs93vytkCqevrFKLqS
4v7DPw4YvHYBexiKB3e6wXtYWsZ4pc7UQ58+5PybhSIhwMslZHOKTrJfINIM+dlq
hXzAM0agn2zqX/O9k90sJVXZBTUUAeCT5tcjhjT9uN/4fZCxkJ+cpf0qGBDhzgx+
Kg78udl1R2NK5O1TZLLdemntYkOteZ5vkg6+TMdNDITj+Btv2t0R3ScDVUaWU3YU
il9hHKr/n0ZjCAsqzjx/g2/+BTM7zw0nTkX6mXB/odUhCquHv1Oy0Zkpx+ML2Sow
bQXd/R1pYCUR9RF3I6mYqjTdwNzhgT9sfOaMvjmqQtVCtaZ7VAatZ7DnRjnYytBp
AksGrQe5mz5pu6pnENwnVM7wffeIyjJp0OAROd6Mro+hWIOBX0/9prscaXXSdc1F
+SsjpmE5tsWr4QSbkk97Sjl100CoS6beq31sa2PQcBhJnHFnpvtmHjNsu9FBhsA2
v5UXE9ezhWidxJTQy3gGByP8zV4ny12fjH3ozNLtJv/bFdx+5P9KtzwwnZQVRaR1
hj1v80/zvY01OtJmdaiA1PwedfmmAewTmo365jurfq3ymrL4zD9IeHlg4zuwnXWU
olt9YDdrWpxekgvw86CE45Cde3CTDhFocwg7FuwPOOeubQPWpQSZatFw4XJeyScx
yACwLhjT1jnLOwlNNHsOTRyYQTO6aRVHDunfdIEfuX7DcH2KkbqkH+p/wue7My+z
oGLVl/MP0gk+AdwLhk5V5cJlvPtlI9mL12OXkiuOlgj+jRChMJFO0To09ke0yxGP
Lvq3TajKkxeQrsoRNAHuYXtQUXOa43NBxdhJLGqeL3RwZzlXHJA/Fh/PjSgWHyv9
AJq48JaqtpLO9l9hgRl0NDBzhHh6IFcvgSuBVE8TSzW7N1X2+5ptPYU7QpDKc/Sh
FfJ7ichqXSnPanjJ0rigt9sTiOzcaKhUGO/CX/mmi00vn2rstrkKWLrKT7yDNceN
2Ge8Ef08z2j/rvYDkuj9q2vs8IqEPMFtXuqmLunVQ05Rn2+Oi98M0wpRkzPMF+Nl
0S0ltsc0MHE9fCxK6hORTw9ZnbhS6Nkyrp1mHu1NMZoAkvfDUkX9hlhRea5YDgwW
rGZsEXlGFjB9woVqGgPAuBDI431q9R2m8vXhPBkJNYMbLwf24fgZEQgrTfxHWHzL
eZKZR5RLVgDagoj1avz+UOWC+DFR5e193fjSfo0H28Q7NKvpBMf3xII5ni+39HP5
T+CTvxzS9TrFs4u1u7EIyfG4vxIHHVOe4VQ9rzViwkmyZHeDjhJdajDKdoqIL1Yo
nMN2DbQD/fGntL/zb1tehbiXuNdn/0Q+BQNFmRwxIOKxrq5+FK2CdzGOhpGIVqum
nrWJOXwfD2gVNvl8M0Jf/i03Jp9oASj2bhjpcb4r8nOKmzCfqMeECNEaWMahRGuV
ltjYgIuKZwZk36HGHzMTLLhfMA0+hHuLv/LR0z6Wpbb+RwOZUpd02Oy6N8XPuS4i
RhrXX7Z9uTse6od2fknPyjq1Kno1KTdXQYhyuZdnxnyN1TOIIGhyvOnQuhPOhlo/
QKqHi0sMpMbixvStvQ1nlM2phl3Dy22TVNaL340KvXM7i8pAZm1Y/GGBteurEp60
VySiXX/EKrvFSraQw48lS3WpoqHIHQXK3KinHQlM5jkBdgmdHnmR6H7LYBraswtH
9z1l3bcg9146z4jProewvHg1Xwq2zSyOTW8i9OuNueqQ1Uv7Q9CzvubQwZ1riMLJ
cMxbRZeXIeuBAdIHn7hO7Uw8odSD51se13qNprBISy9qkGvwk86orluJFqiGjOY3
qb+ZV2m26DsVbeIhLsnpNuOgsJuJgNnreMyiLUN6WQH8vUh1QwgtnHf9hIhr8gg6
ki4o8+V9k9DWJ8U1Ud7eFKi7oilRZl1+apFAhojihtwYdJXvdcdbSVuESYkeUo5G
mvfxK6vTacJzyuqEhaR9/0D+I7vS8e19esjawdco9tDyWCI2RLkbP+otLaAOyhKT
OFfrr1WbwulUWVAi9UjyQqN/+sCGOPMezI78zUc4wLKgcbto4oM78Gzs/5mEcoyJ
xsVmhOW1lmGgBVkLX2ViUprDXVKBhVA9UhqzwqWAj9KdwKS1FkCJazW2If+PTZ2d
8170w8kWR50auR2qJirHtmp5itbDwPGr1dlhR0Bzgxbi0W2UiEJ8bf6zSptoLmTa
p+/BhlP/GXtmU6kxkTuxtcgP0JQNh+FNsTDnwxLWDusVgC8wijSyIl4ADwNrCdP9
f0k1p+dlg/uf1CsJrNyZmjmXsxEKZr0nWhAiFhcphaLScRsVZSUQa6KnwZ8OdeVC
YkIiTM1VaINHhb+F4N8RnlGV57gPwAfq1niCmQNkQ1RQiudIHMy4F5Uo0GHXLkEp
TkLbx8tWLg4GnqNJl4gUgEyac+a9nEmFtxdbFqL1Mc8qE4bR0Ti8jSq445PWib3r
SnZ0ad1UAsnb6c0q1mOT88V/DLNGgbdIOu7yvDYmqo/x34THQxfErbdeCeFRxy1Y
dgOhamF98HS9Mh5/dgiO5kadvmOzhgKUsDOOSkMlVIRw9JfXTF7qbjNaMH1sVpSM
/te4oXNvD2IWKg1CmvmbJK5gm3eGsH3mbMR3ExZdjOpLcafUEhb/DUcZ7+sJeGHV
RQxz53A/aTrQmtu8DDLa2tG9aVUk+t/hNx5qK5WRlT9qfA/3vsNbbLaO33yGlxls
JQCIqKT3OFaEG5K+9jn3Yn26JA5p6PwoWEkz0C+vwv6L07EXnMt6ipPL5mGaU5Sg
TvQr5BH1ND4/OzJRY+ud9q90rwY5r+DfPIiI85VRzLvEEzc834PbQYtKaRThTcQc
/k2hnN/5VLHKY9XjOKhh2S1uLYjbr4/WD6KPUSHl0nLuVKdrrZRIVxUfZ7dYU8Ur
hp983BJ/dpJKKncITWyrkr/4KY2LBEk47oRKBD2NA/IpWCnnb/vbuAhLLbdhmpaj
sfSuuy0M6imRYVnnu2aubbR0fy3UgMrtamasHKvuHoJAQz8A2cBWSOrtuWEseNw3
gd0WEkuPY6Rd35UxTJBClmEoyrZPdsCBNusbqNoY10eNcLA5+ND1pEIYUXPkG+AZ
P3h8UQOwtT0GfUUielQ5re89vgXbaG5M3SUl2q+0OETr93piYn6G39Txdt43c4U+
aQ4bi8GkJTI7HoXX5lsClFn23RA8JbPkoH+9/E6FE5Z5gbfRxK+Ku2Q8y38lp2B0
LiRskhmQUNM87NMtUkoF73Jf+oi2LFrdu18/SQhOmYXjm9dAb6pv9N3OWZ8U1/8N
+PGNuf05hgwmQq8+Ea3BDOompfLbBS7MQ1INeoGKx5u6XHBZgoRdEVcy4HHnXZdk
vlYmolvUyJbXAqdHNHDZG0b9YZzEOvyNUg/dzeZ96WCWYM4rW1xkLPfKI5CNmIZV
BtKltFUDMZ5dvQoihL0O4CPdcmfIFhPgoqviRSLJ8FRVCjBreCbiDuclCO0+tm26
iqnK2kXyDEuY/uLUWCqSkiuJY6ldgiTLmSx0Hn64LLdR0xi0d3hSKEsOZGxT5koj
nTfMQ0nwfqc+x4+vEIe18XGjLyW/ypqyqS93mnoWeOExbOxQuyvbqQA+Nqk1hsGw
hASyeF/oS7SbhCndKfLxshGldgHItILkaqSn3MBtPdUpWuQR54po53npXc/SFNaW
Dxr8fQ4b6jywAJJcE70O3MdYOJR4em4hAtR/7yeSDIX5A+IIBGTtmTUO9LI1YEeQ
vpB3VvkQxlDVh06vYFjQme4fNlwzC+ZD7+qxuKvMNDBFsMR7svTTSKBLLs1ZR35Q
86M4o+GZQbkdPoTaon8YTcxndWf2eLPe10iqjMkV+WTiO1gk0jTRytWCmnJD+laI
Rt51GSyRlt4ibB40bXMSDOx/PmUS2aqWnHGwAbTaAWiAChdvKkc8rGuc2pBO3roU
+hUjGJ8kIDIoKRL2rkDXB9Mz88EMNH/yvJBmBF/lD2rL7qhTEv+4/G20P1pGBfCo
XWS6uSfm5J/NWSmZZzCw6IEx8Hqu0J8LH0KQdpefNc9HMig4sS8IlAwL2WsCS5TL
jRv8Oo39Z4PIzRZYaclTdYbFkMW4tF3/JaQlvpyTIuvjTGcR/58Fhvoed5+s9q6T
0GcqJ7bCPns3jDrA8rNSjAZ9k5oti/pwlGORLtNxwttXnu/N/TxGcNio9YSJwT3R
RfetJXkWj42xpZxAsWqj9fsbSJxfKqKYQKxoKedQpU82XeXB/691adStlty+hU0V
O1eshEfsC6xhbd8WP3uWkZYkWmv0utO3u9NiRMhsAoCgQmkjWrRCVb68fMg1wX/8
cfDbjRSGZZqhl6Hg36m63Sa+3dPNfUL/VAaoAkIsaUiRWUlv5Ih1TogwNHD63QgZ
8nYyifue1pyIsFjgVO8bnCu3G2zpyXjJXInPLcVVkOH9LINMhoxnhQELUXgUA1+X
bwdN53seREJWDpmd9QwC/wQdDVFxFf0F4GTPhks3MBNpP9+Co7qwcYs1tg4spQ+t
r5VCxZrdoM0BWghbL1TAIM0gqRDH1mfAXHru6NMq6/VcZEQprL2FhiS15wFsVcqc
Wu5YqU+Fbw/0vjlfkBF9/HKzCWodbU3OmCpIZMedJGACO6MyYoHmkE8v/C2LnL2v
ZyLpFjBy6+jxjgJdhDm0N7Scou0fuXOjVl68B7HURgLIg5hPOXMBCndxqBolUD59
8bNh6vTeEc/PpZq8zM36ngFbP1Si1rNAmS1TpMihdZh1NF9b3RAnkIIqsUBhdtAJ
uYrVYJp/VabvDFKMStxLJMwapMXKwGLEVDFXWosLj7qhqrsobEilM2D9D5En2B/J
lymIcX7WcZwUiD9LpJ7DWvZF4bg+vdtkhomlAgaM1v6s5V5ccELkUFdogkn/h9Ye
gSF3GLh1eC7GP1TFa9yZz3i5q8ZyJPUFoxFgHCGN+2a3v9hyAEQBue06ddevFbiS
pE+k3eSZCCI7i3MWGiFZuA4+gRwFpSGshiKP8EV3tKRQDrp+YVYkqT4uXXY+GF9G
Qb5gEJALwFLgUz78i6AUUoowKqadEnz9lfVrCrtz8FzQqIXRXImYBsfrstTpAl0m
Hgx4+I3dbKL1Ayr/tFbXODIzZ3pQieuUIOwTJEfhj5YNkFgaVgAPD3C6mW+uicuz
nZCYoF/OTTJE456N7rwUX0Z8Zu8fjDS7oVRGVzDfuL7SCLomBTo9CVFlHIIvD6tN
nD68N+Vk3imSHJDnKJN55QUvZcn7G2vEY1P6phcbuJvFqrORIb5BTamrmTu4fFwB
dBdHHC6PXv8t9U2Erz7oIkk/gEPySf3qWynVjk4giowL6u7lx0kjEDwJrXw3aZOH
DMjY2x0/fXEEOyCfkXSAwbZcy7sCfrLSF1iW7sNLbgRtpYcLgBNRzJ13a5bFLk7O
DzPP2wGjp2uybgQco0NEu98VfHZOr7Hc/KGyYhHIjLSGY6elDTA08MpMBbutEigd
mZ0qgCIvFVZtV4tDis8sTg0um85yqdjHxgfXsEDID9LwmJBwCOam4LBymMVQX/eC
SzM2+Wo89kW0dAivVtx/ZWvfGVGI2BqvS9UE/ncvU88YoGQZ9DSLhmHFb59QnTUw
s2MmoFcHN8yfmPRtxTbZT0bnJ4njj8iFQE74n69Jy11c2Wt6piSyno5OR7j8QcJt
vEPdQUBzLF9hG0WwvUuoVdrsirfhcKO00Ts0Yc47REFWGas+TNxHq3iGTDsA/MkC
7zStd4B79EGt7n4m4CUBTT5TWsCiVIT94PElQmNPnEAuopB0q8gR6jfEfzB2ceOq
PP6eqR+sMj9RR4HReDjSV2EEdyJTg9GGSX0eUR+ujrRow5UIBmYAeC7DXs8wMR+Q
fUUixeGVHTSEKLm8cViAQ8u7vhRqY0mjuBa3ArHWcVhdNHIntJATgTwb5ypUjnsR
hh2X+Y7RKwfcSXV1q2IBuWDfHhV6fVS4Y0GeSo2iHTFqdVUnjMPQWvKfIYWquN/R
UvZSx2pPWvjszHZ8rJuzj5TflcCH26xxZkA0r93IX5gFQFVvXgmpZ7PltoYH4Ios
V0EkIDkAqVSjisaI01xM3l2Kll0izRKdCoLsrmkJ0c0s9zezz88wmbQPsWE+kUw/
VOLl/lKXnW4K/5hUJddXTUuEDGLRIrp5itCDsk0QmZSDsCD/KgyVlWIO9w70LLUQ
gKSWR2P39gyxGJg5QjQZuY4+ZnfImnVqU5u1ZDtCdMjdEWJlJc5QeK4wS9oXb+vU
jqwcDAj9YV+qmViM+MZ71ZwjSVFYvWLKfTwrPvujBpgyvBXKHuoqNjs9nkjA0k8a
/UaEewJc38aS11jD2mmhy3aNmSKIKG91WZUIgEAFJTuIlH+hO2ERXT6My/aAomNC
0q4PkRPjrXTIHaBBs3VxG92jGBFHdfueyosOl2t3g2LMRsbAX2Ai9pt8L/r5zo2h
a46Jhvh9IqEPIUOwUQC+eJbaApCsJUcNWi6nzW/OvoVHdktjp0X6IjyiDWGz5clY
+iahYL7F1QhrwngjaLO7VXKr5DL0E0CsqriyEE+rJJgS1nmCZYu5g+LuZAzQKk0f
zSihRR8dw8SSuiYC/nQOtgr5JJvrz/NzS2oAaVA4/00whDynuKeXTVJfiXxT1MTe
sGblyfZMWBrwAiaYh+olMKaBBiEXFNChJMIZyqBjKaQSyvm1bNAvrO5zuJDqkbI4
ILyU2aREAyOm60EQUVUP2M3Bscw6obp5uxyn9xDufczVwb8Zn3AHOtGGM1k1dIcH
Brs4OjNfkHsez74vBqrkHVaPZE6ORVaYPXCUyj1Ee4x/M1/iNOz03erbCTZCVPvZ
x3nAjGiXe/dFrfCIqzxGufVLZxxMZ8EfFcXRQacnYB3enlcrfURYooN8JK0iQFLA
ApWynFEHwEOzd5WrmX4twHDg+cjBHwGXw1FwTb1GfGZUCTMmTok6XkHhTIy20LBD
DlPXnYWG1X+VVRpk2woIXLxmKs0aGXAowjAk4bwm4tziMjz0hEXjQlTmb3XjTbEl
LRybQFyMQRSLeVE+W57PiJKbjz2oUKGUg3D0zkUemoheG7XNZtd6Zx06ESNR/IdW
MLg9HD9GN9tPLT2HeOxUMOgbRJjFoTNgai/Fnc0otaIeHAaWM8KoAJqY1oAupBUZ
UxxWzYK2OdkVt8fEFrcDp/F/Mi3bd0XYAHc38THhcPpfyIyD+Vpj9FSmnwsBMkzn
0T7jTJegoau9sONVFiyx04jyJJVOGflqsF3udgi/xInwny8mhEPqDFWfim67y0A/
BHDivKn2a3p/kfx8I5SIVhmMstx7L/5aE+SPsGBMAFY8fel6Vma9rLY1Tc7PZwpe
vg2XHAAaumE3AucvA2EbKjnRukXBqK57qP2WJvJLI4RqjtFnzt4k+SGoXxGjkOJG
5b1hi56azz4LZPZEWkrij09tSI/kSG65A+Wec5d1YNJwc0R1QK2LzrqtXRISF9DH
Mwa94d1pnQeGPA7x6urqOD2NbseA9hZ+4DwhzEc2Y3fAtbFv59rMqwtxg25k72Iq
sD/PnukIicO8VNFgZG0e6+jExXO61UYeMfSZ1e0LZqFLuAkc8qDJ/sQrhFBumiRf
0BKPS1pAIyrKrtGesfBBPuutWyGwU/FBROnklii3KFI2c8NZce4w9LTeVpdPLWKa
A5Qn+igFIXwDdbxBJ8WPp27chhZRgcynQfDUPiwl9j4kFMg/aUPN1vu9CrrRL1ks
ichyQuwSSXzwC1P1Rw6yTmWXZXm127Fyt432bDLsyPKvqU6SxEmoGvUx1i+ZqM6B
ShrzHEU4RXD8NC6OUUg1W3Tr9yPE69A5LZuWc3H4ZpnRepvsyxhrr2+At5qqHjAF
pzBKlieoHGaCSZg6wZpLAgLDn6vY5ilLg3xBOt+bcEVcjW9GAxOTD1tCmimkJ63N
QIKDCSqhvJItq2y3KN9D49WxU1sWOztOZQW1UQaaV6OSyXUQuGE23S+GwW0mMJmF
YM/naKb6UPBhZLhuMnFm6si77Q4BpuzxThfoO+0oYfDlL+PGkLyvWYFI0XkV6eWv
80JgtOWCDt9Y3iNy6/nQ9S/1QpzqDVwvvGQTJqtadOBP8OT4C2VRDdcO2Xrf9/3i
GaECXSxu+lJAMuzRztdbMJxKNfYusAETX5ye6ENYdBgzeZBgjAxk5EhhGqazFCDZ
zI5evX9W4lYRNXoKQOkwPuOOdREah+fgKX88E5iYUxoTu15hVWrDpg/df5OKT56r
gZ2VGYYr22DSR+olbGg4HQhhxzDMknGboMu53szw3ZoITRxs859fuFfRX7zwo9By
jnUanG3rOLIW4A/gTsaz4vZdWCKNlfxDkfA5Gq1mxGT8Xsxhn28TFt1IMNLcjWIA
WWGuKad5p0IyHdZgRjvRrPm8avFxjQqYYbfiqkNnvIm82NLvq3xW4swW9ex5YE/8
oOhA9xybBB9HzWp5sqnK9QVOJmZOUu2aYeAvxtBaUqqrgJPSnA8j9hC0eN2FoemY
F+iia46s0Dyo9iJBCobDhBfKikw+qpCMn1Mklxsr79h35+Zr6doxMkEYph64Znz2
vdb1bUVkMcrIk98oJuUfMhI8WX0cxh4FCWXp8XUa18l9kJeBqGN5MAac3npVcJq7
ABye5128jxKlstA4rqeWtE9DLCMZssrQhAxTzf8VUBsSu2oCtdIp4pTyBWU6eEJX
yWaQlXQGe/AAfUOQYHCdJHcA3+Djb1VSK5D/Ct1/IHBL6s/HuvIWnKsy0WcoRDF9
ibO5ZasWssid1GG/cr0Ba96/rcLOqwgMJ8LxfQ30w2svMe8BGdfme2edPYxoZgYx
JYEg9r/Cy8uQ+ZLCbJzcgrJoDpz8C53y0+j+jRo+Rh/Ud2NNgoHnXkv7NcvFEDrc
n/BFSatUo6du+lMHKuRpt9rqh8pP6yXv3gXG46sG6KGhqeRSehT5A/cQ+IhuNjDN
6TVNzePzbaLW+9LAjwEezLWUHIdY/3jfhvYxscoDiIceiLh9bu2AuW+aWYpwxpc1
Ce0T5hPLz1trOS4ZrUmbCQV7oLnFIFx7bOflV9vyUIxOyRqpS4n3nqRhcJJ8Vf8j
6eKGkVOWZRFRhzyiqliRbg1sNsvkdqgcTiSrsSLeG7cn58q5myNRF1UIBTBQubi7
S3q/Xp1LGVY2cIH8lljrT2Iq0XUvZER72C5oZAjLpCOYt2t1OiWtXJTLcJk9PhbU
vzl/SAo0XFPs4vjnudPh+88QQ+6AtsabdgFnIhAlzZAnyP3MIL6pNblby6aV/ygm
bgsmKdYMbUgPHrQM0Wqv9rkHUJ0RBFFrHeo298xMdZ7mLzNVpcKyq5hDKGS9W2eh
88nvZl/0DTZIk+Eg4TXiT7mbYfN7TWbE6rFz8xQLhvr3+mUutymXn8S7DyLH18Ev
JRxcQM5GxX7C00oddKTnkq7daMNIq4jhtgBK5XPmoAI+iHK8enAyIyTPaOEQGQw5
mLarmsRO1NX8JcmzHyzaBSSHEl+pZQvFum/oqE3jKpu7KjfuYffid0QHx2bCNNDZ
5eHZxy6uB/Pi7pTGp9SWPSwtfi6cKCUOKpsMHRc63qtpinHynDQGJiHYLkEnMftB
tRmelcXVOCX2O/khUR9E5pNr7K9PVhzMDg8o81Xgbf4Ds8TVYCfUI3i1jKp5L+XL
JUKDMGwjhHpaFopmDfTrl2xemmQ4IWAQHpHgBZPFh8tToOXOv+3VYXG8EyGIZThL
9SDvP0oZJyU/qKN4NpSpfOCKCC576VhHZBYMOkp7urSB63zZfQNLTmuaDN0jEPAX
7KC2SOcpNixxWVvcGJIqaY5/npBzKypJmRumu0ok3bUeh8bwQEZ+UAVkbX0zZrKo
fWh7sM3hTUv//F3gXfOvHxtWIWsqU9ccWDp3x5p0iD28WGKYuGUWIZeUDjQcSUP1
EJ8B7uelWgt35iTBFcgNNLQF7oeq1xrVxquaxIR06knmY/dS5oQyOt8PDrC2vhmo
oQ5O0pVAFGcFKep0qTtm4YRPJH2SvHnd7dvpyK5niPAKJuNntrpc+8+GUnHP79P9
4hVsy199qudSTcNnA5Kp+s1ojEm4kaae0Iatr7JnMGzlnTaiQjTc/JkyJI+oVjW2
RPHFa73M+lq12AUjFsKlWxBO+iTo048YEbxj1fhHvqhdK4rQgzydBoXFRqQlMPQA
bo6fnXJl6NSsQBMHf3AvYLQDdIWtVuiquyaob4EY8hQLUVQbZSSXD/URTUuvPCyz
dNP1b0JYVWnPZ4ZOtSvagDBXAfzLM4H0wUiDUoJVosBnCBipgloK7qde2zmGaRRw
vDQ5mOo+XOcbua8YXYRM7JdeoPpSur56jezVcqBm10/vPc9coJASgHfMrd9XVeRC
U525bdBJtGyDcrKzLjxPmYFeJDD6crMxsDJ2QmGSxkLA3+/xr1M1wmVJ804U/ye4
MG61hGqLLlzVQaiUT5OnEeXFGWrf3uk0diGQJPSeFKo7A9F8Yb7UtnqZco+LWEba
ULJzO9IXrh15g8BEIA8s2LN6ghXEmrncLUJkg5utHnyFRBicweFawhHjBxmcevq8
E4IOTf6ACLZ3WMFeVOT79xeXMUJfZDoQ5ONB7hwUNMx2sG54epY7DjpAblVKG+CY
Ze2z1YUjGGsmTldOaKU3fY3tspip+x5+zMMEH8Q21QPUIhpCQU/6nk1wKegJ45RZ
YSPmLdT6wvZzt2K7bUFy81KpFHiywiYK0Ion0kSMT7yihadSicd39MIgw0NcKvJj
xh9spC7gRGA3Bglv9T7ABh6u5rX2JsFLboa+Q4+Qnfzg0tKLph28PWq/pO8CUVTi
GvsOAyo+a0u4gGWdIpA61dFV6jZIaFiwD+8F2QfRGWWHKquxcDNX49m4YQ/Yoqlp
J7PHsDj5lk7uDF5Fy6YQ/rUtC4UYCLmRQI3CrdvWzBokCNNg/aLu8g0ytdYDFRMZ
OSOwvFAn/1+K0YSZdTVIBih/tpRtgTH+u9vTLrhlNJgD1j2l7dwAeGBSYdqA8nWZ
uJ9Pv2ZEA2nJJt4YZC5ozBmzuvpkaShUZHSmrM9p7ENFRKJagUu8TyR4aVpf5oTB
wgU4c0rNkrSkMBShRqGtgNBDjwXwKb/pr20o/MBIND6qnOWyVR0uQAOJmGrdXfW8
8/NPWJ8WPJR6mrdlUtCZZaFqW3mjHzYAxuho1PQB5MlcjhRPw3ZZBDx2dlqGSAPo
78D7FmwKPE2DZneZwGEt1q0QMD31FyQasbNOE7KValgB4ClMTLjofJvrQR2VxegU
nAr/YQV/6fggrvwVrfOcnxkAkdVfufDDiepXIv45qaM1g0eHKouG0Bf0BvmO8MyU
KJTJmfaVWg+grQDC9plw6lTwMz7cviS0ndW7+9X5K/rgHCpeCdPibYwb3bdRNwm6
sbHDBvumvq2Md7SL6Lgwt3SXkQHH88dFB134VJ0wWD+A+hI5AT2UOTey5MN25gdQ
G3E15HQlCvN3QjZ8XgKhT0JpfuviyZ3ePNlQvp5LlnU6TO6zvL7W31Ibrgbx1USE
lvlpHukrnI8V8TTa3hstAOig7GlEuqyHyRYY126Ia3xDjMkWzSUhESjjnB8U0uVU
PJQQ+xjj5BarUk9sUAE2NLSJF9KA0pCxpGqUH/ZNHAwml89XEfxi86LdTkEFqxve
oXxdZZ7ElTF7u04xRCsAQ19oWwFRDnLkjcyTm+APOwENuuxaD5PzqEv4kJeGmHES
dbQnvfz7XA6IlAEyq6EfsXSSi/gb4I4oaFLOLmqVtwiIMAJ2dqAJe/JOANBmXdS7
YOsS8Xo2WkQX9UzV2ngc+koWPatJAJ2BKQLrS8/dAOIdjsgvhBCA7YQeDE0lmetL
eL/vdLdUrBX6SrobLH1zXAKTDL0dCBfcJfTwtq8s53fntc/tGX1qt4v3Rk9ooIkn
w3Df2hy1knx7n7myeHuKqF1BR8ul68ZHzoKiyR7qgrIRHyDqU8Atcucs32kgylM6
+OFwGLF/G6Yv6jYn9JEl6PztWsurWHQrXV4RI+fLGlFpQ2qgtreeWSjk7OyEILdY
jicRY1jWGWTJ8tW3sRkM6aGixJ7U4X/uGaT4IwNuB7pFrT3WyUihnHz5Ycw8QY0X
sQ5kLmzkwIoXkAuCbbJieOqrWIFuDLUi8V9BgRnnkRUzDiMBZUgXiEkBm6GP1XrR
AxzW2SRxEnm64Njgrix+9gncYWlb09k66rvJzO6ya4b5H2+35jmrJYNI7oirokx6
oh3Em4kSCYqu+m53iF+uTbQeCR1OFT+fGZCvOthw0YezlnWsvgN5yXiUxjeA1clW
eGin1RkRhTvMWceAVxazsty2GEn1gyLanCyhxhQxdsvxjRNskTH3fLY1b4LMWb63
bQTO7q0XD8qhTvAGNkjDGy0eqct8CCFt2ZUcLg3GF4t9gFBBESMgTVIjg3ukBOX3
hSAtpkpqL4MpzqF88RIaxDIsyIYxr/UYhxmk6d8gmEOycoJr24lA5es3BtlhYZU0
qsunxOpt9l7VSZ1l/gKj1gfCyk3gye6N7x+vPXXOGkjqCCZzO9QIZTDd2K7WPBU3
DMgBMoj8V/mFrmRe+0guGWru8LMybnZPS4x2TY344VB70ccJoELl0Nv+k6Ymm1TU
yh0R7ye2JEbMKPklv5nurMRunFBtIdExfDY/1ZN67R+f4xem3fgJ+86kdPcwLZFj
XYCRSt+Gt7PJQ1sWMBAfBIFJ9SihDd2Th7yyHmXevfNgFzEW8wsUwWYnWDqf4FWA
tzChi89HjnnTMS0qwx75FAmAF8NDARmpBPh0XSkNZsW1hMYir6PdrmUDgEcQnvRm
r7HuRUE4nbNk1L5Weo2A3YQtdO8kEOrQEMCry02cZjR/7Cqd+fmxymBIGoMHXs6F
8Zg+2lqTlYVu+IzSwGOMWLdo/UIvahkUKUPi1Cbe2PVhIYf+gGBTTe108e5M+Pyc
pFIDgDF7OdAyZyu+SFW8TmDlkF+rh80HwyIQmkO2GPXWcRPbCk9EDHZXaOUqFg7f
KlrvGLJu/ZA4ut2S23/0zTXl7ej53mq2rwtRfpPZsaQ6kr1vzg+h0xNJnEwDws9G
wWCOImeb1YCI8yCA5DJL/3kHaj1z7YoV4xkIKbWO9/YfIeO+JG4+9y61p9fxVfK8
o5vMJhdRzGgh5xHOSy8cmwPhFN4uLlBRM6ENA93W9k4kfLU0nwP3q1/M2K3sfQw5
SRxTL6d9yD4MCL+LrVPvPhchSk0Qm+yfl2jlD4bhH67Et2374AN9+NunfrfenIMT
0gDSNw8p9w9iGVllymvrzs8uB62HHf1WMf0nbvwj5D703NGB1bJuSXER9Segj+M7
vhyHKCeOZNwX5Fihi5iRfaUZE8+iAyPWqOJzZ6Tf/VA0zLsH94counkUnmdp5ua1
5nvQyPijVE3zLGmv6b8oGnMNmVjs2U7LhFIWBFXSPCFwz/5j83s2E7fcOrEBdwCJ
DkGZcY6NR+D2h2kRUvbl7yGSuhRS9wlVEuhkIYez8jwOIXhTGG0U9MKU+cnI1tcH
qxzdKtodIUsWBTs9kxIMOBk55JC4cQD0Aly45XxxFMl3MOguW4fd1Imjm7Ng9HKw
yDQak+Tx5FkOT6xyd7i3+3xTLr5pMeAjcpJbFswWQ7r+5w2vxvc1HMRtNWEE7ONo
AtjtdB1Zw52EECvwhp+LLbDUsA7woQ8+HRRlzS5mxwm9q2+McVcQWz6xNACiBySI
14Qp6GPNMF+58NCaTZaC+DnbtZ/p1J4ATO7AMYkfzqfN/Y/EFkkRxS7F8DKFzISx
2l0yuuscdtKJlCM5gBesrZEdvhWZnS5VmVmkF6pWyO/MpB8uCQYyTAT1N7D3q2nM
kFxJKDsxXTKxY8BTslL/9pASIEKmcQpeLJ8pYIck7MLvJaiQS/blRa9C6Ag1Cg5M
/RWt+PV3aJAo2lnK3XwrJUa6DMWWYl0FrZnGVqrYkKv2pDEWbJOc3LFbJt5BQT1s
M+zvYY8E4ohsh/dS6gu5h3w0wQKw3lz0HZX9IT6EGMpQoPDI0w5Ywx7SqRQckiDE
Xclj2pR+azpAPmp5oxHSom7HcPlz6FeL4fk2ddHAqoe6X4GgsKte84SqK5BtP7n4
cR2UMrSAqg1719X3TSQpXeR9IbNlC2BOLi3LHk67Bb9S5tf5uovfX5LNgXAsTnYm
/78CL/MRJlBfZSZvynT+yXt60DOZsaXadjuv3kCxSc85634cHpWWXq6WloMNxIu5
2wQI1V7InSDKm3tAo1VgEMEzON2+SXTihzZeXeQKXslCTsbLVeKblzjtvhKPAIkj
P0gP2+OMI9/mybXYTKRWSiMl0H2Gv5aWxuYUKqIOkbqLXItsriUgUYFYjwMe5acU
aRwP9Y36VcxNCKVHw4GhjV4yOxYHbDelfI4zavzj9o0NgeoVtIRo+QEhdw9Ga3dW
DqsMPSua8NWz7QEt6pEnxNKVmAlDAruqcaLLHrLRjM+6aKEiYprez7KoT/Jdtgb+
iWp47nRrQcUPEcrfKcE1MFoV9/7PH5i/6j4rde37plAGirPcaXKTKqlyjhgF6s/p
qxndu12bfeI+mH1Id9uyrV46zqNNkf9ELNlmPq2pmpO8WJ81OngOHIpkRmJTWyw+
PYjKcdJQI6gn0gcXsDzV/34VcdqdHG7hsrprgyEm0TWKgs2nV0aUzL0PZjMWqvub
5KQ4hWcxQmahVGflaBIMOAYfPe+LCqBNgkaARyQtQp3v7NmkzgKcvl4vjJjaWi0/
Pn+gzaw6r9Q6yFkzOijsEChkRopNXL0GSPMhsWfZ25SAcbrLdWhuVA8Umu+mFPPt
UNC91RRBFrZ3O2k9W5DMYa2ZARmFpNgJv53oI0IP3XSulvfoEAI+Km6qgWkVjldc
OduXtC1j5I/rXZIFQMxwU3ndr29Sl7X1bcqCg8C/g8fFmJf0pjR8zrKJ+Jix8t2Y
EDzTBeCRRa8ltjV37V0M2prr0ULbnHy6zGYu8KCxmVXUjjdknIUV3gvZKJ1ixN/l
2K6aXPjH5mCYJJ80pDiiwdXzKtx2pJ6i2YoaYxQwxFXQkH1ZFDI65KlZBSMQBkQz
xgvDo5y9BvsG8ebhS+YmWzFjWbm6sYgSX0slbg+A443JLdr7iKuw3pymuEAONSgJ
5oMg77o4AskqjO8r4ooDZQv/ibKJmJDcv67k4txWzH+Ely/DZ/lthfJa1SvBjsXu
hgb9vW3PlBksJs5LzwB9yp0evlCFJKs1Mr4Bh0ht0ido6fFL2ZJYnsjz1GVV62Ry
lXdtVN05gMGHry86n7o42RhKtZOgULAvd4G+D+RCDIhc+f+zMn2ja36NgLd8umDt
tGKHsslrq87bc0QIRgvYSYQAAUrYMkIsSVei3CROs5ViGhJLPuGiXTSyD6Gd1192
t7tWDNZJWZ6KsmLd5WjevWYHrhhNQkc91pH4sPDP0Z0UeKMjerwoBKOmaHO+6Q2H
pvZgU2cS8V0dqv8KmfP8+p/Nn9NX8fqRJ9lP5+tWEtG980z9ASrAYFBUl7hcRomB
OqY5MKE+x6SjLUDKa0/g1hpjDgpEMVzl69JDvX9gPF8QipSuIdfoBekoy4+e0kgS
M/PuDKeWfIx8ajDi8tqmO2Axl3PSPRFEseEmLCYSPa1p2nVud7iXeOTSMovzrPgj
cLw/YvHXhu5SHY8iYXgOIIxN6LZ1CnGHnTpgIKXT6DWBHYl/1PtFgroTA/kngJk9
XLispn9Q2ikLiTAOCDU/DE/p1ECwuPFFrHgiJDP0sGNORzvvHp29bKbIJmmLUfus
NhCiGcwD2tbasKLFrSILph5MN4PCvjQNrmUKsR3FurIFccWSG5bGzTZ3DfVcwdLI
iDBsLdP2qZOh6GfAd74YkEC+TFHziJ9QK2WdLKcjso7AOZFAH28/FEqRx8iYvJag
mbu+fEfcuUdPaQ/4G/Ws5i5qwQATc0OK5+ciTBUrKHtyWa4WSA8mEkio9JXBi8bB
6TPoqMB3S8RZddDB/ja1FeUPjx5I/QfP2CoyalgfuMQyGCUNg7f3F8l4/VryUE6P
4xvNt/fLbjm9cPxlvdGkm70DLkZPSEsNn7X/f2KW4i3wThdIyhYyvah02/P3TXEe
MgwN/CW4kGTrLnQrRVdxJsIUZdb+UVxqJyIaXOJ3Gp+XryzCgIr86UFMX2ntnF5w
fp4+gTXrpL+3ltyL5KWqf554Hl9cguUh4li56LHFtOsC5laLR86c1F++Zb+PCRDk
VPaDLCNgxlSxyq6zjcgmqXUsCO0lEkcpkxxtYuRa5XB7NwOHMNSSxs0DRC5tsswf
Mh1pn/fi4n3XcPHqahTBGrch7EY+F2cydCLl2DvvwwUkUnhdNp6AdwMmDUGLkNu4
LITS3nyHqiO6jsW+JDJ1VMz1Mu04DQSWHC+zTfdEmTehyInrgs9zB8pI7Eo0RJAD
u6guZDjLq0qx1CSz2M7g5WWuvjBikxjuRikzx+NBXgVHjo0rVgfjiyyic9p5A/Eo
5jhpBrOBP450NVdthLSz9MkM7AiC7nFUJDNjXagFaxpPmHFLKjFbHWNDDiHWZx0b
tynRSRDwKngDOFeWdLrrXIyfreT00J4cRf7iEwyiGKTHIarrwsyXXpFwnQo4xLz8
KRgMAtSimxF400NrE/9y2AWJRIxQAMWNthRiuIT0mvFhoO3D+jJLD+si1lQsP8O7
no16hJxyyD7UJ+okT8MdsgICBFG0Lhgodotwnvb75DlyLQztgFHB+wWEC3jK2Xrj
p5FZn9dkV/ybM0GdalrHNM7EnXiQu/YfQ1px5HiRlRRAoVRtmMJW95zYl1LKCP0K
McTIOP8E14+vHTQDvxuUMQOQoal5tp0+jCUIEOs9mclM71kWpiijB0YRpxXIvMSH
KEtThZwkAqCwayrbeUeOFvmvUA5uBoAdp3CZfLjKFQ/YoPkjiTpTHjEwbB2Vf+AC
zMYX95A8bnMnbPaSlEYPQTVT3A9SxPxClHVNyYv2UgjbknSAU31EuMA71FLPscs3
QT9kBCEWzLPQDDbmZ9VgbaFdy/3S8M85sWQiquLD5oZH3suowcns4Ot+ul30Npuk
Ez/uv28AWYr4zENvbkwAZb7eYpEFApAOX5JUsqBWSBzZi7tECwWlnYugL0+IY3Tx
FacsRyJKcCFEfV/eZKDcwfU0EzjG/VRYYSb/ZPREEVu+0Ph8A3OTGPjbqMmVC/Wb
FsFFfGwyz46wuY78HiZBq3ojq6htKoI50fgX12sepnwNkMl1L54wUS3/DX2k72C8
opoV13BPYpf91EHt9FAWy2JlPhGvdVGaMkcrubi5BcjeRRRNr1wNbXUk6RqbRh1n
bbVjuNtAvHm+tadfa/n0qBamB0o3b/NhGLYPQbk6JOZ3VydAHyW6H44bUyCzQFVL
Mkg93kBUfPGmhmVBqC8SxrkJrkLwzGMJy/FlAApbAgdOeKs9cEayWhitLHtqvvSP
A0VcbVvTXkNFQ6aOaUo9rZ1CVAes1L7Jx5w/V5xwQWdkDivLr/YYgr+ARNs2VQdg
2ecgulbqQ3qLypJnhxV6KShviO4KuZ75qcUYtKAvsARj+XP9rPGtg9VbYsfyPrGD
R2msinT7pfkzZMUkplSuugXu0B6vS3i68RtKykd0M6DQexlgAhA2S+MCEcu7hIHz
AWQRNWygLqhYJ8qkVeXr81kl69iDyGh/+AAsXCpn5aHNigdQTTAVdlh96/YUK1FB
7jD1WgdOiklDbXbX+ymTyAkIzZ5Ca5b/Mbrl6OmxUwH8qVaTCbWGvpv3n/LkQAWS
lez/IOg70gYzFrMaZy3fcMKi07uiFpyEZb8SH/nx0CkifBalsUZyio+NvFk4KH/1
3M/PfjE6ODG2U8MvWIwBojQCRNkAVa6x3cg/U4Ah+9KdwLsTKNDcoGtbrdK5kQnO
pkaITyJwL/gjVy6rcHyVEeBpJmbw65pEOraSqJ8H6lPnltS4SyLR/yhTD+WhS7Em
RL/UK9F+1Ebc9KgPCcwM3EO7r2ndpHgJ6SjUmUSJEvuDCmBeA27Y1y9g+nyajg99
ht/H/negwrRkfVvsihG5hmOVlu5a9fBSc3Qfi6HxDq85+khTMnDerxrh/tGl/CGc
MvlEymt29yuhLtUOEMR4R0OoI05X/N1lB8UPE4AAJDScLJK45P9jDkyUmbYaDtWM
fPx4czSagsW79z1lvFl30sIJrNLQbH1mHSORq9LNLUBnvcAUbWkNHHehQMOHO+bf
zsNDZ//dabABv5O4MxJyoN/1diC9+I0869uXgvvlyBk9D6dkIW1YgB14azySq8+8
6e7KBG3mRZElg3bNexJLW9xCyJm9cqJA+KgozzQE5sd42IMs/T9d74s9p1ImVSpU
ePwF0urY+CKsxy/V2ILBn8ovc90vj7jKmP0AMQT6hFRODWMh724HbhdZSiQRpmIo
8z6+CJ2GrnYL3RuGAlyZU1Eh3awXzFdsJHLxRJmxkveyjGKqPrKadSbcH0kvoZa+
XQcBLStmfpT/NwKbYb3hx4U9oulFISkLo8f3zfeKW++MP2GLNpQM4ptmlcqtbxVa
w2xXhJLBeweaJbgUXtsCw5A1tlNzgwOVM3FG2h9+OmuSEsdBBBZp8klJ+QlikL8W
7PJe+cEev1d5ce2238nYgzDkpL4MXgMKqVDt5vncJ7i8wK22VzIPavVQCL4Uv0aB
BIBSSJZkh0TGv67HUmpjRfSeJrYq7N8Z2GjJIaljIH5oA0dYt0TIFi8fBjF3sSIm
g0bIWwkk1W/nPKfrV1r7ydP+mFaIX9K9d5mjQaV6Wu/33MG79Nbrzk235qzsHK06
n0xyE8/44A8wuGwqZQkHp1ui1U0Ik6mJWoX6LAOxCUo0wmWBU7hUaKmqORmlkhvs
0OjlvKidfTl87YctRhs2luuV4NHlomFx8hkWuOofpeIgawRswUFUBFJveRw6DWcr
LwYqQaxLGDl4U4rZuRzDwUyJIFK9RCjXEp6SyfAVDKehV+bowos9jZSIEiWV+GQx
KZGbze5cMjHCZ0S6bVfEftBLAGHFS3ioj2R0FU9JUyBlaGSgorlfb4XIafYdOaD6
8GzYiZ3szDm+GdEUGQ9fNfqnUBCa0x2mMcpuiT1P7lo2xA7L1TPwl7xFqVeL+828
ybcSK2IbfuYCAVzGFIedFxIMmLMUdFtRXqQ7PeLYYysZqdSzsNZsUDHEgAcensie
R4EZpiiOedCmla+x4uCLMOwMcTF6R4zcW4wNWX1sh4kiWLjXEBky+KAPBg6RLbSq
n3HDt9/Iuqufl6Qlg3X0oGvRBZpvOpYnSjIHli8c1eoahhj2d39L6jyxgPdYf4dl
T5xL2DXC+cwYDEOdSQpkpryAx0/W3k1VniZ8V26/nrSVIrK8uRDyu85ZFxw8a6Xh
a1fqmieZmSvjfaaNSMp8I4R5MdEU22GgNhmGP5CEzPF3sw9tbbkvo4u4qWeUXFhB
gVsp4ETM14rseG/xjTf5MUeMac793GLk0R4BjAZjReJdNEp2PNCS8Qoo7j1g8LEu
rLtn3iUf3v+OhbOcK0SX8X4vZXdM6s1U/9bNeEDKHumXBR8wyvjgy/4bYs14pun2
YZtv8yUWBIjFVPBTnwwgo5a3HRysGRRCXRTN4QbbqzE78+oYIHUMjadOVE1Bza43
Qog1f9cR9BlQ6RgwjOc2xMb1R8BH8y5V2rufQYJz4xTUguintNeE7ehTTP6nwmdq
VqO47nYsFM/hn+rRZ98/U+JSsM6fo+TaY5UwGSUj/htybUzogZOuh9Si4Y0/6T5S
qlVnFlW1iNZGZGtU2PZt8SfYe1kVC1I9RinwTP1yRmrFgqBW3Q0i2snSp2xoNVC1
HzRpnoDNgL4CLUJI/vwPF5gUT2rZ/8joA/u3jZKi1GjF3FDht1bpJIYUglEsG4TC
ExWlr1nnoWe7A6lBdiqyrowVJkzljsaG7QmG+7+OFqCgNHM7Cpix4qHMfbjVbSCE
UzgIUsmmCmxZP4/TQakkYMBk1lR9KpvYx3I8rFYqbnoSdD3n15WuN7hfZJxiGMNS
cjcO6X4MyRUU1Dv93HZpHpvZXs8fylBGK+CjWaC7bvD+2v9+P8WMKfqwCZ2Ts8Kr
Andmf+iZ7vwtTUlIiAXA0poFUqoTi63DauKCW62T7S4RaXHxSYA60ZAIN3OH9Vqc
JW1wWx56W1sDIItW/Xv3HLncoM9kF/OARBaTT2Y39D5xiNFQU3Xv0cOmSXuGrbxe
VwzVLItL0Rv21jMIXgbOPC96wPONlBhTXYLakWU0KtzHL2PgYPhku2zxlsq0a1Qt
KNcuwc2TM2Y+no14vSFUlzmHdWhEBV5aRqJC0dgHTYgtlVbDucu3f4y/wEC5WNPN
hNcwln+/svRyv5dYRFFdQNacmewjGst4/16VazHJNgPJnR7P6nAhlel/rEi93rdS
Bf3ARh3eWNNRBcZki25NJ6M1/boZx4xC/d+uMeX3lA9fV2mzF4J4TK7T+ooKDVxw
L/8PWkWfv4sfd+u/qXmlsRCSWiPgpfaLZojm6RQNJmPEtUPBS6BWUJDsKX7TBluC
ChHHM+F+/z24xs2j9OvOx41FvxHCTGQ5NxjUA1pwgPkYMXDPjqGr//S2P3Kw7bEt
HWlftpw7BNJ/61IbOKzVIIgerhLn7WweeOom1tzw9odJi1WhLc1JyCkujcXEAgxZ
LcKKGYhFtYbJYPthHeWIJkUGiKIZ5vaCpfZhX/BjJ9t3S7PWsOBvZl2PK6S4GI4e
D91kocidXxgjHNSjRj8pp7dc5ARpgLFq5/h+xdAkryv7uzKsjV9VUwC6ttI0772c
2gHxXIS3I/oaQsHrGYlxLGQHF+cTaLQXwUeXnOOhUPJCOWNBnFkS0e++ntiVYcC7
YWDvxQLyEHpYfBqsccTTv1mr6X+eKfwvVg+uEwlMHZf93zR7q1n1y1PUODBF8Vll
KNl1LU5SVYgwh5Lb+gx+0ewqmtYBokeLnaZO4ZS/0LqwTyKszSB5w7w5jPLk0RNQ
5UHXq9bvclOVYxgAZSBOeL3HQ+9tlcfB5Mq9saydOw4OcmQFdb+XAhaWvZ96Kcu+
U/xBM/pGf0qzur/961RDt9YJ0TK5S2hBoIY67djs6Lze//1hJSR0deo2Ck+ovM+z
NiC3FWJBLGGBF0WTdZKupBGpZpnDXvC5x206+M7vqqXjY6mO/OJCQvYM+yhlw5yX
CmQNY30HUp+tB4FKw5jdVJqqumt0Eja/tePfHyoqIYxt2IKAk98TDL+e5HW4RXiK
swg5ElghXu2YlmlPD3jo5G3wokGn1lCKWEp6C9mPyE5DB97nB2p0aQ8WbquIyIyX
ggKZTaYWQW9M5K0ub1mE2vSVcra/USqGI+I2g6SLypf3iMfDchCdBwhk2lC7Xvbg
48pf0E88wmOTEo+Y2UoQUDVRxw7XjVnjvxoypWJ2N5o3VmeaH5+U72P6SylVn1sh
lHdTWbdsXS95CuJji4zwLEwtZjD0JaqQEThlkkDWuxTKfI9eagT4gre+UAsqegur
sNZXRC4JWCH68CJzD24brfC7oyoMzOPDvBm1rF3/bEwEUwdTPwi09IqbvF5ZWtgi
+hHlNEclHPS3C560Q0fj577vfmXkOmdiztk97NwKKMEP2P0jBlHvpfV/FZPp0tpo
8FKLbxq/BVq0gGg5fiNCbgxYUwEjLnY1yxQtGpODVSMYl5sjEMjoKs1GyDRQIYuF
UH1BLOa5Drq8DynwMwiQ5FoOT/cSYHSwNytgMWofHvb/FQBa4lsQRNKcQ3JScXjc
LSP3DOO7LarYVLMF5eyymknAPqsmTtTP9tNyE6DQ5HxTR9Z33Ak0mGISNWjoBeKU
Xv5BlkufnqrJeSviudbZL7MCbX3oX9HWNDdzEjhsyf1CyA/wbm001P/D3wA7Vrvu
I733vaXB1LPAMocv1N3Tfm8ZZ48kH+M51jApCunig0KjdXnHMF6hWVvWK7PJyNH5
FrruXf4GaCaIOF6iyaMGvfKizR2oHv2gR8zeTEf13XKfvRgaVqER3TuOjlFrdpe6
nrezxDwKqJM7FmqLUJ7moN4v+R+0p/l3CwWGntjjaTUATqyaPcW0Q10U+puTSOrp
+FnMugrQm9u9wmPu+Q6aJEMuKZRRTxoFt3tYejpTCqutC9TcYzDNjk43NhuM5PvX
WI6TbRHJWq5vRiQKWnoXegRY0wG8L3/aw+ZXq0KjOr6NQkl9/Q0MoMnKTzlQkzUJ
af4r76wo1d6i8Qf1yy1UN+VAVv51S46ciPH1WpzNHhI7DirvoM7sQJJdEzJ2Ldgk
XbdBeN6Z7WV8m5yDbi1S09CQpYTa+GGFfMPjWoar7KZVdP2l8lWh/Fgq8CXIQI8E
FJTVcF4oKYPJ38042NLvIMPUNZKDRPQCHKY0aOXxpFP4OjSmZWHVkfMDoAfEZxDl
5Yt88GVHXy66LMLIt+cq1bkPtVbI5KeBEk17Uq5wbTLgUvn/l43r8pY/WIMMumlY
VE6wgBowNAdMhQr/Gb0fACkbRROXbnQ6TwJc1L9SgI9ZGiFaplYz1TTcjJvt8qJE
G+OZmCzMWg4u24OzA+ZKmEWzJweDEuLr0tAfko1oJoU7EOnGG7Nxmnc1iz68+F8E
WriErWUxIHMq+p3I3rQF5COj27ix2kT0xcVNdeYVEvieGSWg8selIOCZRpeEQqRy
hjuBzoewayfr6cDRC3RybRKWyEyJXL+O3dydnxtokVzHleZcu0Qx/9XuB4A3003I
PyCJX2+cR8xL2AWAI/Nk3h694iljmBR8PcHzyvj8S+8gDDQYul+qpPOz69+aSj/c
uQdInbd6B9It2835eldmcFHVYojxgw8P5/ACWCAGeOW4crFibgLUkzPeGDdKr38N
a1pPe9GdFcKpFLOeXRMpinBIQ8sjBC9J2Jm0q3lACfQcL8H9W9snrq3WrbZ4HfjJ
rUc4eKoKrg0xMZjCraZGCetEPkZ5qhoQ3ENqr2YJ+jo4AA/eENBaWb02qQHAMZ3V
ood/b9frqcHIpxtyHojXqyn1rykqpKD2ofGcG/kB2JDqtWbgKJoqy/fMdvp5c10n
G77drOge5IPgFAjE2YJeN+4hI3F5OGMZlV1iXyKfqYfx6qu21SzDSII8m+fOkLUE
CU0FtcsUIXaBMLj0gyCnD9xCXYflMVr6+cTb59wUuD/PhDBiy0OpBrdmKAKIfecp
HH9e4u7/XMlydI5kkJKmcVXlh0xuRXkhKiiKZa6UVreNLaMGXddoI8wGIY9Fphz6
9q8xmqtOaHlMTaBJrH/ctUBrB5jJQ1iAX+DLjGic12i3fEwJsxFD0UbTlHaqqOIQ
qt80NBmE6QS2wPK59i8qm4fJrGrF4BtUqdtHDKBu2anEWzvlSW5zPmEAopCC3tWb
VfjYMQTuX4sGBK0OmhvI6cGau5m9KludE/XeR815n41c+Z5f7qXCPyZUydRDprvH
Wck2QoUjNlxWIczQM+EpoXngwQkvFZiaEiKVZIs8W1ALGQsyC6UU+GjQd+RvLQNC
HWhaIIFo3CdH+6+3FIcXy8AqK3c9d+kEy7Cv8AZ4woY9Si0vnKPlIb/dxaa0g4UQ
NNzozqtS/Emn6c9/NxYjpCVjXo7Lt9G0oQObJBxRSMecrKxMsXysoVzQRznzLkrK
v26+zxfxqzUb02Yzq8R6hfcqAiZyPAW7CqQZ6FeQjjOwyR2v21vdZn9ImQQxkNQS
sPy4U7wUNJ3ONpMwmJa+v1seQqn8pRvTxIXeovCZaaVXvxIHjqAgoMsrqa42NLkn
wddqCpEMrr+4206kBsxq0ma2toWg/fyCP5fEYN6jwZZnd5rIlD2jIjj6PV7gUDVo
drjq+jus76/jERSTW4edqpYgG5I303fCvkWMVmnhSWSD/YlPCNVyAocakVjFSGWj
PON2jPm1oy98O/ATT+pBF4HdTAdCqMKjy1UUurN2y4Yvj58Zbi6B5CjjS4yp8k6F
WxUJo2m4jNwtIfBq7NzUeLGUc32nU+6mWaRU/fPC1lq5ZJqnbrar6OSXrlIFTdkE
EpBArsTslNvUdIuJsDtOqwJwdG6Dlyfa3JWuTqXtXLonF2qVMvqB/iKamFJf50fI
uACN8LM2E2Om1ea5PPcSFZbMOXtzFuhEJDgyXe6XHWsVDHsOJkPevp1CQtpbQrnB
I95t94uo6KNZKBerWlaEi0Te4pheA29y/YjF4Fx3sEvmhUFPgdytIq6tiAx4JBuz
fKPGZ9FJM9hGyz9FZS6b0nOp0ZAcsZ6hA79qwQbSeDaRs+R7Cuxb4h4MN0iLNVUb
CJxJDNWHIwCd1ppbk/5UyKJHchMbQQ7e3tvwsEFmQlBvlyu4Wj0aGeCbqfBuwvcr
INMPW6SEODy3E7viA2CZK/Fa2a34OPl3O56giJjsDM8Q6w72eF4P9RCGlHYsaCt+
/4djjw8Uz5f6dZFKHVy5JymH9atqJXO+zOQi8aYu0D8k8KLsLrZejZiaoOdCpZS9
9AkFuyfFDi7+sw0KFxP8XWcWugTsUy7zWWAQCS6XNDxs5PPQijKgsjMbYqzZ9Zsl
K8BpS6pyVFQrE5zGBkizR5brqS4cjAO3pRauxvV/8QhCF1ViR9BMT09bkAZAhitJ
TxXnJPZXlfCNd7lMc4f4c3bM/KX5IWM3LpvoHdrakLnxtyjqZADMVt5+geTnWrOh
l8l2dTZOg3W/LzOity+R03fGbcLGoARfeGprnXeiU8D2QW0fhDiGRoNUYAqDIfD8
/dEVq6nmNVRyeoPt1PUDyjWxNxnwpI5DMRJH0iKDYxmnZy+M7UvXFC4ZJvVcb9Vk
EOi4W7m33pU5hc2M2AcldkShXDovQmUEY9/pfC3Xe2LwLLlZVmQmiV6kzM64g/w2
rIIig7ydUSA8p6PLztCL71LN5v6XrdNOf2Dmjb4Lksn3DMj5oXl8cQvZMaY00+fD
x0A4YoE49YOWzKLG/6UNwAxzLgrNFEj+hj2ALrmCsKocv+q6C5/7+DKBvV0ZwdfM
GAu0NO3y3qAxuGPdlX05z9ZbWhAhcl6qbM89AXIIxmE1KDY+2o9FMoRUyFXd4wg5
mBuGEFiFfniVo0lJ+vdpgWdd8rXe0Q7OAL2Kdnf2Voe0U4Uo0S4uTcEunF56uIAD
lVAqYfRcjWWK0Iuzwpj5VKec/y6NycsGm6v7X+WSbPrsMh53aa6U5Y6HkcT6xP+w
QQt//Mt2fmEyConD4RZhz3HQC3Fcwv0mWQH1dwR/enP9STU+Rpu7VyeP4rTkcmLC
BDvbbE8Ne5wti+//9ozzLXv5LROxbd+sgQADAaC2zYX/GfFPMAGIMRuAUo/tzoEg
adgryBam144E0tiKVJuACFphbE76KFT+L3JZ8ka2icLfcNoXt2nyPl0xl/A0xQr7
n+JjX/dSbyIaGm+ifjqyyp6HceyNK6mARwMqpjAjPmzG53HGPQaJo7iolvjIeC6Q
0G/iC4WCd4Q2diRGdI8Mw5nJZxsiKvHOziuGon9gAIL9qdz1/Oq0RH4nTH08EDQ5
2sIm/Qy0s4pkOadBs2HsAh/G6y5EOvofUSl72a0crfTDip/6MJ9qfNlYf0uwJgGU
hfD6eVSWehgT5JmeybAG6vidhTrG93LQYU/MHQOzPvcuRQeoewmTOWUhWHkH4xnM
3rNesKexjPw7ctM7X0yRx5D5TDUGuf1lkPozYxnsx6+d6Ho6N/LENtpHt7aC+YzE
I4WYONqrkujV+W3iQfXjNrh8mjHmYwTCDSjIN4R25p5Og2Gg6qRSXXCcI+a68wRr
Mo8eY0UbPe15WsJwVAVOFbqMNChTOgLJqaWmlgCWOwRXVefe5MR78bW62OOfdLSP
IV6/uKvMeePckqXYWzTE3wkQQpEIdkx+ROz3QB7r2qZeprz7N3m5ta4klPvJrSBg
/XSn/TNFc8+MU1+WHOovZSjKa/v7EtbO3FVmjVWjkJt7YaaEcG+gh5ZChpIYwwzv
Deabiqwuc2KMrlr4B+mPTUZLkx4LzDhgUymh6YcrweDS+rxJ+PlFaYMMakaE9Q9J
aayVGrvwm64r+3sIf09OnTvJWDn6rCf8fcCot9kHy+OjSDTued3+kcPrpBlrqRcG
qNuRUAnrtgVOg3lQ0D9Mwgyxa/jYjZkXZXoy1s7oQWiJgcKvcJB9sztP7fZcxn4z
tNOlPD2vCFfNi+g2ItVUx2jyOQREKxzIbKteL3wRpHagIsXX5s1aeLcVhiCrbCqt
Z96gzyhAy/PEfFEuK42uR3XS9Vsm8mJPJuXm8ZPFvLp/9Zcsgol9zcq20RrBF3TP
lVt3xm2JmoQkFwJG1ALgOXRyZYGcvfPE8DIKu4Kxqq24Q8hYETZTG3llhcgcsrlL
QO+2IFH94dHeaN1uJJ09z4olocAPJxGiHnzbfWc23TrctVY/vKCOAii0c9YVx4ZG
JyxTvCOWt9E7SOLoHKo1hxVJ2x9UM8fuqI53ETRZAKQHrmRdO+VUujPIk+exYanm
HRrqgLlMwbHYVO24XbsHiR+eUCmcSxJctKCYk06HpppnNoWzTZitdWJ6sS55I+i0
SHNb16r/VMF+d4/CGQ4EF+lA46RdveimPVY3SX92NnENOFsos46FUdAlg5YgcgK/
kCwLiziWbHmhK0ui/3U2sLzISHvfVGjTyXskUBWsMeqbnpzcDKwYoWgOjnauB+AR
e12bsrWipaODjbVJHhLnXK1ICZ3YCscsTC/SU0LmDs7GhSGUTgBL8GfNYbEN4dN9
oyx0BWKnofpWLYEGxri/2hav/mOQNufGykgs3967ysP+YzoEUaDYSTgbvpfYwjJO
hkXLnYF+qVb0EAepWt64tNcMe4j+1DJklvmipWz1qSNXnE1ybUolCzKyW5bgRsJX
kNQSpEfciOo355LASCNQwSvTMkSLvizuPnP++6nfGEclEQSBrPlRtB0NkXzQm43q
iGyWE/dGxvPmQq2zDMhABpg2FGSLd5DQn3ZAQhT+Zvj4g1e0Zynk7CTHNhaqTCQa
cF/D1qxpI8IcjVgJd8UI1M5zB6iTumzBF19wSeHHvji7uruzJrG3Gkr1m0j9/JZ7
j4Kp38FYIFeAGewmFQvkXFCy0tWUsbNV1e93pFwOlHyv8VT+dkOHpw2fy1AlegqA
sblzDRbygeA6wZ8sDcy7iMnP/+nt5hPO2QVYHBuRg2rwBX+JickukhnXZ3fE9DX7
CdRrG6hVtXIWee6QVl9juAlQwgUTUaXEGhINifo7p1SaCc6NEM6Qp+vcb5ipnAFN
XJjmp7AKxuhUNdU4n1dKEIrKKZ0ZYZGiRIAm7NpCWF85UeCfLxRQolhXBAyPgjpP
OUNzVCRoOA9hGRqmeFVMOov5bXgnFeNzTDXYrELQYKwI+UswzzlJQsRJgsVvBMaM
+Qy6HbQLJxEWZwpeHrJR7OhIZIYxD4L4ZjtsbM4A2cIxhKdGy6zfA24XZVPUtPIF
eU+dHxqyNmiq+HLcyumNivhKYbrHlojROVN62v8PKACR9k3F+W1xkzBlCAre/PsE
2GoUw6/1ilOGFcnk3+0szALVFfyXi5EGaj7Ehl3P3Y/x5XtzjGuhTuMWPQ3G4Xbj
isd6/98/c8qIaZFWeOL3L0BkKccrbmIAhLZvS6KMAKwWRr/nulXjFOsLD8D+AjB4
9sUuYv/D3BTfFHxJli1aOl/oRiUn3gZEmRXAqQMnHbhzf2p76pvkghcBChto3Amc
vG/IDPoJlw8heDKusQIez0qid3pfcmwQL9Dcy/N+mA+juhAR3zwmzB7V7ezh3/Em
aGTKDxuRr1NP4b2KNJTwzmeQj1Gna6jALE/2BcwGrrAdLFWrBALPA7csI+a00YXx
jsFsyYOISnkEu3pdOsl3DETLZnljnknlzDzHhht+Ogpe5CP0DM4LzJTgffJzIFo6
9gQ3DNbZ6ppsCXiw+Dzia40wrtvgNFf9ZtuEEE3nS4yN/mGGY50gQSH40KsLElHz
grBv3yShUsRVmQmnRAzGSiN9cOOXYpP5vSKPTeJ+bobbaysIWv3pK9sALpUZlSDD
KN1i0cuffsoumgSRPv/5yYPCBZESyeH5txniaYw0CnXrlpOFg2Dk6J/KOdCUB01L
AK91nboQn9PQkCRVcx4nL4a2AZLySpO77IK1tkUJdMDQzQ2xsyXxq6ymdp0P1AL3
CCBO+dFlUpOTD/P2C7Y8JZkp8J8iGJT+7uFO5VZBvyyl/jzMTmo0aVySZWZ3z3Qj
bcObW/RHp0DXMbMR8wyiioZW9ksW2zKrJOs39Pv0q+s/UZE5Mo4Ufo1YKItJ6la/
9AuSZU2Zjokez1BDB/7IXKMLqu9/VejUgcOd1qNugkLZHZ3O8NaTZgMEURihO5n2
mN63ZpFcxmKHQt6yDx0P2zVJPDbjijy6k9LiF5cfZd4jgwVkTeMQZoR5mpkzx09/
O9rhh0a2NkTdtst5yYhyFvd8r35ozXcWbxAyRYRC1PyO3GTdnovNxD5KgwRpTGv5
msnZzp/jT+EgP0us2iKabIko1tHZnEpDT7xhINeTGOkF36bDlQBzDMeHxnAFi2E8
O2UeQ1YtWGjDBY32XxxC00n5sBGa3faASgHWBQEUklXQkqZAYx9/vBd0/vTzB37a
n+QtBpRdNmFyCP3RsSJ0RBhhdGKQ5amjqBrmOf+jTsHtnMTmVnnkaQq1HaapGeQN
DRaGFjDCdU7bVTyNqtceM8I7NfNtcHwIM2Z2u/VCys/4KWfhCF+cwA5d6aJ0SIOY
9Dt0QNKlmVGQk/oaWdMSRxZ1itUkaa7s80dTgzEjG7lihbakhlul4+8BS69a6meQ
MkXjBKhjhfCxer+eOyzl7X4bDSUFkiuQ9MDlI4i/0f5mpSqwYUuCWxNvbwFJcbzV
Lgj0lxAXt6RklseqUmjQ9pvtWLtQsoasrmmunj2hFuIwIfMdQOQvIosrzX1EKRgK
9rl7XNhXOnIPar8puBaJ1HecXlSuI+kgdqE35QKokz7NQi7zY94U52huW1sv7vN+
zwwlkmJz620O9wwSw8Ck1j/28cFcoyCRXCxM/4BUsh0DQXWPxLq+6HBPyWG8xuJ6
K4JIeXBEqcpIyGR9YmWXz2tu8s++vM8pDpmSaRaKW1BzPTYPFulfLM0QpTnVrckm
V7OANA1myTLZQU03aZ/l1xym4gnEibPwa2ZbuTK0GLQtmkeCoamUXeaurhhPkZ/0
i3J/i2PJTjscWYUV6T65dXPmhuw4ZEjxu9QJFwZAremWzUeaBHAJxwOJUqq/Xfzq
Vl54AjVeppieaNNaDtsNnKP7xNQ3eD5atVrOAKH1/RDfPCJSGPPmDgNM4kL2MHtC
DZD5bNZ4FKjze+NYcwQRVBPAWUTQmo7DYNHgKqJK8xZ4o5cSe/6NC65nyOWBDv4O
7DQhjBvWvCDExa3P8JKn6765GJaDvBymk+tG+mC3WtIGyNg4TZDI8dCwyGX3zcDD
jdBGW3vDanf95kK8vbptJ6iUOXnB9CAqxnY2w7L5tY3QZt3BBOWwl/7vsnM44ZJN
8Cu+y0J1CU/FnObJ6+O0rSVK03JsOtEYwZS2MSdrk8R0yQfVfSZBETfEpY+jrjYK
r+0Blyz5lasiNvHAnUGXnyMJtMl7Z0Febr06MtarjVuv1Uzbq5kl6qaMZAwPLAfX
E4VgABZNPQnp6yks90ITqylQrLm/YgdBVr27wSdoGwW9EgjKyYoX54PCIXb4Hh+v
b3hEK4CIQtf6UQniMpQZefIJtX19buMruoRfVgBFk4qoue7kJ3drw22Zi8I5+TJI
W+cGNwBkwYQKaN9plrdle7EV7yPEnh4KW/goknM2BcTfxa+bjfPYyJJercIUmUn1
iwfZYE/BL00UdATW3+JVSMeZueAwkwjPcgZxRrrYrlM5Bsk4cU5BxA63F/3HDHsj
3ENZMzzcyf7ZUZc0o3ghH+KXX1tB6/b1lkKb4a5OqrQHz6VisTNlF9OEQ36eXopH
8qyGiyEO9Owlh9AKVIr/qN76ENlEZCGXp+kO6t8J+RxCgpFrIW1oxDVCuGQovSc7
hQXzrwEFhSAv1ODxN0qrEer09hsyKVRmvgJDCaSNsvOoWyeeOC0c6i2ZSVVD8Hv7
VQw6aRYI8KxFLOl5GbnoP2kaAUuNFp9BOWLd9uUV/cKTIjp6WWa1VBLE1QNqdza0
K5FMfpgleeEEeBKBT2t4sktnx22nBVtzygWKtNCB0coPP5DlG/IPzBtB71eG4pr2
oxptioHofJtCNf6Cg4cu0r4JiON1lmbKj4+9btPHoZkWSfpXXVyQ9uoSCKIXH9dQ
9y1C3KtxKS93OTzfYvFRJZVcUT05ucb8+og0DYI0zSL+S9B4x2Ed6rl1C4QLkci2
fKCLo9ECI+FYbfEclu0tmIZeZrU6Kwq2/zLJPlysK2w0IyB+KsgBHb/59shgH2Zq
BWwHaJKevDy94JDLkzF22oTFJC2HX9MXJ1IMh+H2iT4rfMvWM9TS+CX0vd9dhp5a
9WA/g0+c6sDbSDeQOebtK/A65QYdRD9F0jyyb0AM2B5ReuMjk5N2Y3B7A3sNLWYj
Isd9ozLcL9ZQVoKpuKoNDUHiTP4+4vkoa7DKAuW8DOjUFQKXxUG9wcCeFvAZbqkh
179fGo33F1lGtbyv2U/YCJVxIUZ4KEA05XUGJWTNEe/vKTKD4fcq3mG0AdjNR1sn
Lf/j9GmDGfVp74MVtEuyyvYzrMz0MeBYOxc/ZIhs6Y4mn+6S3RL6DIxTcClbyweG
+b+/BwDOgm5DbfB/FFSIQvaQt2xTnYZzZA8tfTmZs01CpifzQDavVx2wG116TP+9
I0yqKdw1vaM0E4Sb+4rEgLGkigEDJ8FMjRNY5LTTvt+ah41EDRevgrgj9vAmg/JJ
LLA4Iioa5qaTEY6qiTTkH8u6hjKtXxZMSYGJNge/xrcJ78R5mDJNqnhsccY4Ujy5
esCZL1Tb8auwSlDPUKDxrjcXFHPYByhpcPXGsnGtSRCSREUFaB9GchmcmsVpa2cn
dWGcgpTWoHCg8xm+bQIxXpZLX1YAdqAzanyboPnMFwrxTvM7pTBlUb10pTV4Ug6L
7WHEDTT9ti/KeusYuu7NyRHVqg46WptmnVIiRBYi8JFWxamOEG+Tn9tvGc4+dkml
EiurZThmO4On2IlB/fVxBwtOFrBe40Fg9wJOD7/Amm0fSmB1vLofFY1d6Wz6gIL4
ISIG10CJG4lr2RwkZtAIC0ZQbJnRJ0d+HrWkzO1SsWsp6KlUzWTtqiH4o3cYjDc0
hLJYFebLje/YF/IaplVJ4cel05JLyy/Tqo7qml0QLIhQh2MRVhRQ98gTrHj6qFdG
UoUNm43HoIHuQpQ3jtA5ncKXN7ZUnlBgftb6tCAyXxpgxGEpHYzB+ix2hB6gfcKT
C8zgVUzxDzfJAEn7iw6JV/SlrFVL7jWiq5V924cHaOSq6qEoR4uV+HXl4HCdrhWG
pwiXo0qnu3cTRRUTkkwkI25HrgRw9h/e7EdCJ5kalEnf6MknUGVyD2712otq1DLb
NIY80IN6sQPQiX3u5HXZgL0gOricgBjloUp/WQkzL5LiR2s8S7Z/1Xj9OKTP62Uh
APKAop24Ko9MtLAUNB32PJQLvcMWGThp6wFLsEOTIimH5Hh83eYYozyg49Gzf5Pw
M4WnkPV3fOKIHRTfh6ANF1HT57LW9HfpAaSqx7N6l+FDZgeutqST8+Q00nWQtxPq
POKHCwU/pILmIM7G9fdPYCwkV0JiPoQdMxDjW6RcM0ili0U2ROy3Zs++4PvsjrG4
ZX7vdyF4vEgZ9pNChSU0FcWnNUAf0IAELdAsvlPx2e+/bsx7ymRgU002T4JWJOcf
aIqcRijFRPlQtI7JamlLdKOtyzwSNeH4Z0F55me18qu4N64f0a7utsw6NvFbY5oY
N8pXC1SnMUlRJ6fa93RtJWWYQBD3XrsxjGTtfWdqoB7W4JkXwChJBFATNyHI6pKy
rf2Inv3fOxR/Dwa84Huhx69ocoaG9J47P5yiMzdv10Gd3InSRAAJLEBZWCx8RID2
Hz3EOJKWUcn+Lw7T31z5dfaZxui46FoTXCczUhqBJxy5HIE+ctfgxGZycL4VadFm
hjJ/xQLU20pABFioEBcik1pcwc/McTjbSQHUHWaHipmKTdKrdY4W9S6jo+2js06J
JLnoBLW1gN5Oq/mPDgeGR5IcglEOT5THtF+kNU3czrjQ3+OjnUXwX6K1TzliguZ5
z6FQN95dKHt9gXqTTFWeyS5nGDuu32mwCGsT9clJBrEg6H+oA0HmFLLZLITORAH2
9HRiOfrs5x3LnArnhUn1qrH7wv+H50SzXlgNte1NQRB6EL49HdR5h0p1VM6QrObx
1dfP/qCeQor5UM5lqcNbf2E9ik+ZV5TdU/DOOPDV+PdR2ki2PTREnwDD+7cjzv4u
HyuGTFXMl+mrt4Lm0yFV7YCPfrHn/1vriJ28QbDD20UasGIG3nerFY5UgA3WgZc+
pCv+Ex6RkO3rZ8i+m+LbSGtJRYMvDItIpWEWHbl8j88/iMXnP0ehJjn+DrkY9/H8
1qXeUSkR1W9VdRcnSeOSXjBheWjmd5oW3HfuYGfjYQDpdU6DjRzmVS6ct/kKydwJ
cV2+zCbQmUrNEvbtifZ2ujCvw1cMCN7utTJQVnsqTDyqToZxB0P9zxqf3sXv7Ziv
Jh4EJg6jc/EtQeIuzPuBc6ot59J1LnByWPBjBbgopXrkYRfqZB7vXhAze8Np3p8r
jJvvaHl3SyuOxNFOvqm6WAn+NMireJjef+IfqpGoc/vy6C/rqEFV7sdW9Ra36AgZ
tb2yvQUp2dpoLGVGgcUcMZg3htwVzUMr19VnuZ/He/Osct+fp91xiXcXQfnG43E5
+IfEXe+ZO6WvjlQ3SbuAWoh6wlwgRdz+f53yXSo6XPoj4UzbPuzEJ2myAlI45d9x
U75NPsupPoG3u5Xq2LzjnNA4R7ig6oMTDQEw/vgZ0i8gynsqdMMTpaEYH5KV42Ou
YfaqjXeu4n2H8XLFAjNnDGCdwn8BbOsYujeIvpTG3l1X5l0yafTuYHC6LPkapszy
ihXLuquwG8X+y/LkFcfmYaaFdsN+pejPyoizSKgfNkHl66iwIeiaI4ffGfzEioJ4
H4xuEOA4vVjBySNFfoKaVArpV54y+OdZOT1dZFr45iXB8+Ko+5Jk+KJbBjh2i2Eh
/RYytm+mrHj0FyahDv8VwdY0VpZ7Aa6cTu2Ab0gJGginMjpHDIbIo6qyqnD1lI9Z
3QxeQEz0vRK8bchzXBHadM6dtC26iL0x8A5YtwO2TDC6LEJyKM/QiC/FCnI36VvV
0vWm/DiP+31jZIM6ftq6ojBTcoeChRZEtnhjg4WZXmgLfTiJCFJCyNe1jJkV58Lp
l5tUpV8Z09i32AAvtYAp9z9fNB2gHp0fAqGaSRrJQQqHBQ8o3y4hTh4hx+SzORwU
LPHMl4ial+77KIswQ+U7i0QpUnkrU46Nv6GeWMBIeGtYD+lH8YuITvJP/Oayd5UY
PXSqhtzJ/C77ZjlipOg36dastdYAUvwEShGEQRt1bMe/y7dZREBU+B26wDZyyXUP
qcjQ/eTQyfpP/xOQte/JRPMqSy32w/gUH7C9xXMFQUPLrohFLbKmvCzvr+1ftbmA
OrFydY6Un/XxzPZiBQzJEYWXfNaJEjXmkDEcOgZfCIhntqPJ+UBJTn7n+Aw+Rg+g
GN1hfjMZakDVbRiLnRLs0w5V5q659bjDLmkWlHl9ksNEKfeOnGY6YgkSZaS2z97I
QppWZTWCSkielel9P3YbSZFBOxf99b9zw188aWGC5WTx2ex9SBwlN//2Cy+7yA/5
ef5UQKN+MA8V7hc0SZwFSn6gZYwp2+boGswEjLplzoPjFXNPWw9/YTUpvMtc1eru
WJP3+qcag4fEwE/OPjskGf2Zg8d1t86py32VyrwxXHgthzfuKCXgjQkfgGU8djAM
r52aO5wCo19ZhmRe5hXUb7v1b/oBXb1OcYU1mlrTjy2FxArTsxDeRSby6E/S86Uo
YJpsfNzM1LgQ7OykOPzzb6uc8LuA1mx8TRIm1gMZp3GSvv3/am9IfIC3fkjCSkSI
Ls6gxyfEx2xCtsEN6yLe4ouvt6RecMKOi9qKXCLHfwcoiqWJbR0TFQHDRfjfZqEP
smeP8FN23XXSz5D44PHL2lsIMw1K9oIr6pk4KTxyEmo0AFCdcl5bqqAeWxI+dDHL
qVZe/Hs+GW9kHDt5NQXlosBVmDJxCowij5IzpIedpgs+Etz0+T8Wkeivc3uYzzLY
UMMPNtr9xg93JI/wzvlC86TvOuYzJC5HMxypxdjaXnrCBctwcPMqpaPsF18s/DyY
k87VTmVOxivpbnJoATkrgwYMp6rMgBz4t8qw1ZubueYnh5fO+VAZom9pkIy/gd6U
pMOnOH7hFnRuxnrImCfX6Sz8/fkkwerhGfeYMMwUvvAFfdZZiEpYYfjalzS+iIn6
ktm82p1x/KeEpHQ5B4MxjLSSS0ccncyXW4Lnv8swSTgMboQRIcp3k25CIcpgLVvU
hslx9T3tAcBt2hptdLS3yVnZfQ/spURlfZfTofS+eXGsHcEbyXA//0yRBjPr9DSj
JiMZGMVlK27gXdGciaivome6KgYPbQ7f5hKTvcFCvOMAtTngxf0pv2HGTbXZT4AT
oNgaO/5WdbGyG2a2dCVqrSHwGYHvlNb6LGA9RAUHZ4kmNsOLOTNxgppHzp/P20Hx
/x3mP5/rLnnr2NvtqxhPKpKHeGcRHFHomtFlzbiCtrRk0E2voZwArLPJnlxt3Q3f
P6UmDsbQuXAKRKRvamFKvWT4IQpuqTamC3Y7UhnOwOBycxmuQ5nwuGq2Wd45O6XZ
R9zIfOBuZvQFZz42zGNlZ54juKzBE3ykMXFImvTJUdHBEVIchHLruHu+Xd60mHEe
cydH+HbOSgS8HlFme3MYA7j0bBAt8sGpF1GnJK72ljdcA9NMGExq1IhzJxpjwR/s
OKHyTj8B2s+3tWy155i+66kv411MnHYE3NoFYDoN8mM9N3rfYTvqkYHgdKQ6vjmt
HXqzj23z5JpBBo2TNioYdnBm0VlE7joEF5bqHNl8tlL5BW/sAp76L1q8XFcTbz8n
npMog+RpdS8oqyjLLEk5zx/gT/pAycrj5I/xicyZtEGnfqwLlVdOe2SjmakskzA9
I5MqpkERzlZYncPRS9wja/CQ1mN2d9zJ5JPH67bCPyAjDSikYkDxddZ3c4uFdGuN
T+lO8gUwi7m83PfTumeywK9LQN8JNhhfU8iEwrSfbsnui/0vZs2dHbmROvVrJT4Z
1tIgIqPZjG+kGNV45h+9T9LSpDOf+wfDgrKEljNpC9sTZxoaYtzn8fC4cqu8haqu
GMnalSq8VC7KkqPGzF98qCN/ZOQ6n/z4q+DYRgwusBZh6ub3eLdfSLO/QNGyzTqI
36hnKnE12kT3jaFQQt0uNux8/U2nxgcnAXs8xQLDoa6Y4Vz9e4MJiu8oYE0lU6yA
L46etxLMMU2gOyJDw62R6hKii3LEyi9SwCOYEY4kaAc1MqIarqPdhg65lRbW5zyZ
R6lWdgCAuxqff3Q+6Hu/FmpJ3RQJ33FhGzTCcwM21VC+YYCltYbD3netEFcM8nAm
nJlZx4Mdr/fvL4KXvDfn0gVpOzSFFaXCqeNB4sEpPm0h860st6Ex8ySFzq1M57ET
1f796ck/xPqXEz0Jk9Rpl1pr3fdpXKTywajKh1P/deEY9ILULnDrJKU1KMgwPsbV
1Rd3aZ8V30Ty5J4NgVIGtg2eYZBlagNA5OtPLALREUUW+9U4IJBU5DOvvF5X+/Ab
ZHqsiD5h7BqsEsNb7axqunR8cfdpqcI8u+BNZ1s6DhtB/eylNhh4vrsolzmySX/B
0tk/40kpR2tvgMwuncKLlp8/Oay02DjpKK9bxZlOx5WDPdc+VBj9RdwZCGHzR4nL
dw9zhui2hg2WdFwqsJbAo0eQkRAUnqjQl8/XCZXX2T6a7RqlgjwfC1V3fY1Pzl9A
P8zsZLlHSw+IVkNm5rO2pN2+BkSUSESfGdauAuzWGWr9BxHcWAiVfkdAvQNOKw6e
Uj7zBaR54bNU0/rpATJx/X58ZPTatRBGj1A62U0GyhUM36JWCWmS2HVHKYOsEske
HpaJXfXBtufkJvT/2AbrQvr2+YgE2ZPdFqtsLpLUQYg2pTXH+vswxTC5izrRvBpc
JgamFFlqrO6pwMlOr1Y1ZSyGGef3Ox5dgeG7AMK7+7xKNdTqMy4HDNo2jAW8cZPu
B3lrzZer6pmBMLLQrsETqGHL21gRvgy8EtWGe5RbF4Ty/PtQzP+WrULovzJX5mHD
bu0bh+68+Q6E4On7h9m3PWA/R7kTbXjlju5kEx9BtVxpYBQJJ4kGuO9ARkZxpWJO
aDfBilmg0+b2jMpcA2VwNev/xVw2lkIYyOc3u+hMx1buTm5edTmp4Gr+7Q8eZmh0
8hk3FBi9yZoVsv6Kt8o+9tK/YsT0kI3RI9EHc3JEN/n+hes71siXXP6TsTVPGnx8
DofNqCFo97d9qIGpZod/s3Sa0WIZw7jnzwC82Aqg7gSN0dF+bRERRyg/JkrByc64
nh6gxCWv7uaFvnKcg5UFVo86V5S11hoq+5gbSGjg5Q59jmdsJxk1cdRLtTqLf+Vt
UUxGRxCfEQqkdjsL6e8ReF0JlAZW7vbXEQ0LpAvBrpafmBKO2YWSM3d0D8dtIXBk
YeJN0Vxei8/VmicH+/Jzu2wSBJlzhvkLjD7zlPx9kx2SrMf3QiUjFzFhBE3z4R/x
Cbkuzdnvied1URVFwZNez6yxdOsmKc7lfPy5S9A4kBUV5/3zp+RWE2i1jKefihNX
4AJNjZOhVf1TC7oncLdn954TN81wDMu0T1iqCInMzX/kCLVvlos+N721NI1fEzy0
t7A+QmWCFOfzVRONYh0XGC83IWaKfZzBvqimtRYKqP4RDFIgc3XRpxFDiiVUoq2u
XXPrFu4R3ORfJfApZu83gXrMvQvib1oAPIomZSC1RLurnnLbOgJqOECOlEyikQlU
JgD8STV4WMEPMT6MyHYTWzKL5Yln8mg3lDlz74d2U8xmMGDlY0VIY/GmRTRx0ikv
oFylZgw6KAk9zec8/zTxWRDoo/TGXZaSXwYnp2mna5o3xjwPJjkmC4u6tqyoSMSh
LPTv9yKAHtx5xAothQ45vENWuwh5mfC01irdTnX4BD/84X1Np19QqeNkqkpYRrSK
+JzOQocElQRwsUoyNOdokV9qMSt5JROH1lK1PBiZnj6zqn7cWqQt/KIqgugc4t5z
0sqvF/l/XbMMHyY0kgV5DwI91PltuxTfuJ8wHLuJfhre7r21Ci0fyLlXB+2cm20i
pJn48lpuItIgNT8xD6Lb7SpZZrzmBoKQLi8as2OcL0xzImfEAuhLyx8EUQBZU+RO
UsLDOXrtbolJMoIluYsoQFhJGDbIONQYLW0+o/s2NDEAoNyARX1N/DLvRc9TTtG1
Jog4r9Lgsl7DVwPUlbj5w33YEheIK/iq6PR6yUkmLR4aAHXzrGgkKHo4WLL6p0rV
NCgxuNJp+s1vH/6Jx/wq5Mw8YPU41cZnDc/y0YGctgKxgqM6wByLbUjU88wh257H
8YAVeEA9sva1iK0LVlEgD3fKELuqCslXpBbhbPmiBggJpg9UPCl4arPlNcpToVyI
9mf8nXxCp1zaOdTR/IEDqy92iCwM2+7TsNtCo1BNP+/5L667NpG/jmmEiNeUfyBo
t2exjlUazkNuvWBiObC7O7meZSW5QsVXq6oncFg9v4hbFDqTVhW6bY+B8AgngU/G
+Cux3j6mIuT4GOxlb3Rhyd1lqwLOTAXD/qI+bzi56xaqQKohQpQXBbuV3Q6s65QS
Rs+fUwEQChsot6mlDxjJBllncaH0DE4XEDjJuhXEnmThZf/wn5ttnlHWg1el/kwp
1VtbjHZXo+rezTRNCqgdS12B9hEe8ya6F5OeROpIyJmFDKebHf9PC0xlC9GPP+Xt
Cuz+NCalxpYkql0n5/EzAi/090SiKzz/63Rcecm3JqLWd9jOTJoKNhx26SiLj/ND
Pyf+RHZkUL3reeLHODMksUOxXljGKEztcUs3m5sMYbF/wo9n25/nWGpmKGWW5xUI
Szn8pW+MbCqvAUHQzZ4TLM6Gui35aG7KrFHVuyFf84S0Hus2AqlMQl0eSPY/f0cG
nmx7YlT8FjnNfaJ1sie9hCYzloK0QuSJZOpSbHsqi0Yiqfxkim5QmFOzlksQXYlJ
JV+8CH9m5wctWm82Wh63mMCHtyItQOMPzGmKgy2+EjbHOReEOzxYzVw2s+N+hsxt
HJxvBibNigRsC8oEgrXMhtFe22UVF2XMh1tNYNsbWKXhHqv2Sxim6kz41fctjLmI
krSZOphG8N5Io8HYYEFJ24ZemD/FBVUgbYh5ifktPUGHnBi6cMjbRN3eStu1otZ9
nVgVHPCrjEMs1GQnPp6hCteleQpVO9COKRX+TDmovv1GizdzaMywZs2J99pdonYk
CoGUZ/hiFxNqDsg9PkJMzhijFd90rb4MpSeq/xXZNsBdjZq+UFLULla8fPbyZeMS
mW3FLyuBrG8crEj2Oa/Oj+368R1yu5tMHDoAvl8bdAWwvbGQF6eAq4Ak3PdTlDM2
1YhL2IBsIFf8kJapfANjBye5FxbXpecuWTmL2muHo6tho8SovIR9gbq6eStJMRkI
3hV26G1+M5b55XJ3J8eUn97agYgVzg/P6uAbG3lR/zOooPlbuj+b2tvEFnrMKuiV
xPyVEXH8zhZ2pR9sGtryGopPiku6eZWxRJlKBAGSX3YAKDZEDt8Y+GFGJ2u6J7hC
5eSMYLXCnWaiaytx5+DNaN6xqMEMrxbLkvxMoYjsKPQz3ghIdS5c7F5fjjuVN7JG
a7/xOaCM6lf78fjR2FghF6gFxy0l4ZKBEm6W3XlPKRHLMPdOtT/rgwRa8LQ2oQDG
4uybZVjm+uE7Kd9ty2g/HH8qjepxBmNa8zXcLywgjvh/pN2sdMkV4cZuWyPuucdM
VmirOJCQWg+FZkIHX8JGdYBkzuaumzH67dfmL4ecfqYVZ3XkAPfm3jz6YHRD28t3
upKM6wvuzXYjr1veS0VnxUtQSpNNM3O+JZh+Yz2gUNNYCeACUrvaEM/KR2dXHrEU
ps52fx5q4OS/qQ1ar5cvONIzVnzltOAUKLGdITy0IZDBX4APTMgQAQytqSdrc0Mc
96YZRP+b46mYM8n8IwSm3eFCsWSbRuSSbZQL7gNC3YpbyXtsJihnGeyqWtI9ohjQ
QJO78sCW9+NjWXirPCXjhyb9k8KoPt5USqhIIjOlvOIaM1t/bjr3eKhINve31ppl
c1G9w2kswDpNVJBeztDlAI5EJBv7LZj0KVsBMlwY0Ny1HAQB2DkJntlOi5twlINa
5YNyqEYT64SamqWBqaWwLXmelRkh5ZHxPnlLsDs9VtfUvRUwqImQjSvYTG8o+VgD
BS9Xc7dMBFZS/UmpIZD3QvIj+63ORA07k69XlfK63QNcgKl6Eo/bj57vXRZQrzvE
KBWEcpZkQwPLbwjZuaLR1+Du9aqrTePWEmsWWufHt+ddJ8KMQeo8mP78Q2ugmOo8
GKjy1V2A24/CVaQfJSne+wI+OIgDK/K5rHRYrVzf+N8v2UQ018neJdDXJl90FFbM
FbKSI3sjLqyh8frr6sx/Xm/TR4A+h96vAbtMFPetFH7A9g1m8kikzK+Gw+0VHPyR
ZXF3qYBOsaKP+LFo+fhTW9QO+S2D2HuaM+s0Sbt3S3IgIXMA7sgsxKjJYE/510A+
YfmCRG0S1xc+PlWw6YuGOI7QOlKHc7TUqVB0i7CRfix1ZcSq2OxNP8/JwHcLHIcS
99i7ht0qasiLWOUMA9TpmUul+RiFxk/minQtF5Yyfl8TIAfOXaTmAAlq9tUdO/9y
kKMAV6JyUbf4010GxA7JqfTr4tyJKn0VoYuR2f4TGkxTYMZKIxouqxIIx18jOJ0f
6QfqeGNxBxyhV4VSjJhd2+DRMVMQXsnP9vgUMr8BlwgN5K8c4UnuwVDtp24k/C12
klfJJ9qotJjzFNBXO1LYxX8R92NDG6rYGH0ne1EEe7QkiT2OF6ke7WlM/DglcPmH
yT5BnIi6BiPViHBKF1sBYtziSUPKXZjpTCztlUPjggKZ6Rbj3Tg+mJtXtAv6EcbW
mL8/Nau3PIh2dNDodsTSwyY7B5dpkftaDre+saRHNbuiqp2fSK+IhdHYgQtXJJhs
hL+NpjPhX2tU4ss3k+LT/31ytRuwLF86XHbjKLOHNw9JZFd+rGWgOBYdlbNTHol1
Z90U3IoL1k3yUFyF6Bu8Fb4y3hv8cAwWE5lh5MB9nVDwfR9GDM3TVwPRGGL7zQop
ZIcnjtsea0tWjrfAgTK22HM9YF5CSBz2ZDQBEV7L1D1yYK6nacw7TQ+ffmswUSYU
KOPIWf/55r75/YWGDcVnMADQpyFhYM+vMbj9kpMZCx9psQF/sTXYTzj8xVDRmSuR
5WJ1BWIqDrFKvp/wbAAlFTDDPzQ1Ymcux9rh75PiHDPMnnYyN1NZCj5YEh4aRjP6
MAkdNTK9EQY96yXTVbNDaLhx1PV8+6cjE5tpg3jR0MEzHyZKs/BFbZSt/NtCWK7J
QVuBTaaQVyf6d+xf2SBsRJ3n7M4zG6dJTHfgEEr+1j7RIaLvKLZkevcuqxIMsuGI
5RTBDcNI3V7gRAIpgH5h+KLnQ5J+UKEBXG+dP5wYbWovmznGTx3VuPnoFXxFa58P
48XmvxqTI7ilmxKkF6Rwx2N5ZtVK27xBuKkMJ4GudezKEIVlDD7XH0n8odK8voUN
Q3ATiu6zAILmPZl1PT9s8+5iSY673wH8PP4qcic5TFil7tJgS5RXijpuXG+BZJPV
miae4UcWQHbTQXKvsBBWc+/hdPc3w6E/MyZ4r/v7sdEkG2U4yoDeuTH2LgFLtBxc
HTdlG6GJjQhYxUQ5NBZRNEqzsPA9zJx4K29FpAo24GMkYZvsYA2974oxmDa8fDoa
82F1rlgtMcVVdAHo085xpmxxyu6bTCDMAu9MEESrHrm+J69WuAkTPLPdsHFeUcZv
JMsjkl32I9cbDzS/9tVrATf0ECV3bFoZANMy1ODKE8p09T809+kgzP4YsLXbcudo
norL28cXLI9knZIBkKT1aOjTrKmk+xcP2i+fxqUUj9BKm/SxzxZl2f3t42wHZG7d
NPWcLmUahb8EZi4olSaBO2AdmEDMIwfZVLCUC/LV3mXDV+cJ9uOP+K3nmiQt+npJ
lPCWK4a2zAs3dq8qiyhMFwqy8QjFIdk4w4JXrkKzDbQ4F1hAQK26jeLqZ0Bu+Xum
bL3+1Jwbyto4DkuM1dEet9f0bdO/MJPEVk+eYFlaYcmIyjTHM1uhpvHU87cXB0Cy
ssBJ97WbiRpkmgS3qrwYVUGQwheXj7RGDnzkDpkSfAXXAGlKIPzneOPfPsjWSWR4
qKLoOM0oaluduV6s2f1LZulDLg/Xw9VcuQT34e5QqXPSBNq1bl4+vp9Ks1cubHod
47+q61lCA8VtChvNMjDg2pspiXSxPNESUj6h3YE3QWy1EhEUD/fS90ElKV8xcO1u
B+1jftdF/7zyMN65ZAsoOCD1j75fhSgb45qcM3vNwExDPKmdU815t+IRW+xZwowh
yHxgQK8+bESNZUX99e65bjCOIJLmp6xj4X5Xj9WHEQzmAuiUAT40WcAX7/ODm7FJ
Yld1mbw7zkP2k+106OF0b/kGX/MXkxe0Q4DiFCMYwjwrtyYHg/RHeyB/eJbfc3/V
KpSXl/GdHZPOafciyXNIrdbewUX1nOlr0qnvaC9fz+RM7dP5m1lXpGisPsgqKH6s
8+HOwdf2sQZY2Vz0ErjF7k3VjYPHaKw15yUBPLHt0wDJaMEgExAM9BY54gYrFdmM
OesfUFsBCcm2kZiLI1hfErjdkc1rCcyhwGlrOevBmjo9mEUQZ+MvRmzc9OocdowG
OrB3LbCqkL+9r3xYiHrmMzO7jLaDro1WJw1iptR5tmHerkgA/iqmJV796HiXSgTm
rvb8tIHggPypnRN/k2hhYj+I1LQ5CZTcu3DmQzY1/Ne63jdppRuYvcW0orjf7vxm
g1zgXJacxTT0EL3LfkyDFyYC3WhCIB682fVpcTM7P9xuHaZ7mHu5RSl56cb6770j
yIRbxDuEOxJ+mwBAafkU3khjic671yvWeFKWLCgG0xu1f5XgA/gRB0VAdyPstoR5
bOD7Il7KatBBmf4PzPrlS+v0M8HM8ysNI7xW5cPHQAN3pBGmQ9FtBuB3/f52ZavM
OputRrvdHWABWURaAj6KXe8QAZv9350nJDML6G+L0FfSNLHTyDN3aFyqGR0LVli2
y3dtCxhU6SqqVgZuS4OzqqnuYMbZ5BwqaQEMI9CntBMftSMIEXVReKFh3YAzKglA
qQq011Jy7kDNe59ReQSaZUR3XWDtyRgXdQCV8oNv3S11uSA9GPoumrtswbfR7oxW
osOowbC7O0t5c9IHMavd6LeNRtbHhrmtCnPboj3uMKMMau2oFVl4TJpT1TcMu44p
mqTnhZrhq+C54a/l2AYI9DZlz08WtuYDaAwM4Z5ThF5voCrha3f7dInR5dWV/2Rx
xiPNIGpLJ+BX7dAKWDfeJ2y0Pzjmh7hQv4pA/fJJLC/Su4OpewsUXjwstCgdDXPb
zv8yy/9vgL9Xddi2qqb+pGfy++ZRBhSCsS/cUs6wCzmeY1Ujp/zEECFpceLTy5Gu
QB78+kRmmSJCLfzEIqrBuLYvo9nBQ7LY3uDYHQe8BolCdw5tksow0RxJd9v0tYyn
B69icYIqA0vi88qht6zWzV/pmipQKDiOsvkiUUJlugTevoz/7pr1FJMo5CyUr9TS
koCEKlE84JWG8y3YU5T/ccYM3onwBdBhJun1U0OpVHMJtFQdB+blIBCcQLU1z2jW
w9zMjUCdDdeNPpn4VINYRX4vOwU4h+Tmucf3iTv/kJONYN48ngXE0UMAimz8Tqp0
kuC2AjYE0l6mjYDhqzbUTssagB0XGrhgY26TzJET4KBhIvos+PGycvfPYz044PoR
ptiEJwbb3khZqN4DmGvoJ8Bu57dA4CzEGZ7A7SRpXDdud07kt77HX/bywBi7ME82
uTwJItty4HlQxCFW3y1CpkE73kFICvkdKBDJAb/WgcL7Q4WSoQyg/JovligeyWzA
tvrZlWWlByHZ58CL3oxY+x/hBIFiEG/1b88fZfiVF95DiLjfueNK8bzXKOlRo1T/
F8RFSklLZcyAeVv/m5o0/rLtsWyTtM8jav+dzZCOS0sMnRxOPahSed/Z0LHc1gnq
bPT+XNU1RrXZ0YHR0P1OoE+qvH3FFBSAY9cbK1ZM2lGhH8gmpj5brjhTX268T4o0
avbL2V1iOIjPZf+7/pr6HPOdPY9ai4W0qq7oHuGt1w3/aw/RAsD4NmLDGBn7FD46
1LriWCGDNavyi21Lw5GO0PvdAMLOCQOQiaCeQ57C8csBE2t5JPGEzUYQUQaqE49p
ffANLCFmNeQ8wX3RAoiCqFDWuFZ85sZjDxsb7JrCADFf42q1Cqkv/D8oN6mutGDs
qLItcPSeSYcxgGDR2aFe4o4I9UoSSLHIhwWC6GMjpjgNon0qnRx5uO2/rPGKsMe4
7QhC2GZ8qovNWSj6DrzdiPYH3tQ0Nwvxm87K9uuao/qy9t3yxHf/Bss1Uc1vEUFZ
GX9DOkX0GBDZZTJo2mZzKAI+0lFHQ5hVyi+7L64tDMBI8iIaCoUGPlqmrQGFmNPi
lwrrHPjU2B1HWA50r9NvbF0wMExlAT54J1HndU6uf59AenRg89H2mH6YrX7y3qTY
5ECzKXAyr46pw28bNaUnY3eMSI7CM+bpQxe8oaia1Osbv5VYolSKwW1MF8DOzOIt
/UOoOrROuQ/Di2dO8UXRmi79GJpRfdC28czHN2WnYR0xNWQrugw4Nsj2+baPNhj5
NMjXHyfPnUD5uXC00vyh+v3jMiqTLCVZTsD7X11eHZjTCsIBF3IK50btyNOvIA/e
/+WeS1Y/AtDyCL1KjIgG80mVdP2WBIiqp3ns/jE96rWuqxCyHqtu7qI07P+xn7yw
n4wqolgHtUEz3mTyZ37RPPFeMfyKXCpEZ8GMjJ8mxCnvWFVNv0rnhCGIg9kM6AG6
sMaAksxIQzLAUi+dAFuHm2sWAQi0hJyTM0NJgy+ys/kdXQYXc/uoDwvycgAVru3h
vOhRSsPYqiGfpOB5kuU+5/Y9b+98kc1hltKvP641EYsqoDpNWTH93epA2kP2Ae9r
BnfQCr3H+h5ievV1qLa575O59BOFyt7nf/MknPFq1sgQMi4V5SK0/aG4DMSYhPR0
9iK2VFh0XKH9tNdpSHT8Yy+q4vf8BadyCTlb1yl1oFNF+/Mhnkh6OH1pKSl3d0ra
G0IUNfveTs/h9MYmr3Cu6UOE3zRCkQEC5pa3QjEMSMgWOWB1v8JTChjMGX6fn0tw
Zmd9sNIOpui0rRdGRkjWmMbJGGR4lEWpcPjA6Q/zsJW2dczMSRPsbh2FCw3LgOe7
gHaMuuZ8N3aQEmW8RiaLKarf9QKqi6uzB4gOt5iSwDZDmRYB1Q1IOko4c7lsF1FO
g9W3zAQsBBwqazzVBM4kffqnbUFLr3ZogygduH2xS68KkS5e1wtD8btkAKtddoKV
aqBPZWIaiWh7yXLzWudqK8gY+VK8tw3uxFkiw72FU+BqvsRCLq8a4uQ/yww5jivo
GA8BJhU8Pj5J8t6ZBkgGByrDd+agE2Wikgz5Go+rBkXK3akTywZALz8WZhsvKhlB
aAofgs+5lzsrvQOKY+9TdqOSTW3Nglz0QSws74orWzO8uX2PFgv6k20pJL51P6EA
KYpyfqmqEI3thhR8XT2SzV+ekDk23+Seqwq4h9OzMB6SE3wR5Bb6wzj7bCaDnqS8
++ubyVzx01466qxpsSqdAbt/Pym+EETfWEwXv5O0cy9L8RzyjxuTx54qBcpX9sFZ
FHMGbwkz8YGqZJfzAmX7dFhU8ZjMQbbi24CvX4PN3FkSiX6WRSaUQFSOBpxJNO9g
PXdW5DH5Sz4ZczvdUTPyZXk8DTQu74G29Trwxtqd8Bvc8AaCwspGNDRebw52dMp1
tO+SzuMdZkawoTPf08C3aTLa+mYTx2ubm2eM5pD5SwP8CW4BKiPvzB7nBghDeFrd
LpzwXzcRs7tX/4LRS7AX5UfHjjA3ZVxufeIusXysquhE2FMt3hgCkTKFrii+Imrc
MQeJs45/R8hJ+9sz4E3GDOsXG2mAqe+G1CL6x2e1VViOcmstogDUEPlF8FbWPPDu
fyqeUOpNutuLW38BdyjfKgwwvLggzeHnhZJQwrPkmMEdAmy2J3mDup7JhKCbmNvH
K97clmV0eOkhuG6BpDjj8JgUWAdTSErMtzzB4GNwMrMi+pZRVanbHxZ6pjoYU3lD
nFtNxHp9T0gbWCvf4yGHO5dgWYem9ea2hqhqlM4YB9f9plwAKptDQ77GqDYaHYLi
BenKI+ZYdfucdcav2px3JupMd4QHEQWj6eVK0BB7PH9mKQoGUKYdYk4iVUlhcvzZ
4qsYMTrxMh+qiWrKlQoGzMzLop7T1qzI6H6GBVcM6rx2ozfZfa3H27FDz0GlTpJc
12jCn69/0IbPmGvQqE2V5/BZorHLUbnzlfCc5vNTV1BBmf0mfwLJMOF2yuXKu/Ja
bK4IAfXyfQaAuhBM9bvpX8I3Y7Y/Xsc3t6YMOhRxrKeHb0TREvbnZZrVIIWT0g+t
J1aV7v+34ZQb/hCYT3yNws2WBqGGLI0tNx3WPNnrqCYpxf59Gdu/SxmgVbKN70bt
lS6RqjD12+CF/kNE/Ivu/kUa0yLPWAbh3KKlygmK4A1CiDic4xg5fUS6JalMJCqn
j0Qtv5EBLcWvQb5P6DIkV+mja4GTCd+r/8MZI4mDFePhodbIywV8C2M5HUoMwvNQ
cpAp3LQyrX9jYNnsb74DKQ9S0vBgoP3+FeUhPwxlIZKt2Vn81nYEOU0qHO74WylZ
W99O4ccrHSSlpM1rcor2AvkTKF2kJ0J7dYfwatSAIDlFRde1vaURWsihhuR85DI5
LXBLRdOxrG4i6xba+UVL0MvNUgeYHBDERggggoqjkv2TdoB9+fXITPT0oVcvd7FN
VyrM7EiuwDQo1585hnNq8/H6jOEuS85D8mV7S/HNRZX+1F9E7DkWPy71eZ8UWUPY
ByKMq0VijxxZkVRsYwdDZTVtOVWVnO51b1HcaPZm14YIHOFlwV+zNDRYAHLqW9SA
V5UtACrFkJBwy4pI2z2k84GAG5SKKIakNu84hzLXeiMPilY4o7PjsP7EqLMsdzb/
KN4VL2C9i+Bjb6rerTdpfDGejI953DeK4Rr5QZKE6AKLHib5m/qxPSDI/+h70xgE
XqGCAHCHmiUX9NDJDGr5V6brf2YzfvdB9hFBRj8tw6gZvY1o+tfIMPX3Mlb7Gqqt
nvxKMlrXRJV30wVAIRsNoAeVw6VbpwIwrHiVWYCofmkU5rgkV/WlcR94TnBcg4n/
+LkbOjK0JOuJ0LghtvBGDzu/rncwa+ERjkPWZfTvgr2tzKI6f+fbddXo9OPExrOd
cKENAqmcFSX7mS6987UWojf+vNDHs+86WqkwdPzpQNdfsFpOhjlkoJp5NMdWc771
pFlSXnT/s5EdoAjmdwjYIUFaiieqN/d5IoUSE/FGYLLj2Xl/pIQ3TKXcnX9oclWY
iexWhQE80OHclb5KZ0Cp5Xwq8mHPkkmu7IiCbMGsLsmwb86DFWJdr8M+aiKio093
LDlOtOv4wLl8oOnRcv8e90+3RgI+66/ZqsLUnhFjFAj+w1YHAT6D3idgtd58tXeo
OxukkXzLoMDY7lcCc397u1SuGm5iWtVBTCHbu1uAf8wrhkTIDou3neD9fxGu1Cj8
sTE0w0JiFCcX9LYqmmE9tfBs7N6IMxEpE7HBUZ5eCdc5Ff1Ts2hpmmiJS4Cpw0gw
qnzuXIG7dJXuG7kpjbpGL52sdf+wIubc3uHOp+kAYs8rPVfqY/QDibnHh9GE8KWJ
dysprq4Hf9AjFEWus51CJrKlhVSC/7K3GZLu/9z2pG0ulj9NYEM5NA2P3BX6ctwI
K2UA+rww3PogbrXb+0arPABbAI2IWjyh+g9N7t1mG4wKr45jg2nbDDpZDvslKfDU
eTrudbskP0bPhzKndMEXZy3WL412dQqSQddzqi7vUHFiVpPYy/OQ7zooMTjEuuOZ
7EbwgdyDBrSIDKb8v4uTQh8DfMLSB6Wr3/5pynzLhUD8bXQTj+g/55CfKBLiNzG6
0v3o/SMhPzQBldbSYu2Jc3ZV8uLlx/DfZ/uo/aI167wlXejpNwkonlcBha2OTE2R
akGu6RqkPaK2+nbOpjE7zH7KMlYwitVQwp2i+w0AqmOpeG1HBXcEhk15haaljbLK
I6z3y/W4/X+AOiJHNrJ1rQ7tdjMe02jxcu2NXYSqcheyvS7q8MbTz7EBERG7kRFE
sId9RTqdoiouHKpuKJo3r5xbWuY7vf6xXKRYUlpTcM6kW+AyDgYaH1jJdVs/ajWT
xSjUFjodaaQIWgJRhUsvR67r5crNV3kDjI/Gj8omI5u5NuJYbWH27uwDgsQ1J+3Z
HDZF3mWGvaScGT0+5P/Fm74xAgW6xr8knfuSDer6cB/QH5MnmIsu/sUazll/bGnz
MIpb+kSJGUTGWmgBbRSApYjmLxiFlfS3zh+fndmUOE19ffNK0u9zqKfB1lyBhaqS
CQibkEBLbeXw04+1j2VK+cI9MEZHnMwaBTzPaD/ukT+xq12cpieJeQosb1+yocjK
/uHmEerHPak1+MOgMFTqganzz5Im0W27YNwp0fE9/yIvclGWg/TD7GUGRthsjl5r
yG4OSNtqH2cC+R7Q3hSeDEk/RLhq1gJ+gwQIWA6Y+3FxeB+3H3zscFe/9BPmCQy8
CD8DwP/mnnDrOejfZXYhDbgJTPnP/S/M9BHsAD511SDz1DXomSTVdgmoJ03Mi6hY
bsOKw9Zunr19geGFJjRxcZRL/FgwoBT719Canr0cNS8/wGu6GRcuNnI9fkc19CmV
DouaqFG/Gr4vPowZppG44T9zaJIGzahPZHyCIkBufa992O19ZZ7Bz8VFH7ziUNkm
N9YgGK25X6jpMfd6Shat1juV5xxLGEfINyoYfYlX63Gm6+IiqbIXO75WMDq5ExG6
9x4m6Eu8ijpNd5z/NryvFpzpXCovoJPNqKm5y+MmU0Uv/O0ytfjoFR+x2D1OyOGj
tYvqpJLn8LNewsmTsRdpkWZL6m6NWhID19FDZSGBxk5+2o7ho4xDpREr3WZvodn9
m5TWMWwzplgnERIza0GlSmHHMeMAKiGXr3n9WPcPsr33gikurweHQ5bBxyn9FyA2
6bNJhJm3G/RlBD80e1L5zeBoaajpsCJDCcQsyyffclOgIRSArQRryVXvmPBBBlMS
88k+dRTmHzsUmZ3VM4duMXlmDdki1LOhRwWql7pv2BU1RWLfeMo49rzW27TTSGGe
xyr5N5ywCQ8tGzmMovlrz6aOvCyHS3DCNdlAmMrcrd+73Ja2KJgptG/Yv3HVvZ0a
KqnW/hP3F70nULbhxRj+nMIBRW2aOZyiTZ8JWHVDiC8nOmhsL+dxKiHz5/ElYJ6L
TsXv369TKjHoxS9iPA0PpMbTydVRPo7pDWPjhdModKk9xAX0/Lr9RYFUq4lJJSdX
ZJQ6u6b9e/BSRAnVQjrmtqDb+yW54K8IEGArKOJ0pvxiVu1xHmFp0IXKGcwX17l0
a32MmCRs5QDCI62dJ+z0iOHUT5iGgqNcbBuKbzOJFFiwHrW6IAkfVylzehEMJnrq
fNLSvweAzaRVxA5xjMoN0UwvKk5at6Wr9puo0lQK9EJ+g/lifrldeJrDwum/L3j7
Dp0lfumYoaP8Ipds0FZFtU/wDPmTkPjrhU1oUXSjtjjKqReMyxkVHN+FMAQf4zp8
fQj8xXcfAV4Wib/8HvUZjdHc6fJgMH4ikd76grMl8z9pfznQDu2vCEIRSYCJ2J79
p5/iNhP3/O/kn+Rxt/z0qP2g3UEEUiQkL1lFhJ/WRYIhFut1WxPtfBSPhVLfNHXy
4sGbkxsHMaZ6YkkRC2z9nQTsboejpXYYYrsH4rMyjwDbudr+5YQvQx2gbKoWR8jH
lNi/5sGFx0QJ5d556dFEndaIFchq5cr6D/ZdrzgHt9z3ZROA7z7d4kXcZSDIKp0G
dltkayBbqrm2wlzMWXmt5FdTGzVkdDgfdcWLbCbNer8zutAko90yveBStI0dExLz
M8uBgFadHvapeBm3RL7cPRD7mYUYLmDVxFsqJa1MK0E8Ns2bRDPQ9ciBx2PZZrCm
aRhCSRcLxcMXpwdkOMTYNZCu3fLv1/piBXtkwtXiuRVxmMBIM6GSpVwQ9k4YKOD1
cPdCXT65BritKs7trXttR1criQo3M39Mfg70F7Rwbvw74RSHrjchXKCJAe/A6h8c
Gp93Vr12uewZy+McqTB2K01lK0o1lfVIyuzoKdJ9Vdj9ajGecO5Py1L5vDOTDs98
6g2iw+fwm3Xplk1uUe9oTKhaSOoXISqyRoFIBf1Va53khNvENj7mshbDGcSmMGMK
2IfYKiqfrx4IS6BuZw+qYk6RlGVxwRuktMy4Pm+aAcfAybmBl85awQep/CBZo6pj
4edh+zaTpVGbiD0Wd2DP9CJChzY+z4B/jvOeDoLGvtY39i5nLFBcC6epXwLUIZx9
AmwRmmMKCIjH1zhwdCu7QUZM4XkShlg9Eudig38gKkq890IOYSisouTrLMeqVh3V
nGtuxkBEI4dO7L2yhhSFWHPyjw4XkdLgwjYGIYiRWJpo0Aeu+/A663ler1r6v4B1
9DXlz2hQspzbQ5Ffd7WpCXude6nwm3QukC4sAoIpkNhMD5vfaPpsyNeiGNTqwPYE
JsZCPn1t2/eNtvK9h3l8fPhJWSfvnD++X7g9GmIPqEhenV38Zsb6J8f65qcBaOv8
NYJIFW3HGjsFgl9R2IZyNvfJIRRbMoDUF6XRUmEj8aMQc/FDV4rjAgJycQanRf/v
88YoVaLc8AH88h8g68qWKw9jums6wurnidDXuMw5a0/NrxL8Ts6xz2I0/pcDHrgR
1l4w/zgLwmzCvchc+dAkpDWzLwCurj35Exkzfa9NKeU4OXsPS6fAiBZGUMM5gvQn
BFc8twlX1MTMmR5hmoNPFrUQ8MA+KWnrQR8+6mc1hmoafBrLMQ7oZSw604C6DQSk
qkyKIuEx1WKk3jAcO9GeoIXJEx+SEjri7tb3LgPvMxyVWJT3ORX6dVcUsK53PoYe
eA3tgu7w5l9Igv4VjCjIuKjKUGeorOkxtp/Bb84rXik8LHTGdwgjObQx4HN5Oj5O
1Z6lvNYxjmKCm86z1K3BjyjCYWK/PsPlN2qET+g0t1s4qMReTMvwDhkP6qgR5TS8
nvjZivPFQZpmr2cH/cz71gd5urW6G+8Q/KiEFolgjsxM8oaMFrWm2v/5ZWXqdmVV
aGq4TnaXIbSflx5hr2lrkvd2Csoa5MTsjpfPo7Z2bgAgxpPUWFCKNIfnRcrTSGcV
g0Nrk9nc26ecsiSZXa0BZF+GS8hGhPzlmFoxSEgp17wE1PBVKLD35jkBF8839u51
r6c8gQgmMAsgQHyKGD37rs+h3lXsbimU+P3DNpJtfst7IIfS0cdOHPBTAPQ0t/ZY
jOGFCCoTLRq8R3YCxNlvkNky/BgWW0NDdK4cjY9cIFrrvNenBGPxidnEywLGp1oO
cxMbhr+bKQ+xJWyxHIKPQe2Q6WcIS5U8PI09+W1JxHVcz7oUuu1EwiVKvdYRe31N
zmITfzzb2PChvPNbTAZMbjEbK2cCl2cT73OYRYRsSDsz2C/qAQBcp5PKGnzFYqmz
jBrz1wmIuvdmApbx9pa4sU9CDDpv4fAVmAZb3CF26aqsvPzlGRnF7hip+ZMdaJrQ
8NE+XjBWEcjkNb2hhTf7/UPFsSS3DMOd+BVFfNqLMUO1Hl3+jqJL7L0wYqYEVz5I
KOo6GCYl/J4DqZMUGyv2XUJcrjPQZnUbzXVu0FKAolzTDrdIqjcel7tQ0bXypR8o
nXH3mXC4PV1LQJCDSt3opXgmcBx/1UJs+5zlHTGGztgHC4Kf5mi7r0u8G53fcG8L
oj4ex5pPiSuwd8Y4XWIgs3vZ3E4sv6JgpQDsvp0fhDWNLLgvnZmqJqTgPXxaOV8q
xCu1FjIsBWfY4xLNSs/Tl9r8zrMpKNZ77olUqDbDI9yhUnR3r0lF9yuxl0bI9Kxb
frNaXA/wgGsWpWuZTlCwuCiImb3mjm93Bjofq5Mk/MSggUM30zvzLzcARmCxW+Fi
09/qqTzFAv3ax9Ob2tWM/JHbdeeVbG3vFbTNRxa5cogQueGScGi9L0zC33RwcLSs
/GxyUdKqdgekEHi2uTH5qsCg5wO1jFiG/b+TgcN2ddVPCaVazM0hU+TF9Hbud+KZ
xF6h6BH/f6uBjrYT5r+NMx9C9f/Mbs0hRdOGCJ6kFGd7HzKAmhCyllcRpEb5NAvh
1a2LCDDmKpSH/xJxSScXHo7XBa41c/9KVi7IFFSN05EK6v78a8XvprMo20QcVeI1
bLFGMnhp59qVYYf08hNypHPUx7/z952HvFA213E7LQ45ZJRE4U1hLu8LBBa/p77O
fJVOre4wkz7WnK5AONOXfeY6tF6T3IIncv7u2CenTQySvkyzy+ikrY5zt9WsfarU
6qtNE61ZSYNtkhz5sNISe0X66P4W236uNyl+EjLSLkE2+8eBAxgmoY4ULcIZSwsw
SEzOzM3HY7oMGmCZha1cK8Fmdv8ZIN7hYrICELwPr0HTpxciYHbVxpq6NDrjnlI6
c6KvS44y1FDCd+SFXAI31HTxnd/f4a8gGJ0zGzqWRl7+vnEzaIKHBkX7wan72bfv
pac5qayKUVbpSPT83e+AY0Yy5vgdiW2URhlZLHxLTYlsG8vnxWNbyMgZlafGre8L
ycCEtROaE5Qc/CWnLY2eakWsQ/5drSOl00tY/7hY9e+JgiDIzqWUtaldBlDNIlzX
z/AKGuf+fhJ80AoEQh3ql81Xlg3QAZ/9wn66P2NWSgD2Ddtsmfi+K846dcD33nYt
lPKZU6Yhe8Bs3T4BH4HSt2MrKWihLcHmlZW3CoKbjcjAQoD9W71aPIGxyidoWQmA
9D1zovii7JD1CSlKll8YLvQ4G0/kyhlUC16ZUyEoStOl1QgWM1WcQxNayMLashCb
5OIX/9GpZUai3UmJ4SnKBAvJ439qTtSwAhEbljXValpW0AR/Iqgfq6EJi13HDZ79
2fjNy/wGaQaOCGRaFjGzTtirkVjr9dHmXTwOoUFNVoGXH5xQwNzi6qMJMjWjV/hY
q2EE8/sirD72l77yMS+qK2eHmJ2UmLJRLSYSTH7FQbOMqV4Jrt0dg9svDXpWpu8w
SFO1YKsSopTKBmXQwjTO0/Ihen1Uuwt8LWW1WQdbzL/kMtN0l7Hs+G/OnIY6cgHu
s9VGZZ9W0HumR43NLpOTApWMs8o2FKwF45y/TekvmDWWL5eh1u1LcE/0jeOoJZpE
FB0RG4sQvRqn+B/ehYG31Ku3jXVf5oC35Fwp9W8ZHzsNNDcRu3RQHyYEApDRunk0
bvgBmFFBQKNx3K0XCebuOaE7+0fEOrLH6tQHJP/zYQLfS/lUSbQNznqwsVuEUSTp
8P2pHnrumb7Q5C2zXjOe8byEs+UJ9PjPKjoixLp5kAENi877jN+r1+Vg1i2akU7T
ehfJVJoz7KBt/JZOrAh3oUgK3EfhkZj6TKKsvg34vUygsfbBWk+AWy3x0ysTyB1p
gmNpRBnBdCq6TmnZe3tjdPi2FkV0GBH/dsY25qtFA4rcjfie+5opvTEv150/ruSl
75pSe689fZIRf41hDhKBTFJ+vFXmY9mQsV9UyJBOvw4akF50bNm+kHV3zJjbJ/dB
ogNdbF3RWcSYN4ZSP79S4GO+HYGitAK15TljzUbeCZku2QnlZW02q5UCYbLykFDB
+DtNFB8Sqbpfz8jZhtROM79nUIudthzybd+Mb81acmamzRl1tWdIkJn1oQmF7YmD
c9oL9tJvXl2p/dldPuqiFjCPNWjJiiun+WANlJGyn5sSG0xQB8SUB+KeVXAFi1RU
t2HXRwTDM6EME100FWwKCEsfaOe5PU/UpLQomUftKhcUnXpnNpaCYC4BIaxS7cNh
C5EcPcH/UEWMetg160ov8IHdfA5rZrblGVX3q61v/o3I2NBQfoBgofUPVbH5nL1u
HKEHPfacgMs0kwEBh4Qy2cZNzul0aZictq3AqYEklQhrB9XmiDC+vRzQN5qsZofZ
CXzLUK2uucXrAHtrAGqKDsxVdz4XA+6f157xIwT0vt1EfHDkzDkkpnX5KUNrYZV5
D2aDSfMJz0ULjsphSbnLkEd/79GkOMD1YL3UUYwcoNvPcIngz8tNuTUwpsNt1Xd6
9mowqbKDm24StUT3fj2slBwYkDphAoRzfDiW/01zdU1scM5mo+IOnz9HWfRj72xQ
ssK6LO42tvmrUvx9tMpgZG50WT+aiQVPjBArPsMKEdql+nh6WX1U8towE4cj46V5
6f6evZ4JmYZhepsKSixD503EpDBm4Spn/irLaG/m+kycL7/xNIDreRKBSdFpyqIQ
E8NsCkyT7ykn4L1iDD7eQsy5e8SzyW6f8nM7V8XjuEmz9aVckEGxIJY6yJKrpA+W
7YBqGywFGfswN8Q2VytliaNNQ7gPVVUUIoqX6pcBtEMSufeIXbXuiVCQKh5TJ1nB
jRJJ3OfUCDdBPakYmTTEPdI6lBvaaT23cZt/5Ew8r04QMWoBUJwy4G/7XSAcVQHf
Awj+OAMTJjWCFL4EwWDyoVPo31iOWGSM1wSPzjOO+d/McXD88eSv7FzFg/PopBM3
CXAHsfmBWDe5mBc+EAbYN/JeBQAJywOqr5PU090koO9gmdQBM55rtiDVKtX5Tg+m
uvBPIYvwUd6A5kselAywBtHIrTfLCQt1Go8VoumYEWtcLhF8rK0mZeoi8Q20Fpc6
wWKXbvJ3hk0zpQ3HqlW7usLxlTGlpjO2g2bz1JTrIqgglBjpzEaOXXc1raADa9Tm
ZlTw9gTUkgayGFzdbVeEYvj3O0oNMMaQrsWlbvFqYJFdIC5p7zydbLSWF5D+6RDQ
SFcLuLkeTHdyUUoy9jYO0W+0u7jmuDpu0Km2epH50eUlAhRlQ7QW4ys26myduGMo
+6ZwPKLzLcppv/uPVzbe4RTsC/jabvNQ2xOX2Ph/K3VSRLlF9OEFhFTyU3zTqn+D
gSIkweZUJJJ0LPIN7hD1k1AOE0HBaXYFwIbtoZrvEUhMtZWEpHj1QTuBl0/RplY3
5zo5d0sjdg942X/MZcuYA4Vp84giqg8mdVQ7RqidQPmHGiUSkhqPFEHeNFeUJIDI
5fsMhTYU+X+m8SqPru6G2oykhE+hCaaCke5/NfAvGsh4ckXyWdOVE0O1N+TC46pA
13FpZdzrBRDbzDrx7x0cYfL/yrzwf0DBqjhjiC+9nPhPubk5PN9/ufhFFbcw7rB8
honpA465YHULKFFjhD9Kv/dqIf4fJbOlcZBQDN2ORa/0WpcXjt3fDSTQzYdajH3o
Wj2GPvcBWwhLRmD7uuReEfa36x2LFIF7jIrvHaJYVb8cPvpQrcScNqpl4Cit53JE
WUBg/jwq6t7/s2SdvO/veioP8T+kwgEfrYu2Nz1Ba+yK/K0ujEYhoPgIGHLMjSAi
hKOVUM3IcJrxM5zvbeld2kRHxz7zoeOKxba3+BNxHHKE0OUgeLsgyuNbf5deiOBq
oyoQ0Okk0JqGyxL/NOC2+nkdFtFr8r7A5LvrB3+U7DuUjLWCxegzH43M8lnhHlux
SQVRpY/IhS2bC6uWmW6qg5HTz0xLSaawFrmjxAj5gB56nSnYNIIqtnS49X4svQ4k
pbRgr9TDROPxegpVu4pRYw5Ezq4dJMaIanPw9peo8i6u36cU8m+SQv7f+u/QSda3
lu7MIa50sNdOmii6wsiNkp3RO65IUYEmj16oENMyFzvjxWQEpGl1MsBE7gNPHTdc
myunpfH7BXSLF3kv6d7jJjQbG01/eLZMoFRC7S7E8qnnMH2YYVv9d2pGqLkTrtg0
t/5NaHL/6Qlnc0SN76LH61Ts/w5ay0CmiqU/dtYFJhuMqNWuCZhOvVdU17py8YOO
VZRKGpd4IM2nruh9s57zL3xe/nwmiF7BJqwaVE6woxB02QdNV0qQqjVPp2Tgrqb9
nFT1Z85zc1UNfX6XvKbqd8KQ80ogLn33z16QgM+kuEjXgkWeRN7rUp5jldsg+kX3
mxBZlXN4a50IWQ8PIk58DUods1d/8PBYJ9l0fkFLc7+eyU/5M3R5qRRrFmy1m9a8
+EVNmmdH6nwRc3Yk64wh4D+CtYpyXH40/nRsMvq7EfvPNaWRZlsFue9jQw5/2UEJ
CZ6fSYUdCXPUExdOODVtWy3cj2wg+Wong9qAmk1yKIZ4crguMOoKK7mhJM2UzF5M
oew6B2a3ho/ahF6Cx9IJeAfBBLo9qibcijbwu96FJ3h58EobsB2yxe0iX0CtfOTZ
RCsBCzEXcbw3+ZZQxWpPK7z08HnOWsf32St7EYSs4uzKc8vcZbSPdXrS1bKnEZQ1
NMn7+74H7vsVdwiDupe8CyusiZnYiz5l2sYFULOchHnf69tE4WB+Jxws3xhufL/L
DjDews9/WV6dHN8hxw6991qCrONJQX7H5TBqLWhUnUhyCaAd3AFEOSH3vao5crdk
8Zxs5R2Amz6C4b/SBhh2dXbWt4Z510KSIf4XwSBkRRXVeY3cwxgLn4GsJMQhTlq8
rc9sAUpBxFRvTddJpLNRHxoGW7DVz/i8m3OhlG7VtaL3RYkl/+Lj9M95lnGzSbZ+
9TSsIhAnHkpeT7qMrmg/IdtqjGz2d/Q+g/B7faR0HXda1CUlxmk91qcyZB+PsKR3
OupF7Lxq1MUM6A5CZ33KLUEssQp6MvcqLe1aqgYCI04ngmfnnGZHCDFCKwxZCPZ8
X2U8Y6omu4kzmjgL+sGcJQhm49IOMO18qFzDja+v7bDjjRyLz2kETxuuwsJSixXB
Z7L1pTVtNb5aZrLLWY/5El8qQIyM0eL1wS90sJ11C6cHszNv7y0zY02/GAEL2bBj
2mBhHqRpH8t02Rev60CjnX0Jf2fWY27qnEs4RfMWWde3f7sNfomNzEQ9Sc3VnPdA
ES/cFMSnUQil3gCWPExRMpUNjLbqPf8agfQED5UpxUZIUA9L3ZDcpb6NO1T4x/jY
TXZ/OWchPD/3p+ZvWYe18nkZgVIDQonIQDCJ2ID0NgAeslyFY0QdMQ4wp4eBf+Xp
dEsTBkYPsYn9ysUdu4/WxaSBgqOr4FuLFWp2F+6RpIZcpwfEg6pJFoPqIgyX/8kr
r6zPk+BtsfrqBQ/ABj+9ivRIDbqFD3wwpRXwOAXddqTeoxA0PbB2v26LZGu1Uc+R
e/8Nms4OReCx2KelyJxYtk2DYJYngCXsNJRh9dOgJwwIWuIGwM18htKS+GaDKSBx
8pFpJyr/PZnSG/AvdcYftdaaFx1bNS1GI68AUkROZ+Lu4rYWEzxz/OD2hRjMPlFP
jnp09xeFDzyzORQoiFh/9a3v/+TOk9GxMPrrApiwjyNlrA55qvxEc3r9mUrNMIC9
gZX3CmjLujumw8Ov5W8JxA1xLA+SwloU/eCOAT9bm98ZpMFHr0MSy9XaidQ5ER2i
xCVuDSiC9LA+AjwnZY43mBq3v1tS7tkDr0lQ5QdLiwc/RK5bKpCwzIw4egl1XkZ8
RH4ukTJCXJ23zKL9A6PyObhAvPoRW9VMQu/qXS/EgDMpddJB7pEYwCHizou3MkEf
d13/f+eWkZEXOLWU3D5AUyHVGqKsDsfxE4zieycK/wmwH4eOopbCPjXc6DIXbVSP
tZWkhJ85MGdUCYpN8tDzBQejP8FSuuyBNz5NSPtXuPBu92F1Hhlh3gni5JkIUFiq
CbKXNbIDl9DaqxpwUgdT9FZ1XASCH1dIuS9U1MKJgzGHckoVNN2VJo1er5wqa1tP
kFFyQlFx4LQcga1B1gCrY9F54qdG+DCKUIjfjeK4D07jQkVPTREtZlZm1Xz7V+gV
4J2kp9J+iRXAJuhHISPaHwOtAq+Y/+OhOy2tfOqrIBzr56J9weGZDVDfYPEhlTuK
qCeU+22Vany04l8Fa7Ldf9KZNECHwmNUx4rNTbobUe3xisvF/3uGaEi7F4FbaIpN
xfFnVqY/9WJhPiqhQ7BrYVu2TaVnTfRQDGuPIAGiFDVebn82TqR/CEFUSwTZPPd+
lK5/v58ZWwSRJugu8Hr2VF8hEAUxd4lTBOrzfD2HENVqJNNpmOlH+6NsV2c6OJzT
jdrkgTcCzqKP1TknvK6Ydhh2P3IZkXxAyPTXs/czVZueFN2khIPRYLAMf2Q2SM49
16BDhhMipICsncVuQ2PM5d6oUGW0z8OQHaEYA0gRs7+Ze8YtYmFRm4CXzYsFWHVl
Wv8A8RAmzh5Y1ECjFWCdCeiwC8zvsLpeu7hDL9oHbpKNtoP09lW8ZZF84kWpakh4
x6rIU8rRTbGtKHnLeHpfw/6g4yvvmQ/PfM834y/wAwRieOg3INNS4ZR55lns8eCa
0G6ccgHUe4sPPfjx7JvWQpImGxdY3bZ/SfSFKuU5aKPgyJs1IEZ1+ajd6ZQBanhV
CDNNCRcYy+igiLc4BvD+mZsyWwHq/l0vzs+98gxZ8/qzrSKUTMkk3aDkMP8ZsZa6
nRJSYUjSt5nnO2KGB8O25sZg1SAvRQwmT+/ycnqMjBJ7jHq6ra3oKVsCln4RIzCe
AEumG//Gkc/5a4XFKgNuDuPQprLr60FJOzGnTPODziSndz+slrRi0lIhCiv70EoT
gdzP53A8flZ57PIuJrE6LZnGt6MgLpia0z2r5IS8YK1gyiVh6sQgg4KlEYrrEBwm
m63haVZIhbt/IBlQEhx84hFA3XMtt/ak0C6O9/Wv7XYp+AQpFQOhOoMqxpfur9yD
H3iWWdTBU/fRbLs8CIM3dEdIOue31bPXdMsRzXViKzzn9nuWgJy3EpR656+Fo7nS
N2D+1kYUb3nCH5dxlHb/eNwwnmDm6kJAOJINbKhiG84P9p+9+zQCRQGvnJr0BvMo
kOEP9b89+DTunRqzMH567NE3D3gI/Gr0LWJ37QNU0hI87ZYnr8RKNEuabA5MDjWd
DZu+RQik6g5CHYdvoShbcMmyDKBW3bE8mNKzr8Z8ZtKFET2k98POj6JetOuna8jQ
KFP47LFa6KFcSugY9xi/TQfWllDX37qQmmcDgXI8Zd5GxD4A0ca/jSlYLjiXYJSO
bea/J3g68iaaME5xaizfaG2pOz6+9tUxSjiy5wtb/PIQgrK+Lpg0fe6RyqIErM86
gzdtPqAYdwa8VZAdu3kLeLVn9+lHAlfoUYsTN5J9JeKIjZiIFyA0K1ZJUGarBmrb
9Wz9Myi347z1/zdBN/6D8AmBjPDhQI26M3ai7DonjJQamdjYW4nrfJuKiXUlwdme
C997IE77HNRnx1f0cLDvJ0bLCSbvqsCtgSjv0F2LGVIw4ArxfAYnkJiKNN73bWxm
v4H/CDFVJ9cSNPXoQu23iFcZJ+UZKeRGM71Zk2MMA2/SMZo8tsO27P1QykS50Sf3
VSHPxchPvo9m18x4+Z4KR8AIwvvpMdkOSauljKMH1pdBpq3tzdHVsOaMjCaHCvth
oflpmZpNb1IAEoTLh80o6JYqYF+M77dAUanysb5iimMbP/L/P1o0Fmv65xIFxct6
Z0BDpiqgjCDTqoFmx7rAhrGiu43+iCrDMgn+HNVytn5omlGK+ByTBD1OF8Bqh56v
LDIA0LiWUIsw7+z6GntsNb1YCaE98i2qIO8Vdo6entGY9UTR45cPBhzxwYlDKdVP
KTTd30bOLkNDX3bmgUJGb0Q8/UvRZ/fc9/2ndJgEig8RdK3v2oV26lzfPr2qcDzg
MEdJnVXELI1hBwJCg861b8Kd/79czUw07yNQIW9fKvKSbKtuimXc0m1cbNH4LSsu
GuiLrjcpAPCrr1QNeYIEWgsYc1Us4dyPYB0XvVHmi++t+nNM2yNuTSNSodQZ2QOD
zR/dqqqNtpW6R8yYl2z2n5pLRIUo0t7Mdscu4kGlboPVUKzbxr7EDZ+BVkDPE7cj
mdD81E4DB31sF+4nhVj9dWtokxhjZJfDK9YYFoVy8Y830Sh/ku6yU5Q2K5X7fwEO
gsG4uEeV3EbZXyrFx3ilUsYFH3oBbh6EsUgEsYOmTpD5whCDj0+uLChooOGEAOrb
eZtAxiwmeIbnbOsttNV+BMejST6p9TAadsy6nTmA/5k0m0JaM+KcQgIQ+YIw9HKl
YH+ek9rOcsqGNk+2WYoEx9PZ1cmBIVm0vrtDI94ChPdfnJxNyzqzfHtj3WuC/odz
RznbRyWzPB+xHjEYeDTyZuJgJ9bTZCWIsLkz0YlHpTkg70j0rCxkrBREMMCE9mhK
w7SUAOm5+uyVJ2g5eI4XICTzQ4CdEZ1AQHPVf+Z2BwdQFyumRysuyw5jESHJIMIb
SsjMhZOWpm8LkXgBmOuY+KB0V5kQF7CIw/PZXKsLuf6pqgQyW/LdY62BX2XS9Yv8
xQ7fuvC8deQLAMWbyBjXMYbItqloWbyonLWEMBmiVPiW29CvtwRWO4lNn/czbSN+
W/x9JzAXfheugszsaMN2seZ7czEHPZtQYWv/uYk/hptZkuDipl7lfrSnRycGYC53
z/bT3CwjQG3PwjiK1fNjVjOYjSG6x7qVYC3Mz9J7lEOqUcPsjjRwzE7KGj4Ya4Wl
kRosGjioZdsIVTU5b5tvVjtexzSLZDMISgTJKx4I8qySPQwvxwxZ+bOs+OeiCSG9
ii4u6xD/L06Ej2Nr+uaqTYVubqWyFw+clCjVRItvv3YU8tZF6sxopfnm5khUAcCO
UdWwxUSwkzhcwqH7jg07TxE4nYaOC5zwdN7PjxETIYgXuabiOVj3hg3L5G+vPP4c
xcAE7VZ4eQynrf6XfYLCatCTer8kArtPViZNjTq/UnNvYHqj2ewlfgLYuB7oJSAf
S565nP5VgupwOeTtqvLVeNzg0P4SdLcKnyhQhK0NBuknGWNuyBoj93wPRoeD6xAN
d42Ikbo93KqmjzozY2MRTkQZugz2jY7vNvWp80aX0/VOWo9OggqodEOSuO/ec2tz
zLLNgoCUYkQ9WZXez2EPrYqfqGkSSAhGolKoBGKesjXSQI3IiQIsoT3OaKuywLWd
87DDvfZkwtWIqVxDTpN7EKR4uu3D9yz9lrbJSKKxhN0LmpyEwG9Wy3DDJrunEdlA
JDsO9FV0gTIemfjdKY5aqor/Gi+zfR0AIHXdtj4PiDRoJ0rWK6NNydE8KyM9h3CD
0vUoEZUMb7RaG+JHBj89K21n2vHpvijYzXET8WBQNP6rQeCNlvADliYo4Jodk8fV
o3Cw5vYU2nngtCKIsIgBxUVIKK20jDPKH+Kj2mNp11R9H1meyJeDY+exST94RMCY
oU5jivGls+ApN+j8iv8qnpjuACHgKIIznzH7o/SYnaO6OsurN4fBqRtMgTyEVSQM
rpIrVW6HL63gPs6hk2ZRMAVOhfsPW2bOYjVx8GUtEqzLi4N0Fj7ObBmqdUufO850
wg5lNvnnHQr5bFSFxq9NPra2sMPj+cZBbztdg+XMKWf878mO3ktDdaM68S/SJ6yR
Bd+A+YRLyCl/sXVBtswOpGxraLX7gH12eisQxSWkI8cRALjfQmIT339yJTnSBiqb
UaW4ue5OKKsQze5EUIxKP5KtYzWiTrjAaoytdtMhHkPcPSFuNi9CKaS1dvGKAxws
CcKf7kvmZLQBVBo0QX/0nxDTnKyhiqHHSUffNaEXdvHfEBBppaaNHv1elasumyoi
eUYVT8wpR7yq98AWXe5LHs4gIMcbbWklPpHSh/gzndPn1Ecylcp8pE0AQzN834TZ
KLz/G7PS3ngUeWMLbtuEdVV2HK0vGdAEYxzT5PIO7MAxqT32DfODBCW3Wa3Llj+M
finAWiw6YOLQcs0kBopQfkBVP3jsXaQ1AGIJBwYcQnAF5UehdWI3vl6kBeYVyKWv
Ar4dqo9N4ihQ7XyPQrSdzyKt+O8ilrR+zsQVw6w72BZUabmxYoTo/llBWzyuS5d4
vej/Mc9XdZu09QGubp22dxc/+tZeg3GdId7Fl97sQt2wygxpUX/j8IlwiCYnAboI
s5EBVycPwQ62TsNEMebNRcsPxyOwaIiFcfJm677CYyDTHDM5hHsYcg9Ge5Nxm8f+
HPLbcG2mQN5hc5cybSH/Anf91jixd6NFaA6OjqJsemY0l+4X9F+ppywgq/Cm7jGM
hTTtMxqOJscDQkVRcxPfkNVRbVT3bTdITebGLulU5RWcu4u8DhgqQq2Of5zsicGq
nr09u2uf17BbmgdJc1fr6i/vidFli9bUkmgNKxVo60pTEwjhA681XTsO2fK1oHgh
i6F2bg8Ak2IMhmqGVGW9ZJPXuRDDRon/1JOfBWry39icUa7JSopvKPVZ/8uAn7kx
aIpbwtBZC/U02z0Y+BpGPTxH21v/9a56C84qFBqF8F82ALWqwo9PWbtBDGthQWSx
4K+wY1dsFTfVV54TnwfJlv7OpMSiOGdHBzdzO0XYT0SU9rb+3aUXpTNHo4UIGKb1
T9FRIiZKeYiwD1XU9a56nMUctAzSH9yzwM9LERGBdeRIjWgE+G7yNJ7J8BwBuvrd
31UPlQnowrzzvBsPmZCx6niDQ7Y0cc54PmHOfxU+PmoH8MbiOgS013ABc69lp2du
OuKtm3bC5SU9Mx0WWwN70OizKcJ7zsPSbnnaKMaxCoUu6ngmTQRTthloVTlXuG64
Gc8viUb9oD/CH2H7sbZB8QhQpBqQHZZz6zDw4NI/EhRPv8+4LhbBoBo0gkAtcIZl
+aOYZkoRjd3/R3tUrOhzpj36cGf0gSJ8lC9jmjoDNSzQc0rZxgfoN/qYhOth7yxD
wMmYXYKaohoOYSJarvhtPdHW9yQW2bnEE+skjj4yC9w3NEcFUnYRhWzQtvXN50dD
M7l8ktWvHhcOZtU5NxANHOLgr/2YacfVJucJyQ3UsZTpHk4sXatjlJlM/tiZWIbs
Y9TpLJGMTm4LZeQ+HcD8M4tv7iBcrNlZPvN2nGlgjVEbSbfB7a82fpecfwdeOGt+
fEEgIpsa1O28hOgKA2Bq36sp5+Cy7+sQaqcD+1bz+jkU68whsKmFdvMnCuezkvZk
dQ2BZdv2L0uzMpVXMqJhFR+Q/TyoWXySnIJ8diGvTm4plCHmSNE1lyCl/Yf+qncT
FZKIBgt+C//fHFPzIOIIX/leZ2mGpsMBamjFs4VOpCulVi3eYbN2G+eOMZDKYxcF
2PDHpZpQzwwQAL5dDdwazMk9lvRnuy+KJQolqoFVOsOtdiN8tR79+SJroUk5uJsM
9PBMBuSJOsZ5UObv8Uvbf9pa+6PGgp5BaCLbeBuHnfe+TjmOLtb/wG5ih+iEiAZj
7oc3B/Fsl08E2/wzcsbuNxGhxeFHoyVDEcw4rBYyT14s9npD4tLLZOT94LoG5mA8
q67F+gs3wJiV+QajLBuZMoSFr9wziQTdOpR2Sgs/Bpc0nqo/ME3p+lE6dRIpsW+9
QtdRavxPIqcB2+rG4AABEtbB0WkhsQvUP04qXnQjhz5eb6+f/Rnc2IrXv7I6rtME
gVfassYU8EmSl4i22SNzha2tp2U4QSEN0pywS9gmVsqvtdQcnI/zKRHxw489deJp
/2qvp532j/iVg7E8jNqdbTYXjveXQgP1odgPUszPL8A73Tq0KWNZNtQGIiWIoIXj
8fydezB96mctCgLXn8QOXdKO9pMrrE85c5dVxIfsJ4709l0Svk4wgwXGqHJM0Isd
/5R36U7WWMyi/41MF0JDigxAUwuJg9DRwbnudm0akikxjydeKYCfHAMU2bCwGuAf
oXs6pIAk7ItUEGizTWP3rBO3hXZ4Y7eyrWFWG4hnPUqPRF77bRQy1IdOzDU7Ci2r
HY9lx8xavj9Tpm0yCTOXEK5pquDYKMSOCeaKbE8fvypo5wJ5Eto1ZIm+pBt6DVmf
qzNtDYqD7L/1e3vyV2xMLXL6uWuzYXV2bSozpwlxiOpgVFOGbbqA0q/fnEG/v14u
Xg37PEnZKNFQGK/VDYsJDuuDJcvCXNs1+Nx8rjEq9V8wqDrxjuf16LYsGcjEF9+/
lnlsasNAtdVMIlBMqs60Ud/3e4WbZtb0fxH1HX0EUt88mEQldKlA22iQchf/90uG
WlOhrqUxs0m/Dw9QnV/cIrQiLcGuyGx1AKdYS513WLOoq28eU6eAFd7SrdMhHmCW
B1BWQkuHw4y4CcQ1hWCSqb7fEWSgwREFWB+I2BJmXJW91REl3EpDjHZQHwhqsNep
72+cubZzVdIH7tIVqd2URD8WNRRREj+UOYbdn/zCF3fwZpu50+GuNLccuaAJLQsx
5wkX1NrljdwYo/lFEA9WRa5TJlpdT+nciETCwQEsL8so/1c7dQ3sjGbpBIUUOx4K
XoG38dIAEDSNfFcLZcgGsggcp2caeyYOZBpYu/MUZAkblUM7618rv3ZnA0qrpLKo
PIRcGCbh8V4rHcQPibTd7XPjKJs9hBO+ZFBtk9/nuwd/cUffZJJBQDrD/GDyreUS
6+j2MGryMai72Il0sNdSCw7Mu0efL5t6woEjNK9gnC5vfEZRXTpFVkhNbo9sqyNF
Z0prANIKQRRC2DlGvu4YzjNCLwrSMg87RhkCLW0Le0J7+V2MZxmaLkgrJWauILnm
BXE3VEhuOF95PsxFP/uY8uL7LNe6v651QHwIgGTf0WN0rS8gYeE9LWILYllzhXtL
08EoVPk3PB1ibxm5hA3uj+BsHaop72ugwvOnpDdYP3ahOExP5iNHD/nnDXFgto90
YtXNopEkEx02Tn4kG2rvpiK5hl4k86ZJ6VUdS8gTO7v+90jdfyKZwrNkOubQSUGx
oJpegT7bQ3wMPDmklY6fqu1mcZePFYtb+9UqHCSyGFzqyLYgLNnaWjnDFo/3rFXU
DvbRp8WkOViH19Q2ob8I6VOYKqn9V0YrzMePkMfT57wulmlNBYFNsqVoFY9xVrAP
lfvjcJqYIqqrLdhhWsP9oCJPcnGpUfNk9umRQlFSyLYgySQ5RrkO6vw1r34U7oie
LvzFYrxWdyrLSL6lXIfszx96vrjm1dWYzs2M1qc+DEpwfHFk7xABUkECY9YfAZU9
2LJzx229SY+ph24+2UE6Mhh/egQNP6bxAy+ZbzRc2/aQ88xjGMRepeOG9UX2SPd8
lz8fllbZdZvo3aG6vq2+1ACUjw6G5MbkdfXtmfqTAc2102CQY66Kyxamb3w4ruh7
GNYVXg0s0U1gFT73nh626l9ogR/e6s4g7cIn32NQqMqJ+2MCXEpRJlJH9yV0I8b6
N0M0jPfjxLAvADJvoLR0G0pNurFubfbz0tlB3IWmPwSguEcFASXWV61MQMpkNplU
8ncHWfaCJkI8tS8KJva3wp81TkUSKFv5QZ0MFNSOAzH86gOVV0VX4NU227jAwU0j
gfIglNYxkWmD3yHKDgUP1ap/W4pzEQTAIcvU3RcyeY6r3icaLpib3jjGGzbfKxWf
rK/V/54eVdvCsAgiFE1q2zmiQv9r+DM5JDrdJGbxXPKBErD+XXwmI70stSyPvJya
WFGSz1k32wuiubNHCJ6lv60tgU5QLpqJu8w5WsSne92T0qx0hIyWPYZJlk4uR5ri
Kc8LkFKGUmHbtxzSWohTo8N9AcOHW5g69VW9lQ5Jx084ln0bvhtPJgZB2oEy47wX
4ejJthD1jwUPIpGQQsNopstoJwTAoHlkJE5sP2lW6ZzJ3pxu0rCX47WYiUeJVRSB
Xq0y+xcMel+0NWsUcTUlthW7dWkcvN1pQwh/s9KL7ds/msI5Rr+d0Gg5CJI0FDqm
oezVX3eS+0UtWZ3/zQMkRmIYk6ZAyWozMalH+wBPQJB6QiiZAT1BoAr02Obtjtr/
eWUa32jC4N2Nz3tb0OJzSWqj3I+DgOqwKd6Kqn7wi1f0p7TLGocaBp5i5AiFQsQa
YLFXoYe4K5l4mqdwqTUObOiq9MIAEIZlhwLiAJkq4iVt82hlZv2oRylTeUK83iW6
++4FtzBrTYO47uQ+/nXiTzutIxTlg2zEeBtN601fnh+9qHpDLxfSdsXXh8W2nH3L
l615bKUNnj0n9A+SL1V98OJ4suBesuQRA8nzI6rde860fBnoAkH7/MqIGdh+Xpw/
wVxHGtVGAf6rXF2m0DKW048jpQZGV8Sj6g2UXZCKiediqNdHEJe7l/rY3uJc+nsq
/thbuZqnbDebnbLibZUQaBnR2ZUILolXr4efvfJP1m2e9eMF3ihlcKSxarPtsro5
2bWaquqNifieP1kasaZPp9D72Ovn7OppHgs4/2insqTx8xUc6Hwt0nAuCHIdxGUC
1zMRD7kPs3/EPqip2vCHwY0lEap6raPlSq2gXSDTxYzKlFd76nh+jr5x+sraOR2r
2F7B1xTr2jnrhfSjVsc/sIUDAuEcp64sOsM9VamKStCFR0LQ0KNHM/9FeNU0ol3Q
drM3WxEhQUgSwdchUbxlTpNNp9cq9fWwD9wzvcrnC1ByRsZ/pkh6FFisT2jvjc1u
Ft4o5nCtTwTBlSwYaKEGio39HXlPS5D+IqeQ5CG7pw+xjlqJD6qYwCh6yefpUN6i
f3p59IL8jgKVa2V98eNHjz9T48JD3S9SLrBTCl/4Yr0CpGET6AQUb2Wfswxn1Uhf
BwFLkiLMX2imiApUVNykJfkvagFUdBq7o9xKgyoX2iGn1qd3+mlSzNOj/LN2gHmi
g010cMXSeWEUi17FPrFAhma/yz4n55iKCcFt9LYDVy7CbQVOcE0YuGslL2ES3ivu
Qt5wYNSVb6D8Du3CrYG1xPFK03l4WvJEOTFnTS+CTfoAakFK15pJCczzePasJvSZ
0ocPWUbRcqWckAROxcprnzaa7WAZ6itja9u+jGPf16pQ93BuONQbi3TtRvuqqHLm
nGMwFQXx2gBDRUTQrW8jun1cbT9co0lgEkP40dJxFEkYweSnnbN0CE/+uwX3bkCF
o00678Sl6R6P/DA7p74zusYpW2jhoigcQ8TDmymfvBH1DRLtpy9ZAy8e+DWb1TIq
eeiEGKjPnQb1paeRD3mmmZQ9cedqkXXFVWHhrl83PmSHtAdUIM7fhDonuBxmc63q
vfmW5+X2rkysfkMgrL+B89N0Zz/40r0sPXqigZRaWEVa4DdgWfCNvJigp3ewJsEu
koyEWkTRG/+E0WTHIgylE61UZ3kGbGY9B+P5MbzRM/9tHZwcsn3/vezacO+8RYbx
cMlJ9/boDhrKrHeITGkF7MfwrJRRhwMotUPISzNSSz08SbvnoVTWY4lli6QmQzxb
OWfProVyylLFmTOT5yszY4Z7hGPnTlY0ADnBGeYSLS7TYjPNgYmey1lW/1Qy3ilr
dPjfvlB/Ek21rtYloecFldT96b4hYAwLDO5P6bbZF+kDjCr/I0TNYpcCjGtX2zSZ
TdB3HgZkFK46/hOCNF1fxOYngTfvqOJoe7OqJOIHE4RrXQMfKWZmLrI8cpC3EdU3
SNp9Z3zTpFgXhyac8vfhUQ0xblgyWiop2+YvDGBGbzOg45hkn882UlLzD2Xy/QTR
heXBAp08j8wz6h+dVvFRM0IWUh+aB2UVRTtdIwL5jL+oCdS+e0HKBelmNACnKchO
uS/SFM9nwhu8Nci1bGAFHTQuK1zKXhpVFMFGlRT1LtOLBN/hJ82hiOcLmRBISECg
pLiQt3xNVUGSag7Pl90TTvcL5iUcIX55Kk+VBQ+fNnJzbX2QiIYPIcJ0cdY+/f+A
7rUaisaBsY6f9xTMLZLjFMFOIUHWzqBbCgZwpe5GHkkY9UcZWvxX7FViNcwcTkWV
sb+eBBFUFyaNbObL7E4AaC+5y+tkKIOFI0qfd8SYEEmls6CTwBz2YP1PrELdsJPL
xFv5G2csMMQ2bbsYxJYmm2maVir7UXKuhvl98njNMTrraHo/OiTB7hA9MmdX1Lxg
XfaWO3lkTsrso2rlCoAgFjrzDjIx4dxfj46JJiMGhTNLGNh+k22eunHqy5yvDEH1
uLevx+LkGJ+9PqFBDXkrISyoeVdjZAaKqPNG6CHkMsdJUnciU6CnRFXUkkGms2su
ovt0wNGpEFAqEPs8p1INYkxgKqWwWs++CHUXsjKZ8TW7aYFjgejuFtADo0o8c/NS
rpqkWkWYY8TDMjfm54s7I8IqqSJvcyzu1mbnWpohM0NDeNrD2QGQJ7bAGpg9OzDD
oav9j4XqMVrR5CsdX3qQcpqEjN3IW9k+l+FXZgMcdEsolBTqe5iyOpMbj5olyBRT
3GwIWoYrPvJfTDCZqv0E9XyV/y7YKjer0DckQoy6LXjlwj2pk9qSEffS0BYtFwa2
Llp1vCSMLDvRQdf0qwxnGOQF1lAkXRQO0+IC2MSX5VDwPnJxz24Iml4357LBw2HB
LX2d2r9YPk3JeLAvweFP7yFJP1vKUR2TMxlgFv1FZ2zlneBZpT2Z1K0sOwAAk1Qx
+WaSTSxCs44fWuXxCXtO5EBYBAkA6uK16C0t+c2LlPPKjfnP3+/2lX2OKKus3oLC
im5ag7hWwD9HuTWqhYKBotrTDr6IzNZu7WLzee8i+9THQsDHAfejloccfDdD0y1K
h8B4JCBsSEyg49af81OQ2a0UOFJ011Mjzk219DnQxxVC9Ej0E9Ejjb88DW/w/2Ce
aT3hOPhBl3rDOnePjcu65nPM1Nj7XRP0j2co6aN07r98ygQSNnzCm05VYKPu/m30
F0O1Q1fDgehxFD33TID9zXwL6CEtGATAoZfLNQ9Xvdz7KZXhLRYluZFFRjCR7wg2
p/diBHYhpkXuQOjRxUBJ7GcPPIU2ikzx8t+yJYs6aEgSzbOGH6Jl1CGd/yfF61rM
TWkrFzDfNTxxnmSZHvFE6UtXyteePx1O2HNLzUNEAvLfaLmu6XbCROGmlonnAlY6
DOvLx5G0YZYVZX3VevJS6nl15Km8LTWVpkEmGDcT0fTPPxeSIz6jNV7MJLaiAXmt
EOvTg5NV8PA10pKQlHoCY+YCCmhBBYUbmkNox7hSSAPcEMue8PfipRtJVcc0SKdk
kRv0sLG6N+Z4m3b2F/7+rLk6ky1pOZXx87PljWiIZfDzkK0DUP5OpSTjsTaYTnYd
sVHLI6DRR45R88twqjc8Fcxkk6L2wCs+Pbnw0VnuC6VWROYFTNPiHAxR2QZT+D1m
YdXtU/yFCVdKyMxlVMqKiK7iO1Z7Dd2F9Pbo3DZtQ4Jkxx8WEgkCyRf29/3msQdo
z8VSUS20UDfyhAVNUsqIhBzYb+ztCt7qRXYkHHA+SjRxU8xj+Wl8poR+8e1aZZ+U
pIuFYg7MN3JkbDzVgAIiMltQda/fIy5eG7QlSEWIB6nkSjAQt5tj9HwxVelJ+ZPr
jN0ToW9Xzey2Clg0qNxJ81rwx7u1zTxcJK3PNHF1G1PwmKKj1fVaqD9qnSuEXKwn
26KnN01Za8fYjY4G5NF99CPe9dTR/2x/0WWCQiCjMP5aDtGriUEiHXFiN92UZqj6
ZEgckLMElxTE6jLwJNxxgKETOq3Q8GIp7WTSo/b4+AYloaygJhvvCjtY/UqTrXxG
SCML8C4A+8qbmF1ZbpIsD4RzYQb+SqBQK/T54r0W0MK/s3ep+W/IIC8vUVcu6bVP
XnARbQ6At2fpZt3q3xptMCWuo+reWb5OI3GkFTIq0cqYJPBUX1u1O5+moyXc0ZaK
WuNkeVJ+95/keqjeoAHk0f9halWe2dS9NCILe+MwyvYZVAKTLr6M5ImM2l2MINPM
XUldoD3XFZlIPwhAT3nZd5MST5a7pP2nhIyiMw/eqk7Uo26bVfCiJqDd7SRBgF9P
p7Fbgv3bWoiM1zVPiJ1IvUzZMQhuKXBueYLg7phY4iT85nDGCHsyhgE6vctJM8dS
uyMOTqHVZEf6M1upsS3+8a7CraEBm1x42K4PvMXQQ5lYm8eVH0N1U3mg7YaCX2Lx
tfekZJUWWgUDQXlgekbW1qd7R4veGA4A+8Tyut2w4mjzUt3YNMMX++I3nbpACrLF
QRiyeM9I2luyqAGAZn9C9mTfzlRln7uy2UI5zCKA/cUjtJlHPIDwdP+LBNw4uQaP
XFDpgNCbI6+GcKBSh6i1ltL3pDiEHRtT4Dw8jDRuWN1+gtfo6iG8I9IQHko8dK1v
ihMiV09mdY0PsfYKvr9q8QaL/1JyNMu5IoZHI7PBzCvOQk6SVIyhcq/zjfyrxVZm
zBzBipYZIfF6v5OerywFH/9mze1FOaIrRpR4FGj6BUQ/rL/ZdQsQYzCWXc2qlUnp
puP65WPVfdlnyQIa07VO7eD7kZz0bBFswhZwTf62RznKOg600AiERLmM/KZwSrR+
z4aNl1CXexkyz6NkjTj6jtXKTywHL/lF/uLFPyphpSCasFfCYG1I/qwXznrfpsCD
QMwCSppLUrtiiDfsNSdZrr08NaIOQQOxK4sNZV0SXY1y86dkT0VWnZMV8fpIb68N
XDt2ZIqQOUv8FM08f1vCVvuMXxGQwtbqCaE4ruprogZpmzCd15tmnWtp+PnWvToH
V6l1diaZA76oC7d0FyYFwLNYGyeFAq+GgyKo3PmeNQUhASBy7uZQWXmSehWRGFhI
OrDfr5XS1sJjSB7tzF8A8aux22BSO1hIy2l3T0i+SGo5PHvhcDzHfm5sGY6xVfsC
qnlplSxAox3iTDz+GSMEEyzof2OOcmG/mXLbVXnzvdgtkVKRwzftXIdi7+g4fVwb
yGHKR99fCNA5kTANnzxhWR+8568kVJjfdFE0KMrzSSdQ3phQynsC/PMjB1QlU50q
RlTxCe/LwTtVrD+YObcovKPdfvafonA8exTElQRYLqkPXdVbvVyzXCM1L+W7Vxlg
ANUPyXotDCcABnoWK8jvCzcpzLj1CJw8YkktQljurm3+AzHvwh6aR6HG7eL11YZR
YwVJ0R5JZlATuQH2BU+5AZmZ2WMxPcG8VxpS1tCfvDj6KRBZAxaNvaUZcY2WAAuj
S5mE+5N+LN7S/Pg4bmPBcEx9iC7qDRYVWnq2QvE8RUGOGIvx3CTTlGkzYbl1sMsy
GDGQlNjCadihzzG6gIp/Ruk2gRX8x8vkyi7j5EyOMUwwdZniaIWozXrGJShDnD1U
Am9ykoZtpkdM57gKjyae8QdByys99znx4nndB1oiFEwURGyRfMal6Xn2n/UuKu46
YibjQUzY2wq9cdE294WIjT3ufE3U6cGR9cNVzs6GLqfKZUvJATQl/Fdh+jGwrMC+
+WSW1RP+lq6nQh92kpX/YWZhNu4hDBNUUqelVePDzUaZdztb9ywGPq2yRCDGJ0Vk
oFWLS967pAYoWJgspWmlnUPH0nJFcSb72mjYS6alrD+rzlCX5WBULA0COIezMLYo
r+Ct5CHG6nzJ2kQcEzm0AHll77mrwx8lmtBFaUebiBuqnHZAoix6MK7W9m33jjN3
vqo690BFBh08HZEio6ZRyVpRWIP1lFGclsct13aOHY7qguQm/AW6ssnTACLQbFiL
npwjiLwOVYD0sR15wBUQ9BC1rG7kFOgLo7iyMc9ytpTz3AuXZq3qCI859FNPtlZN
n6f95xZkmDDQEY0viWi2Xw3SgqKCkiSaiOSE5Ycp46fw7p2YHUMslP6gTy5fdtah
Y0B/zYxscAPpMkhZPA0dojiBGqblUpOtkahmMCKi2/aGGF4Fxu0lAjfKY2G32hWq
PEl/2RFdDcfGY5g8myRdv5UJNKPvWAH5MXq8ciVO9fTExw/+4DA6Wysi3dZl8BBQ
6uFTSCvvAdmFBP5LJZHwynqfA5RIWKhRTyp5RAArnxqmBqFdK9Sf3P6p/kJtzTnp
8osLlyRXm4/os2gXv1QFSnPYkrr/nWzFLfREtGHNbVpjIniSKxJIICIEeAk3LdO+
UZ6AhzMF9OWpTduIIfR00wZre7d+gsBrpLEX9rTedNKdX7j3K7NhucDA80w5XMBE
V2Gl8vhUKDmCrn2y/vyzPhTuvWSpcgXg/P+QGMARfabhAGy8KEk394s+PoeY+Ox+
cPoQqsSWV+06db0LZpmzz7LROc7VOjOaX9jDNvKIPsp+sWxIQcmvAl7pnD5rjqjD
EHy995+PRJQlH6NJlREpA2HHV6tQHITbSHS5ynJE1ZIGFMMDq+KegDXkawLUipbC
bu67dHOFNsZQo6TnF2fNj8pdSR7fXEehVPvxg6XC7911aIDYHCoTeDdgYgeom42s
GfnwPbbIjm3E6gqNU0qHJ//G/acsycdC/xJyHyUoNde5hjulXuuR7Z5mqmXnaKK0
QNwMQEz/WUFIoe6H6XClHpIG2sNbsZ4JxHJaqPd896msi+FcYaxQHBgYbTckiW5R
PiO+1cFMwGAFwA+8Yhtrr/XM1Ma/d2lgIJw2Er7fT07hA+Q3bnd3dq0jomH3T/4E
+jQyxkNQTa3l0yNJNVS9oeJmpBNBBZMyMgS3/CvZ00tqaEFvz5otSe9sGFwPf6Uy
rdG3uuWT+sTJ94YoE9PCX2HIJtEgvZaLbPmQZqVoZg5/8IxInFoJE/i23ko8c2/P
4qQkgS2xmuO5XLdRvtVTKNuZKuqcJbuvCNVqs56nzdzzVb5rDR9OFxeBv/3BdK2b
sB/jeo2hr77RuGTQ71JapLEgwkLc6Tj7hROvfu4K2wUcCf/QZDFlmmGssjLZ1Tkt
wj+4jDdRdMeK29/F0BSnZ9mUlPR5MbH9Juhk8X7BLBFdn9gSxpvfD3gdUiUAhmCg
s4nw4cJ8rDti9FhZNEAJ1/W9jkDIHPvEkDnuWMDV+mZ37i5uBLNGj/D20WUANmAi
bxBJh5wVx1nCRQY3m829+/LniMrU5qTkFzTEVA9A1yRsfqWXy5W+rrQp3jdgYSHQ
tNb8s5XFDXCWE4aT5QNVriORq7Qt+9+7vRaSq2mMNoEbh9VzMKnV7OszPmwF6c8H
VU3+5fU3Z+VObVaBjW+f1ESK3y/t0s0SLIHkkLLKoWmrsHVSi/WqCiAEzWG3Q8pN
Y2SOy5KOdS1JBIK1kf5DkCcGVeiUADvBoMJVkOI0TNnRVUNCBCjaVoENFnRAoBUK
GWAJoPWuRvtZzbWc5+/RqN6QMqoOzzSYh3xuYkrqnsurw3CyyFTpFlg3nlpbqTY+
O7w09QAztSHf0TnSADCnoiH0pff+tdb64zdjClVCzh9M3yly+Z2TSq4I5rOn+xpV
csn3hf5Cyoykp1tmLSeQeUfcX+L47VRhTgqhPqWyMxWg66QbGhb2YgTNyo8hmU+O
2yv7nAUcEjEdIKpJ9S/cSpEe3rPX7CXn4wGIRNfj/6t6WOpGEU08VXx/8Z/QE8MU
C6Qxs/36pgtmBTsHkZEOh0QYrI6ErRzfkM3zTUa5mI1SasOLVrRHXhQjfqje+Cxr
fLKWBsP+mkhgqWfL9sAq4aNHMlnzJ7NQH/+vlLmX6YB2bg+0YwdEGnrZqcIsND4v
d7AOxEiN8axuMKHcFLZxmBLHAKBY3fdlyLsDQI+10+l31J0vShqIyapXX9x7LwLB
QHXfbslczcXpx5SIKcdgLmWoyq+BlrcxBkrgUSfgtV/ADcEt+iWeA6q23CfJEoPC
uL2cPERl7auO0oDaac77zfdgDVmfxc/wpXvLSL3/DeNKTHkrYEdS9IKSrDOiPiEi
mik5cpnr7WU8NAABFEaOtRNuaL0308pdI0KzOngjuntZETeFL7OH1m9a0UIBS/rt
XbrRYAvxF8ySkPo+ipqGQEyZmttu5MUGZC3YJyuFMr0vaKp0uD0I/dVe5wXmvPhw
z26Zq0ym3O42ILY+q/pNectQ2+a8e2c8GbwsatGg+MZJDTsveSGs9oIf8uFYiUDe
avKAVskgS/euAjMPvVOx8fmC+3+oR+wOe80NqR/cMKIB+rANWXQI+wrZhbgApr8e
A+5zzEQmCS1JqADR/8snVjW7XzxpUcMK9Y71Z8WolGJu0HHEYW5AstpOeieXPx4O
NwwzKhQ/QAcAD4K/AL7onBbMrNCR1HOUtTxukEVFjY2TFSSEK7PF+YKaeD0BpovG
F0YB/F5TciHGO1aBhHp3/EwhsT20BgVT8YOT5vA6o0gleuqxFGEbiibhracv1cVD
q8C/X8NCq+UfnIDBKMBV+d8FxaSlTJop74sjRcd0Slts4n00TuzjJav+Q5+D2bUt
CiokXTTCr+oefSw8AIHuDiTaI4Xp90ZZvQoEnz8FAgCuIV92t+KrUE1ybPjckqkA
VTko1Ipl7gAODdGYcdHJJxjwvpq2OBiyEIIBVX1E+eyp9j2cbMelS5ZwjqZpgPUH
lB7dhEw9j2YONBGGOSc8Ob+bSp7mZFMjTT2Tlc/grYlDIDPlgtDS5My9msMUQXYO
mR0xsrbQYoOexJ4A2WhIbSHgerWtAiTFhPwla2DKx+/GO2eAVcz/KV9IWfqFtLI9
hDHs9Q47ZlgDxEf9NitkNkwkGUGLuvlOrWVQK97tPO74xopXFJdQGHjHt/4OK4sY
w1JeWGnKLqiucffxAp/N/YUmdsdtopZA8x13hd4MxKulsvT/qmVQ4LdnQFk/HXjW
IynmjyXOGlCHEszeJ0Qd3xjeIDKuSTapH2XMWTwngvE9hqWnjheL78irvtHfUTcF
FWeaieUS2Jg3gu2CpoUIhogIXw1KLBjSDNqzTevwtZKmHjnyTzGjKobmVYozB5VN
+ZScivLSer9J2GtTSU1dVz7PuFVYpZtQagWSqgUavnnxT67zlIm0E2X8u6mVmKcX
1hKJEKkY4v4JaKEmSRPnJNxuIy2qbUiGBJOmtiIEiJMxFJau/MOS90elQ3BCCHRm
0D9NFEnmKChdVeH5yw0mvb833NiXWwqNb1ZnMYq+bSdVdiPNXxH4XwnJifdiOBVu
0ki0ImO7XKSJXnw4cdIu9CnJtActj7w0sKjrB8qjZQZ5EfXDX1X4kiVNiFi5fEkG
sTxZ1XWow6Je/cmwIb42VgdGSbKj6BUIQOgsbko8Zy8EplOI39q0LAsPJRv0IzgW
J7LeV4FmkQSsyahAwyRP+4thJ9VOfzwcZS8zB0XkCQBqdTpTmymAr3EdUKEAA4Ce
fEYxXGrbQQ+5xZR8H1VlqIXd/e7MnAV54f+K8xAx99NplJwHLpabGHlQNWm+ugLY
4sR6549Q6bQp5WSYt2V06nKt4vQncqrqBezGUgd9qyt5sCfjTg/AzxLUEP8Z3eUw
izPN9xOX+IkkBc/sZlAz5xwLksNmu68ywjKk3SsudzOj/v/v+1U7O/DhfJvO9HF4
36rQCwJK8eRbgejCNW2RAKQcfofzyS8vAEiw1GaEM8oJrTEGv92fGsWXS8TmuFJq
roIfjlnv81oThxwxvcNQliBTLOqf0Owc92SrXlEScIUF0/59Q1HVtJeEsEm3qFP5
g0nsmvb9qmRw/rGFRb/Ag6Qs6XJCJHI79GWwFKMsmRB6C+TpgYZHOwhsM8hM9wGb
Ztx8lQ0GwDHckw05YG6lpNobmZf3UIv/kIDl0pWftssC5zCuQ2WB3IzYU0oh2Zf2
SX5V6Zo5AR0TVW4LHecGMXKDLGD7KnWUw71IHLUIIgFSwo7RqwKXBT3myLqAio1F
dhcCogR4Wo8nnnLTO0Fc8Ix2IiKJ8O9v2gzaBu0lyDtduYuAtkw5IlKHN+lBS12u
cyS/2a6yKjIMA1ZjvvmqgmcePLnM0Fuj1e8qf0T5WmTcCQmpcxj7ljpPP1j1x6/k
dKaAA4/CU77anByDkL8ULNdzbVgJqLbguWbxTSPMQ8okESnqVkRvfi/ITBGXh/t9
/JOcsN97dxNmdcer+A2BOlJj50n9uRgcvmhLLBIvut+m14hno17OD1+rmUoJNDrP
CkHJXgh3Y82dwOkc3IZ9kKBzL86Tm3QMcnrHx6e4p5HtBkfXLhUDbgQcVJ0d1OhT
o9JWEJ24q67PZsG0Df8Go0nn9CZ6BkmjdCpHLrbum8Ab/XEbD+n9/ttV9c61qTGV
COfP991CurdsXlE1j+L5DGIUn5EaXw52P+NB1n7xehMrP+vb14YqlDSatwrDigfD
Qp+60yWU+vPjSDfLIrhyKfLq8svUGTpS+vmyRWJTk/lsFCqqqFj4unEO9cZBVBBQ
YMCE+nANDVe3YyeoQxpSaKcjryrlhnqriZFDO/B/UovO7h8vGq5wQ3srYFfq3ESu
9jKxQU/aTh8pE+zhn9nHn7wwQTajQOQcEqXD4uQD7Lmcrpgdicl89ZhZ1xNpV5u8
arWbEEC3AscgqygxIb4+rJv2u+Ww/U2FT2m5Tw6mCYs57RMfbss5z64Tv9C3mDzj
A+LlyWsPEzKHUA4884/28w70ZVl8NubMbdQmWVqI0KhPHDrhuVWhFtofYhPsEas4
LgMV5TXPHj87ZTAbNQLHS03quVHHUsULYYJGkXtkj7Qgi7+AfzWYAMOB8/9t3FGo
doQC/NZ/40Ho9lCMqSDET4DF5yY3a+tlP1jqAmpRPDUuBZX89dVZXUMlvsw13klu
gVo10ws0rpbeMELu6VqMlWatE+mleL5X2mqIld6oQlAjc1cp6D5cdLRFyC43B3dn
q91jtPSz/VdHNvVt8pB5EUD2bM7iBC1vmLoHGNpqWV3pixAppo/hY5vKgDUtKvHa
BpVDPirRXjcbaD2BbPwSTMCuSN51rYCi/KPFgW2blhJgQIuHijiO/7BwClD/S5iF
C+iXY/zM5WlFIBMeurjhqklHvZp2EoqFWWOH8UUjXviy1GiEpfjp9QtJr0cBOJfs
0LbmB1jIeetH/lovMJVxQCg2AJRtGXzXZweepOS7Fv/6zzOihiM4c4G0qGWsWJ05
+Jk3otjU/vahUB7SmenebcBfTSN7PTK0HI0PIhh3Wv7dswoh+oxMY9v2Be7QI4Ch
Vx9r6y68yoV9GSJOjC0iWmVmLsxladHej+FpiJQFAiFR5+eZUlMHxNtZF1cD8HsV
8j32o8BJBFlmLDHMkfo7Ac5BhJ+k1rqVu8ZPwEIpSCeBKbqoTENoqThm4cokbXCX
b9jWPxUKLeQZMkEJnXJ+8qgx3WEKFqInbhBdvF3TbvX0PrIBESB/EloXjoH+7wse
dLuQ2TEiu+jr6QtwIdeaZdcs8QCsIx55ubSlpXeNd9Wav5a9cAoTpIDQdsTpdrYQ
Cc5FbH02tCAgHTsh7RxJwxY/cF2FiqLV4fi4obdbRS8qGUUYW4kAb1/GtQLhI7le
A/kGbfIQz1kLyHHbKlBDmWyOBYqzDi9n9Tbq1ZzEYWjDLP0vjp4bkJho0TA0RvL5
OdfrKWzFc4Bc51Er3Wxr+ekLEUFbMEbSP6KMsO0cW7SI+7E1+07D2EHnIccTpkfe
F5oIv3IPA+y6QCGXUUAxEfpVoOxb7W5+idB7Nb1sJUFB8GlCr4qWEQRNXB+5Xhlw
4s+LvVhA5hnMxSHOE4xqSztGfcXaoSCQODp6ml5ITLChhKbliqtUwUlYDxuhGX7k
rdTJCcFRQlcXFVCat92+vzqOd4XbFD3gYIZEBrsaSEaLhrk4GqEBJTrNQnG19RgJ
iPSg+zU2CZJi5peGf+ZQh9ADlMu9y+ussm1YkUA9K5+l+HW/JAux1nFEZg1Ljhtv
xT0rOAeAhsTsTR21K9r0Y9boLS0twl9OY+p8pWiSXTSWggJNSv/D0nZgFv7RdRpD
YZkmwEscFT9HRf4cY1byFAsZf/jg5zGmNwJypsmYx/+wqzDek7hL+Y+AYoaJfaWA
+6fCAQhA3kdzAtILO1pclrS3rwQHq+s0ggqY6cwUkiYV7Neuc3VYkV3yaL4y3+v7
w6I+vXKkhVLIb4alqJEz4Xtwe4lrN6TwocRVuSilDTkUy8yzqEFM8jkKqCSxIUZv
RSSlukpd8EcRJNPKJqzxVuD0qkRiHUGy1toJNqSKI9AP1SlypoBkZU3H1twwDNMH
uI7oOMUIgkv+6G/poKJiD4JfYia8PXbfSrPl5D7qu4orHofsBqIEPM3SF1uOkNRe
832B+GSjZKX7TD+aff+BzBiHOfNldVHYx+FQS86hUzhFM5kQHveI1Ts7D1F1IbAN
Sn4JVf9TjbrsfXRgf2NqTigbkX5gAMxxrmYFynokoYb/8HiCfFRlqh50L507Q+7v
a/ppooi+2rGMmr12Eox2wbcC/VO8Um0SUL52OCcGkgQfFHLLdtJE+rd1Q1KZC17n
FInWV71ebQkg+HbFjPuwkAJZC9IOesAdmIVJZYNOlZ3oUxzPWqb5WnhhqKpm1a7q
8M7PzzG3F3HRWvOwh4AFQfToThqobyOWAJHUcIguUZA1rLHJFVNDhn0ezmR9dHnP
+QF5rhDAzDNU0vzPYTSAS4mJvG/jGrmIabLyYR67K9W6sQpmkodcfZBS1IcPozUy
rjoXQv8bWIdIFnEWlfB40atvqFBBa1lVk3t+hTSSt5qtyx4WJg5Kiu5560EMvL/W
ZdwGKtlnSr1Df3O8QOHxKzt+qZSYTWXbLYpMLO+iffMfJdfWFYm7bkTjXzey4Jmo
vPf3vHr1uaTA4iXMgyeDEQy3ZihtkTZMyAnlMUaFbi7tCVuj0Cm+IqTMTIeclsXM
dVNkvklj/qJFCVlhG6UXQp53laVFpoPqrAHnOIcTu9h9jihJsuY84WVBkZW52pFV
emn9SyA2nUogBjE+iFUBNx1O/p3Ag1Oso2kHCNCvXyY7VIRz7dLo2qM482I+gz8h
z+8Nk1VCKd3mQwK+xkW+/8VU7yM5qNE/eeGerPPL0g0dnjE5JdOCuWteyh1dOvEv
O2BQveuhjxRmrKSZJrFLfwDT9rGPhAQmpcu3CJuLFOEdrwecTgunLoTchYVMOHSm
CP3k1m1x8apFjZ9tRlS3C3ej1ae+VFzBaut9x+xuwKDpCjw/NGW6TizMzY+4JMcA
2bljVqYBBJi1YDn8avwP7PrZmeoHjFhEjpDEnYUssD2yoF3j7wZEOentlta0rAiU
gpJ3VAJWycWbjcWloWRxzOZxfRqhrEXqpISPaPeng8mjB+g5B9fZGbxYyASKmpAk
tj5x5aowkQU9QdyaFzTV7fW7I144uHG1XIy/rOjTE/A2jub+yNCxPcjDyzwlhpCx
AZxz/fruScrqskbllcg489HAvkSK/yaKDsb4/xbCNVhG2fZpcY9lMx4ocMWX5cW6
QTaSOgq0eYQW6+SBU95e+J5SVijZ5e7Thjw9rgMwFesn5qcJ9M9ot4KIDyNIC7j/
9D+1mqUcfYJBKmEM2UKiZjItzRrrJWRtHDIEkF1tzSkFVVl48ueyNN9GzCy26grq
YeK1uXuKb/lg7lusohL4JgDpgm67BFWZNsXoYIoOaPqhdq0yvNpBjxRWdPcxTnSM
0MRZzowqC5DzE22PXICpQ8ungInP0cG5JWNIDwUuSkMjGajjgl6xO4IKrOKxo2CB
gfn01ZcuTUki3YdHyG1cbkXkw/LYjmYiB7BRVa2LVAsLhMIrMDBwLFfVSAsmvm5v
shiIcavKHqxSFhiy+2uv/0M45s4vlIbWaJwoK+WCoVPIk8pS785ZcCUvy5wFIgJZ
SYbygT4DHXczygol8whqWujyzQTwBjiCkhMC4E2B4k9/bifA+7nEtezHQNS31iQ7
B2P7Ai4VuSLj/bdPYYaGyh/1XuUzhoHugSShNXBVW5VEcKyNg2IXEogVnodaxmWI
BVuqaR8r7cVYktzgpVvQMG0oJK4V1LwTcGXfaYgjuygxcOPEtHDYG0sUkdUN7YNW
Y8mLhEFLSseNIm5uUOAnYz6IxD+IJvF6QvjHDAHhMLeEVEKDz+S2f70sirIbGXVK
JXCM8uaybAN5FSvlCHWYapN6q0APMKw7uZZqUCcbUO4e+6pT0Urvtc/82RYKVIzI
3AqU85hVkoFnFkvPV3vzFM7OzXF7teGyRXg1wslw+0vOWtChRet/V3S00TOH6uqE
VzVlPA6d5UZ6eJ9MbxUR7AMNVA7MQWavstHKtvn7w/rm/hlJRD9NtCEErIh9CSQq
VVERBuGNL1gm5Zz36MeESqTYrvcBlvJ8I9krjGD0Zpw0gUi9aMArosQ98fDFYYXX
O7FLkYGJ+D7O907dI+GOR8F9sKSfNXOHGHW6X9C9Ih95Og7sbX3Kq5jRfeHHc3vS
5khMnsvl61PYcGsKyl/GcA+VYrqZF2N6QCNmkq4HF/n2Gm0833DqUEHKLXBSNML8
OlkzA0ajIIAS4RxV3J7oA64JZ9H3cfbyKQzND6FEr576XSiZG63X2KYhd0C0Kaq5
H5ubg+6i6HFxV8hDrKH0+ltirFRNf6glPyUOoUtLxz2ALE515hxfuzW2AAQiZASq
rMSX3/ssSBfnQSqmNH/YhlTNZ3iBS+zjRZGoXltJh5wkE16a45MhWUnUVuuSQgP4
Hw35GQk3N9DPfdWNZlRaHl/fIFh6qUNnqP1NmlPfbHKF+XW8rnGyXmKDH32acLcc
ZFUavoFxyVvETeYBlRbt+EQg3dMOSVLSPQP2m6cYzpmJZS99eo3alg6JmUdG/B+x
y5LW92cGhkJFTiDOqhLO9GYtsMh1hmtw6rlWmT2pM8P4TO+r5cmzxvHAGBEkF+EB
A4LiX7o9dckdvuKflgX1oGiwNAKMqCeU7klsGeibcJd3kpdTU/Uvs8FLU/emQhAq
xS3FDWZTr12YB4zTLenrgtNHgN3OZgBYNeC8Drh0OwwILXwPpI65E3K/mm+ZcMfk
3pY63c/rchClxKeUIHGgI1mlWwyUeHbu95/ar5K2qZ5RwhTYSqUWSq69ml1wGLSz
aIolRgJa64nz1XW+2nrS31JmTsOmMNgEXHTGN92bQwVUKAYariDVmfOhTJDwYW4k
ZXgqJuGkVbtUKNjSyhsKIV/BGNv08feF+iYw0hvVESeuUX8fifw3GXOjGdaSiK0c
eQVUGtZw7NAr7QaFi0PR/X7sNahGa0vANjqCU/w2KAH5+1uOHixoJWwKaNo7IkUz
dFIrGNDgcU1FG8Ym4DC/5oJjAP1Sc+LG+gJzXkXkkzJzvM1Tr4kfya3zq83PG35S
UtjBEKQJM5ezQF3hnRaiwHkZU/KV+P6138e/nFDI2LliwkKSrscvU6C4Xi5mwgk0
jh8E60bL69QWv1i6g1GXf5AVLkAlHSVG2JZTkk37keDZOPkZuyHDAG7ChsN1MWsF
vpbV2YXkh3DpNB+LhGypncbYpLuMU1Gr6owPVB3wHKDEbiewRsJ+aNo+k1tqNLT5
CHhqc2800kuJ2idp3zlcmX5HaMhcBQG5rzHLtCA3HTS7UhI5E9bTef7GdFUlkaGY
OFZjFXFvEXiifBwrKCMzHwCB4SVevddkLZ3YWzYqby8846JnkLK5wh/4Qu0rNMsG
EMCvyjC8LmFBjTN7NUVqekYhAxBV4l4qCiQuUIoLdO0YZgn8y9t+1KHEFQjYKiWI
ds95M9mWsJy2qo7ckEfqeldTM0lPxfyi72Xo7//B/smNoRyfo+BnCb9Je2lNAk1Z
Oyal9f4EnJVoi5+ahqVVZAVSjQwjD3TW2C4Fo6pSw3x+RiBCJnQPZPBZ4klq6j1V
BGi1xyKEIxpTONXmylzaXspV/MiPI1h5AatVgFoTGbM62UqsvFherUDcAwHlCZPV
glF4dbnL4Z2PvYcv+3ZAICJQTCuhcjLwLIhX/ZoATC0b7QtOFfo1QIJTv+PyQxz4
3J7+RaYE6L3v6n06AKfpEZsDkZuLD+p1szhLQjzOvYEOtVftUg5gKkZzBo+adxPm
n6WA0VTO3q2jYimBSmAGLo53XmOgaAIrQO7SgkOdeqXnzkGRj+h2tae8YCX8C0vo
3cxFFJvGFMyJ4vL1Hqm/I8a045xr0ZTLt5F3Jha4A1kFGsMadL2lmC2hvkknFVl4
az+AgZk1Hf0aadjj0f2GucY4hICKNHOoPXBUYlfai3iWkEE0HHEl4kfmBX4MEBlZ
zyJGbZpAFiuDq0bYeKQHH5Vex/hFftS7sre/A3cLFNMzoTl+iG/nOisOdOTTJzQx
KCu6zr0FhNH+wy3Fx6WY7WHx3bs+MPmFoICvyQaoKIOoFhis+7HhrRcFubJDWdrS
WgN1DuyddXv74wZEGxd9VzdGgfrkqh+ISl5UEy3QmrIjTQZb4/6ABOfmgdMYf+zK
Kc+HascvbWZUO2LhiBdQOKShD3JSSof454nvvMrydS6/I3g//n/kp0siNY6KTQPg
qx5yFY5LcY0ZgvppmnA20vZw7GszNNlPeyGlqK1CL5pehjIdSoOFcH4liqzBeGNY
l07O0zGSL2lbO0UGlH906KzANMHKSw/sSrbEZLWId5rX0KEXieZc4lBp3ciXlJfF
EGu2nXQMSbEHl5BXUvj3LLbUHhxnvBV+4uq6wRrCkn/Cc62fUFuTINhsqftIQljT
bOiq/DtgLz0jjVhyohIdYLsCVQc93peUAdO4oIwI7NbqqqB0Bz5BRcu14b3WrMg/
j/TduKpLhiwEusD5HAA7U2Dr5pkdFLERGJ/g0kimfY1pTAYl6ZDknQAlKMgsD9XI
wrOvxrGqrxyuDT/Dt1HUMng5ZznE3z4Zehy9hF4ftYYATh86IT+M6F0G8bQ2JOH/
Anh4Wa+s7aXQ5HoFJ1BFyVZY1XEKPpotO8/KGYLCx08+BuCpvE0TSsqxORIGBfZl
3a1JsMN2V6KlMHCVe/x5SlaLs3hKGrZiLbvm1fxqt87JcwEVvMqqnh6iR1mI3xc3
aq+1idzYqAISrtquRSmUpxIe951u7DRtcI1Q+OVraAOgFMxzuRpBP8tQg4Dv/yW8
Bq2Q0+nr5iYggFSupew3h1aWJsthDRKL+oX5U8HYrkO25cFrKcEFeRNsw2oMIQKt
m1KamXn6iNHjTvmP4RhRLwQewiZYH4Rvaj5MROBpArd8hVYMklCoy+ILPPbkhk9F
JUzf7l8few4m9veIyhZC8Px9Eh8CSbvuJ70+d2bNRG7103grkUkZ42CPLcxq+kUy
B2uFy41af+VBhAe+n3s0+nY2JIKktteNjjTLzR5FjQYr6Q5fCBxIcTUJeERRefmv
4PQViQtgDns01T8W9fW46F41O4MHyAflGKE65yfNN1ZmNpvl6ke8O5Qa5tpY819i
93NIHddngegNb1EdhrdFPHpkxKmc4kAp5p+piXkslb3Da33jJEjGLSjpuL1t7+BT
53tMwhu68QkSYvaza1pMWriA/iIrH4fENqDFcuIV5FzruZaxMItYrQmQFKXel94w
oVQqf9MqeqKVhYXlLeuSATgxGs0E7SOXrgH8NHpsDRx4jdLqQRjALV3cc2ek/o73
qHtwbOrj1CLuKfrEk1myAKHYYfizEk1IBVE2NXnVBpGXFzQLHy2nSZ+sbYusw+gR
zfpSA+0x4YYm79tQzMt+OThl+0xywFz9RWlg3D0a6b46s2kfAaPdDUJj+qMM/4rk
nFxPUW2IfV3YHl62Ydox3LVkj9gHKdQ7F61VkCmCPl/TVJr3imZi6RCp3Wqm9Kvm
iTFyJoRtUPzVJvwU8T4wGblMaOCt6V2n7AB0dTd9V5YBQlLsRx3x39+RDqEHqRZJ
XvwMQKKJTCEbWoybldbYHltXvogH7CkVtzzutqR4uTwxyI09nuQqjB0Y12Ncp/aW
vwspnlCHfC7CaLIug67+7c1EfI5FcajzSyJZR9IU7OEWNXI3LaseVV+3N704q/zt
/uotqg1uRkFvZihpZARbU0IXfY2XoqjvmJ5fTfBXWlfc785RMfCtmHMxhsyA5/J7
1GDS8XniLdIX4Hr9Swyf33dmBB24VLJGv/tYO0U49+97Pmj8sDnhUubrJCK0lmDG
m/29hRE/wShYw2EnA87RQu0JadhX5bEmjhkcgCVKf3EX8BeHEEtmZU+YytCufykI
xgEawJtdf2hBa7kpoaG15pNPnSoDWQ2KgjedCHzcGYASrod+pXkXv5N5iFHzlTzr
DtnIp7zVo2cYRGoRYxELFimr+p5/yol3X0cgzTtLiW9HArg3AFQk2z7AMllaAWLt
k9nJkI3UqiMGz+7el/bvtitK2APSJihxIjFKZKqSzNq4t2/aCCJoiARUom++BDHi
vx82b+KWHSBXcQhYH3OaNY29PPtxVuTTD36aH0JLAXNS+NZfJ7uLiIV5i8UqlxjC
prdvKsmKH7CPCqOzs7L+HJrI9O3/LShdF4K0xaiUtS9Q9K8Oz3MjJ7qq2L0vn2bY
zbr/WVGppugkJFmlb61Zbzagy8GYOTvz60vh7rEHwFfCQnK4heeILT/Mw+/lZD3a
/myPzC4mqdHiHv6PpQjJslhAnuf7xo/+ntIFBjsr5+XzdkTEg5oSCakpkPSELBbH
kpjJEziI4q5rZJP9913JAFzkHJYWksKFz/+m7GlsfayBT3qzU9RX4Jr2h6fyx3sW
fm3fTNgc+lZgnlFW+qANVgpv+yLSSom0WbFI2P+OIhvL1vQKfLUPgBLs8umvBW5l
PKcIvtwDOSfSmvTMu+7F+1xqcMvNJq22ETjkFvPPSVITGoTwoO9l/l5NaFbmSt59
csZCN9zGH/Sqi1ezaz+27W96zsDgckxnqdlTEzGt+zgUAlSb8Sv7QEufa6jmO732
xQd0iM6xqEK3EYiti3qXxETKhxj8MeYooJ42DzkCYx6LZTtVYQKP+ESfhWMoqZaX
rp25Fmx7aPCUidSQzRjANpBCqCwCltZ2CKh6Qjq9BgMOiAOJxC9ZyPyH0+kkUzI6
2Nawx9hgf90SGSU/mduWpfKlJdbTBP2wq8omdc1aVhA+gsnYRuBxC2FASiE4aBdw
QJBFZ1aD5t2nDCb/srMqUF3i271v7VSCDKjXEzm3krU/UzcPMjpDPYmf2TjrgV2N
vmV0h1ZxZqJ6NyngcgRwvYj1mCVkhvd/vBL0G3igGqrisdK172/acwrg6S2yv3/2
/MSCImzrmp0qnPdAqZw2dRR0TMEM1qPrvzFIXZbTzyfpYFzQgB+kw/wM+RNCC+zJ
HO+8M13mB+p/Mff9LXTj7hg2v7j/9rDb9VeFfRJ9Dov2wD/nyJV+ReN1OZYPMB4r
EjWuKkdg0h4EZovDUt70Vz6kp/K1FjKqpwrdvwMzjpOTQlnxmKRuyoqFNP8biOal
GA7RljK5nPJGMSb01DYHEZVaAKADB3nnRDj7E0GVcs2dqJ4CQGUBt0YjxlwiXHs/
VQqAqC4xMNkXyzlzL+eyYEYXkhK182/TEcyYTXAaXkMNffO7GWFGTf7MMBN4rnUI
s7fuE3RjtPo77WzuM/B6IszRTGBHM4w/maWNfWfonUmiG5Z3Lh+hY0woAaEjJUh6
RqTM1LS7pqE7JR6Kz9RtchL7oYDYyedcB9qCDjmGqkN3ak2NkXcLFjZqgX84/oeY
qiJg0tCsieTaSKaaPjWkHB3rJ/bPIRwYlqqMsHjJ/EgeJKQ21KjpxBHEn75MOOrt
EMAaYbEnu9ZALPbqDFxjHKsEes8wmoI68I3V4lTl9BIEzas7QeNLdkHvVbFoNOM8
8JJyeNJIRi1s1Bb/XyB7mQvhkhIM6oJ8hzn/Jfc1A38D1TQXBAh5hnfeYblo80na
gyc5lXRqL44FTu4IUY3sSkX6l8yGYRgeto3uFJiV8BB5C4NuNlfOtGWbJa0t6NV/
iuz6222+8qJ9gjfy/9hxsCeLxL/tegySltGetUUHuVEx4x5MRVz4Z/9dmypzOlm0
gxJr6M9btGHKyrXgKRVwMpUXmP3VGXTdssk/cLltXsi/u5nuJSkkVfGpbxIExiGN
HIhI86EM8UbXGMoj2x3bAgKfTvNEc+FRosiuDxPBR07xs1mfKYH0vX/caQDElstQ
YuSYiKpXv8jhFBjY920fwrZaQwCBinKNzXxGcOO+/15U0w+3wJO5PT9Mc6NcO5Vd
HGmJAXQQhPbdcUtqEupa9gdJ6y6Wsncdv0EQ0LnGF8yZrYcWJ4hMGo+MbLhJmI+i
yM3r5mtV7WntjmTTFz7/6MxBl5P3MvQ/BEFIdp9zVUEMXx/aFj1AV6l2tPVZu10Z
HjcMbc3xMf8rp7PIeQvXxZUbLHujt2heXzOt6BnkUBoRsSF1P/Y//wiWLPMrjc4y
pfOSDrUkf+ONjr2OF6JDeugo4tPBjY6O8ggLd1mYNljvwFzu5qdBlLUzIiw2ANbV
J9wClMtm77dpFIwGo+VuSA3ivF0XPWRxClRju9kjSroeetMv7kXjWLdh2Tr8VYm5
AeEQ+RMsRvjXYqJQASwhtKWKmi3x3qkYJQHLCebArPwOrkOVOeZkmQ+MDCWhQJVC
ApXxMo1sB1sa4bqWScBvP1XTkCkuxdA+zYJIT5vpiQTZPd5gWO0MeHrRuhZ6er1i
MY4pw+cpWGOsqrRLDBnyS6u2zR4sKUs38C3CowXZ/hzAwwTCjuu/vr/f4StMoFyu
KYMnbcCdMWwe2Si7LzDDkEw9qmq/EUxMfm9jH59kFAp+u50DeZNrRAiCUof/Ygyw
UJDfpX3utkoAj7D6/F6lHAPNutSQrqWQXXY3Q8IEOMTArnOyE/3rwpHdX3nwKKEc
uMETMZvgKiH7AhObAMeJ93EjlWNz9BZlBzLeRhV1xULkExTAQKLDDhTPSdDEdBB1
puDVlYHxc2CvXNSiSVztA39qdG1ml44qyjXXm9cJSJwS1FjU1yFkYiiKxSNFuch4
eJiipX4lVVJpRs7yPn5FDcMJ4kjYuH8pkjY3r+w5kDyl6gCuOWoiiYLXTgI2cRFj
PIdfGoiySJqtnMwCmSVJVQRGqZ94PmKqhH8gHKD+qgaw8dmV1dsQ+nqToamzdAiz
Tz8fHt930pmq3bP3MsQSWRvMgaz1+K956kb5NIs2HU4H2PU1+KN4MjUOPZ6CohHq
bq9T2oXw+pa+eCpSigdkJXgg9cotzh+VocxFfVqi+tqUPKgBCjNeBS1nneTg8yda
+iaTgfJBU65TMxpUt5PgsCdDIkvtzGZMB43WQhz6lJ7N8211nYQVHakA/7TW+62U
pDIb9st9+kxAG32XVfrc0hrv8Lom7CLA5gVg3ZPWCIFLRWMoeF/jdHCpugdBMdG0
wL7r81ACvLf7KUfkwuPPN+GhwGcFwE8fCbGpTrQ9QXTaCe6SyJhNbabQlm3AQUhB
iXiIzyo2e62AcV+DGm1N5Q33UhMdf8NvZV9hYJZdBSewcRW/DPAcAabN9C31TXDw
RVTCbCqF60OYqVfkuNYh9fx/Zwv2IgBXq0VnMgCH8IFDtgA3DTCy8iPzGIoZkdsS
/ZfeeJeVHUiahvAahSEJin4dGYL7ez9dj/FFF+QrqlQRUS4ZXtvedFDQV1F46QsZ
0TQSWdiwB1KjFAeqfRg6gndm/bB3kj/P7XyWbOr31Rtjj6KoI8Wb549O46CSwCyz
6qpGzt/sDgD4GC9DS/SBIF1w4QM6B6wCIDmd3vRp1lwCdgriWAQCOxXjDZFY0H6n
c00MhybAHWqijTjmZOqNZZW8MU5fAfBHnBuYMELyIy1777fgBJPnoDQghuGCYQvn
U1gBTJbS6qNOaQVF8vR2ROeB89s4cGUryP9RPv1fRbv/bXII3skSUaxQOYeSucd6
JMd4WnrFoJStRO/NLvR3HsIwRHcOhLms3elrzRlChwnMphN/lsHQP2uQuUHtr248
8OoZ9NG4h2lbvBsE1jeY0hcL4C9B25iHx6+kgHISX79Q1dOx2vz//epSpaTT/Jr0
CVxVyr2jOBusuzXRBdvfz7AMysXfbl21ahgIzONKcs2HU/gEFp17wIXpechnO8L9
95VLyQmavLRJKjPU3gG1oLSSzdqoYAd1Extv7F0ccnDjFPB71wrXT2rwJFzM+h7Z
je4h91uhH4ZhU6qOuVUWSarmiYjyMe7M22hOyM978Gu1J3mDrA0DT0H3PPd2etDf
hv3XNOhyGRsrtD92LBMJeBxdhWMQkT0TuD3YOUSnyM+ARKS9czeEtY3e7aUvk1sD
nCwlL+Ob7P8DtgZeSHrcLilTp1tWTMwwjbkz61XKy88f2B1nzfXKmCOBehdZVjNW
3512iML09HQi9b5VKf8ZHi4PokNdP28gYkw72KUqUI2UvWVTVAMfmK56S1n8y/7A
BNkvXM+7USCmE5QCgyEt4YX5YcjB1qQ1p6rhz2miofbuPn/lBG4VABe+jOAJ2uN6
VlzbihzZBMg0DZwTB+e/ggVFt9lw0ETUu4edbKDilF+AimMXOU+AGFfpY6Vrh6pX
trSFdY85G7pkyW9xpUqtNp+KDK/kbeCCBtovREhnuxgEvXKVJ2/vrry8RguZA/p4
svueQ8X+MOIkOMjlxiNYYGLDKh+JyVs/qPDeht96rBahQgY4oFuE1ldbnQTu7wpM
uEzQdv62qrdd5lK9W0I2+e25XlenfQkK6aJL0fpb7xHeMSkIFGHlWAozNmN94MGo
JtEit3OBGTWGWZgvL5WyUPpKNaMOeeZMmT7IiFizeyvhsnBJ0ltDC5wwthie2DSB
uduiYXNO41vKc23IdL3MkETyasRInIaleReYgRU8GneskcbN2Ag8/CXHBQN5+k4G
SM5tm8q4EC2DVOvzFmE5Q+wWWx3rShC3kT26+lF5OrX4uc6UUhEKAYZZGcdcLDb9
5iphXszOcWCfLoUrVC4jU/yd3O2czFSD83Lyke3O9PD0c303nQX2UOYnzqemmiXJ
ooBGyjRQDNTG9LgNuMn08fzFhqgSoNx4V0aPLEdTic9/EC/Wd9Mc0itaSOfYyfV2
MO3Jq76K8UWNJqwVY5VfJtPMcTUesBHvmuXjxYtfBI6J0oclRZLPlXIxgTw7wVB8
scXZrsApGYVEWEb32FpMy9DqFt+nAVJwdHtFVPO2xpfPI/Rcjlylhocj4fDHpVCS
Y636/x+qYUO2c4l33PGVWywsmElqAMy0kJP8NVovRlQI/TOJCZjor9aegjGv6NA/
KXEZR72cqv8CPVthapLkvEw7sQGFV6vym4AI3jaY5iuKlgzKH8iB55BPh/h7rVFN
aAePZ907W6HaPq8rMcAGiXcMBUGpSK9VdBLS395+pLkP3WrjcQulX7YurTSSU/eg
o50bUBO1iHzpGTu+W8rnemxxsMONKfjSpTqP5n7rQnqeWBhtE5kPwbL/Z07f5GkG
B1M0cMO35fjYTIAAlpN1W7w/q5pIQS2VJYww2TqN0vgITJPPpVbiypW/j2A9XRB0
iMLyaSzXUx9TbJlKZoLF5FpJs4uVtkMw2U8hYM7DFQzn69aqJjLEDK3Tt1Vk2SxH
Cf4DX+X21wWQozwk0MtVD5T00fqRiKyHEQ2Vbsh86br+/JqOYpZmVBDzrHjniLCp
r/jxVTpJkBlt5/xy5ahPfU57vd0EeP0hriM/XmuRdvz+o0GWh6hTuG/usdbx7S3A
AUMvCZHBCNsyTjoUMHsMXFNWsSAVir2aViB7P0cPiVSkw3ekyvGVUGqqWMu3QpjI
VPK9kZqqCDY1InZvKjGPkV10yvXEot+aL6wwuujJ5KWFNBhcKZJZhKZ70QKb1HSJ
Wkmy/hKsq7bQ3f1jNAREz3boh09x1/bL4t0/B1ho0wQBtDTv4LbWYmwHbM0wVSEu
CQp00WJSb2z32gT2qpQVdj6JG72CeK5bE2w9c8eORDKngReEHxmOb7CL9cuNH4pN
cViw1nuRaqWgMCESmoYFg13e2ES8FHEbbMs68qKxGCVsf5PbvZ6R1l+v3uW8qzSo
s1ZApkjA3Q3A9IkB7C7XyWu6oV5T2eTFYAJ7zcVv/GceFi4heXZZL/0VSTkmxekJ
6PHPhbKPVRSVOSiKSMTEESjczkTObil3KCbECI4SBw/Lv6Xb/WMFIektWvF4Bq8v
5YGOx8YZwFC2uLCB7bOlk/p+sfiB9DqrVMG45of71WSfrNQG0zBkJXABwBPd7KhS
uqDk/krXMcMWBb9Z6DHbPgeMTdB/n0+3L+Y3h1fVFBf/riEtJkMgjHz/VnlfsSVV
tXjDBNX6uDlSbqDazk4W2IdZJiOTqi5RxNLT1yu84SgULOpt74oISKt7+zIJD3PJ
Ztvgln6amzyw7rEcJqSkq+cF+fDeCm9/1k6joFJvxIyMeYCbK5FHK5A0KJ7sL0E0
1qbLXc286oaeq9dSS0C7vD7pJqQw2OS3p62TJsRNZJEM/EG32PXTmedAmdVnYntx
y3nCrqfphChZdlNCozX9s37J5Q2ulZAOVv19uQCJfhFTkOmMh/yFEbslJ4SYuJjf
nG2N/pFU2xCkw0pgBDvSpQibz4ztRGBD1nZwXpWgMXtMH7yoVDCmIjhaSGgSTOs1
k/kMY/gLOTaaRAhkHIHiUXT7ZktZWq8yJR/x26LS5SiPp6kQ4BXEUrUrlK2gZ4yZ
Usq0grj3VhnZG5hCUtEgjVT2gsihq0o3kk/xm4+F4V/ZH8ht4bRE3wABCNOQ32pG
eWa1e3jJBrLhG89IEPXsPhyRLr2q8ayXI62ASokSAafrwQ6GDAU6P5I0RQi2KR1A
TyjH+uPA4s8vyd2tsRHI83Wq14xTysO/9OudwAYm71j8KXzJtM1QXLLFVn3R3PMe
o9KEJCEyNfo0RjKswyvFDeIBeciY/RQXa1Lggl7KzlL306lJhmj0743UfwkS7v7j
4YsbKqxiOg/9jZVle61lyw62op7h19NGU0cR12AatOelCK7u9zcgejKrghjC6FPl
FOrnS5YLlXpbxELzCfvlsKMAF86vZ3ieys1ygOr8vHir4W6dUVTZ7H4aHyInphjI
B3t0F6KPe69Fqp/uYTJo35LNJ/ggle7sB7mP8m2wgwLBBlpLq85qMB0w1ofcmPRA
PuaQH4WMmrdjwg4CbaMUQLpnsbrd7CQvEOXT8mBAXuVPPbQGrpLH6JJOr8iXTJpK
ZzAltr5aeU/5FDga+mTKE/RAfHQH3eyLo0ZRB//yujFzsPNBH3GOlQayJg7kxHrS
bmDzVmRw0ZSriw4ecUO9M+ioUkNoPSvakzRDWLmj2o0a1YEi95jxh1vlGvnJ8LrS
yfGV/lQh/QUfUFbt5hM2i2aHxumkfUpJBKjXXYEbFm7+e/a5lLN32ux64BLhVFgl
GPj4v3PtjEhjfyp8kdrDUsFpX/JPlPK+Bxrkaf3UcScRWxv+2P7azsOoTolBEYIq
JF3xa1rqDUPZTb7LoIUO8sfIVVfees0BlAJrnY9Dy/ONgBeZcrNZsJJqF+c5ZP1s
vMs28idz1uds4l7ON8Y19JpxYlY9Hqrq/BXatb3OO70JesO/aEPcf0qe3p+gj9O9
38sFyrzdt+ojtPVyEz0pWfS+rZKfohoS8TN4r78XPPPumDPLlCmJogg1+DDS584H
QD7oZMI7ImDWLKc/eukgxdxaZseGm6CYcAcbFL7ESWO5jbQBVSYopAS5gr2IAyQe
FpJ6tgzbv2sq6gt6jkVvQ81v/MN7dkMP6Bpvsmmh6kQczMPFbOFbcYQnOVvuaVRw
tqW1ndwbDAa5lnta7gshrHj4ipJK5AMHauV0gb+vfU4j1wv6a8L/XCuPR7uLPQzv
orup432xaUwTxKlSJFGS+KaWMk1GdzjV00wIC8NSNGJdEL1/YcJa68bIW5ObhQrX
28kfkoMhaeLpd1GJjxrj8T5z8Bn3uHgmrZbKRiJyA+F5j30E6AVFY2IXCiSEDzCa
eajN/cy+FmdhXP5HpBvjBQnEWBZAEfyBwrFKXSpLZJ84BsW+K9+iIdzB1I8le42/
LQc2ue0Sug1gyR1J1XIYwU5xNg/yVQKmMdrCktmzeqw+MnJ/We9k4e7iMFpOQiMH
nGeDX8AM7cJkGrFHUIZNpMf7rFwjBBpr65IpkP7FHYn9RPbuuVu9F6FP0g7/irpr
3QR105AVYiv7G4pcPNqD40Pede6ImxmfUd27ynRIjWiZU1yED4xwdkoeA3/9b1Jj
4vfLJJQA+FJIX2HnJqV9QWMf/rygH1vFJeRVxVGXao4WyJSOqsnBXrne/RuFOAbE
/H0dNPU0YoZE0S1gjm5A3X4/XbqXCkTPO1J5+EdIHgwpU2PpYdEnWEoyXkXweaHr
j8k4/hbKl5oXc6hN0uERBwaONEYBdSWXqDGluSuc9qvZ4mNEJu+uRY99p8m2SQ1U
xF4U8nWvdZ2Qs5hnNwzZxS3psbx1RAkxe4DLz8+xLC35Mo/8HAsha3HvBpA3+HSC
aZ88u259CYdq2E6kwtZGNPWND0KKtwPE3chCp/LwZiyJwtDjgsQtn9Oepz2qcv8F
vacrBWYInStDbTh+7XaoGr9uqeB29hD4eoqRt2bpU7Og9VuTmhe/Syt9zopxI4KJ
idJDbFI9maYA95X+s9A3huwNuRTDiWTPu1S6mI5GHXp5YnqlUa3NzgfRWem3hNAr
v2NvnYaRPNs3dd+AZ51UdHJEkISjonHbHYCQZRowrUOM97I4AE3f3xldrrlgITfg
aULv207Ey1xGlvdVcUc1Vc4MMAYWkY3A5+37tNx75t65X5321P+MC81AMdQpLbd7
gIA5JidZMb9BZM9BynVzNCaMbo0b15SqJNe24/GJifkhX7KKrMnbnfbBTLFQUNlS
XzuwABlrTjF5A5k0kXDpzvSmLC2IhGyi1/fcbduyJzTw4DQL9rPosSO4OyD1ghnb
E1GXjVI7Od/nGjVAtxpv7cJCnVw1k2TpuhRS4xs6rbMQIO4nqO9BdN4zPV68LbWt
p3qInDW2lC7Ovs9fLX1H6AoL14Ea4pRlp1Jxii7I3hXAGENAOjenz/sqFGz29zWE
dfOOob3Us7KLZoSZpx4zL59hJreP0q7H+6RGNOUsBrdKVSi7AgdHMXQClSNH6h5h
EIqB9bBR5Xjf6JuUV3e5/gEkd7WIJvrn3sWCjTBiELUCtq1id0Dq/kxokM0AKBaC
JwNkjiQHqyZ5gj/QZBOKc49uie+uvBP7IU3V9RCxczLUH7fID7DlWor101U5yTYE
kyS9Uaf9/Xo9ImRgdtIdLrDYgf5Jyq9GQ9Y0/kKTzt4BQMXLzTCApAJ5FJqK9QUI
/SyKnDmwZ3pB4Ogtocj7YagscmXH39LqQWrVVymQNT7kjB0MzHyqjy7zDYF38BwE
FT6BoePVGuXbxUgy/NiLaEYDsu+V9qx6jQqJRhBDo3sLbxng3Dw3VEUQBw2eFKC/
U8ppVumgon50/MbRFr0Xp3kRajM/Now/mCc3Mm41Gtgqu+tSP3nEz2fdd4vIT+er
IBOPkvwp4P9DHps8/p9GTjGo6YdQXON0Vb6liCueOQNH+o8GHbzwsgAM9oqGW7Zo
iJFCY0ljKhpZz8Ox9Nj0frZQgNcVsZtNirzjb8ps74ZZPkZfpZ5TnTOmOgykWHhC
eTU102YRGNRXebX2pVtHVraIYVoLgIpfC4A/b+0zUUhY08urN4FKBww4STT3TPjT
m0FKXQ70puCAkW8T/MgLvVk63OEpU2u2HnVRK+PRR608CnlJWW7qTXb9c0QLZwBi
tb0glLB2QSPyWg93s/xANJLf0kVuHDDjV1ZkB+8I+9laWKk67NfZq/hPw8Z44xhR
39iLIfDNap8v+vLBMQwWOF0htTdOTM32VQ13DQ5yhne1cTJZkuBB1O8yte21JSTd
f06qoiZJJX8sbxHxR+4nWh/yp4P5pLTrsUyx8zl4F9JjIlA+Q0tBhEmUnuVmytJH
+Oc19CG5ERsr/UG5yR+v2P7R6CYcTycbxdgWNcym4II0RgLAzH/x90gVPm8z4FVY
uRJ6nLaRtHDFscHh0j2Yewr4825XzvAeM/H+bU4ax3WUgzsbmerkLHPjDEn/40uP
AA7eO4RQjLmk3uKWw4o1268SMXUzjMTlBimHxH0s1CxPfCZqTIqnk1zuRd/Osks3
61ftddrJl6QaNblE6ccIgAF3f/w3VW9ONzaTTlonmpgIszeEvMIb36DHTKyf0YkX
46O9SVW9yXzhWcH6C70iO+CDpIVMTANDhvY/qup8MhIPqAcNL88X74zHXubqE0dI
IGtJ7qO/0SL8d1+e6PBEnXhEca1o+YoyFSWUMwbvgzjuwiu/gl2Kg0dEccRZTGtv
U7+h0I6MpSRivpPrvNrNclZ5otRcLzOZTd1IPqY3auO/T+Hgxght85pjOAwJXLIH
oVM37WiZO4L4LutT4dRB40jDKwRVhKfwx38/fRqEL9AoTfZIemJlqu2alizg8sI0
YLW2Y7zyv2122A0j4wQzSKvTrh+/u/2Ao7FsMFjbj6oVCzcaYAtZ5Dm8PAa0O2I3
CMf80kvBIPfwlIYdvqkX+NDSWzWNLL4NqFxlKswe6BjnIjPfDWBGLRXAExy3cPVH
jliMXFk1XfXnrUMmF9+erveS6v0t5OIN29ZUnnXVZF03lqvjMCPUJiESIPWOlFRJ
Q9NfcnQ8AxNBU4JVy2BkeZt+6nPDyv8Uz+jogGV3iKf0gac9SeIwm7olndjC3cul
uIbLuqJZ5AiLvIoTkmAJOPWLre6wuYK7TawO4sORbsYRVMbx42fsaYrIqCz4n6uP
64dec/3eRYvl2paZG3p6IzBbTbYdrFZa6nVLC21VvgR4+DWe9DMFN4nADeW/iI/c
iYLzyBx17GHND3gakJlblbsdm6TOUl5OHyHlJcVEt36f8gDUtD479qZCYBazIE+8
bWF3WTOr/fIXFdKlL8x6ARS60YtRec0D+qgVS/JSxSno92IpuylvXS93v1Dalo6C
LImt3wizhaDo/0KpX8L9uojQCNfuJFISEd4I+ev+YDPVM9jw0NQZAPQyMudFlb1m
fU8j7DfNXeGtCeHuDDGk7cCnq3DE1NYTL2/ly+ZqUK3YcQd2S+IfZEUhVnbXu/HB
7Zy5qe0OJAPqJtvmfzkyQOaQ4QtpO/TDyVSlyk+8FWNuFbppujC29+Ydup9/eJ+G
d0lYsDhdusRWtSMuxvkwZz8hoyLf9LJmS9IoQpJqqg05vcKlWIrfo3V3L5DQzmmi
FwHE8+ayIE6XJlG9QgTmAGpJm/WCThv9JYnuFBwnMvLEdqk1r5AhJL320ygLxLus
rv0mLBXCa/Yta27FaLqqnviHEP6f4fbhzLZyrd8tsyywarrCxrUtek2CmHRUUF97
i/ZtdoLCS9hVpEN4OTM6gcxYcFlS5XUGscDIGySEX2SasBewPgxbOW/g3xlAqbxR
6jNZDtCSTgjCHJCCzeo9yQNKUdZqPriyTeodRx28XCf2j2fe9FrUMgwzok4/W8VA
5LGHzFN/wJi/q9NmkKrfg4QIcqdRPo3L8wQkJd40uvYVd7tapKrx9mX4bHztPjEy
MJw238vcEflBWUgzzgT7AJl7D4TzeU/BilkE+w0dKLhHxjpDYF/SWAbK/2J32dvw
C2U28tbDX+aVYcP1N0I7skVLxTBGnxMU7dUufp+5DovK0U/UGibPf0qwSmDeNvqu
w9uYk9IK6W7nGWN9PqLLHp5r89O/02NkdyUMN/CliGVxl6Okp7ENV45UyE2t01LK
EQoAskM1tU5jumXz0HTNpUZiYmHXIzM/H6ARk6J5FTsAJuzih7DK11ZMwalBgI1H
d4taJHzTowoN2f4/oeP+ux653M1srldivJu8F6SSwl2yeMfxDEnZ/Nyk2RQu8GA9
LPUGrqD9Oa4PyzmEuC/D6R86R118NtK4MfyPUsA7Xir2x2FIkWc0PjP2PZCyzWeb
Hu00M5ZoqTeLt/OaMRdJKaqmJk+CscHqPAjone6g5BC2HUWsJA25aFVbKMWjYVTp
jolA2eJNBjwaHrscFEqpdNMZaYBNxP8bjOSQbO+bWnB3J4j5HBG29Lb5qk5xrh1F
HBUTZEV6BIPyacRq+R5ENpmrPv4aOHdVKSwPqTOjq1fSSHv250fH/5/JB8PI5I8N
IFsJ1txEUHyEeLDr0f6HhUVRUHHG3B9bDXjI3dhb10XPRzvZ8TU9Gx8DAuD/LCiN
GBbWgDDzFK4NLqpaKmlauyuwYJGZlvqCWhYGH+WoDYp6Tfjlisc66W9BX9I7LVdh
dcFsUAnZow/ptYV2AqIvQ7wkTGUQw/JngSlJ4xkJ0jL4+mf2XL9vq3GZbbs4RcRe
bihD7WSgzFyhT6+WnZYPQNmVKZPW+5zXfeA1heV6HUMtse4ApBq19t4DrPR3phqs
cj1Og0yBxIMAYewLP7aG247RGjZ7HfSygLcM0PPxxY3nkJaDODKAKs/Ie0bJ7n9w
OW5fdBmNg9BJjlZlX12wBwWJkQM5oFXrjuB4XwlIqnOOqcoFrFDUws/tv77ej4d6
M9DbSKOAqdtvwVSGyyCFPqBH+YKqdN95zMrPkthRjJii0gwRFlWHGFJjbjWqDNKT
spTtuqRWGCbrvuqlL0laGPDyTeAQ9CUqld4LUBM3prsDKTd6sdq5hdA4/6v15rOk
UTCq9Y3hl/F/WJo/Qn3PnAHyn3pkNWrZL6wif9362wuHOYRuNwt3QEijEDaXQn6p
qcUu5X77H7mYG1CFEweqyjsoRBzzeOy+LxfKuNOrEeYja6PALNgsmr9yMlkWV3Dz
AbSbBWYdcK1JXePSL+SPUuFFrYhUgnKppgOEGrPqlNVtFzNfz+MRN8YYOxHvRabk
3E8f2YfU9b6CUkBXK28lC5LHvRiUVlS1JJjmoIEEb54n2jazSJpwPUum/kyA3jSM
FZv2mZzI83r/U1xBs/YCEx9HDwbYGMkW6QwoSwVmsid/OV8LLEpX18GgnAbBoMQr
o3NcVKOLPh7UMLHJTUdkYVE4c9PgXm02IJrE3LtBeAPIA6G4AYvGY5E+3M2gbgCa
Il1yUg2kdAr/MOzVtZj9T3bBJTVL0IpwlTi7clgE0tvT4RmfnQrxbZ3SMuuMdhkA
qJ5wlisAi/pDK6l90NLOG7WmjSBtSjrabwQHyWQdQNbVCgpZl+n4lnwGAt3HO5fw
A5vbH1Fny7oWckuA6uFgOE6o4+U7X8Oy6pAqxXLryNXZQBFGfk1CA9wUzMVx6nht
uOn8/0tCFc6eKZAonklJqyQO6hTVNQbFYFIZVnII+1sDT/m6+E9zrI5bGI/7RE8s
gak5OLIN1yrOj794zNOf4QJZ4kRI81MD8ofh5ueyYFRt6jDU9/MAzDWBJpvaPoFm
Y/Qqz3IR46AuvKARt33ZZ7xsEyvWbHNBR/sR6oo61fubeetQFjhFxIVJ2NCd+X6d
ZPuvCPaLGTXtnU21w/XdAIIxucHk0HKsdMYDDjujrsEurx+fZNNOC8irEDfNQSZM
pLfqQzZpp4i1zjz/71UasMqJbvGZ0Jz0kCOzdH93gPw7uJuQHU8bvAgjRChW7+1z
/xOCb9OXkLCE4uLIUoAN7csR11W5xRtjB8B9Z9YT+Psxk8zhB4gJIidoXGWvXkcN
WmMhFxEc5z5BRh2Pl+fxNCNv5keZdkYMn4DEBOaq7Niwh9qehpYzGZliY1viK+9l
UTOvwobX+kOUHLknSMz5fU87P1ButKADMpFzTxfR4AguhtlpZnlWnp23x+EZJEtE
upmQQHiM77+yaCELTbwcRa9q9f+pD2hvFYE6sFoFQWy5pC/ieXlrb50XkCdegurv
zV3Xh7qDpzsjA5RolF7EFU92yXa0rKKhkCro2O3tvGjJCHb8Gzm9lm3hw8fmY2cS
h518rytIT3Ws4UHDGYAlF6SMVjHsNr/qfXCadHHPIXRhgjjCV3h0RaeSMLxzFYPz
Ef22XJ2xJ1XiBQdYSn5CO14jao6G4V3zW7VvphvqsuipFifDlaODALQtKkup+A8w
kA8mF4k03IwiMKhnAGHgCzmcaAy+dF46uPnsktvXJyDJjRNJMEYxj6DVZH0Zl7Sl
ZlNNK0PopPzfaMFIkHjGIWc2jYqKFc2RCMN5KEkthEA7z7kiwNDNlpw3M/GfbuU5
s8SBYubhhB1kTr+dxh9s0gmDWLQEeDT32GwhakeI3bNQX9puZDJWYeRLeL+XRems
wadzl/ZqEteKDeeaF8Ac4q8dOiSDnrBGIVrWKOh48Ruayn1kIgQrbN+zkzqPqkpY
pLFUO8XQgN5OXJWoB3LBfm6L26b2CfmJRI0nKje5FdMhxUP1xAIHHpqYzyF7JaQI
v6VeHAlz+MyaI3MKIBH7P5g1FK8by33s/O2onMwGdB3QApB2vjihzyLxsVEoW6Cm
qcLuZZG1JaZFhfmkAbwaggFsVqHJrCXpExxgdx/k00xXIbFuJKOEqK33JKBC66x8
A8ThZ8U63wt7O+IuQB+8uQgbainS4bS38umM2XEATZs9PfFzQVXPhB9iQywzsvUU
LyWxOrEEakvrqiNSMvCjooyQ6o6rjSIdk9LAY3rW1WAY66qI16QetlSm+K+mvoC3
avXph7L/X1qJRElwRI05KLlXgZvF2rqvaSTl18+pMt2wF2h7osTEOINTvPUMZC0n
yOJU2l7WFP02HtnQzM+VNH8c2PcJpYMoGpd47vZzc4IembnGeugUdYdvnBMQjymx
foQtcO5FfGQI0JYU/pswF3cszkNc1p76G8OrM0lMvwuCYBKKYhScBsu1VfuVgVVn
LbG3o4cS+lyar5YEO09uD6SKahG+WyYT2elLwSVaNzSJLuihINdlvzteNxDoJpKf
bq5tCEQ1ElhhezMWAvVhGtQrC2OgM0qbkaBs6KSComYqeziQBRDS/R4Ef9fdh2kd
8sY6bjt/lHl02lofhoQ0HXneNlQF9DT3rC9WbpgQmYW8w+0hUxNJRK8LDigvev6f
hkfY2t5vLa3w5eb/NNLR85Yx20G6gGk38X9sZoN3dzoYTudjUEcbVBGWCqU+IfCu
L5V2nFm3WLc0yo4kZ6ILVSqpVDn0Ly+S11UDDj2v9ZCH+bnwwqmCq2ijuSksbukl
ToBl72IjIrPDyG9eqJ1GPCQUjnHC2kS0uSe35QDStpZzRy+/C+MnPDTPCqIpFAXF
2qQFhZSiosxJh5Fxp+1IOipsbrarB3+H5KLtBqkpIqBiSe6OP60+nhCzM2b9ilqX
scdrSJWCdl1M4jgCuK1nz3El67PxC6Gi6zPnx9fPjkFU/z41IvmiZjtSwPT4tpRu
1gg4mU8Rrt5unBKvt7pGc2AXGz8TNfLRV43+9Bw129At0Pz/UR8ocSkpFPfhQ59D
mM9fKAyrkgcLMqfam0pqipxnI7Uwxvc0WeZ0D4201gsHMNWGIQIZKGV4GNtnXv71
1NhzvZPtMO+1fTA+x98klr3fRJqisIJBfWoNJBZyjQXx+iEzuemm74hRJuQ+LQqP
EplveiK+eI6JFcWDZriMDaIkMVXXHgbEGlpIP/AiDB+YLkDQz9yOu4uYUJSnG8IR
AHsR5FGHEGNr6eYfy5pm1E9iPxnE/6d3rHBHD7pYtp9wDqo1pi4mfK2godijcipE
dL0lqSFW0fDGCAWKuxO2HKqKy9als4IBVM/oiWfnoq/7MqqUDAKiGUYfmnrBynu0
pIK/Zp47cfxJro78arFjMlmd+47GfB/eQRjTUMa1Jx3DI1xLv2op2vbiMNmtxDuk
pIqjieeyfLjqCa1bS6VQn/sdOWll7ta0DcftT3fvLB54LI9uH5J0YJutQNmToQso
Bz6oERvAh4veXyOvZd6uTXaI897CpUbAa36USObxfGkZA0llBvuaxumHXW6QfUY/
BkVBM6ilMUI6E2Fd3VSGbU1Jt/JgSmXZrplCuzq3MKQt8E0Rs/Zvi6qNJ3jvnTMC
5112SqQDIK/2yFMDdmWZNKaLpewxqD4CtvvK9flzh3SrR+dItT9ktn1C6y/Q5Yot
DrMZSuU4+yMoW1Zt1qZrfQYBhP0MsUEeGveHcUMg/Br6ajvS8on49mR7bXFWf0xz
BA+zZq3S30AHq+vHsVm8W8dmJJVVDKwPhCDDRF/59aIlpwi3aaX7b7VVxCVht25z
4Ya40sbAFY9sCE2YfE8XTKLwOpBdX8AcA/NP5NsW4sReA2Mv4k+03ex1Pdx0w5Bt
Ig0hkArAgtdTfo2+XqAt1Yfr2lVLjfwHkr74aHd8vAG/wnLQdUNeyiqfler6VTcB
qTQtobGxVWE6VmzPFSJ4b8yDOYHW+h+eePMPYOgvPYWjD37Kg2xOQebpri1K2y6h
QbBLVLtb9E/vzeHXTF47pP7WPduc5Fau7TZnS3ZikQicdRGneZi6DCZdm2u9Pw3G
bJA3W22NFAGjP9RJhLC6InjnTwG5x/JKT4toeMEaEYQUBtM0Q0X92PWTo6s36Zgu
peTJIH+/ejD0ZAG6w1gn0PDwMhwWMMSzrzOBUtq1u9YzO6CFEIfc3kd74JeWz1g7
I6a0FVBvezOOJmQLnmc/ccowbdwSK9HDkmRhc96wMOJsgaVoTX5eKi3+VLPRAuUm
phySsYinuACD+vVHY49fNVqNAt4DYK4jo178wJtIRzlpDAZ2gpe3C7RhK+KrpUAt
pA6nLhjycOJMBjIzEBZp3oI1Phqd9+zH0x6WZU0b8KASQrS7QIAx3lSE+YURwTaS
OAAvxUsEg9i22+r+ZGLNVMWwikgitihlNFdR2z+Tr+Bf4q8uzwg+/hR+2dcxbUkp
XD2kYpq393syAnUuwq4rpw+yMr+kDE89VJBJTTLZu2B89ewHDefAOYQSaNcXiWnj
GCVm5Q6Z7zO7/Vl5dYYNuE1xT0MYvpD5mI3etTbDny9lIRnPzagu38NJtZhKzWLK
agXLVfVRBO284xIUTXuCg9PGG/QFJ65MxwdeNBQZxfuZtkSFpvxuveEViSzcVHQB
3z+G4mZHY2pNBvOgUN0KtjY5FRBMuH/hMLaW8+fmWOGZBDh/5ypfAzmNi7WHT5+K
1eZXYg7iITCpO0eCAybqgHUzWmVQVbRzwuxXAToqlgu4bZHkEVMmQezJlkiXL9pL
5ExNeQ5ShMV5x7gxUm6R64+BMHe4JwAzYq62CQ0NeeeWLjBNgecw9Tgge/6Xy4cc
NTva6yLztsVEElx4QZOgHJiaoY4HAYwxcJn0ca4iVPqYlgEj1WjvMrEy/jDsDy+2
kvFGIqpjWDHr4nLz3FXrt9rG4OoCArVt+mzC08LdXtiW5UfqXw/eT/JWedjfCZuD
XlzK5VDFMjPZOwG85cpapLuHuLQCuH7mpAs1EdathIs+YksFJ2MUuxyD8pWDOG70
FbXbhjLEtQDY9f2/CcwyLREXXI+/wrXsM0IweO06K6NTDAorFHPAZ/PDUUx+9w8d
Lv3BimAhgqcWrdYSXAoUxGCnomuWz10II6yK+sjvVsJEhJCJSKTVjFz0zvVW5X0b
unUkl3li8Plw2OAzCCJ+KfVjdjWuqxKN2BwldgzjEBFBM75q0DDPrm5F1YziRn/E
2ZEnHOFSQr5UZ5FIGnTbQbFXtjP9Qtv3C7iIXEpaUGmkrL25sB2Jj8JNSJp7weB/
b271lLJvr52vBJKlftHDLX4p0GuE2uS8g57/Cvh0rtVtAjEWGmEdyHuZLeOqF/KJ
qVHmTvyYY5CUVEsxkNTpJezdHW+z9YnPxGsbC1t09QY6Rz9vwdmtioLhHKfErvaa
3GoFvQhBylsgc3y8gEbl63vu9YtQ7exGcCB8JSgmnCuszS+HS0OyDQmmJRho0XfK
FMsN7oWneCWjDQJpA3CfLTfW2F6QD4nv7joJufnVvztxV54iUGRdb/+fmAD8ihE8
Xm7Vpf+GkI2dOg4SX90ja2QxQRjpoChguH/JgdUKS5ASH7rLyha9EkAEpL8MfHhw
CPDqHg3TSZ2PQFULMRZPHnNPu1nOZ4EEKRIgc7Ge8D+xOJA0oRoG3uh8lyj4Twba
EmqEtmZZpQBACzMDBb9bKtK8wkaGHvOW0+jxL/VShloXU7zXRI0x6365znyaLh53
xGZVRGaK8NOVCYTqGafH9GGztA8S3DTtIqbVl06dt6hDFGACOM4jK8TUgXYRySRe
S9Js6QmErlLju2QywIXDn3f6DfApp5Tdw/CoTN7wayrTnSGA0xCQSMwsPVWzCH8m
gqZ7SQ9zcdW+ztUtW6V39nuhhDPEKDI1IdHxZHt4hI3w3PvUjn+sG1rQFI/+AnRt
TxB3+pvHNOX4qCnmxef+28p1FYdV0W/m3yPJoWIpfYB8cElbgOyDGfk8HYoE62To
eLL+LnjJ3tn/LxM0pkO+u6oH086RkGGotD2SVV6Idil6mWVoSRx20Euh15uzROKq
UeZ+fzQ35CpXEdKRXFesij9nfpx09p77m7zR54hBD/m4q3RuYs30mqi2uUt8S2fU
vKLEaYbSMEWJF6OhO8k2mEtmF+R+w5pc+UNkOZ4n9StYWUZj1PGg7TyKwwJj9pi5
/G+PS4e3+ks7iT4q3BQHGjxbNlrmryQjPMV5aFkZhtUYLG81rdg+Xjbd/zlMbEhg
bEG87iSzAuD3Z9LNMvSg6ib9PDNtQNpgHpRrnyrGUs1E1vZ8983nnfm9d0NWj20o
MLJpLSu+OIBSFFYdVjkGFzlxWnr1AmpFCIgEHYhGfLOduBNW4akRPZ5PI9iY63kE
xkYaw1Y0v8WvW76sHP5D6YfiU6Xhb0QDi6O5JzmncqSR49BS8XE+fhpkZWJWVwx/
F4yvXDEYV8HKze0nAbtslvVQfte1Ky5HI2L2+9KjxL6qHJx6IZBeAdZWE1w5oFsQ
VsQXU96HtJ/EI6zfrAb2BxMLPsy8Egofmv7PIYYX5eWNVTggQtEa9aSf+3yLfRHi
6Fy9QidLzAtwirwoGTeWB527QZA4ougX2hGI6iDBAb4tE5kNTqfRBjG9M30935B7
zxSwJYxSUwppqlLYnlxua9lsRit0jDue/JuY3r9D+BHQyNRbST9D/lffVzVAGe0k
EG6/O5NpKjV3/v3tNMjTWOZDjLYXoM+1jsEiHr6dNHpewAB1MyJjjELqGPlcezzZ
yamYi2og4KACEOb9WNWRUu9ouRI5T/CBqZelaUOGh2bhjMi797hGU6+eWS+iD6qL
wLkPrzJ63QwRIsNZc4oTsIFDS3cCM56unGVYR1JFCO7ZbqQD7bahJKcNw9FkRQdA
hoRBBb5XoBNeOXEnUybeJKjQ8VsPCPX6aSCb7FnvNbxUpIIfwRgdJj1+OMkYBs/J
UlE1qBtUN1cuRv6hM3eXGmI/+QS+LfLk0/KBvvUzxfk287NonY5d5u8oRUctOB/2
FqMg54NRRTeZ9qPgOBE14Zczu/Zm4TV8VCW6a/Bs/EZjezJK2qNe5OBM5jk/Nv8D
/M/ITL1IsPaeJrxVwizuVxcwHErmIx4ArAi+shTNwOAEg24Oaek9q06RluOxX3ar
E4Rt2E61yVI/RhKVv2ckDmDUrDYTT5Gt9TfJrQcJTul1g3zAYf0DemxLI2gxtyX+
U4AjqhUk6dkfQD3ARrZzJRnEb0bUCySu9OI0k2GLnOeB0zrz01DMFMohSum0RJup
JkKAsHc7dL3oFrxGKw0A16+tqL0SMAhFWaT3QGO/WR74Kndf6EaYMxaje9l8UVkh
GE8XNqjXtAqrqO6Fr5V9KulPNCa/wArc0amVMNp7BdegxHM1NUVG9yJLGQ28Bcjs
GPJ2LmxxIz9iwRcNguR9CZtIRjOfEsRq9bIqOteKYbW8mT7v7YfTd8GAJkTwNo2S
eNCszCOE7haCywPh2RurwllwGc9FxDoxOkPYwJfvib6PPW7A5djKjVVwcqV2BrUI
efiRS4QHoGS3TJxIFtkA65iKNEgbJuV/WZ9Xc0zjvSYtRvbsD+oqnDsU8IJl8Gxe
T+9GuLczhJ+CclkuXC0sCQf/+v4oI3lR9FZNthOKNcQAKcjGrtVtaLVYTNrUiSmt
yi4dxDny/lr6pPvs5j7WpmwgeIa6WSfAaQdxlaLGyYUEDgtg+EWg+IsumqMJE2dP
U1JCIJW7yrj+B6rFqUCkoVWSwoHXqMGlIo42+SLj7urSpDEMMnWoqBMQWSROgmwH
koTeqMKaQASQegX/fqwL67r4R8vE2njib0SMY35VeAY0/wqh0r3SG9XQfSMj6XTJ
m1U1Ukflyqa4N53XmtbJuNsDL8zwTTuqASdCBLO/Gau6tV3Sha4BlX3vRfdqCVuD
cOSG6aPMklqPSTF/UXzNrQgKOQA8sIWTa8DLGQ3AVTT5owb43QIkCW9gSHvJzQqw
0zVxXUYDmJK6nJwiALdD9d3Xgy3IHFAamY8VbYesRZIbJxzUR/4FpdnjfIhX8Wea
JmDPUSGcvsuK9ouU4SXCXtX2pcpj0j04uDg2d3NV0iDxKku1diptuIgwbtNVeY+D
HAKVkGergoQmLAXmgfDpD6uTbL26Xjm6PUwaqlGLHSAY8gTKwuRklpNQZCzE0x+y
0mUOrh/Kcd/CTI/xWQnvHbI6wA+UDq5AbC2z9oPRiX5i9Gb6wag9x/qZdBTIYE+l
0KmErSRhQd4JymQMwSbycsaeUVqUQ39D58z5JHKOZkXoTk4dLR/O/PWvLKggdyIi
9cl+Gn8NFMx5/wS7CRqcfVcMdZZk/XQkyT65lbKKB5M5xg5a4VEs9V1tHTj7SILW
hzQNa2SqLOIeQcCRT8VQwmVACDe64J3XPeByNgyNhOcajhjlFYl9TIU4Raqbmf0D
2Hy0ZpzwfzbvUemKAbqdLhdz8KA1MCLU5bOgLqk3mF5uy9y03lAuDN/nlY+sCc+K
iTaXYdazkgSu4bDDhYPuhFXrYJDifD3Kt7Q3WrXuF5Jy/DkWWCoyUw04n11CcK77
0vPV+UwFMAdMNiqdOdKOQXumB4T+vuydi/jk0OmgJdaEX22UilCLmIBRpTaBPicg
Zgxlbhwr43myCBZp3paVdYnn31aC5/fojuyJ6yAyQJwCPSR6YHv/Icey4lA08wuo
QcwryiEbnZdY89z1u2a/ygAsBZoa8LPnGXF6P1sTrFUYsJQeSt/P1tX68jVOGY6o
8lTit/Zs39/yjPOHVojQ6KqWkXnWJLvj7dVG6PqOFzjrIQ04vHMKPDXJIZv7R59w
yw+/dGMgYwphr5wxlWcEQHWySWINR3OI8i2fYPbhrk8YkYjzsTVbLSiCCqWlnsb2
rDe9I6cnEK28jSsYZmMoPbhQxGNgH+xJTEedwnhtj/nW6TY7fObp8ZxAUVisVqnt
Lw6U84+QBen2wBmEwPnz4mQJv4SQRobViz25xBzwuCs7sVcxERsOYDYQDjcp4HaQ
tHIcVh59oQmBjMtRM/Y6PEkngAnaUuXuVVQUf+aaZPfMLOvHZP7zGj8/HQAc0bA6
azb4ma5aQurg4uzXWbBfUgeG+DZ6IqbWO6Y3YX9Tq8sE5qtuCPtEToolxV9oUq8m
XN9oyvfXrNTW2969CtmYvhR9pn27zotspQqxnNzv5ZlMbYy1G9Q8NzgVmdh+3Rsv
VkJTz95RYrbSA1/b1iNKCZOiOqImHfOtQwWDoRq65nwc6zp/cb8P0I2EKieHUwz/
Mzf7UcMZ0C1Zkx4rUZ2Irnk7iPVWUHO/6u016zlY5pG/10tO7KXe72CvUhmj64Mq
cZmwvsO1dO09p8qtZwNovQF6Pr9+BH4r3Zu3X9TQoIegDUNh+ktpP6vooPRrZ65N
fn1ZApoZh6hJj8279MQYcyNahfjgR2XtX77KzAyz3icQzCXaRyzSnX2PeCt/uzQd
S1nIYfZ9i/LBIMIjqk1R5sWoeD7uhWqE8F4zSSkwTkZGV4tWhqX71K8xAB1fPl7j
yN/MopoxUIM/1R0chmwXFPVbf6skLcBBLCsmtd9b+8tAR6kV4OVXeSQSH96jXU1H
7KIrBiTUn+5PrvpbdEqddWpYq05lEQ6yxnUlA5HfmejE74BDng7m7LGDzLrp/io3
0U19tU9i/GCoT6vj5HKsw4BJvBfg+xLmJ7hcSMifzq0ChUtdFd6ecOmrZdoDf/bH
5wk3kF8vJBqIivOahSTdCGv9Nhk7NpN/vhBUMc/TdUlU/c5Yh6lgNe2rHOpAav9x
FbQe6ryJ2quk1hPs2Ud77skjNiwTbJeYf+fVDRDlfwhjLQaDZw3n52JNqJcV2AYr
gV5UtREVFhh4t4XCDpCdTAksboRLvLdYpWD+757fR3lQSy5MkhbXkUnyipjDBxdv
ST48wpv/4EP2WYT8A8XufbE4/LeDkxlSoZ2uPzVNroeiDpxqsQ2OhKsHjOoNj/bf
xJvUZgPFBoHdoZ5dJmMomapW/vYkFRsPVCmn1zycZqi7ti7Ms1LiWKq4iZ1D0dZ8
hOhcrJqWGZbS05/mduk+kBgMsfgCR+MdGOm4XfSydwNnbtu7zn3umNSAtY0dtGtN
OLETYTba+ZaMZItLucQRQbrAoWKqVf1vKlOUAedbeVP2zvgx1dbdrfSyDkze5Wo/
d/XZAfM+OHmSG5265xs4xp7/0GDWWjOoTQJ8W/F5whSTuZY96bdfEbDZkrd4Gwa9
XouceyPpRv1G2RV5osr96vVVUNkoBIpyiE/7CfZruQc7jbKKlN2+3Zig5IhJiw93
MW61ILZYLUdmU9JapcOh+rcMJIDsdLbgzUxOYTIlYBwQYrpxzdQSkTOO0YgrySGg
6zCiOdoj5qagbyqnnYylD6tGj9OIQCDhmYDjiTd/dFMekOrUmsGVBP5Ofrll4GZK
2HNm9R9ZK0GzJ+MEfXuB61MEBs/ClfFtgTK5HOAdGmUl8+LXc/TSUpInUWd8PyQO
yBwHnSkdI957GKJFM51SBapYKjOnKSjYixUfHK0ejNeBqvTHeMhlzEVgA5EamlYO
HZxCMCdI69BbqfeuGwQ6MC8vv4bbwIWL4H92bhvN4gylPh2kiawZwfRIdop1g+5h
A6Pi5/dObDe1ojdqCpx1BU7RUGLYpgHLCN4xgy6LBC9BHB1J54KZ1Hrfhxt/wbTa
ABO+qWawXq5uddcgNMgn+DiOSh7bsjyRdPfIMHDE9Mrpb0z97GlMZoKGLl64SaRK
VCCJkBPM13QhO1WrlrqQ5em927IyrD/H6cqyd9/7DsfFKsLmh3cEBJ3JfcleP2TF
EH4zSdCJOmRNFxf8c08D46Wlq11HSCgU5UTowR4re7KrZzF2Mku+bXBgOtRJZtK9
1PAk11PT+meg+UidldC0+AXoLA8F93qt1/PYRuhTlQq0V0ATWpvefjrH6KsHQXxf
XaZcpiEX9RVTJ5uix9wjDeINlxsqbBADX2t2oTS+nVVaNgYUPQuR2T+TOTGV2xC+
BDsmveESg3AUHtV9U1f4ww7ltr72lWXN4YPb3utTDPtqFhWpKzEiieb+ZG8iJ9AS
vLWC44HHjWHE4mVff+kIrmNkUz7jFs6MrYTSeluTvkkTFgHzmB0K3uDYInwWvzMF
IDcQZOaMQEIDaDQlRIxpF0Oo5nu1D6BaRvfFnxOZ3snrIyuNbetBxaGvRbHMQTEm
GAkdiNbYqFpGb6GZZxk/Qs87XfhASTGxjYmcl4D1OEfdSu58ttT2r4jKEGyra+5v
lu+3lp/z4q28F6gs/oTtsmWg+fB9BToCP6CCWmPvfbiFgKgIPWhigrvL1aH84pY4
+UuDZ55orThaNm4ifkopCM9K480lPAM1u8CHjZMjEqXoQJJQ8DGADj3a00Dna4sV
ab00U2sgsjXAjSr8o3YLj95OtWsgoV1KS7JOhiT313Fvg0f6qdoqD8Xn0MIyx6Io
V2s4y7e9lD6I71oWLlUQ712ZtfTcGtxzftJcH9eAosPl21Z9pYmt05ViLWetxjji
THHyNcU87v7oRC3rQeSWL7lmrAXDIXrG7RIgkrFpnGt3WPdZP9FXRr5WpeVBJH2j
Q0zGwwNhYeWQ8FG6sQ804ZUhyxcRlTGu5r6PpDKuDzJmszB6aF3LU5Wz7YbucmBG
1jusb29pSCdswI2pC1p8c/1TO/1jBZNjOt7J2NH6ql6VNlziOAd8iWnsL9ajYlTn
fNMk9uevjUMofhM/etQM4t3sQ8YxI/H/KKEDjNjqDVjhaKuCHOMRaTAdCwZHUCW3
zdYKjMJZw6jm8s4nT2cCLS0eShxYlTp17Uf43+VYTTYQIjSItHX5Zy7ScEKWm2YU
+EjI1Ih0xNUdeLsu3tblrTiAzZ2QVRJDypylOkEijMdg1HroeJzH3ObAmii0ygAI
SllDkK6qAyjFH/2M2mTUHDLH7RWR9AKA+aUjPQKiCb4znZ0AngURzgBIJP2hBahS
pOiG6PifGeAruGODSAnWVyft7ussOI2SBKPUqkE4CvSgZ3LRka1pR/vMQPorf4bq
Gj8WcZdQs2WuRUYO0WKriSDRP7Gqh5jIrTS+TXVQQsq2TKWCGe1tPESQyplsYOCT
Ida3+lJ4N4NHW/FM7dCy+lv12sYTSLyY94zHXCQ6HLPmpfPB75ow8wA/hqRcEA2K
EXImpI1ujwK5vLp/JkMUPdjRV5h8rletyZ4foj1mEPoeHAMArrkLi5oqBEK/Xdsu
inHIHHpucUf7mu2osKB1Zq80hu3V+wF7CzmDuEGuLtlzuyPS7pn459GhomAk1JZc
zefWEpBpsV9wwfkcpFro5hUUQT8GEHTM9XI2X7qK8z7DHJekJcCtQnz2hTK2Ez+9
YCqMJd8ZvCmhONTn84RfWen/eOHqvfZwbdHhrNOdB7aY02pvdWkbjpVoyCIDx5Aj
bsl1CdPW9Pj+SZDRVVglcbfSYqvevqa4fKfIMwOrasi6kMeZYN8U973aDM7P81nO
2AQ6iUXrqZ9HEwcWhOX9/CB1eC5Z/AqWnFp74z381fcbOCbWgH8Sd4FW+9Yj9DHy
UuwrAxv4qLEcUxY2LOfAoAikmeiBep3DJAQUawPZNw3KCIodxIs79zRmy4SoTtA8
EHC50y3jASQ3PLhrpHuKKFiFE2lx8DqdqxKrcq82vG7S209FGzG57ydncv9A+2tK
Q3KTUj8FrQPqJHrICrW4ryLNW7tG/fd0Hw4CunMmstitotguXppHS3Ma9qqoMpIv
fgsQWmlNJOPCnsILOwV70P9AAcml6ILEWBSUxRUGpYceZ6rdwH5lABjMX2cuzDP8
L81swcClRrnxuAuArZEV4fsysXSKLKkswL3zIbRIjMjBDtjCULU+Tsb3nxJCFxky
tyOxOhb77QhppSDbeK4PSgZbatM4W6jjR+sHW/gjIASvD2toSetlQQ/o7wY2f9Ed
3PLYdrkJpsz5/aaLu+fDPlup3btIRjrkFBQiGLCD66x/jo4hNuC8N0BEFfiGYUKQ
sqA+49z/6XEp8im7gozF0pzGRROEhF6KGNd6ndUdO07Uf2Hiux54v/joKi2pu7pj
S5nx6FKCjKZVAMR4PosBisurdOCic9cGsulaOD0841ttL9XCSls825dQ4J6gUCOZ
Al82CQsq7BwTFu2o5RaB7ESwg0LSWkxM/Yi0nVpctEdNm9WdIAknbB8jAcIktMnN
aI4uUL/e0/r462jUJqGuO2zMfqpHXHQr/KHEfFL58X4LxbdHqXbpgF9Oj04YfT2I
LP2n7e2uWPMi01EykhCHuMt8aZZaJY7UiAN/4zUqXoXWqHLWfy7taDbTjrA6bDUL
pSoMOBa8vV5SeQVEJN1RNKh+55zX0Pa2m5g5VCBVTtNODy00EO9M6quLxcFAOErf
3TomkfVcpzbB77suRFhczLDIVimfaU7YSFVCl4RU1XeI7j6jKps5jHT1FKI+tZxB
X9m0S4Ie7E0ZY6e0auH1nun/GNjeMrgBs4Vvm4/yIsCvQqajrx2RMzvkbIouj4sX
eBJHLn+2T4e5mwjwYG9xQeWlq+Q1YDMi2ULigW10i1RDv0iyx1yfps/yWGtLfWoW
fVy3vByKOVfcDDOCztlF2jXxsflze4QsophEW/BbdiiAP1IfFNyANc9R7649NSJu
n78qXKTJsob1TDTqpk3XepmNnwg6d+VGohS/TZ988D7x74gAASXbNQS5U4tS9P/a
qycugy4CO6DnsmuqSfSmxy2kRHrylTwgDV9ueaQOBfCcejRldO5qqpo/B1imeNyu
Tzz8HTLgOuJhxAtZP5HTARyJLH3EEdOREIXRb8NsX/tIQk8B2A2DsbTd7XpsIbKH
HTpoAJYyoGOKT9gq6acs/+5kpOQuK/qPYx9dkrTjpN2pwrYQmyc5WdIkrP3hKKgq
owP54YpXXpuWqPXk2ca5mHM7pAfci6Lw0Vm7SNrOaYKq7HwpByGIbnlZcoww5Scv
C2CGUhqiShZbYVv0lIN4IjSUEthbPFUZ2slR9pUz052TsJ6at18fSo2aCf0kjcSl
4ULSSWtKwKbOCUtZw/I2WyY6/lq8z/7z4L77T+HXoOscwS7qu97ZNM4ggds+6kE4
K6u72zOmwUudwagO/8i1NhTYYr7rj1EyTwsoHZnVpfviErP8NQ3MJNkH9FIDTzLo
e1I5+H5Uw9Ba6IMz/95PZVXqiTY7dsWwuGDfVsnRo89urb3FQgdAT+NKLoFYDu+n
KbWSjnDSON2IGhNuP7hKs0rK2xihAQoKNKYekwTvbGqQsth8ziZnO4doWs9wu/La
yZs4hEutWgn6tlJ6pfGp/PE8zwSp4Okeiro84jEs/L+PWgUf6mLNOkCs7IJxe/c4
53KsSZQFKYWW0iDrxMAds/B1x4kfT6ZRdWTpVmiPUG4KYw9cPVWGZtDRjnBdPV37
swwKEthhPdExAO83vbhft3AM16dXO6J+rVrfoW6EeYB5EWLRVzy/8NQyu4GiEzt7
TOyhLfQo54Q2u2GSQQWz78ccF147USfg8FXii8eV5R9Cg7uFZ+NiJzURK3ig3MPS
OPb0XeQ6qKruVy5/q3G1Pdc+0ivtlx3ocDrPpcDbKXSQT8AlJSOJK6xtuKzuy9Ur
UBg38C7UsFrX6hSsmJGPzijPF2x+InFkrN3Z4EZ/lXzke++0MRR+mw/Q/MvzAxoA
VAAb0GhZ+dt8hMRzDfd2Z5XJAjzNHlQdCDuNN7i59ACn8e3HnMJZuNFu+YdXtGkl
70P7zTy8xuPm24XrfIbGfXxewHhrJyzyyxJSoyo3wmoVrn8IEocRYKumJNRtwu9q
YojwdS3RZ8mT4MsROWVIj3/gcxFWzoyPaHe4azrmFlbURgSF7AHkSst4aA/iR0z8
jnt2A20ndO4h8XuTQIguj/rDzXG4HU+h3gpdGqeadV1sl960cOq/YJv8GiQdwhUW
ATtIwT9xiZIxiEvdprp+if5Qt4RiauhZgTFIWbs1vDWT/++D82x5G2vICerLE5z+
OFW02bgP0zMRLytFC/0+eUy5OSGn1qt2aVh2Ep/Ql6jysgSodwbYEE4zmyGijklK
GMIbRH960ssKMD0L1NbFJOSPvNjCk3xwxSG8xqxLhmDSS5UduGQF/IAI01cBgemd
DeiO3q3y2+EmQLkKy2rQJnsvgqTriQrXI3EpMwFIWXca/KmrouyemZ7wiUIDvMGI
Qi+d/D+dcvHnbPWpEbRHqKeYntoVRTOKEQXJKd1Dah/pmxqgEo1Bw7IbCb1qYIKa
Ej5MNFcfj8RHV3gwgq4sI/bLkjAs1p0SdCmCk2wCTAEFnBmMg7wzntURFttCIGY5
QFBHvTair/YX0ZVxbPuijGeaulJvqh9DksPiz19RkrdV85FssHknfjouRSUDOrmc
YcH9a26Gfr0irZ2/iB/50Houv6XhizMTB/pTXXwZIw6rOuxOxacnj9orskqRf9+6
viVkP/cqCeQ3YE3YF5mWxxxljoAfMA+ri397vuzHarP3vmHz6677aOAPvwrtc0bC
Et0G7SBWYm4wtHIWEvvXNjwOEzbNyZSvK9KfpyM0cQMjP55UGQ2C5goNotSl6ARh
ep6FQyvdWHNewKWAmu9SDkIDBzmizH3l0h0HKkIjZxn6Y15oNVggpVg8y+LSDPrB
zHUcrdCLWmG0sAKtHl0GqJtf/PTRcOYxsuprFNIz6cWl32/z78hCWSAkk53D6ugn
9wckymG7YzqZT1JZ0yPnmANTr6ZLN2DCvRj2ctODbP0NKmdbf86o1BdSQRbKL+kQ
f90wZBZ4Qi1uIEmqjzxLte1V6KnZfYDp21jfxksBi+BJRkF0VgHnOqryfH/lotUX
fRN5TFAufYcS/NWTLKORtNWMut6zVV0Tms/x85apVJkznnSaaBJ1PzVDInwm/NiD
ZWb1vGONTJGuCrRR4aBWOaZXe2IWtQ85tPdXzxXgVxoDXTzsVIfkFryZ0N1wEwg5
+auB46zMFLzbLSa9yAxQum5C6qPw0//EJLQM/GTC6lDzaXBMsTX0mk0YVpCkTiCj
wP4KIHYeNk5TCNXxrXwYheyDePsqUjKSp274tsiEaxoja4NWhkzyqmmkFOESqLVn
PXg/NdAibrly4mtg1te0V5N6zJM6wFmRH5g6Q2NOO3g0Vc+hu15e9tPDr/0sy4Um
cLnsLY6ZiPB9OQyovdQ7H1ZiRMTTp6Dru0MC5H/LEKxs4/+LSaflSm8Q9msFHYJf
tPZPlP6XyiKQlISxAhSGS1tbIurStHx4Mr34VOwSLcEYIofBGIppDNLwaXLExN6L
ZECnqJlDwdjoqEpWgY6tNzBdFqkxkkPJsO6dD2Y/aeqS9df3UpWAUjr9Ygw/mNGM
xX9WRX/VgTYhoAadohgDOGuuH/6Xe1lK2a74crbwNQGf+cWJQcm11+9Tw9h2Pk8K
wkyUtg/W67ZxH4BezFU2EW6B1OxrG5cEM8pHB0ARSkXugyNWKvNqvw0NAHzLd5hn
KgWT1h7PJnrEcvJKZ67nEcg63ScT1Rwj6zq5JqgcjaksloLQqk3zOu/ypcJ1hDGR
NQmtZWOs6n0Id3zdmYRytudOqRXINS8cXOaCBAWmPTB4PL5IM4b3rSiTwO4WkEYW
yoponL5SxEhXvD7inomRLkZSDXlId5VeSSV2cfVJdQs+yy12Rq434KTuk6sbLtA3
c1tz76Sh5mC5xdTObo3N0CrwjhXhUxI2lU0U09J2LC716U9aGEPT+BGLgigSsACp
ZpLD/4I5ZAPNqBHAfT+CsOODjqTrvaayGHC3aPubVUjQwxhNQnKkIdGJ53b+sJ/U
2OrIBmJeWgHiaMHrcpZ/vy+BkNZxAia5u4wHiVdfrx0jOVZ4FeRmI1Zw27U7F87F
oUQvqEMAOUnLlAXq+6aRfKG3Q1yrX30dpW7xnFCX9WzfxqdMWNpVGWFbrAomPxRZ
xj39ijywfa/PtgV1UtGEfsRaWEEq9lc5J8pk0AcwLzDfG8L2dhiGlji6FPQun3vn
fHJpBl72EGAGUFNGE8K64g+64Q/37HuBtMy3hs/rgLtdsg721Vxu9E5aQUEE2s1j
Cw4FAbOUVD8qvmrxdkbGxlwSkitkph4Sskb0J9qFQc3GLr4J2CVHTS8FTCuF2wLd
sc6eNwYa3AC/j4rRJx2bysSMy+enxsBKws854EnNNGgGtgZYc/AUkIvsaprRfc/P
vXF0sNl4nF1zNsCQh4wKaIVvK2HwNxWriO23BJGAkjH+vC3JrTNfsWdULyetqpwf
0CMxE+KscUiLfsNGOigUY5NUMNhiHp0wOgbf2qt+B00XVHLopebTVdENnsjN32KN
6Zw492SRr4a+kradpaT72HobYPeyrJoOfUW9F9jYuqd16S2YmmW56mEOr7ATUR71
PIS7oCvfiCgL4JB3vivqLtGWKVGqJ7NlZoGJVVxCSAWpedXlnrcEY3iT1XONJiqZ
a3lZybcvyTQmv7dKawyzNhTkvflkb6Ue/P1LKN1NOC32NKKTpctQPlB5p/xAm4Js
vUaqbkcBfxxJZnIGJcTmjMyxtcwQ8HnYL6l291pT4oTRTQVukfa2AtxUQMnz0jZI
O57lrna0HSubowNyoOdACWTcMoT6UdCx7q2Cl+1bCYIG4COvmFHwgXnrNZpl9bOi
ffW4tk4hZ726SrQSm2Sjpropferkbur4JNQWLG05MEuv/7idbUeNsSvIcTVqR75J
JG8/dyIUGmYgCqSdnT1tbKI9WG7i3QL0cWdOnf+0DayWZj23+rXKFIemvie6tgqe
FAgil26nY9HTHkp4Ax/p99pQj7k9rQrtjkH9otLYWw3ucb8VHQFdtFGU2sDeVhBQ
PGw1Ohl7MTw1vrcihy2dRvVzGALCEZmkHHpP5c8CWpiZUoQmj1+P6aMfaXnBS1Gv
R6e2DxrLRSoee4iUTB6o49V1V5itncttQO5tStYX37yQloTgLJ5OsRRqSGTL6+xU
YeNA8JPzaVClaoUHVdNto6lVCiqeENoWt1MHkmOLkkU9aMWbYONIgkdlEBa3Fcka
6nYHypUdx6xXl4y7tvfs0/9Ju9zLvgcBd1Z9F8uNVm6JpURHLr5eMlB4vtswiIzY
mKHh9by5gERPgGMUIIa7SWUQjKrChRBFDjmJD1XzuXNvlPp9CaLWMA2SjSdLm2M5
OwWBJNMj/L9d7WOZJ7/+jzn+teUlnwx05SeA4UUwSvZY8RMmza4ZGqfSp26BUn+X
+HAKec591JlEnv70OzRCX+uESvCc6PL3fctCYZShW5KBqIsrLkjp6xs9gQfjUeuc
BK3HWvbLexaUQt0RilHfOTBqL42hcPpceUSksbAwfMbugdLHmgn8GT2s5YR2j+r9
tPabl2Lfm0vhPh7gcL/zu1okoPHZF9xE7XomioAP7FUdC+P4Jp2gt0uAtU73hZr7
mtRhSMdfbd5+gndwjRM2J+pWJ9hZmYyo7kKN2SOoCwSuKciN8xiJAjf3/y+COgvF
tLh91vvCXUFV78QxNbu0Ce2iwMxCLPVOKjxX7Yz7YGsiSAwMMZA1bt5hFUMdjCLp
6MS+0KTu8h7aGGCG26CEHCkvnr6aspYxYFVT9tQcd1/7DtmS5mnQNiwqw5crCBfk
Z6fB+hx1uGsJfl+pNZYb0orhIwbO2FSJVANMV7QQpN/3W1aMHtr6F4r7EM2VdcTR
9u5fFe749yGrHP+PiQzayYXq1kV555/VmNwKA20KTPXUrlRmmn2vuMyjaiqD+ldO
QP3KoRbtlK6hj1U6ITPa5lNUjjgBuldVFfLRasrk/eoqOwUZhd5csQfAGaNp7utM
1jFCWmsaLKcPBv/diLSAQFvdPXPhrH7X1KCVZcn/Vksul91GAPAm85eEIUp1FpRP
rdG/vYIiH+doDgYgv4kJFLl7GCWs87hLERFefxfjPwrKHMTLb0g8WY/LrQnGIHBn
f8iTI+9SewkM7USLNgsWmA7tEfTb2foAwJpfzgG3X7JAQgv0JcnwUyTox9cz146e
NJqt5LJqJPsf0WB+LwNfjArcMIxpg19P+6LKHtO6UKPs/VR3fYmdLunnMvXQDQD5
xy+gI4Tg0muPCJIh4ortkazqt5GM0V24X1Y8dOnKt3ky6TZpAOQzZd+CBn7vyLYn
wPWQsnX9D8uMXpWHWO0RmFZmtbnRbmMK4VkLxPB6SmOwjt8phvcNUlApx6fn0j1G
h4IzhXfv9CPalUaDopc0HvVxdagDfRWfDT1lfMWLNzSMpUx9D+2D+nlDR+3SF6m6
cCh332/Pu+Dy1R/MUYvCtNS6nH28Rdy6fAc29NGUZbIToZpunD9FMZHg2gdlWJJk
2nVON7rAbnm8sskZl78TZhjPTBAGJFp/T+l3S3yB1VS0czrUoF5ZFVO82YFNmlXs
Z1PPbfrX9FwkUc9y7mtTgDFnMq0UASzLdiKJkrnlHQEOGEFopPFqKO4+ffsTh0y+
KX7qI2j6EG5lywiJCECOQcRT69ow2jLANHXjmz/pfx9VVZ7oYqo6CiPRl5hT2dKC
BhUGzQ7r0hHuVO4pf266XQyq/Bz83eI+w1ktvYiJV8OoEGgADLjbFTcBCKMBB0Rk
g/AbWcp/QOX8IwuIFrM3HqI/xVZJ653/ymnpOPnTV8r58ANq7T+TzuP92TS2zJNU
wNyugInNoHddnpoFcLc5Q0LsPm35iunqglNmWWZetAi+3H3CB0unSHhOwZVS5tcy
ZKBbOsXOfV9QE8Z6zROy+XXOCFrwbDQ2vbVgqY+M+fdmNPjwmckADq5GpCGR5emX
oW0HY7cnPVa1ES6C0uf+7sdfJYZoqEdnKWem+oHaXgfI2wnRU0dsn0a47eTGqZz4
7IwXV01fuz8usfTO1Go3ssP+Vo2fd69bZMNBXRf+EUYANwOggikMJIXiOdJTvocl
KBEz0wqx7WNpZUimpR1fn6HsYnJPIhNBGBhs919Hzo7M4xNMSSCffCZ0UH5QPsP1
x7dVQhs7Rl2Htu6xS9M+SA6bVjgSqhkFpOv4O0QC7ojHZFjgIg2KmSvQEzili5m9
R1lVJb/QxcjBeG2In6VIqTySXkp9c8CxfbLUuyi2+vDpKEif0eP6eJIfu/KbjXly
fzGQhrVLvOI9Raf6P9lcvgNzhVXgTm/ehdQU6p6vJtrz10uXsozat0zJxLMF0C+d
dgnXZycag35GDEFRFyk2U4pxnbIiQuEoxzDmpOd5rwquWSdQAKkrLVvFyOwimCBM
i4aEdxp1suXKFJp1fumi3bp+8udvm51wDoiuQ8DCI5LiKPSsEd+z+WwLAy+QR73i
uyivG7mBMZOGr3N3cTIwb8nH/Qq8mGwhBo7c9XNSMVpWUogQW+0NmNcl7sUKdS2d
cd/w0xYsyOci2gOmFirZyuCtg9WVb1o8Roz2unbprUUcouBWdyZ0HhPu1Wb5ppd9
GnSPM62x+sszHiunOwBdu6a7PkbTAQHBjLOwh0fYhf+OIOuysUDc+zfHULvvnx6k
Kl/mYEH3SyfOuEvu84kExnYFVXUWN3iQb/EZQqW2JXKCHV6N90XPyuD1QcdZ370h
9/5BDXFoeUW1qLartM6tXiYJ+6ZGG5umUV4NR1CcWE4IwzaABTom3cSazlO2Ad4t
07UX+RZDQH7LRl4NQEacvGaqUcb93a+kDwuKHxzFr/EYEL/FQlnpY5hwv0GZN2gR
DpEM5rWes8cpKE843MTpmnUIrzeH5NWrHUh8lm6vY5OdXLkB7oDR15jPHOdeWmtr
sesn+yrK8M0oOJYQOsYL269EBnBXmJWsQ5uC7ShZAjKkIK/xRR5d7cqx/PJA/evT
kwGlP3nBAsROEMT7xuOdVuG6TmmZcz+NM65nbp4EcEvgKlneffMYYROrmCitoLzF
ElsvaqzStK+eLeT89rnIXfI+Z63uOhARxv2rax93MykL6ncIHVNnypWi/NOuiej2
IlwQyAIq7jI0yitJpF6bB5VWJpTAWrrKbA8v0UegYJwfton6EOWRcHYhH/rM7vOu
R/twZbjEHST8tokzGIwAC8x9rafxcZXw8oFHRG0OT3R2SSiFhjM9evWisPcEZc0T
WDZ71JusNEutbkmHb6lkb8/i/CM4ti40v3fwTzVtHE/D4WsS1qX3QQJEdgeD5EX4
NAFEXHyw/RGwjEGg0iWdB3mGaEo72X1Kzi6KhyHiUHXteajac3B7kZE+5dCDGLr6
vzYCMkAwssc0Mp2G/ab28f4auvnKmQXrUOBhMOkDQBw9KR0XHDbkyNjOQL7By94E
VxWGrd++ruimsIWLpDqlJ79KDG7f1t3LVULWQdt8UtOSpV9evqFsGQn8Mk8S+H8I
qKhpWIgCKnDUDxufOiqxSCDq+/mp23vFFhldQzNQZ+U5Kv5yPjMFf/z9gKUM2v8/
hfYkBGWoIA0JZXK/yUJMOrdH/y7tYOJXJNaTl3nuX9z7c8OPdtwoHJYLWej7xXC4
UFzptS4zt9GpQhkr/o1KuhNrgGaFyzw4aU+Rn2EVYuj/TbE37d+ymPCmaSJIoruk
1Vbhir74gxlYznpIJ+Z+/fcjpQdM4luV3jDOp4TPbbs++M7lPg1un4MrMS8gMk53
TPXum2f9dIvZKd+JvLvb8/MZZPz8LGKERqHOMGQm2tdPL96DyNNx6S/tCZC6jUk6
eSbS95/8OEOsCptlX2GzhU0XZvKrxz0uM4X80iWxhWO6e8lUQBwFs5cLP4ES/14t
5fHakt0JcCacTqiwDrruY30V3dbuaGB8Bw9D+FJKUW7kXpFdlooJskM2gfk1FU/N
HNqslEQ9oWaHp62vSPArC+5nTNT4w/6YKdHxFHDTxW+yqP/y1082X0AKV+wiq/Mt
y8OAcow/J4dMSGa1WgqSYH/Kgx6QhKTri6cdldP/52PF+EI4wRgKaMdZJZRuAtF4
BZwnlHrE3e1g0AKsIwObJquDaFHTnGIoxD3YIFlW9D446S6eKsiGQkUFB0bqKDm3
AZJFCH+eEduhfNDlh+kNEYo909XFoiftlY1KeCEamwBqFPzt93K0wzHV1qSB4TYk
tfD8xzV7UdUFORptXDCf+CMPqBv9qlFgN+qD9B0L5VaueOD+1URJ6R6+0foLfPbB
7LmITMLzqc80OXPv/Db+ZO2W6dR73B2LM+LZbedBdEUTFMNpdSdAZiBHtmNp2QQH
k2FfkulzYZ3463QltIksbHqZtEWnJ3s/4tj4Vh0V3qZaLUMTAZQ5+NC4j9Kki0l7
9XK+LV+vc//YnPWWbEhrp9XE5eO0oAnnF+7rEvfvYxJXmtfoUtlKd3WbBI4yqGaa
yxhhFyOgoxGAQqH3JVKk1AjNivstVn3M/WtOZ+ozKtMntmz/b6WBZt7uF5Y9MsIX
nYUxrSZz9lpUteWg16wa9xIZMMWkIrJ94NWUDVST39SzQuE9xCbcG648jljGnBC5
7rDf1cB0Tnj7tRmWcjqK1GnH4g/vBlpCY1PRwKfnD5gm6W1karKq75GUkC/LyXb7
ozC+p3J1iOxPYpIcPo0E9ZsFUYxeCteXzQ8PhSnS89fh9ZqrJp3jZlWFI7gpezhw
qTr5CsgviG4oJ6Z560fk0o8PrXUR22xnBfanGs4AsaZQRRj+yi2SnCo51ktOplY9
R/APv9y/sKKzES9Q/fm6X03B735JQrUIrW71wrX1tyMx/1US+tDx0BC1ZJtYQghQ
OGj3l7z57W6Cei9HASAZWgWamliV8GLtKVcv4+DgsMr+Y8Dgn+aOoy8Wmb72RzLi
txbnAdpwdS3vaJlIY6XwS1RhUuQ7MwRm1zahJE1EevECTC8p0sGSp4DTYZyv9ZtX
+rQ7LNbvjA/X/dJh/jByU7jC9kUqB++xsVxWoJx8Rk8TliBP3YHpjqDpbXc/v7Xn
fkfnPQi1Lzo/ReL1txwodO73SSi5icKLFJWN8mjwZkIcLkHQ0U+Gmkc+8b4hi+kw
5eDUpIaGQ2gJb/WQm+b1mowtlHsRHETwxFTvWNE7w9S/Nmyi7mRDBnbuVcOKNMvY
lDyq04EIdjZkPuS8TGMBAbertVs9LRaP2VjG4JjaTzLDbnR0jytwIRPjIXT1AkUZ
qXzK5W0tcHes9K7C6HdKWC0UY0esZvBigKhv/To7qgzpQaqTUVROMh69qc7ULPNv
+FSpFv0g1qvgHAlHNEPZ8kLiDeqk+xUlIxjHftQUjv852C51tk7viSx3A6jW0jLw
DpZC8XxikwzWvM4VkX2xlT31L/7EpD70L+AOa8qutAc2Jcbgl+xoBFmMcaFtq2fF
n+CusAWr/KQr49g5c9RlhHwvKP1TQLowYt7ZWHrtrzFS21YC6NmWV2LKcHH1q3I4
crviy5YOZs3iLd+GGInVznhf+IZCvjsvuuTY0BxatRloPf7YKCntCCrCS6hxKh+b
xV+VqLa8euuAw5rku3oAbIem6O8uK6w+w43HGCkwFjqrRf4JcmzpIzTAlvwEhqgo
eKGS4b4Ret7QeB1ro+ffBQdgPr62u1PFH0R/F85HbuxQIi/+lPRuJxx0jCcLVGxF
PzqvHZShgieSgQQ+l+2ozx9j6iD6v84HhCbY33F8IWnuWOfsCzXz16cH9mwQzpHV
zTVTt/OXE3dr6gwc6sELGqENg55D5Xy9EHznxREZLwQbxil34+k8RC+wk03T1XKb
7AwhS67ucmEGkY8tOgDtbdEv/beB3SoNlfdwBJS/l4bY1UUjPYZs429uH0L83JIE
3FPrvKHnw592opUrSxWkBpyREZ8rhOb8TAXI16SMXLF8AA5VVxUixTotVERZ1paE
EPS56zZ7gK4be2q85qzFjRCVF+RTvlX5TzhOCetA75+4vumhkCznQdUrT+cF2Z8q
gbaWD77KDfhJeayAro/ZiXmqDiU3aq2WEuNFm5mhhPhmjDse8cCug6dTyjCdVUPe
5PW0tyBWLqCW4Y6w8GY0VizMx4u1eQHnSRuI+oAKaV/PFVeJzMTR/B13znoq6FG5
ub4MXFSiezjxWLxD7J26NvV9TXqxVsVoaXGUYfhKfvyfUkT1XaJZDsueDwUOT6Ky
fVbgOAgltSytTT6Uv6AnMVMG8RICsBo8Qs3BOCazx1MPaTxwR4TQGkB44lONwzhE
rQxXMZEJtojP8jrcyVHlfLQ6Ekwz/coRrhJexKytLkKcnbT0jFrr7LftYDvJZV2N
x96UjTfPSwsgtKJ7TYRSSbjM4jSnvF4IMnECOttLfs3shsCK1fygNwYMMhe6L20a
MCs521oJyn+al+F8G4wRiMkNkesxvAhK8NSFNBao014D2yoqoJ+SxVeO6YGW9JXR
Ol6RrKFkYwnPKpOClxjnWtUnn2QdyEujYVHDVrfqZE1EGDrPo/fa5o3yqESlJfsK
D3I0uhFfQZUP2kfUJjJBtr97vAWUxyj+1L8b4ntP5u9bhCX1TFIwE1z+dMxuyYx+
ecsB9uE6Z/vjPFt1e//Jy89NOnd1r36RTn+NDlLVmVDX2/t+KVIXrt0kfV35LBkp
5bCjYf4d5DuGwo0HwSy0QbOWmRkcR4jaG9tiWVfQxJ5/65NFTcsJv1mFxvm8lhY/
aeZI5Jn1cFbHlSwFZixNSU0gCrTzDgWHIS0nbBzSM+8jiOg+qo1p35eP5qyL4nzl
qvCo12strXIpdum/DamNEa/x4u5jLKX2k42waJ6vs379nzHlSlPH/aHaqVRzTCJt
KJVYFynrQmaKsJhJlwHrCs0g9bA3NtNEq4YqgpFpJxDGKoaoo2HlMWbPeFdniZIM
oGczqpzaanAUW0irAoFPgtDpakUjMCKleaXeA+YVTI1/Sn4w+suIY8UYePx3eg7H
mBBwrWTSMnBNpTbfpLI+FSm5nNxt1wUMFFnis62+Uv/cZv06AhTT95Yt3rbV87dK
ga1exjNtXugaJtihgMTO/L0TQPcr2iu+8ikMk8QMTFwKq2F9nJtLsP1fErMFymeB
5gU8HemJj3GZaLXvr3kPl+R+gIyHQpg395OaHv6VnLfh/AwWSQxxRkV+JZjg+30a
ep8qoSdS7RcPUXh1P4zXDnZ7Ry5CL+/G4lT7bka/mlCjxen9rnJVcMAOKTZ59ptq
Mal0ZTYd8jwz/hUL5K7lWIBUem5ED1skZ/Ez2UQciJ1NYihCcCb2CP1ux9znL324
IZbIZ3WK8vAZBuv6uJqfWTKvCf6ZjVpI/KplFTyzUgmheyJ3eDYOD0XalCt7yEZE
8Qb0Tkb6p2ZY+UX1YWHbxceqAI0BBeVJJvSB5s601IygG1aEkAssxdRCj5NZ0dQD
qmO8AR66dIqpg579u8fQSbASzL/SUv8KNsVNcyrRD6+gtHcqKTbm4mdTxhfwaA5c
aTPdG3GLUExG/nUtFVIk3FxtSVkn8aDmJYM+tYhq7m+7B0+nxhndZxe4zKyyNdBQ
mFBmAuiQ5yiKMjM29R2dpiwFhohVlc2bn/q9tmwmuzkTSOUO42+pVRDjjf9AntwF
Q0IY78Wju1oJofFt6hfkKF2WF4FI+KO3v/85DqoiUEyqQfAbaFpsEfps5gb8XjPe
BZxEnVs1KppyE3CXk/1qEoW9DCoHG3TevsT0U0Suvowiob+wnpfhaTp1CzMm7G7F
ouJS3KnfDw28tfY2v/0bRTsuZvhSHVbwIhKBXciE3A8ZJ09F9OHRGbXHXdeaMYTl
xAuugSsSQyNJ+JtkwhehEXliIP95AxYOJ/TYzWf0j0LRZYav80vhcUwn3AnLODwd
hj8Z/+ZxrKcTlU1kQSLgSHKWyUGq01ig3n4XeqPAaQt14aibgMlfkBQANYoh/4Ga
k5njzeE+VhHU0A4TjgEhgphTnJwzjHrPixsIl7iG80tlLQVA7HTm1Tu5rvfRFVkT
A5YsB7Oz+VXMejYEBAkQ0zkyMGYvuA4ct0cVEfNVq9nmV81ryXXN/niG5QR3NnU5
rF4jkuLMAz+GTSTJSb97a5yUOeocykosElHHTg9Atosh3sPNNlpswu/esF9tdRxp
/fVOtoJ8COecvFROAOGeCnBnBGm4XpsEhhHEq/k46Eth3wnjMGFd7Ag8oiEakRhb
kUSyerEov4erQIR89wPDvrM5R6NO9LO9TX7ARqsEoFuz2UuNH+GfH8xq9k74BMRg
gjQ6W1RI07TyooYxZjmtVFHFfRMD6/cvr0GQw3eHHvglLOfzVduwp66vtO/Gow8v
8BN3i78A3I6h3VhsPbZRLmiQuSbrZDFFMR0MrvIurmT9H5EguXoJCCFlRUX+za8j
W3oREcrRRifTFgta8oZ2gPLubHvzsm7US9/n44fdAS/U9QJTmgBRA4MTNYmcaGNL
Fn4Esv0YjtllGP5aqLY4OSqZUI3jc0x/Rk2uj7Hvj6QT/Q1Wlo8pNGYvyIjNoIWW
DCHWPNf+/uzLsVVP13TeYJU2vrBFvbhlAHQynMz58U0eMmlPectrz7vKucxmP+Yb
V4Z1KoAI70Bq9LTYQsaQKIf07uN9/uKUbHSf1eOIaU6leYanq6+bC24xDFOaMLD0
OJ+c9wiZZy+V5ZEP23hLpRtSNjXP0RcxzGF3YK7hbrvorhKeaEkpR9rw12RQzB3I
nk1DgyI4TP4AI3aIGBsOVvJcIDGEm2hSFqrH1RBPguGBt/jxG7SzzFj8fGm+UuRM
IeNjSJlwY5+YJC4z4hIhPfOaDCQ5RnUDkxeE/NAMpHchOoAT+LngqELBL/mVmo1w
TTWtT/dVnDL2GFlrX1nzKYki2OC4pZdZiaTrmVf70wh7/JUjRnqpyU9UfXffbHWa
jKrzyOarSl2tgEI+hLsVseKNNvw0KVXmDaps1Iw77yKbZivc0eE11rz4WuPvbMzG
XO/zyhPsG799iyL6dcjJu5k/7LqCsdaWP6xXL+Irsbl2+L59MABpD0N7UU57TiSX
R87xvMWdhmPsXkFOcwuT6y/uta/NvVOp7tHd0QjTeKN9Qb6ViECaIoDITGHkmDAd
f/TnmWoRabAosXHcF2yUUans6Ayq/AhGK/ajE+1iAscRsZei1uhlEHc5pRuEWHqj
obaXItiCipin9wkxQvkl10ZW70Zte3jDIx9BrH+GHInp0rQYIOwxllc/pVAWu24y
LB3a/UK9S9NqIG3P4mPEBjkU8KpPIV+/mF663HhNkGygvFS6xtTrMRxIIkYvZvfH
f1QTrmI1EJg+eEl1nVWbJpLhjWN29twLZi6INeDzpCvKqfxoBuw3Mwztii72hXH3
hnwK3wDFkD+5FA0NtnE0GmiIz0Tl61OqP3dIN+2He/POQpt5CFlejyiwYOEhe3WQ
GTDkxwwuMSqweZW49XDF+Ss02XrxoAV0LJoSrAmxTMUBfHN/GaCxlQutemxkwW5M
eOoxHvM5zcuoh5vjKfHD+l5h5xbJtC2STQEQojgttmfux7pN0shsWLflbvrUhRSJ
cbNdaUzNXVIrqUt4JOvGVOobL1ddMytdDWGzo1uDYGglWO5fPWw8gRNXw2HlF/y5
raRZ+SpARdxYTXmVSS8MOS97zsr72SQUFWnWUmP9RIEzLmZ5PDh9ms3H2eKkrqxr
j/Lw5Yn1DxDUSH7sf59qkr2lBIno1EmxBM19ujCmJESgs5DeuaC7UjxIbxyfy11y
vG4qDiYXApVE3ODCaLiGBgKk672hPFiBDID3oy5yNyLcIJno41c8n9HOva7zP4XB
AnZIaBVjtAB3fc4Xm8/2BqCEuCsvHLyCoM77u2jMx90b1aMQQsAd9rA7eYj5iZ2b
ZDcJdW+d89k4fBzL+2v774mckIbCWv+Dkj3Xdccgi2R09Su1oPh8zbnHUlTxyE3v
VrYsz9UezEjSSjKNjkvb7i+KV5BL6Tzg6B+rqPy7QYIxAjFcdmTK0xuOzEaNrbgi
ArnH3uVVOeeQ2gh6Az06K30JZg67IOWyyOYLPOwwoXkSVIzb302F/rooQMc20i5Y
mRuIY8JUdONEbTFO0+xAD3bnzx9PNkgxDWAlOOpdOVMt9pbBT4WMihIoBBDRO5hZ
rD979O7Ilct5RGz2oGnNHJNQ5JfeLrya2Vu97QQxjYhIrXaZWL4ptszO9Q1SKQ8G
Kc5xeeb4F37RmDa7Cpe7CYRIv/zia/cA8guNBtKdJ7Lcgvi6DkTl2qFmlYQZkKBU
GTGIPkm4GGwyoC0oWL7pcOABBDUxXNDynSKc8Zi4pGcNckkCQM2AIQEVXN2J4v4X
gNsLdczGX3447MK2n9EjSv/eHd4pYGZJpCzBZpy3gJdgRNWsRjCCoIGT0arX5b/k
qNjzZyvDR67OPQMbzNgVMjsi4Go67KcwU5LK8SdJyXFiSFahWTf5DX/g5S0Be6qj
wUo8iJGEOMslzWtvFh92W9DUzHUNxzBlj1UL8UgNeCNIQ0fQ0pR5TFEdxuDT25DX
dKRghs4IegRqt7zYjdvB0w00v8m5kjNWuIt3Igw0XD5R0/DO+Ps2+bDfWc9vixJj
Yl2uOY/cl4Bmm9IrtRAjwshe8igT3jth9I8XuRLjEKTJ0hN3s9IZW0Kq74oaEfDC
IfTR9Yq2HtSTvw3HcilRrgS2hjev2eAsU7weZ9BletAQU4wpWnci5ksjP87/eMY0
cTGH/pW/t4otfYTqZCwsz7ZF8MMmRsyIVbi2hjuS8GFwi4Y/NBswqzxHBk1rMlfS
wDu9eJNtH0K1FoVoEIL9bHssJREgWXUqRLfwhTyCVdx++UR5p+zFtVLFXJQ9ArLo
9Vs0XrFOdADycgW9kKefQ1FyfAQlL2iW2/aNqgRfeB3nwCFXYXbqxsOffEn0TzxC
3MV+JI8LMEZeDbiyKlQDHszDz0ctX6/C0VChWntV31Ilp+qtFPg3VVlx1roAEdrp
22xQD/wshu0AjgEyGDvLh44QrFnUx+cLR+o/zsv3nZQU3vva8ItQPsdZ5I5HbTLa
ZauyH5PbuQwb4WsXo/8LDbyuX2mpNHmZq7ghw7RCLYf/1NB5N8qjcnL83n/i5tpr
Q9buWYd55EpU7jdv3PCy7dGPt+H6OEGxQNgQI9azg+hb2kZ+E02KjgqM+ofbo7Q0
NgH6xUGPH6SX5z2CQ0QCTswUvDtRGjiS1igil2XWyyXPywrYasO2YBs8XvqUwpX/
6Tkw/Ly62yttsU2QdP48HHKTWRkG0hoQfH4MsibVt82Z0zudrx0ZmK+CZBySBK1p
9XhXLicveJxIKKg8C53qES+TJ5/T02pd3eRhOWKsLYpuJy5He9MrvSiFPr3q0p/y
6gE+ZS0IgcQJmmADA/P2doDNUCvpIUs4p+ChUbbO1vfIa4uB2xdJJRrIWWMZUP99
siARorQLubMW1JnR4fUDNSqHtLd7dbwhw08h7DD3wRvCgQazjE1SrIF6frM9xcI8
IUcg4G69K9vVMhRlQXCD9AxAPcAxG6F2Ur7Zo45Avt2KvFv0WoGYvDTAyb7RK1II
siutwIgb3HXZLrFezLBidZCPFDk6Jr0bplduOG6uiR13+VleuCLrKf4gBFkithsu
m1zjW3K1g1kgvXikTfdak4xYcZyu+C2TtX2xPURQHiD+7RwWtESVvppbdYKwpfL7
j/B+K1kAfJRqWE8yLV5aFZnIhBPnkz76W7TRP7v5benSF+vgNnQygkEEy3LlyOWk
MFAAuhLc/AArbAJHVVa6pDevM+ZDgKuoQAvLyMCLTQpCvmWDQ/pHx+u1wo052HrL
Krj8s9ArJZq+JBe5gkxyUvOoG/hhDNfpU0LDXr8ewb0R0J6und9PaXWFDPi17Hur
0fQlnCMPtbN5IJ8F9rUxc7Le/4K36TRCcfJlZhVvQQhQ9Vm2Nhl4+iyxepKvb1qA
hr7L9bAeUwJwb0FRn496/lkO3yAPdIsMnlU94A6jjUVL6bOkf3olfbdNp21epkVL
PWdPChM1o+by3+vp+DQZjGNgjSmjNiZBk6VLEsy6iwrusXhDQEhjt5LRKDJ0gNgV
ab4sQFQihrykvwA1hT7pdWt/yEpNQBhxWdcSdJ2R3D584MbDUDEzvzVU69Jl1DmM
xNmSOogsYIbCSdJWJUVcnnmSjAaml6+Y4NvgQkOJCg3n2jrVsi9zPZA9ztZ+Z15o
KZanndbKdJ7DFUB4bZk4MxHnneUJonDWb2n+VyrMF08K/sjlKENCjsoKyAmhN/7K
ZiDq6UcdVjrBWPUTB39lOPKhpvqEF/Mu2bbiKDv0ZeD6JWLxdP6rmWNy3/8RxuGz
9K51mknKE4Babney2MBVBN9zHcK7Ak5MAWw4VZyHAjcyEx0WGRbss7C8e5aa29li
9NDuKArJQ8uOWFiBTC/Yv6ct4neefLN76W8sVWXwYL3DiuY+iRdD3NWEaqpjowgf
LWM8qJmI9bgvWYZXJrG5R3v0fz8j/Yu5b5FON1Elyz0bZBvGK9LrzVtbd5jprHfA
pFGtaUEi8IBkL4IBAWjKPuWjsOzmXztpqSnXQzEwnAhRcCJJMNrr3m9Ghi4WlQ61
zT8u2Qar+IwRpIpkD+CxpXK/+ZwpZfsQ7IB1vZffr6l9zEty5e6HpLcS4vXFgdk3
oWSrc6SD5EjmT6V1jAaldwNTHjSzviCiu3hM0seZpKKK/lIWYj515Gf3Yvj0lY0V
e93u+w/xCp5OTXChN6svDG7B3csC8hDcj9TLtmk6TxOLYupmqpoIZi1m83sKGmEu
H3DC5cCNHTd0I6uzXmP88EuyIOIXZBHxEcE4XcGjA55ZtmkquMMu/tXzovu3r9lP
63ih64FLQVqYBNGDbPgXlF9wN6Rq8pvrrxH2OAkYqW9uPnCz0wX5IjTo1GPbF00g
fQvL2lRPWPPUSSS0aEwpq6hjYW4JT6qLVCpCIKbEIaJ4f1LRmtkWz1p7EIp0BIhV
Z5aLQT7IadjhX/6wufKw/HnEtTEb/87mk0SoF+Mq1YPPglcmrJXAgpYtpv0lwGCv
IuFaRxotXsJepdpzd7fWsKhUSbz6jTJ7GtDoUxMPNd/iAHyjfuA+cmq9IEbaZqZ7
K/eO+i3/1/7sTD6F7aSkZv+eDPaiJ2QS3ArSEa9t2OF4l9XZJFHxm2beSzFqGTVI
qjdyJ3huurVosgMinbNruGBDoXDpybj2QoHDvRahnnrpdz/+Oz6WKwnGYleDuEz/
kIL9+3e+jouOKdavd17C0KsU9ylzcLcQCDTy3hTqlnm3t7jN2y/Zctyj/JRnlrwR
/zTPPQo2YNXVgR4D7qC8nqwosA1RMoHhw28BYRnEXODwFjWpCta6M6zx0IN6hRQm
OfzBMQRFIxHN9ipf7uiMBWxdB9I8aKAAzK6TTxKermIBjCgh+gXXAOb3RaySdEx6
BLWf4a9qAhnlyQBCkXZOGBtQKd3sQ18pIbWJQmQbSORbHcq3jHc/qWzKNvgrMcmu
ezlosGEs4S8HXJHHa+wIBEmDr3yitQaFZfdFUMCXo/SwXX6JJhmmLVjK4IjUf5M1
yvq9N0fw1CulEQzKqUAtEN10C5nVPhGDpiHBvaCI3E35xeCVvKCElFsw4sQqaFC4
BoaYNJXZH22i7RdgbsANLPa+fmZWne7Czb8DWd6avNl740uDncMCuWXkVOPKzZYO
UsPxgAYUIt4ldAFRdJ1lG5W4pjoD4/OsDP20iz/mVNJssz/kD/diqSuhUQhXHBwd
/RWaKbjXpA3A/geZ+eIyGYnucxkd7qO/9e7pcgINknC5coo4cTtoRVuKZG1UjOMo
P9XBK1UwvTTMMHrHElY6OB+a4nts/TW5VZPQ6pTPSai64Fx/l7tsvw/8N7I6mj2l
Pa6yM8yf8FrXRtjcgzW5F6pDNG9dm96eFzeWAqS4iJmzK3xW895dmL+WqX6b4/ap
hzxfXv2TO/lrgcsxvMlRGuiIkWvfBdg+Whf84d0fXLMwB2zI9Dns7izb0BGKgtBu
/7yWWTwFnPEJ2GPdlUa6PoXB6fLLjx3TU8SlNSjLPxSImGAzMoJon/EGODy9MpLz
4EZi0jYHlpOwlColyvLXTEDExu0Oq7QzAoY325Ww3j+/Jr23TKVArngrIijCi6zd
pm+83YYXIHsLoS3e/8rJiF3RER0JG6gOnPsRd0wHr9hMbpBcr67M+OAybfZyY6Pj
XUHPH4tRIyrhWzU0Oe3uvQ75nL5w6mdtM2P5pK4vWsm9myLlSBldPRW+1OFCRsCk
w33d5gZrFN6cQllZYm8Rjz45jOvUmXz/fRY39ZxcwBpEY9PaYlrr2/8yCbYTUPNE
pk67q5hkYIBCWPNrtXDFGGAD+N2VnfUH4jzuTce0wppczlBWkIDDVoCL1uqUKzwj
IsD21H4X/ag9OjUFCDNDvBnAknCt+qwxKytqJTrLWEwFtmHdYC9nfTK8XNp4C7QQ
3/alQdwIJXjw2SEnWjX/2zROfb3mP9ONTUrypEjKysejj+OumO+BQ+YtUDRZ0KHb
KgV3H37dNg8umE17GsAdhFmZPI93s9TUeY4yS5Ekb4rk1/5N2fmI08iU0Kb0ZNJS
ecZs0Wit1zdF8xEsWc4rezZp+XmLblZXqad1Yr03imZ/aAwMjAJ5us+rSRufk4UE
xMbeW1/1TQthYe8E4+HgJyj0vOaU5AY28BdLEa3UDD1EnUojL2IUWrqscxA7TrOt
N1/i4OELIVtaECGXYF4kgZqt6oKiKUo4DHS+ydRfpNTUIZbMD1gxdjZ4zqTm89s7
yynJRT6PcLAwD4SEWbHTqiI2YhY0hh44F0pzJKWSeBingw3SH6/8kknuAeyMvOyA
rZW0Px3gyzshFg8aCW8t8aXwhm+2yVuC6+WKCE6LLjsg+LUoFld5KAUk0KOAoyyO
yI4VxaQBp7eoGVXaZ295EfczoBLewbKDsmwUh9q7g8cLR4uzjjVvpcyFNVjKVb4v
014F2W3lMx27qoBIbi4ME34nVpGqN2rTxSGjC0XPFKo8m6ZNUbLVDEa5FY/lzJZp
Q6jdmuKepB0u/kqZVpaBbxje9TDJGKZuyCwQ3jfVI+wguv0lLuzaXBziRxzG7X/v
aqk/+kqr1hsBEGaY0bXpsdUx3D7xvpL2zTSgpUieOmy3ZboDEabP2hgLyX4KXzeI
mTFFARUMuDaadnmf7TOO8gN+Pbr0cKWkRxR1AC9tOJT7e/rR4XEDYJV2QjIakECo
SM4gJ9Etf/KCoynqLTJpluaTtNPvBdYbM0ME4d7Djv5VamIemMDV3Ce2XQbHqCtz
R4wiLIV2jNZwXlEaut7hbl6AAGa+dxHMDhHJtlMjX3l8/xu1t63oszSKPgtD6gMd
mxQB6ED70ZpAk76GcGY1c5y5cGDHr5zUqz2VHTNH2dAXhfVNQZ970V2f8GNcvCvI
1fQLN5AB3tyV6fZvg9c5Y1RaymUKx2sNRwoQ2fkR7lV2icYaO1DfVltgQjnVNG1F
Lo7s3GvrwmOZdKnAY+hmTZsbJgKtWN7L+rNOXFfH5DLc02JMhNWwRo9rlap4GVj6
R8JHJsk1IXTMQFcp+HP3bOEN5/MsfeB7yeWK9eqxqaaZy/EmwEpFfvjRPZUofIiL
RhaWk+hGtPXceFHEdveanGVxN/oN1EoNxBWDFzWQ/xiqA0lKABDw0dsSoCm4kWE8
acJVLutdKvSjW6VHS/eGAjYUpmTxvAtFKXkyXnUHmlhQjqH42u+mmflJosLe4Irj
2hzoEQzOx9oNZjE6OCf2juV1J10Llmm1ziJQO5EsaBU0eedjntKCfWVgeWn41Q13
1Xil0uEWmrMfz5uPJbn/6t4q8E2aUkL0xfhy2C2FWjuQZOaLEm7Bz0h50UoYJNqG
+YG6mXLUXiN+giK5ZDbeKC/35Gy/TiYAkzYdzo9N7W4KvQWH+R75S+mTWBkarmxs
Dcjr6N1FesM0pdkYJYdOUF7jVBH6em+nn2sxCSUbaxvf1pOatzlSd5bB/p0Vk0XE
eZpTKApN6enoNIwfS5tkh1wgWyM3jhchhcfP2H879iVzvSYGM7aNWoReiIn8Qevg
CmrpRFhPZu9wGGUBS6x3NZnbjdEVvN0AgGwAyB1EndvfZeABhNCLtORNvp20NHTm
XUxfXomqrwKAaAJk/3l+NM7PyO8h4ZrklMg3xOjBK6wPzxEkt2pI+v9TMw/TE41d
azg+VVkwZcq3zK65jzho0ty1Yx5FLQY1s4xQEzWhwOLJyapZ3DvA+voVngps/Avi
hybPG/7O7OgX8iQjxU3VQRQL87hohKRW3hWcyipYi0gair7FJM5euq+rTyu1rMp2
9g+PH6F+Ppn6Ejj3DTQ9dnKy59tljkFOpPXHCtTtKtFmNSfhE8gDHDpObfCeAJRZ
70L4wM3LMevzO6Qgu8KlF92hNtDoDFaOkXn8wDhzjfkWTQjVvnqwqRde9lpWGgjt
F2TUpJ/fgWQaRvqNuhpe6tQc/ORnAL2wY+/RiDrjeQ0VCTdbahTtY+FSNNBaLk03
yDxEnkltZv44j56Ok/zyGZJh5vGi80DP+MD22ZCuc5i+vvfzQmxHyZYa+SnFUn93
5//p4piD+L+0ixNr2YVl3nQPfge0uSFWGpX4bUq46W4hAURxfJzaRBr5Y9/ZjMB5
0CsXsCJr0SdhaOV830lK4nbL2Gl6S8bzqJ9uOuQVrQMCU5SHlCnfZQ7ayzHrbHhC
60UXK2q2/n/G9/24W4FLK3FUtP6HvZiuihFQIcwwc0WSZ67lE2iS0LPG+NRxM2Nn
LeCYK5g8rZlJ0pGYtG0+J7NSA9dU9Zg1M2LMw7AeZGQXDwYz8tsZ6+KynJSRYqLt
6+RFwFveoGU2vwTI6LiSwCcycouXsEmVWXPNXWjmv95wimiPfFyW7jkv5zJJ/g6z
h6pcENP84IVWCun+3+vDuZX9N6Am0M+S2iQCNv7o6gAGhuTMBh7TyI1tdK3+Fkqu
OgYXhOA+21vM+t1WIJ0NP+L0mSbjo+t6YJ10wZD5NmoUmtjH+j5uPNNFC5Fq5gs3
D56EtzxXRNm14aQ7AcXKdckp1g2RYf1IPKKLW2+/KxeSnBR4KxXnyK/TQxbFxJuF
33QPG+sxcKKfuzK71jkjj7bD+Z3J19pV/3b0KqSbrfsPfX61V6QyNXIHrvtwJ/sc
HoIgyHw/TtDdP8Km714uqHMqYu+nZiqRghBbsY8qdYW20JMX5xTlWUbQJPIJ5oUO
1moSDyByRzX0B77cYqHH2ohH3/MsmmsZj818w/+i45caVVKPQqi8CNiB4V5UwEc0
P7BAJ01W55hPlAjt1+K48sTBeCB2TG2QlalJMC/GZbCHz9Zlpka4U0n8lsWuNRvZ
P6o1qN+2GAQoXs5qmvpQc4/kDST/t63gf1CfSsXzmqhK+I5cottQtq5bEM5/RAAH
4MhWcvX+nIlNQDPdP5IjmfnyBA//hwJ9ajtzG8n5IvqdRt2UI/7KSMY8Jz6JhKI1
FhFNNdpMxDSP6yBgovIYuu953SRTuMOUZXXO4LCkcCIZq2dXC5FiJwEWJ6I/yFh+
xwmgiagxj2oedDfsx4rhExfnUdoY0utukbdPQKe9UnvxGzHn9SKqgNe/Wx8a0vnw
DQGbVCOgu/EjrmElDrFocvPvtcAeogWfgqSaCaMER5AyO3tvk+kpGrojIGvb7l4f
Cla/i0Rfj1ez+QFQy7hsPpTTPSYRsCsMZ1lbETuKOBdX5sVX/FjgUis7NtiUu2k0
3rnKiv4a8+M4KS1p0zZImTTjUccqK28wbbWjO2TwKKe4VFYaDJKVrA7e+jTR2sMY
2OZ5EyF+k7rJ8MPDvPusbQlRXu6LqhixK+HEwv2Iy+TWYyrL/WCcZ0n/phdrlO9d
P7W4XqgYJWO1XhCvIUm4K6FRS+uF12tJNImb0SFsG7lYqAtHSO2kqmyS7uUwb2vD
fXI48eP/HSyptV9llriV7H4CX/Dgb4oyp81qUWZQe4qxYugweG8eVqnIAVvypihT
8zfWBTWNIrcgimU2JTuUyIUCk1EsLt6nA0ukINshcCc9Rpz5D2qnBUWeM9rshLvH
6IZPmKBFMUYZ5M1sDBIEYYDoxbJyasu/epk8Q+2Di5l/fZYSSoQePYFCb/VpymmJ
hhCyWmpa0xE3dqZfeYYGOe0OPdkrLY3burTSAIUKca95nrAcU/VtNqGfMQErXaX5
HefCRy5qu5XEF6mgT1xvL7pS6LvgzzFIQoY3bygQGImO9szRlOYCaKAOreFlfg28
wkCYYc7M0WEumWADnVBgqu2VaehOjxMzUfnVUjyxOjjnwA0Yz7l8RdDsoMQxEKSf
BbzxGyORh8jJlNNzRP9jfY7p+3i8MS/znEVVa1SzO1xO5fSKIUiZf0CtHq7QP+Ui
mB0KsvIlB3DF8udcLpqY9lWeq4jUkSAcC6P4cMw4abUu6Bnl/J/4XLE5LGCaI/Um
qPoxzQ1OEQlT3OvZuoqDxOhCBA0d3Ork/WId4mfiBRKzsWUgDdoLwfQ+JJSq33ek
busVoliysBkt28Jx+dlaFC9Dk0zQYzjxT7ttT3yMFiiR43XJUtdCDEKjyxgJNvSk
yd2Dzrtx6PDggKJiPeZXxqQPFI70/0eBTiIlAiTAWO2vA9+Mel+8c4QfCakA3GSR
VHWKbMu0HaELnMOHAYFujrvE/ODDBpoWWFUNgCK3jYzJLskEo7H5ONVYnKoAeb9E
5Zq15Ah1Bxp/rueywCQdF8IRy1ZNYVTkJr8VX+VAJuSf4aU5l3j3HjhOH/pS3txU
z0jNu6L9HGGVdVg1wuRuAEb08mDpKUz5Siau+1EtV9QIO1UI3F3Je7q6zr1+hYQG
kTnMZnbK7Akq9WiaokzPJlPq3KFPGI43HuskPN/JdMvYn7OYD5TCO9nK8y2yS60k
KM1yVyOWMhBHLvFqHLOqc0oPtLm6VUyRtdaAeXUmmvZtoZ/Dhx2wvLVVnFxj9XyL
AOjs8xAwWE6VNUhgAEMKVJHdVtD7NLht8e9Nj0/RaSGtmA+niQEpsZE/2QC+GdJ7
MH6fEAbejTX7uI9mLknG0Z7SgSABEuRPPC0ld6TLpkp0A4toUK/AIutnIPnrzgBP
mFjBtz1udyL1oVahjHTE2mntktNgkFpX7yy4IS3FopJBCJHvNIhkuVBDpMcpFj9n
PrGUTVyt0M6VHKZTjDtJecYr1ECEW1PxZdv678DpkefqRXZfmedTYXlxGM1/a0Li
/Y92Euh/shWTyPByRUQwFfoQTIEHLspAlWwpLBfncnOnCI5aSfXUG/tsL0sP6lZj
FBU5e864QjSULWsM7CgR2yN4lm1LARo7BQ7HcFaUXpd4YYTM9Z+O1LFHQYzLrbyV
LfHAB5AXu8niUlulVXLmhr9RVO60r3l4qsmW7WGgIPNv3oqqoPAq1Kldh+YDJ22W
WovFzIlo4lvq9cZzJS8oVjGqeN0vRQEYEbYQj9QikPkXEYFoTvht+RgT3DrNGsoq
6DPYGBqW7MugDlXN/QKM1bOPrQtRU4lPLD/3bpRAaK50MA/zuyzkjl6B99yau4nv
MascRUPWNNu4a8bVmNdTfYxPMO5GCAXUnOQYuWa8HoMk5hPw9ONibDL+5RBk2ZgJ
nMe+RyuGFXJLtTR8RD971vfPkT3gNtoGz1y0jE/zsIF6HQ0Episx19yQrSBGSEP+
NDosrZJC7OYKUY180loQ17wWYBwfbx46Xoy/BhafTvJuf8N2WQGp1sLkTg/FMDGD
b8bOlPx2c2yRIfE7iJLGZD+b8SKdI9w63Guw6hKaqK0z2ytHRcRBW2VNkcwUY42p
XbykJPWEuRa0zXUc0+5GAfkQMUy1q8yajPuY1YoTRK8y45svyCF9hjrN8NAKXM1r
AEHV5PBRQU2elsqERIbnPYsdYdOC0StfgaAYpAOtwvaWTOm8UbX3gndZyoE3sRdO
rhWoYeTFftldvsVtcn790jKUr1KVvzO9+1N/2fJIbiPQJXB4kdKO5h+TGWz5ir8r
4oprO3kwD3pUVZrvT69Ut4y1f0qx7ydtMft+jKWRgpZognhtBgGDWpBq9GEY40ef
2e957cpdeWHpuNhB/Oxu7W5K2Yj5ltq6FvBqQFJY0DGstkBJoocSkKBZKA0YKsQO
pPXX4wqEDO5FMP/BY2PB0948d1zfnbX1+sQCEBtfvqanswRiEopxVPUEUUvJM4PI
x+uc+PRVIKvF9V5tUtHqHrNsZhovdN2m7mlYWzw3eQYHVQOCS2g4CvvD8C9TXkF3
7eORYQOih0CbAstU0VNaaZUiIkaWM1UB56jmPkPdiSGv/fAypkiUEweMQQCM04JH
Rm18FDe2OUj4ImuBq1MgOY65yX3pl0d7iknFBNuqqTrA/e9Sh5bHjcFh6IPGmZr2
HtAJVq9H0pVWVGUYZPb7N8ckPBXAiy0Iiw7RGX5bX+jXly67yIdblHcHiM5ztrpp
cBqDas5ML4+RVw/VpRq5lXcAc4rvvlFThYYBunNCbNjRPnMTfBohYxQ6guaImlD3
HMnbXqDfYj/CvGWD54RckRdOFgM6wSlSza4Hc047VhjZJqKJwIkq20ZisxnhWwTW
UqlxhGgGJ7aDABQcE03UsYU/0/jLBtmx2vmTL9JPQ35h3+UUqeX72u/nkXzqGx5v
s5aKEIXK/tQHU/E1QwkadSmTHCa29smZRuDxRcPhiFFnYjaPgUSD1K//cbiqppgY
5AtxWAIgHlAoTP9nTlzTUGj9NjqeHqICQzbCrubUz3mY/Hjdua2rBZPJjgtXlTZx
ozy4jEiXgBaXDxprNCGLRkpofPIj2NCBSqgX08wy/9Jzsv13DNG3um/SNSNBO3Vd
dv7XEpZekGNWwKv7voAwBzEXgjwyghqPEHABh9j4dllHwnvjNLQkWMbCv4fgoJq8
pL4iDbJU5GkrHaU67Kx+9WuBHjEnOVr0xLfINUe/SNhpsl9Il57jUawCgMRlxxXj
g1jLcCYCoru74HgHhPEejCMEqrE4ibAiGwhkCpDww2P9Qypi2TkcNj7D4nvBfAnf
ANN4AByC5IMGGvpqD/fCV/uNQXA/euEH4t62mAt8EwbCXHIl7IXp71wureQGgQT5
UsmAP8a9uk+jfHsKQ6UupBPWNuK5TU+cM3Ag7DKnLGOoiiQXMOcjGc4YSnlNpPIJ
aLWjjFHrtODajsI6iWeWiA4bSGT/NSWxrJG9xQqCRo6qV9eQwYtsY5B5aSTIKYMN
HbTw1KpFHMTfGDM/IUl5v8bm+/IbebRot+HP57PVd4DROWjs6nwCs/HlD5z50/60
rHME2YPP02mrHEfS3XL0wuJeuRISEzhh9GjqYj9sIfSH6wAWiWUJccnzDvyRDEMb
lSrVPxUaTtuedfJuHdxxSTZu5CmTB2lFIRKnsLLOzgdcgWNreYGQElUrEman9nB/
fd3gR8QHgS0LRwZll51vu7CEUCalwhYgtKbaH7Gi4ABf9ch2xHawqhNqmTSrvFJ4
HhcGk7QubFBxX5sykoSLXCz2ZamNA7RUK0pDSKjxmFmNtiY2f2irG5EdenDrmV2V
/+0HWS0RJWwuhbdko8MiTydDkRL10Pp3sMhn7+HnJEWMFNJ9E0AHPr38uEWL+ITu
YZRlcnrx1G6XR/xv42rBl114hvFFyKn4LxSoBZg0oMFIotGOCcvBsTPyGiWfUCJA
Z5MwRQHbiuodZ3EyzUZNyt95O1Az5LBkzG8ASZcEJpdQXnhcgfvkDpyPTeX5r0cF
rS0MbRpxz9fGyA+hoUpj7wqiIS0IjrxeRIedNrUqYcCHVti4EBHpK9/H5iKK+SFX
c1wRHDdEns6Asyw0fxL7d0/fewktI/q0Hbuo2/AWPe8q5aq2oS0PcVlf2NCXNwAI
PsY+9jcDSDKowm/DxvF5KhpY5Re2crDBXZYdAvlYuW/1DOiDQmBPwm63NTd2XnFC
R5HwFOdX1Yg3Iq0I5D7ToQFXIMEJYS5DXsPSm4WIAnxLgvdeWjDiBL0jARwF3Bpg
QbR7+XqwESwREjOM2PmspzE9YCMCN8zk0hrCApAzufHr+keecLUTMMyyFigALjJv
K8pT4JBUVQprkbHZNPNDnwMZlumJIheCkCvwxCPZO4S0PnugPLIlz2eZD9DJtzIH
W6mHWeoKZAD01PyLDdjWAUFof8rh1hW/7ht3CVDogFTiNur6hQmflBvicvLZXk0P
sDQBcp+jKeVVo8FCGgDVQTsgtsDkKLSXWIhNePOiTkPEiTo7XYAGve3l2oaxxV93
Fl6vslnfIw77MXAJLQBojrLj8IJEIsKEghaK7J7H2lBOlMlyjfuvYYP6AmJErKg2
bvm6ZpTyrKgxeiIhomH/UZMXZIbfOs8nPKMwfDIWrr5+bKrm1fm1gv0hKQDuI1G1
t6FopXoumjL8CZsX/SL4CaenLXJyAY3ipKO4m8echVccf3efQ7YvSvdH0XnXBG/2
X4/fvhiJkGsX1HhphVJJ46vnsmIhMCZU+wzue+SS2qejrILDrWQkw3+IzfqbVMX8
cx9iSYsh4kJ/lBkmD9OpwJMiS9MvTIgwCN/WlniRZy6lZzqUgbbZC4JBRmWx7Yx9
qOGRQOi2hNNrneVN+gnR5ockGU47MJZwirPtVastpPE/G5ZBB2WkVbvldLnFAVAT
SaBmdsh8dDhCoJjfCbeFCcd6YREM5LCav9D7L9H9dd6Z1UYZEEsIFVvGUMq3IzEZ
KG5jfJv4eLetXcvQCQpzgooDdyiD4IKd9Q6kQiw0sW5h/SGBaH9TezM/LcCRWgnY
5+DygVarx+gmURtPvNtx8CWfcQRhrE8qPXldocx+J6OU05Fuijz4WWeNL42BVi1i
55dLyRAishon//1G1HuCYqnyPfh4PXJeAItW0itvEEw21hoB4eiIai7Zy2BoktZg
TWYzrqpUR1rtJ6Lnccbavcd+eKCF05idygEYWJpDfa+fPNN6H1EVqzMv7/ahTC/F
+C6Iew54rvJwsXqpfD9L/eVP6trF50XkE10nQZToafIYGYm4Q0udhxoolkxi073e
NsauJEdMd3uGn6azr3f/xEDiRFGz+JdgH/OC5hyPu6V+8WbpnYAIWUyc/RSbsfZs
2p09Ter6Cgsd5adFfR4Jifk+I7oBkzccK5PgBj4zqlOAqay/JAxOl/Yj2W61rGPW
eAjeFnFzuerrsZ3lZVry6ApmABpsb9x2fQz+YmkNZPaPe0JzYnlIrOf+BVtdgeu+
ANIb32RfI5uBEJFh1wgr9WOmz7wU8I7w50tcobi+qc1Z6HV2ncz9fD0Al8mvY6Tr
UCciZhZFh3mqlzkwwowKplZ929Snlg2Wr9Sg7bX8uGktwMFDq7vqPhAslNUwNlHf
fvo9uRQoB1ISzYHMEvnluq5vpBVj8y8ffXA/IorE7pAH/RoDsjt58/GJgDBw4OBS
/1sPdcdfTxplhG/ppVi3MGUbjTf6ZpDlmPwftFHk2RAkC4vtVrzaczjoXp9T+xgv
NTvgzzEpklEuDorlb+ygzyETfRps1LEyYeBz0Xa+vERY42VWBh+Uk77pvkoZgfU8
u3hz5NNEe8qFQbL2F0NszBgz/BTxoI9ojvw3Y/hhNsDILAe8kGBwyYVMGC4IwV5Y
NMGnt6Lhml0kSQtwTxysOdCtFY+y54D7N0hg2XTAX/8HdgnqWGQgUj6JTPzSUR/k
iYGfXlTbuXffVXw5GwkDHg17/4nIuW4bp6bDuriWIthRvqX8pOT9uEr2pgUSzqeY
zpuTWoZcadA0UBf55MCXJe/5MGfETvsYm1qwGmkKO7J9wA2YUp6kgtFqavHB8+Kb
kJoL4vaKgSTKgMIdNEeUs30Zmcp8mxi0cmHHl9MgujPSsg5CMu3sFjo07SptNaBQ
zEASjcuL9RLp7hz4w5oB2rI1kE0037gw9vKRLBoiVn4yt28qpXZJ9ccqZ7YJ5Rm8
47g+opPQvhjqUoTtQ5nq028oR7fga83GJCxkWakQgbjlnjS4nSGxph/4KRyf26tq
/IDPICZKPS1bIdgClVhrsQ9OvYI/xz2KVLX6bnTmS5jdaXouSN9mMpkrIIiu2Pd9
Ndw1W6BZDcVOC8lkctuNercbu1q2UOqKDt2ojGxCMvwWfXvmOJniMwWubTwKzRgT
zf6UMGqYJhoYr6d1ZPq5Ps6VwAtICmEPpzfE6f0jdcT0RMuCF1Uaq767A+mHX857
6/T8xtnvmAdnxcfaBhnOIC4NFJEbr6Z3v7b6XpnmBKy4MBh18HHxrytu3IGpgFel
Szou/3K6t19SoHjOeFNX88+QsTGjIX3a48o/y6s6Tuq5MxEZBw0UQ5q2kobbZkpO
rkT4NvxFlOCJNC21wMrx6r6AIV4utvDLbsrcgPniOqxrDBmRVhoxO3FcOuT8iRLo
cUo98GcpImNZwNQZtJRf7sL7642WMa4vJR95LUsTpFlBRdPkBzD/n8t2MVrO8MTw
14vkSw8XcDBZcUelnDZabFnctgplhUVL6rz49wYhGjkBSLhDoZDJs4J6yNW7ZNJ/
5aWYWE25W1Tzs/1EruoynRYQsGYPoriFf57j27uU5lxxg2/P83lVjFYO5EI3UP3Y
GcAFdLxhk6tmtxP6J2hX9IBwlaiuhhb6kZtIoqHD+fcROLlPW+27E85sD5RK6iZB
c5AiWSFbdq30HFAQW/Ie30gQqTXPPnZ/QRP9To41glEOtkEsxbgupVqn/4D1Xo0F
UKD7xQklDK0LzuKLZ88XUBob2M1FYqDQarb1Wbv4pB7/XXRezQbZiFPy/SR5lj9N
7Oyj58sbBhGAHS+bX7UMG28fgSrmSYYTYLxLajs/M6q/tX72Kf3m47Wwkpn5czvW
Vw9tU6Cb92gOspIxwkYX3i9yH7jD3mwTz73Lcu/7+GfspACRm8NeIJ7HSXSMascB
cNd55KsQ2PDwIWx+biBNoq/O6w3hDcqYAZJOgJRWNG8miiO5gmreVGlQuCVyFB96
47/hP6FVkfajTAmqE1ccISqLOXFJaWwhuM2RWQ46KOViIUU7VjTT60IVsFtDl4u4
uZbTD2QovO/nV8hfIVCkHz+eRQXFGjgHUAfhsnf3y6pLLaeqYZ27h4vDP+RGwHjo
xWNcw3VKaPTQ2H/LU8jZrdPKVUP/OuLlIzL69PlmmKj5bGRITze8OyWe9BbxNAzN
bBpeZg8cjznOiO0ZPDsZ3LuuiPWqZSh/RlNy8VQwWLD3Grm22txcFOU0duleBo5E
PdwexqvFOhe9HCwP75GM6pOgdvRwEPndN1SeGQFwTDg0U7qKHpLl+s8xDDgt9dWN
7yFyDg0PIY7v+zjqjr7AzzNHt8771Hl3pggK2qSCQHFz/oMofsYoYs87AbVGTOLv
37kpWugpCEBAFlwJY1sNQR/2rFULf/tW6BTGDKgPq1dCdUbFsT80EURM2vVuLXQa
Qt+Nh5xlCyWgeeGtCWafVbQrUUR36k8mKR1zawHgdVUgTlxrwUuWg5EF3rbtkGW6
jAaLJy7gk1a7i1ZQ+4w9nO1ib6ICcxy45nwBB43NDLQ8aFlyOAMv9KPMnsNypRIr
T8x3Ok6kPEejWqo/EVBxVW0nznU2TP9ZGd9NceiIx1p4Z5IE0RdVSRQwPCrurhs5
8xLTlzhT1MVK/TD+Db32X9KIlWpZ+Z9MkZ5qm5B7Lk4DQuCNxipih6DRoOAOXni4
plRM8RoWWIkhGYJsUEzZht/hBci0JVsJmPnqGNInnmhHNcV/1tV1Doz10e62XXSi
CGuXdH8NNvTXVVNPuxVJryZNq2v54AFUfOUBFnLvmUav9/ecgvf5DGDNSlvDp3vN
pVfLrmcLPAdLBXwwdQQ44tKmQSMSERN41XS0u58VUoXOFxNRIsFVO6tg2Qrrugbg
tT3eHNEL5s/D7tEs5zV4KcKKliEWACl2W1gY+iXjXE9zcKYGlOF3NzesaskdehxQ
CPtoSr+IH2gAx59HPL6eLzAqMW2+65cn+8qOrUVb+gR420asNdUafUOCoztPTWBp
6WUvM3Qdu6R6Bq53JWyFxvIdch8GZWQ5MezS8phw6ECSmi/XvjUU5Y0L6Y3MilM7
v6932YB2fHQe716Wy3n/PyJD3XQxjoCIiRrNH2Sy2dac1KRY94gXxdDUNGl6QBpF
GCa4zTc5h1U8ADP7WYyuVHpkGrcfS0PzewTW+SvPuniPb1exHKXmwcgnvr0tFsBQ
W3M+CQLtHQbPzwq1q2t82aMSv6oFpv8/YKJXtI6jGZzxD40b5tX7UCdpo5H0JguS
48j7HyvZVozUcOUCfHDfzTdw8hCBseE5R5YXNYCXAzbneSgf61NO/BzUiiRyiS/+
riagMF+/dhMVQNsmHsVR3usu0Wv6y+KfzVGwvcgQH/MhvgT9VSF0V7P6wI1ufLp3
PDVrHeSyvJ7yKTsfJbPRYEYEAJGGLd5Mh9rwB4BAZB3bMNqCaUE3TVTEohPTlNaU
kG3pMSOfdoPwdHijkK/JsMSltUaSLi03vuYiIgNhB5O+MVRKhKu50Vzgx/UcT0jt
jQIneSJujwY9NG5VRRyVqj2DnIRWn9Y1bfvdwLO/AhkDDpcWGe3FyftpMvHkqyge
xG8BdrmPEdiavuCZBSOVHiCJlmSquTq+8jKPKxbFGohAhP5oSYTWi9LNwJmE4+Km
3mYMubhrABq6FTsg8lzUxFnp0OEChNj6W71sqSQhsEsojGGCKZF/YJ+uFnfOZbmd
eK1819M65xeGpHt+FmD+zMMuy5MofLTLT+nTWz8acDpRaS3Co1wfyLBXKmE3RW+/
y5jS+s0pj6G46sfJ91vZCd2LOPDL8pBar+oMWGEz2MI+fYDMC7R5J429pKvp1cxL
rFMwAfXUgTzfwc6FDj6LRY/nkKbLrqcFUe9XFe8lDtDfvVtgodnpd+X8pP+HHF71
+bd1fFXXaQuqE6Z02ogp1nqh+yHA0R1dAzTIh9dtwXb7FSbMSnXFDOYHKAv6rgCh
pIq0WHUqaLqcfTCf7fzAHEQG2Zmsdcqj8O95wyPr9ZrKwe5OR/yelAdnIsVHc3HS
yS+MsrOCHOr+DDF/qHH36FwaeUNN3Dweo7ggkJvvdzvwe1/FG140omuOgB9c8uPe
PaAKvqGIRL+nsLQfykuJGa4A0/AqI9tiEZXs8QprUivodaXImqqt8WyTL8S3DdIO
SHi9jKov50NV5TENEXC3JWuEg0M6AtIcHrbYXD2w6hxkrKq6c4Xy0KH/DucwAv8J
8XnvTOqoJp9kEe3z4/hVXL2xK+N+WzyyCQedj0xV3YXJr5DiDijtDBVyEQoedfv8
kwOQHg1Ufifj7bK38h03+2WIpMYRxH0tYVXAz6LGtsK0cY6vB1TTS17XrDHZMJsz
jkziu9QCDq4RRLE3cdNaOVaSP2tonJBYd+m2t2xJMRlhyVa6j2vpdjg+YJ8iqFJq
7J9evcYIlftBki02cSmmaWslUr+KNKa9erSTACkvSBGIR1/YhLs5+9gBbkFTlvnX
qImsFVnwkSuPn8Vc3iYYU7Bg82ycVo076OrrdUu766mKzxYCCon4reTovC+j9x5y
ZzC+kmd4hi+3+1kaZ5klxL4DyChjcNgYBjsFVdzLRkxBdU0iKBp6OnL2lRFFJeZy
Ek3ONfygh3PRMkUnswtWdhZh4XqZwjnOSfhqnVYhu2WPF9+XpX+wwxDYLxg5vjnN
njpGhdm2Npyhn5vbhAVdBq5M58g9os9d25O1TB8BHaZ3AOivjG+PsunWbag1zOmW
/WCZFj14lHH/q0bzkw8Gr27Dpz3Cfq/xJzatvAHLIOhzcB60xL92W4zwMqt1hkx6
Nk4utm9O8yzbVuUa2d1SzoaNHHaI3HzTBpifqs+eqEHhiV0EMkQeXZtUOywlQIfy
x15xjqhk2d4YfMDmudou00u3j3WqH6EsUL9gxi6+axw3OlvuyhRf934eU3tWDo05
kJ5q7UI9zLS2AMZL2zcnRQwn3Cm7I8zMNS3x0m8aGk8OM7i3k6+uWz4bVtlDnwWN
9oTSez/11kkj2KkEbnuY3u+FcN4FpqyVZTsadmkuyCRxIUK1yXbXzNq+V5fSrjJm
Skcur63Pt5nLSXVilLL0Pc2JNdOCY4hvbHXEcKKjuE1JAnOQBmcyDCkXqJ7I0j+z
VC0lL650w66Pnsya0eBW8BMHyt+LnVMsM4Bie44Zb4VZg/tG33MH1wnc+dLTpzSd
rja5Ol12hZLeHqYb13kONIBI5oGofbLgwGca3cy2g+NkvTUiXJAeElyhTowTBbMn
n/O0sZ365ZRHxH8wdZ/9vCrR+yIqP0WDE+2hqoL8kifB7IW1V5nHs9x2/AKz0tu+
hDGdM2WZu1UTIzxaXQ7DdfAHETWdB1tZnZIGqTapqRjOEkp81sZQzWkt2MD/BHiy
EKsZ6MG/slbq0q+VKda28xHqnnuocpcAQnQ/xBxl7M7uH3yNKqD5bQsNttq9pQ6n
jgHtg+EuLaS2dbGPuDPQ/kNNQsAAMd5cLhFWEFJffymrWC1f/UjmwP7cD22lpb+u
2DES/UTXqWozG53CXVMY6Fz/PURGe7YbuTxVu9qj7vcrTsdmK1lH1NvljWuDbPV7
8kkPxf3IVm6C7Rs3xdJsZt8yZaDuaCNKXqp30cnLIO9gTp6Yd/VoLMPhvMnIwwlq
fDl1MkJ0rWqVXBia/CR7pqogjwHjDCMK4gCrMxXfRz36o1nAqhCOjdE/+jHVQO5t
m3okaJ/825ldqffDUomp1UF35J5vN/Zk4HOrKjWp5YgfolFJuA4ICFh5NBuVYFux
wJrbU/aLMUQca02WtlTmuDkkp+IodLN7yVDWxYIXazVuWdZXpnvBkVC6w7+fkXf+
YMKoHWtPYvPWJmXwl9pYZNC5Or9uJm1QLED8pv+WyiKHkF0fhynadeSaZwJA4meu
4gmJEneLEC9kT729D3FJuKfX9HN3oGPWfSc545gPXrKbZ9FdgMOKLJWNC/c7ksjR
+OTElGth7eB7xugSLmDshgKAzvfIgscGlzb7EkmxzKhCOZf7IQXvzNSd8s5sDPaC
zCuvkYeoXiYNC9rzEble/J0ZYdlrkwVWQQhIJiz1lzo6zIDDxrxm5aQWulyN4asR
1kLpLxM+HgisS7StdlGKwvlbdHhik3aQ0jP6ZrgJb4N6QtM3zUPG7Cd6AMhF86Dq
Gtv4//WsKGeqWRB/81lRlNf4HoiRs4IGHlPMji/WHaAAfHT0MMjq/uxb3+Ylk9P0
rn1RGrwgi+zXojGLi8rhfFkhWkTyLEBwVTCdYQwkPuNkVbBIO2NRF0XoejgKvqfv
kYJURxm8p29gpJT0Qm97vx6aO8XbkoKev+AbWq654dkrgjPwZwleIhZP3YcsroD9
4+C5585p8wW6Glx/lPfKMnui+hds58dwYERssgnMHrl4O2ssnOqDvq6sQ7NwIyV2
CilYA36sI1FcWFHdFAftgHRuLu64NipyDjABa+7SDoGTfENij6jXfCzhIhuO+pJz
m252AQ5RtWcatXJL3Y5Jw9Rk/nABmXppvVJ/u399VWnuN1DdysxeTMd+lKjkoSgh
5+Cp0TXG4GG3yNn4vTK41zFoggbMjDGZl/YG2D8jOPq47TfaY7uQxJpaP5Arr2Zw
Tl451Of1scLwyb2aGMtKqNOyW8b6KPFn6FWfIfwO6+GnOa/RtSm18tfbhtzbDbQS
RYOzTaUimTArIP619IWh7wd3eouWAkep8wVexX+YW8lsq5qKg7p5ZJZJc9TbtrQW
4p7cv4IOWoZX3dHCVJoT2pDfaWhDFaxeDcx7bxWXE9q2EjAnjlSvJ5QydPIZ69HU
jikUkQJlcnb1+8uraStyIMAfhEOZwgtVIRa7+C9to8/Zr+laffVc9bwiAEYBnSqD
NWq0t64PnxQl/emOzCgNSwZIadnllrC7+djEvJAVBfTzhxVGpcG1ndKSZg/BLMGK
KeovESKt2pfChOrbaRnMV9RjGutwKpqd5UioiG9NDb0QzZ6TnPvra843QWGgthWH
aOuv38BdZgMHl1Bi1AzjgL2EVTldEh0oQHOlZCEJ8mPqBaOc37qYwgE4eeE+ofWK
O5wGJxKch1Ugvq1bQAh8KVgj3pOxph3CAycRo+KbVYV+ckPUMw/ApDEShPpH6kfE
XL5JvQJNcG6kU0Ek+rbyzH/oe56qBb+Tq0EFmu2iU0MEcH+YDvNlFj8cWYfHvqE1
cnsUduKgrCuwLtfid1UoSc4+UkS6lMfjmV/Ogc5MkPaXa+2nxzIZMCcQ30NqWUpM
/4xB0Vequ1VyRCSqaCP0S8p6VpIYasoF/0sk7z7/mI3ZUleNa7LeM2FZyZ/BVvrd
cQ0RCU0q01HP2ny3NOSgBOdnlTHOuV0mu7E7jWlsW5yZt9iQIr6m/3Q8SbXR8YCH
YHn4ZuX+jMIENgStIum6cIdGOsl5D7+rWmMeYsgISufD38YbxZUP2rGKya2Gx8yd
QkmSnQLf/3WMU2Gknxpz4XxpXp0NHfh+K88bitwHG7ZXYFhAdi7upvnIjxlScgoY
dlPzyoTverN+WisLH4swoo5sI8uVI0Eu4tnSS/J6Xe7DdJkeXPItgc9bXWR7RQch
AsIwFOgnHubC2GYHfeSTrY+K/Su01bTfoAgz5Q6wzeJNN8wmAb2byL5AIdy07Rri
j3GV7ViysowSmNqzqM9G1HwCPW3tleYsir1/+85K9wB8Eg1KqUtPvf4CPZwTv1U4
kpXnSAzOmIBRQyC/aIa2oDagIBzM7AvXQyZKeN90uULA/rqrZtv8YKYYaWfvzD0c
1ZLJxfq1XPNeMWzr9UIgnFKHkEBDa6DJ72HstAPmuFjcT6kwBjsRXF9J6Cl55Tfm
njzUuUmgzXvPrzcQds9M8wAfVOUkfwWlJX2Nutic59sBpygxL5g3g9ScqL2+4ygC
o5Aztg2QNny8ENYnRk+zlBl1oCCEMNIjHb6ujmJdLoa5506q+vVyAQtuDXJXxMcS
shtNplozkvmRKXwSXp8bqKootqDzz7YLXzISzf6dGv+gsIRoUtv75t+AXfgH6F7H
4hw+JxWXYhIVujkxo2twWpONU3DitpZ0hlw/twQlWNUPjIQ54dxcD9j58swZ1LLl
okXBeStlVOi5XC4CVDW0HL49eJoj7GShxb2M8wgujZOJees98cUaDRjFmm7FggVK
fFj5RX0LMnP3+JrUXxZNGS6/DSY1Q/fjW91245icfWVeDi/O6HGL5E4mn57Thjv3
PFP3IAjo4ZvidHcbj+wj7ZSVCVezlI4pKww/2Y0X/smOg/Z+Bl6alMSyy1jAfGHw
qLoX6jE8yR0d3tcm2FUGeYFMwoabdJX9LOQ9Ttay3lTfMd5jEqVYb/eB1ZZsJ0yQ
sl4OefWyckzYaU8EkKhgQsf672c2ZnroK64+sSDvBeRXQCwGDl1QDIT3TkRVwdTh
yamK5uMil/y8VixAKWJpLPF7lfdjBfNWMziHJ9VJiJtW7Bp4PjC4hzieD3BgxrQI
U7QWR1NZYbR1TioW3bfg4Jxq4hy/MsKsWeygYXAAWrRql+W5viJmsozv7bMVTRPh
0tNm5iTkOhFY4P0YciZbktNmdDrx6Sr3Sbg5XNkKz0zvU0nQI9MNHKi2AyoDBSfa
d5SyQ0RNm/VflfJ8C4pkiR6GrJKh5ni0G/ZiJI2uQ3DJsFtCpZw+U0c/iTMfY6zr
nGrZj20uH8sPAGC+XxvmmDt2k3t67bOZF/ZA+RGM0Fc2tLzjc11/P5XJD6kkSw+R
KjujTdN+2brRsn+81DCu/57a9Uk7LgznGba/cB701f1y7at/iFLQiyDxVHFgUAHl
Z7wcPfRKRaTzaShY6/zPwcf8v2IYgO4Nc+XG9tTXT1/akjLB44DKTdRJtNHKAgo6
M11+iv9bUXKeFudmvnuv7DRG7itWNZxvpTj+/cvDkeH6KNqYfEKX1HOne/0vXDs2
W9rly/cmwBCDlfQ93so9sXlX7xDlVs1SQDms9rfioNoctkHvdhoeMbDv+iUkmxsT
K9sZtP5eSL5NPUli7Jwjb6AL+3KRuTBeX3Q/Juh9J/EhaO9XpST5VOWncH5GC7Bv
hBKiPEmnR8hJdCFHyeBjsKjIa+DwPBLOnYjxr/zmXLzxPUSjBO9jAaLpy7Dk6vkc
MQUnYcCQrv83ZCgP2/kiEhcFbyum5luDUoopvMi7Iq0D3geHJJgMB0RdFwrZdg4C
Z3W7NzBLyeJxuGTvX/IYyBY3MUByB4OhwDohUp9GNpFhl978k9eQ8L6cGFV+dqni
PyI0m5AciH/LIyIqtmp2u8/PKB4kGXva+VCKh1yXFFOFfUwA37IoQqa4QRPjhvHp
2sy++nuRgbonUinuZoZ/p3eRtspYRA4wJRBpgyact/XA/nU0Q+96LhbIz92rWrMu
0cMJBXA4d1jHFOxTi/VNcMl02EZZQLrWZ7aH/9MoAkAfym6GKGpfg+AnyQRDr592
ycjwR6GprxB3JNhTLkv/aSn0mS8Al3clqAR8rZs6zd2vjfFZGQCfi7F8bXUCYlkE
LnLEd8+0cr5VVnUI+AYEPgiOzVE8JDuhvfi+EFtAZHRztNklb/emg49UKEVV9CfO
NtCQE1b0qoLVQtjQMN1hMpSeMEA0hoglenNEFuzoCVbISIChdhxQt5SQpC7c0Hcv
XGmStZyndsFoXOM1nr2hdEniwtRgmT/3ATAOYGFNgYDhQeeS6mZjopU7l2gW7vK2
GrXdVP1vfYSx02/BdPelCEnCnlaQQdGeEFqv/gaWgix0AVpksK+voUatfcu37tzQ
aAQuVHy7M/cEMDKja2FpOdKWlhiGtYDeveUZStDZEC8OsP3SH9/H3eVwJC8wDlnz
WrOoqNExVI1I4PkDAbBeyze+86R9qMBxwCPIutieSAiGakQuykGXmagOPwvIlCpy
r7N0942ABvnj5OHO/pmH5CHDyDw55CtZsKp1mvgH+mWkZmK3lYWSPoh2SfM17ijM
6Ebewf8yodeDUB8xClqfUqw/lAze4Da957aYPMH8eqNKaSsXvPhXYMc6OvPy+7yc
L7R/Wz5uTvTuyTSuxcDAXFw9XSZ56z+EZEN4Amc0+LMbfkNVTh2uThs0qaOMycXL
v+2JNPKhNyxU+vNePhEUqTezAh01Hhn004928a4w4cx5YJJ5+VeZyFuZJCjKHJyo
+IHWihsTttaYFGKt6W03i2LjQkvJK3fazjRJY3+u0Ain7qBAPaeC4ShlWH1v5Zx8
4HtahT4AnQN4y+FxcnuiVCqBA39ll2RVxmV7VQBGXtBXqmNIxcs2oIeGZ1sKCPvM
4yBArlPT4a8gRthkaHzjpUuBTyheMrO2Y3x54NSVy0K4N6QqyEZB5O9oaMtoGFll
1sAaHAlAtddc6JVm1cwvs/uW0aSvm/bGQbObj3l9KU3/8LQP66FoKg7EqmAE/Brw
UM4DuPxqu62u0fWbQ3n8qgsJswXwqy4S8Llf9hh/S4V6cFgzjm1iikNh8GBCN9by
vEHS9IoT0diAHTg9ap6eKoEOeyf2a32rqqLBmo0sfybOnQw6Cjp1G/b20W6bmZj5
Ie+MWGxGMd5xRx8mI6qEQTsON0Xl176K6aX4XTlQ2ZuIgtqyV6zzmOAs9b2npUbr
wBUDUtNHVAi6XXfLsEMKQed1TF5usmpt2vf4SnckjREWL4v8hO4u2Fpk5yduD1cs
dj88MlpRIfWPuNcH7ggR03TzNtzsO6aKlGhy8pkxPFnSjrXZk6gjyG6WjEPo3vpK
0Dzurophqga685L4wMv5egkfFRMexBOdWJQhM1KrVBHxHKVT6r+dj3b/zPuPj1Uy
6emH5IDOJ0CbHKpJ3roHlp641kcHCSiCWqY1rFgo75Q44jAO03pfatGZlGMle9Nw
i2a8ROQorrwDzm39MXMnysSAsbVJleWb4nIm6uTyjxQB3JNYPWpw1Sv3jBeHnzOG
M5jKLMK78zB16QtgMy310uOY3c6RZmrhJIh0Bxh9kxYI+h5RXKn8SoEvu93zyl9i
YzyH5Mu5PIRekSDTi2IonnliYVl4T4y5CPgzRqDfelHjXuLhK4R7nKr7z1TvgigA
+ogG7VRhgEoB/CTarNznVZo/ePW/K7LqEKS8VaJM0xT1C+bUjJ7yKCvNannjFcFG
bQjy7vu8rV0P12g/a9A13FDEaWOqZaFqJK5urQp5UgKKSF7IARopA4X2Tz2TCnM3
8fxQ+hOR2cGr6IcEz/ai4sal12nZiAFJRQe1zb/WZ7h5USoTDu+hytVG5guj6b1m
Z2KhcnaYjp+HD4RaVWd56POqw9hygsfYPJrEBiOfasnGS/zXkJB8tANrsOIbR/m5
Rj85lHD5V4ytgC304btkZm3hQ0Tb3OCQu8DWfe3GbLw7cShCBCYhgturSsX/jGN+
XaXVAKf9TWEEDmTHgMl73x4CL8aiFK40UboOukpIk7y4KjiLxrGCNGxfedKctJGk
hg5wznE3j8F6jN7JYJA5aN0c8Tl8P3uHxbSXm/GC6gAa/z0sdLTQO+L3JR6YBN2N
rvCo0/qF/0+3bHdgI9n3J7mNQFmbiBHYLqWUw3t1VBSKF5TsB4mwDhOpZ6Y9Nxpn
WWUog10ocI6D0zNX2ShW9y/0cfHBkwBDKdEqWuN4YjXDK7AcGECLujK23Rldmp/6
QOO9ynQFIHq9xcpnNV8R1CeqplbCxctUO59Xif20zmQAZlTeity4r7EFOeFxKqv4
6EXhEQbSQ7pjIZpcjP88yIHJ7DV7nM8hE81Erh5FQjmiBFuOCgfY4tu6XXyMvusH
cMwibILkW3nbky8GFEgMbr61rQAmUotBVBfMMAberdC1MK5r3duQHFOSbtxyWeLP
hwTWh5o5bm4THIq22g8zUQipAMhbSX579re0HuS31KWbGk5YevxHxkhacqrGYKNp
KvUNzlewk3SRLW3ZtqB4MWvQFi4rqEaPzS38q27XrJZjDb6XUsVE/Gn1VJrMBd5S
OpbcDMtoG9dfgYWLUDhrZ0KEcmdnx/oRcKBjsoH4HDR7vKSxsL8GrqG3ff1kpKPZ
+Jh2Nn6jrU90NwFFrQNBVs+CNstsuYkHoSIu5cjEsOqXiGqlhZ6lqfonevMDrmsP
nn6tr52wTuawCTg4uiKQtFbMaBWHVrhln/Wo769/YMJ2Zh2uzBsRLPYs9pmt9UR4
W/TKSdmNI2vfNHHjLgvZ602svXsGk3VmNOoaBjKnAVbV5vpXgk5u9knlA+3/3Tst
Kjw7P95j5asYOs/Cr063yQGpEqGevt3ecKGdnEggGD5Dap3dAI1bRjB9H6bbuCZ5
K39Ll9XOi2c8kMa1wFvgghFZl4X5Ijz7wipCXUsouvMnIxj2WIiYGui/hm2LM3JG
xQCBUFgGyhZ/iPKPP9lGdb2H8UcZtUAF8QVCFELCtlQe0IBwbJFOZNVs0ozNW9DU
7DrfMYQUBJTg+EnXvullES0SeFOxQRHz/xN2YVHrr2Nc2d5bptiZ3fUHCq/pxhOQ
BJcflfM254qeqxbyv3DdM17oJZC3AnR48MRviq4kdEhjLhUi39gEhdjHQyclUq4m
17QyM1MbLN2nZhvZ9SSKXT3nt4NEyrQqeyYghhyS5LVLWhpXMWubTYjrAWam0kKF
EVFEQkCHnc0SMXczeyvOonRgt4rwp8DH2Se4TFYMDCpobmZZ/YJFqsQxqsqrQQFW
0vLWjEfJApiYQGvXiI3flvMIM33KGW7kKFpg7z2IuqOAQGIEtFTe0moOj4dcKGVC
drIKMSIxLpsyHV11YV1G6kXU/fzeRO6WHgutGygEKG2T2eu7khf4muteG7sQyUUr
UfLzcL49bMH2UqpbRTLVkJTJcA/memmpA8WRkhQv8EWS02lDjeyXZYveH2Cf3zCT
lC0eUfNWLsuriun972mU/JyKWDF30KcK2ZsCgr51Ovo6mR3TUPtsE2xiqH4vWhPj
D+Z3akhRo+YF1b1+zOeVuY4x5Ht32UjGBJVhsde3mfK6lpsmZ8BVg3bTHeG8yWe0
qb00NSmfAhvqkwunxfjpWt9hLC+RGhfMXxSteHt+QLhSOceTHBsa7rfnNHoIQFDi
qi8gxAjjq1Jiol8JF9f0k9RcK9TaEVGR6+w8Ro3JKFKMHHvNl/9hC54vyyuzJbVh
hyCDs9nmnJuKKi1nWVt54lOBVs13F6PnJ5tFMpJDsSBqoUi2lXW+dc+9bp/glAsS
S0gZyD+h9RAT4nRsV4+zBLCaUG5N9S5wrsbBIjBpr49swWlOJmSBRpLDJmaCwbJH
CS5+XPOXQvcF1Bd6Yw7cPWV4EPSf75FXlBbKFdK77UMmlrhXlauJ06FGY24qFwpy
NGL1NBYhcEx1UUimzFvLXDJE1Poqt98m6vfEE6ljSnXM+mKtJ9DOQK+M6S4TZxcL
88cINwXNBdJ81kTVmlC2gXChw/G18WcWSZPK37sziIqwf8fPA366CIhAQ/0v7ufU
dMKPFDk0NiOWM8fCX8yDTb1agP1xxIJJVDGdm2EICXv163/r0cgK0ooaUgNMilSw
Xo5G83z0ukCNPTtmlDnuucEmhEaQxe+wOAyblllzUDtygboWz3MMyMOaR7meXmMo
Lh3amO+TVPk0pgAJy+L8NyxOE+pAUlhTkhlN3JJ+V6yKCUpwFVxkSxRkU2ZBxcj2
gaHPSJA8tud4je0tFK4HNkI2GwYaCB8MIDesAS+40rLfiZLfqhJfLixK2I6/ppJN
8A2mN4cZUp7MNjQLvAS8PMaB5f8LZ9yqEIPczAaldbtLG8S17noujhyi8MOjZ00K
6sUCuoSWIGCnPeLU9HR9S1WdhBGU7AvgkD2sWK+NyEF62ECVJ1HZDM0CK3/ivmIQ
/1XFcmeKrSu/EME3wb6//NlhtusxTF8QjyIgYci2iz7r0vayLHJL4dCfZIEYYEY2
TNVZOxW5aUyoIyj28v2Iuqk9tDTUrrClTvFECDTzvFhxFGM57xZsEm7eKF4lzQEK
Xj+uOZv/F19ljI33V1KAw0X7jauTi0ZVSXh0vE2rtk3PrMegh+hiIXYSbQTCro4H
lhlDq2McOrdMDeRQnZGOVQJkzqd8G9wLzLmiULqb+JbsPwdkFCkT8OpzG6y/XD5y
4Arrph5pGYplGtiJog+0gntCcQymh09oL8AC2cFJChSJaZ3h10XZLsDAcai4Md3g
Kz1mGqu41OcyiQpOHB8+vlMHsA/3D0mnZbJylwFaX3lT12p9DcZ0/a5ARf/oPmgz
fN/OgyLKWPac0JiMpyDNg6MF67EQGnHI+/aL42fGTRgHB3K5rp8I4LKrIqCulIOl
XS7I7KfcmqFDiuSWoP1GAd+PDiAxhPbUe61TpKhOnDmQUnYobbdRE6OC+kdbxuRq
7YTlgAl2eyfJJKX3GlA+xJ/lzhVqvWoGM3Zjpa0EeXCWGCbXt0RsYIUnzgo+LRE+
egfi9UIIPdoXYdA3vNZlidQfPF4Joe49jfxyk6JQ8QXTh80QDqzs0V6DY0MZwbnj
s1M/3HkrVb6WR6RC4hUmSOI89TQBxhaGX7oCIgHqW/1yW0nK5kUTZJ4Tq02IWfY4
DELgFfYLT/2O81TQJENI01gld5D+UrpCbT/hA+SIxly8P4H/4kpL3QcCzyxHrCnA
gb59S6MNIOczBJofhaZYzhZgbVo2yRNefQRA8qjJJsKDAW3RU8okVTrctNwxmhho
T+2U+189H96J8kLPqWiztYI+xzS3vLpbtAF5O7EheYZm8BUUt4ppTtUrAAScQO2A
0ScClqFF4BLMZKRb11NlxWijknxyRw9yIaGYXSFvQ/SmNWwlR/Ap9x9ZSPjCxuZ2
MZ9TOTBZoCyVubK39Gjf2jir+2YOzwCHT6Ii9IZEouQ+nYxE+f4UBdYywgyqg7AS
v+rIwBbQ1L8KTt4z2+ZdyvMyw4xDVA8BlhtSBWG3GpMbATgGFMdgkNYeDcY8PQQO
nyHJwbtGPz0B4QepSxV+P+y1G5BZ8HPuTburNZlL0NB7K2CwuThk8k8PUmB+MhVA
k3/l1scPOSrosxuY8BUGQsZ0gn0SpyfnOOoTk5OYfXLXmU+5XDsFP/DYD9Kndrwt
3tS1ysW+wumyEbldVt6trJi5JkFFLf19+ybbUAELb1IwUIswM+WPecXGHmcngZNL
bSsQoUlJEq5/P1L96dA/boUsMNQDp9aU9QbZzoR/jyNvuBKNMeKjANmWnQ6iZDq8
b2/Vy8kLMq5Xgw8gEXzjO44rgagUSH8uNjxLyIwtw/xWoXZnQMxMqAKABv1nEywE
kpgodtPi4f2Y6D6W8xM5HhmsLjqj39GXbCRJI0Tq0E/EbBRHAOrkNU5totzoCEye
47Yc8ddvlp5rKE65485G7ah6idvLm2h9je6KXCvkfXCc1xTsqmWUOf2RVbFTF2Z6
4BAYEi3gEKFk8/xSSMqSgYoqsvMgJr4yz1vQKvxqe++VEnKf0rlhJiDblccgOMl1
541gJtSbaqmB74eC4GX69DOID7ZZZ+LX/pFA/q8pSMEPXu7B/Zc+Ez9bou/fYXyY
8BQ2tguQ9t64ehnJ/nZHoTmd8ZdeUaf0qWKespcDdi4Pl4zH26Y6k2++SKWGIIxD
nK5lo/ac1DOHj9gv763rfMA50+1BhpmmffcZtEOQLcWinjzJ6bLEfokBt/SPckra
pFOaUOmLmdb4HacjCh3BPpy0q9lWzBQ99VENMXOFgS0hVmxtRVNHdbb6ErxPDBbF
rINtMnYyyvzytFCZ56OOKscCwgL/26uJ2PsHaOKBjpq4jmfJOuEdzc1TCeXR9P6O
mbHhCTcfvfj+nxHODpDiNtigrtQircP7coQTVzGWSFILfkoxjUk9FdZfxCxkpBI/
hvLhvYHn/I2yfj4l/Q9xBAwsZ44oiwWinMF13wMBJ7b+JoIM0YmklBMpMFqiL2wZ
A1/YhuMySLIUcykzrSvjDFZzfRW8rjTGQ+fU8L0W842FDi5sZ6L4AQ/pbS3aqvOh
PvFbGOM1HdoE64XudGssIz6csQjmnQGs93QVuLz7lt0idc3C2jc38YjGWNJzVW1N
uCCa1esEcsWMyyd0IESuuijMJkJM21fRqYmlXUZldrOI0e7CLu+esOKaYjSrtZGL
XcsgLM0vTlT9WRwuODVJvhsAGQ7zsvwJSojtBrILyWIRKGo8eoHqZxF/P3rH2P6z
TL6J9da9fRADwx5orpmC25qYbGgzuzOe2h6Dh8jwmF3ekKmfYSed+INDKegGgT9a
anV6PLJBJQ09W1lxWcxvjBg19BkZE9qF4zrbn2vQ9zEjrxZG8TpCR7ccGHwUANkw
1X3ocnt2NCBpVYxSHGlTOKvzKJl2U72WuiL//aIyo2SayAYqme8/rh59nFFWSq6p
dR76A9TpQnqdnOzOAB3WA83ROr+KeoGJ0Mri/SVIiaHuA//f0U4uoo7iqwdtHmKM
+PKRHhlpAHDJ984Ur53aAKPkUhsWRMLN6PqtVzvKjmZRAiYWgdc/53yIPnTZbNcx
nF1roz9Ckyu/cZLF+0C3J+LK/8SljCPWRPWFi66FP0JWcX+t7F274ix4HjFsTvBk
6IFpbevOF6epy7eUvoPwv9zW8Whg+PaaCiVSvrSlQpZLX/C++ec9l7ArS6ND5mZM
zz2sgi2x5kFT8TZUXIHVAwbzwAUOS4GgQGHMJ0pvSb4sG5xUcf0RpLDbC6t4Dit8
uxwhL6pCnmTk0TIVuYne4VO1T4ZyfmAutH/dDH6i7IdT/lxewiu1/4ni3IhJWTnA
rz6YLBPMjHWZexpYFshw4KvmWLdPEcXfKuUH9dBzroKcW+dDJmGfUgwq41Cvz4/J
141XYgXmVExkru9bOlwWqEyjU+F67wnmqmzihaKIv7ohVPpiRBBA5Psya2MjVIgj
+0P2/6shAomyOQZ17pcVOpX7MrooFJL1UUzXdBpDhOck4kBfNP9r9rgMCgruw6K1
D5fS8WeJLCRL3+7JzwiXdRXSkMi2hTHa/gleFCpcAje9408AYP+dbTZKBECEYdVS
l7Qb0cCHTcmbAePJRNB+dc4q5EMZZUrxblyEhGczfBATATdlGowslyUv5aPE58k7
Tq5wdfeflOf937lehmO+2s+fpuPjAa6FpFnBtd1ERWB4RC1bX5Jo/wbZP/Mz+o87
lKwud+cxLZ0UbRL8gaUKg6DgDu9Oq9MTKjB9XjC7idZ6DUOpy/s4L/BOhnB9oUKE
WRyqvQyGaUDsEOtAQ1l32i9eYvjOS0Qr2Iu9APEI4Gf8jWFc2SW1BGGcRvCU/X5G
Z2/MWLQD/jHam0J1aPKdFldfdfU/96alihsqrcK6D7qVXPMjSIFIZbrWYM1A5vmX
GrYu/y9ZYG8euUUIaffffJN+TYJUeMx2lXKrkX29v3ntrsVMjtlNzbpC+mIfuPUr
FjfGJ4iEZs+isN16v670MQ94iMZ3XK/OTi7ChwJUlnZTLTNrGfhme6gF2vJg2gqs
UdMlhvhWlbT4N3hyJfq4+OX5jOwYma71ln68zITk8tMui4oCKXLqMhv4dkP13sPy
qAhKycGZk+kld/wTnKkOfrqnCY8UKbBDq9//9IFPubl5jzo5eNJCiS62xT6mkRQj
e7F5IMtTrD+WRJ2S6Nd+xh4jen+TWB/Up3+xQRPxSWv510KBnsD7A5NTlI0v1or+
BRBlj3230J6JF09mqEXOpAX+/7tKLaF1baTXKvxQkfpz+BtiyUGdYtu7m2R92cOn
KHkS3wsB270xC9/kv4pKSx0ZMVpLGl2vEJ9p8hZYIACfS6b4cczIisCx4s1bc8YR
3fBXo8gzLTF9H7+WJOYBBzryiu9RtLnGsMYk8g65Q5B9S9Gzcd4gK76uj40pISmM
TANCOTp9sMf1RBCBSxS3ZqcyVX8z7VNKuukJKRFa4buJIORzjfD0ahgznaicnTVe
xvCd8qS9lF6FP6Us2rstqcuaJ+bnLMuH0C+PNDgfURULKzLj8ETl1MyISrJvyS+C
5N5xTCLvM0NcvGWvQs1txuc2OMXh1QlBvOOmTgTuDxCyyOy1DjAgR1tIwlxdkhE0
dmUt6eBB0LwShgtHRhL5mu93XBwgPYpa0FcNMQ7UO00rDqV1oTCJyYv83OkOEzkU
5rw8MJjPkm+swT49RANW7UxwSX1YwXUn5c5Fi3MMHeoLb53qkH29SyLrnREc+NiD
05V1SxP9QyxSnhvV1413IEiFeiWrVHKqVkiNvabndzw19b2CdWCdi0CbV1evABOt
M+cSlKbIIJ5kemgzgo0ZuOZ2kpi64dU6K2xqrmoTfIX73Eo/SEBHlbpGQZjyFhiU
lCPwq8GDwSra/kf6N6/BMwNYEZ1BI1Yjr9K/kzoxa6Svldk2xJAApVRyIGWXsyPM
EOsqJlRj7znp7yPTIQ2hAlNiHxlUU0nkErSFIwk3p6kOPhAzrv05ASZ447ZJvLr1
Y+pOWwdyFSzR/zD9RBm9SyEBVhHRemGr2APoLB+RCP8RG2KzVlsFnYRi4Gr6mDVk
jTA+sFmEp+R6IeZker6YYhEPHE8Ec7EIOn3XmPgkfrtNCcx8R/NFOsJ7RdqvYjmp
vmoP8zNOHWFgv9KqDvo6NXtKr7D0dz646Vo4+NAsFbI/3YT2RuNun19sAmLwvVzI
NsQryG3PzWhOtvrc//i+9//3kgizA6b9T1zrC1geSLiJSeLHQaJEYIreIeEUTEdv
WIxjjVHGiShECCqv+ANl16CCb9vntXuqYA7Hp1F5v1kyDBZ+yrtSh+j+8lGPt4Zt
IDyi1xawxFYp5CpsAOjzHr955G5FXJG6YB7+82KfUttlPp9v2n8AhBPHrR0bMWLY
UR7ayzh9Fgm6wRsKjq0J06b7Xa4AeBbBZFjCMwukpKQ9kp+fvTabVCcZ6bVzkpjw
G0E+2sR+i3zV8aoEyLV/1ye1Woo4Dwr6N3AKPt+gDZ2U4B0NlGP3gXyKDQ5KjfMV
C9DJZMNlPKOy9quxPR6zLqAUhUvAfqv38JF3mXJci//mAg3eUfY/mEkig5PuO7Zp
UekaFgq0VaVpI+GDGduE1a8Zz1e6Y3AZq4/YGL9aTJXPCb1qJ6W73JirlIh568jM
pVT5+fIqdcuoUZX/yN46d2NQceInOcWBrO1ffBk6SXerPd8FPMBipRybN+VeRtDw
sMprt0B3US4ayUD/iwSzVL7gg026KqvxLW7krIpaCq96KwLRKM+QhGuTfNHpu1iZ
SQ+JizM+mEt8/6bXNuz/wH7UZLWgoEPdReV12iUU7hGNCDfuBS+WOEcTpYBAfNPc
uKZgIeI4NalPzfo2HUe9IeD4MpX5Phf4z5pR8RoU8Vs1no4sjkGI7Lm+katzJdEP
TGDSIcIBrHNxi7qislaoihuSuFBlNxagtcp6fI9lQe4FRU+kzM7HSpzTKnTpybba
0RpwN6xOl5ebpoBzTIColVOiD5ynvjSEI3j82tX7qZh7U5AEQC2ZlvsOOKqE6hHB
lhijTY95UvlfXxLYR3+t8NunPM+/igNT2OxrQVsdIqFHHZxJLEsymwX2JOvR8z89
1VZWEVMBZR6O3bpFJjL+uxvQjfRqLVhb6MbfQwHQNYPMAIIA9ie2f2V/3FK4TpCc
yWx2eeWwKPO28AZ6EGWk6N7t6rJ6TZ+inWjcEAYvZUpOZSWV9PmybYhodhtH+/b3
p4X7yUJJzS6I7y2mI4r+jyplczQWPqN71RJv/pRNR0TureMSfysJUkf4XoTAe4q5
a+f7LsYPju/2rQP2tTsxZH7BjzofTpQVLrNG8TWhcWPpK0yAziDTBAyX0vk6YXTi
6LORTm1scAsTKUWsZmNly45rhPckATjuYtjZjgX5+pWuFGfLe5nTXBX8MymVwWVJ
wDG0gQzl9xxZuORGD2nwHk0DSwSkitAOJMhtd2Nn/MY05W8aCaAzO62A0ACSik8l
VAyqDuCX31GjJHBeZR8MkLYbdCYOiyPXuti0/Y5ZI+WoX4zj6agckY0IDU1uU/eW
+Uc9JpRhzh5S5TNfQpsKGyx5bHnbEqzkQNIjmUw6sOnGavQ+4OepsipxspVcHC7I
vq5gYsTzmvl4E/IBI2zKVKmfqIjUf8Y8oLHdYThOohjvsFHpsQb5xhrWzIsKlox/
Oy2GlGLfTh5VHMccdt3jbqpx7Fe414u3aaudpVUZPA+FRcfdh8XYPNNxTiwIKfyq
HqB1ZSzhmbIKQzR15o8WaUQpaDyufGKz1prCSO65mlL3uAgXlSamSOPlk1SJV9yW
XPPQ2P1KMVFeuvg3TDVnqH+ob/1W/Ch1wfIwFyryf8cIlKsYhvCgkLHo7mdXMMuG
2+aLYFmxHeyrMhfBpDJlxUE/OzgxOVdlJIj8AxQVG94qepSqhptqMFMP0xHLIang
eS8LY+a0ir6xmRAocgacczUZ+mrm8AcwANqBc73aXVFYAJ7Te8fWA1hjYQ2QxxDa
617a6fjecyGBJM1xXCkxty3dKU/r1dfXGzimrC3P7decfhkvSos9kEUmzAJcfzZ8
8ijxUlZ3HzEz7jC+FuneRrNIoTyz3kzbZUMyA6CrVBTzY4YKxmWDD5Cvv5qPS32v
W+muiFB717bDixq9TLCU50wdXv89WXRRNNd/Rdp7qo849jLarbsXzhnqeiLl6PP+
chphldyTEYMzyl3/0COtale3cQMig/Zf9wevpxrKB+e/VARr+JT0qtkC9/tblvcM
dgQoU294WkToryYYqrYlZ1NFdnBT5Fa9IShBlS+0ubwkXRtfW0T2b1EVjwfcmo/E
wWSDopQ4+DN9TOxILJSCuqYxEFHl3rBsRApOCx9+JIchobgkGV/LNa0/WKdB2QVD
7VdBncGNB+k4HiscKy/gsU/Ah5994UQTzG4r25Wz+eOvDO/7+tzI79AW0pdcdWuY
OjXVpBkIgYMojdwuEm9CQKZTUYYTYGNDyGomMLbTJ/KcZla3ChX0iXigEGdDYU+0
PTAc4Zg1XYtJ07PWLxb+dD6RkKd4ZbMb3skQIOzBzCbHAODbHN7RJW7ODwUxSj51
+VzV8Xx7P2GBOacgX9M66oMz4fq4lCe43Q7aaKtSW4gztDMmJ1jqN1MRJsWBbUCx
hxo/OyPUrIV/2PUdnlnSgdi9bHmbY05T3NpCsPjwpeKdJCjkjVvj4rN2uAj8lzrt
DeyXshUp2drNRRBMwo5MgG/Si5D4qYygA41TGy8d1etvuPQqiWo8GLDAilK2ZJ2v
836WCKpG8atVUAqqWo/SvgOzfYPR2ZmrkRrkjC3iUGewfvc1ig6ZrIRgUx7bMJ0Z
lZiBonl5vz3jT8qhXkFFmGPlfSMVNwxbzPdv+pv74NguMZQ/Uze2bHOapgdN82lZ
eHQEpM9Jw2vnyOvRuoH/HcON2Hle8LR14XVQln/wTwAehlXf2HgvpEO14l61fOtd
p4t/0O8dxYWAI1s54qWBTF2hUR1SPGE6EQhxOhEawIWHl3fPr4GEMGmXYD4kcjtM
LhNK0h7es15koHHwZIUJjexje/XtYuBCFxQNgKoEnUBAaBm29yf/Pk+pk+oF2kfy
+PJ+kttmqIVSvwRFB8/PWtLd7Q5Vg2URkIuSzvjv5STdVECXmmv8SprzZYd9Vfiv
zti7c75pa+gE5TLh+yIS2nv775CjPebBGUfbY2IRsbLdD+okKevyeBskeCWrr2D9
275pExmxH4D1KK1Fj+dFbKh0snkcbzJmko4F5u0+KC5VP19tNDLZmtVloaGBPtwC
7nhe6kVYBMIUTz/evEnqSZAI980dJHM8OcJxKqXkGf+Wv4sauW93Ewk7jPyzmfGZ
xBtYv4mFi00Viyj93HDTPKXHkglpE5pyCTR1lh8/VPbrcI9HS42PghCi6/gvWKUo
8TyBtsDtkHXD3g/7UfPJ/pT1F4tViT07TUmmozc1o5tK5JwOT+VIXBixqG4UKcP4
7c7IvkdK4smesO3SHZ6015C8BNTZqnD/bVuheOCoLyxUUH57txUhcTZrEOIn5GlJ
NByWoMNJL7KbNes9Iap9nTXNUHrZU+i3YNH4ZB4eF/00Gi077RPLOSu5ZOtUbWLN
2W4qAII3iwtvzi90iy2/1I7RuIkCiyOTdaGfjJhCb1V30yzcMPoT6tlzX8kaFeOD
a/NTGK0tPXV5KLlR6EfqnZ37FwXl26fDLS07/MGlwzS36suuPRESs6teCuN+QHDv
oCn00Q1cfNbbihQ/idwf5r0nMU6LjvPgYyDVE171LxmtmWx9dtDSS/TYpjjzrF71
+xSfzPtAZ9u5MZYwX5g3yJSvt/HPiri6MdQrlYTuBGcIavpSZCdy63Hq6ljTjvlt
XDr318qOzBQrVnwlNXyUNv2Or6gEra5zqpSGnPtmfei+y7X5Y23lr56Xr1qR6ZE4
Fu91ssIQbKNcq5T2XGxxqMzVASjy0npGOnnFgWtFXXDd8XK/eJ22iF0G8gDhJoSF
OD8SwLt9fTEGMCo871kWUJyS6y41yRcGVzd0+FMF5b9WEPFd+D4/rLHT0p9zsKLb
sCgrztB4W/B2anosugck8v4QGQ0suMmJl3h2nJdY3uvzUqpDOzJJPakWFhZ+HI35
UD0UfkYjV4lfgsjCt+Eb5gPETEKKoQIXk0s7+k+PX44gAM7USYwYvASE23Azr/Yi
zWBwKnTyfRV5oNrItneHRRLC83vIZWJG263GBEG87EIaSWU+YtFIAtQqblaqi/ir
SrxamPycpiWZ5cp936jFkfTrK8FqXhm6g6akQkQA7fx77uOxZt+0GPZ3gqZaa+cd
jsOZ/lyUY/eL7AyyeEgNZ+lovV/HHidGYXzE8oif0iK9F3Zv1MQ6DXLmVM8gD585
HILNQcmt2LTzQmXldDcAOpNWUyK97PG7XSt85FpayqxjTePKDfZxzreYR57kZDaF
Amas9oeNDnkn6eE8t2rsFetdG0ckJsLiWKEfvA2OnWPx90NvBO1MxiK3f8K+hsnf
s793dSfd0o8NqCxUhyJKEtXDTPZCZBnsan2TWBfS4AFNp3quZx0qamMnq04eJY4L
ckEC10lWNmROh2WuB0d8cLh0BBfPswZjm2LpzOux4QDbdVWHg1WJNawkoBjIYRw0
ufeBZhNQva9Y3rDrvunZtsZNrrMBFz0PoEcNeQevuLXHb9MD6JTlb4Udz4TuH9Yl
nqsakzQA7idVGfqlfW7h3MwPI8roBHbmt7L+T5/4UKsxIkp0OMQXhzr+SfZ0Q+WU
oiLPp1llXDOcuX/kEHYrr3WeMQ+560pc4mr1kARFEbgeZGvGoQCpn74Pf4hW0+bR
UOh2ECqgUuQGkvnyx2/WGOQttQEl0xYoglFx/Vui1qDqUf3/Yr/iQgwnG05xFGOF
A1NilhtWm5D7WmviBgRxh8KXVjCe9zs70OxJjiZI8zzyX6rQSoQANldjDTiPBKH0
qHXUztfu59wBqrAQ/WHwaP0Vf4ihE0LT7MmsheSdibuxzmOu3cf/jkUfz18UlSEl
pHA0HDVyNTPWeJaBI0GEWWgmUfEmwm8C6w41EZm9KcSRXkyABWZjEdfbWtkCdK6x
zYnu5sKBfhwHJk8OspL+lja8MXQR3d8K37SfrjpBqYAxxXv7csUhSRAS8vVbJzQK
dYryMwgdanS5lLZuYoHrLfureP+ZlMV+uykYXzidgS3eSkcj6Mh2vrU4UHYakjYv
sfQtGbjkKrAPahY5815z+FsIHx2m7pCIzMKD/YQ5doVfWIRXsWS6KCPJVlNjBKU9
+U43ZdL8gZ2SsJGeGu856eLkBDZSexyv+8x9gPdWpBFlTQoTqmEZ5YYYDvbbnrx0
8GrWCEmsAMs+J6xUzVEd9dzDY8smGzOGYi+gWqTHpI9WymZ8juTW4ax0F11kfwQa
Mc5gjPqDRHynYBuoBA1TAoXyJ3aFTjpsViidC5xH0OkOz4tV3hWWnSh5bPCT4VQK
rxHyoWNZTU0XDBJ73jH+AXh67PotEiuMpS1t9cam8pVkIyqYjQDzZusCYxpC5RrH
/7ar3z48/i9cF6H4y26jiGUnDxuAdA0hwMywBjBAPl4JpVaY5fXMHlJ6FlwNjDhC
7JQxQn12/r3ZVCsmhRo0iO5nCoYT36Bnnikd3J1KcvYISBwFOwFSZ4RxtEhxDIvr
a06ruJ/amXdX98BcKN0tYhZx+hJTJ9ZOjEBMhWB7YNbaBlb77t6JzE03ulXC5acV
PGmuFj30VyY4w3bAaLz/pzthN3f9YdXZ514LBy52RzXLvmCGeyF8u+C7a86T75j2
XDqW/ehMoA1hCzTa0it3v/eY+DKTvgeDjhGfWOvQgfWOC8eElTAyYVyr0WQ1WEU3
jBTqWkCTCEtKjlbm89ewaph32C2LTMM4RKv5IDJhGYK4zzePqYEaQfM6zrbAV22F
yCdPT1Qw2BiGeLucKCf8UvGg7FMted7vBQYVfYXtrvEgMpVpijaH/O7K7NduiMqV
zo5v+KWTEKPQ1IWdMaw8o+u3vUJjm6ZYwF9AAZ8HdCYAUG4RP1ypzblLwJRMs5Ac
4bObQ11yqAI1+k0UZWkvp3sXHh+ptzv7+2DktFQPXddH5tlxivk/2VoC1gtmp5BR
LBO+Zvov1ojqJtSF2aoUwWjZW0LLOmgx2cJLmdBxklzQnvx0xTtW3vI8csOaFUdm
LgRVKqmo+IzjC1sivlIJK9FS9ka3fyaWCaycVRL7zJBJW+LxgiZDYg3SPYJDLPLL
OU9puz3SPRVJ3xbVMywryYeb1mF5R7MZlRTWlXeUeHKFK+hDWfKUmAXRNFqoXvMW
9AeW7Ifn6k/QPz6F37Wvn5ZD2FbEUmdvWWS4HPLIzDau51jF/W+2bYfEIwC1SE6d
QZ0NkktOo477TCccCgk0rDbwPGk/fGzFa4waMfKTwUnanWGb+j8zmg4CLOaNG8Ys
hxo9anJMoboBJatxTnUfBe2rjTdI81183nsLYKxGxmHnvR2Kq+hdzs6qmsJz0OlQ
pJNcCH1PQXhNyj2sdPOiILGMfbBEH9Cd8N7FqokO2bEoMkuACd0XCD0wxBZ/zPFZ
0QhdHxHSpVVO/deI6N7He2QkzQvRjcM6Zgcs5BgsyURgqaxiAwoqPlU/73SNvghN
pOEhKSyepGC2MWn/Vr4NrIPsEPAZEcCs1WWC6S6/E/52q7agggDbR8mGTWi3hKq4
B7zHRYF1ldGDp8hYg1NPvDYUqWGq8f0XhGMy1rLlM7TonE+MyLvvfEd3mH3nHNNW
RB7W853Nihl0BnH3WMWTOR6hDjfj3qFaZ4bl8qKbanm7a+CPTFNjghq3yOKhiDLV
HorTwxcT1Iv4vH8/k7N44qtPKPmRxhW2FSRLBDB8s2/DIAnUOAIvEJtY/GxnqMXt
TliaTAhx2blYyIe6+yeRYTSB2A2sMdhDBZBDEjDNe+rVNdGob3yqd8ibWBbLQWEv
po3n79rncA/6voFM6MC1rLqY9PuPLIsHNETTkv9JKNoVySiF4hytjNdC8mIqIR78
RBdmrZPOkrzBqEgfQPpBspBsOe4a1sgbZDEo9AHl9j17vSQHMiNVfFX7db59P+/d
tiMzMyeQKVXw2YMAHK+42EDGSl2zJ6JZf2FZE1SxTN7t8IqLLwItfCztwwxZltxi
MgUhkrFBb5FF05rerB9CbYOdUlDBcdquHehAhr81/lPBe+EXi/G6b+qUxTiMABZW
5LR9pGP4BPozlyd8ZuKD34S7iTDKxMt+1b3JJymoWv+ut2rjHwlDgtaCtSf1jxcP
F6NrT7fXyYgAnuArzrLeELhtN0xyJSruDdD/ABDzEYIpenHrOE7eHS+GbYYFAesD
sMsxt3eWQfX6/13xYFuZ5mVBXzzTiFvj8VT3VHDfPDYDOKdyBP04ZEJ2TSP5EvWE
SgafE6qMZkDF/hJD3R1TL7JPVcfBLPkKnmUXHezFE0pLwbF/byb9EgGXR5Kmp+HS
eSY8j8GcKv5jKO3/E+/ejvZwj28tPL4f9HbQbKIaQTgn6fBLZVW59M27vXVoyyBx
AFicYy6BUwofrtwLkZzfTNiFftqZ7BLvHT+zuRufEDvzifY9jexZX6CQNpTgGh8u
jP7RFwXX8lSUTqUp0TiP6cbSwLrQ+53RZovAM/dKfmZNw/RwyiPbcEqTFDblIqJO
IeDK+djja7w/GGkfOSnMidd7qqOftRpMK9RYA7S1kAwhXTtgJy6zJxJSfCzmHcol
BnD6w+0sPDYGLUpaCSVt5nS/3Pz27nhJgzbnc/FqyLQs056qicjhm/5ODY8w/G6c
xAZ1gdjxQVspD0owBp4uowFrYhMCHe2OgDACSc73b0LFHXH6xSI8afHosWyuDQKW
LZ3HBjA6ow7I1VkQndoVoMk2+AAfznMjtPbwi9VWRSX3l94nQmVSKdOJr7S5ZVrN
+fkuJGxkeJWllv4YUfGvtvXYqR1cPI6iyEfTX/wTHuK5YxX+xgXFZ+QfB1x1jKTC
vfezAs6vGhdaxCSa5QP8BnZgbDFrzLPE1iLwZxTm9ORkY2blgtVQYS66c6RxbM6G
lozkgdx1k6f02/Ilyw1JXrwZi2FUQMEEkOXVj52aNwBx22vR3gnbyoZNOWhRYjip
a8UH0+UzQo81vpFUiSedtoSL+eD9rBvrR2O16E3q4zsFLEUGquDlASi0MNo3dM8Y
Q1TLPKmCEhskGhDSL4+cRt2I80QCOSTORKoZm1xR3CH9FsBJmg69fAzIuveLGYlF
S4fSJvVREEjYD0QBJuftRwjh1mq7kzAuyHOoY8xpGiATAXF47XBukmIA4xuPLFpa
ll9oNvF8p75pknFOLDOsYkuCMsWeNx7LfbKZsZY91lxvfzEo7jo4I64TM3UagkOV
QRA9YpIZKPZzZeV6tHscSPvldpHI+Fk5d7snX+iCejWUc7nVcPJj1/ToSLMVeonz
tlbGLBgJuG+BhFSGBau/25SK9jSpWR9TPTOD03MC+fEUbqbEjrv2YmHlaZONksHx
mcjdonZaHG/X7PU55403S3tBSKA1CKiCtRWg8JIiGX3vxkS60y+imu0wN/X8Mmci
8Du9iH6fS5lF6avOdsxeFihQhoNPj4mmYgJqueGUdzu8J1PupzF6LljhHS13jbk7
/2qps422TOyKT63Yvurire6x5xgEbBHNo5g0j6PqsQmFdERcx6HfRCnx1PxP24nP
XcSNTNL5JDxhz+K2C4XKxgA2PoU/8FvjCK+fNbTx2TsJwZwLyG45fdWOEXW6oqzT
1FLPaGxG/3YjjF3kbO806jQ368V0+Q0v2WOZ9ukfgcP+c6bc3zuz2/wxmRh4oma9
R9p0owV8x59T2GVXWtzYigs914G2JbyMVd/8BnjZGnkwEdyBE1I0mn+MwtowlnYq
+h4x5XUyCWUkGDz+DYdnSVdQkJjrz76eY7k/4kZMAmo4xjtdGM/SHx9P3MCIAHZO
8xBcWxsVKVVAAr5nssk1Yz8e8G/5S8/UIyYjKG7oaQW+M870DSpzwRU6rbeDWPPY
/5NJ8k/q+QgvOBwvGqeXg0Di3CbND73ZUmRFAvkir2pn01bItL05k8/+vDAErsjC
+986rTc96wvc9Ht9a1dwI2IdOcyJHxZhbhY65z1OdqnpGi4c3PrKYhMetEGEtQ2j
Cy4FHAH5mWEEuCt0RLP8lKe6HvMlsPOqTEtKOPmXl7st8vG07co1eLyEm2HJM299
ASircsRtJhTLTJuUCV22MwonHClHTSi+HTwv1zqgmLsweyVwprsLs0CY9Xc3RMJf
4gulzi6D3MRqisxV2SJd0r+CiGkC7k/CYPDSerKG9o39fSGR8vAGnKOJt7ov5RgU
/TGSuEbqt/AXwHfmkO7qZSJVrNaN0Zld840sMsXIMyvo11so/+pQ4cqWK5jtwMIr
bfZmcb/rX4lcM//i5jKzYmEFr5pJoLqtOiE0vo3/vQN5aftmX7MfvsxAK0+Iio8k
NALVLLVtoUpwviGz3EXBZOYhvog63BYFZ6Qv4cEWp/Om/ET0+PFzMgpmLuKALE64
w2WFFDuOQA4qyiBXslU+wvdug+RbIFZbHIVgBpDzvUmYTljZRQJEvazApHYQdK64
anGDoVuwR8TLP4OvQZGJ64nkwwgvtIkfkTiRK5/gkMM3fsapIsbe+0pXkVuo6N+B
irkib+up2DLCW+li6bs5S8yRrtgH3sAY1h1my5P7Qe9tOVa234kkkWqJvZ2v3ELo
XDCldrVUqKay0bf2dtbQn/aht3ReLSPUSim2T/WUiGaeVfRXaDi8auRQMLVysqQi
eGVNb+Z58cjW9F+AtYwc8j/LrrTpYtvkcJVArs/lEYGoWlnBijQyTQJclxgRV4yn
9biJs2Z88SREP+AUbCVNuRfstnDZ1zTKuJ0u6xp3EvvEBwOGbmO41iuI2qTsryBX
s943MfdW+ipYknV2f5qet6BaP/bH7hiRNJzKDLIT2fcNjUdfUXj2pmZEC5LmJifA
W1fkanhW8WCZ/BLfXFYgFdxwYt1AsTa+jZQ75SsJ3+ZjDLdBqZwrV1E7rpRc26K2
cJZhxep6kXPYTwd8ZeT8je0RZ9JsBnUKpgYnVzk2B0gVdjJ6hh8t39Cwn4gwXBcL
u2TXeM14l/NlqE3aLStOocWF5E48eEPMrmw/kup13OtcCyZpCPQ4hGMw6xIlq9Bi
RC2vcWwMrDhSmftbQRgxYyQ+gAmdMxomIlS6YLOEjx5GjUKw935FzqeNsKgrEyS6
TpRphEm2emrpB5/ZhwaBfjEpq03w12ALsOQ59Of7sUZpaNVpPxbRgGDaC/CbGr24
s/RX5NZpj8syuVn2He2pE72BwslEU/Qcr4XyMp5SKZ7Tecdx9KIPp1Io33k7OSYL
At622FAI+o9DO2zkVQJIH3L2jd2QyqgHXarXbDG9FJeocOVPW9zsFU3Po1iUpLRO
KE2yZx46aBX+O9CcDKZnYx9BaIwXimCq/Lu/J5dpQzMWjJ0jm/0g2NbRdysy+CET
OweM0JpW8pPViVQtVUc18X3BhwDoyYxQceEZsARcCgxfaSpX9goFprGEs1GZoqVz
QXn2koRUS1CS9RJ4kdV2WJU5eTSoZA0mZhM0q740Agx5kX3wA3FG5skwUAEKjOcs
xxdBvdUyV0t0AkcmOpxtpjTsrt1UwjQj9FTT2DKSOzcuxwM80NcntS0jmnJOJjjx
9N6G75Usb+cp3/62/V/YRkvuxmHttjNagtkEJw36dvw1jO766HSBFKeq3UW+wlGt
UVON1Mz3dYVUhREfxvcqoDxHUtwQdIC1iFvih5nRJejwUAVcBQvsoAGk7j9e3OIr
FQ2+4Ac+p6NKoB3BxmUq9YP5eHf/ikFOWpSbOSJO+skvwKzjQni6kMqxsly9OPLx
E6qN5RNHmvBajC6eOBLcU694qqNPXg1gze2nQGqHYn98fm4eC7JrJtX5drxEgkg7
90P246wYCjuVt0fc86q6RcHN+51dcSH4bnAf9gVQK13cS0Pt33UZq8XlCFvQMDwT
+kqMkVoxVf0YgvlAIue6gpR5QBzoOGNiSuPmQv1EjVXK3qdA1ghl/CDEDZy/m+Rz
fQNNfyOlbBhZFq3oC0mhywNhR7pycv00iXcoGQp3tzfr2IPvCLEqv1+rt4SR5UWS
eXCT3d+T0V1WoC2bryifvo2ichVygEDFOcZJMIjtGghehH5+fswo9umqHIyvkTGX
lnJJ36F5mr8uR4bl5mP9Tpi9mzdSmsiJfJfwXGY95n3TOqRsDMb3x7PrmjTxVhvh
ItdLWxwAv8RmL+uwi/DP2/qSkYf+PdNxLICcSk1ok7CaSGHZ69uUG7n0DzakeeXK
Cs/i6t4PsZiH3ADF3lGdS/mlhoV+Framh2ekjJCX8frYhsoAH77BZDt8z3ktttM1
Y2abpDWrDk4+SErdNuC4gSF4qyaLQgdzjYbqd2GNmyLYRJYPN4Rvy4oa4QeYabmy
bbZoHlbuP59hj9hmjc9yFbR+OgqpETy0MJQAIFg+HSH4YuVSN8ryjaHaWFhkkkX2
oao6Y8/L+a1r5SS7YCWaPNP5jhG2TzwYIxXPdB7uKSnR90cXF4/2TFogvbFQHyBS
MnDvezymG8Tc7FR9setQy5TZ00I2ktdMGlMOa1EgfxZNnP9YQEf/BB92c7M3ivei
lbi/qV35mPG21WU6E7VYfw4w2TirGXA8Hu5Yfn2Q/FDLyW1WQMd0aIcurr3xdxdl
bHRoXk05TWyjhdlJkM06ht+a26x/JTrzN+wS/NfWDp4xie9J6iI6ACZ0NxwWP24q
QbJ4S+qufVU1XYo1CjVh9BO1eRkR/yfwy/Y7Qnj9u2KE6Br8eUu/lNh9FppanF49
9/jQJeOMBZV7U5l03QsjhPwAN8apIUGEVy5Zai2BWizwhCFgdJASBLRJcbPj+K/t
F93KtTgNt61IZIFr+ndSEtW08stviHe8w48dGu4mRoA8aWubYbGpS49M4BMMkFzW
V5YBCfCgd00WPKM+RLQum5XNrkW+1NnIjxeNgzW3YVg/pHHMWleSx/ao3wKsRZe3
LFrjnTSe51rgW1tZETPE1hRQk0WQM+x3U7g8zfZWV8ND34CojOtXKj7huxGu4Mk4
C0bQ4lzw5+MoXGTH+Ho2Goiu6Xuc9t2jQfbgojtq2Kiija+QOCW4G5nfY8+nFbFy
oN8UGn1uA1lOMfwOKoVVdb8guFZX28tXIZ8uHRDWy/ofcm/PB7CgMqEL57DfFGRe
esoqN4ms5XygHHJXqx0H8lhgJTgay8b3qQVWnsWq9U6DW1+TASbtLrXxMwYEE19x
9hcQN7nH+NcXFQxOW5exmaQ9re0zLbFjwZ2le7qkpr0dcqN5VtAeDpPNU5HRccys
RYPEUwwtrXs/wRg0K0CicJLQgjVTkeLJrwZ5pxPb8stuiQXiWwO+Q/AJJifuR5VL
lFAzdv5v8W/yZHYJhQudqaJVZgb67ZN4NMvnE3yWm9vqd9n8i6GmvblMRwRElQgF
qjBWCKFM4QFbwSPvUgbn8B916DD864PvEAZkBsCS2Dtb3SQun8Dl8aI9QomRRBW3
ryl8EtTmvh+phr6ncwtlwCJ5asdm+brsLkbtwBgxCt36Ar0QTxMd4agMfxLQ4jKj
drGt8gAV67pI2gjGyufjycwfuozN78gKUau9JBpl39Jf9KzwPGTAHp8zADQ9Scpv
Ekj++1C8Uw7VaSeIn711agqyAHfIBfcHEhOMhkKkUv48TKAeKyACVi/DsCH/OL3a
+K0iaj3pMM4GEu5qoGuUpwdtYQwjkGAysX3BnZZ7L+l2OGsIREIscCO1BvRaw2Ap
xXu9Ekg1WSmrm6SB59MsAjW1xU+Xoea5UGpE/cjbH32pez3hGz9zQs9lR9nN4PoI
PP+cth2jJWWwC2h5KkJxWPgGby0ZV1EoWjkKkvNA5bc1OhkeX/667szjl5copfG6
1gMh3z1O7pmV/19YYEO0Eear8sVISH1Xk4I1sk1IF/eyaGxO/t0gA3iYfTlgHS6W
lI7xO35Za1w0BGnnlgikZkXZJVLO/qoJBzHTekfhJ73ptIqhHbRBWooOGSykVRTr
t0F9lyHvamXnJaHkLSgRg5Lje/Dw5BCATTJYsKiLJPd6YsW8VNGaxvVuZj+eCnRv
Pm2Ilb1Bf/r6t5JOtwKYyDNmuTEowFwP2oPANn/6eOmVt/bN3/0nuCi9nMqFCKwI
xOQaBHZ2naTtPyhGoRyzjAs7/BxAHG9hXga0aeLAlrceaHGU1I0gfWmuxwiW8Xlc
rL3PKwyejMMvEtM3GVnXOnIs3GpG4GYcijKU5v8jp54ZqPwOw5BlPDUGlFBrOqvP
qJmZNZ3V+tM0WUiVmiBUPBhw1lgRxSm2FhLOHUvJjU/wq4LZKu+b0BVGQ8TIrPti
jCVw7M0rWdPfVfagu+zEGMERA5/lSOdr0dS/42SQVCw+sqrmzDude9+OXyHVDw/Y
x8WjhgPGjO1O9UlI2V9duRgiT40ErXsJJRezyd19LEIqGwMEtgPA2C+LALduKE46
fa0Bqj3ScSQPbz1hy4OXQ88IVbuRhYidRTDC2+gBbvmE8Ya/G8ArLVO01EVzmbAu
vFkr3aPrpNGbNbx/w4dep2nwVjocZKaHNg88yevMre+YWSZvpEkIE/Cqsrob5Owz
t+ruVIJvKbiDuXRtOgj0b4BDpVm6tRdgecpgjUcazFIOt5j6YXAMIW0UBN9ZtTL7
VMYSQJUsAiui66nZ5ABu4SSTswWTh7xg94/x/w0cu2ZaOVNJqOSnNe8kqMMdR60X
d7xEPDc0KfoMHoX4UrJzmjOs7o0nB1taCND/iyYQ9GcKLOldzvcC1n5cxS/IhOMq
TQKdWi8thDvb9y6jyIBwYr5J4MDWJL7B62bDbBD3KMdSgaax1wLOyPmR9WB8xXyl
xjrDqqiRPQL8RLGu9kvJKe5gv4JBMGNHbiX9dUzntMEi5WRHGkxkG0vCeQ6KdE76
DTzhFAAJ0yyd2olQIWtqqwKdvnblXOH0NnZGSo39Dbo8bSIUD/SzsK2y3M6x+v6N
TjVn/4H1Jt3J1b/SPf/wmHLWLpFY6Wc8tA3//VNXHnIP153WO1yA93PtGN5Iql/5
4MQEolBr90vW4qqsdOTggn/+GUlCgc9rNHohPcmyVAjsLt8Fhioieo25XLlF8nV7
GC+pMb3FiaHSfPkhIiCyqyfPrgO8JQ3vkoNTiDd1+ewiGA5NsVNJu4DoPHl+1Uiv
oPPJ8jLcWQ7cKq0B3qY2DKBZjDFRXe9cSCCeQSv2iVOYrwtmRa3mRxSz8vAg7xN2
QUFwktLr24E7eFB4Y4qdstRtQLN4LdcfMyKFKpBVnrpOILQr6g5tl05iFNIY/Yai
iH0PFB/H68nGmL1cx9RB/k2kc/RSnP+X/ghGwQMEQ0jIV4hnhTLRuJE45xe1DP8Y
FAS6u3RuMo2Vo/Ivjmb9joITDGAZUa137DfpoMklbF5vjeKvckmZqevinZn9+JWT
C9cxPAFthGCydf1gwqoDgjdvfWVR8Ffw1Td2KEamhQ8BdxYCkMWBytPoW9tARq5y
luleJrTpjlJmmMZOy+eVAuJq+xN7mYBkOOfx3xrwca2SIyLV2RYkSPaDoNbUdecm
aLia2/K9EG+y4jTkdgrAk3mmzYaLxp2rOOvjelvSY+xgPvAoSHU/zQt1CTjWj+Un
wMmiojdSg19Bom4Zfp7KCmJqSkvjxRlqJlZ03evZArTggcMNeNWiB8mxNBZlJFoh
CMy9su3znJtgItBGqfProW+8Jj17iYxfiC/NCjgXQwglFVOMKXm7SGTtE1VrR0c0
tBgU7fLXLYbj/0cyAeEZ5bQ/gsvvl1lZO6n8wW7qApWr0z9wt+KfuCECeUQKykPK
MlLU+SaXF4its0h4XkimFZ4HgE2tATPZUkAGUyZWNmNYoahuXv2qloz5/0Aml1f7
mavUkcNJxyAJvvebyy6b2whulSGU2f2Eoho/d31skrV7GcbbAA2ngFLaqTr67FuL
4trDblO2XmEUiJs3VT3Tag2KaV0hz7z4egV4Ys2Vq+bW1JkzaQA0pMyYE6WW4Fhv
b9vr4iEWtOq/agupRUUWF7J2/fm7TgrTt4x0bGHoANcEhVUopDTd+Envp/cwDpDX
8dtVxNgEyM6KctxSGG1/xM/dsCYUY7lEIoiHkf37ap3IncIfNtifLXlnC5BzaBug
d5G0aRi67qpHTr8fNGNPu8h0/TnWNwI865Ni8aLnBzWRPSYSOonHgkjAJidFO4Jq
Jf3dwjr3ilAKFZGiqyrczUzRHT1v2sgaXmjSLGdbYLekPrX7N2TODEtuuoMVO2Uc
09SYARHZ1lZ5iQoMcej9yjAa3pMRLQwe+SKtPAPl/evoHpsOCIu4vMxkie1tBDYA
AzQ5Q28deySjuudiUjde7o0w4D6n52EEPsPoULeEFas/BOckkzu7nQC166HOd4QR
X+5uDe9UvlI+1L6sI/4oBLoFspBlN81CN9u5Wh/7hdczE+XNAvZW6SNWcVhKCg9D
FOmXLbRgNmcLCCX6Gc4TinghREOMC/uCOijkMEi2kdd8w0MsbJPZe+Jd2lytg2vB
OqlUfOStbcfSuhpykSxQTSafBtuk0AFs7BQv0VIVO3NtqLrpdixfX8P2E7ChNNVt
txVkeasQo2vHC0GOSkQJrHWYakAwtZxuVTHpB50DgjyOUlVNJEOritraPaOsqy6M
cB3cWfobaZON+NT2ju9ufTdhp7hQHyybPyz7i+2NeQ1B4HvekTrIhIwBiY08XZ6i
ML4ej7wKMdizG0ypISxfW0ejV+kxuUCMAU99hWCuXt7ZYx6bdstZTvDWax/OivC/
Y1g1P9ixhLSFJZwjnPQLC0e4Bme7AHgM4HVSUuDXslHPkiWQC4hq4kn3qaDQrIYX
jEoiSETxB0vqKyNB93JGU5v52L23MEzhoyGdZUZjklZ12R6ZLbuPnVJoO5zXGk7r
IooJ5Qp95YYdVz032oEQ+rq8xitZUTqi5G1w1/4+JQvEFQq7ga0epf8QAwRiV6/2
ssRuU8otERHJ7SDA41TbTBL3yQrQ8t+dZCqFoTrTSSEoxr33BijPPsKm/XWspIcc
vCpBQ+UP1LLVd7cmp4sUap5hQSUJ45qCpz2Y7qWvxSQYFrsPqRMKm+v3tLOmq3TO
pxdfSQoPgejM/W1koTomWfnFAFEELdf+zu7t55lkMTCraH5YmNherf3lSKC2P2j1
fcljOkbIHa4685UiBZr29F3s0zKGZNbajfVhMsCDKWlxGj+CVZOlkvZDQDrT+iPW
mDvbdRHO1Yxq3qSvWWZebvlatoQqXWIw899xA4r+C59Z9aJ3q5NjVvX8MKywsNd7
WzZ78A/g6fwI46/ufTKNOzSjbGwv/QbOalLdXEDyD+uDXwrFX/J7E7NN//LdFnGA
KOz+fFPiORm7yBmVXuEHqxWdYzDbPSLWBy82Dr/xVQjZvLOMioxyhSY6wA6eBiJb
yeNE5sSnZ3yJnnpaaJA2NqsT8E1id3F0jza+XIT08fj0QELAWqOFj9M0xuCZkPqv
njwW7T5RujtIYGJWNeIYH5+GKmygvHwoW/8rJkvW+W8UWg8thvPabsYxntGT1Daf
AGIimcWPQJGOq1H2FDpATKkii5QmOgtYhcoOMEDWnTz3Gw/EDWhOWr34UfWKLZxO
r1jb27HmQKS49mGuNHNPSXwccLPcX6K04dUC0emTPwxQhJKoDHhSbmyDNFqjx50Q
T/YuH2Ugwr74UwqaODoI8berILHvWJiwoSbQ1k6OzAr/SFds9s9uwOzO5AmbmFAq
js9sq48/PXjyIstUxh8bGuflUotFs0+8Lr3Bkr4UR0CtaxKEi7Y5MuoT3GRiKx/a
tyKCoTHJZQK2BP21FbDiPGyza1J9P2spfvTfM2I6xL2deK1t4Lmx3NLzXHpRsMFm
xhrttd3SqacqLwWBuspVfxGhaqZzTyOjCYgCXukDCqgdFLd6zBKefbzo1uMtGA5V
6uW7qT500giFzG7VZvkWZKnTddn21l65T8OrEDqyL+xrQqG+LxRsH/Qi0f+LRYpd
ZqX7R6NAY3UriuD0KalWCIOI6laX6z5y6ErJaSiQgopOs+FhaKNxSju+UC2r2+hB
QfdZbsGU4JPZ4h6PYd+kNTFO2dSLWzKW1gYZea7dnN+hKW2eSLXdCTvzM0R4d7sK
NA8gJi9vhZrKxBnwPEUvDsVCxXK95Be2eHIwfmp0MVPhQVxUcL0mNt3IQUwHmwj/
OVkhTL+QHwuzmE5iGLFljCPUeQSHIuMClKsLvPrIy5k0HMrbj1OpijQTz6C5O6Fo
gdjcI7jEMGgc+2zFrnSq9wgswKoJGZO5QiNALYtl/lBedB+PXjITgWAeeYzkVxju
mlH1jwqXxrr45xWWyORQaZbtMzN3z5eokhYIq3+gW7ioysL9oebQ5tu6tB5rcqAf
TgoFkRu8nlOhOodzYSEHtl4ozEIxqRdI80hAKJ9vlwA1uYeC0q0BTtN9TevY25gp
w/eSHKevK34J2jPryCwMcMd8D8/3LiZ1BWkVNO3/fwi4+UDjDDBPL4DemXzLQcJ4
BTwyrKn7l7Q1pTk8g4KZNYC/AQQbz1dRCgL61ebT5QvUHwmAKzyFXhWMosBpHLIX
5T1t4RNmTRNwVmB0D9RpGx9dLy7/7x9Jnt9yk/LJvpSn9n0/4eBAkq0hMLvz4T/y
Sl2JAkUku9gsb+mW/5dCrtUS7zCxyYGJe4O+0lNzhKTgkjE9SfGpLSJLuUwAPwgK
dNgtK3sLstLSmzS3Lz26EekwyTu3hkgTRywLulogxJQteaMWwigGtbhRl9LmLn4J
QN+LxkW4EJyus3/maW2B+W54bCx3mJyXtqu2rpkUD0Ntp7wWsA/ZbRDNosrY0KKc
9pE9m/rkGW+FUkH1RS+1dhNVtkE1wqM3slfvszUkj3xvG401PstW0A9CV0lGsnqf
FqI2NCPDGwk5JPUPyxnfoBPx3VriV+o8LvJNKaPRbj9b/pJNcWiOit/PWCg5OYLm
E5HlYY0kSSQ13GkclpKQPufJ+CINjBmIysheksV/ML7dUun5IHkjKtqkzFktrhnR
KQx8gZxrGHjgpGz7a1s49Zip4YhcALJZY+r/PhpzoQagCpGrvuCPCTPsmCc1s1/l
DpICRyuk6l9lyn0IvnDcHNg6X0MFj6/u/ld/b3sW8MshSbNpq4v7gCaqBoRtU5t3
n/GgrjHj5btCphgHIOc7NL58M/JnjR2BqDylAZouMFzZeemoAb0DeB4Q+ER0hgas
s6f9AnhUS8L6xuZXbAZkdULEFtHPKEb7TwjwFfj0T/YmRU6uKArW3OdbQwasPpLU
b90jKYMag57NaNhzfM889JrAnTC0ERgu7V73XORi2JQZBLOkeQscDgFaG6ouALgC
OXC2MFksycvEZT2kFD08UP05uzt/sf8NSlTI8mDFJc5ksWJo07IXZqNsBv1uUKqo
vz0DAc6v2vk+gy8n0TWVECD+BUkzBSfQ3HYSBbL0b/M4qoNqm1OwWLNBHHHQfQkY
LvVToBI/mHgupBdBuu0aOxfttie+T7XyrRxG2jVZsdtvvREBsq85fjf30QKoaDKX
kDPIkOJ+LH+ACn5cGsTBNX34To3rMxGFxCkkjw2xBzXNR4suEnc+vc90chztyFvd
eq3fkG8F4Fj6WV3DhckmqkiBcXCjTA7CQUEPC79aPYr0sibqOv9zELo9O0dUzoO6
Vx4HqXtSrCZqPhYXDW/lRtS4fo/kIVA1r7HeKLNkG11jqJeawrbidqB1UwY3p79J
62zG/KNoNqswGhx4Az5mylJAnU2gUGN+KOzNUUbiEdDPYtAa9HeBp9HAZb24zdtr
J3b3w/FMF5zSLMZ1xaI0vg8os4SVjRJZn8EKDTb2CpHHaL6ADAxWwvU6jBp4fxyr
ObBnThqYaNw9EIlfvJH+qdxLrBxWvU4pocuhNEYwFc/hFeApUz06JAGEBE7i+1Xs
FXjOC49TybWQjs3KWa80+Gm2b8wNi8ggRk7QKZsoTbkfaR0/xklLfclH0C86HvcR
U2Gq3MmNUzv82IDU9RPDL6wZZteCZqhrtM4d3rw8sUnvsCeqWQl5HiWVgUfxE/gC
tVGzs65hGWhBXXH+yqO5d+hHveZeyDGPHDIzb4xUulZJxvL4Ydd12/ShjvA0A2XY
grnCN8iBu7aaV3HQnDHRpS+2bRC8RSJx3gqXxJ4V4CFGD5Fi+ASUVJV5wbs584Sy
B/B+mUkqfp9aT7vSutuF4nERi/2UpP3TADpF9BRhNYNw7Vl5dp7gXt9sw/nP8P37
QpR5gJmOlIY8p+Km+KCk1+6CKqtouPbPjgG/z9C8yCB0UkjuUxuZES3KpBI+820d
tCfojFVPnPDlRuq7XoUxk3gAA0z6H0SDADJWf3SwVUetZG1CI5INFljxaRJwbskk
axxTnzg0g09Cz7A4YyGv2B01WrttQPfCZQYUEbkdycTfHVV/iEvAc0cnKKLaN1aU
9j7/kK1sySuL5yKeqxlq9Ltxrit0VzSLYixmilhpDrfPSgpDXxWVWlQMwviNTPhP
I7aaEelydhsGpXqNp1oPzk9s54yOKo06cecplLTGjJu3zmSBoWu+5LoneupJzZwd
e6vGZsbVZnkNtdf4+PHA+i77B4BJUXszrlwymqVgWCpdmpGccT78rTr/t0A3hRsl
yUrgxXjRrdWO2NvWYa+52n9AeSEW5bpq0VhO7FA4q1ZjcdhffEmt7/BxVT7wxgks
+aSV0P+bpo9RdRkSBC/aoiHaPgvx4V6COFbIO2rio0wcaL2ERrEw+2Z+4VQ9mii9
oCQ7/MnLzECgwGl5pT8ioGGHYv8ZngT/yOT8eWT+jFkZTyirDd5frm/IkW5cdVcX
X/KkwjzxoKFTjnQc4NyuRh95w9CqyybfoVQjC/U6sOH+eSE2P6woCvTcOO3M5tKU
bXgnFPEBDbUBQpJuHOKb9sB6twIf6BdUkS4sF376bTBuQd3ULOyhDohZZLcGS6gR
sOXZQ5I7w5HRhbMeLEqGqr9AKvN66Yo38Q2YR3vWfbFnL1G72Gi590ZK5C0Lk3C6
iG9w32PkpiIfAhXpWQM4sRgjt8lK2J6n0roDO7GUniqsSKjTjGMCj9PcW+TroBs0
6XzYy24iXJ7Zs3cZRtXMEnaifYLg/ftUE8t2lB+tUm5Cc/3/9ZDWAHHQgKTYA2LP
Rwo1jvz2CKMKOR9TQWlH1e+UIyK5FyZyqDT2iVnplBlIaYH5XvkdcdwXfgShIx08
JTYvbfM5up+QbqtndoO1L3x7QoqLGSPNco+9DILj+BbSwUFqJQbiD/tBSUqO5g8M
8bAYqWRI2Dz4y0hihFXioJ+/3w2jtx8RS8/5cbvFebAZDEk2R97GkO2sbnlbG9EU
3XXcbR9svMpz7PTDxsJWYVXZwa2JQ8ootPTIycLDtRc+Fo50/yl6R9XcWKKdvTPl
1P95BpTKXdNptIy4xVyST9qmswjdRPCcxJKUYR7vG79nnaD0fieWERc1UTWQcRpb
Mx8wGeyTzn9THjsO4pK4STOOqzjRHGEZ45tdNxxdDtHamI7wPXFCIPerTb/l6R34
1mawreO+bGia8A1xdJ0BQ49f5GTLdMvvv+n+3NCDXDZfMlaQRMpQWLKOMGU8zL76
4S54TBZzFepRV11eMZEWyVqJHmt6NYNU9inzocm6pt6XPY6CKdHI5ji2zEHzYT6O
AaRyQ3HSyYiO3Y1HQXVn8zMdZx08QDl0KQO7wyIfE8HaYMteE+ID+79+nZU7hS/D
5DUdJ8Un9++KUAReMhGR3oMPMJwo/HbPqPS84KLuJvf9E2fnLXZnOmuKb9UErsp2
nJCupwZbwhzhJLHPL6cmbzu2UjC6KvScnqSY7Sb83tclEZpuO0YQNXX0E/5uQOuH
JV8AkBr8WDEc9oeoQkcpz2FSQJIRl6Bnl0oxcQLd8XN5NCJPD1DtPGsTKlYMRMFn
7Y/ixUyPVT6nUoF2Cx6tiLjrXf5tirjeObkP0S1K/duzERzhgtoCVvURvrZGarsb
8A48ES9XqQfF1tpej1Q3ru/EohYMo0pQpjl7nhEUtj8OPXt43oHmr7AfJn9D7jm6
+sfeKzzUO8iNyBlAKT2IlZs1x9pppJVhnGhyC1U9DM5oyJHlPNtf/DV3zIurwWNr
VO670xFY6iA3wup9R7WZN2zSJTi7T8YNS9nZR2qN+DpfDuTGMjjG6AwSJmGAb5zS
gkErxZO7K+CANN3f3dI1HzWvbntlLZdzN1cXLd5uoTrDbDrvUpDZbASyLk/U2ioD
0ZHxgi2RMXh+QFpVUdAqGJraotVmN5PVlMqpm9Teh6BYsuo/h1M4KzB6V2xm7s/T
HrMc349KpTtCRxkuvvoxoc4ih315MPxuVMiPL5jb2BdsTQX7+yTojsuRrBJ+E7Ds
5Zdb9pbrvUwro1CzAqG3phaQFfiGbrq4x8v6KpNUdcsR4EuhEja7aGfwBwPodF/Z
TX6HCmnIfWunZGM4wmtsi+otqCSg+kZ1ulQf1dAaMNEt0O7ehHyiQ6Ag7DYvJNqo
60x23hqehq05uhgTv9AGsi6MHWksARPfkKwanUa8TxaZBxKW39WIdKVKKGRrDcRb
E6pmXwulyuWYrPItJqvYFnpwj1HqH3LZrGZx52E5JSFR1VOn5YCXgfYs6PvQXA7G
TdKWzk7XcUM9EBcX2+GiCyN0tjIWqqeMsSCKE7X3OMJrGjUDFiO2VrOKH5JTtyJ8
D7SYfVLjOfeQ3yOJxz2o5xazMVe/m+3NdT07/0KE+INAY1yukv4V9+ezF6lkjm2T
HJ3mPinLwYq3pXoDXn9HkYFPxKdQ+lQ340dBqCiuyG4RM+Vpra7/P6F8VJcwpNou
yej34nIF76M3IwLCSQHpZFTzIHAA1DndZHT/6YFGNLOOP0deFt3gOpXuJzh+KdXK
nuYqYOyntq5J2eYl9EicvrfInAjUGudauvDIYhqXIKXJeGSGZZKxBrFRZQFA93RJ
zSmmdvZelcY2Qj7qFt16imW8wd+Dcqb5959TmAsSrQg0X1fHzSJk+p5hHscNKPY+
1nN9VuCo/jqBDsgVLfZea/5azPok0+uQxqJVQYg8R7g25AG5gosPhw2TOo01mT7o
MRcB4yvvWi7qS4TW83CBA8uPxdHN98wAtQ9ODQgIwSjqkiR+YlqlxcQ21P9rLL1w
CFNb1rsh2hITbhjBeMVnRInIvNLk9A1NQCnft5tAQJQEdxHhAOcsiQZYeJ8l6dSU
UhrVFaeohjNKvM2/Po8jtPQOUBbTL9YU3xTe51YdIUTudg2K10R+bntEA/CWwyoT
WkgTU9VMo+1Vt/YebGX+VW23xBe6WXo4z+//SKQFSTNLYTTWvP5+9XC/EwvS6Cu5
xmakdu71/oQWEUKw0IeOsUYUJbH7A4mQAwsuEdhHjZJbaHx5S8kVs2WlGUjh91h5
5eqthipr8v3zRors+c01Tar5Ts2mNxFaPFtUSbQ3oFgAX6E0MlvZZOVv986RQEzg
9BgYbWMoI30d/LXek/VJRy3u/pBoCwY2wCXDyBnj2x3aVyoyQfTDsDISul6JlpBP
PWzp6Ur8QBCrrnSoyAcmvQ0ezY5oj4fSPHSEmqKUR0BNggcipYU/LRqVS93krnFx
1yR9KgVnuzm0I9pZDG9cqjyKCvZJRUJtR1m2bpbGEpkM5xuTw2it+k8tNflxRAfT
vxFGLDXMb5GZZTfpyjcQwJqABTzZ7JwvBJ9JWbvseNHl8i7KVQpf4hhiIDD1/7RL
hHUrhmfUqjiIwx+bFnsX2dwX/mHgiPeKGOLJdD2jy4MdrP6gpfX4LILO5Kez47mm
oRjlcc6xRB8li9YtlZq64GuvdDmwH0lwpSiXysH2RcrPw5XRGleSvvibFIN7BYyg
3orMKm26lLV1hCT61X3tNWFdjvy2WLPeAqcEO+sRN+Psvd7oaOQAfbkNKMA3JZIe
CwrN0mV5gznXydEcqTFMIl/z1UU6C/njwzSXC/PyxDh9VXvi7suUcA7MYTtbvRuP
2z2pj5DSq7L30mSiMvZ0SbIE0uBoqpoi6u78d89XY4lvDh947PPZs+6/y0tH5LaA
xZ15Sy/RFxX9Cc1+QcUZ3Mw3xEI1/Pyg7iJM7iWzGdaPHcreDZQl/kJxoRNs5T9k
DthXDtMCX7XlNL9AAf98JUmGTrV/EezrjBZZJeQSC9LfGH9mz2TpG7jCrLBAGqtG
WXmLEd4EaMnMqcTa+pSnDePo66At24emqCqH0ZvaGxpAn9zLyZfVBfy84OkTwRDk
sNuF09hvpLxkU7sL/KKVlVJPMWKauPblFsb/bg02PVEayA3lltnM4W3cit01WPi8
J0CFCTsN7xrjMC4ANk5VhBM7OBGkJeu9TydvWIOnGluSuXLDx3L7/S4UxviwNwB2
LqTuM4GlY1uw16/uKlPQbNm68xFRNVxWRZQ1XVIPdWl9I4KdEnM3mV2xNjL2RpyZ
y9FaOcWuNnD9sYBhsxWLBZ1D92ZI+kMOQ7bUMzT4h4Ox8qKy5da4rs7t6pVMwQtg
TpniGNUX+EsXBfEhXSj6jva2zw0Da3/KNioC5eHNczXTJ67mw4YCAxJQI4cBUCsv
FGalO5uBwHL5Ti2wYpEupizr/FJs4fZ2jrLbInzPcRo7I8VEGkUsuen8m9GYe0/n
4F1Rx/aML9WLXzF9L7x/jzX9xzjASbNs8IQZ1nJUdayT6NMkQ7KkJWm3ki3FyVhq
oIzrdVnF0CJK4v1IDitWNCZdsXa0liD2UFwof0TxFq9Vsuag6EkSy7s8ThCIl/XS
Elgf+02DRXqc7PAOEDiURWOQmtAj6qEYDe2+aRdMPXs8TBDlUw2fInnUTBIfufl9
kUauREKm0ZiTcAmjVF47dodUSazKzRJUxcUXPoudrmHPtvGla7+si0KSuC8oglLD
NC8MO5p37BSullF4XDLxsQTIPYYknvTPlILofbX8/n1PmAicH+MQONEyDzcipTQe
kkvhz5wbSa9XaRTSccUU760jyETYakCCBa+MKj8Ur058pwHg7Z5rjfFFSuCbFnej
JeHO/fzdMquUE7hTQ93FKOHHtsPv/GDmLhMIIT32qWDFjSYmJssSSkvAsyBNJSG0
ntb/mdmgUwlspQ4WTVu16J+dWeGiwCuf55gYyAQaB2qEBosHFNDUdc3gXKhRsBCc
Y5t8HZDHW6qKL69QRKu8j4Yir4MVhwTGWxxopKlYeIsDir7sf9IMGq+tkiPybiIh
jUV4k3exXiUWunED2TeOHphrmiDMtkdJfnK7p65XP16233nZVbfI3WN/RjbfyiT/
lUn4soLdaMvVLGJc+BKx7XfyxOM/uQUjp6mbEKxJnpG8lXhvdLSGzpEG6g7NaZFs
gylwtLnzXftglcpJ8nA/SVybrIfbNgUK/duVCVFRtFYpJww6/RFa3DhJ/CtEe4i5
NH2kwWJ1RmMj+06LuzXMis9vFyd/NYYj4VhpnkdwQIzb5UrFhuEg+euhLjsX95N9
Il/6xIiUD4cMjgeeGQ2pJniECLZgDsvM2bP6Pf69x15vD/WhQSwSB0JkHNHYQYlF
eBN7xogLevMotZ0k3U7s/gvkyMZ5hSUCBtegwNyvtOTUgNUke745rbY6AucnkfKa
tuXg+nQ05MaV1Y4JJJuqiXUa2zyioHEcNurxbQqOhsCOLziUHfCweSBpD88RdB/V
iv5ASYupWW6k7dpQp87L0oXOQT/C8BfK2r9xogxH26c/P4HabChrV05yvajOf7Dn
ecYUdirJO5TX8xC//hewK66IY2YliELkSeMtYWI7ywwQ9kBlw81CcFLgwjhgzKCY
4RqLfzJ7TsiL3qfG75aoM5tYc/CR9NCJD++LxJZwP2e8UmHe/pnDge79bWXyhETo
b4nYiPMVNGuVwaX3YvbeoniPmeZfPY1Cmp7Rt8vxqshG+gCQMAa7mrMvb/4la2px
/kNzfw+t2TtSK7eR1ihK2G0oMaqCZz7dEWx4F3qMz+1tqpiM9uQcUT4CaArLH5Ea
/rw+1+TE21zuSo3fqz6ZO6uhz3WbKHnOFRmn1NHAM/IZex/XRk7ei/fManoCUhzT
BckTZ9+fRCMT4mAnLhDSwHbLNjAfliRM/a3/enH9oMa7H8w3DKZACnYCEVZvlQHT
LkwD1ebo6NCQhpmbADzSgPxG89mxH7CBvCKy1Ei+V/KCtGHSH5mxvgXuNqLm57ME
JjezZyLDGCM9cDoDAVkJaDIPHD7gjtf4jzBwZ1bfajySYQMBfj8Zzx7vUNehk10T
aVaQpYKqVnFbt3chcBKOdbIObyaChI6ksCGLtEkvj48k1yFLGStMJ9qS1uG1hVV1
RHIpdS4ni5KjmRCGCrHWigfS4zhhDq4bOP7AugwX9wOh8oEDvRSj63nZCdpo1jJ5
M9GLhqL23O3WENVjhaApeQEPxbUEPbd6dfN/qDbD0Y1VpkQLbDVCu6FlI8l0aBfu
JI3ao4bbX2xERhGJN9jYy6tQH9NsYEVWhAUEeUNlq4QfkRpG3anDX229umdlBDjq
l4d9bcw0UIy+ygrA+nOFfx3PYgdK4rJnkxh9iilGoEJqDMv9+rFS9DXsFsNBbkdU
+YqxMyczikMyEFHmE1y22W/F6QXMa/8zel9z8Jo3ELsgh9I3wZ1T+wnlvIAs4lFM
0sKUHgAPE52I5G3PAA2mxovlmjCIUVz3OPW+KbfH7Sy5ZjFol4l9ZfyQpV6Bs9NI
3cjGuYmuRPgWyP+Ct2LWaNnWOIjbvZNNBPDP83tKewr31WK6eO7gvYJpYDaDXXJm
aHfxBQPKCTyff+r0/c7ufjO36lUL5AiYurfFmYHAhPyitB78HsJP3ABby2o3jhbB
uz2Pq2tiQuBtzZiIgHeOw5GyqV14HvUD1vpUbSzP1jMvy96Lr64g2DKBJ0PqxOZ3
Jse0BIaDOnCvjw+LnuQc7g5nBUCcaheMklAxR/1WlLukeUu9s+n32ZVjVcqt6C1x
Mg5btzLr3mATmgH6dQWtTCFWVF9n7Ky7QKXyjENp36YCfWHV9ayoXAqCYuP3Tbyf
dRZ2oYwKaljc4jGs9RY4ts+BpVqQAgQdqm7OoKGj2P3VK9GdoV38ppfGtTtwGjui
w5UFRz6NTvNwmAspZGVRgh+T7DgXjTZxP2Y9/0CXRvdui4Q3JZOU8rMs0YsaYb+2
gLZ3L3fo9895eQz+gCOx+OolT5JcNlapicvJD9K3neADiqpjl8EkPYGoOSMKSdMp
MDC+dF07/G+4nNF+ff0wkInfKn32/uBw8eIAUmWuk8QRlMemKdvLvXuLjVNS4rU2
0bMqOQmvqvIeDQX43MewHKPixc/z2MS0hxnxGthHSSYsu+ETrSaqm3wdl6zaOtFz
lmU/4wjRqvxLOtQouHpiN1eWtGabn/R687C89WTeKX3w4ThuAPxwu+GgkD2rOpHy
R9bRj1IUoCm6k0SM+P5IbkeDycl1bCWqt7eEU5AYRG6ld+W38AUfaGLiLQFqQu2H
QXXlQlkkr+Y9dx02XS2AAajUTrcnZk6XsbpkCJEIVegchwGIqpqg7aFJpWgkLe7N
nGbqUvNoNFXI87PqFjJCPNg0T25D0mf+8so96JfI8tTDV4x9XrKXl809yKbFbSZb
bDE/lHOm9heAwCZA1o2Ps4LU05V9ilK6QAXjWycSFXZ0g2QJlMjVqGlaSc2VBcnt
e/hSmHcUm4ELGZjPv36schCtNoKhjR1YbXbBmEmwDsSfxFBoJZVoJY6XvhNutEch
fxxRUc963+Fk2zjsVLz6MHp+hORJ/4RA+WyJaUQfEL8u/8sRscVYlY/ztKXlvLcF
i1P0d+68Fg+IBcEMmUU6AzCiNm7XcXQXD+TMd2I6AHeJW2H3Qzt1KH7kX1i6m/z0
aptLICEwufcskTXtGkXYKSyk+Yw1RcJe/UO5IlcByNDF4H1oY6pAQb1+plTI/G1F
h2W9IMAqGbxiODfLmvMHRMzyHSwXK3D2kKCzkqNmfpI/YRpf1rXpjNrh2bY1tX14
A7zXCSCL7G0WFBkKCsInxvNDvwoS+AAdb4R2r3jvwgt+WQcTb50JHMW1fJUr0DMn
eibkdu4a2PPihIMEdJwyMRaVYHXbQ00j60VewMgwUsL0THGL1nk73sjc2V6KPQZx
lZyIKo7tlTsCX/AIpD2kpiCgrdCHZcK7F93uMC6D7P3twWzybmgFwIEf69tLldmf
nQsCYw1G+9zyms5cj/t/u0ujLkZa8+tjwLl5ze9rt0+MgQtuJ2KtbYBIirrCoIMv
50RlmaOZpZc8wvahzVtWVemBp8CfY7pgmlCqr9kHLJ8+Y7sZ+1qFII0BF9Dr1ydI
gxxARlcJd1VQKT/kmtEyv3rktiK9uijePPEWy5d5HzFHavtPYHxgc5bIZtZVBmpg
brJ4mlWlJepPWqd0a7NYtkrs1tTLFnnYG9cSvb9lqnfw+kzDEeGpCdgbBYkgpFmv
QfWXZaboNNTjz0TH8y2Anion96c2ALVw2v3BhJtUxxP9bBoNzxo7Ft2hDnIQkIne
fU6TZFXEqUeM8qCi1FiwwSQyGlzmeYVjuXGjv/mgb3TzPZ5b3JLu1BdNbwd5YOz7
2niG9KzrUL92MILgQqfAuDYA0oh2MnRDG4JwX4U0RcWwP4/ue0ptCw0CYBiLNTtT
LbgpZ7nCs18rfQUY6OQ6hKmfWsNaN3LSrPtpNv6gQnQ5ibZMaaI7n9WtaixaS4v/
S6CrpiM4HLKjXd7AGFaewjahRUYOIi4tDnpyi9LfhCq/huu1v/RUQr7Wh+WSGkab
2EU1NUo3PpaK2prQo0e90dyUx9FtQNnvHzqNFHNEOWdTOBnBRj0xsVL3Gffny3A6
kh2ASDzNaJbLhdsKDNgr+7mpjXonOo4E++MGgaD2dHVbppjtlcgCdub4nVFBVsLR
N3aqWaxSxdG7e5/mUH1MS/pGLjivMQNTExgxED3/dKclALtphosgdzhdc3wW30lu
MTH6a3I0MTTJbmREm2RwDCHmc52wlG09t+3rKTFHfDs5l7RG8Lny5Um0lfWSOh/Z
zYZY9XZvKiYKZj8I1OsamKX5UYg1Oo8Jnc57eQ6B+krC4qNAOEGCpxyd/1VovuVU
/9bSiTnAB6MukTKlvazKoFCcOFKkij6ygvuGn1PquAlYI0y0VukObCcl1kE34dM5
PlIkGXjcl5FZfm/fA+fQ20dVc947R3Gte2Bj9AN4MnK/OFp6HsLCTHFFVfUXeMyv
3x8j+IRCaacUL1ixPaNXDvnovGXRPEgM4XeKaVOBt24dJjUasJYP73f49CNFowbp
0av+6tRz+GbrXc1m7hrCkeGWgnOrXvIn7Hr97CsBbkNilPcmallE/0aHLSUUTg+P
TWy9IKrWnzRC/3wzGfBM5UdivV8D446wPdiTLzATfeptyTxVnOJ+laSOZUBMbLiv
i4fDYwMwraYitHP2NECKDJSyb/TdLRahDOm2Kcq/O9w19U9c1tS0GbHZzfqUSnx2
p6cRD0gUB49ssP34jDj2sAWTc3vq3KnpRE2hM3M/M4hiAduvgbuh0Xd4coFiJQFH
KD97jQfbT7Vp5SYxg66coqK2iNgpn+BIA1QmjzsTy0QKXo3CpnCmuO1S15+ZzCZs
q3MfUraS/RdDd5SBLh4d5LLKc35BQsNTUJHcO3qzW83IlOH8CATZIWOQLoqSiOyD
FCkhWXRALiDFwfFrHeeY9uquOnJN/n/hMMIshfyU8LqV6C1O6CkxiGuw2wgQsDAE
rKbwSGZvn/eqODu5s7HTpwdanAQxsnEM8zmzTkfETfOfrZUPURXwpmgnaa3LPYsH
SfaAWZfjhxFxxX+zGlVr5HulB92TSdqVXximWMfGYx6PPIjymXD7BWyIsBA8XXEN
RxQk+imYBjyoPTuV06rmVFZMQ27SMov0Sd+iUa9VSKAMfVOo8L2aeVJ/BNk7D14H
MFHuN200bNgKE+Aw+1ONBLQ8l7gkpSEroo/CU6T7eOgazkiPMzMUJh+7MfzuKqqD
9G8PbCClm9ohCew9fwbI3orZb8Slhwp4KhmR8VLr3b2r1uAt4SRNNPcgGyQ0IS+D
TI2t8YhEDncHUGpZnhviysfiF0B8/nAwhbvemVHHIqt582zgjiBMXT6H19KSfTa7
6iNSYnVxIkVq2C7RCJUeNrNo+6Q4nMZL8ML9ZTomQuaeAxlBL0JWZ91FkOjdjlgD
KFREx9ej63JK4EgUeoENXPpVz7ptbBCK9sBR0N5WbVJyGCdVy5y62gsk7/IiNZ4i
4gRN4T7RpzD+Qnvy87xanak9IqEJ5rPGA1Q+Kr84gfnG9mcP+QYAToeBOOM70kdU
7jnAP2xoZQ979emtaPXTCCJPbLtRrsJ2aeqFvlOHI6l1UuGza6dnD284rD6F0WDX
ptS/k0JYcG9YbofMVbNCaqLX+oCtpF80u5I/iZlsftuom8OIwoFBv0SntARKwX4N
WlwcTtEIvYW5gtZFC8SbXJC5eOBqpGoFAZZbjEpMYB6aV8EtUhBiS4iBcUCHTnrQ
c3TVXyh6W2N09y5dfi6fYmdp18bON1tZJHalFcD1tUsTqZpLF60ZJAjJuJXokArO
5QzCJEq0DrUrt4cUuOH8WEolSugrM+B/AqptzfNjNa2qEE9T6qTsVmbi9ESDs8BF
C+mkAXnuvdM3JH5ryv+w++6txBMzB/3ikcT82LWPUdAVSAJMTRASnPxWMYwQJWTQ
r376WexcDyaqBNlFvPLLjrxt2j6/5ALHVg/XNYlwPy38wfhPXRJvOXJHYAfnheFy
ehrw5AII6iJNcqaZI0ZVz3Nyo2+rQm6UNCOtM/c/GfcYEZ9NI2MYtHwzlM3PPkoj
yMgZjk7mWm0XLOAChro1aOtJvtt3AQcyZ8w1UMtC2esu1cBv7JwTxM0FZ2KfUB6X
U72qmsAGfGrNc3q6l6cLprSxFtnmnGOS/Xjyqd+RjLgbaBl6fDRHv2YWIIQIojuq
ldfrya0FW/+PvMbIxiScAd5IsOHETuzgZKvuGIG5kTvCXvCULqe35xOdHjaCtSTL
fP8MLtD+HK03HvaGGxk6JDyCvmd37iXrnMNrLpu8vQjmxDbIsx3z8UMbZjKitU4Y
aQ4dKZDoOBXPzeN1HvYmF8AVNeKF61Ocg8ukRJeWFF55cPMb+qbtG0Vz9WBsYTSE
lmvHLFx1Rv084UbqTfIGdWLCN+d0/HJyX975AAYyw13I52lF3xAfv1orT3G2Vp4C
5EUeat6yFRyAM35tS2lY52ZDynokK0/OgQYffqT9pTCTOSdQ/ovf55UeFK2lHz3S
s/YNUalhLlDlQYqCUzvyhUNhBFD4Adfn2405L2HsgXSo67d2S472IVGORxv425mR
W8A7mNqBgZXQl6YGc/v/KQ1xNbB5gBtQBFps/uN3gE7lI9gHkwm3VzQHqguOqSZX
7zeoqjFli/lqyNZRqq4DFMJ/XCr19CrWWPA3FghZhEeOHkEVZ/tT0LdhX57UfzHC
dtxrIpIw9jDLCLyIlYAnaeeIaUEykBVHMUvUqPLt8TajLv6GWR75EYt+btAsxTHg
J5oEewM0QOQ1KYXhBBeaE+2YS7Xd+Hh1nIfBQW/xujb1nb9qDGKuyLecK8gzbcsi
RAytKcONaTS1dSxuUMLT2tzEni47+zZGdtMskmxZLvuoIRPNdgSxnC543CBd0GWk
rsYoP3mlQdfXnlpHeP6lRHROtBwRMne88HHrqnfkzcIrz8wtHJph34IN1/v5f1vO
88QrIloeFVm+Ag/DG98HVcBk7lhK8w7VifImKFv8k+tuHxQvk6qi17P2ET+vSYTz
BvKygFdQJwR1ggb75kNnOXcKFJfwnMZmb7jqK8bb5mKCXsJHL7olFm50aSKi2cyj
hai240WXFss126853RGlhSBOrZo5I62trcXldZN/f/pU78lDOifX1OQ9FoIQj4ZL
1j0QhHlGr4IMgaWRuKR3cteosMaaq7Lm6nFDw1XJpKey5CIPDTTLThhrQ7LVaW19
cqZJqtu7XzTtmoH0jE+XnCc6CnWUmw2ihH6umm+p2MrBn2JbXvG0U58dwMKmGFlS
ZZEvqPTOuxDpAdq725zmH0m235VbUbI3ruKuumFvQzcaX8kyD2NUHluMWsA8DYb9
mJSa8zR7mStRfsQzTg0ZLrx3X7mTaQ0wHlgFWmGJBbqkWLu3Lp3BjM58bScEGDz7
aZruyN87UP9SmRHpJywgYBp1WKGjF9ra63UQEIyYNCcLHuVHJFvNx/PlK8ghIxNq
vywcLW3YL9GnPplUDpQS+n9oudShFEas7Qa3RLUwxU8gGK+1nj3C9QEIRxiOpDRB
hKHrGNPzbwqTU3+QcRz47rT3EUZdynKmJ+XWXSyhzSW5TSxeIwJiL0+7mlTUdsCK
uats5TQKzmh+qpQh1zCDv056OFu4SP0f5+p9TjICgmgCXqALUfh5gzvlHLTtf/LL
wEbmNBaULJR3Zhg4RWtVJpcB6Tl2q4jWj3A22p0z2zpwv6g6os7zDh/AW094rjU2
nzHfxs2lrt8XCwPMpk+Z4BOR7ev8tcdvo/6k5LTgB4A+hq4AjgR36XgyH+ZRg1aZ
7rwOh7Wt9HcgQYIaQlH5moCjYmPlZGpAg4j3BuCvES6OtjnXYlUKWZCoiD7lP9Ck
l1ZtQ0VE4Urm639nBINWrnD/Ca6fQ2PF1FXGJ8uptmkuqmEdAoEUCC6z3cFOgeVx
eS1Gd8keww/xJK9xlAiKqIxH0LYH+4Pgy1nj15fffiB0Wf4Q7WWESEjiQVcw0yrI
6TNqyecokp2OXW9UIxSb/7UVoTKUw3nWFGNOwAmRrRlBpm6aIOrLLRQJv28gSckj
Mg7RXWGEzDjA7Ep3+TMWHHrCjUHTzbY45eEGnvdQxkRar6IUp9kos2g22G0Rp4w2
e0CxlF19KlLmckNyD5s2XlxCYiDFsxBrHpsL3sl49zfe82Lgu7ACXJk70bU+z5Um
fuBgLPaxyQxnoeL+Sjx3pL+XsbE6+GweidSJstbFMfF6EEjgiGcK0n7+dLrXavPp
2OpXa6Npc9kgIb9HKB/c4nkqbSn1zcssJes6sWTRy1FIRAbAiijCkz8+lZAZnYro
wkalL14jlar6fne/IWSsmlVvhgv+dYT2iR6J66AkHzXHwU4bPvMkWL8fcWhsxq4z
dEyoXnm2KT8GClVYYdwUg1HrKSKpsZMIFEl6NuJV/5rP2XgiEiF5FotWVKjFFxdm
jM0jqAYKTLBmWTpHt+UXNvCs8wBdFQCFdaucBGmJZ6O0webNTvaHkEL+MIePQO+5
6RIsFsyoQ4rPil+R4hAZZCkaWI4SjKFAoNS0A87KEHoUVWuA7Pc7Zw2yoH+cxZDZ
qd9HouyUF5p6qDsl36kyADZCz5zXaTeUQI9XG/XcuRuRd8OnfHWbCtdlq5t+P+I2
zn4jFvqV+i1AoeqPXnIJKg3fhp9DfZ6D7a3A1Px3pmLeiBGo5DS41bQRwGVtGIr9
qoaH+CiswO41vTb1/hGMQhFXL1XHpqb/W8XQ105eOnaFuN+qWCQkHqkVkhgk5Qz3
qAVg4+xLIqj0aemGrAfSQCcElnO1DReHIq/dzo4Rs9enF3ZOAqRueYLuVyk8eiyE
6nU6Nb3ekYyrw2uOQOnzSkoL7wvJHZ4dpXkss6yum+p+w/b5GhJICY2A5xdDZx0J
w8z+2SP+12VXgHG2KJ4/3+NRb2CrtG6+1/hDRm0+U935oTOnkJF2H8mS8kxTAFAG
7eust3J01FUwDFKieDvP1M901+FOvGHVD+vDNzMNRPsOFCc4Q81c7PeixoSuNyD1
onmrZt6YivLbDQ764JirzAYkwbr18iJ4HjIM3Knn8XWF5nc+N0+nknfNazbBW3HF
mynDsyJUN9AbPp21A6D/Buk1XUHE4aGzDEELJ99m5FLry41F0wYhp/AA8Ikmv9XI
4UssLCeLJ/lh+2rGPNVU+Jkwd++WSsslQ9FowR0MmrV8JV+wQkv5g0aRuDNy9K1/
eFHJNrqeLdJHptoyeVQp3G/JGZmfYPv7ZThH0zNr4G2fxzRUuR7SefAO/24V0Vf2
TKieUK2nvGmHU9BExAfPZmFtKTRCUoWLAgL229pWhepNCgj/yafBE0F0TRoPzd5o
yRc6YTmxZ7Tg2y/OYVWRNhXzoFV/G6VvQ8KZS+Qthdpc2iUxsICtFdTzVkSN2cLe
HKLOaJT0XqYqe4cF9q8GNihUojC5FsxKU8rwMEuKcooMFm9udhJtehYcn45Iuqat
zwrKRAP1EN+AT6A3d9LHk28JbbtmcxFpS/yPWLtWVno9bVxpM2QdBMX4VLEzaJTB
f5HlWg2ixJhZhBij1jjw/GDvlIwn3g5pist95UkWGjMGoHs78WV8m7tvvPNLvX3V
eRHB1gS/qczuRJQasHcFdQq6G7ENpZLK6S1TZKpZQJcMSt6RhddnjHEjMDoZvexJ
5BwyHRYnsEdPBP8HgJiIhGTJNYWR5kHObIZbMkREOtTvNl1HnPbagNjs+k16AKMK
hMD2AES7uAEmkiP+4fDSZ81hqgz37yyWnHYTsXNzWyIKsXg7VzEjVPUYZuIQLAuX
GLHiaJJL/CStKAbVuM9CA7nyf+Brx9pXktRQD+RSjlvCoSNS8+sAYJuHgyQnzz/L
9mzsOeecf8NrNs4uCMTn2WlHTtfvrI7tua5G4mg6LRKvtVgpOl9vQnD9QUpHxBcK
B9/qIMr9F+fZ6WvvKRm6UqMzppHNSgoTrj20oKLsPK6ie+N4Bbbr4mJ9/xNj3Jj/
JHPBsYYiRqwzmI4iFim3AAZ4EHQ1ALkVyEopwcJEo5IP5XhODvyzBGuGkvdRYGUI
gkNJWKqYJ/VHY62pyhIcmC1NycrKbbTCQ5zKXFI2qoR/5SkQZwlgJLo3UbFdR0St
y7lzAreF5ewQL6+yl8h/PYWh0lHThlUa7/DHHzrpB8mkDDLWX3AQ9RGD6Y/v/YVU
VArI79CUh2oxWI6x2OAm1N9auQiP80C+YJA7hYQenxwoGBO0fuo68Utnay2WrDim
5MHchPEDL7cRpq/82yMH+RSNkf04XtaM2MjgEi1YqfMTDRcWpiFjoe6YvqwKp6UP
0BKBnLcbN/KG+KaIly6NAFrsKjPIa/G0JAek9ALDgvBoQPCXdd9IYxKxjiqnomjW
5WDKpwrbgQu+v8k1GEILnnkY5cnHdY/Pi4odOkn7HWQrnuYI8sP25lKzzzLCZtMV
GJ8elHNZFCz4+pi0wQ/rgFUcB/VHc+PNFtTlM02d7TpGQLM9IFx3iq2uEDVGj2Ni
xXOh9c+SX/b+CZt0SR+rNV2JuD9hS1I95ja0HXeLsY0OZxOZ9VHdNao7vNNAEo89
b6BLSr3Aurv00XZzuxka1GNVDqb3/PRWE2eFU14WDpuKhSzT4AirM91i3a2WW8Rv
z5iipe0Qn6FBpEypr+DAljY1u4TPdtcPp6rPG3l3Orbwl62GvQHwI87wDu6tkN1v
saieGd5QPrBU6pV72NfrjZNG7Ss96j9vnr8yTSEcn9dj353+o8REzcpV0/b8R0bI
GyGQB87efxu8QEkquLUN+PT13wZmgDLYt6idLWD5V2sLVXouEq0WogBBhWMSksvN
KgOaUa8NFoCCoi96EUIRNSAcFYjyUTQ7e/y2Ma2XAB+kO/uoAlaXiBqrSR671uNs
VgEPuyowV/Ulcc0sITsysa14ToGT3NyfNyZXMICapLlRKGbDT3nU9COdGaC0S7i4
4Mk6eXtgS23Bjc6Jx/rcKL9/HADiDOevIdd/RcVt+vG6Ao2bDiirQGFexhSE/vCO
lpuRDDFe91F3NAC6t3Foo1QRLUOf+Zfjqw+98GyTqhmjVeyH67QXNR6NAvEFsfcY
ms1LYhuJkjgFpTLGnfApahkMtxbWpkYqUxrteSK/vv5EJ0Q7TCkFDXU09WNsxpMt
7D+7J3MK412H6/sm7MMk/DFs5udXnJlFIJqT3gwMMT1HkxNVWzfMMZLKGYb9gEwu
pvqFtzXB1UNWf4e/zZmOiRL6SNgrxDBPw5QWqDrExH0y8X4fsAPkxOXXGz632iRl
n1xIH1ed90Agxq0Ap7rid2wAvIeeSrVGC0s9frtPrVC9E6ju2p/nhHjXH3BqqqmA
gq0wUcyPyjT+UUJQRC7cAFzo9sDvGpgCCYveoyVUVczhmVavNmqpW+QEhHf1tj/+
qEJ0ldKwREk63FNnUjxlr9cyQWzRPBWc1KX1LmcIa3ParglFgWe3MnC8HjLkJUx/
Fk4iDgXcoWZPQb1t9LwLDXBGZh8f33/9oUEWFJyCW+2CZyIJxhCPvq/+5BE0DuXu
OusYedtU2Li/t7oLTficKhmKGLmdG9ixAonPPKcLYJimSvX7B3qs3U61Us/e5vha
y/tYtEplJLj6VzbtVrSQqok8CdCsmv+0+Ckra8Vaby3LcmAf5nJWjairD246cJP9
arO0ZG5CYnXZ9/b+G7zdfHQqidVC9Yaona/qr544G0lDnFeV/A0wISWf0BtYWP7L
+Xk7eVkutKEF7GDj11lHa22O00Hz9ObsD/5HabSl15ds1P3ufZ/F6Qo8mG4SJ0kX
lHBZ6vZRGf1eEOtVj2JByzdr5+wuZc+XquOnpL3S97tKYaAd8ecz7xthWl+p7Oge
hhGZvuIKk8LGaWDCS20O12DpuNpymMQ5yfPUPO8S20Twbcge/UVetqKndGsxGVhk
ChlzuN1c0yW5al6nV6EBi+vXJ+8EZ6BnfPjfArSrFyPOoOedEQZwPFNZhpOqAMIO
UR5kB8TwwunF1k+OrPDbEYMbhVZ1NXBk8/bnKyek8TcmVg2jKz3atW+YoqmDejkb
a0mgZjurRpuUUsTVpC7C4Nfk5IBsY0LPfafieiuDbG8ji6Q1JOujZ2pVQ8PktCcV
3ro9IjcYNJiVyrDxVww0QYvgfKd1WHidMqUHRtK16C0Vy5yNbIRhn/7eVRAfo0XQ
meG14/Y/ouOA5f1gpMtaWQNjrcvOUpeF+3Ppr4L7YY1iGstldZkr0LjgNO090vF3
TkMHonffbwGsBuAmGVZTQ0/EUlMiSdIYcuUrKNDEDdhgobFvrnZR0KTzvrjFwnis
NZEpVcu2X5npL0qBKkO8oGqnooHyEzq2dHAc6/4ApnXsfMSh1yDYae5yyNhUVmCz
uPSPAg3R++t4bMB68r/nsW4jF77xC/53KiWx+i4WYrdiIAa9pqvYBQ5DE+sPUyv6
zcoH37p/6JmD5NpeHJD1ILuqdNK+FAovhIg5NFl8jcLhOMF0f8P7LNwLvDCVTJV7
8A/PNC9+PLQIl74Exo4vdt1Yb9l28tZtqLQQkcd8UpdplFurSvrpSL4t/8f1l3H3
71JY2D6iTs7FjN3ExAAjP8fMNAZ6Zw7BELx0xwxRUEBtMrCOfQXKVNGORrux5Cvs
tjAbsL9v4a5Jo6Gg+HcmC+IyKslOg3DCNxFr1gqYmkPJW0ge7Iy4b21mVqqBIElp
rw2iEBvh7/hUpst+oEzSS009ZLqI6OzxWDrX0I5xO3Cdg8TvAzSLAGcBx+QmVHxT
OJSwQzIv8UON7zLtrFdcQIH1PaGK3G3fZEAkDJh/1IeG1QO+x7G/pIoRVlagD9d6
61DAZjfSz4MAzU7p2+XjN77mKkuIBRIfeyg6e9RgdDXKAAnDD06W9cOWIQGuYQ4O
y70/ms5cx029IXMScFvRUoGmJ9wDg3m3mKrXbQiRa6DLklW6CXgbBoO9DlGFDIrd
DKNZCybRBwuZPRxJQSxITNaO0jm0Xm6RlbvLcMrcHsLczXvi9Kdu2aMNSfbXDP/r
Ln0U9yTGkVpzJzUfPNu989GWM2NLvKYPWjYc4w0VBtSWUNFC6PmHiBMGyVrSoHna
jrygcs4Ytjlk5XM1KEK01BA3Guxe3DZD/SaYA7uWAWoMgrVXcRTG/Bo8uFJdX2ob
QEai60U9rrcOzypgs76wJ9b325F5LlWcpOjD9ELVwsXfzNO/WRckmwrYONRxsdIb
ztEHqezT5htwsV9QIgvetI2TTz/xHpLIfs0T/qTjJdA7iy17teZ0R55czk2+sdV+
dyiaDcLljFAX2YZ6MWQiUGDTGHYRCnuqcwX6xxtk1xNAu+BywQ+Ob95em3lJQyVb
Igf+RdQvuM0hNDh/mftWkowwN+ZEU8dHazRNCZpHrYnc+sk2ZIQYmJxzalRMTSAZ
32XptI+UnEo+m6wrxhKdSaLugbOEpHbD6VHM9IloziUbkvQUWz9DnYWi5/ABte/o
QQ9fnxF8V3u2IYe6vYgkpIXJxMfjffg+7Lx8LTkYyhy51hG8xDUIsyVgk59kRrdk
lJ1f3qPTrr9h71fM5q3Ms3g1+RoM1W+o3NwQID48gK/jxOoiwNRkQ8fwjVQGCP/e
o4xkZh/rLAZos1Tk1SAXfKVW+4Ic6P1nv3OIuPDAR1URpMajSOS6Te6qgEpLJnWL
sy3xWbgqZwrDe49OddXXiwYAGQMdnV7yQyBW2mC6KJy0ZJFVDkwpv1ST2xAhw4Qq
jrUVR747EEAdyFgnTuk4hlS/VVIguNh5TOnfuZBkrtVUwtxMNxtCF0cqpeSqUQR6
8ROA8s1BrM+YRI8lObK+pH3PaZyAuFJEq4lo5hL9Z1waCHtCbvtLigvFZrAPsRpn
PteBMXi2K94EgmD1ydRJU7zQVPpOEpIyMhT31CCxeMiflTKI8C9eJmbr2n9RnNyx
3wrcAHvfsL2DLqFLC+zxdq9d58oGVJRgkHbol2hsQ26Nn8RGDFKK2QWyPCzrxHKk
rgB4VY42uXj2J7NoaLYV6Vc6+LM9GzO0rvGM1law5s9WTFW9Endzmlu94L2kJV2c
XMuPC1bAykHhHmWAYPK0bPimGAEhBKkgAUdgPbEgtF8i5DJTrZSV3ERm8MHpS8uM
+5hYhE0dv41LgT33n/0SWszsy8olEnK0YSb+8WvRJYmUjt6oE37F+D/BquGLYv9d
qxOc8Gz7YCx9OAo1gYJ6N7Aykt6XtiDBi0DbqZUWw7yP0kGVNIscU69zX9E387wA
1T5QU/CTcMVUj2ZIzxv4xNFf2YZaKTiLVfzKIWqKiMgWHURegDwanJqX0t28T/57
C5IpHVxavAfq19ewje8zyFF5D8+20Anw/KiTBEnM9Fcl01BH6y05xZBhCbR8eVho
8/aiATMH24m7IIaixifAQ9fdNIkmwFBraN/LZqOc1aQZZGJ3Dw0ZwmuIxT7zlMmB
9LdbqwJwf0KTq+nqIa63fQMTGHd5V8h0ClLnxC4jBstB+9I/m1aAbyQdZHXhes3J
k1G95LPuytGAC88KryZXD8DKct79vU4Vmm4rWf/RDt2T51Qak1bS+/FiTwxjTGNh
k1Do6lnH+Z93NeQlVt1DXkjnxyWjDYDQbj0UHtP5l3y4W3mxNGgwV0XpofHgsZOe
mXCPUbbLPmKB39Ms4uEi4zzAlNl9AnU/bZB8s6JMtLVrFhYK9HgYHpXDmjMvgC20
O70PF4HDaLx/LGnZjWW/XI3Zs+b1u9UM6CqjDk8tFFSLhA7JpKvIbfVVT7/7q/Mn
44dRCRo+2uNwdQA9zxVNL83EAoYOmYcw4wkz8W5eWVIE8wFHwocKqzHMXvtVM5vw
gdoSSw5WDNIW3Immmu279T+NrLV49ttZOuDADlQXYKf4PebdPtfvkFbDbFKg+lvz
0yWjvlv+27AKwcXjgUq2a4MQPPG5Dk+4nWhoT/A716vRIyGq39c4pSFKi//z5E1Y
2VlHbcw3+Rtvc1mxaHX28c4zWdvnJh+HakJ9UYiYHo//3GGeAoVPuMusCtn3DaXA
cYnyz/kuIgUVASl14gcwTeSJ3QH3PGMLpk1S8wJZCh7opc8vdWheSrr/9Im98YUH
x2toXpL34E+qO5Ti0+SBCH0HfEBW2V+SM9xbAX10MQTvdMt+E8ZTZDrLvPJXoJNZ
nveyjg+jFZXB/Xmi1nRyiXdwrTUnTBR3tklMxX7bhGqtw+2rJCjYrMo5HUNyZ1pD
0Z6hcaKcXbrU1/9NtpaTqUSbVypY3b1XskzJAmhDNFlWzl6qjaMHfhFls8EGePD5
qqNKWsAdMkEFbe7Ji1jeo04lCmAohQl5/S7fWouxO+J7SiCSQ7DvxDSTit483Ork
kn+QDZGVnph5cEcO+B8kuSabu3xKvUQWA4k+cUdA8I1eE39izEb4v9xvuHD55q9A
SoDFb0z6eRQOztY2hHyQ3hHTzDPbNBFe1vUBJfddagdBO31Ems6jhCnSBPOQkipS
wf3J7b8ePxlaVMVjw5aKAqQTUs5dSZE65dL1is3iB0x9g7ZV5FHjsa9aot8vg5rq
gryRQm2ogpKS6DOnEpoUlEOeAZUF0MA6ZVLLY0/NpEvef4FinT7oBLNgppzZK3c+
VaAY5xh7GVjmQhBOJjdAm6XYq+FcRbGy68Ab6/O3IuhjKbuIplX/ucZpBRKjjzxa
Qhml9AxoQM6SyjB33YmaAs/dNQwDNpYJOfVcT25r4FEBt58qqFxaP8yo+yqEihv+
Y1+VN8R9jwJnKTxXd+x/KUgJokTM0G5dcrWQn+MYxecfpGLpEbLTeemkXU9q7kGU
SR6StFM7niT/H3drmlEPpWtPyeMURTGBMi7P48lmTPQREU2mW9woI5g5cQBoaZCr
Dv+GOBLmieUY+U66KNCXA3xCfOWMyidTDo6c+Dh/TZC6MeEfDZFLdq8DcZ12uBOQ
/bY60zY1LXX1bRs2zi3Oes2Xa0HokyiuJqo8QxfHPYDLSc+8gKLS6abnzkxJEOvA
OBGgDH43Is2rSyM/ceNtUrK4r6agItrOF2zU1pxSX/bFIOIq4tqG3xRA67iBcyUa
rYKpBiZxtWp4EhZXo25dpZMqxwozC/uhf3FXTh29bxyqs5lZA6ULfHx5y7qYxfD4
2hblECdGSUSeoriZc7pIY20xmabk7YvjuZyvItGSN+17SCuNpKMD5ZoyQDPTueJD
GALA9EhqC3Yr1OaFw0zMONNcxL1W/dhFyJCmYccVNVGyKwevn8BqDbl1GPnvv5SG
4Y8gCFD4GPEgJ3DRQ2CMod1aCaYE+QsOLpX3fcgSsv06PlGKSFkQJkze+o7BbdyZ
p91V8i0MhCq7Mbu/XI8s6tvH9k3nCutZfAPrgiieE6ridKhyXeXHFdVdv6IwJLyN
lnaFyk+dWH69eKVOIgosOfD9ISQrXpWXgJ7xkiZKglF1MiCdT6jt5OTem4xmd5Dt
1yLHkcYLZ4kpRwGEiNdIOZuVz3btpiX3RyEs5U8/SPXYBByjJxmFGSIEqkuweglC
dpEe3dlg+fhZKg3I+u5d/+rwhejmyN/zmssUIJ1O+2deJ7B/Zrm6WSMaigi082zy
eA2HAhIcbGQdsideqCdQ2NH6kMS1YYR0amnH5VA2H3lokiGN3izU0/wRgHJXkF4Q
mSM+s6/JlzHcHtW249JzUBwy/PsOESRrGQ0bqt4dXTAp0uV35mHkmOJF+khwwFPg
ulugEvef0TV043vEGZ9t2j9QYT7shTASy9UjZ1iPULiibepuBt59WChLsjcz9cFU
hD6m1mn1VLVRi/9ZoWI1fRTlNt9/hN6cV0pHeHFqoA1OQOhM0GWO6iuzZZf83BbK
/QkRuH8LAvuwZNgKL1EfHZp+A9DY/gWj+ykj0eQK61/ZaaaTm4qJUP/C7ZK8iy6D
EvsVJ9z9uMfpBroYIzSlCWJDE54obfKzP9vaLvj7S9AdZ8iGnWzaakmFoFX4+zmR
rGpELiJaCslv5F2aNj+2wcox1un/gBTj7xA3g7L0WHbKww+ZMxa1XNdh41EIeAPg
VwZtJJj2VP/F8vZiddUIoA+hXQFk/Yk1EQcZN3XJb5O2H9H5ueB7ToLV+27J4iGR
uiBFPUX9wJd8MFScfNPHafs2s8HVOqciciv4YzQ0hV8LrGQoa7BxU6YGmBlMPD03
MHn5APGqvr7uu/EmKbcT2Xc3qvtLDfHAlPl8JT2berWNpWygxQwN+CS+BSb65BSS
0P4wJrBHShrhge7dOlhKW1IJ7omCCiwZQsuwJOBiwaDldNWCxMT8I1mXg/bb1+N4
/98jPYVcUtmawkRwnqjw94SMss6u9FrA5ECbVzvGmiaI7FyjB/vhnajDHTOI7k45
+2mJo/u15KAAwxtjdiBVd1bOxdZyetgJd1YVPwE8BwtCYjW/Rhw7CFLkEI568Ywa
rYXjF0uqpIPg45jvB9w0Krkp5fOzQ3f5Jt9reyTQl0eyKxsDYlcac86tTfVoRhW8
Ga90cvDPtbrHKb23C2wHEtNt62Tv38GH5mQCOo2akA0uSBc54nkZ6jinjFIvvsyf
y0Y7Rj9aT8hOU66+MBw/NjLGdoT3dE3aHMt4LKOI8N5JWBJfhIHK8SRYKPIK3iCh
io3yFDao3Qu+0ZUak6Fi53j7Kdz383vz8YyIsnYNGLRoToLJyo2Q+7inZGHoeJ8n
mWb4mjJ9Nf+sDCD86Mrm5gtMw2bYW0fkuzqg6xSOBwNljSn++1x4U2a/jGD4I32w
UYcq1ViP1J14XU/9SGsp1tt0ig6HWrsiTSv46jp6ib6a3FSg5ixL7NVitwCJI+Zy
GnET0ULtDoYEXvS2y19zdkHmei6dvGuyDlD1sSmY+qqzou6uGR16dt2htC3V7m9I
61ZPO/00fKwWKiE/m3eZSsQDDvfQHEoj2QQI+apvwY2+4MTaT3GfsjbSSf636GV6
OazLjBKavk2YJ8iynxw1uY1qRBRztEhfSR+lGC9zLfRw2ovNXJz7/GxfBHaDQjSz
+/tStkCqpbxLV5TuJy0lf5tefeyZhLamIt4HotPkjV7y3w5aWUYnWD3LIggpjGj8
cnIIFkWf5/j18qXyUImIPt/Zhhn7+uy1LH5XcxQ5jdNkrcly80CJF7S6xjQyOGvd
AZKQjWKNJE0ATvyu/bn7kqbhWC7OAqJ9ebl9+9y63nNsKv5RV8s3Os5Sg/3ukaxE
KJMrRUQR38B07PcIXuB4lJDuju935dbbjrSW8z2jPwsu/35oXmWvmFu+utyaTpPK
fCNaJ/pF6ikRsChwSSksQbF1Wiy5fAsAKp7FJoTsBw7cEXwakJV58O9Brojf3TJI
cPVUDlbrUhsXHBQIbYDSR6qINs8CdoYtS33v0suwH72QV/AMEaNFgaAFMEpHH0UI
0L71f/yvMMnJ1VXzzBYqkNdg8VUkFKoRC2aatbNpzC9uziXFO2woTHRaXRLgs1Kg
aKD1Wb4jZq/6B3dn24F5wjx821olP+r/9BfPGxNDxrXhA1kRtzssfblhAo1jOcyz
gqb6VUEE6aLV22FmImrcjVLlHHPpkQv/QN2MFGNcmW27t+m5ul6U/xgtqdg+WfQH
0mpIarlJBAEWvtkTB2/3qYKFWFZHhA0jLjduGvJVR4FYq2hWVtMD07huGSO6n3Un
xc5lO7uPXFXTpjkKkpv30GPaHuRFJtmg6j+AAKPSxxivpyyAJ706H81xxdMCKdQ3
xkLhy8pRPUxd+APQ1F87RbE+YSydjYLjEADSykf7lz5A6vggpmRx0jzGgYVDXKhv
I/0inQiFPvDZyEO9ZGnutgXImL8whjcLTi6W9w0HXUjR3ZELXKfAqzk/34DkwhCf
eQmPOd2+pxeS7x3zctibF7wm1SwONVGXvQh2oLLP8rBnVcQMo2tJsXFw79ZvNwUt
LjbLsPgcYV8CYy1S06DBdzf/AtFDhUtmn3T0UyvtOe9ijsZMx8/t83oVBx+8n75H
tp+5H3q2Qeu9ckQE/CIOrbMDCXsCwUHDyTRfHkVoS0xe+9R0kl9MrzRmBJHETCUH
UGoFcazsnP91Lh90ffKntQaQoKugZTMq08Kfa62ySmUl53XCz/U4kC6WyGoiO2QP
LTm8LLegAoNMfgmaqXilES5OtP081+s+jlwuuRy0GMwAUTmBrwGyyJxi7BvUFRGK
8Rxpak6U3pO0T7ndcZlOrZOqfphSELz8H2fWQdby6qSjP4ZV4pAayiw0nK0cN8RG
SW9ho45aY43X+wBXi6q9KPzzWdbrOp2pnBhK8QF8+7Ik20mlVTqnP7freM0bQBQA
c+fWzpp1i3w84Tqrx8xl79vwRv7tOhTZv2FtLXbNVa28n7qPNWoOn6NooPn2GiXW
183LRv7TGCWJietwzIUFKXb52tQaIKQULNBcl2DilTDi3lQDWYBbnMCNDbYC4bsK
pimvNYJ8jV09TG2KZKE8+QM2u0UWFgBb/s7+WLtrMb7y/7FfmYQIBuProgfkkVNy
nfpE+IBH/UJgsLp2Dr9c/F050CoR801Q7iH0uv88qNgIi5qNusfhMhWKGhILEqwB
hP/ouGaxYdGVc2SHrDhhECE8eNF1XCNBKCilet2DN5OQ1Opl4zXLzc+83B6smRyl
L5kkKh/eMh9/lKM2/+vwNC79CUCNQnRUQeh+Q+9TPLDisEiTmBXJsBv6H/x6jlQu
lOcnXniyN7BA9Vkhi2j1iXTB49Slj6F+uFtNPn+MarN2shRnWT11o0mBj6xlux/m
3BTo61+7G9n6DYl+48tCpouy3bMX82QUzSXIqNh+ncAv9x9GoZ1gljHpWmtwG/7W
sHb3xVE0IpwcBk6bS67Efq/RYHiggtMNxaqMrFy9QSkl2ipMibnpWnnRusz0fmId
kFkcGNu9/8i+yoEx0Wx9fGcBWdDfLbhmEgaFeEwRtTbPElheVDqO/wPcQLcBRoPK
dGM3Ia/0qV2+ZpSSnmseEkMOS8a98zOhHj0hes4Xfy5kycdcRlX2pVbIwGZ0tF6X
/w/l5U+FABp3g6Frqwh5W79whrfHPtVSlDv59xgMK/xN48pdjdbgxg6RboRvkfSd
NdsXH2qB6T2m4UUqeJanUCF64PdvpBhILdUvHkul6EAtRpo9bHI+zueX6glZ/EUJ
VSVa9B8th70WAQJbb4Q2XnZG0KE67Uhr+Eb+MuG611DfUVbEEElLiJMKOOWalWzB
XQDOUi53CkRzXzpnfXj0uZ9sKU7MTWU7xTD6N0GqZLS5FkYEapNfUmv21dEqXFSy
hT3vR0xBZAvmY6xYRvHO0Gbh1eQDkawb+2oYDcQGdzOExdBHzm/bC5cWff5iqg8W
EIUiCbTmYt9BOgp0QRojJXLsgxts19Zyg9E7OhlirrYntEECWLbSkTcn07dlYgvk
KgHVkCskK09SHpx5JsaQDhthYVDXVKIlEzjsIwVGdLoSfdtyxAt0Sbv6fbfIp5R/
JFCvGJ+JT41+LZfAoOp1MyhLqqrusWVXnCVHBJBmuxs3nWNNTUJ7g7bHjFNaaCSS
yQf2vp7FneJ3hYB/PhNSLgEzCKWScK3QJ4TjZN0xdajOz1TYm7MknaQbZZ6wCazZ
W2QHxdMepl8EyXY9AXTR0R47YGXzqDQ6qtQBOoo/f14mWp4Ce7lxoOUlDAPgQc/n
/hnOS4XLBX12v0SCuLS/IH//sYn1+Ccj7SxnXhyScmuQ2zR3eIME1ypEsc0q/HrG
taekPL/7rFDcEbVv6KDCgFltQL9OMmKS93tCNSAUY6as8t+p8lspAYYgd8aNC+8H
L3vtjxYf8YbE3/uXyfzSgqxtAQT8/q0FWjuFEdaJD1A6sOJCOLni7yuAYRcQFik7
oI0RLnu8IBbgwDXr1GRj1kUCNjHcorGqCxsxyqRhA5KoQ8RnlaPhl7ajKiVrzBHO
bL2ron2aJ17YWvyWPibc6axgqVTBn37uSRSSFn3Gvq04Tx8xerWfsDutfVy1jM2/
syZlNZZZBh6NrcS07HZ37Apg8UMHmnfLkcFi9+P7wqnZ2DDLzZEvgH+uFwXAyuna
Ya09QoWZxkyyCRLGwNxAoTrvA2c1xzrHlh6intVxQlCzWDnH72GnOGLI1Gfxm2kL
3uwFL8Y6v/KesICMf3kn/TqTyYIhE6SKtkyZtUosK2oLQ412KjE+bIJjREPBXZrw
xLV0TYUoOq+Zf/tqYxUPA/XXcIJgUuISUZXIsDgoOVd04egCG3uHkz+x4eUFlNG4
tItYHU5R3WVj+wN6ewMQrdV5ByM8D1lJ2HbJaO4CWbHHtr9ARzJHsOVg4x/kWkIu
EXW27PoSPkYl6EGTQWZXavLvx9wUYAyT4Or6//hbGSIb6K2JLjkdQYKFsKPfLDQ9
aUnaXFvMSTG9m2kgY5RkC7L/er0yUUniWPjC4AUsRo/yiHTXBUAlGQJyvyHm6uSF
9Xw3+datglo38c4bkM46+RMALLYWxj8ifBmRD2hUfnyrKpxYdjgunIkQR12dekHQ
y6cjPuWU0g+rEu6cFN690qVW4hmHU3oD7Oqdk/zeYzRhbtfIJZDWIBwrOfZZTgnS
U0suCGV1kT4Oev87rAjYSsvQ9BCY1MxFw+a3QA9Oo+QbxuLeCDHfUizUeUrdtJd2
v4x9peEcojahQXJDPRKP7bEK8aH04vvvsFm7lbA/D6wFwwBB9QMsD/jFMOs06gaa
JmR/Ncf3eeuoPg96sXmsVxVfhdAZ+qkVHDQcaQAx1a/S2WkEkvwncCCSbB6JDnIp
peieL/suwojdbyTqoRAhL0QDzRafk6g1wu7tlfZAT3jINmkpfmwWoNj1dnfjdxfJ
qgyEmK1T2GKHYU89vYyY/H/b8AYbznrONbXU7nASIkEWAMQZYKA58FhYgX91+k0X
yIP/OhVgrAx/e1wai4jm0KWSST//hG5r5WvYpyNcx/8Zy6COfVvF7WwsR5OtX3/E
7bWBXhCXPuQELD52N3xFouE5OGLG2Z6+fcU0KSFbIdKJNPCI3QTRZmcnqlQFTVqm
2podblq7RCDHciV2mT+bWT6mV1cZl1z6fKXhmNJy2cvo3uq3HP8HRta7PcAn10ts
v1aWUseSPC7IkB4zcBmKBI3l6s0v8X/Im9SjEaQFj6PCbsFH9VXOmhGV9I7iXfLp
eB4t0+46lN9VCUo+iugm5/c3STzhz2qSJJShiH5MuJUm4HHt5jVgCQrFTvwuvxwS
GsgYpghKB3t7CeAhUoVgGHJBnbU8BBvlWegqzIGCpy/2Cngs1r2IppSCiYiOl+FZ
N8vzpFm064pAfeaJXWWMcviYDGrg33fl8ngFC4h8fVX+kz80K+UA2ihd3IQR6a3o
AoxR0Xc7z2uE0q0chJ13m4zrh5cvyOF19dRShA+jQkx1jVGNRJW0D44ICLKdsrhA
8qC5feqoN8LZ1GCAOkUYA9mXzA/75m7/0zD0E7lUN5VPCmVooXmotN29DM4xdiWb
HW0xLMK/bxTrfh1wGk6NhkobtXa783MCVkIUPlKKXMN0dCS6l7wMUskPMk6Qb6eh
d/vLTPvGXevN+f4baz8KQkkI+ozRBqN5Kn6wSca2Lwgc6i1PvNy0sP/kL+QP5UN7
N+pzsAQgN7UmQTa/ffs654b+jTzauF+TRbW8XH3q3gahd8As5lHmWMRN0mhETcIP
vzK6xtSCdM7heOcMbASbNZjR6YEQgv/RNsDSQdtsH5q+Zu4HZXiCRSqXSYes7MvC
3ME46ZGqISnLBOTkJoqYhzfk01siHtLsk525FQfaBNrGFPNQda8YzO/oNsx4QBRd
9ApNHkWEEkRlpH44sc5s7h1o41I2ZSoICp5DpglXsjQkT+IpTHTep0M2k7LKI+om
ajNoSpYLaDyhReKGKeyPdZ2v/IDlkX4TG5bn/4hz/fP3zzc5MFp2E9eDKzp2UKPg
GED84pk94CZVLkiR7e88LOHDGN/dDj9GlW+rJQ4p2Qo+IJQoU389qmmQkxZV0Tm5
CJ+nQJPIeMV3FSQMwttE/q73heV8jmPn2jWKWebGtOYL9UnkmdaMZx+QG6pH9KHE
0DxQwM0smsA2VJZ/orah1/98dd7urHgzTkP5qcVtqXriGwgt+n4r322menHm+Pvt
UFCGWCZ0QnuniM4/uh43t+a/eslFJS3s1nQoRhihmvicX+xLPg2qE4UklwPFUTeY
apUauV3We+XIWDR8147AIvbP+ogeqr+0Ae3Dm7UPMT3Ct3pwz/dBGn43/A94XbhA
Bn4zI+xDVGYxt8OjGJ5G68wEDOZOn0Gip9pMvC1HVu3ZaeNCa3EjQpNTZUMPWsZj
rt+B4qgazQ5yl6DlvOq3oFvrbVSYWKvlEey0UcBUv2oqrj9Ynh73BzhbPN/UO1KW
X/iWA32DZURy2h3vc4sy+6mLya0LafgpW2l4N4C1kdlN/DWRKX4BOdSECHFJrPyu
d/jQ5jloxhC07C/KcmOHuI7aMesUnj8iOT5pSr7hjvmYw24TWHroCKgFRx4PZM1m
joCxYYJt/vYbpA+WbLCyWAcY9aMGf54MoNGID5X2oC7HNhI2qhY1sW4dZWUsdfhG
iNz+n4tUtYsO3gAQz8jFaoeer7eOPKIIfyV9hJ+c/9yZtfsHwUxAZm8MPvgC9Tkc
IOOMMr2RXfbmzEAxJjweg2HEjExXCqNX4wBOyOKnsofnO6MEk2rbn4BzEC3Z0O6W
RBu/doSsLOpvluMitM3eGaNCmnWOFfuQKObnxHPyCto+aDRW86JbSbmdjVineusc
6gtxupgypPA2y+Gk3pGOd4GPpl09XEIIWsuIlaEDGt9qY6WGxPl/BQREMT0F/Lsj
2JveeBp0SJhqQcH/l/srvd0CEq+CDo/F0Aw/oltIgZS+dKDFEdbFHjm20s1ast7B
MfHWoz9+I3q89GbwywdUfaxA0v71z+6AbFJg0FMmiemsNi2SZIlql3dWPVbFXxXT
CycaADrNY6QbBejqsZN2P8DHr5t9shs0z7IpIHhqe/T/FIVRX26Mzl5xyatDeRdJ
kI8ZuaNyeHt80x2gH9ZJlBRYAmZjEGeA3CQBOY/mDVH2o99IahCB+Ozz8OQN3eOy
6AbjAC87d7hGr428tGb4xcXWir4zW4FTIWLc8SCxwF4gYxqJ0dqleuQD5kaA8MvI
wBdfCVRog4xhEvwGboPUFB3Qr5u8cplBt59uGBdydt25keIKc5zZNGw2C1y/0/8O
jwYhz286HGh1x5R97JROfIGrzoS+GEAUYmSOdWuGpI3AvkrP5D31x/6iMoosp4uf
HzSPoLRJI3pdzl+lBY9JBOyzrp9QN4ZJ4qhgsX8aqHg9Ap8s99LE5/Uywer/NHjr
5BUwm4J50/1w89a0Mm/BX4cES1Y+g+vpQx2V16OEtX10zWwYe4MewOLUvhmlUFmj
0GvNZsPkA7eDd2rVU6BCBaQ6KnDkASm66Rxff5zskbuHIKOkQBPLUrDSHuRXm70q
e5JbuILi24pwGjRGieY9JEiQxYIaTfYAGjnBZ9VzZm+Byqac75k28VpGVNqLP7Tz
+y4AwuHF+22JbSVD8nJq14SP8qs6A2kDBfsr6uGuqrZesQc/sNaY62n1KcQyNxi/
+J/y0VKgDHs3TVyIY9NUV3EmFGfqY/cvLdwXxeiJT8qLS+Y+zIQLcYBfLvW+sgK7
af22KU5EBlbGOHV8sK2/FcF58FsJpLKNYBuj7tJGROQxo53PaPUSM4JphxghZUgw
CmGMbLP+vN1xs2gLjUPq7VdtHx2G1PHsHjiJe7aWBVRlSZFwvh2XNi3TpEZ+8dQv
vt100UsjBulUz2NsBTDrG358pzCJJ+y35dWzOC/bSyihscwLCZhwH4pj6M03Ah5S
o7hYgpWRkBppHtnmjoDs1C4CYVZIsIqru9V0Y5Z2ynLe8fE7wwx+9KOAIMgKEgW2
rU4fXRK1Dp38jnnAQ7/jWjsIGbuC1inaeZfu+G2bAO3DnVWq2wJxkqOlR7CjUf7L
xgU8edtPJIgOwY+pfjpcbh0VoTj34hYkHlCux9+VZ5d9MG/UdRaGURvTeptgLWkW
XPeICRG0J5VzdGg1jQ33udE412ZoLxTPOXBhjeBKUTGQo5Qf0Xa8tPVsqkBHwHiw
YjfIaRL/xmi/yjy8flZMM5rm12HAwBSe1BvQrxUWhOOXNAlKvM/0DsLGfxI24OUL
AsNyRT/vY/+vz3oAFFFJFMMpLFS3vLdaft5i8nHPQqEjigkMdO2PuEOR0r8re6nj
fsH1hLwEUoqXb/ZLCZwgeyYdpZjQP3rqOWLzAEqlM+KXnmbf2UAZx/HFrbKXXk70
2GmRNBVa7tmEgIC/7HbGCjuBhuUdMmTvdMg1XwAHrucDr5T3xTOx8pJm7LQFI/hh
h9s1F/W98peaLGHptFTdaGeYti8H8mn/o9zJ44cPFEMYIzasKZdi7KHMaIDyYgVI
ivEkcu0pODqrrh8gwGmxiPKwkxEF8VMAODmaMF9nWwGYOtAAfQZBJl0VV2+pQqen
APVxdC7cVmGnITCaBaASlNNGWAvlRhu9a4nQfaML3suEz+mHzLHO2M2FqfPYFVCg
0S9cO7rnnL87lkPJY055+dO9Qy/psiIknExOIpZo1yFjSdVcg+DxlkynQnfrwfGK
lZYlZnP75J4jW3yhlqfsKndqtTtr9aRHHdeAxRGYqfkE1DaD6GV5AWTDS9sFpUkD
57LiaBGwe+E8EFmt5SMioehg4ASXGAgRm5kRd62lLIvLyJV2tKXRBCApDTP0yZk0
NVm0SZ8iPxoikZ7NCVXbkTmJwJH5gnz68s6/5w8MwapLzevmsk7+MWOgHufXOjKQ
+4P9OkNLo3DUl//OPLa4yOsL/Jjt0tx8NkfaR9cg4Y5XnVFlzsfEsg2+NRByWcSr
OE4wY6plzIcYapvELjAg2OXK8CX6I/nQoE4KHNtflPbRDklwDzJcTHSHJUGtFBC6
ENUMe2rzT5+Tf3ZjTktLETM36koEUDPVB7Anmvwoc+EFUrb4CIoazOfr5YSkJtdV
jxJFR6+snGS2mz3hEQHtx9vfuHp3f0UnwqXD1oLOCuMa3Ui3DFwjeZMOqoldK6KM
J9rQrqsStfiIgIM0Y7RAQSS8DlL/hFV7AUcHEmoWEcgEEAVlZi1IgvgAc15+1GL+
8yVVGj4nIDAcrmwA+5wb36WJRh92bh6T4NMMgslLJ7ex+r/WbEXiGx55jTQ3m9lw
4TubdUkBdle7dDIMwuv5zUzZU10CqSVkz4BDiVRTcRxpWnCt/+kLN6DgEjcllhkt
S8OrVkbtMcI7XHU1LL3DBp/jaPH/px9BO5UgGyJ83YBQcbwKcYpBDJvbN7To0BJy
sx6M/vOWDuRWLmIb6J5hxA9hA3++F6UyzMqRKsv4t1GyaAX8YCS6mFyiMuU5PMF4
QfeogHhQ8dE13RwGCAXRmuml9stCX2//kjgps+amJPWRwD6EO5smnFlBZ3vuM8Jq
Pr88s65SOPaqnxVdion+Fd9CrzXtBp8PYlSesBxg7gm7LiNBwLR9FRvO8K1Oez0u
yPFPcueWzNQJ1ClJysJKuR2TD02mBBGRtglsuQ0LnRS+KtJaP5++H91E4eTM8Ji2
cEUBtqtrb/QoUwiotqUN3/I2iBhI+H1Bd3rJWV738OK7DsoLbbegT5PQ0jFuHaEH
bWZtzLoVICbXn05n3nsGGAKzBvDPcyUEIekBYZA4FDVjJMerriqXd8gwp4RzsXlp
/7Z7tG70GtQTW9sC/JG1Wd5EsT7WwFv3LxG2en2QJF4UScIrHduBGfDQ1C1/yE6T
OiCYuhquteCjnfN/FkvJ6Cway1Q7gi0X+QXelibppRfDNjp5il2mADItHABwry+4
4kBxk4X7IRy+0GKzqFcyUzxGycSJXAur6m84qI2txko1biOzbbGscJMdOjS4DcZs
JUqgrXECycAmSVHbSn301yCzojZE0ZDpQvQRxlmxWcCY1gdbvJfkPUw4a8dyGiZK
r01VDCjDhc3KXydusCuBdDFTR9C14nJYJzkNNjeeSGZ2980RK3Y5Epj3r2cIYhnN
/j+tarfDslKrog0NSMi6qua8biuNxnz+shwTtT7I6tTLLrJv+8Gq2UHoIn9nQDFk
zvPUZaYzhQgX+6iDo26+vwlzX/A+hmALmJsko9/r3gKPX133Za5NXSOtsY9vXEib
Gd9R1hZY9L2MgV7ebJYC/5h+yLjtGcZznyjcBqSK7fT0nOSEKwjgHnVAZRcUYjxR
gOUZnICL2bVnBNI6SvYLPY/ws+2dHGb664C00kyEPYqNSGNXLCwWjYO6ZKLCHPbz
FbdJJyG9ziiLpZtB4mYaC79NP/8Srw7wboDngUALo7k15QkuqE3J9BERGdh8rPNk
xiGlmJVIbnpHwBjP1XOQx5taaPXHhyOL5bS9GiACZFWvoy6jlP2pKGTVdfZrOgpB
2ivQbBN0Y7cgNtN/eIELQtePsuSBjZQozUHwn1DbIZ9z3s+glS3wAu9ioVigegJg
IIsOgCnw7euu/hfkJzeHHIuZBLAYl5r/PNRmu+D3QikR7YxpYCpczWQ+8Hn4zp0T
rgffb7FJMgJLHYrldMOTe2rJNOGxpokJdBytPV9iplMriqA86gJjNylXs1kgQgIc
JafuDESvzPsSe/14FzAZLY6E18u8VvOhgzOqnyS9bkTxraRNSY+xPo09C9Q+BNxG
fedjlPDTnhJoAuSciZtYqubRzAF7e4cr0p16GV4qcxWSiS/8TInLlo93pApiCRei
cHA9kTnDm/bKVT1ngVkrkGcWKFtoUPmOtpQf+DL9+t/I+Ks7U2mZeC8UjPeShMhp
QWtdEyOlVHB/OgNmw2pgXe0N5CN41x2HFRU9clkol2k/KWiS98+Nt1OqXHPDGEgt
dfXzOYTMdzvpTmmWtTJE0fvj8ZtxHZtJSfz22/GzyRZaQ8O66vcL/WIwYQCe2U2s
EucRIl1gOK//WlSHGvR/KbPGGQrh0ckebkOCD/xTL82lCu0DAzW8Y5Ylwc7YGF09
kr6D2J7TCRLA2fopySJqH9FatIPlyHJxJeUEVGOhqbyJVHHe/wUM21Yjmlr/CuZs
cOrEUK2QnXFHdJO+talKAPwmnQEaZRmjcX+InyaEy0uYJX0Upz6VhteHOpoFdAoK
gU8Rp5ADMOd/zfd/HJ+VLi48zxCfaQLuefFafW8YtGPRvj/1kabajAT8TBBF8hBi
yZT8rHxuieX3tx88ModgfqLmVhRvH/ng6DL24vsv8ev5YUMp7bLGGMrBeUuCETVu
z8UAospTPNaVAV4fRRbLAvLXe35YuK8BcixrJBaDFQc+VFAG60WP5AkIo4gfkgVH
oJM2gFusxWAB+7zW/0jLKGVz9agupLBTukc5CHn8OXoE65MXAKc4voDQaYngiwgI
CiZJ+/RxqpdaAC5/PnPUNif0nvhLeZl137NRWXMUluvM0DjMmtTWeLHzF1pQ0g1n
8jk1thEohya2x156nZC2hSRMHZ4h9xw69xG/nNDFiiBO+Ovr1tqHDsQTRif6v9F/
w+3b/lps6Lz1tusK/OJF7eS2T19eWFjtoWQMSRkSRWP2PXHEAiuSBaOxONVzAnrR
36D42bgMhE97brSrGDMoZxxCoDxuIt9bg6/YWc/i0bav+Ny/w7ozdUB11KnruC7j
Dvqr8B0zmeAKzw/z5xPg78hkE3x8zJGLBHdxd8seBdLc5IwQe5q87nKF9ZjIMXsc
YVlxvyN4Mtopx3fn1mPBv0xGXV+/xxNoPPekBybPLnNFc+oBKsoyBtjc6gPGxo1r
pfzIGweU/RmzWRA3I+Utjx6VYSymlDs9ZliU6Z0OTLia+CIb6w/w1u6/+R9FtEFy
3ujN3DBDtQavTozBS3HL6h1X96jwpMZUId2nqqff56BgtsyQjeSWjcTbL5f2fXCQ
zSoHjm0PXpt28vfWPC5CvnZfuiacjNqPGBoveD9CGPC/3ILCBtMJUbLqUimkTu+0
nif06nLbE18vwBDIhLU55scjgMuobUaxkqJIBComzO3aP7PO5SvIKnYIZXOVPxWA
y+6Ggqf4g7iF1Jsz4YFfv1oHI6VQegxGFGA2Fq0tS9wPx0Qq6W1CfvI1hrm4KnjY
NuLG5OF70VCRkowsC7MHMkSKB7KYZ8V7rwPLWRvMUCe+F/I2ndv0/Q8nfRz74tIw
ZUEOOIZMfTWINmnfl4Z9ZhznOBqge2Hz8SnmZXt46c44dp0lpdl5tcl0yR0iERE2
pv0E7hxM/Tzs4hZ8XwwDwWXaorP9aKq0+fXs7hZd8MPPzY4E5MFOogWS/+sQhEyw
U8Ff1MnOyLt1LoD9rXmlZhTRNKv78ZsM0NqOD1qiid7Y7MWeNV15mvM62foPVBHm
4WjSHhosQGmp81HuWQx1sBeLSMXlWi8Ra/dpfrJfdDL/4Od3ktZ+UKEstHnvIAtO
4qPuk2uAL48vZoHCeeeKqDhFzlp1jbh6VmG12El+MJPpVMJdvoErc77luLw6jgzH
m+XtUrBKINDAnIrj0DnfH9jFS9I+nun5ZC3JTwdz2K+fHjThgBrwDX/8gR1wHkiP
vCewQc1qDTeq1hFeS/JUADLdPLxDTnbVTSgkpE93NR/ypcIu4PQsE7Jyqv4WQFjt
70lExC2fLa6L4fkxP+BwABa+QkDxAwoox8fEM/lnBV/VxO9QaRFLhsC66NicnvBx
P6ZQDBkaJRLIiNDtpVj+bwoVzjeIsh8LqmnDChaKum1By63KwWqISCU3ZliCyF25
MgwPAubclE1WP5XKH7DS8dJhD/fMM/qGxh8y0Sm3kZ1H06sH1C7Q04AJYwt29Hh+
Ox/wYEAFXmZAQBeMVtq6gj/3S9bq1wzgq7/2rNQ6Grl7OZCh7IxE9GNARdm+MC2b
t7I9K+yLGyTDfw11Lwf93t1Xw7mgSC6CwGekV6/R4DrBUrDxXWYWYiBGAsawuQ+T
/GDsIoUHqEKbfvse0fAAeDCrB24Uom+J/QWJ++sA1yIa6VxhsO1K1im1Tv2rIuvO
NMNfBudTcmku/cW0QCPjPfyVj53CZuxdiWPXafky14ZFpL9HjpwU90JEh1zh3xGg
CRPubTp1Nj68dcvkK2QFddytIEmzGI3HVbLSgzvVpOpszBnPEQOJ8kZaXSpAUJfu
lcSoLGWXbMCwf+hbgtPMGgNVsF3fJhGkKG7ogf9JLEITDQ5bb5kltlJyt86Oy2Vg
wR94gVfp3/jLi2Qd2tLBTZA5Pe9/bdmA2OgVFLC5fk6ykxARrzkXgZt0DekuvKjM
oVjNRCZYJruTSryQuIVpw4mCnL/dzU0VOXv9Jo+ijv3ffJUxzL2ydyfdBftDokY0
hkfLqqHtDSqiy6cxUFCrQDfVeqEZoYbqReEaCVJji+nZ4sF2v/zet6caMvwjCsnh
ePTjYMRmh/QuLP7HIvuwJ7RlhIlXwFlrVjMDWMdygj4h8Wvz9bMYlcQJTkbn9Xy1
CWikajYyrVsgIf9bRx56EiXYqAPzNFW/DNls9C35iYV9cWGpfWshN87BwAsdgSrF
S1tfT5+ZU4fiP013U776Dp+/LuIb1JbeJnis7F3mcMzLzmlL+to8RVueKv5z22BY
AEgZDPPrER0/8fO7X+7N3msVLZNy3CYXkRWJUxquUZbH5JXCPfG4uaaKZndLRjhI
pNocQyyQl44H5VmXWEt1zbzJde1zScLIq3EaxKc4pQ7MdUxMRGoFUTKvNuT4x5AX
G+F0ivLFoFCc6/Qj1UGTr0iYT69Dn+MAzDuFdB4G4QMpZDeRij1shPXCAz+TRUL8
mJMS0YyAkXO9WKIZPSNbEnkcCuMet2LYbFCw9K2+i/sM4OGQilFycyhptkK09kGw
yPbUs/4MdMyngy8ft4ZfIXmicjXAL7BwvG8tehv4Fphe/xsaz5cbD8Kv6jlT3ZyD
bPVTRPpcM0arKGE+hVYa6L0I+8LxAxM4HD7N3WuSmsCDHNMvH4TJ0sZESghX5II3
Arnz9iUKTpJpG/bGTqvdrlBf9vHrzc4ledRqK7SG0dQjYL83cjl1XgSkV5R9Xs12
KjWcIrSrG8I4AOPUgrTP+Qc5NvhTZ/0xKtcegax30WjX8WpZp4RGtyQvCXZsms6r
yYSboKR6i73XCJjNFWjEXYsQ2So8gTKQhCZE/P7cQ4G/k25SpufJngf43oxim2JV
AUG4/Iuee89kBxgIer0I3U1vGsCXS9eJuFYvpXhKSRbFZZTnA+nRNBqEaBN73DwS
BzECox6AFKrwb/6UpaZxDjiWLAxAmp5UPucc7/NCYVr4tGJFdLt6Eb0vkkKXCsrb
CHzLV5tBscTfTbb1IpgpmpOeft59yjpTkwLkeXrK9lqXLdfivXddyqCYoQHa7J37
wJPjWatY5wzy1f8d6Jtt/ziKisNjoi7QFoHaeEbT3F4r/y4/3IrBt41Eo8DugOwG
s8lrp0QmmyUZdS0JlcKTn1PLxRZr6FYW++eczfdyfAkEZXhVmFh/ng7qXRXjbijp
iGGLynBJqsH1Ksl964S4o8cbf0HpmYQgIXaDMIXuinggwoAkq4gkyM0u/Q3QXuqY
dAuWOdvyNfyqLm8a/ogQw1eJzZmAhdiNQf55mFjeee8+RSmccDPGuI5StX/ML+rH
HYXTEz9aHsMFajh57UmuzMAA+Ya7NHij/y9UfhN9nNYn+ygfxm2ttLXZnp/Ss34r
GLyzA6zQvHtq0l/ZoLw+ywsHNvxnrEUi82PKVZ3YG6zfNPIW/xnN3W8xrafYF2Ob
lX/opEPy3F+rN1Vvjf81gb62oQhSMkhI+LQCMM2GVUaclmrN2zOHd19XOnnSxs2z
O31Yi+PXPINRMLiF9TOhhx1U3q8vNkW2A8sOuY2RGUZHjg+7LauvQMOlTZLAYR8J
br8O185oKmBlG8nWs2+h6Q3cYja7NkzziLMslm9KxR8DagxdLs0P/pmG4Y+Tag60
OdU6vmD3yjC3vJAifNbHGmRjnGAOTtjfEojlm7wEI3l5odPbXpeWcKywDHyBbBAu
zxVwsdBPKXmrQpXZb+ktMLnFYVtaCkwHysuhepJiv83CW+ruOqRo7dbLL7LB9jVw
chxYFrdwHUOqDOMJcBts3akDhv2hq22WT9GLuglMO+ETfswe1cd7KVUQ62HCdnzF
eH8fAbSqn9iwcFDzWTnfXS/ZPaJ9VyXZRNqo44+iAXofsX7tQJd6tV9EpKU1QGXk
DIjXAVOV+SjP+PUNMYHmj4/OyRajnmJZsSG27ofIlajQKwipcaNR31gwHv2jY1o/
yst4adf0ijW2vhNUIGBLXFJqo02gQh6pAw/GPjyE5pb9Yv3TdD1b3grCbypHAbt/
89zhYEXzh8FK5brs3twSiJRHWjKgOoYJVWEeGtUbU7oppAJ1xkHnQTj1iLnfv5+N
HrQRhgXXz6tRfCj4ybUt/ilM8GDd/Pb8cVuQuMag9gZgCWKJcIBVmZEd1xRHwxJm
cbqafC/lzn7e8oqm3fM8eZEiruZZiAI15IXV2tFnIweki68A1yYJx97TIXfBls0y
DZo/VZDcf6YLtE1CcaBHUNsBl0gUwTokdrWQZ6eCBmhe929eEGExfbdBjM6XshBt
NENGPOfCukzoXNuzPaEJMqeYvpIS1ewfICa4SbjV14o6niKuG43SsHcpyKZoFhJq
7NEFOevTti7UL6CM357xbHH3/Imz5ODvB98R96is+uGEm88IBCMrj8QPMgceM9Qz
uu0iHGp59I1Ep0njorO88Gw4IK4Af78zWRXlYjgWUiz9g+zvfQGDaa1j2rDpUiQq
W4peE3HSciGTUkWESscEU/UWHd4P+J4PV1kRzUAIpX/oDiVul17C4GjaHVNcZVFl
kqp7jEjaNc5+0ErVRu5+PygAJwf0XcW2DTc5gRTpIWN+jtHdFrVBV4Yqv4sz+SdR
c13JqNDPX91KPChtaIIKp35LhUrwRoZ4KaNY5g2adB5zJKKDci8/tmVFJVluXk3T
s/eCHe3bnfxZOf3MYnKDehBxfSLgekk8Ht6PyuQZN9okLymPk0a79EkUgkRn/1ny
cBKbDc9wNSYCbonKeymprRKhnpvDVKoKMwD+P27ZwmyZoEkep0H0/93kkZGVQZqu
zZ48TbT3R8YMwUNzEwsBavjALKZn0agVUFe/5MoFM0s6cLWwL85Ze4YKijC2xMH0
s058SYu7dfQHt2q5ZZAbnaFxxq2MYOuzdz16kORxVVCU30L6pqeBU2RkqO50C+xf
O00fpB8YjDMETSoZbpIGfwxqYoahymodzQW/n9vdi2IVxN+2ldeZXuU+QTGlSuhZ
A3qG1jI9wp6LRo2kMBVXpJphfq59Lfs0w073rhIGYkv+n6Cej6xAjEe0oBMYBnLc
QrvxDLRntFDs20TC3ZsU2bUxpdGg8THgOvYntFBY8ijlOFJE2XKKuc6utAYegEC/
mL8h2Re5jkQU5TWa2sX1bTU0TMCySATUjgTTxNE62dlMPn/ZbSSjf6S7MM+btYlU
zPllT+3pokKR1GKsBIuuBD4r1kNcsptGxGionhiCgWWlkXjAyCHAdXzG9mzOMUmM
nt5CP+cIiwKNkZrI7/lVtWLzCJcC82pxnTuK5Qyor5ZXOqxjB1wgNVSpSjDVM15R
UTiKoDpkXGxh/+7gXkf6n/6sm8oqxuioylCWZKovsg9Mv3htyjdgLcsP5nk8gcNv
Pnkdr7PcSH0ynljwfoY59z76Wj/W3FhA1l+I+mFnodfu1vwINmnEDQzExCv94Rdz
dtGycc1v6DTNAIP9jbOi9tpY1hzQsBdtLtrv9e+HQ16g2YZvTe80ecDDiY4w8Y8W
ov+A3xdu3BemW2xl9baqhkrl0iLjtZTIIKa5Pawa8q9rJfKjpRHyCRJEO+L2Ibq0
zCTWWzi1QUzBBMXS8UEhfu7aNqBirvMrp0rncCd15VFLNPoAiylkLPyaNGrfH16t
gi7NcF2k+BnDAhQequ5hAGtHJJw04kV4Kur0v3UBTJu19afNuD8AQlf7xwY6eLde
ha864knQYCre6dH0u5jqOBtw397AFEOWOUyUkkd+x2BeMSi01qrJ+xmXnFS0h5+C
fxZjrW0O5O3sQntO7a+shVZw1yKYqVV91fZSuH27Twjb/1JcHXVGGuzlvHie6VUz
+baPSXNdoffsLe1AA38TBoI657HUqstkHaGTCdpcWxKjaH7qQSOqgiEkiSqdmusZ
6jLgzOX97iMV3rv59w5yatSDxBOXA3AolGzXaQi1LbNw2zrPe1urnk//F/Bp9ftu
PK1BqkEs4SVMaxOBTsBDIfZ5ytyrxzXzwxfX1Dcua2ziQEyLO/J0YOBpBdBWoq0P
iy8CfAB35BDgHg+LvMbKnPaxX4MHYt1Z2+hgD23UovvKwhW/eucTpnFXWKqFXFDp
UGTWqXAASp1WlPka/xw5ZQjpIpH4TBBUpYj2lNEYuFoKdwkUwCsDmkSQXHg9MHap
gZ5RGTEJhNq+vl1mGzBU3JgYZ3izTBbDLV+Hz7LGPNTmYR6wpGltrypudiUQWF19
KnFhnZShQzgesYUyOPcVkSer5sha/WaD5jG49PBbgebOinXoAdtSCy/lBMEUu7bf
YUPx6DejiepZ8UwFRL/rXy0xUSvT32PpXz8rXUqnZqC9gKB6pvjmpL9rq2WJZJvH
JZn2Sh83RVNHZTxnukNMvQrE34H78CGvLrjkIrpUHNIT6ecFux1OSYZdK0fTwRvo
Hkzndv7AKzPc4EyYHTbQ4PyBeIxDx6OTPRbXLWsQZQX0d0MLD+ULHKppsgestnRc
OZqoSX/37RVdAd1+FlcWMbNxif1gXb2qvBVSH0z2SyeZ+YLqRejvEpMLcXyCNgpj
nWtNzI9iIiuYJZRs01tRjlsxX6LLkJuwDDhyf4huY0dYwdxz356wRgixIoO94oHL
QEHsfBiHzVP3uEczuJlynqG2bUweiyPlaKx+EVkcYaAoWhmz7MgvMxRIqe3fXvvI
XGsTXLQIDl+WqZhHi/Qhph+SeVXaNVjRoHeCTr08ikyUaCW7DxrW1Vnq4zeOlfVZ
DD7JtURhexwuxF5CUVBibO2YCd20CnzvqPi0wDLf5e8/DhreT7khj+tFgAvpI9QV
rduqYZcjvSDgH0FJX0fZDqzDR0qvrrP2P5fQt7smq+s3sRamAvymtc6qIiJzSU4S
24EW8mBf61imkVw4GUpUE4EbaMc/9mS5EfHEnADmujNnTUXCQEd4JvJ4fTEXPZ/x
G/yAP7qUqT4GSvlLVOb5fGbiABtHb3jrR4fhuUJ6UeTtBI+RCeijscNEfIuGaXDN
o74NiX9fK4c/dQ0PAxY/pOMqkC+LiKMm26RIhmsVHc1ea7gTaP+J3uE1xcDyPtTG
tr/5fT0n/ZCMOfbO0A0Vns3lAk6d4/z+iyiSrwKnGjH9wMg5Cni3tJF32icMpd5Q
qw+Ijji73WqmFvDLeHfzM39f5Wvf0gq9SsRDIoFJthQV1ytX8nXYgEdw5aWPHG9s
D7wJpt4RNk7gWD0hcfDP+e7dMBAaQ62Aw6rjUg1ZuFdiNtl5nfMYzeUj8VYcReIq
9+73Xi78g5KHL/8J5WfZkfmzY8NlVvWJc61o1QNi92iX04gtOZYmqLAWUaaJKg84
tYY4JNBqB+TlcpjhcHFlRysKujcfNa7bgQJanfxtvUWUnZqGx7pBrao4XdSZf7Q3
826eFwpFlWttvU1OQxy7vPO6+GLC82HF91+ykPCxz1a0pzZqYP1Ep8ZCcyATqmb+
NP7K4f52wn4Jd+6abSvVYeSUT8nq/g1HVD1U238iCPng7yy1L0/k5C3h5pYaa/Mr
IGmvDt0ieUOR5s8tevqac0FXaYx4MTbTxCAoIweG3NeXD7SZVxDotkvsudFl95ZW
9upYqilQG4YrspmVn1n2J2/Qwlzakv7249xczLd6Enl4Y552Etj/xQSCZgLLpxc4
V208nqqJu3RDWvQMLS465FKsQHj5QUOoMX9NN+V9EZE4O2RHBKOX5Eq9myHafFl3
qwFf1BtbNKmcEmZ5OfcWfBlJJ0VLk4SO3NKq3q8x9+erIDiXJ61rjcWlroeq+XDg
PCCKeGG12yr60bWSD0EqJPm6Vu2ZyyH2W0JwDSCqompEVuYKvyWsvbE7qCBy14uF
PclXDqnyIKEzB/aA1rsLYP397qNbxnavmNozsxW84O1BXu+ZlDfDxj5f/GzVub2d
dMicI4usgti6JlEX6PwSv8kridYDKyHfZnRg+NIogn9QIJY9xz3NgL5bLVIyhWei
ig/T22XZMQWuZRcBobCcG97gYC1YDYeQBTPBamLgdB5slyR3hhQZkae5ycnJaOov
mmKHXd1ZFWK4NbZamB5mVduVVM1hkCGwo9vuaPDwH8nyr7ypdEl/Jys3QIiPTstO
UukGIm5SXKlDOOiVkTk4CIH/dy6MSLvMtbUMXKQOZaBpu42Qr5s4Ahj435xOQjo7
x9YkcacbCBTXhgWhhCsHj1S51p30lSLq2dlEyGHpdqkAF2fAlRIR5cc9BoRMhez7
fApn94rwwL/JXcPsZSXii3qXmr7u2/NIAKWFdhnybDgu/YZw3I7WmaXWX6cEOPyQ
+dhupFuMZ68vX+hgGec5sUHImsujXnqV4GUWeT5wveYflWSdqipU9OKAWoLRwtiW
MUbb333Qlg5e8F7vlSEcOm+bZsPl2kokKTY8D3fLzO5V3SsU9q5xNet111LoD7JQ
b3wXi7+A5Se4V2awzhSSoYM9IG2GhehmYNvOg+BmXqosLbUaSWjblKg1bzWpsAry
6gthukb9Zcm4XgUbCDoJfVYXd69FGPteiaDxBVo68HzM3fbQ886CzeldtXjykUqg
gYJBw0QLmqZ44vDluNclZ1gxoDiuxSlv25/lRJXGPK4lzmugCMl7qAA3kjNgzY5T
yCNyYvLlvA8dBXR9SS7MSaONuLcZX3RqwW2bcAbCHNKeEdBErNkQQ2xJauxWuyQP
HlMXoqPt/LNY89kxvYRug0hjdyu1lT+Hjr2Zt1DOlrHYNgwOCRW29+35C4KFtSsz
tfouObpp9mEo8cJHD76oDZap3CEMRcTGdAgVmeKgQzZWQJ6xI09wXULi2KF+eS7v
BJ8JtL88F9JgQDZ/PGbuaPEd87Q1mmGSt2H19nja0fRSoBWmgcywN7ynVc7crFtV
Puam+BeWe2y+npa9F6YADO4FjavrCr3mZ+kqfyEsXRVC4Dh0xsmDh1WpGBy2VgAu
9RPOL3B+aSPWirFAPQQnccLDcVaZFQEU1pLZf857Mo1mh1yC3q/9DXemUUcrQqSl
+hJh1ObcmHatM/iPiJoZPI3RlPf2A/oNo8iiItGkCyCniY4Az4HI6h38VV5NmkCK
8DygOKK/OqUcJLU5VVU2Lpvm1GuDOo+gGPn3b8NoGre3zw/LamYhGs6sNoVdn4Zl
uKuIMKjiYhhx2QLEbwLjitk3bNTEX/rT1VsouAUGndkdWho1xOKYojAqIiIT1oi0
KzJyfS/HuIIS2m9QhWMgJPxhbPHZ3eGF2q3FTsypFq9/yRx7+RF/O5OsqQg8uG/K
SYztsFaML3mQ87sNdj5iPUJrXs+8BmO/lb7WAIOzdW6Xq5CYGiWtcOilzt6jA/VP
/6Jgvje2oZemgZlw9m50Z4ysWjAONOHclHrALrjJwEdTGpbPpjglUTxNcjfapWdO
mECiMfBFvsuxM/L01IlLRuu10gU+6PePXRQDaK0HacrT59UUHs09OQDZeCDfSKOG
Qm2HAUTqLNcQLTtm+MoGa6ywumJ2fo0Ju9zwdfepjJZdgy/26LnBp/gL6cKjscSs
Yd15tGgHTYE7Q2mbz/H/ubj4t3megl03X1r90kWY8mUtQ7Tw5IG1+1maFoVvUDal
pBiv4J6xcO63Ui8q4f2a3tURdj/MzRiNKxHVpQkXut2J40OOf5uGhQeKAmv7AJ6f
IBFQXdNJgKwd10v04doCPwWxml5QgmMbvPi2hjkb50pD6p3eI8D35CnAxI62TjgF
mxrSp8oDMjC0Z7cgQq974zejO+yWSvZawUqyvg7GM7PkZY7gfZa7RFiDQIjDKUnA
mq3QbqXa1Y+ArW06IBSkMKtj3sm8ebHfhZIPx9q4u3mRO70fsNSrQei7b+VJ/LMI
1l7sLNKjVsdEkFMysbUqQfkaW/wsKq2RXpuhHeb99BmV4XwnjKbc2OtThkbTpfdb
riyHnMOKs9Lad+kI4mVrezGfk5AFnDTxuQbLoNJ7tC6thPY1BscGXBCh+R12odtN
jCMNkKcUNZmbkVotSBly4zfixX85fBKe53/ee7j4OEyP8oMcYtceyASdUM0lNejL
Y17JjnzWiQJxa0b2TqM+etAwDCCHAg16cJepsk0syvG4NeFBDcaudzH9QUB8Msso
5qrpddzA2gU4v9VgTtSLtmk8WSP8BUy+TjytV3ifuRSCE55mXAEFr19G6mopuxkP
PoD+vYmigAiiK1UVWz/VgwMJFKnsCcg1MKUPEi+Bukd/+ne/FKHQxPf8oMxEATCp
qxer8RIsCRkY6EwbYwu685SSUx0qTsNVLz/FILBlDmGtsI1N6xy9AiIFaEDHw+8T
0NcZ6Z2+JyjepAtZEgeBVpPeoM/YGHKAXDwk7b6ZGotAo99zK9MHZ8cemnwIKm8H
z7lERDR/9gOMDZCcPkhnHpaSHprbPnjx4TFeUF+w+mgU4mY3dX0d983VqY+dmMPx
KoH5L8xtrlVvnCL8rl4BwWA3YY7O5GPmPtxnWLSK9Ey8Hs4NsqiLfl9H2K8bWmZm
682oUA23ObWox8ckttBQ8H2W6aGmOYyqEkZ0lmt78l10X2g9TdiVwp0VfXtaNOf0
YWtUQhWhFuWqq/jlinWDllxOmmb4WnU+TaiuRTDKWyX7tZhSn3yzmwdw8GbjwUip
AFJGmra/VpJ7rokscnmv6KZTsTW3Ue7JIqQ0MQ+QkLOX15CdCtssxmeUD/1TAPmn
NMX8l8el8kyb4O1bcjOb+koFAsB6B+fCSx8RAktz0ONDjRMhi6pVgycpIRgM5Pb8
gAAcYZjJGrIqD1SJANmo6Bt7+/3ltnSDx39k7lYvju45xPw0I0vnGeyhzMVfzi5Z
pfxazqBTx0eZ1L5igpYEKBv5CcEnmtrCNW5GTc9JKqxt+HLcByDhkTK1uwUrIzoF
RozrKUOied+hkUBSHAxcVt/OyzllLmAMB+k0oteurX+EU3JMS+FLu3sreXIzCgKg
CrdFm/3lrNr9ldDs6Rzq21AtDwUnD0YGJU7OSACya6ZkOmRdiH1G9Nia+lZ9oRyK
W9GfVGxEhZeXklLk3qWHGp/Gtjc8UaP9PUOHU5Agp9s1RJKcGd/1XGQkNF80739C
G+bgp3QVIZQSxsQuoUqxZoyX6K8pAQsbdpbB/8b6hjUfzu1qx8DoHPyAuNNTjxtO
/cAFukoR35Zd5EJ7FLgV8Qt4jQ3quSOVIuSn8ZbPEwvUwrn5yf6zKXDZ+aDzJ2Po
ml15OnMdsMFkAifhFuk7cWb4GithHPpu6Egz0OGBGenkjLxmE5YSUEigZEPdVHbL
VeV2xVaQDZLDkL1MyGn5vGz3FTc78MkD/PUTQhkVibl9deNedS5o5h+QAY1L9vpI
qugdasSNvrPpIlhQ1PpfGNParOgO2Sh1A7m8rB1mVVP86WIeZMnTyv92qkLeV/rw
rOiEJi8G//ZFXpQkDHxI8dU/jl9L8WHoi/7qKRBewkqLsC/3EIUWc9pXjJcYC9l/
ieDAlZoc2TXxicgAILbaUm3AdEeMrKcx/9Li8Z/9TZMz06sZTgdgOLy7PSiy9WFz
D9ffGqb85mgiGhYrxJU+1aZXdsua/xqX23fepp3N/9FWgqO5zdXC5itoLFEPgPub
r2XM3owfR5zjQ3iqDkarTc8KER7LSb5e6VXOH+pALn6ifyZXt3adDsj2KXSYyHFM
4VTCIb5WU12+9UUvwQENknGb6HyzQsWzjHy9hEn0jcM4K/P2hOC9AYtei4z3NrBp
PVa2TinBDRBKhSmKjomWZHk7BukaBbNZw81EMXr6hNEu4aduL/hnulWTjHtaj1+m
aYgTZZjvnRtkZLJJ35R+R6fps3jI19ti4WPuCWNI77SQHQ6J8PICs3KXHO+C0ipV
tA3AhLJNA4MLPtHRowZODsge4OXhFYECChILK2a+rtih6DOwHHpGN9iX8Y+GK5tg
eKefmmUeQXUVMlkTKOM13Fc03y8W3QmzRrjbdXbiEqdzECuDwLJDKhkPajFVzknZ
Qbr49eBkZ1GcUZhY8C/F20f4jGYrxVPspnzFPi6R5icw/Gm6mHQ4kCtjuOOa+n03
421wYDGBNc3NeiVp8HUNAYUf9B3QxPjb9NpmH2wWIkLfLOfMmBOiknMU6Bp53zRk
TuWzdvb8IKrqiiRiJJCUj2ZiK8l3klZKD1TFFUkRNWRIrGpgZWgiqoMGcR3SUkca
sRvAG67OR2+WcNA0b2iXiDLOhbBd6RSuD82B8TEsYUS+GsofnEwCn5jaTwsG98LN
l2+uYbdDcrLqK/hH2iwHHbt5hDEL/bDAwLqv1dIV07FcZDGCOaB2Q0npxs/hM3/0
tV5RlQ++ntSAwrYsr0mldDoJL3uiRedOfP0mzQwt9gRpu82t00WA8ecQojqpMQSI
EOlSiCBK2kcLWHwRF43y0e8ln7e8vqRLxkC1HYSX9RC9s3LNbdfA1GhXxpMuVW6u
SQ4Tdq1+Ug8pkI6SBeETaNWsc+UG+MPMnO6onDwLHOjrhFtzMPyCe7iKgH4Y3/kb
rA4wLsypdauE6UnqXv4lODc046w2DmwLa3vnlObJcq9ZESEyQtAjrZRgikzucV9u
ISeTpANQmkKBQer221mrII0eRiDwvWcVpMEQdGrOynnpDBF0UwgKHolf1KrbXQXM
UMnU+BKPwF76gaF9p8WU/ta04FtZ44pl1OUxO/42xEBGc0fPgIw8OrmntSNTlz7L
uYaeLRX2cHN4TLem73FXbgYuLh3lHptyWxJtX3qwBYA3Ra+OhaCIWO/pxuQxhKVS
W21RAiQwLrIxhbU8tlIEURWP9LZLXwryjf6TwxfZu1zN2WUdyb8DqpZ/yXMpvwG7
XnxDusO0c11Yw65eFJX8i1JmOMC80lgU3uktLMsfTquZD07K8hH8WivtRLbuAop6
DCj3grdp43L61i+g1qmN1ptmgvAVlxGVOhGOaRWSKUYhghT1qg5JiENLfKdIlpdg
CZScXAVACDjKH39sZBtbMcBZl3KOwODukGpxsL/Yq6ZUaClNa2mD02b49W6NutMK
Y6KT8854Sn6XPrqPmv1SlRNJ8zxQn2AkZCTQLCi2UFVDpa18Ir8tNMvXQy0SN3WG
uJIzo1naatM3da/aW2mcsyfnVWU5E5N32h6PQfXg9Geq7lROTN1gdjgTYDMzL0Ia
OO9vjCM7NJI8Ygp98/MIYN9ZPK6lBLrolMX7rs4dUjhf0x4EZUpATthbtZFPXZnx
+33MnaRmmcexxg19f44VCEtde7A2pGHaQLFC/1ThKM90MPOcsudpOmt0OyB8OJVj
mksXZ052X8tSInAfHgh966gpxEgiZzFWg9u3vIbQM/e6yXZZ9rxuJwukOv7euR52
gdw4/be2rhh3gT0htuR55XUeVvdnBO8/CwcleJSlxALeXcw4GyL16D5NFROa4bsf
DSKDgq1uG4SewZ2z/veKEF3N2cxOgX/93N32Etfvj6bQx1D8ft9RgFGNcXOOhOp8
UZkjMnuc3mVG3h4aH5a1XCR5zSmPQeDaKENTRTOuA2kSI5CJqaJZCX+DGEXaN3DI
ND+OyDw0WlRlr4tSNr0dM/RuRQxXQg3hFJz3jfC9aUiODE2rXC/DfbtZyJ/ZzwFX
MVXjFCVURxtVWbnp9JFBrq9xdvLR3LpTZ3fY7cBF0MsWeReUqdNAosdsCCRnqe++
VZ9ATn/1p3/5pPEwNtlxhde6r0k9Me5SE2J+LESir3IjF0tPSirl/gAnpmQb1zDI
cmXr62YBHwuopa13HuGR9jR8O5y/cFbJhvmUemrZwyHsbINceJ+SzO9tLwC8Y7AZ
Sd8owekebGB+HBBHvQJHMALG8leDPGSc+Ft0UEizAb/3RRxaXjMeeW/TVhEZf+Uu
ecmmWZWwg0JXyWWfyHobQZu/O62WKLV9bHHb8plDFRlU90x8ycRDh54ITZlw39Ei
l9tyifMfaFIuNnKbHL5i3yFptiUyJHoXLcbyFW6pdG2RoyXkbL8hZv7C8o3QeGq/
O/cyJQoW9vvnPMf1+vvdPrLjj2FhPJ2hHEFcbcXxk+iVsPRmV8FgZumzVLmyfg6N
AtcLPVD94wwTcyHXvrpI8fuJKyOqzV8Y7WazVY/2IJ3peakJEeGxHi9HLP0XbuvI
j9VruWOHsI++kD9vkIl5iuK0C+cDdFQRa6GY72IVXu7agpD87krFYLGnETbU9BNA
EByoVr16dhCRfoAVj2RoDVYgRpjCjNve+pMBE5aZX2eRrqXLnB/59abDCzQgcoNV
Z0PM7B1i63l/W/08mY26bjYBRcpuVatf8fxTqzG6mHu0TWhSw/ereYGKhFHNctvX
v5CAAH3xW3qhHKoMIPcO+GiP/eNjL9o1XLnHGKn2A2j2EJdMdd3/C5I4nKEwmI3S
9n/DAcjSetAwMhGVMw95VfCN6CiqC5b0nzVy9w80x2I0uvM1bMC5uIFunFNG48LV
d0gNQKqpFc3bBmClUNmTLY2tESy6xdn/ZO/p0Ddz/QjJkOTs1EWqC2bTXLJlF8b5
0/+Ph/q/Cat5twS6Avrer9ojknw6kNUP1TnilYXOD2ncZQe89nEODPWAL02UD1OI
DUMTNM3mO9tOKTQT6PjE8EUNCO+2B+9ik22dv03AUIu2nRswPJjktBRt8q4kxu8Q
1Xazqf31vicqB0qL7yC8A545/UdLWZyz9Sg2yTZoXEecRP1P1HlhmpI6Ct23G43+
3jy58RhYvy6uOuyGjYK7ItOfyB3Cws8DMjzbPqG4ZkvR6hGnCsmgxmeY5348SQEe
NM9qLbR7dyJeA1O3NaGg80auekEO05JaxyfWFnrNXsbyoFwqF0HM1L39HEmsnUeP
bQ0mmjxd+8bMmE4LjxIwoK94Zbsq77INgXUCyNRDZtH/6gMj7m1PC0njYKqht2nA
Igeh2yrWjUQnQ5855tUhJp5lLraW0MU5om0F2+jZ0ba8LNahzP4bw+pcV3vpyDCI
kgW3QSBPiBAp4TWSMN6yoRCgHP1DD51mQ7zi533Nd4H6hMHzPaxkE8dRIT14xcKh
URfGrgzoGqgvsusWKfkq/lDussr/5Unyph4uZiYazkf8R4w/yGm4JtGAgiy0+Iyg
DLT494Ei+z4S5Le1HzImHFGrTm4ZWrmEcJydJGhoQojfB+BghYv16CNgbQ8B+lnQ
Gi1xbUUAqknCK5W+lsKfPwmVLxOYslCGMTu4Iu1hZga8NH5ArCwyuAEgEla6PAXn
WGvHHKKVDYC8wtTWyiV1vl8SqPuMHCGYxAs1T7Y1RUGjAN4Xjy1iAJs2g4lS3XaB
YMXkDtMUY2B+aSado1/E14AHJFgsvWuWNiLQ84Dh0xtjCcKGO05zlkv7C2uxbAP7
enCWyVj4H/WizXNK97EF64832BYQlSVNVzh8hs12Ci59j/hjiM9eFwS2OztPOXAK
Af3YQTy88OyBNwgGl9NmZqAe/bG4mmVnTMR6cOXaUEuYkM9nP45iYGRXqAHd0SpD
nL0oxRZ8o4SNNubjCyvOzb0EwPvJKRI4g2egIsyA6GetHmHLusgTFQyO7LIvUt0K
LHINcMNQfxsVP/GRG7Z8yGeafioGOYcuaEhyob9IOcsfpmjEnpWV95HEUo1wGDgD
ibI1QiYiZ2VmQAngsz1g6dgnSRq8kQGAU7zLRRgR16n4kIhgkeLUz8jntnxOL+/S
jpTwjlHJle35RCWOyePCW3Yrh3gAndDVgeP6EpTj7byKJ5x/stW8gP67cCWkK+96
vx6AITiLNGS7EZ+iEU47uswgU4GU+8zRYQRDTk7ycCuoNC8nErTbTpt1ddFDoVUD
1d0qdb+p7kSyBeRZdUaYF2n14N+rfeutdczGv/MuQh5U4stsGATFJWR/s8w6nKrn
YVtQvOTIvlJ2/OZ3nZq2oEfSv2YKT3XtmhvbpFNWPFA1v9GSgJStdRwf/L5CIvmR
oBa+pH8FUrP7bS0W7IC+lhORn6lM/lmZY9tMWwBaU3LdgVW3DG13teS+Ni9+0Po8
Xmn27V+4QhggLf9W1uCQZoSEVGPhQE7H3VdyTJB6d0waFxh2bw4knsS+kSF+/sny
mUI/Vo3/SJ+gmYmqwqp5xHWxWkxJWizUiMNzSznwVShj0487D5AHMdVL6eWs0Bi6
1KEi5Lb36yRTJ0vgx84tivWN5w5GzlpGe/lHEL0pfeaFziuUNru86Kt1ZPa8sVms
dNWqSpS5BwbULX4KfTsZisJ7TvwEFpDpsgjyytNCaX1o8RtV8QK/vwK3IRJxV8Cp
rKnwsryT595wYpmIRyCy4uRd078tmUKxj0IRGrEGPheDlHx5vNqLXPSljucWxBZ9
d3uZlSi6NUSPUZosP5kTRrXMC4gEEN7sq56mHXJ2MvY4UOBDHuqCQ9ZCm6IauFwu
3aSHY70OS1F05X0THQWLpaJqAlbs6vYmZxuT8kUrQ0A20ITePQXV0vEsent8JBkZ
tVJFQut/lTyRPGEPVKFHAtUnQiJhxEMAALdp+JZ8rpNi8TK95Ee+8uZW/ruoaub0
IPuyg0NphAf+FrL0TznjL1wjBBHv6AkeEJtpk72eEYUMUqswPw8CR6KvHccUsdSC
kQJNUtliepJW0LwwtDsSHYao+YWMjlEyWScUX9jLbCFps/Wv9Zl+rU7kz29AGMaq
DQnHervM0MofKdtEwjYo4T/LqF4yRF60Uolxhr5BNH9q+hNA+Dx5LUt0Gol2ZNZT
UEmJK5wjZXALkou94ARhiVn0uUZJnF61k/217rIm7omcOehBhL14VtmEpY7oSzlA
cR2agbVb8/bGJJ0kP4bvdZk1BivNsljHBAkJCyFJTD6kN/IErOB2J3L0ZTmk7wEC
tPCXQ1vCbufE97OieVvuEH39I8qktIj6RiBHKGVYo33PNPst3vuM7nriLvS1d70z
rZHSIKXnKQqGGS7wbfejtVjxUlfws862q3BsHRzhuWiEVHW5L1rIRoVl0S+q2UyZ
CMtQ33QilyMMpUMQtVzPRBl1WsRURH/OaBsHHplLdI8JyTLcfYStQ4bVyNSaLOQi
aKWscIg93Zpz85XXvGmpBmd2lKd00iDsHx0VP6nU7wg8oHoF0A6woNp+nSiRDYMu
1HdGt22Yu0q3QQEwLheQ4yG5Jwynvjh59/uGFJ+pmVVuZc3eUQYZCbUdNvXcLFoi
PwAWHtcqyB+DunvtFcsmcPGnE4TncwOTkmXRUWgHtj841KLBiX9Am8nHtsgCOMky
ZcHUcaeUCExHMhMbcIt2I0gCzdFvMjE3TVmO4y5nLmShgmatTjIrXBjutpkePocd
RISP1c+oXY/HUU28U1qxXW3HxWZg5eNlz76EOUTeChGJNB06ljOKoPppaR5xtpgc
rhIfKEuHy02gJMHr4aEJnJNKqcuu/sZZ7I22x/N7ab8rORqPhj2f4aM374EVreiC
O8nHuAlkAx+/IEKxyv9ncg7/DQPTVCekYtyRZxrWzTzJw6xQLaoZXTmQrV12KtE8
bqqxprY8b2aLSJlsZlbC4PvtNTuzlHH7lGLZRlR0w3cPImCPh7v/jvGx8rRGu7T3
D63qllcq791KcK5Uz8d3RlY9S7UyavQqlhifKJ6akhxZFS2Zj336iapSzkGGy0uH
4bwcsH6JHln8w+oRX3I07g38b6g4luy8HyJTQL8V6oOTUI+ua+16+1fzJRSNX4Wy
lVPgX4i8PPDLHZpJGmbyID3MGc7XSwTCOL/tm+5Wi14+3prsUChfOaDxDImcdiHI
3tJ9/0Uj4WuCtL3YQhHsvPsReeS5JmoLd095hNUAvFkIL2VRZH7ElNv/xSb/Lab9
YB//OIVbjgDwaCIhoWf3R8nxFQ63j98c0wkxdMD25a+SKpo2e/f5zcJ5OAnPkbUN
Z2a832bWduzAOSFjYY+pREj3nItrW2uEy4GGUhGEawz21Dg6PAtkBv7u/kVlFRk5
+00f9JLlZ+Z3Ye8wpTnN0z5SYRPRyp5bdiboii6FMTKN/9dNTqlTh6qs+PtAk8+b
u5S4RoY10QazOauazgUqcoie3gqfBkf8GfyE4kIogAwpooBAfM9AdW9RdFD7ZJrV
OYrOC/X84MnAZ7sZQA/B8FU5LDw0G8jnSCVztZm4fXpGucsoaUmCTXoR09gNMdow
nCHb2Bs9CptsE+BnWG/dKpbpagTqrIhqT4BtmWshdanQPz0TIWg5Z7PFVlXpegKr
F+EENX2+Ri2e4bdM28V/+ylgCNMSvFMfBoskrbKcvBd7xfp/pZPwYR66XkLw/BEO
yf/sCsqCZjtEAqELAYpE8UVF5pdjoy1cLpXzbIMeIPq4HP4Jw9kUvaPKMMKFQGw4
DPuBvHmv2zh4SOuVnY0VaJ/PRgM/t371UyulFusaqUODSHaGzQ3dr6jl2iRFw0jz
FK47tNmvXpe/lYu0GbrFmkVHmI9Scpbual5gCzG0SHYO/8tZQ60BRQaIghDBPiLE
JtjJP7z3ouu5lUDJu9QdJLCpsZ7/ErwX8u2Db+eMHrbCan/kr7XSg7pZSw9MURrI
q6EMT7st5Nfg3bD528wo8kVIPaHuT9OmODEDuh2iSSqehQRYlq6xoYt5EO62yZH0
TZxVGeTemh5hlB0ZOq7kCaNhWJxTBonourIVCPsfGZ/7lY4rHC4FAYI77Lj7OR1x
ydSY1gzpNRw0SLHT53ufbdYBpRIRM5sg9PiUTVgug4jYmLcNR2IPUmk/BSPYolCi
86Or+7U/VTAIUiR2eKKSUySzwAuf6AJPSpjmJAAZGnmGVKAMsS4ZVQxN0XSMCSLG
H2VuKeOKrIaIX01CD5qgNf5LzYAE6Dh9v6xzc5rUZAZmQsEwrcAQiZBevOzJKsj8
X2z3Exb19eX661Z5Vs885OTy92blLZfMDxkK5nOCataFN0vcYEh5gwabM2VhjuT3
cemiB8khMXuwCmugQPCEP7Cmmv8QXmvzAGcwEGzyudY0yHPmyjNXqp6sqjfo6TQJ
PdUiLHrFGByRP2f20TpXWs9pmhStQYPnJzK8ZMbUXzn0nLV6dOhI1p0H4r8l0AWQ
qsgrZvRjgHsi4hDHe8fybJvmJxMhJEA44q+/yQcPp6LdhMl+aQyqMfAtVvVArPEO
qptyaUrxrUMH7tNQNGEtvf09SY/xwbrkfb+iDdqMjCDjSykfMeBzMxDNGlnPoBbK
by7JZMil7yDR/TiUd1CTJMvhmZObiWyoQa50WHXyk2H25RVVCpsRQXgkykvBtawc
BJO0wwn6Gxk6CRBHaX/uaJ5HbNw7LFIUcSf6hHKOG0FPfzgGmJLX2jGzdQpzeSia
OKvSuwAg+1EWzRyUOlThnwSqLWj85VAGRhHe4DT6D4ETJtXiL94XpGezkPoR95q8
0usetp0hMukG5Llqy2IbzT3JarODGs2J5A2Im/ilOO/YF7zyHp9XvVvOxFpvYGXK
6pkWCE+1U2L7Wu2pLG52Fhv405j9TuoIsXyFgzS1BtAhktt/8NGYu4ue1k4Db74Z
7wB9U4Tzq+xM82udh9UZBWc7MAQJMsGqsW+5Tm19ER88eUgFbwcdGeDQ5gGUcDaR
qr5EP0+I/hAsF0WmjlnxuzEY0T7FfYYZXUSGw22Ci6Y/3DyNqOcawiAqVacyDKbT
Ex9gVXfy/5EsLWFsAtHhONNRtFcxKVsHOsB2vZwzpqeU0NDOgbVxTT9LqQE4S69F
NrwoqBgAAOpR/+WeDpoETGQlH644VYxwxvF2FVjIRPsSQ1n8QZGKTtQgETOrrco8
m2skLmFv/VYVtDW9LKFbOn2rVkwaY2mUIN0LuBbM7suW/ZjFwAReHcSp+K5Wwq1R
K3Lx/nNlr/Rt55TQGHm1eYVj4POBuJmpyMWV9oszjb7LfiD9xO8yFJY9JhorYMQg
ainQs/fR7i5bHlVqggP75RsoW4sXQVS4rQNM2bkU57T1X8T9IkObnXdjNBXwe/2t
zoVEMiRna7H3LTru0vXiURVRR1I7wbFEklAutdyfnbMupkOvGcdAFyQwHgWTJMUZ
x1KpougG8SqJOaJ12dTf7QxF2oawPFuYcxZtt8AesClpv+NWfN44QcXQx8yuyR5F
KbcT+x1vUQG2hik6gTP09+0HzZP7/ZREIuUxmC+fwfIlVVm3ZxSqTI/gcEpREdwO
nVde6BHDEyeQDIg1cEuRrP7Ff1pk4ywppJwkxgKM30N5drey448ByZiAOwuBB+X3
8VKsjS0NbfzQ5MLLZWq2WYvr075GsuV7/2TJeWQtjp3+SXptCFNbxa4s+ojz5MwG
hY/1THRU7LvFTC8GBvPOfbieJJ8LFMNe6TNtHTkcJXyHNvAaKq0WuEp1b8SdewwE
+rjqcY9n734aTCd8n900GxOYX3vvbClma2gURX3TR64WdmWxR+cTST+VqhA8mJdH
zSB73u7BJbdR6vSJAmpkGGMkJvRyOcImeU+nKgrCbD2Fs1xI0gkfypbxwZgyyVQX
SsXG6re7dBffdkID9l6Eomx4hT95KJeVbnvaua7H7zMPiIASCDvo605/KJL9gAiJ
0yrH8gNEpCUmqshk2+11M9mV3eMVN1FllROyHpIyP7W86m2cOC5OKuERXdJ76WUv
kktY9golJMyG++dkowzMXD+s4C8jg229L6bojYYn9TmvhxQuLkkUgP9lPhEF3uDT
GJRFR89Z4n6zMrCy3ZOVHnmd5oqJ4v3kxxYHqFTONVT7gva5UAEdM7PbVz6OlT5E
gdQETo9a4+oPUqzRRgjXxyUtIwrtu1LjyGCS5FdTDXIg5q/g3otkor1mZW8AwP2R
wK1tlr0EqnI7wZG5KA4qh+wLd6kjZD7iBJ86VZDsoOzX1hr9/gEXQKXvsV8PcKkS
kfMWE78MMSsBTQkClefo3Ez272+ALQnXwwgj2q/OMy3SE5OKN1PUApLNVDPty5cF
E3pKngTpXBrleC3GOYbl9vR9uRcg6RAmHXS8s509th++4JwpuW8beeXOH/ViM2he
YoSWlqnLTuGC/110nNScjnA9FbSyNIyNQbl/JSTWVL1tpsDyazOHKtjyCfK4402M
Bdc6OFM670anGYoAyyTdsaKXs5rMQ/wY9xkyGyO2wLjuu9Z0f60BOELvSBYV9DMS
ediGK/kVKMz103fImJ3Xhn/mRDPbvJcYH7zo/bo6oDfCnSUUqJbxWdexO67pe92z
lR6PnfeH1svF4NHErvx2Jd5UklWmwJRKbpyKTsLu5x1dzfei1xdVJHwnl5T79Cr3
4lGP3YC/nlU1cQU1zAm3f5k+QRUb1OHX2ylBwrsCe1a+BIg7Gtw0rCcgJX4NXAQ9
Lu0VvtQHvzm9Xe6/Ph0rbIy59Nid9shrSB2i/bpGnnZxc1hExb94vYBI5+uoufwf
99TmQOIVziisMuaQ60ZanvlPGxESGFb6T+EyDFZNCDs6P9DETJ0RmLMZTbSF1R3z
8p+oRao2F6ldehJNNyfD2DBkqPjzP3WxCcVuUFa2RJiIdLAbtMGLbljS2FdnzcJ4
NJN6SbwEUHvpy85JxI3Et8GeeccsqRyy9JI3qWSKkF1OC7fVCkEDxHrqZEAwUi7o
Zhb4euwLBN0hojDadcuMVcvkIKJqU7KjTkxlqoihEQAdsBjpplRPR8nJOREItGZE
sXIRD46UeCM9fXSK1RnznSTp76YdNq4fDtPhygUnqExvwk8Qci0B9r7623ywIE6H
+puL0JVgcaRVRvIbcnVx2dqECvrrb32KfQys3XoPEI/+5UQniA35X/Nr+9mvk2V+
3PYnHxvMHOZlNe+/A+t8A4J1iBRThqVluBDAYAWqurfZP1kh9wa25iu3HgU2SbhA
RtPPi4V9c4uN+z1xaqXmJHPxx+rj/BPbwe1/3D4H49aReaaXmgW/9VWwGTi5q664
HDO3Lk7WfmXxGOkFAqFm+SNKH5UXxhDhh/gxj7EUXi9R4bho0ohnmDtih9RBkTpW
4Zjyg9qHOI2YsFb063PwHS5l855Wypbuk/1Qz1PYetnquKZHAXCNIliQvsOUIGzg
eWr1ppKwNPQh7VAsQnM3/TdVupLVbwT3OM7RFcpjmAZSt7LNvagDF8mv3Y0Kojo6
crzm1evobTpdKaqodw/sbY6FhICe/5vwEWiFY5XeIQZej1p+sRYGa6jPCWF+x7oq
gTX9aA+sHLPSBgCtehAkHrRO38m2i/0DBnwnOQWNzupnbWObxNvZ3vrEbgXYxEpZ
hs17vhmROnPYxjI2wWgbAOV2Y2HM7v3hrjcY2xyQel6TgM8REj2s6jTFiT7bnv5u
c6ucIiVSqO9Pmi3UwuEbtfOf7mcf1AqngqimCx19NqVFSiXR8k1JAUQgTvIlo2Pn
pjqqonqOmom9Yt7mvMXtXospzOXjFf9AVKY91UK/wOhTavl23mfjgFm+AE0UEIhS
COBVIfuKq39l/EqZNoMDn8vI2+07wNLGeu+O+rz4mmiTwK2AZYYpreD4xe7bVp3l
rQc7L48NSObgHyVm4yUQ4nRki9eC8o2WKoRDr12Rq06EiSy6jc9F/KdQs36RQO3V
n6b2UDb/6JfV0Rjrf88ZV1lUQR1jxQIsKHhvVlS/IezCA2+JeYoaDoLQMn+LAo5N
KUtzSuPsQMtbEXIfagnyijHmCRr0ugECrdX2LOvnCqJGI1L2lOeLulshuuQHciw2
50JLfOyoGd9bK0YDZ2SjrqThhGfg2s31k/bi2IYa2vI3PZroKDwlpryua7E9RcRR
tvZtrcLv11jP+X+4KuWWl+04gNrr1pNDUh+wXVSP+mgKkisRwlFhaO7q6yHwOl9E
fT/Wr0XhwntjaPNSZGTgXNTZ/up+vIZfD5qIkZ5FU1oSHS+bIUwiRsompcAJMlyg
Aaz7po/iftYT/fKyAlSqgen1eGP9plfKM+dbM1TurP3c57DO7D2DxW9rNdZ34EKV
pdcYnZlIGRwmrbAiGsuiVP8HBqnc6ildlhdDVMQl1Orpq2uNo+S064eel3y53bKU
ofFozTxMvTEqJNib8QmTMPkur7jmDnQ5vNRfKjiqgnlSjs/OyKHndmttkWs0/Ji5
F4bZVaiRRVEtDkN7xTameMCm5cY/aNfuAlpzNd0vRJERSjA0jw22aRdOHOZVXhNl
uOLDOqhfiOuM35BRkSDnGidHMEPusfN4Up4Aq6ohLgXdoN3RQM7eeP0u9LClFR7L
4PasvQa69A8uZm8zn2whLo0S71VUT7tjObLxMcCD9odoGz3kOpPM82QC6hDPiX8h
eG9Z6yhOnhzoSkSWpKchYQXbRAY3t9c7JhKrhPFa6jBlPowVgrEd4NekPevKlmoq
fy0UzR3ttXcbwui8bYA3j7l2ML09+/5V0FjClJrJ1ePCffxVL2Smj3hsTd/OtJVo
CRa0nbKS3s4d/y9PsPWKEbL8SOoRcN8aoR5u6fLPbeo7MY0KnZGxVB+pejf/lyNB
XOl6Z7A2rfYvJIHdWQYyBDOOe9GHz2G8EJEL1QOtPELZw9n/YpSsEqamXliBkoCj
HdzPykPnBViJ1ah7Ph631ek7gQQ7btWNZ0ZhvvbXm90eIvS7sa1Dd6LmaONjJAak
lR9T6vtOEDVeMDLhp5mxJ3VYYezNZ6tG9sVxDDe0MXG+m1LE8+wFdi3JGdpKe9nD
6fOrxdAPYzJdiAdOU6E2dPP894w7injfrsVLl30yTWYysgZWBJydKKXAMAgTrN9V
390xQP/o4+dyr0WFv04c1Lxe8XA5cBCHn5phQSwOhMevw+0Umgx4Zo5Ez8SXEF1T
TbX8bdIKqYHG3Se1jBUW3unT1FJcAEd6Obv7D/fpYQixEJ0X41pjA0VkFDOxjqHg
b8pP+t96YxY+QDFWEyDzmflzBxlGbdd9FSBW0TF2RttNS+bS7A9P8satvxpb9Vwt
H3mjBLLsj/ZJEhWX5Y5bbE6WGcbGHDeJLjx1P34VKq9uPYXw+Gc4PErEzIHHzuFu
6hHYrXEJ78hG1KQyS40N49/zIX/7QoXKvBHfR960xesW9xvMe2omMameTedwyePt
RXL6Mf4MgJGy7BlbuBVvVSb9l0qf1eldGaRbxu1RTHIhCjC2zJv5ZWdRt5ip7n/K
j/FRv+rbrWMGqlFVfpsAcaYbdq5xZgGdZzXf8rVqL4NdLHlCk6M9h+9HUsD39Eop
6vsv7SKTRcBVyIzcZJy5pOotDRfKO3B9tV6SEaim6mYoNLFqtW+O14pOkWr0t9pf
tnX37rtjKk46dU0Lj9mYzrdlQpJFooPK9ecXkVb1RgwUdCMOfQzgX9WRkWsRZBwG
ZOVpAUDGSWf+M7B7LXknVevBr/Olr0xcreuZmnlQeHu8a+fIrJggntBFM6g/M2nC
zW0msncMIY++Si/CCkOAWxGh6WaCQEYulih+GTAbrqBsSjGch0HlJbLZo3ku93q/
M3a6GeW1NIWpW+GDRQbdIXdvnqrQS5mNlU1R58nGdRA/cwC7V5lkGGd5+jnUK6KK
Ijk4To6lYZb7zCoEitUCJAX3PRC3r4sWCOM7AbxWKxGXsJ4FFEQxiGIpSMauTkZC
daQY9X4Vgey8fjFnBve0lNlza85ePu87XQaTK2UoNtE7Bc0I+FdL9MZPCIBQn7uJ
Ihyma6B84x7sJDX6GQ01PUn55coRthDFNKoyqw7J8SJyEpx/Jbya7mEWPGN/viup
ZvP8nEUhH8o1c7Ni1dGn6X1n8gRNj33Cqn4qlwYyXV6Myp8dmAVEmPANmJGkrj3T
/2UJwq5UIKu1njH6+f7D3Pmr6Sn5nzKEq4TBfW1fBhBOHEqlZiseg9KFVEdCN4TJ
h/k2doUh527UANHVOGGS8Z/hpwd4rXMI/frfAHLsEcCbaPEQPLcbaTP9g9DsDejz
9hgGYV7ZEBvS/PuvskeAyPM1f8RASZkSk/lQdSXX0U8ua3ldTZ6rnTeP9FewAEAq
HNxji8tT/1LUnn30f+XwSqlJNMOAR5xpNwJwty84JBq86GkJdl++R6KdoXXIycop
gtuaD2tu+3sSGoyGkmbooFDroo1Gp9bC71MhM3LlJU8beft/vpS2rmOopMd8grh/
FGubJTEoQUqkiHcFvdOfIUM8d3pn4m5IkOJZDmOhHeyZ0bHOpQo8XWhN4GhYjtEQ
iOxYUV9h9GNhBdNmJnWfAaRIggJZn9fQzwjjeQp8bVqKQmbU0DPeIg4p/Q9YAIf/
jdGqYkT+WJb8i56KdmSGhcetouznwMTGTxg4+chXm7Ie3xWHM9FxeIwwMFGfDdDz
63AzJ25/zqu/7abZIQ1Et2bgp+Owxa+HqKmq0T8zPtSxVtAzjQxsAXC3E/YXc/jj
UoErWi89sUX/XA0h5gugHmyJStGdnH0x0/8ZThA1Rs7uQp0XhiX/C6swPfQqd30P
eWVHhM8N6Y0J5ZMroabwyjNHr+9fw8ibEugh3AnQlZpbT3dg2eMsP90Km0Yo+kKI
6JCTFm4y6gcPSR5nSMqExMlSO+2pPZj1kP348gNNq3m/vGaKT5fWoIMT7SemjuZY
yU5nZTRU/0z9kThis1McSz4ah7QugvCfMS7MbwiDcR0YFvN9LM1ZI14Nrk33oftL
5GDW89X3/ix8cfXz6MEwGpObez5cxhsb5PoDUnipdFc3q6O8gD1xbFCiKGgt7fkB
74Sma/L2z76u1wjXyQtx43ULVUKWA7QqWMAVBwcsgGL1vPMFganHPZOL8/R1wdFA
Vki0xojSbx3eVgnvBN860siszH7wcARlYJlzO4T2Lu6EOPv/ruFnysRVU60EG7xy
Fj+KFnEbCH4FL1g7MMQS5yIESgbUZffYczTDp9fdibp3hlLBXVx2lpLanSWmxS1I
ILRcDE5JDoYOTEt3AZSp6FJe1C0NKW5QflIC+nKkgLbGfmPHKInjqidX9kuJkIMC
VGOyKoUrwg2prWAHfX4ESaH2uM5Xz5Uhv09eVmDvlX8zmQ+aDjomAAzjRCgd8NiS
Gl+Zpwgq75gGKaooIHjtME6+X5fSN29nE75bVrmCeyZb8T6kvm91DuVgNeNRYLqT
URsenWkWL3drHClO4nRglPt7DTn/hnbIFGhkEneqg0fCuMN0Hb0roUM6dQDGoE5H
vG7kbmcpIZ5FUJE3JM+p4hSquR8i02M7bq41QYE2u7gvhduhaFcM8wwkLdTWFa7X
7tkBL8XxSRlt5GqheyVuYjZd6cXke8ikPLs9WLnV3u1+UAoHvFbgHt5c1vbyYjVZ
aH+VBphGX5L2sLA7TjRk2M9oX/QbV+SrLvctFstxVT3j+2mPFrDfCAC6fa5FHS9A
50JxhexkYf/kiI61Vpc0Nn395iokoEPS/bmRKNY9AoO6DZXCjm1+SLexdeHlNjlg
YM0se7/mk0rh6CdugrPUmXpetUbAEIw1EKyNaBX+3ux5pR5MAmMnVmzIFkhnSC8s
QVcZUhqfeMMHFrx16ArhTJvwcAss9BRaCelYw1s1DutpRkVN5EcDTNjn+PuuUEle
n84m4rlOfXUX+QHnzTN0juYs0km06d5etbSsvw0IK3F7eWD2Sspm0hO6BPP/Dwdf
qpA1OZ0tUSl12JNC+VXzqDfFxTiWq9Ee5xDg9WWQ1L9ls7qlPzi+kRWDRQQf/z1J
ULuJ8xwawXZ01zCYrcCgCp0CZXx0+/P0bG+1I5z7+NB0AKkh+XPa8NUrZg3tBj9a
+AmeSvQ03jNO1BzTGVuLfdoQkk+ta/nspQ+1YyZFaSXBqxS28nZkbm0XE1ntfWXN
LY+T9+hwmmHrXDdz8RgtzDxdCzNADs8OCpJE/vYz54Rrf6QarlU5Xxib2iDnjJEL
OAFqI4ao4n79hoiLsWyfeUIbC7PcrKS0N9KF6pkUaq3CZ9oT9v9oD64FrKD8uZNW
FgsUcG2JWa/daBCfOSnGzZBXaXeQWXcUjOb2fYDh/+FjE4yo1FONYsSxiph3n0Ux
vr3F2XU8pIF3Y8wc7GO4Bn9z7AUPoKXC4aZucQRwF9RDlnIPAtuyNDw+fmWi6ztx
mfkxQfzBP/B3c2yYG2y9HlOHYrDjj+qrx1SkqjWnDVwxkURa8tn8d3d5tJoXeEI6
lWQnrNvacG3BebMVKjnTyzacjrF7f1t8Ym7Yf3sLYunOWzT2ucaddVTVnSQe4bWo
5OObL5wCdDoB20/DzdhVM61766GeUn86wz3n8+omD/O8c9coXnghuY+LaJG7AQkb
a2bxv5AbVBwVsRUxQIwMT+RZ6SdsItB+F+qZj3dbVhqBmCwAQcPp2ukRyiwrXFqT
1qOLWU1a28djhzG08JrVhkWOYa4OBLjs6D1xw5c1N3uHA1dnVusQaUPOkiz0ZumU
nnN+zRbuPxKMPIvuH8uEbUPjI2T3373L2vM1dgBco9z8MPggWmT5XUkBLup5iKc+
aDjnpmNRoyUsur8CN4Z9Eq7j8hScVmORnPAF5Vn3tZsTUzz7oL7iGhLEf9CkLfPi
5QYEvjLIJgZvciG3KLuRxJsSDwi1MKoEs8sBOgUe8uJhX/TRPoFisqP9+DCZK7Ro
iy6mQe0C67au2tpIlk1V+4bmQv6UbhF5GhopzAuRRrKvcq38TTmdGQnudR2E5W0v
JrtQ94MQX3SzZmzon9Rmyi/jfJpB39lJ9FffLHBYTmzSHpQBMQEVR9iL5bf2b/r/
WtGHOE3hRt/2ItJS/TwqnDBDZFMUzJbG1O/YU/0ZizHdBDwfXU8V5rLf8ASwBSoH
Y7N3PF4vYE8sZuLPr7xLGwQPWpGE7UBzpzktzRsTSiNHyLHsglKqgJzpcgA7Kbuc
2mq7FPcRF7BUJVz/cGyK552B/MAwwdKIxAw+j7o7wGZg+tyjerm7ynzuuZEy2uNo
6tEHq/e7IXQ0H3ZlfkgJ8gH03pyk1jm81qXJRY0seH67cmaKWAz/m/yNzmA61lUN
y4I2qsq743e8ELkYa71YOiSOrL86eV55V0MA0fxyOG5jJx/eq8q/s5Gt1rrCxQ2X
BKEJRNhgHPU+Px13DU2uDAgCl98LXCGkQq9iItz+YvH57v2WfLYy0PKOz+L2MV6J
zVykzG3tYs0gPDSRF/oWh3MX/DEeZmEmbThg+O4ilz+hMIszLDArgvxtwlWDbU1Y
veM6iOtuuwtKUSbkTZ+Rw8XnqA3ew11xzAzNlMZ5big1Wb/zDh201QQK9K22QOgl
ViKZu9YP+1dagyEdOhq5h93oNqgA8UsVYeH8Ko0iyETeY4KPyTObvVSf+3oDy4gB
4Ogn5aWA1aeFnl8Z7egX8+/UjyqwKNPyB8LU4YIJPfbY8BqePOgqvuwI1C5VyI/4
xQS38gTFdbHkZYoDRvgCkfYBoII3Bz50Fz0Fc7G56SIYtCsbApvnkNnD5U+7YvTw
ybCvuEjlGeepPIK7AavXAOo3K/qVrx7phM3UeYScsE+pkMIrN1tXypMMcliA7Vgq
k0Ngp7F1iUuqnEqIplwvKWmG+4pzCSeg3WgfDPEHQ9lLlwkGiK9/KzVfpGjhpgwv
PhGsgyW05m6BfENlNrnUMVdrFkliqd5/ph3w4ka3eJbvZJdlB3tvLW8PBZod0xjK
6TUwwmEnnqUnx/K6u8XXSS4ERJIsJuIUz+1S+sfv0aGpTH1pcbJnhl/6BhC/vwD3
z4bxLmNDWZZl4AYRjtk99zpXmwj0XfDOBQAE8qXUiqcjRyrvtXnjTmzQAtOQnmXk
puQyjtuLSrKMR0qL1AjSYm+grpwrEGEIHMLDkXsjRJ142pgw7NdKIhOhKGNH715X
d61vjbquSBViibOC5BW1pWNwizSG173Uox4mpZ4kNDEuLg11oXKmbG/HkT43m0Pp
Blg2msJqeVFYfsS8bZMcrItSJXwozr0PuStn2D36blcsHDrMLWkYKXPc8Wg91ztM
rkjG6KEAlVEQb5xBvfdTj5TbjC+OgrmGUVUe4ChhVb34Oe6o2T402Fh3ueZrJnLC
qxvsklVj6h4ayJc+JhFY/HcX18diaJixF6dAfq/kmjHg6ofiGtF3A8/GPKxjb7/x
pmqg5/O1URkECBxcdrQs1EVGPCYCgYwwY2o3Go371AclzfcdiKJ5gPWeO/sqytw3
866j9kpSkTYjRY5WTel6Bo+gNRL5lezyLmyfIhdhgP8iH74ghNSCpEj/owLnTR+7
vaAshlVk0pyZ3HPTprFF4MdI4/HPIUHudXdCTbkhu1mk5rqz9m5ySjDmxNIaeTkw
edxV3CHMZLezW06T9DuwELtkUJHG6JGkrkIhZSiMViwFKpU26C1/W/gyHwYaLC7H
+kLxOoXxfJsANZMzLZ4Hv857wWU5YviSnvMlP/f161o2f4/1GEF+YnbCe88wMvJD
giIGH+frQjZxS2WHhYtS7ZGJQK8XbdMqvRkyE8Ai+cTvGt34OBfEsCPN/g0aW5C0
f8OrzJa8LEidGllrkG0hPt2oljJsRvqIZrHRxxDtDTtfpcNuIQ54gTIH+tc/4Ynk
ljaS1qlpU23a+6xDwdJp22ayh8KNLh4SjHmV/gUsho1jhTrM43Izcm7Refi1dfWN
mp7h6wpRmPmJ+YeIKKPNjl10T8SlCQ5pLRQjl1FBXCQoDAW4LtcelYEA+GfJyoJX
s4oh/8UyT/OMSMNFksq1q89YzL2XMyttLdEpocszBZYXtA09qSyDEQoI5WwTggPf
7vrx2CLwuuN+fXm55Jf/YHy3clsdr776uGoDwSjlDQdKQI8z4kH1Palbqv+16znC
3i6cHtBcM/dIyLv7qyavHekm2EKY0sre1Vm+LLOjcxWi8yZNiOIO6q6Sf7m9MtBU
JW6XFiM98l/EevuOCDST7/Zmk44ahrngdTW+xgRc0EgPaAWxdcu7sO5G97rC0YU3
DQBRCGY4+hw7dC5jDrPcxQ6cOr/J7A8BfR+Z2ocYhnz0u83F+sm6BYSmG/JErJDj
fOTfNi2It4z34vjY3DZkyu8+vDt3EbLKeRyXDnYc+jdhGlxKML+ObQ1mDNLwn2J+
iAXBphDUnUbYIYRhaQuYjvyfuMbRh3WYATwuC10PKXu7fBhomBI4v+HpVatc27GF
k6z8cXaPXPOKB/Nmqwe85yBZ8GMQUy4PEzIU2ySHTJq8LofQXjz91ABkBS5O1yEN
pxoMSR6zUYb5koI1Tzuh9TIrmsPocBsTI+Rd0ExNi+nUZL56D1+RNBkYQjv7zS0M
360gACSwlzygpHvfxiDD9jPOKFvQrA+aEY3wVWEyXpNSZ7vR9YKQkFUNm6veH2Bb
iEEef66A/rPDtu8mS9fUDZcjm+zPOto7pOrc5W5yM42j52VXgselpgocRRQ4iLE/
1cCKYMsL28rKCg96BzR7QCjZfPZ+OKTGfX5E2RNVFmBVcroUVpgDPhc2ctLX00qO
YRDzKLyfIHS96FP/uZYqCA1+B/BJwb1zEOJNJcnD89dN8nomOVCd8Lfk0hT+bU2c
6ZmEH+YturhW2SjtZeB2vgXWHnxhA2f/1c6Hm5EyHY1ZFtCcFrERHjRbHu9c4MTL
k3oei7aYbI4+A3y1mT8DbODfq0+rbgQSa7e4CipewIy/nwgE0QldOEOuTOJXuXIv
mLSYIIRTSaHatPZRHKJgANLizm85sYqPdkJ60Z9jiOenMx0+k1PrRD7R2fLVwDRy
p8yycgqM93nqVj4qKcH/kvLOj4Ieu9Xm3Y8GsUfaqXbix7lo+F5gzjPJlKotHlu9
ewpZBaf1KlYqK4YCkn5kLxBnZA9tJA56BsSoiMfVpeZfevq+GByhNGb0KanTIBVr
f5o5mSmLVu4OoVBfSrvp58JZ6cI2XSo46pY0IVbvU2HAZjIEh0a/Y1n++/PeLrcy
vfyYf34PbFB6S0H470nzm4+9LwCj9P2aOCpUOmRNZ9ZLCKyuKG6DM9JvdSnE2ws/
Y+6m440q5Z5fLZeo2TTwfB6W4bugdkr5AhmLwRlMTvLDpyU/zAumpsnsnDv/vsUD
mi+i/xbicGluumVtdMaa6IXc6euAaRelNbnnxK9iTkTOiiCvuUvMCkj4eqGa0/yZ
oh661du39xcHuI+5uGFVbifyXPSiaSGFcUOu0FHNGPsSAa7il32STygfkPI22EQk
qLJtq7+bdM3E5eHu2S4Zey9aYSdabLqIxt8dx3H3tlSZ6Go1jBCYd9e1aw8yX/nt
097TS2hMJaJAjl68nRhCYqcrVfg81wpzExjILvpYLiNBws+JPW9KT3jkD4P0txe3
PLNLuYmr10zeh1c2zKW2Lew6kXlT+jnCU7KYtOOzMH7Xa7R+Ep4BcOortqjykeQh
6lagqTjZPUJE2Gx9rTDKXYuDd0dmgRKw5Nd+SveewIJf6IeYUpm2Pz36FWbX70iT
NbqcTRZYQ9P5Zq7oSdcxeYEu6vUaJPtdpbFZOMHgL80yRpW1PI03nW/DKmU8mr5K
EdBBP7AI7A2MFbYB7M5dsqvgv6xY46VWN7LIKlcuhw81IFCUYkk7YXuj/55Eql0a
ut2NINjtXxHtB2YW/X209rjkrM+mF8PZM33HY+FpLGWgMmpZHlzpLsa+D9YjUBbE
n/5P8YCKh+Al8RUZ+9mUy9MGuxtm2q7DWWfQ/KlZ45Lr9JR8bLybqwXx38EcbaFn
XDOC8jXFQsRDdXd8RInndmqa98TKPqtnZbR1HC45ApfiCtQlDweIjpIaU0NvY5Fq
u0W1vsxHRZqKPdIt3I5KtjqrfKKgerP3VRYwNsUeHuFEWYSwiVVM4RrCFVpsn6OR
Bvtvp5vvZhyitLsB1t+XwWVRBUW1Cn5o3jZSN7bqyjZXqM88IXyVMipaXXm14BuI
5VdY+g76rkkJOwq3m697PJQHyLclUm4a9atui13SlpayeNXTinzkEBNRfoFvjSTM
xqUAwcRESw/XS9d8TWux6opQ5uwsf4IPWfJMI3S0cthtHDz1qftA/9XEcZ3XpQfo
q6i6OQf+6SGHYgXyJ2cG0hJVnM9uxgD9wCOjo6t0bGBHgnbBZFySDSgvqiNFiz00
EWsS7z1qFenX62vq68Uu1u1pHsZ3ccUHcQc30zqLnyGu63pxQ7lctKy3MV4jl0qZ
wJsu4YdbTMgKI/HTjpMAKj2rby11ijdeYFyi5p9hSjONWbrE4CiER5wsduUqxTgh
iAeQBBszLIrsseJe3RQHi/cueRRlnAK1BuD9i6OrSTTVEqkig7nnXC0wu26Dw249
qm9bnq6mI9697XhqAqfu7olahFIbUTuusTNkPPaMeNVsk1Ejuybt8drCa+X7DuAj
lGjCbhx78TC/mBY3N3/OeZd9CUFJ+Bc9ua4g6Ts5pAF9uCxQ1+JWckQ9SZ4mDTcu
yaQAjTi5LxahZLEeJpc5YjwrCOlq7UUtqtFlyqPtz/8oZRppiHsb1qiKAKMpRH+w
wUPs2F9b+i+ySVXehJRhNxYv2lHK/xBOcy79N3zR/YmhrrlSdFbrxDjZ0IomtTab
Dqm1diOtkJLRHWeNko+i7gV2rcgUvpWxddiAKjuwKUTSD4fQ0KUCRza+nol/GiOW
0CXUW4/h2028/SU/GIBiYeSjT63Sp5lKuhNZZhGroRiqJeGqC+mD20IHKe950Dq5
IF7ycQkYHncsm6fB4mJSri+Pg/y1OpYBYF29dg8xBu8tYlGTGqGXXYSO+9a7oA6+
QYbUmAOMNkUlTa9rj7R22ZWYWl1BG3tdekpvCtwMVcfTRflKgM5gQxGEG8fzgHXX
yhCkVFNAhQUCOdasqTc1x3EapC9x6Moel15fbu1xPT7YcU9y8PMkVFUCByT7/pi1
7lYbh5/qaX6yaXlIPmjNUxxqvjFVxaH5PdHdUkVnxoxcjnCfEpJjhGpUxvNfxlN/
CWiXeKqnsbPDb78uUo1ROkVJ180q1MJNbiKPDA1fiHC2ArMAsLkgLfgDO3gr+LKz
lgkxSXh6RGZfDrrRQ0QEqV8WmkpgmXqUE8/v8f+T0UGPIoCdSwpHFXyBOcLUK690
HhGX1A/t5i68cn9SoUdUKwJo74Kz8g4MUouZARtjITv1g0rvR8PvR9lveq2hdnYu
58O7+w3FlVmeTsY+X62J1lNtXWTUaw9ikERSflrk4qaONYzbClykAIeZVLd/mBMh
HbmTPyl2cXYR2FBqYP77Dcnia7hRq5xR9Km9DfwC7PrY0c8YmTVANJDuvjDaxFTZ
UvKup6EQvWdTS5nu8RObgrW5ILXjesKE72xVeMzd6YB4M1UnMNLZrEHNMpnUANdX
bwLkRpYFHoZUH0bABBWeZ3/+t/uN5A7PH8uk0qvf1/slfcLQysRW2oRV61Cq6l9f
ieUyhNUaamv6bCG/fOW3/DZTRoaM+0z+VBQdFhPQzPBiv+DwhPf653J+oGNhp+8M
amvC4xLdrTiC9g9QokD3bbWZHUyzvZgjwWAJc0x9JmWe4bu9KIweh4WNCcQkNo8o
A3xGMYcjfGxiwTaYxyx2HfRXwIT74I0pdNTGBmNP6TMwxwDMsQI7P2ytRtM45BYW
GV1iiI6l8hkBztZOrKk8py7zjxJ7KXutKPN6zBraRmpa073eSHGRe24tC3OEVrbl
vijC22z0Xo0B9raedVdoaP2jqaBf6OKaPoXx5e2/YS3wt6bV2i+VmgY1nXE4cj0J
AB1GLBDGZx8bsj1Ta4mYFpz8WbF6c/Dda4PHB+ct8Rw9xvINt3ctftj3M/y97a/5
n7e1ZqB5JvcluVU9Rz+6WbQ3PmA13/XQFoG01AC0D6WC3CV1uwAaiBEWUd4GHOpo
LJFlt8Lat3JbkigHFN8poFBJqQAdLHyTau0nInJQmiDYq904v9JSIhsF6X99hF55
QbsJNFbqOcWbkwZyNV9AfqvY+jVekoN5tYCDpt1G6ieT54XonQQVbjQg4I+uf5jz
ZS0KGYXja+dLKquSIw13Xqx8/ks9NN/+9tRJILj/bVKfxAgB6tZVIEC01NGOI6en
pTJvXpvGdWv5vOceYorMTM/d7b/I2l+w09feLfIjf4epdQ/Wee1CX8ouhagf2PNv
Nw+R7499LbNEcimiUq7j4DPoHCyqaf2Th99Er/uavmqjxzO9Ubt+9DCiiUeTATQH
zpd68oVLvnKNKh5weQWbXbE6fTq4OTTYx5035QoxtoVl93ibMY7buzI9y2z29dmk
HIe4BD4wUPDPyAJYyEhiTVdb8ZHqNavXhWmSCHtlc9yyNr6Vw3PG1Y9zoltoijIg
vgVrjsgqrzLl6LX7MtBEGSH2hHUa7wQ6ZL+vnUiwEKXxmes9/DgKeyB51li4+Yzg
Afa2AH0fU+TLYExbBa0nzqZ7TjE4Hj2Fqg02jLrEwWePnZM2VioX7raBJyEVwFui
7e7GKD7gdRdufFTbsSTUUqk2CUtXyGn/JOylVIQmzUMJbidXmFWvPLWuJcROP0hf
38DB/CDQmsN52X1q648UlYqg62szHCY8yb3IbdUd+hxIRgjB9seJmT4+2E478OJV
sN0LZgZPKPeyMX4d12JWJ8RBIKVSH9DDHQJ/OVJ5cgHO28Ylm+zpKqngh5ijeUMo
LeJwS63/fFsCOLs5++dh+dPrH7XHISLHiXBLKj6fDRvcLjOVYdcJOEm3pi60E4OX
brN7+LNZJY0VAjGNSYVdgPm8PcL33jr+dcD/+R+7pkDZEO0xd6VEephicyM6KqhA
KKtibcNKx84UqcCupuS48U4T0scGHZRDCnGXU3VFKJB4I4EnQWY/rlBY4YvMv62y
ioLazf6VtkmwYncS6nojpidZ5Ll5bI66rBCHY3B8p0DYbFXiKem/D/7cE/yrGLiQ
pymfAuenCk2gcDIfzshaOnGDXwgyvc0LxU2Ka3qN0BkZsDoRgaBUP3BCupl8GoBd
yWmcpjOAk8vKki9WVegJXxwrrjRLAx1VgvcmdGnaRSc09+GAFImQv3gSum9TjCjb
4PrIr71MoqzZLMKEKx4QBVNxZKQp2JteBGuOa8y+RHpjyJ/yk+r8q4KhTpDN4R/m
+V1lDLVJausB51OsunWdSNcIqBluCdVPrv9B96IDvoRYEvQs9uv4SLP4GBD22XBp
OMLFanXTuUgYECyXR5242FlO2Uqguls5Mi8nMpRamjFRDXGSxqo/83dduFcgJKqt
ggkzgOrTUzmhZJpGvhZy+LBtDWE8CRsGVwk9Ob1/DuU8AkvumjO2DEzl7tRbYWx5
Di4NhUrz+bmAu/br+DvuCYf6ZloqIt/nz0oNS6t4O8tOKwQ9mN2qfPGXvG14Le76
jV0Hb3kxh2SGfA5Lh2YC3XWMV6r70xTU0R38lQNM4J9xBh2gRS0ZGKBDOAF0GbSz
IhRdHQoevEMwXHHxaS7B79k6yzHGPxJvFZ7RPAVGtyMQ3xvJLgFiVs5LWQJTOWwR
usGde9o/RCya2NPTZee2ZcW4aAyFzH/lAS+2i05HR7dagqADBLgm+qoCIYVW4kBy
CWCqR/vgMX5dTAv0RBeEEEUAlZiNj/qrSpcU8/x8T+rbSxiPWdJfmH78b6ilEupy
5qee9KDa+NKwdt//CxLffoy4eA+XD4H2OpRI6LMF8QPvQwVVdvOm0XBznBQe3k7j
rN2DveJT+ZClT7RiSUX9SpBnWdV6XBjzWQ/X3CwW+xKFNaYXQAwkleKwj+hTGfp8
gluK9CbCP02H/pEwuUmq3he/7Mq+zKWfmGk7pRA5/6FA8Vx3mr0mZlsdIwPRYniS
+saBtowDwSwqY3QzhTP1nvNbTPAF2E4jk/yc8F/WyQC3VUVnlPgPjMy1VArj0Yhb
QJ2/C/qyd7W8tlmWdTdsnYMzYaso8L7c1tBKLel1jwCUEBezWRP5+czQJ3J/BKYO
vbLmidg8WD17pk/Znl4PIa688o9aNsLNR3XrgrOuk4lyTJXDO2COm2FF4FHLa40d
oNfQDOarQd0tNAadIHWp7FxHoRsO8RymFMY3qlCmKk5QzSKREuU9IGDb5e4++vXy
PjBBeEyo9IoN0QDo4rsG3U5mwq6ktk1g4S69+bAawp9MlyPCtuuRV9gngCRIxHwm
3thqfJgGaAO4XzpbGOUQUe+prYaAT8IEcxf3eVFp11JsNl66gRaojU3XEfP3f/mu
kXYRBgIsmnIndEDEa2tO37gpJjrYg80MrHl4WB37Q4WY47sqz+vpECuIWvUVMwRD
E6ilP6eycRbjXx/ZrXJQ6wpNekiMvyXIvv/F7ho0Wwd/RX9Wwr24Wapvj4I/btLn
3bAhBbUmZyDYw5W1uprj1qh58oNgc4+gW3RmsLAKV3jI7qUvvlq1BnUrrz4b55j1
8xyPsIPu5tTpiVLOYqwx0jouTaehqSRHAbqzcwyp6bzaJ1wekc6MFfxkuJpMwAU/
ok7bg3kUnoTC6B7o7BTvljWIADvBxtXBU+z9nonVvq/7K19nArZi6DUXbyPiAr96
AZKzmo5hTc0vuUHB2ZGOvd0GOmkePgpJqeHiTuzMCwSTzObkugPpgCWmXLM+BrM4
jY9nK5v0JEiJ3zcz23GOiBSQZ3MYEBcxdkWge/5VpYZqdnb6E9ZfY4UX7yDhM0sn
WVVbjk6CAcjiuU8igqw/wchPfHlHvBEBhET9eFSHj+DXXnleMreOHP/OOLtuXBzR
I7g1b3z4Nuv69I/z5QHAzBN1VAvXa2g5lVYSctqCheE9+x0pknCRKV6GNja5d3dP
Yf0c6iwHDfTOELudk5jlWTaF9qRSnQP8cFSCPneHdk7uSx+SQZh/yu2UB5iq9jaR
HIQUZVGHpQNBtjI/zhPHyFkeBfMvkA+vseFpZdKbmzxseNefIYVlATuc7MYqHU+t
5bgZswmRcsEnxj2qEEz1xV2kHdYZfAn4FpdIcrIJCAf6Kdn7JCrhi/6LbtaSAwuQ
6bkYfxi7oZ08qpSLLJVgVrVouRVu3mnW/Rpz37PKvuUDiMWSLn04nm9xobLWEx8T
HsArXi+HipEbNB0GCMy+LHUxyMbRKV2rAC99aa9XaYbv88ewMqPWqrQZV8Eqej/f
IUdXd16KsQECcvq2kH0mxL9ZemgDgb68FG7+Kae61UD4NDVKXYzbValBeZmMTmla
SF7fsjFMWF61g3GE1InzVtdwr5x26Vw5Pmj3EsarlKXe7n5AYko8va/vrLkrmMf2
g5daXHtI8KwmTGoGfikotafhq35ry588yrhxjRYegcx/iGoogPsp0SK7P8QEANYJ
GoPB0v+tv/KlxmYiUFuDWOvqPOnVBKAc7CtWZKWVm4xZdEw8xdVyjSlz0lNwg+HN
u9mEJ9nrktjZ/XqJYraWFXVbKgtGxRaRyBsI1HajTPmWZgt2XHUAntjvJuvcPi1Z
3eIN7stJFTIQmuDwD0RS90E7AbrE8UK14KFUDpDYOMuZ+OHJiAtfQWemTRpX+NF2
TlL8hRPzA6dhI/2fNxszipmNA22UKqNohibGx0F1MDzwtu2RBpbTGd0Aue5yLEVY
Rpq93gv/XOsLq3Zzi4r10uAFwDdYfM2KPQ9vjpgIWco6Q2cG5h/ZI6nJBgaPvrEG
EogndDJKHfObFEi2dqYMQkIScBqZgJh2Mb1SrdZHj5F4jn8ifHGtQBz0pa/92TNg
KBVADRmpTvWLr+0wJlhKU7+IEGJyzsG5Z2tnpbeCEhiNeu4sP0uh3XBvzixRTbHg
ADZeFJc7aBss28iNg4A/C5TPZsLoQ2+aca1s7N0XOSPCsViRcBBNts6q4zY6s2bk
0BlbXrL4oArhGdvAELn1MiK9V81+auzthNu+ehCnWpYmR5pZHi1DAYci1TMQ15vF
ST8E5XBcnwnwyBMTdeGwFuYTqiuCYSdpxdhBUVNGXbHfHadl8VL4O6V+5MBmokCc
Yjj9NNzmFgTvQjZqgPOkpi58OHXiEd0BVMGV71lXuvQwNRtbTjf98PFhzLpC66yd
N/R5oQnbBs6pMN9zHnqheSIe7PXZx69brIGDZb0YXwrvrBHkpLHHlGuFn9gtqdlJ
FsoV1u2O7PGHofD/BYJzxwCekb+St8vr9TKedoczKzfY/wWnXrfUutzkti0m6Lpd
y0+8tKVnkCiP19WHZGwe/mw+vGVgfQeSpYdX/BwgkDtg/8S9+tr8N6m392RK4YtQ
k4Mz3h1Vo8u063fFvWGMs15sdAi+QQtbcbNUw2FGuJSPlixHXZ0nZaNV7baSbNs7
F67N8/xsBGAp1nWKLae6ScoEMtffovgF5SZhNBN0gt9Chj3Ht9utNoIVXaPuI+ny
t6zJ0YFufHGkSr8Q2rHtAsAFtMMt5xXgfC326QsDuoXnBwADWvoimVtam+5/fer6
V3cfycxEc7ScYZT38ggz4GorK+nj2ma9oc8TPOltJKJQTFwaJmWCJjHwlgKl/PCy
u8Z/ifBntsFkf8s16gqFnYh0jBqzY5tmlWTvK/6z14IvfNEQK8mgMlv53I3B+Pl8
XAj8fe8NPGShEkFpuNar3bayC/vu+alQononFSQVCI24yxcHCSTgiu4lfe+0WvCb
9E35DcG+HWNfIpNj3hUtW0lMThbR1x4NzCTsDtdIFco1KoyODrX36xsSk0JQmx5k
hJVsh5nBwzVWF7adcA4PvPDUhZfEeV1bldR/Q1ehrTtyuM+vYttvZJ/HJwd3C0Xw
8yw2SNFrn86CVhfwiQsuNqplTpfA4UUeIRdDniktDjJv8iEurkkmlnDBLQKc+Z4M
hI8XDujcariRtMWgKKEbwgYDtebTmPzI6QSi7uQnGD8t4DgPpOxJ3X4u3jlwWdsI
pN195eO8YdXaMHWIfDgl4Mp9FhKmxUvUyezmCMiKsc4VoL5kkXxDsAA+LW0dmuOq
1VcLmW7JM9sdstwoJP9DVVlu0bWB74HdCoDsbUA/bHzCx51mykHNVOWZ+AWKzrh4
rEjHozdTxHtKQEo/N3YsDuTSbJWbqrXt/VHwP+C2As/lx/OQaAQZAER7NoTfQCCD
ELF5X6v6I4byiBVXmueev0lpnq2rQOynE7wTPEnFAfNil/ylSgYY2K7Xq1ThuVZM
FkRbc4WcVJdYzPPsVatqy3L7zxB4F/fJb+2wkVvsY2nTx1MXd6ThdN7zJKdEkby7
H95+zNTBWFtPm6TMDRJ/RDZmOsAvtGUno+qpJU9v02Gfcoykbw6hsqNSl9fLs+hP
2a4eEGiFqi0W79YhxOLizdLhCDrfR7ib6YQOXW57dNIUp5IaImcqgBvaWzVEZxVD
0xlIrQeXi40QfKBAUm3z5g31pwvSscymrNu7LfDNyhtpZA/jXof1dhm6+AnuWslV
JM7X6tL+fjFec7ZshVeuzLDJA3DdKrhV75xz/CSZo/Dw9CY0ZTHuoujZ4UuXY4Ce
N1JBrYS4QssxzEOIyRf52U7/yJijEzV2jDH3HgRGCdDP735xkAFwl/TlE3xPxuHX
RCd6eDBUkq0ngb4FMTjsqeR66O4tLJRh9KDo+XlxQRm24mJ3jWvM7tS0KBBS5AXX
NCHJkkVgZfCyyuIISb+AsNXigDNoSolGBAd/TONaNEyG8RRnqopRLLJra9ByO4Mm
5Tr8vkU/aoXitj7QhZKhlAkXDRustz1UaBAw2mah6+dt6P119PbaXgbNO0vmROlW
0n5Y5BC4XbQtA4GgBYXhA6X1pTNvIkZULg4ZvUdKcL+EwlfjzOthf/ghm3xxrGoL
NvXAMLflgguT3O+xPfU6rM5NgLpSuqi9HymAZMPdlxTgRUpaMhfHHHdxidGf7J7f
0nZEwmGQA8ZIBBG7bFeONIY4x0QvFtSxm+8oKU1rKVrcvpPIFDMuhjzaOQbGhsCW
Wnf2CyrJdoejWx614dUEw2bzvv+QIhhQRB2eC+BH8CugfNcl+AxLznKFlPL73SnO
dGeiaA6X09LdEmhnXcTxYGLKq67TMDXdjc8d77BQtTgvHSAl2x+2z2nODCy4ZRVF
PIF1D8L9xWvB4jnFqZFMZwXwBnMl9gNdI8dMbz92+RQ4h4Ct/FuonqZaedraIfMb
E0UjU1kT8enj1ucC30TSC25ni22TKERH4vDZzCQMMU+Hb54mIBGhETk3txeYgg77
ix3EfO2ALsPXRlbbGsqc9G470MOUD3E6vHC8EbaY/n4k8j7zGKEkibwPijL0BRtf
Bkym5cImO6uTIuzCEeoHJRkYQX6zmdi+ixsHhJulRJDpFVVflHJLLTkH4S0/c7CX
DGsuAXnSyRKK/4EibNRmYnhpCIzp0kJba3wrx4RM8XZxpYEY8ehyI8Bnub7aaXIw
0yao1HIB/AR2IUvYB7GOkv2GjwX0mj0RMo56kQnq47zk3gKlf/djos+tQcoDA6eC
0O4j/GT+1njI43oOtoz/NjaKmTlUjEwLM0mEW1tEuEaK71Q2VjVoAOxzIQL28Jjq
8h9r1/RFHIaoe8z2fJOBgW+OH63poc+6FpKj2gt1tTTbMSnbjFgnV1fRuUQAxJG/
jxvAdiAcKEj5lorb17TNPVZhYZA2TI9GzB+sFKbrX0xCFEP97qdieI6s93YZpZt6
Cz2VyH4Um7Kh8MysH7DWBLCswBkk5JFkJSuV3DY5o9vn7y7eiNLqNd3VGaUrhuvV
CXBXrjMvSVXzmRMSiGMRg+L4L89gHG0FsIunSBlY6JdHTaXRhg6cyuMQzDaJMhuX
8ymQDUzWzms9tNiC95mbWtf/x/+PBR+LjhyuAjzV0/gDALUnmaGuwcdtJVb8ilE0
J0HBMYhP1SLLaPYNSq4cSTVmSZIuMYfh7qOyoDtAlZMyciXDc53YPqnTaRIYxNT8
Plydw8XvmR0SvEAeTjuB8hGJonh0pjPNpEKxTpgKZuPx//+BKW73OElKR1oDoU5Z
2L90YLyRgPc68F8LXjfAWX8/8KH5dyl0+M0NvwYgsJ/JSbzq7vUbNgvxEq052yZS
QNwG/aj6Uq2EcM6UKo1uUZ+fYm16j4TINM6zNYZCWWmExgBd3qTOHa5F0sB+CjAY
TNiGOJa/bCf46sROcSjM2vYbr9IOBY0SKvMJEaQLfvLplf5udvajoYkMsdnhge5k
0KS4AylWHOlOpsVxWw6GLl7Xm9NxthgxV7/pyRasTNdSZ8y+hXaSrmfsyT86h4VE
045YxOoLSQzDtQFzbv0xigLHggMhne8tCMXfIJE95fB/IdijGqHpDPTD4LBGnW67
dC+rGCjd549v750ubgVh95rALNDZElKhIGmDbuGqriwOagvfzgmfoIGwW6QOTB57
yALNck/5cpG7F+DbYo00/VmIaN/qa4elKdXUjfQ53TbsNq1Q/41RZ+rUnmlqsZYi
wq8ksO0hvcJH77w06QsfyGu9S6Wmrcny/WivlXu85MdYzstEWJvDOEoqy2viLyaU
qzP4L2cD2uoSfy7G7wuSvPdABuIMUYGKjwzL9ZfzB8IEyC4opPEjCw4j6sRojRUX
r84p+J0sVVM8QmaAhdXI9Kkt02wH9IiNcS0aySJUhP2MX8ZMtsUqbJncz/JaxkGy
aaE1yT71U9NM5CfjLhqG2/+nmzdymMThQ16KHG3U72X0tYEr9s8erVMMafDP+U9q
bWEzIqHaVxKsw/7eT/0JYddJkFMa7t68Wx+Wvp0dxbKI9KiwDgkAIma81HN90iuJ
3Lp3b7KN8c0UtBF3W8C0SkyfGPK4nU8rJTcv5GDAYpVusfArQGyEOX/PycI05aHZ
xQBaptjNQJcPxTs/w+BcMzfyJ1FeiiXKrCZp4YfEBuyhsZOrY9FETt2uNqPaJuZv
khmWFtRmZN72I2YHwoM2EoDzugk+npF7aCc0jKiGS1HczBcz/XXCBEMq9BsSg2wC
fspW++zNhKNq+YJvxBauC4jpGXbkN11yR7Wit1lUHaDja/fHqTSQ5uQXMe5Fp3Pc
VuSJboNCgpoK33ryP2BPSmL92oCt2mleBC8yZVURXof/Hpg3lVD2HMA4L2hN13Rb
aO4hPQ/lcg8avnAWTbP8kWJCpexmietLo/L5tVGvFkUBjM4tvQx2Z/o/Bk/zbpMe
c3udR4/m44bHLav9W8SMW26aba1Z2sbnxlMdhJ6eAUxOVbRmMyrqBOGRwh32jc0D
i9D7pou/hbZ8ljmDpVs18Fj6HI1elwv0Ug84q5t63BmJKhCB4GZrRXPLueKP9/2R
ujibDpTLLBMxYzGfnwHftNDV/bQyDwIBpnqKMWsqjhKdbe9FVhRdJI3/giZqI0Z2
9eF874ep4RfYFsMHFlcc+qK2keDSojDnEi15dC2WULYzLjqErYQlSefF7r94AZ+l
S9g3JC+GNmMkcOz7rn2fa25QTp47y2nxlhW5cL6LAmJKVvM9NI/xvr9L7BtLnFjE
kTvAVcE+Ng7u4N5eyRL7q5LFstOSjMIHef9ia8mdagQE0rmcQUfVjIPar2bxD+cM
LobrMvXuTjbc3sTVq9HCU7V7hTePnRdD7kvvAh2R1PSB2aR+Z8Uf9o8Oe52HdzX7
X3QYlsijebUm4BkPMfARicsnaDEkGqScnuo1ioN68he8rqZPBlDBgjL6QWGzfZNr
/FrdGim7viXqUZJQTgARgj4f5X9k/Sj3uEbK8qzOM8I3hxR99jhtaRkRk3U3n/bF
mSXo3FawbXmQ4z9d72+N3N5++78bsIEixYsPvH/sTtV95PCGJOU0BQMzbEJwnl+m
6wgF1Ac6VCjFfHSp7rSY8Oo78HjJ4ZjhAFzhsYvVwXTMr7Xw2MCnQa+4XUYo7uBl
KzBvS6KEJ6DlWvtPxwjQ+YY/pKqIHpPDAOAqHFdPoNzee5LYJZBJXcCU0laDvlv4
Jqn+6E5W00P37eTnHh6MlKoXHO7r7MPGpmLsO1ZAJDrBWYAIu0EWe43RXKXeWYRo
gyNG6hC3qHbr+uNMyN6U+3THjc2TefHv2dIAAMlu/XUvKqJCHTCaMmBw/wyM2k5W
858+PSCLzKsbLiPvYr1rX1LIJyvIx3HtHhG+t2naOsj5Mwkj29Ymra9+VqDGuiDz
fHjnnTUCIBJjRISeoEcgEywh9/c8nBAwzY+PYSB+FJrtm7FqCiqde5otrMwtbEMW
JWzrFRZJuhUV+fySdBxdW1QkYQ4tp7ED95LG0iw3FKGZkh4AHX4nrXnfwOLQAek0
RDlcJUKDFquxiWgn13YWZzkE7EExcqc5nLZvo6RVGPyopo0FD7XFw74gondEj1AZ
ZkR23wNv4OYDj3J5/hm2nldKpzIXy4D7/ZM0k0q1RHkjKA/rkmj9krdfosuLNALa
qi9SE2vzDEUhhW7JVbZRGqW0wQrNWtPGmsCH+c7vh9qwqBwIIZPQ+9mwn1uC0I7B
18r4f6uCXWgfRSH05UCSgIU8y6Hw1bkkxa1dJRSc/MQYfQLVq0lP16saGjnWLXEv
wuxCPwMKa7iE2K7HwPZCyWgoW28iVS0YBovOeCjlHQf1F+8barsmu8/tvxvh4CL/
S5IgNlFGAz2WtGQp2YoPNKMUEy/CH2nvNM+YedXfYAzb/0X4nvzxuCqcQKtfN+zK
nwZjnVwVuQjkv1ISyP3sviTCzpPcvWWMP4XNLTwSVicz9vC+3a4iqJZlTwSKxCrU
ciMuiQ6SlrIIqshbHkWdwYytDYZzBFYhze1K3x38uCmdrAlc0B56+pjb7ecRZkBk
prw9vpLDJ2HSLj0Bq428XJKnj5+YqlBOEoFcINuuOt8pQSK9b7VeJGCnMYk6ihTT
bBhb/hEKNXNdEEtcrIRWnFrhxp4xwhvX5tr6zgccpKxij6DJHd1rdNsAc7vzO4OX
9EC2uHGQcU4hUgQPPxIPVWlFYxYPWXktOwabbPyTFjkyuoyEnQ/oVriJm+vdWTI0
LSg75XtPLQQy55np7hneoYgubUVelc/c9l2ooz0sOdV8Xvfz044/kSkR5QUtMwEX
zQfb7hnBSTL4vegByEijhmlO5k57FmC+QX55zG7+LmhdoPk+4EfNbXIoC0yH9J9e
birCOYwLJgcU6VPRV4rh6Nnt33X8tyEyvTjA+DVts1bRkE6NcRWgnzZIdanf3P0l
r0kbPUbKp35DtgP+3c4uAIniFE43QX+MG5aHFKxG1inEiPeeng0toY3hDhqpCDY1
kiN9cnCTEs/kDFVNg7rgyh6vmVFuhUsFsKQ34hQVNQbkMnr4nv9mknznAQOQ4HLp
FG3amGuTfiBPOnH3pMJlFU7ovNEWzl2cGc9TBvP8tj/l1zUlKH8SwmYOKnlWQt1B
ydp7Xggk2fz4ax6v2Gjxq87DOUDQ0IfkPfXnQbbTHA1wazPn5YaPYFODksxomGzJ
3q40X1eEdeh5YsqTOwjli5p3C7NP3i1cIcRmiczTg/UeUA9Y4S+ABzAv+MGJQq4G
FCEnITNa8j8r24djYHq/keFH32ZKqBgxDLamSzkb7zF8laplqLzt/owmrcgokhDj
/YBFvtDkkb4jZxvUQPY8RtpCujAJ30ZQIx8s5cs0NQZiO286CtQzYQr0lWrQQb+Y
6auNW7HU8tJy+gSX7GEt52OnCQPJjJxBpXivb4u2bdUi8gUS5txY/ysg+kj2ao/E
T2g3N3oJyGJTy3Me70eFAmRuF0X43TqibaLZYfqST/DfR70O0ZU2/x5J90ykj4Sj
a4I864t4aEzr0wRv4/n/cqU5mvGQm7KfrQMuL5PWY6f/BZy4jInTrLDt2NlK63JK
ui8O5et4ScMCm8uCkz5SUkYkE5eoL/EhcFlzZuuxiHpZGMzNezP+ZThuKbDP4Wf9
F9cXcfdb2YgzjWc/UF1+KVI4MzSGN99I2nf/r0FHbOr593FXv1ejIhGDFNzSpurr
MdGfGbkDdt23lYyoqN7097UfXHIsZHudU4DxJqWcZDC0pN7xvx1IAiYDvKTxNi6K
uluc6JsgOe/N9aVzjIEVoK+cGOx233+nGRS8aZFbzRdSz63MLOcMMshJ/CUqt4PA
tfwoduhXEolawOI4mCAKoD19MT/YF7+xIFB0VtAdNK2WiAy/fjUw9xj4khZNjoai
hz3xQOItGKVFStBPNmOetduoh2bIscDGPc5lkOkDNuBWiHMexuxr6olzUaIZ9O0n
W08WSNtAhLKDNw7KnfqiZ9GArFF7zFfJyQBYwOpShqdDUNy8Q/JcLhIkShlDsBg6
h/NWtITjVHbgmnQW3jzMF3ZLEtu1JXlMHJJCxT7LfUNQnGzYl9OZWV6aK1wrBnPj
/ca8RapnF1KSIoZ3BTHEme9JVz81JyTTumOUQqE7TeWjW+1BpLRNecQKZL3m8pqK
zKqT4quCfFGNPF8SVyhUyxTdF9G4KAee0Lta11MervTDxvwHIPM/oyw1kxEWBC3H
2Qo4tatSLst6xiVntlTTHaTTS4Tpej1WywLn1X7cLQ5lT2eAd6FCqJ0MQWJ8U75S
ycAXgD8p4sJ4O+Bidfp++FVVW9RiNkdGb0vrNB+dY82PbIfjogqxwgV32jrr6z5A
Ta+sr+/lDeeXlnejSnZWXO27Kj9BPcnseS3tHGHB6/t6f32mafJnc8ZEGKp/PSMv
oRAk8MWXc/SIUnCZq3OsgzwD5eR0F/x6FL5KwZmfDhbqNnEYauuO4JlWreuYMHxr
Tdmc65YfUJLuGI1qQEynsI2kcBHwkjgZa3Hz0Gt8zDS2BCi/M4wuODaexrsWCENO
qFprliCxuK2cS5O5XmjepcRANAhwj4tiY0nAzfGmJqnUH0p1YbGgyssc2arXw+ki
3nXQJWZguNlemyxnm+Eb2D/CWssNuxmpcWfA4I+0U+nuvsOF7abpTkt3JHysco27
8sYYBVs3ZaPtnd+IbAbLDjc1p4NGTXmzXo+CW9PZLF4+AGQeVPAOKQB7tZD+KNLs
5Sz9Ln2qwsuXp2t2w1xvOa6eiH3o+xvc/GrgwjdC+aTD2nfUavMTRa9d6lVtLPRW
SpUkWDdu43kfoIrqwQMZOBzfLrBzPUmn7VlKQF6duUmWSh8jAg9/XLBQfMgvSxM8
RwbBdjSfy/pXTFVlSrYcWaEvfNYkDlJrJp0u+k9bFyb9IPCnO9GaOUh7jsxn5bT8
j57BXKA1ZiXCzrenDZGpj6kE4ymQxZl4b2dNUJjg9j0pewQJGVVRKeQxX2Ol5j2x
CNtzKlEXiEfEYjMySt/0g7iaGUaECewwCne0+XlzK7SU43lxd5YEL1ANOjFjd0QY
+Te/GI6tVH/lS5kKyxxxQB+xA6tRL8TJEF/Zoa9JZf072KWaOtA2YkaBQptjTupB
z2CNaaZQL2rFD0oKla34zJLXtVfNT3hYJM4+0FOfvxzShluI72O0cQXCNYX6X6UM
756eOGmQ+0rS5MEIPFnttL2b3U/i0e1Mb9v6u+dtOI8et1BULlPBrzx4s5drzjaP
d5OAFV+Hoe0ySvl8qC3b9wr+Nj1WAtr/qX4eDfhRIiwyXaPQ+sNIxZZTztURl5Sr
P/H4hUToJKE/UlPp6kV6vNt45C7Wx52NQWJ8TiZvrpS3JSadx+zPRJrMYPsT3WLr
OFPPBKNNbW4vulpd5o6PnF9nMSHU+So5bTUs2g2MSIJrY9Oitx2ea9ftrjfKprVU
CXQs+9pDOp8uiw+wQd0aFKtncZF++kifC4SuY3keb8kTuhcn4Ife/WJBhNWv2Gt/
V70XpvrD4z9pkBeciJwe4aSNP1THPLtlwcEKZoEU/KRB/xTIn9Uk31piwfoxPmW0
4osXwa0ioG2xi1gyAASZuiCopsF5CipWKXYhTtGIcORvewlubHqiLbqYd6K6B0Az
r9/f9WiEyzyVWvV4ccvYisgQcmFW+mhNR2Rfd6blFEEAtRJDyH/elEYpXQj/8qLg
JN5s+lDgTkRBF46GnxV7xS+SOpqTWnMqjtOXFeFq6640SBP2KCdWX8YRY5S7Mymz
b5pukFt7xfSiGw8aSPNEjDKI2RfGcviQ3+tqkZmUPb4dpDIq7Ugx5uWp8hbYP6P4
BvCbr9/33LSZLl4giKc3ZJTH/3sbflyqYGBTYgXt/4aKXRmsLYWgDu/POGEB7eKU
HrqZbnR6MEF91P3vD24PziMIQEWHdHBME5x+iNi1TGTm2icPKXYsOQCf5Nh8Fmjf
1ygHL7URlLgx8PaglOcUlTsI1269ELWpc98Bs0jjY7uCGMXMjK04vo4uWxPRi7tJ
k0QgaCv/mJ1+/6i2rSj9Bp0fMJOSyjtMBbntin6wsZvB11oeU93w6eWyAbgtfTmw
hIB13w4HoI1CSlz+wU5oqacpY9mbQc5+kHZEazlFRs/abXe2UwIS9lfv3Sye2omQ
ARO5ysQT0K8Az90isEIBW0cVX5keIPjGEai7jhVr7ZkXHehrQQRgm/LopYbZS3F7
COFKsjbLmPoi+Sh4Yj6HMnDJ9D3/94sMIjrpYgXiy8wau9c8z9vDZk+GIerlGzH4
xVa4+mDYx3BPXVoEV0VNg5ZT37Xv0xPMiBpmSehRqXxN4CKUJQRYvvrUliPBYZD7
JLvuhm8or2WJkonbQCKXxzNVovFdH1XonlPuEBGhPR0d9ShNHjWpFaR0tLHMN79f
rRhINQl9meLtiDMgOX4jvN3Nruh7Efj+df7+aBFT1T5OD7NfdDrlazOyevw0CeuM
7xFG/GhteJXeS2fDqglJfEuBAafksdZS6qwl97grKODZ4ABtkZeM4G65rxoSWQcG
ikrrMQkrZw/7i9IkogP5AO0rcYEyF5/UhRBcE118rUxE1gGHuALPtacs2v39AdGJ
1KjsBqVHpYGYkoPSueEc0gN5ehsnAguip1KMqSdNyMwhx+zhcr6NQLKqaAb3oyLC
7Fg3GdR9NffOMTgHcgT1txFu6070Wh6MAf0Yxodd11kgPXTUcN/BvlF66SJew5+e
iD/wyXyzm8R9DFK23hm92PSZY/BZVjP7Yh34V7vyHd2szgeG7BFkuxo+qgSwK0eC
VgxUT/NiCncVnH4X/I/nxw88bTZYXzmNevtLDq8nAGjPN3FRXmrSMbWO2q0MeYo7
kCMpOFkERHwYWsK5vaVkDPq/B8yA0sqkIREyoDZMWXbLNR2sljxIAiy3Ui8W4DMQ
T3NcFJRieXCZyR7vEh8wjdoXOxVxwhALqCzgQtJ1BMz4/DeN4VyQiOwR9qa0F6Fd
uMDUsgLlqOXbpeLrXwgDmnGs11xa/9BUoshINlwrx7rEKxKxWTZgT7azhzPO58hc
cUto6xSIGcOuAcqgDRDIf/+UEHJ/0fk81XflgvQYMQ/FliHGrIhJxLzORTlSsPsi
x3eDWpGCtp7bytrh7BcSR7lqfy0JLleNWGl7NGRgD4nNBYbhS7TNC+lZleGu+lCc
+Co8segOm21hNnDVVf6H3nFHGXfOA4Ri1nQaxfqohiEmcILabhMEsy5JcnUvJZAP
KZykyb6pW0hmgLXnx6UqEAx6a9W9B1VESxzInDQVqoXBk9BkWWwNNdNyaijb3mw6
QNZBEus5Tu71WYpY93dg66tOyIhiZg0cpNSDEPFY3llV05kkStoJEHfL/HdCN4WB
oE/9HiftcBbdaKZMwdKt6dkdMr5z7zGIZcQOjZ9UplHNnUSt0HNvDUu/c9GIPoA8
95GxjnANYiAy6FWm5k0cc8Fkg6fvpBGRwz3TUXLR51oM+6xef9Vh9GhnbNPbIZrj
SbaNstFUp5owsMDMWunn/IEE2LZL/fUt4f4nhT68pFJ4jcs76fqKwW9It7kxXtS0
pvmNEP9vV9urXOzUhqlaevhGG9sHQRvoOrTm6mROaiN4XDxxyf8GTD9WSGQWF72N
mK0wIbKQ0qJiaojoi9LXz2XK/gs5LNy8q77Zc3unkngBio2vW7A7vWtac8mW8/uw
bJ+A8q8Eb9017FUCuDJXRTxw/R7oIpisN8y79TgMLmqxqNf1O0PjucleCF/D3uaW
hZh8Sqa5kBpdfcfwyVTGZjAhEWvLND6Er6tofMtqhfraRyC/lGOlht+w+3JZfTyK
dO9OZJywGuEUZszq7V6lu6jxKLocJicrE0LNtU/i6xnNa++iv1QN0BKt9z+961bC
+3eeqInX9g2wUpZSUfWMG0hGtcynlbrhHPMeM+kbXBMJQYkG4bG5NXBYgyfLNmKB
OGQetQikYiILNZuM7ydCh0ycmFlOCh2dpoRrEoe/EN8EqA6hrgSOjs+eS56qnEQr
gEJSQIU0ZFxsgRrOD8e91maP7JgyqFpl1599TUru0WxbQFJ8mlyxzQy4sIK3bpd5
dV+Q8Luh7uZyov0gEuYUOeXdT6vMov394WGMekezOZaKCOYF/9Vrq5SHOjFR+raX
RG9BwX7r8IadPsqMPrgz9NlchEW59xnQytn1C0rffgwvg1l8HWnJvwMslEtybsOa
eyDkCNlfCLhIz2gctEmfzM7rwfW0U/b/QwzvnU0GTsHwgo5pjQd5ocruZ0F52Jq+
/Zfr41ZxZqTF9dH1RiJcurOAddPM9Qe3OntKMuohqKBb7N7aDmcGUUFeAFrrpyR8
YYFaEo6YXUjpLKwKkzPEQ+KNNgNQf3dZ/BM0w1gXwgxWqN83CTP3rpTqxxh8zTHb
OX95DWe2Dh46FrXwCDteVHKTIs5tShMEf7tlx+YdOiOwFkMyGVvAbnR4+iYLnZcJ
Im5kYdukx+Q4MewD2XLWWbXLxeuWRXPCO1Htw41PUAg5PWFlo8gvB2LBJcEiEC0p
9JU9G/+08rL/zD2rrWHVUdcbHTfY9pd7ozSIsyBgIuO/uOv/fq2nKQB9SR7+1zV6
hsPZ7i3A+VqK/RAPb0ktyI7ilTPGzJwj9CRfM3AYsgjpTATc0ChxfBU+bFw26+RI
WA4HD2CGpkV1gj7e24SCfGrNqaQIQDxpNiJJBIOs/jgO/luB8rMMjzORx8UqgUPO
Ibsu8V5coNCOjciILkx4NQILKA8D3D/mx7s7aCZSAtT4T8GUqijDd8pDZVqlDoCh
vAlqdmskSZW+5IjEHeXvMShgcvZVDIqjjBEHbwQiAbIOvPE7k9dylUnQGiVnKV8Q
OL/aJJaJAiff4Ruq7j7tHQgs5VsQ/HJaKtP5Bl7kI8R2+p+A2GtSH7rMAzUOFuk1
8oIVG9/g8Whf4LBsjWwVQbw3T93xFC9jh/Q342vQaXHXAinEKroGtrzGo5trLbgi
YHZTELOsflQpNxLuVH2qESQ9zd3RI+/811OC0+T8T4jAveSz26IdvK6uU3hK+UhN
ZqcSAiycr/kEOeQbi6ZFLVFzaeR9txzxml5sA6Wi1fWWslf8iEb/ToR8NXmTl3o0
hpy8gfFai82BwgKixqL9sdgzyWkoR6mwQHkd+8/sFi/R3qoZR5laH0ioMBZs7ry6
dzV3cwZwz6XaJ46chhqSBR1/spP9Bqs1xKbWvziTGLTIBL5F4je48CxQSk8udX8f
iXsGlwuPv1scZRstzKHh8X0vOelmhTwTTyAkjW4tR1E2+uEzjAqzE18tSF/c5i6z
S2Ed3+z7pLzwaYOmpZltz470PjTWfbJ1ot259FM8KkSPZi7mDHNvtZ/vek9GHO4H
dK2DO0XfFfvHKBTzdlVCPDpFFXqOqc6+SGY9OV7t/PhDqn1ik5xhmIIP/9FosaW2
eIepi3VgoWvgPRWAJ8cyvnucB5JQrUJqM+R48xu0CVF0FOkLnYSJIXFHUUzEayfn
sxmES1UvT9XFyAGBkwZ8l2RoLKo4BAISH6dNerdDENwdGk18qt+V8BLcRW//MWRk
yYvTld5oZmr/wSYOKquq8MSUch9HY63sTHAgNr2+Gm9rfttHQmwYjYXNoY2vBoK8
M1onh8BXDg01RSZhcYGIT3widm89SN6Xcl1K+wKsZ5FoS1bvqx8igYwwhPfLaqvg
3fkGoUwP38ws4TUfEhyEGjcqFQ9bEkcUyVODSmmHiS9Gx5j2ibNa/1i9Gll3nPhC
qBN1wzoS2c8Rc8Lf+D8v6MPR0gzSJ5PgSGt10Ofz5Y1HOPcySXdBq052Qe8o1s+g
Mwr9vppPfbOYzIvPyLgOwl8kDd6p0+8gejJ8V+p6Ao4g5ReBLvNMiHeM4lcidJ/4
sFoTKWcntMETIfyfVOObt9XXw1utU0LNKnSMf7at/lzTde7oPAsFogoJwPU6gYxZ
BHH9fF1Y/sre3nYuuLypmPW9dPjvhG+3dUX47qUnRG6zGMcZIk2kizFM2rGeMwKJ
M9m0peTFiRhTx7bfOTNGYwB9ZFRm4phLVQvG1AIlTUJO0KMG8clw2PzAbjUS9zuC
1cZ6xokGVjTzKNOwtEYMz5HDo6WcLEiVZcu00XlHBf9IqKeQRhkYlhMMl+DSuLn4
K67V0e25TxxO8PuHj7HLu5mi22pgxxC0X6fQcno6aWHO7hWni10veEsXxlLB3smI
DP8DnliCPGt5COwtrILmby/h7eyyvQ7kCtcSqV0e7pl+ZtbOZ+lCIqDzZ1Vium0M
8qIRSTRY2NUyF6I90AUGx4IF0fF98eaB/i3WTo4FEorNXhSSbS79NKq4eHHVY1Ck
D8CQDLklDH6YLHiuxPTdD0OejQwySmlGQ2AEXdQRooTWgwH2hx11wOgGknzyaP5z
65OUwogGO85G1sTTgyApk8gSJD89vLIukW7Rju8smA4XyJBA81+0KF9lh/sWpyL6
M4+9g6+GAm5m7Q4HHelYs09qeVAlucDwRfZnzrlcBHJZC6t8rHIOOs6nohbJXpzC
VYm3Wi/J80d+t+/ltqfzF/6tIoFYJfcN3R3XXq2PmREf2aFmZv3pbBwzrY6TJI/v
7/Wf+Hj7NOOmHf9E9WzxCOxMHIilDwi+hoWK75sJr7mVqsSo+yRt6MHDUU/R+oeZ
5Qr0nOXwIFIyTeXcPpA1EuPOl1egovqRNv9xzQOE2xgCYzmib/AdNg/lP0Qx10/p
s5LaSokLYFkOVIcUvhDsOCI3eWqBL17p9s+Ebh1RE93kXD6R4bsMTa7Cb2X5HXZo
SrpbfZ2hen1H/dlTIjq9pUoyIJkrkKa9pukOWGqm8lIfJnZwDn6P4oDlgYvqOzBa
GYpytOwatRrdlZrqN0RvR6fPQ++VUhS3B/ALjI6XqpOl8/lMCw9DLqcbpAz+80av
06vCMCHnc72aiugVDsA4sSkEPGq27hSz3m/EJtUohW5H5axWV4/muQfNcmUjAHRj
sDt+rcu+OlmCtQ+axmPuV7nnVvOg9ZIuzkoUoUHk/OyzSpJTYdol0gThULUD4id2
IkX0Ns3HzZZLVHh3vdXqebNsieAqJBWWgu3tseX1GXcCiAj+yYUthiUpG1zQ61IU
zcAXTEmks5HxyV7aU2gbXB2hAL48cBlsTO/au57oFlP6vCmPxocbp+bONEdGzdfz
G9sJFYwX1GbABWbcihgZyNaEJXOeevFFO15aOvv9uT4Tot8aXDilqbFeM9hHjWdO
/EiYxw/Fkwhh973QgvYPu4tS3wJOsrrXQXwGPAXKJ2z9e2QnuVj263+LomTJUGwx
az9aBEQrrhu5JRepU2AkNtPnOGJ7fLdIEPUSUvfgxEHbpRiuu4X+O1XVQMqlR6f5
hVDIVDpKfrq+ELyXGjsT1mKKJOkUD5S+FkZY2+ryoa3rv+wzkmeCXCyEnwoGcGix
ySB0lPM44Jfl9zMYY0yo7WHfzQmUyGvpsrH6rrd7xbVh44oPPnsRuStvf8IR+mbE
4r/wQVuquSFwxknPfWViSk9Yg0iQhBI7Ik7r6tJZ9uxng6HoRiX65MCMp91RMgw4
LtDQHKJcqagYSVEWHd+7GPgfb/iJ8cxkzlpOQ5YoXrJOlnRzFKasxtcBAnMDNw9j
bTjQgalIR+ldpeKF3YZqvRcgUC+3tlcTT9whhyZyf05xEc9DjlCxS4mDodfP+Q9p
DhWuRcdkKLultMhdn7Wij2oT7Zf/1JmLH2kQpFiBqit8xOpRGvCvbg4nKNZPwtqT
nA16v9SiK4aH852auSTR4qWHvkawT1cdY8WmgoiffWrdflKXRh8lC2SJIWhVPjmx
Gra9PwofGvobatET7hgPAqNzY14fC2Wk4UdQfoxJSdC8xtU4m6DQGyKUUl/16wwO
g1bLfyrWg7M15Gh7S4YbJuprDugIEWNMeAHVhcdA8I2TJSSXVc67zCVLDyJxFE0H
NKVqNgi/wM22aT/hB97PFINeYTRXYExPgNvdGFpb1N0DQuByIFzxCsymk20UQXST
h1Jf3zj0t5GLLfCdfNqFRNsAGdvdeLs6QLeoJZ7NqrcxFbpC64Xl/4655W9qDETO
gBgsXRmQZf0yIqVbX/ipaporPbh03lvrqzcSduXyXwPfsxTORcYJZGm1qnweVt5M
uo6Qzeh1/v7Oji6M4o0dN2a5G2dA0BAj+fX0aF8JHU921xkIOULcqvHkTSidBbGF
QNEfqwXa3SApogMelm/awLQlL7LhCd5n6BQnRVnXI2kfpPvkKLdcRueUjlqdUhc8
tGWa7KjNR4zfAbZ+PQ8364K7ZBRfI+CsIgpnZvBg7sv/4ST0GD+7aXQ19G3RcJrj
GVa60Kk4CwzALYouDMjN7Dvnac9NL05AubggQzazbiSdH36AslPgiININg1kh90S
7I0Y10bia7X91etDy0ri0f/br+RZOtiuJF4xeyRiTIUcaaAu/15oyepGvfEJSLXs
h6P1FEBewUb87msFhKYGgIom0y0QMG7HLdjtlr7MRnHFcjDUmvNadfrUGyYxsagw
j35odqa+srcQSxP4t9GCMgVTkaAIkqFeiIvWSLH+O3OpfbybG8Mx8lEU74IAcps0
iq9BW5ST3xZz7NvppilfzoiQXjg6jbVZ/oA7Hm5xvPEt3ayMG5JlJHNJhA+mm+r1
YwAyudJkziM7/nxaohf6rVRXPrnplbHCloKRUpVYQ1hSPE/Ka1SgUCm1RgXd4pj/
H5KvK6pW3GCPe97uVO+wKl9IDTMg6i+8w+ewiorRqmqup9sZQ9zIfYT1FQJB54GJ
GzNm5GgfX5aWsutslBuhCxQcwZ5z4bFxvaniSN1djlro2b0BYCgqoORtjhzuEmbh
5tCmqAWJL66/GqQO50BQLMrrXmj0l47hf+zOxQdwXyyuKlodgj/UvsJDKbtBwLYD
agHw7bSKDhSMs3bnfx5nnWfg7L7wxVtpc0D9xcfuesqTjZpcylbnBOu9ymlEzQfk
6uXpT3cWPwLBndjgo+UQ3eKztMxMgWOI36MIL140WfP/sGAsKsaa4m+KgztL7yLF
dxiMpcN7CHfTtNzbChs8mi6wxVdwju+J1OVPzT9Ds3aTOEZMC2rFk5KUlKYDd+kY
9zDa+QvrF1o/O4hCT6ehn7g0Ncic7+Ah3N/osf+LvRd8U9JATOjIKpbKzkSFCLdU
fcs8AkHW8jlSMl3YGPg1UEM9494kPaP/pwWeSD13PlBglJspee4hk14aEMKF79Sn
hjAgSz+mIsit5TFmPSLm0tQuM9arXuj0TRK0TvQb99i+wNUetGqCUVUMmccPF5HM
pXVmJ6EwNxD03aHPzjgO91mCGYlH5i0feVbePjBGJXdxc4njEmmeyy4kfAaRf4HQ
r1ZHjSC4DUH/UydnDfK4Nmqu/bIScYGtoh/0gX+99gQ+ueapKb1yWsE82wZ2Ascr
0bpdhKdhWU/UkbrOgpaZF+GzBs779Zyv+HdtVyqR2hhvoml4alQxHE1O5n4uzzOi
pAcX/JR9xgJn2Yawdg1W3QjFwyJj6Ki4tLYHatXPWO3RMj/lhe9t5Vz4bFZI4U2v
zDBobC6DNJH1o7aCvls5VZsBa6PJ/iZ0G1junA2mXczG3Hqf2qF6kDjfUxC3VyA7
xh2ItPnoVaipovgXvrdCBOH0o8nC6FqiaVPrHIv8KBLs37aANJcoCNy+ZBQJTwq/
EId6qh9rmnm/FVQE8J9zaJ7AMTPdiWjuDcYJr2j18GYuxyMrefOac1ACRuHkwA34
8mzns6a3cJPq55zqndEjqpyd/5Il57QoSfwgYk3edZKhEIt8CxQl52xaGB6z1tAo
yR0sVNiPyodBg6KqtgaCcmy4oeqBLlATj02d0hrOISCtR21Alv5GKWrL6fX2AqSC
ud85xMAx4yx/jVXdzsfLhZF50SMBfVPI+UHHSf7Sx0XEpz6sEwSjm8b4yiyy3UW4
hjQ5g6Jpf2K99Nvzu2bYAx+GvV4M9RzwF3qxpM+vuJPWM2cbhBecN60vh6mdZXiR
N/AM0Nw7V5gHTxHyGTWL9bLAlFhXURPjm90Y3k/0cnc0noGrpVw6pDH02f9hU3SU
MiuW0eCBabNEFj7CIjNZNMFqUfGOISz3Jo9G+m4R2UN2LLT1GftBIxCY1kg2CYk6
W8vhDqskYkX9knsk2o0X/yHE0jjzz6dwaN+ksU9hS08kcl63FjQw6zvT044hGrQf
P+Z/7m2zaaTFaAx6tVZBIfyk4rcOKOyM373SehnBMNxw3EgnACNNwDd4MVnDdGR2
wo2ZL+J1neq4a9ZP5WdnN5gCncQtk2SMbT6lfXRZU84En+9QYH0ipTj97lyL20oy
vQmGxgSKYca4G5JTBvZj5f57RefrloIgEPR7+Qew6hTscWatrjUYxhTWq09FuTZD
/cAiy2KqBy2czbN8HC+L8Ku7Q72V0tZIyFpyGxy4mfQOOHj/2lEJMgHuu0EOe86t
WhnrpRB+O6H1GYyxlze9Go0b7TcO11jMMcV6/EMfDIvvhQmUW0LljwBZro/iebDN
XcrROnHkcszWHapGRX9OHWBnO0v/hHwrcKYwFZlxTIz0MWw3fhvrzgH1sG9aKNAi
oKZOwn5PCGkNei1Khnsr29D+quSrvhY8Au19qPciQdomsLozYAhQYlSnFACeElm6
gt0vpyYn4oghLKrNbCFxh2NC7LTDavLqtJZeum11Yq2T56XjN+qZjfmOUxzP/nHe
9h7WQCjmBZP3vEb3rIXI9qT2lBXZj88Zk3hbiVOrriS1N5FLZA/uALEYmB6N1d+b
nVs4+MW5KPDkDTM/Fak/QWKrgXZCmG30lsDgwu25LyOCglXnjCHxg9GO1XPNHVi5
uSyQLEeX5En1FyNKYw6JxuHtjbK8qZS1pk7XyhT7GkpAiC/W1ehiD0RNiW5KGeX/
rrvAXps8qubXhOIrDxQJYYN0FdWzFIdDv4coPMaOmYTjLzRTsySrESGdat2nPeYE
8/Y+fkoVHJHVAnlybKe1smk9SdF9lgyzR52blDGQuEUrAEzDo0fGClG2/Hu6eG1P
76yIr3uzyfEkMwtGkio/DNdlSqbcpYSJkevfr9bMxsYcT3VSUkcmDT5YnUFa+R1O
oy8651fKu+Gxni0dBKtogS/lhAoevevpXnqtcOyg9X/CoOuq1NJ0iVWd+K+JAZfy
jymRiI4QWn26ds2rlHak0tp+rVMg3pYfMpP7hRapQDdO6aZeTHpXT6boIfv5FaQk
l62UUnO+5HDvsC4uTv5iDSmlgiIeh3T9gDCP2pDHPHZ6POdb+PWYMEkPl93ojqou
BD9GQZKHO8oZ7TLwLdGHz3D7YCTtddvMNmTMOavqnkAMZbRMvrY2p1qCq8ziyi5K
3dMVHmjAnxQq1LnO89ckS0uiViL40+Qj5rAUgyXdsGJHT5qUKpOCUtk83e668ZgA
bV2PKxl7r6gcUVBE4rrkhDewLbubGb6QjughgeakwKYa+Qxtvk9pq0ehiWIMwdeI
wsj/DLL3PNBJfIMiZnMERuEnUQ5O64bK1+bARFxWcRqJIjFfYR1Ip6fryTjH80O5
kDnaUBhi/kJ66BnUPUEzwRBei87GdejX60rhtCypF+q31pjFpY7QdAhU4cBhA8Na
ajCGjZXY0IQtTL2PzJUjjk4IZNwJNgl3NC7YvjM+6ScE48Zur4nbIfZh2T2pC+kr
HRFUwiKJtljERPg6oNBR1HyluJkhinWvxSh3fbSFhCyiamM/nLFw9ZdDRvy1C2yJ
tGFgCa1G+U75G5D7y2vI54tJkzmqAVunGYlVyP4vrMnmHXckRXqaIhRd9/ePeHzn
DxiccSXMkr6OXVpkjX8ulrQLJ03IWwkKKZG+gEpFzPjxxJ1P5R4XkXHd1k187h1P
udEtNeDj8tMm2WUrH2+Yb9XygNX6s7+WgnS/zexA/5HlwKkm+JeK+/p4iOzZCby6
O5fBB+wzS1JgfH4WvyoB7PjvicZ456+qfS2OtLKxeo1kV6zSeiPQuPpi3rNnBrsc
HD1aS/wpX9QUv1Yn6bIQcjmi4+FXhSQFwK8sS6IUR7sNI38fnwkbNBSUfZDNzE5b
NC8FsQRVDqWfOfS1JCD9rMvAPYbCgw/+91fyVeLEAt0avk5z3CGcurcKVlhHwMcx
c93CfW8TZ4Ig3ZgtuIjUIR2aybUR6eOJjQYyihZE4KoDUarIniNhrhZjQe6eiOzr
HUQw9TA5P2WHXRm4BPhl3shBJ8k4NuJRUcn7GkAkgHPmjWX8WlEfCBPh5Wsaw+PJ
cJY0dVUOfHGn91L0LQCprrL0+hgsY6DKvFgDBxyOBLFFece/2bYYxZ8YuPe55GWn
Dqm3YFIsgafrqxHJZiPu3muA+FvgrJAOIum73OGDcYAgXAG04aUALPFPHFUrzLmw
7QjBrh/4+qFg1KsMqfVyzyFCFKRt98ScZ8dgwbKmx4ePZYboYbQxFGLOrCCZjv5n
co67GdiAwptg4wmoNvHwIJb9WFWGV9BrmpH9IlefbdeA2iX5mDDDEKzpOEp1DoJJ
9cXda3JIDRfLg2XE5jty1VuLhZycW3mvuT4O9BIqt1dpXYUV4Zvms/qnYEjC/AGl
oeySi5Yv4vbkYjNbBHsz076FZiVLO4uv+WSHOSj2XJ3QmNZzaf4l249eDySTrYI9
7mDeCLXIMkb3LLaMHKt+Nlq5XeEGC4OoYWK6ijvRBi2BazgnvT/p4ZtB7FtZtybc
OwzpntKIB1Nl2M9qUKPzBhU3i0ttVs4zbKBNvmxSeqp2v4nfHxzBdozEZMKF1NYe
UNNz9FuzggINO3I1BeU8tCZhvMT2otp5VVsbXrMTIDu/TjYjdSuUjGZpmSLJX18R
W9++9D9bFXT/TCDZ1cONQCYCGfXbmBFRH9JxcHl/osvXc7VKvxO4ZaKD2wn0GOdl
D5oIhFVB3kbl9ujkDGh3/9jjF70DlnwY3prb5BS5YT2FbK8bDsNJsV6EcoViTpge
ZP6vrcLmX5D0KopQNqqd1hv6uQ4/y5WaQ+/E7RmyHmvu72E5wnmU1YW0IWYhAf/W
fuLzN+gda3yG0069qSqntuH9GYSao2aURX0YSpWXDvnWVGSd5wRHPf8z0hK0Csyn
b0t281ylNPuA8aUmFrzbD5CwQjgPSm7X6QMXiLMRJ8LX01bp8OmBb2ybw6L9FhhJ
88BonL0J7T4uMp2Gwf5kLDIW6X3YOfBSZEtaOYMlv7cKvENonrbi8BFQrJM8CK5G
6/LZmiJqzgKV7SnlfdvDAeBzxrOxdwzVY3cSmyf7YOVviWPFh9U+c9GFoGhlgCVg
Y9FxjMkx6PGMCM3v4fjtYqRoGkm7r7U7ByYbA9NQvBBSlVIi4VgZts2nM8xEcUaS
YBLBLrOoTNCWBU7RS6ZCI2i+aNatUWsE1jdCjCF0xnToN8yLaSU05V6ma6CoMk4i
i6ZpRnq/VGNm/3LbdtY1ni9hSOYF6T1O0/b3ZYm64bYjG420ZhH/+PJD2Nq4SojP
Cz9yWN54fsqJpHZ+VnIE4j5UlTHwJMzavcCel1TUkQAulgircY6qegJYHtrQ8ph9
UH0c6sQYJ79BA8yrH+abuLPR8pdaMCwl534L3V9QAutIU7QD+o02r6xidz4skTxQ
zo1iOPqMDM4RtskKPZX5njm2VGlXG8jfYF759vwMsbaeIx3QFD9bY8wflAs13ina
AbsWIWLHSjPDYO5XzhBssidTodguKza0Z+RGqiTlp+scBtYEqVGLH0mBYFJ4Jl55
Bg2T44ql8KE9kF61wahOQpYyTZOqB2AjTy1KiOHOBqjoQ2W8f6Mzc8uNEmCd3mQg
A1XKGYoLpnowjItPG4W5mHATVN7ApTxTsE11WkOhLNBBMWXrocN01GPHkVeS0Qia
k8S3oeGTLJNDQL07jqGiph6yrouTa1BaiuXIXqMWuxV6FSd/jrErjyLHiTYdOkxo
w2UqQ8FUXmzPggUmshGtEDhB1um0J+hFF/3Lzj1ynHtA4AOteVcYBlfIZGIN0Whh
Du/Ma3ZKKwHvL6JrFITHBJINPk+uEu5CdoAv92tbNjd30u1QV/pGoNalnxrrRQ9m
D0pZT+x3eVSMSHkMziPLcD654SEvg76S+j+BFGfGz5HjTJbqlNq8oWa21TOWKPrQ
RMBnjOaFNPblqBMzIn/oK6a3bIQcQx8B8IfI5mGtMiSwSXEmydbROKQKwM9e+hM7
dd5f2QxgsyetFI/iYV94z2Py14hwvaGYpAQVqNzOCN0PAONceNpntF/mlLyssQoR
+aJX2j44cBa8oIKrwp2+5pgsrP8k2UITQcGcvelTFuAILe17vNoq7+2eWFYsQQf0
6g0F6Ey84jrmBIeVDQx6owyFnChnc3k4E7pkldGbiDCmjSUYWBR8rKB8JKlUIM1/
hmQwVeAilw4OT5eT+XAT4rHumBwsfPvrPiNwo0gqLVaXZzEu6BqJAXqE0ZgtL8vz
YhKQQ6iWYFqzknN0KiCnIJT0EC1iuYqS6/we1T+AltiaKB6DMxQJmEJnJPOM+Zcq
P/G2Uuq+xHH47HyJgYmXcpLgdYnb6xlqvpqMW9O+C2Y6vPFUyAJdNGbT3AfHXzPH
5g1PYnzmg9CiQTEuxCpDzGTCGr+nWSFpIZTFzoNgn7PsLJYZeISHmTlhcnoGA9vP
IuULNYJgJ3Tfzyq8i25oiyFcoVs+w0bn/qYD0iNEVEet4Vik+hzZgRzkniaxo8P2
SAguMtodZSnD7vZjhwmjUZuE0NCGCWeI80efVUyeO0RX05AyF+QH7T/MTAqRTHUp
P4fA1rPAVubRmG7+7pclpFbYVzPA26/354l8Qg0/YDkmKL4nZqnLA3sHQ+vIclI6
ND/Kd6hSQ1LUbM4qlL4jGDjC30pVFJUVH+v22Wjsq9Mbyxtv+fuqjdow8z4+KeaD
DCfkTbLe+MdHbtZrjpnv5YtFll+VVzydvopCymbgKxBlNpKg8tIcKkeGgvzqCcpu
GLLjxkkE8m0xgxssShwIRB9VmJOqXnzDw/7hD6h+CRdjb7dYnXaym5jFu+rYgEW6
9pP8XcDfi5zp02G1KjH7VUOZ7dQy4t3Yip9uXokRy/UcW9hAsi5t7pajIjWMcal5
k6KfUNbEoryvFvIfddoLPwm5OPfkBQqkRjH2zMnnlWBgsQNO/D6DvT+XP/0EXnNr
T0BQeSMJ5uJapOMd4bUHPaM57RSOUN62wSDvIeNzegoBhDmjFIjgqQBwG6w7e7Nl
dE4jOecV+/FT775hO96w9FZO+8b0VvEGa9v5rkGkb20Sk/J/WmbeC/fMwHdYteoH
6TSh7/KBe95LlXUrPFA0EJz2xcCEG9KvdkZTef49LHF+nNyjFJyg5cD2VXdVL8Kh
bUZPoqNEmtyfhk1Ilf2QnUktKpoeKiCaAdUYLf2nr2N7tuNGpym3iqOVMtGJvRvv
xlIPievXpahqdBen4s51RxUlhHTWmvNYJUjQnXnqr9zv7B5BWD/+DpI+YHcCGAN5
WPPcJARvMf/DZMDPTm7Wjwi94gBrZse9CeiMmC6rw/sRdhHF+uKFi/G+kXMmK7YB
VK6jBvPDl/TDZ+50MjxYyrE3PYwllJB3cey30eAFL6GWW1qAc4G/Kqq4NfdHfR8Z
7wP0p3P2N3RrDTVAViIAt3XSPc7BiE3H40RnSZI6l7jWusyNh/wVRj53aZbyOQPv
NbRcNt025Kp6kDX/HIGzanvyY5QioupEsgoY0mnEIaRHVpG2lVHdrhEOgutt+JTK
Tx3EWDmgRamXSP/S6vPAIPrVoPfOa/1uFoXrV27HnKmqStTBNzywfCa3vZyjYkIx
fhKzjrceZn9UxchUeobazNJ04rJGlD5Hkli4fbNQKoOFOnIIh1c5TItn8CSl9Vyg
8FPfQ2GVq6y7U0KRK9PIvUmUAHmnvp/mJ7qKrUCjH9f9KSbHjWLlaEhQctig4dPY
RF87+HtEweg62HX1L2JQCCRvQschnsHmWvlu/cYYgssZWcvAVM/MZPz+l3CZMogo
PSncPV5n60B9+wPws9l0JjcV5k6fvudnBxd78X+1EZB2SewFH/DwqX1Jp60PVZzJ
woZ2PQm1i5jQ7y+7iYTHpueGNgNCUVJwaXfZ+Y52TuBYvUYgm48Sh+AO1iyLmHYW
bIPzqNKfU009uwqvlQ65mCItjKgP5k32ktfgtFH30FWgWIQRqsxM+GH+FWb1U1pL
Ja3Jx4gr22whjREq1dsEaRcI17aeclnlOEaKsa82oLQA0R0ZB+okeJ5QKE4b24wY
V60f5PHqZ1oowBGC4ov/UDbBoAfifaINx5jeo9g8RavI2i8gvTjY/tQAX/RkMG3L
eaMqbEKT0L3a1ILZcWAUZJGrIP+hdpyZPmKMRn61eUXGDHRZZxbTvqB5t/54mnjv
usugyVJfpuN5bmCkXKEWzbhiwVrBzX6RzgMahpZLWISpwHGCFCgq/GM7zdJZe9CC
xX4Lz6wbytty8P2CoNdSapRZeRX6Wmh/dUu2ukKUxOBeS5Aued496W/TPGp/Zroc
Z7HkgXjHFKHbcQYFXrcpmWP7KLFggeR4hXjFaB/jfchBwLoDd9v9YSky6eTaISJa
csZ4eP+a+fsg2091s9k/Y/L+MUj6bKICwGraxBTLAn+qCxIePSsu+LwTQwZsuS78
cGatvOiiLaw7sg/zaOQV38+81MYqS9aIqR6KfJecXuo1ocw7nC4V5+ypORHpkNTh
iOu1aoiV3MsR+zLC24mlhTLdrGOYJJuKzkItuVfaiPxD0+BuO+XFbHsGzA1+w72G
+hjK50odBBcasnlbBleNzpKbCYtbIW3BdHAQXvlCSBO83jehUP+JCAgldj2uU4sM
Ee66c5cBVh0SVdhSCHzgcUCSgY5n8ARyvz44i9rGKS1qx4jrzraDtk8S3CL+l2EI
FyR2A7nmZTQyw1btbUiipGS2PtC3xM6mjZZi9VmaaAEzooLrkWWx/U3ueNyTJAnD
Ct9A99+DBECIivUPAwMbRdH4McRh9T7UfDQwYd5+wkf2ucOBNfeF5CYX7vHGD8Vf
7fVsAhnEg34wR4BIfWUPwrKOXYIbIjLXzjxSGFLxlcxH7f8hfeat1P5s77u7PQS6
IfRR+bFLY8TbvX73l1e2A3sM6TXMEC86G8vwuF20eynEnojucf0U4WmCKW9AMGwV
0xTl0PalTKXpZZdyCt/0B12RrMe/yX6BZYEi17o/HMkNjhHKcLzd3C4MG/GT+f1K
zGaTcFrXzhv4818I1Fun8dSc0YkNXzHSE2tH4YYLRa1W9EX4HtQN1ib/h4DyRNa3
EYOlInJEd77Puc2FazQ3NCu5K42ldTsEskvfoLj9wVsEVOEqj7y4xK8yE6R7wXII
UnZG0AnWdf/EzSZYmWtSilAyS/k7EgXdPej2KeC9tRUzTqgWb01nfGtR+v6cshOJ
TtWgafHDV9+WkrLamnSA2VVkGTXor1cE1xfUY1apYY1G2ozlAjslLQXOsQvsYIcN
i8GcbQ5saL1jA1mgTdBEUjIcSL4lhRXs+uQwdjiCc2kIKLR2bfl7/PtIfaN3AayB
Ww4Nmn5F1hznPjY3nZwVol+5WoT2Nhy8Wq6jds5Ues1iPAs+r3PEmAJsl5gEXtdf
ywiD88jn2EAaV6mxbnB3FzJ7y/FWQnZFSizmLXTy0gV3zbir/vW6zRrUMbcpqXvc
r+UuD8NKz7DJMLTRwGtxHhi7xpyh41gBayRI7MV4CL+pmu61O7nnEBmNrb1U372e
USrDCkSqabzzEN5YDdyYnv9Ta2M5aYl/+DkwiHfm5TP+N1OhwgGBtdaMF60O2b6s
oCWA6xFaGFAMEaltMKaD6KP/+tcFqz2prP9MdEsicqb/jdVHgGVMrPd2AWB4UwSE
SQfph6m+eFYvb1IZKqA6DrvKBzOD77mJmQyR+zizJKSlNnD/Ik5i9+zj8FQmPM6q
VQBxpyDEoMKHD4AgjnpmKxsG+2pNKvi+7dRlrzY+eamsqtgrSWqTmGkubRbPI7vT
NFSLWkPNwQzcORJC8eMcyWLJb3ftgIzw5DqTQQs3HtxfyZIXYIo/XWd33aFGp9JG
BRDIzN8FOHUwzQghmNuC7JP6qp9IbWMCZvJ9UBinznrhpC0nZ22pO4F1Mx5E86Sk
N5F3wBtWtyHq+zoSSeYhYtemwILgmzuDPUYmLj47XPRYDgsoIxjUbxVhyFtbIMMx
ZACVcZ1s7l4sSToEW2MIjO5+OsRHWlKMGdTlWurOebnz+evQnNJ78TacA96bjLKb
7i7mJsk+8r908iX1KaCvbaPJ0g1x6Uz2CTVKlccouTIxGj6q801LO363fmvZgAWg
4Kh3qMJb4VW/jq40n35pWVbbIz04GA/vprfX2633U7h0w7P7DPJo5b71r7fLdVul
I2vTOXhUJHRldCN5R/RdtYhDMlrDqoZ9Huc8O1o452j8pUwaD74bU0km4cQiKB5O
yuj5gibuZbqMbD2vbY9UN6wS/43ElSPcYhLuhbwvGom+RYJt/WJDBlkZjJC28/yY
woyK7XRT/URG7axwTqdIsEq9lT4DgryUMjWKT8E80rs+iyeM9fw3yyX8tWd4ijvs
gE3rxfuNmlRr0KMzUIQ9mtZdcuDNIxvb+E8rSSiEH8K6/MKCeEqhoEe1QCL9VnVJ
qSRp/g2M0K8g/Xt2QThoJF/KjSNvEqPmmBM7Cf7Fu8VAB35lJfKGsHGbTZB5fIXe
cUuavoECcgTPXLLSjBqyOA/1KdDmpVDmk2s7NI27vPoZkGB38TVN0dwiw/ODlFyA
nmDvT7QN3gLWOWNqdEn7GkFsVRSo2tiZN1GjwCI/P4piMLIKuxn9TDTEpwK9+qa7
emAKsCeJUsoRFjgDsI6sb3/oowmxdNEKVFN3S1r3rGq3wjpLvD5MXvimJr2jNu03
+T0NNVN2csxkMHJUfc2FpV0giEkkjVjPJCICAc/KaKJ8MQnJuXobrBEzimLC0KhT
KpuBIvSVibRp0qKIED3X5PHyex9dgErnx/DuQXcFZpGdEdEukHqkaijOzhl+KRD+
5gHo/UR+DG0tjHgSehs7gyHTmw9wpWWkfucwjanN1eRwRsFPoRKj4XCPEJIdMm3y
IZrYXVxoFl2fQ5QfIEuiwODbqZbJm6e+OIvC+C+y/L3Vwo/gxEnsz1CVZ1nA6hLy
7pjGHRZDIXoYm3AMQffilE+PX0VV/zEQHncWrXVlcpOT/B6xcV9ETE/P1yW04vLT
NV03L7eNFxhNIsCXCxi9YgZS3ufpU5qmziCBHRFNPa/wEDtwWur1BttNLQGB17ap
iC9McX0niiXKogAdzShU0zdQ61ytnmxyVwQFaC9OBkiUZS+C0OtEo9xeEdMZD3+e
0fEbPkbL3axLEbGSqsUgXsah/JJuLKQYM4uO/f86WgQWZPzdwsysx23UPWDm987y
clmReuFmJqN8aa1RvWX8fQuIUlvrnxV9OIzoxA6WKDmsgFdeJ30SDcUVLv18EZjb
TCntYQh76QkzEaiyLb37mIJLE3VKs2YKeJbgbKotwBuMRMM1dZQjf2Nl7rMEJp1G
/rgaTr4mHd5kpb3wgyrGmtB9g+Bl8vPhBMle7Ey+6HmYSVvCNQCYIXkUxQOArLzj
r3UzKKEoAL4SyxVz1vVCSY81m8ZSUxaG6aNINlMOP6mzZJCaSzMrZ94iw+NqDTD4
S6b8mG26ctuEwQFPvc8M/j4y3yZGG5fSFj2PrVMlcRyWUp1TRs++FtaACHqBTXUX
YOmMUnkacCoxxt9ClfWolUKj0in3AUe/xo8HvC2FBl4Av+pSbPWDc76iB9CIJ6+w
DDcjipa9ctjSbgjU/WWLogCouQI8JKXyQh661/gSYtX4b74GunW2Ubwb2XiJhGur
RLDsrcIwP/TwLwd7Utl5IyKN12U0+TNrlSlrFt4WjWgNhhXRPSVDDz2b0fqiTsSr
GAY/FT8C7oo4ZYJzjpDcg3sreIRR+DEfI935DMM0gh64T0gJ8wfh+rxriaiIymsM
5fVcdO4YtPQG9iuCz3OOOfQ7HcGND57e/UHfcJJEFDK+arQeCXuFguhya0WQLA+d
LD8VBqbEYDRyPXNfZCUOICWaOcXSvFF+jP5HUeTID3s8Y18wlGCh/QP3mfbRmKRF
StC8wAblizedAmNrhWX59Ao3itdqvkVqEnLb5+OKsdD5GV/GXcmPr4DXfR2kz1ww
jHLuy5Bd5w3IF8+RHCsISEVD9CArogocO/348Eug/mgPix1zv/7KUbSMb05lDKn0
91rgJdG+NgR4XyYJVP6GUu9w0iZVW2++R0xq3P6An8yEdhmH6RqILR2tQVsXPmzb
cBR+8JI2PK8epcbOQtEboF8ixJwLJVkvzPzRIX2x1/AjQiHjM2IWob3l0w3xgsMe
uP6hsGKeM084+mamqPgpKIP5i3r5Ymsx85nY2Pl2B1idl8sF/Qp6bM+UoBU/9ha2
oihxzOWr0UED4Vh90okF/9s3TfyXAGu7mbhCEUGmAy7BM3k0pXNHychyn9qCMs9O
Tk7cfUmJa6gaue7FlQav0BJia1y6DUEGX6EkYplZM6IYGu7hW67w68eMiCI1POFD
pqdcDeF9cVsFj/bi6QAMZn5LDbkk4u2m1J/8R+7WUxjHtG56UdlfjZZks4VDtvS+
Ni3+piktKsSDEiDBWgfstNE80DMFVK2WB1ImHM6nXVPLWwcxJdN+3khoAqaDAtUy
qHOPJL85hU836e0CaUHzZ1tHbn2uMTImAQ0Bva+ZER3uoX0T/J8AqGjhwK4gr4e8
BlMeFrYmKoXClSxsozicZkUZBoGnraCA4BTE+BfwcKgb6EeDOed/eweUN3R9Hov3
QhTUj7wBRn0T3KNW2CuQ2yiRYG0ahcVBSsU2XXTOozAH3hQs43QmY4SEExYOe6Yg
9uSaashJd8s6J4ZH1wUOulh6EJVTpqkEsaBpskYOgqmTnofaUtHEzmQdgdwTyuxk
4jVZLQDjsJgWijjt3ng7Mgz4CacKV+DowLVQizKJllhHBN1q53gFsuZ8CQBXOIN7
OOhWI4Ph9G0RWdsiNoaM8p2GszrpDG1tosh5rx32C9mnkWoHyx1ftY+xyuBDqL1J
yGLJEaJBf1IcXrf0N6HFgUob3dSGQhHmgIRULaTvdoiaYzdRDT5dlLalcQe6Ag6H
no4GseESXHp1ZeKv75q9NmKHF5+Xg1/qgaHDsnW1c7SLaOlcqq/QvBBw1scD6ivv
0/DrAmHCXIbBRC/7sr9gKQ0mqdhz4wYehVOLtTpgcBIDwMvhY6pB7ZSgR8j54f8K
4K5xo0O8ztUMu5hjpGqI/wEYEzjSJsiw3JQimaR6R8QgN8LQ/F5LwNOmIkZkAJpp
vEOwQ/08T4UMINckBYjK6GT65dP0EjM4EEyJa+ySExMyfGRD+cWdctcPzWPizhUN
5fhHHmUhWBc2MBaU6Cjl3IzO1TvyRFsu+zzt7j61eWPPRAcGCWFS7u30z1uM+Fdc
coDvM0RA76ypUE6FjSSBQ2mb0BtYiP8Mij9eXVWCN8FOKy5Pne13++lSeik2wzgP
+wK8512Zm9yErqWQcQNjd0f4VM5ET/q3ddrCedMM0FCu5cZQFnpMgUcE6slog1G7
iP27fHzv+dlG1KKZ7YLb0g60oMApGvj0gFjuk2mFk2bdTpnuGZG4AU+pWtaEQAiw
QSIQ5PWTqKzrsWxCARHLI5fvc+WXmuLdeMISVorz7CFlQFQktTtBz8+RLUgjlb2C
i0pc2uRLvNjZMk+vMjpyT4sOgiW2ycMCixq3EiOwAnY3vrLF995YPhur6svJVdsB
Okok/0iwFBaeniuHR4L9yOdrkSV0MRkfcLKnkaD5q4EPTf2wPKa5yrAx6DNDFBX4
tuq6qMNQxNDju+lcjDrzaUmS6fCitWy8SJ/WgXK/iqc1n7zJVj0XtirCl1jG4Ghx
anP+XBTOWUemvnyIqsP6Xnv8nid8kA5oqKpMEkiNYLYYKVYeFwVIsU3vrCpmTfOZ
gGEMpaLxHqK2WLgHacisaAMLBzZvisii+0fa+nXKsSTcJUUg9+9qeGjE2HSupsiD
ruc6hM1p9GrENJ87Rcg7VzKtB9y2bNUYA+n5aEBfPa4T5HmM00kbA3FUZ1UhcSGm
VOMIY2VMWkwHY5/1Yc0qe6YbLFmV8y35Me+Wh/R5SHJ0QLz1GdUAeBDUTNUdKVwT
xuCNBJQVt463VvQ5cmzyFRXJAgbg8zLVR6EZKUgekvBNitsv5EZEWFK5u+Vl1lDk
TNdayzNhd4TJYKhcRXYObjZxgX5sfEldMwij308CxLdO9yLjdpxvsAr3nzn2wtNU
TpUVO34N+ohBQa1Vys7COyseRfcUhzW2YKqW1m8FGeDB1XOu0v+yj+xFgFwxT5DE
sUuDU4rurZ7nZOgIOeqC0eq3lEM4eXuUNtVur0NCoGRpFncGg1Nscdnp9/VJPX9K
ucciNwSbLnAXueoo0ZHGUHWlf33/lziXRwJ/rsUH2M/inK5H1uXDNfOQJnAatwHp
Royy3yylTTxGU/CSUJ4K2r64idZ+ebyZy+3Igs0CHtKfTrviz7LNn5AhRTGuRHZ5
+xw/MfdtTyeCHFEu4EYotcNEH2T3M9yQFH4wXCxxEFvkTV3+7AZ7JduUqjfgZLVU
IuwGoxxGUgdd4uJxocUsAzW8bJJe36pFS2KrzIcezOF2EtT1nDUEibxnKVO7/YfB
6/uR0q/aDRbaIwXmhEljhPfFNsn1lSWpol2bMuUCBsArmwy8jeplQTMszZ4Ml/Zu
/98GNgQ3PPXYTpwCaPfyCi9FaV/iXpEOrzcrNhgffKHQA+yhjJJjES+doNQ6vYZi
t+ctr+r0ij2D1AHxv0kecb1sX1t5OekP2j1H/qMEn/ww9amF/Cq0vkdhZeQcVqWh
DT2qsjAljBpTGqXl6pDmAglDTCGpKjIbb5iphqcWM2Oz4SOJMofpbYEqkAbN+aPH
DzLiAB5njhKMv3asS+xlmR/sVyDXyqaxCsfN2HSTHiLVKUq6SPbO+K4Pji/uRVj3
0prIdx8BSZglDqRsfZB1YyG9ngXxz8usqOfE94HLX11UICFujcGd7N9EqZMaSp7W
ADFBgx58eVkcz6KCIHQKRTub1YCsUY59E4HqxvCPmGwCPfoOmj2v4/vWU4ebJcvx
7S8cxk7wRsMfoUHPsE1DtB2ak9MmgzD6ZHU2yk77xJR8KohtsaujKA0bkRDXBqKR
D4QoalZ6sdT8JfRdGGnyKxaA/4J1BNNAsBtAh1Of9ZEM4Uc9oVGorUN1soccBTWJ
U8BH17Hfnez7tbxp7QKbrUvjCt2DqsDgqCJhevf8/L5gzoFDBeVnYXEJItqfPnxv
yl9OmmX1eQr5nuhARTCRnq4bK2FUiwKFDwvw15yr5wsa8oHn9ctaGw1ssfUtnMro
3lXHwvt9Fu1rQ2/Z9xKqaVR7WXLjlS4DvUI8qu6w3ejfAJEefNKKeE2L87iBBvKY
W/GhcFMk7UmZ21MlIFXd30aXLBLp/98tmcQ6O9J2MYUnD51bHyCW7dUuCLYd6Uf+
9NYnWbow1cHPGd6VwJiA6WgP7y7pxLmBIUOiEE7eH8Khyb/watKoOaqhNs0SD7c4
TiI8SRAb9gcdpYZx+UP3M+ZJZuLA1SQYRWXPiyEnvj6XdcQlfd/8K9ia/mFpXpPX
xKLKyKyGrxNUVkaGLb4P4ou6a8EbHQucmRmSPN4a/9ljk0X7EJ6BwenxCUijVh+C
9Ko7VMDQWMFx2Gbc7YkkkT3cQkIlHhatixO2ZzshtAXGT1AV/uBsjYA6o2l8EMCi
r/Wmh/1MDYNK6XrAdRQVc0a6Jo/6LPuK4dcQQXK5Nb8uS5OCV4gGaNtTsj6AM1FV
2GdnTx8UorU91/7FD+KsfTzkZs5Iv7eHuyNebljM4DRam3uI114G9WLCrkZLMaS5
U+6AAnUsifXczQ/15nYoTAomIucJpZ1PAqHseu6owjhdRpMEUg+gyA3fSjzZrfk4
MBB5ruEaxbj0aTqz1vhc7uFxKYFm9Ap1zbruvmzJo5VQSpiMDikSIZgaYBAr7AB7
xxOzOoj0HiS4APSG37HOXeig3OpO+KpTzjA9i5zbfP1hbGvUgwTgYecn2IyIHI4N
HX/PKBtcXs2PK56D6dt1MmVtZVpT3JEMOTQ6pIkHJiKhsvYZy6zefthOOdOM9+c5
1S+8McXUjmIYO0kKMqw+rvPkvp6rqJ/OaJeMBy179g3s6Jhj0iOkNMAv35cVcXIP
KDd+TEf5o38dv1IIgZmobosWX6AELq0ehm2cP6lsRMKGTq9iMr/oKXSBcNWNU91r
Wg5l3XrG+bAXkYURRh0p7z/I4D3+H4LoZzwliXBPQTrEPZM8pa+8sx1HnvWfc2s+
L7bNXsbAiY89wN9gVEWhrVfN9ag8SUFDi1Dqg2aw6ZXEu43LwFI3mYzv19KlVALV
tGKt6jGDA8OFFTW2t14IKVFGTTeFdZETaROGmQJ8B7b3EFkCsrHPx9u8h+9NsqA9
M32Ao1kx7U1u+J26xpM/0ymQP96QlTjXGQ9VB6wdUvfFAyQRLEhMtEwFR49nnZbs
0LK/WKhj3eJ26cWKcMV12NziJUvecNkkR5gJl13WgyLO5Kz4PmofGJm/iCqpW1PL
VoiW+fQaieqjZm1u1h5zOTdvh1OLaZem5ctMM8OYUZ/+x/nk2BpG+2PFNRVOo5Zj
7lbaMppWu7LkUs/J6C/OSTWNQnZoxrGWPrWggU/1ZmqlhWKTTZzUx8qzPAf6wSAl
/S+JWcRjgUVRe5xN5W6VhfhXISU8Gx926NWXtks6aDTHpFaxhvkL8exQib3OsXxA
91k92kxVhyzkOinFzjqUozSm+gXYBRpsFzppKlkYMHiF7KKjhrtHJ1QdDpgcnBYD
GGzlmiZp4BOexdKyTMyniJ+kODxyTnBDt43Rw9rHsYBnBemw72t+D8zHn0dP8L2H
sAMuC/kw8EfRu4BeGS7r0KLEB5u6ctXIBDDDi+wWeAtxZsEbJzTU5i76XMnfDaYR
hSSb0Pq2i+Wfx3izBjtW6RmPzby2Ry26dGlzooMEcFdvfzN60Yii7IiU7aacByTu
B0oXAUo/MyptJMEfw/J/tzuFkvPW/jxC5bmG84VWcx/Y950CjSHrME3zq51903Q0
0e9ArAGp/eYv+xZxn+nlSKZ+CH2QjGQQBPpmNsksB7E19x42Kp1saSjAhW7gBN3u
arQJABM1nLkcEFQU6aNziFd1XBqnBY6t1ZLLDxfb80iL5KmW6PCPP10slp3ppDnN
sMgffQWFj1DoBsdPJFYRYKqQ1PoUjmpU5Ld2d4JF5cljW+70kDzgOMhRRaPomm8+
JRRKLRKtoa6mDPldhNskVHXyzw2LeUsNmV41+8np457L9QW/dohTE+nTz2hxy2Te
DLgPdatCzYtfk9TLZHQ2Wz2XF+78rrKP1QedBBUlbRPlxSnTOT63w95lBXCD/Gud
TnDu5kxpn6MGliPmyv1B/5+jVTOGechHYEkhQbGzmfGoz4k9XVpU62FCel9u/TAS
rwRprLOApvD6kwGT17Bq1d8qGkHyg3c2wgWmJE6Z2ec79Nu41ICBnz5uPW2nw1+a
sy7Vp1850hVCSRH/7Gce1qD9QqyqyU0oLqkRFWl0lRTBujkCfhcBG07hb5Myorxf
POtxYN63HdXd/kfPoRVwryfYqbXhTBYYwwcmMHyjgUfZAGaCS2vEOoXjU8yZ9XM2
wBWsM9D7k37+JDafcneowAVYAqRMX3mnfOoymYX1aJAfcCT+NiNo75hJcyzEB8R0
WMiYHmf67J0K0ncb9I1mFEGLVqdiB5cU8B3PdQw/TcCHczWuYPFhOwYdPUlGgOGt
dUq6L907VSpqA2RutswgbySMxMZ4LBqsEIhpJLj8H/SXpuWvdJRtm18wteCKFIpT
UmdlBkdq8C6azXHR0uvGz1xDZmmseK49Xe0DzRIIpe8zEQw6/fgIGzPOTQMnTnYb
wf24GMDWH5MprUH7B1eTd2uvQm9qTJ2DKU2bhnSR4fnG5o//AxWfenIrqeNGKRk7
/A9cCHyycwzIF0K+moe20ExcBUJFjHG0sy9T+hjzICysEzFl4VpPORJvzElIMr9D
ch8wfDedcJFVzB4+l+6VOnA8I2uANLzSoIAaFMXpJbipmDn1BxTkO41SsF100oX5
DbrwLIlIZbLRrhVOXG9Vix2bpXce8e4xpz6LcmshyYoxobHYd1km00JAv1HzfrvK
ftZTo07WPahTi0wHseM2x6bQEoZ2hlnj+XUHuaIO4q6AZVbnSCpZBht/xp+uFlEx
IZ1nw+lWNbKuuUoVsxTHB3TBQQo842vdZRLK+dLV+lBY3LNTMEtgqZsb7KxDh1C7
md5vaHf+W+YETjZFNjZBKJbaeFWRjsYax7I5c1QMFQFfKrv6TpiY+BECZrJ8uJz3
bXh914DIr+yDs0TQ65r+n5sQ9CHnu9eT9yHgI02d9Bacp11kX4/mQ5BD0VRypZO9
ziH6u865BROMlgzvyFuw7IesioHNEpjur50DFOqEkcbMWGzCKO1odWucqXpOv7Tg
AZNZzcMeeB+YLTkyhbou5nNKEwepL2Vwvx1N4T8Fqwd3ZpH6Y7HbC9cjwWAM6lmo
b0lbg31+gmpJ5ddRpv85E8MKPtH6S2SjgWhDUrIqJ0bgSSYOg1chhLoQ2utPxFWX
isk+4P8R0yjhgLznHlqPYy/iS6y6dXZ0e/inKR+b2iPEmgXwG65OouE69PcyNzb5
vuWcsrc/bsikn2hN0Vp2bxNcz/gYVQP+INwBjJSx6n9KQ/efB0NfeKkLjeABnJL/
h9AG5yQRHKJZlxNqznoi0o7e2vSRlERsMVlkZX44T3Rg44jtTNr34DvmUGkKNXkh
gMPbuVYkA0hCiV9M4Byd/zWMVy7ZP3wSWFrXKbbnjLMOHp+IfzXUAdiYDvDIsbq5
NsDOdFMG1cgK/qwEPUdXi5LVrgwtG0cP3Apb16w5Z14kAjvWC4R7TTHyWdYeiIn8
iQSDDBMcgxQ8sIvj2uIAy+KzYT/pOes43XWk7WWpXhI8svq3/9rl2XZakKAwtAnw
VQ+RpkQWs7Ej3zk25EJ/6xrMYHB5ut+aKzduW5ZKUvDybz8WJcKRIxYITq9EUq41
E6ce8RecFds/2Cs1D8xWaq8ycb7UAcI+JxyQ5DCatfr/3uMucgK33RBnsp5pIm4N
oL3qa5hVmVEDZlQgOQkKto87tk8hvpOj5tzqtZZxUmBkNR1GwNpqppjrWL8x0tAb
hTVaZG8eZuVoYQ8zDhodlBkdbRKTMpl48gNtsHSeHMVs+JR4oJAHUgdOFs2fOjFf
PFLyOvnXKeGYEiXqZuCPJZVJA23+yQWZW8e1rxWVrdTJByJz0tVdKyy4ipFVH6Wg
ICWLyPtDxg9epNoXe10hjybusyMOzPzYkSlXstdo4d39HOGbC5QQ+c6YM/lWPiZg
w/JMsPi8i73GycFDRrf0J+EL2TwqEs100GF01IWv2tzUrcY5SSaQGHIJ609CB89H
kPAQ6akRhlR4DYwi7tn1dv6mZk7s36RCarXqqP19uSFCclcyM8y9+TY+1vCrQG4o
3UmI47DkAf8Q6h+0C3/6AmUL2hmy38IPulnV0pKQNRNQ0HZN0aE+TVFWoVn0sejZ
0oOEjUab9+JhnowuAf1xwD7BJShQpR+D8OLzgDQexf267T3Pz0P7frSbRoPCwI2M
u9uCTtVMSLGKW1ROrhFSi3RiATDlohaSw5UtdhY+fIHAQX5ZsNDYS2r9dW3IVRBH
hkFHIsVqm2yl34F1nOhNqkfl+fd5nTPqO720ZA4SttpVynpZ9e1ozgJrdHSbxr6U
jMI/WbL9XcZndoDI1uWDdRFzrH4yW9fh5CM3/bA8B4DXjndts8+9Xge1+IJjUG2y
4U38N+UL9jzRWTG/6gPsi8fxCiERuXkPFGU7Hxr0KolO7qYAjvbdY+LmbhwshJaZ
J2bss0ebuVyUEkY8txDZjITpjaFxj7hRMGoTN039Q92W3DadwfXcs+aYA4k/NPZu
9zXaSEGuAvw7PuCn9cPpt7GmgIXlALsqEGh6c3vCkii2qvktSQ3WDYHdSusEntwu
vZhFggpgDDRHN4tKphdwwbtog9Q8kN+Q9l3dzbvtU8ZczLuGFRyAW3JtHyu5bi3q
9lffrhhu/9AB+CH76wbohGP3SQCRO3+Wwa4XL2zrTWJOd0B5jsLp0a3Tn0U8vhlz
aMH6DGvPJhqvo4I0zJ1o5/v5Nt1G0SttAn4ByjQpPSaIa2RPAAfyVCBIN6T7APV9
8rVZy8yMv5U8Hr50bacPnHSa7Nw00CyoN/MfuEehz13ev40Boii+iYsPpGxNC0X0
jkhwqGEu9g1X0stq3nIa0lNOv5Qmw6wKP+SO01Nqy5AYzB3Z10GMcvhVfHLqYsih
t1bltANWuTeRV9LUSfqiPWkH4beEQq9SyeS6GoS8xz/zoCzh+LqdBOC//R4zG6X5
SM4SeFBwbCcUOWgQsrJZ4d10B4ungt8S404Dhf+wMUfMC35Qr5opMg8m2RwHV/Du
cn0sRwFnwhfUdGKagerG4hiqfkNhkrk/qjMo0LyQRnhSeP5z6G0EcCUdMwDYcMJy
3+XwR58+r7TXYNzDC0UExa7/Cg5yB3VQfHfoJdwSaXKJDGZmGuKaZE4HpFm760h2
cLiKC+Ty7JxdqF8bCn3pkFdteE8NHObNBe+rJcVyeG0qUhsDNZ+Q+TGL2sFPVXt3
92ogSPQIL5K+isfwuNvy0kvqIO7QyPZOveD3FIL9oSz15kHowZ4r8juR4Eg+WH9z
HJar95Euh7WRJFq2Ef8fh8PRk2ffnSlLjC4QvsTAiW0I82SX2/7IZR1J+Mfnzczo
agos1+u3IV5ix9tTkJe9sLUkAI68UlV+Bmfue1kwjEYx2MxVTjuTHtTXKOk8+YXI
kQ2YwfOHnMWLbjsl05z9FbsT8n/7pFAtxZYTBvQ796B2gBFQniaBK1Z2XaJppcoA
GsWlwS53mPnJMwBAwavPIgxAkX0nTIp5ztByakxDWvF/vpJCZ6CqlmmKHRsP6ML5
5H6pErnYe4/KF7wKHUdYiu3K126QlK0lVjI6V0txciM3GVEor5+biQRM6zEOu13J
ffk7RTJ7DKUyhDHSkz3PzXIVArjz79vA3CPitAgk11mryzv8wFgQlfNptofRrOlY
MZtt4h+5KG9cJeQpWX+BQn63yEfcCLKsk+zNG2K3VxT3NXDq3353GpIToVI3GetW
QAGRTQzi4r618BEe8gYYWZO0EdBSxLj1UE7WHehQl3rB8jDqPDjm38KGgjX30Gir
MMpOyAkIc0p8+0VPOulwQyUSfzt53FhP61cJlwFQbDr0CYL/iF/az9PK/BTNU7VW
r5s265fnV/MZNcmbwYejkS73cWM4iaaaL4HA9Q53OYxz3ii1bzYAy7uAeB/DKAj7
J46ClR8OgZH9c96LJCmNt2wZyq/9dHfglaefmf7Jt/nu4iqyDNft46HCu1BskDkh
j5D/l75MuPM3QEnPv17bqXJhTX0Ok6lN6o2kLtVqgk6TRA2Vi4+M3U61634oWNZ/
fbYXXeZ53YEjkeV32pq7YeRxpfbdS4rxQE/qbGkRq33tf3wF5iwSXV+IsMFtkwEo
25eMuFevX81Sdo+6aTgeLjy/1wo/nMF9X47Pd1kUbXGKfLKg0+cjuY6LO38MqNz8
bIHW1PIH6g4I83mPYlZuSnsWrrb1HAwIwT57a+E1gRmMwLFjzhAsGqULcP0ofVQ9
g58LB5jGw6sFtFqAGmvParf4ojgArIApy2ypFlKbBwGGU99kZSZuXy/6Tc37QNqN
zZpDTgkG5YrDScQDy79CPIcVa0obEo6mrQu+UxqpXhrjPfzqNmse+al7ZOV2Y4qg
VmNET1YQu7y241+QwmhJACW7tEeAqHskW1RlJ8hGenLLN8kxb6OjMGDEi7+zxYoX
F3UfkaqebgCollrIzRj5DGprX1PEKI14DwR7x5O3dQekOQtujKac0wJS5MP3In+X
n0WXv3HrFigy+yc7H9NSXC+LCw+sGhXm7K+3d7rhNqvvtVgquKy+tLQZf2gmz2fe
yu4fg/f9mPspwE4mh4yulbm39UY3/3o98pZw8CdPqfdNK3ig7NsL90xpTUUgjJgQ
tG62TA7yO+vVjfIKXO+BUfaZZFSKhLf1kvGRZSYFQADNn9xOU0QyvWj9qtw96TYL
jV6Gw2CVmpyeTPCw3+NUv82e/WuRtRDoha0EBTyrAUPyFFSvT/kRl2CqzJkI+VIO
zZFfwlVoHXIT79VjRRqwhanQLCf0UFS/xy8RY9Vti7oqPjyAcf/ZvzRK6w37dgfx
kQ7oOqeiKRNRDC60uuy0cvYAwvLrsMKcloJHPzrf/4OexZB/ymsJNbWX47uNXQCg
/ZGQe8fAC9wi7DmMclvWbWtkTYlmeCc+yBgmQoGNhNy/XEgFnBvBQY7fzvBHUypn
WXCqmaMKJSsBIIdsrZcKUzm3A2VitqlTx9ulJURN0yDdr6Pvg8IlZgYW2/i1g1Zd
reb57wcry65ZrRQvZBeQ94wPbEmnSR8c23/PvpehU9KwE3rgZbQQkJNy1nsZhQ32
lvv+xn9MKZXGQw1YklTrb5yk4IFF2mym2c7jq/LTMzSMdBRJM1jxzuKEl+6wdkl1
JgpLnCvNfl5U4acXf3Jw/yFTL3s3zuKIsb94WV2p67t70ErIwH2lM+bFlYHv2leD
bpx/uDBI7PR5SVi8V3opmWzEbgPTD5q6YZO9pdd2/1fDqQLeCMGYhjoGttGS6s5j
ZjL+DbheV+QX1Bv9FAh4KrAwNofLxQu1+ZJbmZdF1ALKZsLAQTxXmtroO3dvFMM/
Q8P1ap7Q/fvKSRAbwSUvXtMYu7nsPbjT9KjEay4b78YEm5aSk90SIynFiyOVuOEp
t52D/4Aw6itAkqID327Rc9mORXMcKKDwj9eHILAikOLBGXBluOpVVpntyDHIZntl
tPTq62mrxvIXz45/TnAVa25SNX30mg5b6AFaiB06kRu2djf/dYC7o5WV05KFzXhU
ksErj80zQzdEPPFsaGi8Mz/ojqxrDa0BsexCkAKlLq+E77105yYdkrtp7n2kigun
1ToAt10d/jiR4mbM2tK6mC1WouAlvg14IpIlADlM2VJ9RO8QViDR1PSZ3gE2ch+c
5VmsQTxPuI2uG/TSJQx3280dti51sVSVSnT3IjYfNG0KBv7wI9pp1Eq+/wurwg4z
LC3XUo0CaQ+XXYnlBGzF47heL/MDkMZ3RwqhRNAbW1f1A2uZ6Fn0ivgiln5RfwJJ
Rz2PzfmSF2sJ6r1hcXohiuLn2Grb53lelG3lMDFb19cYQy4E4JU6JPoaPYZcT9Iy
R1xj3q7xUKbw6iAGWq+PoGu/1mZlokr6YKFiKl4DSkLFk4sMshmd6JODbJyG9hax
noWdXjufobTUZp2pWSoby4+7724+iXmNgBTiV0yySOktUGXUV0aWhFyKLc5TuisU
aKBZcLr8ET32FwY0JvyJdQgfsNPIIQ8A3A2o2lcbDq7/RkVvWczlh/d12udSHRRx
tK4bY9U7FemE/CeC+B1Ndb3MyozB4teObvutEJF9sHWMDDWXzurxTlMK2h0zmqbO
CrsdTQUUhvHo0zXhOPyBVpQ2Ztz3YjeASuV2VxYftK1W3G35KBAKdhgCH+R6E1XP
1Vu4UAjtRcJpwx+FJp9/swEQzSegnL2HgwymUIV3FlyEdeAobCF7ZafnyERqqgUl
qMZhTYOybAEumtBx9Kx25fd5FydJbW6ethyz0GOqikRMLmDWGRbUKocfqOGy42LZ
TIE3gaX2xfu1Vq66t6sEFlCSwi7dIwkMCbLNMugaTwKbYRT7HXXXaFjFXPAyuJBM
TXThE9JCAsygPLvPusRqqObQZ+mwuH4fet3D4eSA1kVOQRRGJ5nve5F5I3dMJT5q
B29O6QXq4nbXncCjIBqmnxid4bV5p7eLxajUM4smAtE6mgHWFbPJffCicjM/GIRQ
apBvBPZ33jcVWGoQbJJ1VPolThjqfpHBCfhznZVI8o2exs6JmL0s7dFeR3efnDhQ
LYd+ROhNZgjoZjyS1m/lSo6tt6gm9IiUCgdQAOQHdkwzherIMw6py9KEK5+SZ5cp
sGw6bENjFshiazBvawfv69LsJgjUPev295nNOCtON8PKt2FcycCe1UiXMiPjZDIm
HvBJcwKTCANxP/Xl6LAgSLAoDxHtPA61fOnVFD6UYc6HSGqy5uUrf6KEuSQX7fEj
CEFU0YzFQOsD3WqSmtPALbuxqg2XS5gqPGmYnZ5E3gRniIUou5KW5MGSXj8QUYkj
JrlWVeQVL6BNm3WZps/zju0zp+7TsjEX+qk3Fa+B7pNcxZIuOz8oOm9IMVqOpECH
XC38fRg89iWdumTaBsXCFMZXB1HYx5FPWmGdK0PuRoWA7/c9h0AebOn8immqTrpe
4+XjMwYBu7QNdbKn7/3x0SaxbRJzA2uSnhoNs2crPtLw6ch29h6qRtVOlT83+qw/
CBS0tA5K3bNlrQjTiI/wnsK2HTR1eM0/5GuTro201aydR4FyY04KX1KwF/X7UyrB
z+moHI8r9b0nr6N1RGR39r4pba3guBr4YrdJTNBCXx/f+twtt6Qaw0TNW8siPw6Z
TGxrwCovN5/9rGXMy4UAArsKO5btNlKdV8Tl0vYThv4KzVajKSGuvQMasoOmPR/8
B3R2VRTrqfuhrZJtsUqxa9zUHDYoL1GU5zqPhjKlkRYp9L6QBU6DEDW7yWKe6Z1o
V6kNZpFmnxC+IdG1ppv3mQCavcSs14RxhQfW0x7o/X8d25h18fWmR2vw5ic3lyxM
4aLJQ6flKjoTMnVEroIWB02bDvh8ny3J2yvn9WByse5fGLM37/uNh08lRkdEzya/
ADt4L6BvOfK5qGxr1IOdbNLL2WehuOXnwLIorroXujoj4zlagMAPn8uo3ERbbtG3
DRUUHWkLuRTblNxeV/0B4GTZ++8fJVmJQ5nRU2QTd2TB0oOM30n/fr+XRPm3vfOB
RGfiluabtjnrML6c/k4J3kr0UT/ime15Y2A8FFSBQcPn2MKi4KGvAr8qoDI+Bb6e
msJ5s3MPpr3M2IPnmIGh3XEWwexkyCGsA321W+h+HGpIpNXalOsE9nHZuMJQ99SQ
N70i5lPpf6P2aWT9NXMqBlSqdJ9Uee3O3kBO03pFTxMdLboHWmzZ0j0I3XllnwJM
IrtpfkwsPjbW8LvG258RPu0x9LsjSzTOQ16CYWTTlAz3Yv+XzNM/31LTIDeKetGJ
/ef+Ox9tzQmwcPgqV38PlMxqPMO6ewJksmpO6v59zfPlfkLfwbSt6k5G0N7vzxRb
KNJMquuigBt4jLCb65LbVj06KZfahPiUtHago7DQ8PzV1ydkmSN+q8o3amqsN+pu
bW96qC0M/dOD6UZf/P1qVUbiH56h5p7gFF8T17BmyJsMAIU/j6vfndE+NOiCJEUG
1UFUABG93hz9lZU4i7MOhT+QeH+adkUWwVPpo5pVGVK3p0KPx6+LNZfTusti3r6J
oHCO2a2iN9fWQXWbib9GSpq9nSFMmrFjwW9nKp9B3fFDDZBgGraOImo2Koc6Jlk8
RjATqDZ2nDePBG1/olUJm7oEgV1EE7b9SWucMQlME0YE9mEG+YXCPC2vkvPAXczd
wURXCtzsFUjYmzYechnFW81Vx7ekoZjhS0RtdSMGI1uiCVYUzMhfrxr3O8ZNmjxJ
QamFlg2c6Q15URkQ2aIfvnJCw1LrJYM/WJHDOavk4MuLOtT7MzyI3tnjDzvNexkd
khQEu3l9yFtPmvMner+K0KhyiWekXIhUeCTS0z1plcUORxVgybVda3GbHNupe9IW
Kqce9CRGBNWiidQUggJMsZ4wLT/kg40cNCTxLPZmcWIvwMBqVRM4oU8/XZbohuym
8XdhXSwKRJSPnXtJhLxYJW3Yxmw7wCXSOw1Gc/mlvga5UopFkEtuWwqbmI4xVbMi
BgX5LWTBVUpbWYIYPLxVGMsTrf0qcF0lT1xxUOww7+1mbrDd02fxCwdwurVe/sAG
c+jgYpkZLV1h8n5evNN8APxqP14YUWf+CmlP/i4qbkHHTNCcVtxqsVOZ8rleWd80
G2r2XbiqHCV4zJc+ArWRqeNRrRHspUXpX5bz4IkPC/+qW8rE5dsM3NyuGBjKYF+q
UJ9m5WvdyO+g1nujmcBTyVTCZlT2OirRJ0lXKPhjpkkVIElLcIIwwu23eWHSQflp
3Bq/z77bhCbp96gbJ9XYbyNpCpo2zLt5QwhOuB17R7gp7AnziOFsty2HVRE/PhUC
uMMmPU64+mXJUKjJNfpCif8Ufw9HOAiz+J8QhpnfRWYWX2Yn1+VUd+3IG3eaJOI6
Z71lwb4/uO6MhIMf2xShW58DX2TlsHGXJvy6DDQo8lqpnIEquA9jNs565KhDvUoa
mxIljSt4rDx5YEwe7nTEoQVljLul4oWvFT/JCoCeeIOVBqf8XThs8Gr/sB7Itrb7
mV5FxjFHyygEG4pCOaJmq8EBgJ2LExeVYV8G91s35kpSm5X1PJGWjxL0O/JGfKA/
mpGsknf9gEKZOMyEV4MRsQQwKleA0p5RyCqTTtlEi4k7buChk8zc2nbh3UCruOZN
c6HldAYyfWxI4homFLLK2kPhdbOlsSLWE3bL4vZsMfPkYLzuaLs6CmPVzbI6XMUI
K7+EVmqdHKNaqvxumh1RzWDNS48DXe+BDEymHe7JGS2WbbcUJ/oVC8i139yLMzck
WlGBrA12uTbxWIoz6Ik3pKRyu5e0+6z9f+Uwtzo8p5HDWHwTR6AAzwFMIFUnCaKD
XTMP7ue49U4JrjpKjPIR5agIVQFBxoI1UuKA/3LnqRGk8tihBGpaZBI1GTXNGXXF
Z3E2DKgD4Hk2uCnJG+oPr260QfFqiUZOEXMvkF/B9K7h5iFZbX6LhCGjo1Gyoq0a
8V0JyUE38c2cllDhPtdVNiQoaggWSc8tdR+w40rYSJ8CMZzSsmICVBla4iDpKPux
qLa84WyYQBALKJt6urr0czUIyaF2ULiC+Pl6H/MhAYPtoPEo6ZIO/tO7WoWNTZE0
XvGlxA5tf7tYbRO3KZEnjYx8s3RLLamr1QTjsXUZ9WGJNZ5PYKx4KuzYf0Zw6MWd
uxWUzUANYeo1Q3EXLOAvBTu38EQPrXj/x9b0/mIhBX/XpOnEd8ayiezHUpJ9hIJX
UJVaO0YZCbf6ajxmu2Pu0hD85VVLNEp0nPjyS3Akfn0e67rLDmS4ObpX6KJiW0Nc
M9a+n0eRZd5E/GM7Ha0fuK8ieAxJ+IKT8OHPulWiqyoSVE+dmm8rX5mGM8CnjlCs
dCkwYINTz9hmrZaGEJ1QdvtldNtdSiAGJDje2dxkmWerwJMBgFnUnCiZXj6Jm5u+
GapVpw38Lt2dEBpt5WQqLfQWFEAeIC51QouQ5hh+nR4APdbG/bXQ0kdBw2VZOf/T
oMylbvr2lhP7lXYHqkux42YSXmwD/Xa8bIKiBsSkNs3bwQGdwrqBSiKRM73Hoblq
zG+/RmRKms7CvPYC0w3/rkv0AvKKOA0AEGvKx9bot1d71pR8e/AwJtY7L/Juuz+y
QtaGqgGjL/VUSkJUFkEMD2fnQ0+JpAy61DwV20lUQitfNkp/xqOgzD+ueuei7cDD
HSSv92AMdJCmvUDwGijEqpo9j0madOz8feYjVIN+8fpOgnKoit7UZi0L/+YmC2qD
qjI3IAJdceyz3AD5JFGs4x7VpxpCGA/zT9xOYIC3Edr/aKVBctKGQ/FKVd7WjDYW
c1PvSnyaqq4cW1lXZYQRvdo53QiG7TwWsffniIYrdguaqrV4ZlE2mYnGBDQS/OkH
OqDFqt63edROwZ89e4hycmU8zh7MzQtMjq503GGCH2IlT6kmDTH8Byp9HZ3yy5S7
jc8rmUtomywo0rSLBzTC6KVlPAtb8BKAdQhMRr2+Hv5MsFibA2Y3Rod66BXBfVSn
LOiRndSMrueiiSuGHD3QsJIcDLQTJACPAEAH8J6M16spCruSvUHYWX/aTd4HDF8+
6a7gYLxN6Gc43xXoOnNxyBt3FEAOTwJ5zMaiKeAg3SiZ7VwkiDdcldgMPO7NQ0G5
OI4rk0K8xyXAgAZgmQmRx4E1A3iNr6u+ItfOSsprb5u9/2Z6ud80TgEPreNqGbd4
PhQMnnLWo6JPQGefNpH4Ak4DCxRs+e/SU0tpaWicXPXB6bTfs5Pcq9gxVm2C8E6q
Itx8NY8qZ7O8TLhKiRNrfplkRqYQIJwZrKdAv7fU2gA3bXYWMRkHqg6ZEp6Wn0SW
TEIutDQwC1W+KkWl5p5C1qbRK/ZKfaLiDfljjeJqsULkImT78GZW5i4VAaS72nX8
jCzJOEsATDmiGUvl6k0vn9MuBuD4P9+csMHZklmOkL9808/QkeYTj0PnGMj/73TY
6VmIVy7Zvur0zOi3RhVp3bQ5XIxJft6rP2Y0KLFL+9WyVBSn8jjUy+LOlXytsAVM
TRMV0DMjqn7dRMD57modvSwTZj1+18WpwQjFDRVkeqpgUWf8ZR6Qejw+aBUztU6Y
QWNfnvbwUsRSUJIC0Gnf5952xVYET2a43HZfwqsbA312FcsQ1H/WjD/XXzDgiuK8
pY//VyBS+1cV+x2Vwjegi8ZDtv3CDXWhUF3CnzfrArYn6YiPiU/fwEesFjcV3svk
cqLawfFn/skmsvP+g8G6GTZkFpwaop2dstupO4xLULjEfL04o6wdOiyA1xSLaGFn
+DXk9ucJBn8y97z6KEFfmgLvXAqnUVyBgxNDCSbkAVM15G1nC01tXrUJOCpd6pYg
0AIWEQnmiAXXI6KD+B0vJ3m9exNb8nTZ6FIPo2JIcXqNopSxXJQaz1sv1fqXgXzp
kIFQ3LaA0UIgDrE+GrfRQ1x5JWTHHsg03Bi6fymmThACod26dVaeN7F/NvwJDRaX
HbCsB245YX3k8L/PEFYJzj+TiFytCuHNuHaP03k8G3jOC83GPgzKFrRwFZ9tBVkJ
jQBVIEUGzAnaUxSNL/8XHvukPzjVF6ZNBCIvfNLLxjCRHt5HCUuRfPBzMQoBHDHJ
bsDNv3oz/b1wofv7BuJEH09fSRFZz4HcaqSCloeMUiyqka5y5BMncadqwaupAW7d
wkggwCVL2opfQNLEBuX0mm8pI0hS4m3rOjKxCITp9EIWH7CbvSGj2qeYM55r2t1e
4SA6YQIXqNGLd9h64j6MAg3AWP09Jve0KCc3CXitHlb4/Rn/i6fO+rp4BVnr7DtP
w3gJeLhtTenvp0RpRw7ISzVcji7aPxFUTTV/S7LIIR9V5/RCKhrQNLYaRwhoo+T9
0UiAb+/1KKwGohvCMXaB83WKkrdwefK9sosSLJFLqv6ef2/R5OOnorRcgJqWRybm
lBhXnu3ecSnYiW5gzWo4RpxVbcu4XmXefH+nfwLge5BwjbnxvS5dLcPZPxPZHOrd
TO1ZG6MkEShyEjVrddvb7wCMkSWVSEl9V6QKR71LMLmZBeWlWngGbRmnsbNiIWnC
MRN3ydDKhDfSuQ93fdcacFt9acNk1mStVJRCnJlv3hS/JQTFvQW+DiHJO66x27lq
7fKVdDdq/4Nf0Jf4+bg7iwWE3vEA8ci1OcfBCyuVPv5N08MTjCUoKHzgtLGuQAQl
xxtyh1RDlSub77GwGE6SKhb9wtHn40DKqN5O+5Vnkav4Xt1xRIvcwyHStFPk2QI/
4ysp1cxsUIwSSZlx4OHk6TuyO6tsUQCxi4UUUU5wXXuYmXd7nhiGxLXJ/GbiJpzi
qO00XLoXpfR6VwCzM1sSh24sjXz7/3i2uKZMzSixgNi9e2a5nvCxiRIlOBXOeosA
moulSjqWHf2Bdv8fkMT/LFMiUPaXSYDVHIla6y65p9OZB6KjKF59gWu/u1YjB/5b
1vmQd51qmzNAfXGDSDYEk1VVffv0ku4WpXy156ZKfg/SowgmPOft2ALKdCGB/iXq
6Yk1XBbsnLhlRYxx/ShC81FFZPTCpZmMpvh1qk/RxfGly9YmBh/t0OftQJZMPaxj
MaG+LXe6IKEOli3Fln0bOR+40NVq9HeDZjy3R4n+9MgEt6ZClV4Mxc0heEv1D2SD
qjY2vPXRmhCTXjPqV6GPUT71J0nYK9zn589umDkMQksGZxSVjl517OZbs+DzmvIg
t7TYWHrz3DarZnAJtloWic07Ju80qGUrfymAp+5F8yrwHI+nQ81TOZJn166BgEez
L0Xrpyt6Ak6of3tFkNJbBeeJt/Da/Up/1luoNUgZNr9m4MXQa/VGtsFYqj6gBf9e
5KwYqWWYGwXkX5jWOPaiY6mbdMGXxsiPMXP/w2kjS8FtEP1Z1M9CTgLpNt917HKN
h2be4hflPbtp9Q0XM5dt61QJQghbd3IVrd6l9xRAPYhePJTAxqrsNBki0C1lls/t
NGJ0Jgfu+9vXsPTb+ZAsLTS1RP/1b/Ya52YcsTQPWLi7ld7RagMS6oV94VyN9y5l
cxChZmfn5iAOsZp+mvBxQ6zvvck0e8o445wrl/nyaS936jgMaU4bDnciRSIerWQJ
7bzyPQDusSgIbamqi3ggxqzcM6K60GMgU5WlFJC4ejUE4gokyP9zW75uGkSn9p5a
Z7NHFePpu/CZI1KBSwWF3OJbtYgvhbroMCR+FR1TCmTbVwa2wT3hjiZxZ3PNtgS6
qyu/NckyMi1ZEp5bAseaCAWuiZXqlSWWOGaC0I+iygiElAL5sg5xoz31b+nKWHn2
bXWGrIgYqvToTReQ0umGUU/KGYChcuwqIrlsLDyrk1MtZKZKpuPjdp16HgCaXorC
5OgQq8YMckIkBaok1euVfg7p7uKeXklfODZWEBU+VjG1BPX2aM07kATAuZBi7ZVg
D4kxjZG1O5wPq6BgMWuKqa+6NOzR+N8nsFfI7dSWfiXQOgRWjRaTMgXQO1O01vSr
+ibgyfL97hMsEKmhABGKegReo33azz7IWGR0/+UjNKt+QIMQTzRPWLr9dvORPU4w
1Y8BD1vtJaoIEU6l53YuSJtHh7mFAv2h3VEnxjuLWegSVv1NFVDwynFmmdgMcCwI
TPpGhdKS9T1X4H09LkYSCt27I1fRdXtLInOsGfXPKCbHCTfsd2+DAHwsYWnAqHUM
weI1YoWz2wrMy9wS2doMxn5veLWxrkxRK9m4slj0y9pjvQ377oTj644ObFSm5tUr
JvDbsvML43niaOfxfYB3QyCU9BUskvdunXz76h6yMpsDpZGXePFdsTMV0+Mv3zHX
91lDdwQ6MLltu6ISM95M+YnO010u/PcrUEYqBZSBbr5SFGhsCZxler8H99U7NqFv
WrFeDWYZ6Au4uR4aX6HI4H6uR3FMIgbkV75jr0C8FjHJH9k3gli4ERKMS+r44zJy
KIu3r3GAAWTNxeRwFmGTa1MndCXWa99JpOr7afpjAUb1y72Fb/FTBt65Qoeott/+
Ssb5tumwEfcVfTXcQfxnTLVcNXXXBD5qOg6fO4y1rrn4lk47xIUPk+Eknx6ia5FV
eMhr00q/q/FEoFej+NvIDkksy4DN3brZBuoKr+h6y04oIpWcJ8ZwjA+ulk0LYbaB
1xJv2xhBsiE7SJUWR4ZODoXnR/oeGQxgC6TXpGcmMdZb7u9e8TDMk6PJlpQc9yoF
5CdOFvuuFE7YqChlkTSCHS5DGoyXGk/prSwcrR/nKKVj8O4w0CK4t9wYttu0JtOf
J7/eroS+wEy0aqDI6PuQi4DzrzxQ+LqUEfWG9H21j5PDVeOmfUjMpqVtMDOoksPE
qqk4Lnnu1WT52lU/W0WOp0OQ1cdBae9QqknDO2hOHeywEkiUflevyjZTjdSq9H6O
5jHhaqq6MMgoz3uph9NNHAhJ5dsrv6ZwAeSO3P5rZowPFALi81O98XcC7jQ4GZjZ
kFJA7mIO4r/mi48yCPlYO8AUXh1ULuKL/pgmhST3IV7cK6X35FT75rXUwa0dyh8h
90mFKGWZep5ytVUF/FAkQK1a61O7IEldptuCsFTjgQm7ImAPfDj2maMI7Lkniyi8
8KbuYz2XqVzIo7rcPbBCcSfk3HYteGqJs61A41Eb9ToXEVTOew+rtgl7qJLoCaRy
Q8Urdv1m5mN3CLNKhzVtauc8QtS58ihLumoWqMvQ3pzjOG9XELQycSSG+zh+W5nD
LKNRIMpqM+u2on/vfedGuid70c7ITJuAK3Oc6QtLjuuvdqYIXbuBhJaruOflQe6D
I3wBtj+f+W79Bejd6vDXcBt0WoCqeHzNrua7G6Xdt6qodl78vjpMqPmcaUf0bpNa
DpQWwHXMJln7lxCGU4yIBbuWNmPmLksyG1FxRuN7NWhVx98wvhRN6Ut6IxwgJV09
NyosiajGLjgdLUJ5BIQqD76Rq3QrDsGf+xU3yds6Vq7/0StfBDDrY7DeYSJRMTDo
vHX56sJqcWIFlC4fULKAMDAX79PM3xmctbyQKWjgV2LeyubvisDfPsyKJXcUzAua
X9TEclCcwhjPEJhgMi2Qg2BwV5/XJkBndG0FdESGoBxJlpeSUxiifNemmk7lnqjx
zIckKB2ip+Ku4BuNN3FoT/Dnck72ZtLVTs30/XMj/0bwzHqT/GcufzziY/pSzibY
uyccugpKuvcFu/KoMlKiz8YggIEVJ35A/vyM5UsvxCBmpTiPX6GvDLr8wRXRG/eM
FPIELQtfgvwR+xSvz4X8WsDWx1vQWeOnejTgTfZbekjX+Y+CErY4MUW4c73am/sh
lFVHesFzxhqKujkvhXopYAYRyeobMTeLNfiSArOOGU0aJQA1+l1y432LMsOVaxFO
mlcnnJc/WgDHxM8V1qXRNj04U96uhtCqKyLreSG1fZFhwVXQCOAfI3WyMKPnf8Br
eLcbFeheOsd0naTOSsjB8MyHBtHEqQPkBd9h3mFn9NsLN5MzTtIpOTAyuK7v0kB0
elQLZlfPdIDfCdxsvgKHvK6Vq8TClWAQErOvttTQ8yDYJKgT6AxPcjU5OH8/AZDz
T6yGmeS8Q1h3HYH+BdC3ZupQPlPJdgd482Ofbzru84JiGj/jNcAM5xf5T3JoZYVR
yI9fWnVh3hy1KoEROJHwyD88aA8EjXhVuEOtvmnlsHd+Jzs2VTWdZsjv6N6cjLnR
Ri+zDbHkFp4+ji2armOuVA0lKCPK3tn0swUo1/a3gwMAVkKnxq/eQvZM3VEb11qt
TtE2CDt3lYfaKw0cXN20+9t5k/A3Fe6XgcEfpC3lzPOFJA+djGLi9M1U/YsoW/HC
ud26rtSFBtDxJWA/xJIxm/fbeafuy8ipLpZwKbBO3fwAgv8uGEulktFDmGncEZv5
ocUqEG8pubdzHtn5Yw0FMQ9bpS1edHa+vHHqkCM/KIFdNiqZM+PQI/TkVnHDQqQq
0k9n+obRBlaGdU/hL7mKeRZ0s2VtTyXev9Jh4J/BILnH1gm50f/ORPS/D1KKb9+8
6RWyqUbTu7mbTbUyfV41W4DU8LqPYZRxhibMT//M+b/y/CTXT3e9ZSH6Kj57EATF
TjrUILT6XDvWxdn11T78loKhZnqn+hy2x821+oUPbo0IxP1GjgwiTiFhzF071Sdr
m3JPkQ7Lq3gMmNY8EqKQvNNoz2hNNERN506fbRDe44i0mDCCJBV5MDRqaEIydkOf
tlNKrDSwmPHtcK1QCepl8WeqKdjmTc1n7XHpDRzEOrbtAr+Xh6GJPKe8JDQ3r0oI
BiXvIItCxB+prmaRU8sTfccxiBUTQ6O/DsFlCtvNrJKurq8PaDx/lt6TzhShIE/Q
OpwgjJyf6d95jll8xED58Glrkd/aYRm6qf4AGV/K5nGZkZJopIovtSpFJuZvblPe
yGj5fTV/Dme+Z3T+HRg7GcnkEji5aNgzw5xscoJFDGfiRFS45Z/OK0lqCR+WUbob
cy/jYWgOYtZhRHrmZ+9+fmnJvbeMvDKUoCa73hXq9keWrcwBU6RPt7ciW/6/ETI5
9yDpXBJPj+n2KUfhZkJowmkUQpaItJcz2US3qpY56bZsGtrA+9UdUCtpG7TzQTUW
fL3v/iwTDiqTKb4uw9v9wFYz9OWK4YC6XvhDjoXPDB3Jl0uz7uj3CCyoZlu8JI/Z
2OJNFF37SMt8Os2y1/Z9rEEvyLfRoNJ10I7At1FL087/ygO02hJhAphe8hEifeVg
pLYZatG2qxTOhMbdxD5pZhAP/Hy/ZlJ02pT3O8s5cW8H8GrCfuGtEf6L6grYI5jy
KxKlreunRqyMvJ4lrsXCWvO3f4i1Ysx2CO7J0GBxvIJ+dVY7C6vD/j8buWbiVGzo
1ytARJfIuXVLnOSWN6z/pk1M7bthJqpmOjQsBuskraCR0gUJZRHmZP5iwLRjxX2q
7gXbsT1TKfypVHB3hpXFEMNqJ/XX9geds7C1lwO7qxABU75RK+nBo1+Sf7y6qM83
K2Hq/kn0nVjm9N+0Ziq7FrElrUEgxoyJkgf1pWBszr71ltrInipml5+t3J5fl7mt
DvyjfSDHOoMbVeUvVtXrudVnsdajO59Aw/J8bbrFvpl0bRDcS04mOq7C5M0D6iaV
6HBbAZg+ZsD9sR29DNT7lTUQDQ9O+YSaDDVO7WVr+sO9LpKex3qf+4tVzD71ToAH
Y//qHzapT6tQ3DfRdFvlWTPbOVJp0cLuyIwo8XxYV+BOaXzgoUF1b0ATD+KFkfoy
5YYfI6YpEHSOR/xSKvxOyIiPQfyTAmhsmnKV9I3RGqVAUtbyG6yRpG+OW9y3b2AW
hC1FA0TUOGcFTWZ2J8SApmxbT3L8oNpZcxeTJj34KJZonlnLoV+aAZ3z6fk5tnis
toIZxQRMbaTDmlR9HW5XASIxdqA92N1gJ/qzAi9v+ziBWxEHmtvoEn8PTi++MVXd
LtsKDAsfX4trY4O3JtPgXLImhCgUxPqENcVVevZEoyA09XwWfVvYX/7xV/AF5GOm
Rp8tUYA3Ym9eYFR1HfHNit3rdCJbPbo2dpmQRDSN5jaEPnp75RKLgTbuLmuWUDyf
DOLiD4hXbhLbv4L30okplHu78UDWhttBo5PT1hRb4lw7iZT2Bo0C6Ctf+Ya9+wQP
6RWZIBMfjyF35ULabTTQ6U6xQEHV4mk6o8pHkrxDuxDJnFZXPY9faMmevpm+1Q8y
cvWQyACdVXudgvAZ4VQ0+4T5KtcFCcO59yja//hhn0mBrRtTY202s0QUEDWEDyYK
mzIeQe0DvsWXaTdNTrCqm9BrhtaKW40YYf4UvemVX4EPBwFvM5OkdBK8ssye14K1
Ey2zepE0z3ik8GQofGPd4lbhvG6eSZkdRNTadJeXCHVIIAjkt4/xPwUJuwPjIQom
IPn5c5zH0YJbTyAmTn6lHkOHHHz35Gx1SW8D9MZuYUNlnlW5+yOi9aq24uHJiW3d
PLqqKeoanxT9z+VmkycUVQAvCjBVGZqVCziOqtFi4WGfdH9lNpyAiBW2BdOT2fCr
9QDVVieqenfDtgREdskR4kAxNis26NMv/zdgnmyMmP3AfxlIJbIXoSY3hFXuIuIb
y+KccItW0cePakqNe1+j2C8KVTX7dePCIP6uJJp9+ZDtBPainphhYYhHdSRcJCE7
GhJxNJqkVHed3f3GKn+2scfpWBcLpr99RmbOi2j2H+G6LpQJ9Osp48BTkKv1qxeh
+f5El7dvcss7D5U85FB1z6RYtUEnArtZY3gcRSAsUkhqozwe8Yciwx1BKHQ9MggJ
XyR1kPaFf/wS+WnTWyAqmQ5Ogneb+fkGrSU2GevegNH/XBzDE1pYo1H6fCVFyNZN
Dcjjb35V11VWqiC4881xRNjejnvKIxAif0vWKpNZ+zNAeoJ65Qk2U1BzasTngGFg
BSvwMZQYP8jdiIhbd2r71EeHTAR+EBoJ26Cvv9PUyopseCRshLbk7dpyDb0lBoLv
JJfD9BbBjAj7+BuzsOHICxqc2jFoxmdyZeD+me42AP4aRCjSyJ0n+YhSucdedo4O
9T8vsltXVliJeaNCTofZvmdLcvghxUCDUcXWF+ShCunivSuojELx3JofBzCs0AO2
K/et0aruhckbIeBAAYcQorg+WsVUSVsd40LxW8W65WLZVf6deQgyDDUtt/Gl1baq
+IdlXKDKK2rGnLwQfbNVikIVOxju9QyWkJM7HFBDZQXdXgeiDVzKkqoSyqPPAXgc
CUCnJkNf/FvnzYrkM0UoqGxhJXrESOpEayJIRgMLJZO6JEg3C3E/fwSuDulYaANP
UT47Mq+VwIJxrWMYubLiYT1hH7FFOW6XBZzo9ME1b4I4YGu7MXUZxbn90iyVGmn2
xYQ75I4NpP/RfK3l17nLDbXsRNsfr+XCumCbwC5PuCT1D0FcqisbxGZ2LKJCkBcm
i0SpkEezjh2edR+vd/3xYgcz695etsXPJT67w7CV3mX0wYzdSGFexhFMKDqZbft5
2Q4y+oxMqYe5xgCNdyX3neG5Q0bA078zy9pLNThM2lxiSslvC+8wcUwdQHVvhufr
gBXT4z3VQLiJrJ49mHL+HeTVfbtvWvYOaIC40glyVajk5jkY++W75KzK4nrv6cUd
YAHHBQljtwCmQHJMzZs8f2V4pEyvcSZntzMnxtj6DSOzhyDctZbkTJuDDRBVEq5Z
waSIHfm8sR/X6GEXnhsqPad8BCPEQ+qaXYCEEYoWTlmu655GODs9qXYYOEiKC4dS
DChMGbxG5vEmLj56VbryWeww8lcaESQBpCPD1+Ip2x8Rr3nWFpdQsTOIanIaSWDN
3R2Zm8l2+iGfErxdtsccIdg72fBfff6phgirX+cRAx8JLuiF47WrmbBDEOAI5YK+
IF11R4TAnshDveZoJ01Frq2pnhRLlnBQMtCDnWEFsRIuJ4OjCHEv64E8TF6amswL
sl1vq/OyP3fmwky7vTPgDyvt7wMSdVtOs8FViX0adSL5APmZ2hxe30tCj0f+O2BR
SQUcFiBO/50tK1JACbZFm+IiPxM1Cp+jkC5ByMlZhpXNfVLEU8aa0/XskIS6L13u
05O5kXqgm69GsMRzp3oSWHTxSBPtF/k4KhHIeK1iZ6s6ARl4f6iassmBTrnfDb9N
JmQfDLSCMC3TfF0+fL9OC1ec7xQOAfs+yvs83OTLmEvc0luV32Y2Me5UYIf/D+DY
pQ/HjRNR/vptti+Fj78qe96SYcX9QDxKJ7oF1qu0tAAzpBAb6OQ+v5PE74z8rMWL
8v6JD2Q2uWf+7DLDnCsgCjB/yRNjv/4aCZSeuPiZx3UQ/BvlG6MWLJKyQZ9mdYpP
8721jH5gXdEGDIWCjmsf2NkDzoafRWGgHRZQ6JxKLWKOT0+SbrgIR0Dgzqozf0YM
Gu12N5r3AtYxALS0AZ7wuv3fAD+LZ01sFP2nGHDzp1vk2lfWteEmB5Jx54ilhXyT
I5u8c+CZjbPCfdRCtwzAgtxGTy7rINogxph8dKMMgUbqyHKv4krprdirI/65sNV8
mQ1ErtT3+f0LwVoeKPyy/yOmmritJoJEZ9ch8WKwW4exCNKxqn+r9HeAPv+KBz09
WOv4pZR8mCW0zgad440ZoHGZDtMbvqyd985GEMH172xrv2s57r2K3h0mBBS00Oa+
zOBlH71BiFRKJBWbhBbjxuiynDl786LRu38QVwBQubFNZie7Dabldann4ZxpSImr
xI7C2VMeaxmrxYPhyMNQx1UX8CgX7qu24qd8WRBPArjHywZ+yvqdbpyAuDrncDCl
Qldzg5szlK9ZvDAKUYMwdbvltMezTZRsAFHwJstYpw5uv8GYBAoA2H/dVpT4IK2/
s/qL+b+tNcSKBZRfzvKUkvxMMS7d0xNsArZifsXOzHcR4LUonXMN5OE8pbGHKvc4
Zw+e91arL6LoyJNks/atoODSOa73gE3pYAlyz9plcV2Dv7ZmCArLf1QYdidxZxv5
20siY3rAqXwBqmsbhuzKp7FcjkjR6UXJsbBYLcIAqtNPVhVN5bQNyutIsPymIONe
0pmMKS5YjsEy/CtcI3b8VYJ8Kxl0Cxdk4otH2eUiV6f5aAtlIizLZtlhSUoAYKva
vDUO0c7aX6SkmZHAZTxVZgaxbEMuWTnNOAsjEFbLusT9UDKgykpGC+NtQnLogAln
GhlY1ezBv6glAZAnWpa8+96Ja6YzPddY9JZ5z0Nhw+1QRbZG0DqhNJ3czAcULIOi
2HtktYW7DC/fWeKB+FlQGgymLalaVAzhLgiva67D3aKHOSCmdvf9CCPGu+0VAkCr
4UPELnEk+veWKgjAePe+SDC3e+09K5hrAQkjRQxW5DCkzc/MRgyCGnAhOAtap9M2
XZwK/Ol81Cj11RwBZ2KmbmAW3L6qBooNSml9x7BGFIqvzFhf80aXzdgR6xhF4orO
KFYo9dZf05xlTC3oATVqoSyVDJfD11g6ypIkK0KW5jvllfj4Mp6SY2C8rchSPSR/
NMggLYHzhROIyGBvtDNljUuBDkkcJDkjkE1hQEohCTYHV2A8HTGJpdfGRTNMo/AF
yXfoHkXvoZduFBRjQIv62bBO++UcHYOixRMcy6PnZoWzno7nKQ7tB9iy+USzjzAt
fU4wsnET5XE2ItnuFgJz01w8agOVAbqJikPi+0fgTRp38KIYwQNnbTEBP0Dd+89Z
0b7efw7VLOYrhH2ldibsRZnTYLLKuof0agVTPmSg/muysqk1TnJc+m+Cv/MURhZl
QjPs9kWGNEBFjuoXEirAZum7CB7DQyEShNng+DS78yf3EALQXwQ5eBu0JHAW9dJF
IF+i8yK0wEGsx/YicCquTdF3/MbuNPkiXHgoHVyTrH9+IH+op6gvliO1kaHxtM7t
XqGpg70p4uwKzCUjFY9M2uY1POzWfuEORrAVBEFWnvTKx4lPCqBLqzr4zduu9EHb
I7wJ1pmquo/a6BErA53I6vuRgeObYmO57GDQbiBwTQlw5AzBd7RRSrYrxYCV1mkM
fklUzggrpv6a3/7L7QEG2+HMZLXCE5aIiunIzoDLXSKLN7eMMNsQSGEaycnqL5ZX
DmblIWqVVbQj8hzPbos92dHrha/aj0tbaK/1kXPQvtwYLGdU7+9JrQCWv3R1RnWc
kHZLb83IW0xCILEKDG7MrYTqtiGZ/oGxRM2EMRkvIUl+RJLtzyqmzMYw21Up6UVw
fyb8JYm0s6MR/d46bUvaZE2vLYtnn4JOTMzH6AgZKnA+hkpZWl1kbg/ZXd/oik3r
+auPoO/u0+nwLjYR+a9L5Yz3ouxg7gLLt60Vf4nXErAh4Vbk8QBI5tS1o2Kl5xnB
nrixBmBxtcPGuEyVS51czktns2AUGkphtA6KLjYxpjj2LOQnnd4iXmk+/PSK1/Au
AHRwIQMNHbOfTS9qDelrisf+40AxvA0FlCY5ZGuoDWhOjq6bn1wRxg/Ct7bOpISs
QtnFx3KgdWVEgGgrN/XxaZlyJn+aUYfVkV8am68eTMNQ7DorbfP2gyOitwPln4L+
QA5Wh9RyiinPuS52O7OBqFWY6zQztGuZOaIoRFtssZ3RVgKv4mJheROnb/i+9qmB
fUtu9Mns7Dgt1Rz8qv8d0JamBZaZKxmVRWKpBiAOYFDyELAzzAaP2RXhZuTEan2+
16HFhUiD15dXg8//7VBuj8ELwBY1jhr36gow/YxYsfBesuK0V6shiffTrFZTeuE8
aX2TMz+Er/DgfQeVUREjLr/QS3hlp8C51a2zkQw6gEQ1oeJ6Qip9+RTYHFTSjcg4
yZEY8E9Q/axdVRaJjy5BnwQqjPB3X1+PvimM2mMEXs6P35fvrPTWToDNRGxtTfrK
W0H0Mi5kym80UkQvwIQiEShEPcMLJzWPQUop6m3mFCcovJHASeul86aRuw5DYGlg
1Zwzi2FTTszpPYcjs+jPv4lxzRdCTJQR7eq8Wj/LkEwEV9H0nBa/UKKGc3+mW0ej
W1QP6Ov4pTm2XIyHhgHcd9+GMi+DXm1Ou3LKYEz/C9QL6ik8++SItj+4EA6xG38p
c7tfd2HefFUgtqVSZvH13ZJswBLWwHzeb7YDy0U/U4K/7HNQx6SSpa83RbDMVLKs
P3RHlTrkakFBWpnk/6l02b/z8XC1SCOYOzHSvxBo+VbctUsmbrpc/BmYkXJOerdg
VaU20G0OjB5ZyzO634ElbLYlg6xqh9W+t3+L7gRQ6Y9D3a1vnoQA2DGXc8YGLzhu
GEvLzlxUocagAZUwdbW+ANtBsDThw4V2VJV+MfaEQvmoTx4dUu9ALRX40AIu7mDQ
656aj4M3n6+DdBEDC2+8HNyNqIhGTuzJ9kXpPg0ERykwejjUqC3TuGVl2GrOqfho
2Eb6WhN8VLu2dk8E3gVNXi/D4p+oTlfzc6fl5Gla15QKlScZ5SWCUaERDY+fo24m
Rm+5TnmrB/iiOTuuGAcGhRpQKuBaUTump6dNzpBn3lUuG0w6bwhO2+DbuB7x93F6
kALqu+E486FBFFyiQFJ/h1IrQbqImeIIR76Vq7vbErzUI1WoWzs8B56rTnZgf+6Z
o3OWCrdVUC2+FCaDyd3ayurgFcQCGW17CWaIw05y938a6pomFkGBcJyWCuig6v6M
ZITdb1R6QU8ksZrbXWsHJaUi6cr7B543z0oAQSqS5XvTcWaHUk6DlkwXVLoabO6J
E3YyJNFUEyOGsi+XlVQeWaO3ETgK8MnDrq4zzeyoluGN9N9pb892B+UFb01FCFG9
t7hSzdj+FHP3eUIqfqVXcy8HAKngDFqaVEIKUk/UttF90vyIWVo2bsOlnaZn9hUE
oKV9rTdFuZZECu9YSQmt+Chcr5zOwFben7ZgyYy3WML2ckVyoLizsrwUqflPIy0+
yYsha3b6shkEuD0XRyan+QUYwkcrdJbbZ5VrXjpYN4eARhb6tJ8D8nNpk8TTUdyL
mrCYigCqUKfjOcQ1YGKS7axC19mDrAF8FyzA2BdGyKJGD809Q3rUzSwDpSvHDNIw
SsLAd1KcVpmFZ5x7xZkxYpzY/0MIbEi3Lp4ewWQd9na4M0MU8y6gleVJz3btrktg
OiC0iMo2BDZe7NP5fS1lBuHFFcXkugk7zqdPxrnTxJ4kOvb/FPHoZICttA19H5Bh
QB4hTv3qAXEbSGmu5e6E2dLG4XYkb0dUP1Bmsztqo+lbToLWeNMCad3XsVCQaygz
jbYSAhtCe3ozFXiEVj2GcnPlKYaMlZ/if/xo6Or/fZC3u+o6d9xC4LD4MolRoUWf
BVK+hEdITHbHmtrWTcD7opchWCeqgmRZjXb9Vrl+N7IsDFObPP3GQX3HCEeQqH7A
bCUb5zgV17pew+heCqOd3Hz1uqmvYEOeBVEV7xA7dz4udjq4M0pwMjYLcWQUmN2I
dNNj0AlAUZI9StNl1wnP1CnGxQyszYjhoc+epAO2H2zFqOEue2UvW/5ciWwi0Buy
WcOM6Y3I+gNGUMdDkA1589zLKJwFNHgyXVG+clSCXVbUvCLTzJCGTUXP2JK3QieA
BrgbzqElDwE2YwNY+0kVtviNqq8VkWEFurpe2qB4VtJIP8awP3NRK7d9cmgWCCpZ
frIH6ihpBzJf+O1GhuNy1Ij1Gby5yuUGGrGd85ZRDG+GBIoi5zwWfTblXw3UnxsI
W0GoJE86o7xyYxqWQbdJo9+/QYZ1+SSqj/umoA2RKMOasQ7LVvDD9Q0fJPmQ32vU
3l9uqRRAqR16+S74JAoGbKCl48+7Pef+cBI4l8/xQT4FrCKQF39ly2UbAMjUbtTB
Z963uxYQ9sjoc3zRjGTG8z508jsdqzsLJmZMZx6vyxLqT9IUcUBbrDsWJ9+YMX1D
OlLFEbZhmYi0PnXELSBWkUs5qv6WBqEjZ7xCPj38QyVoxoFVF8UPGawytkgf7gRR
cTCF+0fEpcO40GlzFECpMmFkIPfm/vxq10qlB+XyayRfFE0QG8NoroXfjRJH6uxX
aIZ/xdWlcr2tebD/qTLqQ6dHNgjkydYgconvQJKlO4BjkFijem840NwlQvmiAy+U
xeCKb7PP1E0LSXLxvvXQiI7Im8qznR7x5ppUcEfNAv5+qlpZMmLbbYh01ND9XxaE
v30+MLHRxXq2Z7Hnmg6+BUpHIpY+wyV7o+GUAC7MHvGZLOd2fKDXDPi21a4+cOuP
mdaHd8cGrlsG9GsYvnlfoUwCXyqWqxrcy2/U5cd3DbXtqzzTxMiHS236rtD7l5qV
f4abEy3eaoewHv4nRENSnEwS80gc77SsR/HbpP9XxjUA8qyQTP0a2eMhJOlxgJ77
ShRT4jJj5YfKRcIiaRo3cH/edfBHRa3H6zmGSS1pKtC1T9e+i06MOAaRUfb59EPx
vcG+4d+86KcOCrLzD2H5hCDYR3o3w7OcnnuaDsxBwe5ahBQv3WTZHzxgKdEfwCLb
JahXVG6+WEWwDQ79EmcXxZaaL3qmjXQiwbA3RpFRfGDODa3xRSli3+C2+rp0TwHI
Hi0NItG/PSfREFViwt+IaIUQOEZPzLbU9dEV70Er7Okajxf7U6e3IhVCDzNAx8xe
c0X08/o38uBNnlbkPSll02Fwy7T0fk5IGuFdAHZB2on/z/Der72+W1EP6GNG3+Gx
pctk1z6JuDXedSzwscj5J8STR71F1bR0X3+qlQX6YD1vi3pdJcInGPXR1YsEASaP
cozGQ6AS9hn/ZaxojSleJ+ueIntTrkhViFyd7RZYajt+cvo9yfCSMnndCYclh2JN
IaJ37StGZsZPtwNzeejQB4HFc2rPfz8RFz6JzHAqYGHCAKNkYksvedUMgpfjz+5R
SW5508Rd7yQpl9iTcfVtNM+lNTM7ynpYwqWzboSyz0GWisq1EELotXXo+P7cKuVP
yIUYLcXrl+bfnYFFbYkZyh4Xxp1yd2/ahaMgLoSWv9DGiO9vobPd7WmR4B1UUOb/
NSNjJi3XSlhxnEOmTaqcnYHSPnzbKAobfNO29pkPXwdmBHar7eBGKXCewzkspG/B
C5zuu0tO9BA0L4imVMmUkfsYIPLBxXXILrlG6CBT4BBziuXgAzwwb+MfApWry8wo
DV0Tn3KIhJzGQYOC3XJVRIMr1g5mC4Z9tn49e/EpFBgjUfeuNtdo4uYvlhi977KU
5S+NdD769DIj5EdJoemGqtA29Wvkvkug70XEOgeJO/fLTPPzL+lGTunEp/DrwICX
PrFuck2yeNeu/hXvoGftHF7+tKPCmwX8XX5LMAp0iyBINNbol8KP0xtRxnWJjsPR
xyhYi6VO/mi58smnJqykFo9WuXGhOeNY7Uoyv1Q3yBMpo8+nkinF6PImwfKXPO9I
TPtm4smqWPMVwov5yH0SetK7JqhZEtytjp6za7s6TpuiBSZoSGmvMJdhiG59iQjM
Z5oqoy1QSOBSqPwMa04ROCkV3qz4nbO9e9V8pX8xoue0rEMgTmaOjsXd1uBL6qZ8
I+sTcYbg7HcZl8pb7+0rHUMIQ02Tx83p+2IGGuyWRlpfaIhbS/OfXYHG+lKsSl1W
3lNRQO9bGy2lJUjKi/aiewHvCbXNpG/XFyY491eYQE1Z9OqWJOsTtpuDxnGUTzIu
aptASfwfCXc1m9EBopuncxOuhyvWodR+XZ9vrvxF5GIpzLJThMzUoR3x1kyRQbA+
Pw+F4/w36DT76YLLPBXs+791v+8JcG/QZk8zQ19oHNO9crMG/sBRV7mugKr3LEb+
rym6BgHTx5ZFtRVxUd4QTNEQqy/e2pbZGI47bIooNU7L0fWrrMVGVwBLw3+JhQ2I
/9OxKzgGMu4Y87HwYnzNrghjMzwNkvziLZhZg037YLRW4lZRvJpa1ICtwHRj+VSl
wULP4jbJyjDUbwqbMJ3B5RjigwdUT1Gx5DiNWBGuQTqFP08/Z5q/JBCx85IXybCs
qm9DBaDqRkAwk0FtLP3GhAIHkOmSYafM2Ihh4ZXKe5YVTKjnqRJckMNpyCkU+e3d
E2sXtrW49nO/9syfuScL6IUKsJWmbQbUhtfW8RUlkB2CYNgIUExxQ5z1F4l3fJzy
Yzu0eJE3M3DcvpC0AfFVvtlMLVe1Z1yIiDwZx3Oj9qyDGHzn4BzWpbyGLxXoChX6
pf1PLoFavA+v5IeRTdL0zR/3PmnQFQiV7EYgEyEom4k2dJcCY65CSpMsUI1kuS2W
rqKXvt9395FqwQz+FECqamrqjHUcet1rJwdVpG1Zg64b1W1PtE9d2Id1NaivO9jf
bx8aLf8wWwRSyT0abn/uyvTqRgUVHWyb2FbkPbdImmhHKbgCQqemZzAU3WChJ7Bd
MtiboRrPBUUpj7OYRp4dL9Ocvvi3VQSXwIRHkw0VQMSFWIdkAQyKpTH+/8Pz1kFD
5etYgxAkqwGGfbtTcDi/FZCLCIxmbso/Mw2rY/ZnBCiJfb0TeLX4Wx8emRmXX9jv
8RrAegop47V3eB9rSgCfg8E9y5p34zqlp5v7oE7vmxkIUYLyB7tQ1NQ9FCfRYCEi
nV0ErTgQtzubtCAz7xT8h0zxwS55FWXa6xVNh86w23cuxVhyCOTqH8fYqa5xJans
bJNnyWw/A36l5V4Wnquq3EUDF1i5YPH6dh3/xcLe9Ge7ffTHcQB6hdV1BisOJrV1
cAyWPXIhFhKjJ6h0fzymfI0mlboFYkuvUkHRtOleCFq6ottlRv2Ttj9OPIKGa5Rb
/o3uGzQUX+HYZfCdV8wvFPgEiTRkpYWSaAOFOMDJNyWtFcnx/9UhFy8LwPXs2W5J
MElsLHYj9ZbOuFyK4tItuJsxuJOozdPU51HYUWMAMPN2rGcHwnlVAsbb98pa5wq1
QygUyy+gD42xI6XdEGh1azrF02gmga5uVnwqukaAAbuhHKM53LYxpGhU/6Qp08nW
VfE5NlVKovQC8vFXzjTPNVzxxkQbZxoPrWAw1ZyFDdQ5xPUg2cFhhBbw2MAo2Fnp
GWlWa4GpyvqpUHAPSzZdxw9EanqNtNpZpMH/5wXR67gKU+hGOxAjZrv67x2YQvaP
J9Qf8ks92rxUAVaQz6zHXqmGhvbrMbYbNSFn3rK2oYwBHYZ8mp0jz2RjMmTrCK2D
0JxXBTlGwILMwHDeg1+aIVKobFGvs8CcLPE99DojJfZtYwK4mXAzZLpF0hlyHzHl
x1ccfrdMjZxlQD+6IWOSwqXwqltsxqxg5k1RG2JNzAeogvN0XK5rduigNxbA34a1
+RAf80DCDHSDLIuEqnHGA5eat4eqSx9nfZhuP6PyIKBHqA1w9DofN/y1CTozpM9d
fG28H02vUTww0rFC63RF0vmiO2HlU7qEfq81SosKPF8mzt0Bq2xWm99zyIDTUAJ0
hs39knM3P+KIMhax/+NRcZwgsIwTOmPkYsOz0kZYejI/2PSpzEHBr2OTqhymOsgy
zBjESvmrq6odmP/DSY2UEooEIP5IBdzw0v1tXxCExzz2ZCeEwqdqZAWch3AG3Bhn
QEzvZHwBACHa4DjaCwNmlg5+hoeKw4Womtbv9WC+tB55ax+tC/5BK6sLKyNdiYEg
D7UiPbeKFnUDS5VX3FDxLSSHwxujLFH/vo/5kVY2osX+ReD2UievdHo0zMU+6xn1
SLSFfJSEtlPgwEKWKAuvOZQXoUhjxhMqaCv1GKRT2zfDwtnjjQ6tVODNlG54hC7p
n4eWxq8J4ry2uNJhAwG4kNTGNpaSjFtELMfYkHfTLIDb36ci6vOjO7MUbtAo9Ydm
pks+2Vq4vdQBtzkBpjmjVwKrK6hC7S3kCDRcp9dD6EJ7pYHn044T+42vUIuJOP+m
EUH3StZeAg79bm9TKngsotB4c2QG9Ui5ngJWE7Htc8hPTt6qYoiAwS08JYVlEBvz
QEyaC8JAiGcx6jSIo4Q4ALRM9is/762swNELn+ERHnfFhczwp/lN4XEl/icQWSsG
YKFj1Fo1tXIeFVtoxmBEHSYR9luFG31e8gP6XeGXWjSunv487piu0y2R4Nfaj1Ss
9mD1B+L6EQgQR/7YyfdwX/mq/EPhO+6T+q/hum4OoF8Ynv0oWe/israiskVWakGT
El584QZvMdQYPBxw4URJEamcCEa6HsFSXIGwlpxHm4tiMjr9AfcSHq9uNfH0XRYH
c310PW54vKpF+m1wFIfrNxk/Z5ZbyWaX92e5KzUxryOBkamGCBENTtubwIb6Sh2/
P8Q8ZFQ/jDG3xX3HEnn4cN+on+UM1OrEsENQ03wIYbu4YVk7JiU5STU3AzNlKvS2
VBmx1EcUEwsVqgoWiYJoCOL239SabBq4zI20vRWi8q6BYcgkI9bFYymMgizds4Ez
k2YadJdFvEU7RQaOrhScH7IXYvhLLMVaBfGwgmRO4P0Lp97IUmWHg3M5287B0thr
8Nvx3d1R9nt4jrPs30NYxNxOLOfnVpp09Rd5qMFigt8wtCJqUaozirhOZ4/u+B99
XuUUfR9673iSe4tAAZDI6tHV/vNObjQPz+ejOH/MadJSIRNNRVFsQcpK4dI50QIt
torjQyUDUSM5H4lUe4F0HUhMEs9EqNpejsuMOt5w9X8/wXOgjUZNBQ9Q3/ebmEXF
5c2T3EPly0FM+pMsvkqJPiEchWM7sJV9Ptwf/IsEfhjoQUFuXGDB37MXwqWhRKh/
bzDaApL5NU3Q1jOW2D9Cn4RC/SSbG5nwsK08g0QuuFHJinQTZiTYp7/2ZcvHVbB9
7UTSxKwksxfhapEcJutsv7U7CF0qqzkrHXaqrpwLeJyttDBf+8s2XKaCs/P0/SJZ
XIcM+Nktq2Bo+yj/kHX/Tot2Ta+dxfY0UiKJfZ/NGepwXTQ/m+FwZAksCuwRTlDa
mgX2nt6R5mmvkqwvAmUSMXIFcVjLQ6c0X2KBZ3C+lCwjGa6Xps2YdWhHfzglTlXS
j4VGkhnZAp8RDrsaomKjDOEydQZdyGQsVU/4eKuUYvuzAtZQKPjlAd5IXWVZab9P
R7UC12pW+0ni3Q3mS2uy6rlaBZpEawzWwV1L3hN449TIVR4UJMglFA/tFK5/oniL
YEfttoXPjyV8A9QumPztS5RBWjHfrwQra5pNOpbWBgREVlDzxqP7rKmyKZehw+BV
593yobSqyBgwRUnhImJZx+F9hlEcDJYn/goTgjvhtn9jlb2RBoua6rgGjnqeQ1Nb
RLyjs/+UsS0HMBr7dkCNNAdC2MY149T24yEyIixghlH/5VlW3vSPeoHc0b/iU0mK
3hKbXZsc3NINjs55B3OkAC3Jlao7cjk9Pr1WAf2SKp5SvaMmnq8RBc9Y/e1xU2H2
27iha6RIhz3qNpSloRAHYsZsw59loVC4oP9ccryP77E7E5JFKmcXP3hk9bX4tJ6E
4R3W2ybiIY2K5w87P8BftO50nVnhIHCxHt8o+7+r4EBpcKDjT79Oz9DhNCmEa1zg
Cp91NjG+nmKCEpIgqLf0NWzJPMMXoMgtc6cdlNxx3eZMII6kcSqQvCCg2LwQmN6y
ph5Cuicnv/F8WsOnxgYD2Lz+e8IZ0R67yZEdzB51Wrumdal6af+4YAqT5pPGkw3D
C47JlcS89uUrL1VLHUELk9gENqe01yHTAmW8gwGS5NUWXA35f2JEwqGWVz3A5iz1
QBRyCaREpcsH5rf0RrltoMSTWBz6D219VHhiD/rLPCpSPbskhMpY59+h7VXe6u1X
WmBipYAD053Lsc7XSM1vMss4jfUjcckG3Hh9JiwrNGyjBbmKZof7MfPrJpfBXQIY
WFIo9ax5u9gYF3yFvxSLsA/NpRPWQstNSZGbbDpiK9L7E6NZGI9Mpsj3SNb/YxrW
51qIWI6B6IPmU1QuaDr5L3t8oz6mcRljAT7FYe81x54oF0gF6AAilzOxItn+TGcT
YrKXtAYUXI4AQ/T1Z32ycZ4Y9cz2YiHlawTR81s7WiFLjTkv8xcs1BaJ45mChBGs
9TeSmJV5utoEsFGV3GZjAr2AUfs9ntjzhhRysi75lCx4eX1W3hBy9UPGsS+HTiRQ
/hDeknsk23L5usE7XXOUA4Klk4zqxa1WMwBbhReIpjruavNnp3sCed4kSLPsu2Ry
BjS4YCTJPpcZZxvMkXEUfJzREhOb5nDC58g77pXzQxvtXmJC8YXwuJZksq8lEgm0
fUYqJrG4M3hTMDxTSwNv/8GBxfFxGHekegfy15zTI+w21gRAeBqVxrsXgCis5x0M
fYNNWHibW5xAtAUHWzOIbK4VFRmKQ32I2vDE2IZ1nxDatgCqJCE111KhD3JzoQ26
cRbJY1DaIuZbQc2dLVu1HW/t+1WErgAbTU5iM8wNJb2zOqjUcd/pNjYG/bCWiUvq
6Sr+xyoUj1QnqBYCpdnWfh99kXGGIFsZOtKmeo53lsP5DP2LDA2WgDSH47yVqo8T
IaYeuqN2IRpKdWWmboZG9jl1c1s1teppkr70Y7SPbnPgIMv234zR9Y5q40HhdW8I
4XJ8GIcpFMD1l9W9yWgONXmPgV/h6CkDKDa3zS8/DHIG0Hj4JseWe420YH6xm/XM
coUm46n8arRl5YFPauQwO9lXV6cwui5nzyJEHgEyO4dAo2eiY0GW/PF6mdXaWSav
yr0JTzZHRUfLu7aNCbh3SaGLoqzKhyfkBrIfv0nWGJaHxO8qmjC8eAt4q9LR9P2N
VV/IqkDgNMvtr1r8uSZ9QgcHdq0T2YyqacfHbhcU3fWk5f4Mhs1Knvpa2/YlQTlb
e+Mjv+qZeKVlJkWH54TTb8TmSMKkeIqFM2Mz7NY1b/r2HeVyG5zyrapIgy27yFNq
1himM8JhU46CpHCDSsh5fcuBbvhqyPw1y/KQidgIIxYiTtXUtFGr258j3PTKfO+h
9JOEUtKr36g7Ojy99vw4akVHT6c+wWQFCEmTdyyv4EAnsOtBGZyjODBYgqy+ykq/
uCVidbUTcdh3ZrjBIiYJys1UkIBDxzw5R+9+pbbsWEe3698SM6NahoNSxb33/GkH
EkcvvEzB77qUh10YsZYoFnwcqW3ruAzwEwXTktI4iFi2p5JcFXnM0I8Vs3de5/Ga
1vS5g7Ob11OmUDU9vcDISZOyy6re2HWEbf4yZ/jVOpDHFZt6CCdJCSeZrIqHtQMC
4JgdYD6eyczEOYC3pkLtAR3asMhVS2fr3ykRJMqT2dTjdarNXhmm80lwiC9R+nf9
/f1KLMoM+l6nCOZ9XnaUXUtO0DVmJ+hutSV//5mGzt6dgYR1HunaKcPZrmimRSGB
JhvMF5sNE7Fa0Z0/7EbQEpjKijipdITS4C6XCwcGNt7M5WpnEggEM4L6ONQlW7wr
pNSS5/uTfa9Kmo9DQDsyy4n9HAawn1mnp3iJHE/t/XIVSXx5/mUWBKKtFz+dpudR
S2wea92KFShM9DHGoceTxJesNgRdZMUvsst0JrTxeDPdhBRLMAB9AHKWAhLZ5IcG
lipiJLxtcpxnNWh81LVmQdl8XMiQ2LnJFxvzQc70PZMBF/CHsNZX+/R1hDE9PQRg
zld3cyyvvYZCRHTmtTUc8G1MOb/ggOjHAQidBwJ7x4niKO6f2V3o+DtvQ8wVPUdY
HhOOAtgnEtT1A2Ust0W1dBiX2UR2vmjiyIXfHWpWOm/vXkJYwntFY0/n7xfL6PAe
JJ3c7OiaFKbR9gAs/Jsl7/A8l4G1BATnpxZQp7F4xMod/EW+L1tUoCZMFgzKja+Q
xgKZvfmMIJM3FcTtSmGJIY1V1TNxt/ZH5B9zqq0GTbus4JJXhsjAscHfVF3RXfCD
UiAymex+0z/11CwEkiwN9ahU5RAWhXipzMic7oVucFLVrMEBwEE23UOe4X0vzvhn
KvnZNxcSRKKSN+QR9t2b396DJEqB3vjsVvBCxAsN3jlbu1211sjTZ0eJI1tb9hei
U0vVy8cabOqt/s83XP0aRnHrbA8mymlNKYl0BB+T4wR0OAkstQbSHexZDT/AmIij
gUe69g53Qtaht8qeSTQFLh6+4GbWhApisuJaNQmdrvhg7PCyqcZywvXQZZETTTm0
y9/b9cp7xwRQ/+70qPU8j1Uq4TozCOkvqYMAmBkWWtzM6MeJ5LgulY+HSf2rMfpm
aqOlCJXyBRMxsO3n+IWc1MXtag2NwPmlYseOyCGcgZUdetI0C0yGe/eoq439jrzR
DJMzu6hiEQiPAAhnkca1SyuyuwWIiIGOSaTMeJf5JBxhjVOVF45MzQwRk7BsIRho
RmiKgHw94hjnIzbHIZFDhBKNvrmhLMJk5UxvxsDQjlzCsjqYGBcq+p/9HoKZhsAJ
mBBYB3u3JPkpP/nN8wiXAkTcRR3pZvyOXf6M6AOBsb1CUktcOv7Bf05hbtCrc2a2
CGF3i9MHNkZQz5OBir4HXaOOrjRfYqW6UAfAmZqlK8bJJvwC+8Fa1VYSWuIBRjpC
eQhSR8Mym0mwGuoSB204Qe4dZQ42JpM0EvIdG54FPTtaTFXy4F7Q6DEUtfWREbTz
HlJSLhBXD8Eh2MZRbep8C2/Y2Wcdark11vyX6AOYysGie2pxSaydKol2QsiJAtu0
urlZbJ27wQYQfzWKTpMOCMbUePE+iuSR8XlJdpZKFl/KkKf5VkiEJDrP4sqZ40lB
Zk2NYwXspbA3fCL1PNsr4i8rn93K+pASw3QjqW6DTa88keQ+e4YQXS4tw/pNWL+M
qYelUW/cCla8ZzWUellNK2zI7z/cHgD/esRzJ/fLl93W3PycU23KrabxTItmNphd
pwo6UVSND/nrgBpZEp1KGtN/Tbx3kBJ53eFfmRhdfRK4rlfOaRaYHo7cmvrv02tS
gJ/mgp7wZ8Yi9Bbgpc2jdFAnM5yDMNTbbUbJldWWCo0cZf6CKXSP/Hb7aOkUJZiR
Cf3KE+ZS+00byyjzib58JuvBZF+lCFIT1eFYCwYK51iA17gLS1LiTDMRWHq+oNt2
MTDfXflvdKh1HFcmC4/HieyaX4dzjAJuCdyjql3+GloRTxFBuUlbTPZaEM8pQcaJ
mqy1CPVI+HgSKoqkxYxSmmnfwyIY7wCLzskAypwuWuZm0QrFqsim1a8+toD5RZvB
1S3bn2ZiNkE+M0D/NgqozXT2oFBXY1doaklXWZZyLXlsMQwETgxFBQYUUX1howS4
pdzf8wlxA6Cktgg4tyaqy7hqgEAL6slakEy5o7/BBsU8ehz0eflEoWBpp/3QAEPX
OT7FGl4i/IbPOkIdZI+3iiNyVQYYy1AOg2px2g9awUqW2yYc2/gV6pB/p59tSjAF
rCY7fK7MPyJAp39i7ZxeZsH7mI7oMcihkINelGWGr/R+cfAwltQYGVCYwX7wW85N
evQliMs4jLXpThwVEnYGVgopxvQpbd0Oyen77oi8hL0+ZRn6mfLw9Dqt8tHIvSUm
qy2WJ2kFCq8GmHwwF0eKVvSGXbLVSVGnP2aREdRgTrBJEgVZOO12aQse3mpIxB0+
PX0SOlMbMIiUkDIxappSVdi9dktqx5vhNaDeGkjD9cil7cfYbPNdEP/6ypcVwKHd
ezCyOi07IW9u84SETb9cQIzaCEF7WO0w19pcOwF4K6y6vmhnfnKF/dVtdq9X3KPZ
ED1PD5ur+1LgISQccmV6THl+kEFuhogSl2x99ve/nRh0A6OIqn8WrtTLCOi/dR48
E8qqmBa0z+8nSb8x/LWfAdq8rKxMQFU+vznhVFpnw+uJ4hijDR+J+7hHCLLJFr56
/P1f53ITANirRe7d2FPFefzHqkyRQeQRchoq8Dygmo4eUS52cfGvs9Rlk1Fe/HS0
Wng0xWMAgHJETBpaAzjPHZSQn+86RTUSBiHRwWr9q4mNgRSs4FU1hLPcFFY/7t7u
z6Uwsmiqn07Xc52sakqJyY+yOVBaBA+Rw7oq/1y0+UxzZC3AUvXXMbStvqcZOKz0
wN1p2/mN2l9Svq5ss8nibGwAWdy185bVuQsUkn8lO6XTBgAHJa/i81nv+Rqf2t7B
ztoH1na6rtogU+aYdZd9OTI6e6bQ1YZggpDTV5Vm04g8BywH1epoLbYi4AJnulvm
Di0v2AhatS4IJqZKF0zcPs1fF4u3WP0RWuMLctocHb9o4FDecb0ynHzf1R4WwIBm
ab0TqC453/lCC05ZiLNe6AhaZLZbIkiI6WnoMWNsze2Mm4Mn+1/i8NlRclmZbY5t
ihndlGe5gp0XNmKW/CjcEmziTj/YxzX1O6XXCdyABIZkr66mPJDobu9Nsgk8x4Ds
ZrwTQMl0yvbhdLgu7T0UTr/JcHbVlB9EGNtU7yBC+V+hRc3t33v9xkHHiwisCfSS
3zHAYTkC7goSNMpD5omX151F0LVYqC/bJEOSmDGTr/ydfQrfox2OkOs69gTfoLBF
A8+RDjYNPJXAaRMjmVK9NFt/SGH9a/RyzPk/4zfl3vcUOav//MoHQ0/JmPJZfEDK
aGNFmKVfCBsPlI8BY6hGILbL9dv299bcDx+uiE4y8CwiEySUaBQ2z2o0UKQdVfa1
q3nPdFAjVfCjTVEj7zpNSvuHnYBP7CL6BZP+2Qr1PV9q898HqHbCKVa+9fEfHwaU
Mk+zCf5MDEUyUPIobrITfCxBO+zRMDFZmmpgHjE0ARCq7OQPCWxHZ7D+PHnsUxf1
eAmzOBSuFcFiE9IedZ47x8WN6x56iNN9/ptDrHbkGunvU/wTvVrQTfQ80bSmjrHT
FbkmHoZmh3H3XuigRDy3qRSPSJmq30MMdqk/WdQjLOc9W/R9iHqHDUSipNW1zK0O
Tn2u6HThSj0jtwPAef+hnzHkq61ZrAe+uo3KbYyaJ85pYhO6grzh4/Gg2li6d3xG
Jsl6LDcs6Lxmbg8+9aOtxtbOXbXdGNrwNrmF0acPB6/x9ObNW93T8K0oQ2mWVz2S
F7WAZhzpzE+Ym7rGo18+QsQvEjGst6yZFSrSqBg1KK7gieuZXDvBVGy9/f5rFmUg
2xeIdkV0KJyrT/aX4LLMR+xCtTpdu/eJauNaZX/5/A2l45XvxWSW3+JhmqFw/0Sv
rJdKJHKrmGrZMyd3Rdj08Lm8upaP9Z6evIYEL6JlII9mPSSORU8yXNvLWp0wh6je
+GNvJIrDcah0YODqQ0nFof5FRhq8xltg5gXNH00IoXMCkE+t5YjFgkWIizqnuoy9
8CSsbzZ5xGd1I2EyJTzh9lMGoakKtPFC/PDafaw+xPJWNOPcMoVZ1he8r4bp2C4+
shKjU2Xi6L8uojAkXjbElEDx8kEa+raCUcoHEcg0SykG3bQhc3rF2nV6hBr3vdfF
bGMfO09AVlqBNREW3z6omH6kuxhrI1Pa9kxvoFFhiAbyArGCxsWsSe9eVUSRWCtP
hwA1vDbwjd+af5UyBMK7RW7BDQQStQdpoaRKN6c/iPWt/wld3LXRX/fo5i/Uaz1f
FE/ZDE0O4KZnxvo0aBdVSNi7ZFFz2HOZF88vg4Ybhf96bOmDyC4ZNc3qShyLTmHS
wVfa3u4Rjz7nlppGOKtbcSwmFN1QVQmhaytYJUswitL1yB1MDVytia9XopLK5mdr
ctqI2SrZOfam1zD4xjZ0C46UL1dl4NKyIX2AUJtT63STx7AywKFX7JfblvCEgECv
//5O9xmr6WbaxWedCriUfzmgsgKcFwwhoguHp5huYUjmX8iNuHN1p/3Tztvls0cq
R2K5YMIkWPvcjwh0nFrhRj+UVTnR+pGfGKVTpClBKOWk5myC/IjQ4sRoCJiAaaaO
g2SGtwyPc6Wp2CTEADqu61Sy21LShFMpHrD7M3t/AF/RQafXLQJbjhdHVjFAoLQQ
a8H20w4GaAm2bQCkGFB29mVsskEv1V/yWmPtU8S0n6FFaOj7dTifQHF/EN9GZpvp
gsV9LEEJTjpkbuDrczmarzhUbOPo0+bKtIuqAdnA63tulO7+JmkwWj+z3vU+3ceL
06suIaIClFYpkU0Cq4DgIv2SAkTo7Q/uZ0C3t3OxcElE5kW/1Pz6gz+CPy3Ox94W
ei7cgW0bswyygG3vnHwrxkzzuyunCszaDdG9tGvt0fd7TE6YaDwbNtfN2yVvjSf6
Kxbdlv7Yt3+wRTW6AjIFoVljlDf90UWw5MwnrvMjHQd8wFXdJYzhKNRR507BFo9b
L+a2itkrJZXEb/9Sox64p3dvJ9HLGGPEbNS7+JYE3H0+yjgkvf89CEFUhW1Wf/SK
k0KkmJVGMOcje/BvuikWK9Q2/+aMT96aguOO6NiDZKtscXDa2CkVe+px9UKMOHY7
bxXEx4cmlzJFIkdfywZLVVAs5Qd/XCT9/xG5AgRAgpy7tbOEH+k31MXLcD9w6Cx8
ea+Iiugy4XiN5myt6/M3pnwGVSwmGrrZnbFaj7ydXDwJXF8zuAijvxUROVhKEV6A
juKIizDO4QySMquUw5d1mRkmnRIfcICxBqIM8GYMcHjpoAfcNeQ3R/GvljLl3kvL
/ZZ10L0xZnbC+02RhitmmELS3xmbSE6k3BAQprRW4gtKAXqqIeLAFt6sLsrwu23l
GNkYOtMOf1ohtiglO94j+KCd+7mtcXCNIb5M0OBT2cpDCpC/+z3hz0KC52JGp4Zs
LF9fXO5YKge2fssuZypJX6uXl6M2avKcrhfoAhR/myxv6aWV3w8TSeEbS0JKXCyM
8i7OwdKCmcIESAJWB2SLnwRsbWM1gPWwY/Cu+XIB8zDEFAuX8MnoUYdPKxHpiS26
tllZbTpAdlgFgsCoZeDcyW45UNPnxC+7NHAwoL4GJDwWFSjxwTuIO1hOU1zotFDK
fkFTc8dMf4tAuHPGQUe0gWcLA7p46yxxeIqlD9bYu1fqsdyWuTdxCmR3jPs+Cia2
dAwlFgE7KNqW9e7LQzHYGt1icR/cffobWYcBI0shnKFj4tcpP8fzA4v97IOIo7Sa
iiQ80nCR6Sif8jsedOX1GScCtZ+kVs9GqrL5mxj7yzZ8wE6SaTYLsRI/POOT3so/
hy0tBJSCzaK6iZaKpwAzERMfpgntd1bY7X8RK1ny42Qwz6WEbDvh4ALOWR6ACMfj
yy+e7lcLUsqtSRYz2W4ToWSyrXkxDjTT4sfB6ASZXMlTECPqqVqo4JdPTibK4rLC
u++FTtdf5ZC2NABGkZXKhNhbALp5DKsaW58PfFhpWHuy7x8EVoio9CaI6csmZj0F
SzZRdd3BP5Ndck4+sMPfGMtyTA0KgLymn86E3D1vBv0PJbwPDjebg+Vx47xAC9y4
qv6rbMQtV1n/1FU678SNhLG+qjG/icXyBUGOJANj2QkVCO5G8gczANKll1FtWGiI
u5i/qW+lyZ2RSXPiuap4CN844SOwpj1qUTHgKSyUReghvz9/2pfkiuFjgomoz8ep
+XhXUNEs1w91v73dRVjmAOtzu47S4pS3s7lkHsnoszqo26LkkVUbn3ip1vJOueiP
boOxLoSASD/Kpnc5WXhBl0Nghsw9U56CKaayvLWuJOMhP3xstUloOjHQXyD312zW
6cW2PnwaT+g1PKbk3JvqEBbbCh4hOYW6zCgzwrkSMD1rNRR13v0LE8vFCC+gdkLo
Adri0iFE11JoZttNxGX3g2z4vHvfihhGhqLtJ75NoCyeoGzWKyhN7FShhjCt033O
zP5ervXja8kGDSos1oKwMj73pLsjd/8aKhEBzVsf79hV+xpbdtefxFaej/pm4gIA
AQrkU15SZF87RsQDR5bcL5YLjzz1Igv/8x1YIhpJb6WNQk51ZpG9n2RtRAtC5V8y
EM1QTO+kEONcXIDtcjdCcrFzZEw8F3TDVBjs8zmUJM9YFfwe/xdXQV2FH/4U3gsB
twnEoYnaW/HkGdYlmHIsjwUsg0kC+2atXADHJHtZxQ40OW3Eu4xliXdWRgNPbJGe
Rjzlrfa/IIIjZkS1ozyBO6dbxwyshQOYGc74xJlYc7iSfe+otHuM7UsFQpHlYZlg
ICVLXtdsa+QPUaL8dBiFqqwqF+Fe8MOCN6A+3rjOP9ujBB2/3YNfb2B9tEQ3MERs
0TY9OMTu3NPqUE4TJPSpsib5Ep3tBLGkD5DjjFJBWDRcqjsyGRda8ZmUGxBYOBMb
9U4CVhVNcN/S7Amg4RR6JoReCLCJrQKvcocxTnGmU8F/lSxYwEsPK31qOaQ7Zb7o
Q7nPIhdEP6fjCKk4e89+XeYy80UGuMPYmH2tw30S4/z/w6aVz2GlgwsAQS858H60
ccMqAqMWHnGgB8V8RTXBm6T1py91JW2Y7XpAArbOucSTkUnHqnp1BNZ4rTjgQ3wK
f5IJTb+MaPM6t6uzQWaqi2tLaJUmwOgfA9XhReI5PqibaHNhXTvrk18SShzRVq9k
bA1tl/kRSB8zN2cvDf5s6LqXzqNMCHJLiOSJ2a6N3rqpTzKa38BfLlvYvEkjYigX
yjkyFPpJMQU/3bAztJh8c0crpcyZmr6fJ9j0z4Cjzr0NvOmC/fO+SgIGa06mXs25
vILiZly4jLrcriMAS7QVNjlWNuTvpOZYtw3ayHJEZJBy70b6BK7oKv9vhwZu+dPu
PyBJCWCQAqYzJ4Seoy3Dqfldwkn3ZeK8ulHKi2Yzx5HWl7kbfPJBTqdUIxiV70v8
dOVzmQM6iYkAL2kZmycI9WhM3XFFUp6FPWW9pkRqhFSXhkKzQpqJ/Kllwdy06zpe
av59FdzN0C6QOkGqS6GYcAphMLN0aVYd8M/O8NfDunBCXu91LJ+SzpPjNerzlVsZ
o14qlk+64Tb99ajSsThnYQaXrDI8Vb1N9X3uDjOSyfCIeB/5Wf1faNwb8W+gLxRO
l00Uqfrec3649FKQ8UyHOB7JKfPt0mI7bHVjCE+Z6Jsr2lr5N1YPPkUR2/PoQtpE
AjDFfgGHC1coBgiEhbSPENF7uRxb/XJ+L49+ohXTrevMk+v3I0KE26EdTi3KNVbM
pmMg2e+nihB7ZNu2ZbezPIaQZVCPLrGaiUKsx9RcfgY4oQ03zupi8urWTok4F/Q2
/KkvHf4VyW9r27r7+jOWTdUSfKKif+lif9Fan61Ys6mwDY7q/dxL8io04JAUZ17u
1qc8618cqybOzEHxslZMEQ/TLUcTR0KFRFpJF6RJ1moSDhBe8lB3+spl44B2tIUJ
ijTL83cJiPN8xL5PmYYLvrfG+rlOFyqxmhwGkipefMdh4NGlU1tW/N9nwzV4mSQ9
7OEyerbTfIZJeyr2wXcu7tBp8V0Vsbb16vYN+6oDO1sK93jrWSwD/rZsJ8XmPCC8
UvnXuEyBqWGmHXhR/DDxVkbsuD3Z9WDBdoJHGuXjopF68wnapokWqmy8piuIaQ6R
dPdeUiC3QvpddLCCVWq9oytee7q4WgC+E5dr5N3aodWCu413+5Q6lxQlKv1sg3RC
9PplhYUIHlNVfgeIvc+in8BvMo9DEEA6WkYv3r8tgB4vZ2BHtYMwT2p1OfTFxa5M
iUdVSmpzVD1Fq4IoKiHwC5G8RVTS9NYKieNgq3W2NJl/GSWz6UrD/EH6953zEF66
cOC+uOj9Z2UbpSdNiRBSz8Qz/vweBrisdX0mqi7tTAzD43P2rpZVh+D76Sl7Spk1
YPZDInxj6GCYUgaFVm/+uizKfy51xxUMksehogIjML5uF+4HMDDR2SmUwI/8VW4O
YxxGgEiwbZyJeOcJDsSQIyVwOFngZ6feRFw9K6MV2HwAz5D/onfVolhCKgjfDsFi
ehmMZsHxWf3etRNMD83q7RfMEokoZOPCshcz0FKE86ZL4SSYXLWgdkj1dQLiAVi0
nTcOPd/VGxgjMPf01IIPhoktZwdJXZGdhsVs2NZz4qh/8OThHFodaunArKZQm4U9
f4WXtgcSHtAgLYZQRNPtRj/C07vAczHBnNRmZzDIjWpAPCkz/qe42370CDlv7wdd
JRRh2z6JshWl24KQUgBgLFi9ffh+rbXrptzQtvj2vpQ6OLrZQc6aad28LYqu8xPo
44RHa+8axK3ujJ1WFxRz8A8IIcX+hRTLsXtenLXWn/oL7uBQXGttDZ1W9nS6yhuG
mqS3+G15ThUP5x6WVAAOz7Q6rTskKngJd+S6G2Dp4kAk68cJF3cVyeHA+PUZF2zJ
HqbSfqqGUj9UwCKyq5KIZTN1fKBFWlIPeWHLWPuqppenv34EUjbx4x5/u/I6cIxj
yd41tutyz5/bvhi1NgVCy0aom+Hwc1NfAJj1krsu0ZfsgtrMmpImD4IEY24GZwYM
4PXWF/JcOlJq44uHOuAv6Tg9aiMoGZKMU3TC46rbn8xWqO4itukF2NAal3Rw2TS0
EVnHSxB65oyd8RvKZAqokzx6g+6YsHVYZjG5YyIOwBbl3zjn7kaOK4mQm0PehCkw
41WWM6uFtfXME8V//fPvfD6Ht8ov3m9RXDgaxi/WRGulDA99QBn2hz1WWkbk7uFQ
yps+B7hDQ+w9sEDna+uMoOaJxl/zuOQSfHCWBj4eo0b61PVDVcUcRlTB7TwE+NM2
RuYlZ15LcNSNc8/Yij8z6wL3g2uWsogI34dSob/UrJMBHiGGj6eGPDVXtJAjYYpK
1LKYrTpj5HW9r33HchsVI1Tk8TgjB1tfszYTKNyysTGC0TArM5K0fgKVmrhrz+uZ
Y7tzLepOFsOn4m0wkZDzEMpwukE4oyxM8aK9axzg9rnVa5Gq+UOxxH7OZ48pq47G
SeP3rR+Wf2kVLozTVYpRIdRqRNEvuQ732gh1R4oN4hJaqBnEUikT3EecCMg8/Fk/
LuZ12LfAPYnIg7aGDihGqatLNdoXI0bqpCjVmYtlBWx4gNgBogIHeetgvv9Va8Q/
gG7g9CkFcS3rZUKsL24SU8ZCYUIqDFxxnLGb9E6aSMsnzQEyXSimQUgCS1/fsOZJ
9Qlvfa6WO/OH7L3lc905uAWAufQLclgxl0kyOCRNkUUsZZxW2T8UhxtM6Mc5+hrv
Sc2sKU0hUfdohCyDk5lk/oZx0aGxaJ0XHHfjS4PoaV3U1kFUXusEF4qmXfR568IY
/WmTB0XEhHWB0pS+UtWvKHXvKUZE20KeGNSsuU8k+RIL0xXtVJ70kWmNBN9PmPsf
F6/Z7Wc8aPZALehwGAGHGQSEHl56tIegN/697eHmFVczuvH5q4riTutcgQ/Kh8GR
zELWEtvOHWuOVFGWhjFIIumO0VP+LAnfvkLOpWGgAtqgxGWxUGfxk8tu34sz/3FT
0xFPJ1Dzodh37eleDrrpYWzhhJ+mtL5KiiTaxLSd//+rym4iWRohPA+D9OstmHE4
70e5Uhn+o3UkBc9tJtmjDP8Q/0o7sRcwgwZKMVvXQjXb7B72UNNbRFByFv50EChU
cZcBH9TUu2u3OfvA0B/Z8ESd8Ps+OglsnDi74Jh8g1MbVoEgjOG6lcq0v6v2HQ+V
fuFyatWI2+6lU11+a10M5UYC8mYqgwC/UBUoSDRT/fP2Yv5iA5NqSmxO9RNj1m3i
5xX6FUYq8RddtJjtBm3pZuI94NRIa8Uto1diSlznQmi3FnaNhjji4SZ9xLyH9qQ7
5kS08/HfKZmH70B0cYOedzfV24KEN0OaXxw6TeX1yeFpYNbtC98jMicdoXanucHl
5uNpueOG1XMzE/b1fMxfk8COVfSLlxbSuDtT6w2q5Op3sE6cGV+YD1jqRJgJFp25
J0Z1LfqQQFp5e7GUWsUOCZXakpetVfYvDIZJXzIzQGjbPe8/ZQwHhWMiMHgIeWCb
+5LqN8RTm/6IYTAKxOBUBXE74CbRlgiaPn0MS5j1RXcfSNN7aok3nETzYUEDDzA1
WkomLQTN4uVa3vp0FNRoM6pe8izAY7myxu5b6lw5lh32VG7FsS+Gs3ApozdiyqIt
V9uymRb0bgb5iyeFCT3KODMLv+FxwxdtHh941RsJQl1Z0vCZN4B6gkndjmAXy/Hi
aBfH/ta6+F/YUWYk4807RdUaD0PmNYSsD0gIOGVNwI83mwMLfVEm8/iH/7QjzCAm
9TW+NdPf756kSAOeOj4xxrqyyX5trzbW7vtg9s5X2ttYPT0cUBSZ8KNavPlLjn9Y
WlfYVV/ZhsvH6c7H4X8htGEYyKF9B3E44wv4U0UX/Dh0jmhldx8ShBQO5ZhUD45V
gSB7Le8cQkrTxBp8YIHcvMKUOeIIqwvUW2T7UkktRkel5VBArcTEbLfc+sZ61gQo
uOVAdGh+jUali/qw84h1JUTqc9U/7/A3kB8tlyEq0mk5eqYBPr58yeMcF+db4Dhk
O2x8Lnr3GBfWh9eulimrBElykDZhIPSh9dlWkIHLsnis5gVGjIx5/P8xjukCZ2Re
XLnREKDHOh01FiFIcXxzuRaBVS+pnANNaD6W+lup18Ho9tnMb7Tx21eimxfFd3X3
ky/6NKDogqX0sb/rsdnQOqR8SZnSO85TvKXG3KnZN0EK+P0o+stWxmnGBuF4EzYz
6SGqkBJuB6Lh1fcr6PDAJmDNYJkyMT2hfYgOREyl0HvsZRodeygAnb3SIL6B0/dm
/aKk/ewIQkXJP5vp81NGtVnRBHWBUe3RCLJyh13AOQxM0ZvnCcxBzSITVtP8UHOv
7bZVX2mXx4SJM2ewkJVmm6QlISxavY4Pq/4QUlotQzU86HQWevbJwKtH0dJWbjuM
ptYwcuUkzqF2XoCv++jvHkr8bnefzkqOB6bp8neaOSwwsk78e6H4jdGkGObDrx66
LXR5YLGRTUOH30i271C/vEOrzQEVayLje/nDprHE0o6Gks9U34/wOFb1VccwxYFj
qk01o54bqtJS/54lMxr/0yXroqTUi57FtW2LL2aE7cFSRPFwb1RMBioxlMmhmLLb
HVlC2Qj4Y7vgfU4lgglw5u+zJMT02ljGSaOE3mJDSg12F4FF0HI9f3fTBdVXEMxC
SktB+Zo7gTzd+3fXPhNadeumhcDuXVdrKR2ZPVMuKKSkCD+EVJ0RepoGAukX8Bog
S6ORXBippFtkYvnCwN7ZLMsloA8LmolfZINnBeEyMDYUZHuYe2BBOmReXatsRn3P
bRokXE+jvXzX3nCUvVpKndxK37fyuZBmN8hQUHUmD6sO3tLhAVqrs1hlDDyyr4AI
c7pmjILDHpgU/Bjawaq8erDlBqd4Z+lsg3Np2p+x+vQcTzE9gP6GiLpzWbVHKjp4
Ba/13dafFJLh0tzZVB3Qf+vY2v17qRwsSprHuahJNtjiQcfrN521Z4xe/3XJTuFD
yHwVYc/5AkwKJFsqro8ZFOH4kB/zJvL3Zp1PRIHm1iu8JdI2Ebiwxfj4hGnaeede
H6YpKjrCoYxMrDfhWuVxGER2NxGVhWP1UcedUDqmO7mKKz+ahORxACBHXMPEee5a
ugIE7xrfvka6SCoOCHOyOKeUbBefYDTrgmXTWS24mxaKY8QuC/+mE2cV8wkGQbNU
rwjic/0O6Oni1yE9z8YZGpgkXFLRPYEsPJE5Ao+a27IrymJbw6PJ0haneNuXe9f2
o8KD2fadkWdsUCffCRoAVknkX8MXIbSwkNRGemsS7SmPGDlyqmqxTZUE0BOCqhKb
3CJi/b9GvbTSaRldFxE1qDCoTFtVnliB/kI/+zZ7QQ7t9RUTyFxj9MznG4jyz1LY
q8E1ybaQYVaYJmYEa3vgUZD1Ie309mPcwtL57hFlH+Tss8bbwrFsDeEYxpjNHG4C
okSpRH9BVP8kI7xSZBhSKH3b73jSTgQZEsPXwMCuEdkcvL0pJmTzLhKXxo83+LAD
dhfANKh/pWoY0V+Ze9wq1O7pHq0HvsCHoDyAX4wade5HtJ6A1vaQpP6MufKOU3yw
wzUGmr++tFOAiC3Wu5Id3+DSp8H4DuYVrtsv/1niSMfY9UWp3nGSD7dJ3olON2kR
whFM97jhS03Xnab29wVRjH5lVIoxU0gYgsRo3q6yDAPeNHwz4jIMAYInIxIS/h/y
XeVynLCUS8FELMYXbQ486CZRuNqKqv+kFSv5Ny0pcvFv1GxRzxKMj2JTZ/axUw+j
/5h/3w9qr1ZsKkVhdAP121pV8DOnkcJJTkSB2STN44frebD2v4cr0QHPVRQ1z+ht
XLncvzCSJhWvfRXtj18kTgTacm9iWFgHL7T/8U7ssXTS5FP6wQI3DPkTA7Ee384T
RLU5P+X5OCfF8xlwmTTjsy7MElQSlxWAzrcjr0ZUg02dVZ5IkOZ4SumjaVoCXV7t
ZsftNDawWwPlOXcukU6OQ8F4hny8Lhcl+cRiQERKHHGUqbBWRWgjCVBZL6S6zV2C
U+8r6Ymx7AihYL68VTfOj8GkBkelVjjO0lIZVSPbH+kTqtYoVsRU05uPSU7prKgD
PwhtteC7JCDTKjyBGdzly4YLpj2U3hoKY+ooHOp0JYXQ7f9T1JKxmsXrxNKtywAT
Wu4dE0KTBvMx+Rn0+Gf6xssiXBkPOqclOuRH/PndRzAJrmFO5A66ZeefpnQ49crP
+MU3swtAf8tGiVyO9+bviJ51tPGcZocDPMnxjuOUruArsmGUK5aWto20T6tL/7oW
2ZTR4Y+1tnf297xxcVdfuj6ScgnaVJKCi1f6OYqubub5PzS8//UE41cCX9QNXMhi
ebFchHrh0fSqKbdLD5JrpGc8C9X51Nrx5sveWoF/4oKR7J66+9+Eco8I9Ul1+u+N
KW1kZ+7HDpcj35wScPKISz7uBUFQNnxBLnjS8AAFlbOLyqWMUSaiuY4U3m7fI86+
sWKfsSxuk4SdwNaP6/0Rysd1Du7HQUOav2q3GlOK0wSiz2jsLmjIZYtvUBEZMaPl
R++RZZGrIRe3PmMtLzThQTYeyNMygLLQQ5D3XwJHxHOKNhWM4wm9kuVatBwTNXbe
eqpwjTJx/R5nTYbWSpM9gSQN97+N+41BW4MlQbvnFYC+ztK7QGyvpk4JxL0w+xZ6
kr98nbpXdqOpegKoWjv75WdvT39WwQslsyXV206I6zvY+pbp3zUlL60oA6XZUHoP
0yN9SMMs5huuGU1EfNgKV3LOGiJnoxrJdn/zxOdiAb5YqLF+8ebf9pmXm6NEI4HQ
S9kCMDHzd3NTL/U6yP8lR+tXQUND8D9j+dlbcocRES72C1OmEEdAwH8G5mhI9bTV
oCcWkvpZ8rZHKaKfDFqwcRDA+fgvBVuZ5g1y0r5x25wwfrP1JdoaF0McCZ+g+beu
EdNeFrmMHCNIJ0aNqS5Ss5apV1M60GfNP+9mVs2gsnTpCCx7dWEUQN/eC8Gu4Iys
OzTcbMweIPV2W7nFpG5VG71v5gnAdTmDS2jHfTQoz332rHmITSpwojdzFQPmUysH
UWD4R+cgY+oV6Wz+Lw5BzOyZDH1mjukrlPox2qP6YbIeHaWuI+2vUQXpaq/qfX5B
i5qWy4ESPRMF7rTKM3wayfPDa0VBooetQXaAKPxdNkpjDBJN7/yJIIWB40ln8yg0
jwxEZKEIPF7nlAvk9duuWSECj1+AXptxqJ8sXiN2B+gbc3OHudoPZOlb1Nqz9Swr
0u4qoovJji+ZVW8x61ERDxkGvxVKbwymJuu+ung0uVWRNziN0sVInSW7s3PD2vuS
GyQGHJO18gHO+Tab789fEIzpDroHd+CRm6Vi/YeA2GCrZUYXY5GxXPX07MuGm1s5
09JcDo1V758bc/SXlfZ/XIRMdotyKLoiNaLa15KdQ3Es8Qn34QRrJE9ti+CnT2xc
tDpvgKZPZZGFqALImcuZsPksTYguiYYQkXBX9xE8zuN4CqjDBxPiex0IF5lMtDNF
x8nhiBNUeaDIdBqI+ITKTkqwzZtxr5KZHgCe4CcXwdaszKVeNtSEwP33Zz+5D6Su
lMXMuYkunJqXfTlyiyQpJLKWwhuk8G/s19qZEt9I3zDib4Yh2ZOaoqrI8Wmg0BcO
QH7jxG40PcOA9CAvuUlfEFFMZw3eVkxmmg5stBzmzyIwIvuyLO2O3ZsAbkp7Scse
uIHWXEY2agh9TcjHKm1n65xCj2CnYRPCUEEdzFD7AxBbuXffX0N/E1Kvaixw8cxN
yvBj+fNGIdLAVFmc9OjOQlblKjtQLJffieGKIg656n/gSuJfQQ8zE3m5Kjx0Vrzu
QKhOUkS1oBG58EAX+GLZi0YZq/aHjyCY3gj/Ah6sB2dewPzbpLw5qjB+LwfqNVm1
SiQI/668dYAoWhNaqzl6kULwQyRDG4wnAHxkNHgiDSZ9LPLefwhauINbjBTrK9hB
5wjEXzOiD28Nj8tKBx3E3Z9+FUqBxS4mIOjTdboJFnaVfwHBNnWTVMnvOdLrNEgU
4MsSv0v7wumzApgbSpk4WbjIONOZ2tF/nKA7s14/DuV2mWCI3gyrce2d1vJf08+j
PKaVVciLixChz7Ahm22zqv9l8OFnl1kXjFpf4PkrgikeiUb+V8uuh1e/geOfbEB0
/O/nRWvWThpTokItCVzSJsN+4SqNBv/I0Y+B5UV3I2E86RPU9PGXicDRT+oFfX3+
fffuy0QyanPnSmzGjltx2IcvdOhBPu8hz8W7sBObtaaXqOQbEv3NRTub3/+CxzM0
+8+/pcUoB4EXkDvGBFdLzbJ1XIBoWEqF29OXF+2GWm3V+O+SXgw+wcLbzQzZfdgd
HTUTpcqEI4GqPpkh0oY2X3s4NGTUqEAQvipkWMGa79FUs0COJOyxpp9mZQKr7u4T
GpuKSHOv60YkGFZVMMqwwmJ+iSngw5/govxBFuFil34Iq+plIcfF4AQTNTofWbl3
GLa30835g3RCWuBEaJ1fy0js8eGH4IsU0QY3l6loaJYPrCNufaL2CcJmKdaCQkk8
wn/8PNG4SKROAhdaU15ALXpTftzEEggsAW4scemKLq+C0IL4Un2inQjPGM4EfJSq
E3HjKAiFFZC8baauewAKFXPz0m3N9Yc2jMixKAZEeIGtS0bOaz6CLmL+gIIyb9pg
Ll+81SQDg8srmYzFOL+qkodgOK8qpbBkXWNyIOjAyIWdeAemseTzvnRsinJ7Vf3L
oMI+2g2jsscyRBwRsFRq6M5d1YovTkadjNkR9hXH0lcN+46i7BrZHX0CsWac7ARI
T04F+ARjB/lWEHx4rMQDjdkGpsICxWZq8IynIS8Vdh+XRA9UMZ7Jf20qndodRxMV
SKTqbkhDyBZMjesMYL4z4HBLAzGC/bm1QdwfKrIW+btlmefi1D2ni5DGVlSynhWw
JPO1KuS6527sxF7I81ahNhPCpY4Pwqy3Q6BEbo0Ehxvv1Mf27vsdNuA/V91RIFMj
O9+Oo7djkXwuPUgui9zGCbGSa/qqYqoo5uE9VRtkZRMxXEw6jm5vxRJ/aVUZD3bd
ajiaHSsbFoNs3x2sJIxi+8E8yQiKcAhYalelyO7acYVi0UcCtWzd/xWwhLEaUznz
TvLqjx9Tw6WHV+nutOHIx2KoBal2BHcPq+lDkW+o/gTzZ04f7FSrjHoK7BDJ8XHL
wOfxQ1tpYGJtOMQyjWiTVhCcbk24PeztHHeBfC7qsTSQbapTsDhpsFt3qW1RDc8a
VVo46SMCqJ25Ek2kEJ/0/EU4MBvZsQ74sod3B6zJkoykU43OHEs/hnKkUrOX5qRQ
Pmo0akBNCD7DksQe08hwLQBNyvcBvKX4kFsBgaYTXziYHUm5MTmVycu0DSWa2ro0
h9MrclPboIXC5OGgKeAdAhN3ctnKo/EI6+24cfzT5R26UsIxtDg2yD/ZZiYzPuxI
/Eps4WXLXx/Vg8ezZouQr8UX2QnknEQIEMfQXi2L/NGptFd7T15Di5+8QBoRVxbf
Okl42Oki8WI1bXs6xV+q2cIXKWr6e1IelWGmEDFyiXpY82ayNAHICFEN1CNp1ZVD
T+RpAk+5rDqarCGPp0UV4NUu1A2tjRaweGw3CeoO/BhRYZUBGIj8fbmYA7uL+7sl
62zvchUHAshRBHA8GnTVFjlbFHPMFz4et8qWWNp8gE3uP1mQANDrQFKr4OVwCqEv
RP7lBwLIG4QsN41a3PLwcetMbh7scykd4leCNcu63fZjvLWuHRdE+DWxsEnY7ykf
uJR9Dg3+HwxW5LiDlaJbL2oBiJyTn5GLjP6gbDulP4AHn8PHSzxV/kxILLqg5UXG
MpIJiDfm4Q4ME9cTLo5UkaGpp+A8r75n1Y0NHAOscYxRcmncGPkT8mLe5am4aSyG
RREbaQvlHXa+X7FB02gp4iCkpraLmQ9Aisbvx60J/fRO3RAc+FmPh4oDRdgEA6vx
GkLsKOezeClI7CGF9iWZijsU07b3/gw8DU7EAPNCm6o36ra9EQqhqNDY5Tb9ZlHV
mVoq8cM8Ofx5KQ88RErWXa5PImqjNLIiQiU5+rsWBYostn+xVk8wBsGbDtAbc3t5
nWMpB6gkbJT1GBQlLcCWPyA40MEmnQdobBg9XZmwbI/dq1uYIamqJoctvR52dfmo
OgDNTAGqaQAqYnjtuwaK6QL9S9FJazy7p2z0yCgo9fgFGUN9p/Dq8FQ7mhJtCwJJ
XiTx4JEmNujgr1JZmJFF4/mCtxftgPNJ4r+tlN62jKUrv/gmKUem7iswlqqtq2xe
vSrW4JZw0Xr9L0g7RP16YAeuO1V6yz10w7Db1p9pfD5W0s7XDDd5ZT5BkhuRRPAD
H0054FbSvtUOB+525i1Lusxtwd2XOJMCUtuy7HHbaxl1QKiHef6NkwEU/xW5ILcj
hUrA6LFEvZrqcpauRbslaztTOTdOyC4d6IvZiZezNpXyB4X28Zpz61NHWOMVSY7s
cfImbVKbIIEnzPAiTkO8iFTKyH/S2gtxIAMQiuxGHpD6Cshh36J+YC5yWjuO44Tv
dmOclOZ2bsWv6MpvNxHdIEmcQo7sA5yU24ytVsIfm0C9eXNHyg/uRP4NWonp+8P8
rQPBttC/HQ9j+XqO+oloMXgcsR5TCtii1w4sDS97XFJI2w8fpxwPLoIu5+I8ha5V
oP9iHTrWA3Q1J4gZxg8mv/uDoJWq+ePCq0ovYd5mZaE01rwZBZ/oUkg3p5C8fR+a
dwfFjzgPHVU6LYlJKLC1ep6lu4Azo9qDcO9o3LBoGVzteo77vPVV8SFwJIKRQogQ
HdPOa/QTBSRw1EQHAhcGxcUQ52MCw/jGpFJP9I+LPAk8dLrUSsB1UKXehHm+Rnr2
o8fkTkdU95qBHJOVc1tvcdqz1azqgvQiPov/YkBaH+i0yleM3RltNYGnSbR/nRx0
zzu9D6vkSROjcxhPj2FRWIVeVVpFdBc2iJMkvz6RvVwrpOfpo7xS0Y6Y2TmeBWAh
vMBsvA2kz8tnMGYxhZugWOwmuF7YnB49GVA0udsVo8WG5k7q+VF2tGjazyPEin0f
AZbTNI20Z3uJkeV6nfNctDNSCrVMXepCgcLXTgT9BBoVSRV3a1jrMcwJrezbFjGG
nfX8jSlAFMfcPfsxh8XwguNLuGRJl5eOHaSilejaCNpTLbesvQC+hdiJ8Rh9/p+J
O6W+2asfp8v043SypDX0TQLZRUTh60NvbvoyPz231/bH1qTOeT74Ts3n3+M6QWcc
qwW22l+62KhNiuvJBt0NPBjyDofo1U3nFTdX6FtouTAJQlcM53uRuEIoFkyUWwmp
hbpVCYxWYQPWcP2Nra4KBXHKcdYS3AhIfD0lMo9CuqNk4ylmD10yagJr/f3OJV9K
1LgSQtSMzyYgXmDNsVaIyUBQGAmI7WfbwmlW80M7lLU40dBPmNwslSFsJDKW3Hpp
8VOdEIEQI4L1m6P8XJe4tlBXtzX+t6ZUqMwOOCmGc6/T6ywTCml7y2JvCPosx8DD
NMSIVCrACx9hRncHqoJoAI6WylmZZt78LH3azy4MNxeNXuPT3k0FnCmxKEbNVxff
YkeTNJkVOZxheXsDPlGfC3EdB63StGorA5R/+XKwMjKFjsFjaka3FxWlWxfGDSFc
LbFLZRVA9g10USfNGtiFiR6DcOqkzm0AKAqQ18QdWmWmAi2fzyCBZ+YCzzPXyWcl
S+A86ssGLkYfTqcK8cjLnoqM8pLq8ZFscLb4G6Lbzah/upMj7H/iAucjy0CuIAgN
hSmS8q00yZOXRjX/wakoe7TLJvh9IlHtZIn6x0z3qhrlrCbqudJozBcILsqlOQfD
2y1R0aHzdUZanv1ispJDmZZgfUh8Kz3RSRv+TB3ZNWWcIh2OUI9vfTU+0Lb7VhsT
R+b+5r8Dr6ReNiJ2NhjyC9VJf+o3LekggbIaI/hDTlIdqqo1Vi2H61IKbJoMpEuy
kOti6Vg8tL4Vgu22i194V+EB9A2JQ0Ah3xzlx0YQMtGwCajkXO1NLq50SGwveIDp
kyg/5K0sBeKOfctB7JqsEp8vgerdLxzqtgs0lV8wE1cdbbz2r1DpXlD1fNG7KdpA
tKXmkjcdwJw1eSz3FyRVu42BnitCbxSt7ScJaIFskq2HcmwGe6JLNu3679J8YbBl
Xep1EaFrYAHvjoWB3nrWoj9Ph84zh23+2uTY5Ai/pr1+aqLLO9solTSQEDueB3uK
t6pYv/oSgNBF4h0r4iLYe0eLeY7BmPnkMR1lXtvIJQfIiXM9I7vSEqlg660VusZA
lCAPkGjJ77Piv6AybzgZu1EEKMIX5G3sj52FzbB8d34CQuZUnIrdrEgfMLgcsf70
2ats2NoKfxQW7cKRCRV47NwNtx/Sgfi7WtHC/KgjNG0fa1lZ3E/7Wwamymedw74F
R2shpZHxQBCgdAmg+shQ/YZC1hAo7sEGecSARAA7flwKo2RyYiM8kyuQ2y3TMzLw
RR4wP6kSXzIMs+iIkjKtzQp9cKFN2+6OgWCbBqWlMf85ldjvCkehYJIdSt59YANM
W3qytfsn4KNZKQGYqmUqrqTbiTpoNEFiuJ4Y+FSG+J2XKiZKfVRG+qOclwa3n1EX
qS5KnSqS+tpJo4KOY5cVQHYM07baEY10n3PQzHPr4diQYHJ9oC7E/B7/UJ6xHGCP
3GTKxtju5nRoldKnLqKVPKjOtLc72fpyKFGS2itLXjkQltooAR/4oATCXXSv3MIC
d6I+/OnX33GJS6kCOA59BRrp++TtS1+fJeTijbvQfHYxf06yzFq3sPoX/MvX3mhP
APvBfcXdXu55O4T0N+f9HXkMdTM+yIvweEq6BBIz2f/0DCiOaRBEASZUVdbT1aS4
0d4gs92yc6z9X8C0Iks5RGCJaRlmo5Ckv6CQ/PoDX6IY469xBYAX87uCtIV34vW4
7cBelcMlbewmqBSzbbK+fbrIHDC9zC1tOId4Y2NoUf7Mm7UwdIpyFPzj5P0FRyV/
50rRBYn0eyaWgpHYv4eVkLmXsuNUTrjzxneHuoWxCqVu03nS+DRuCmr8DGdouzRv
Hc3uPAst53zteVDH5/0NQrO2RGJRrmkaITX9iHDOCzOt1RbHF6x9Tl/6tq8pf3y/
b4iPeUAlSzrZe98TzLYQFbTpgLXA1Oiz7QZ9xyXiSDasSwABC7VBNVuy7Hmb3Yj8
IQJuFigl/1XyRJrpGee2xCHGxv2BHWcqyFTjr/031NFf8zPOXCmwVGN3vrpAEMfU
zLAGVtikf7JfH142R+ZVQoE7oXQ2XyH5C3z4Sps0hAFkfjBDjLU9bAWNvFRy5AUd
8PTX//TrXaNQzxDYVz6peBp7qhcXMEJt91fl1H8FaA50zV9X8YJa3N5qnJu/M0aR
1dwg5SVWWzSDeAInO4+9I4chDTs9EFMZDRoIlfw4ya8UP5dPNyZv3wqq5oZKD20G
pMedp5UgTuoK7dnypwwoUnNwrjDsi+Z59CorFx7quPdZLDuxk8mouuQ8KTnWCXR1
m3pvFlOeP1FTWXIONVgVS4te5oD7Npz7cVH68+B/KvspAGPUNN1gVtqALurnFm/i
r7hN3pdjOPatC66HQjq8/Q9LRzN8fzVopngUrALt+dI2qJqJTYeC9qQWiiEz6X81
v7Jn+nVE8YD7OILrrYOzoPkLfSz/Ls8dNskxk+jX6n8g8KZTuQlNFAFvtoCwCGTb
bXR27Njik3LSDykV7Envo4rdWbn20nZ4O2fKDkzmYNeRPtJcmAvkI2U2TsKQxjRK
Dn3NqZtSzMwH9Do8Au3YIwhl/NbLEvCokCYWwIK7bt+IpoYwMw9cwcVNR/kv/2T9
RzK5VATjC+0n3pfwnzMbHljzWk78IvoYlI+CcMls7Da56A31BQ9qpYqJk7PYQAKZ
R1PyajPILc9xLLiOu48//6NugokuqaG4YykVoE5tQAcksn4CZWpm60ZkgLeKdzCi
HkQ0tugUHZaaNMgQrfqT1IkIjW3z3zSkHJLmrrHEeXYLlBB4JvaMaGbzmOARxSQs
AiL0895/QauVJn98qcALrI+gk2qUZ/UrlVXjDpGxGZlsGGUju3x9muX1ownBYNP7
8vA+ljF1T0uu4mpbB2ilZTJ7mCdCx4Ns1VNK/slfkK+L/tT+j+LYO6Laa/xKvcaP
Vko5x7QKrfb7iZP2P9oOri3TZuEs9M30uvbo/xHickTk2PCVcs5uP6ctSJFJnM00
4v4q1cgiLbJaL0yw3GEMiU/+gBVlEhh3plHmcCAYPjsGn42WMfk24lVZbaNFzgbB
ccFM9MtLDZxGobURHqGoWLgE7+GqxaZ2REvqcGmMiIMdEM7RyGdf9qPQVdzw4ShR
cUcHBM5jc3Cd8m0bjRG0X8JnWlbRJ8SKDlKUvfVMIMSgYRS/WlKXHKH1IKRD214k
QultRd7EnmQsr9h1by3UXr05mLQfkC6w5fGW56WpZpdrsWIvpX+WUrOC0+jTAcZE
vcL2kYSyrhTxsFRyas2arhSO6dG7z5FD6mNeqnD1CuQF7b6RT1t7pEADghbDbQS2
Ta/fl05X5pwUjdBtD4duyZ/YKv9Hk8OM4C6RFXRRTbsmlyrANGSOESh1DhsLP8q1
s5EEqvdUzzgUlu3TG0V8ZqER2/fIA3GpZE11K9REHTx2wKK3tI7JgGB5jZ4Yo01p
/GhXICO32LPFrZTXJeBkNoeAiNf0h+Ufiy2oNmlQ8UdtzXNzMXzbc0qM39A4qKiD
H4MrDm7phSkFkTZxncDwk3aXKwjavdn8BNyeAmsFr7rY5fdU/x6+J3nAV1YenDv2
l8RKBsFdee0PrwBHu9RBa6g2VKrbSecg43AgYehmBPS+A6yABtYJ6N8C8Yrr3W2G
vDp+4FmY3emgOv9ATL4SDSg171bX3vxPkMibuNM2lKQlp6CDwORjmxw+fPcp6IdE
Sa83gKHFBE2HAhWxy68cqJtqi8dKWTj6WX0rUBDL4v2WbB6/wZJuiHTsMDVEhI7A
KXIDwMylUuu/CVdQvTROTbvyuIvWX3w+cYzJCtXm5SbyzyTcYCG1ldDykYNrcze3
70kiObDDYqyqzhf1mkXgx7l43IrHyu97inwQadtTDAN8GwCYq+yj/6TLy2NgsUzA
BVwc6YaDLb5NZFjg3hTssYza5K+/ytOEv2ox9uWDHcSxfZpfKB2riGAqKi+W8LZ5
+Ozt1Z/L05o8lVoAJlciMT2q3y8JZLzJovnzH+mz9BncClQ6QXLf8n76b6WZsv1z
3hdn7O/LM1rQ074yxeQz55t8y5LD6PRWSfMqJNI0vudqrRRHvYo8xaaBc7AFVQ7X
1PstEt/j+NiBLtfNrgujxMMgpsCZxKd7SgHvQOFFUPOn8gWGWL4qiSdWl5LD7FCh
D4mF7SVGvQIvwHQxP7wO8H2WTtdrUxpXzK4fuZZogPLa3tJ26dxGIxpFcEZ2EGXX
zXOaRuEF/71SftubQ8NI353AjaUdyaNob9Py6ekPHZ6Ui74UiJsXXy6Xvav/Tw+9
dAsFrFCxw1p5NUZuHqC05X2Zk5VdFEvG1gZsWPyC4kqXZO17+ztwkFac13hXLW3u
RySXUDy9kL5ZXs8Lt42t02xtgHozb+2nYyOWQb9Fb8OIgUdUI1CrW2zPE72Pe66K
BJJ8S8PtPvsmCGy+g3D8I/vvKq3+LQMs/i+2J9a1Ej2KctQRP8xB2WdRXB9ifJLw
8h60CqgBFf4CZm4Fu12DJnl+vE8PXgEF1VeLqg0YsGRSDIzCBvEKlQTjoe5Yu6+H
Wk86kZOXdp4EI0CJWMvv9NTXAgtmKogGmt/GDwo8efIHLaccXNSI4v5RMCPSylMG
pLO3Wi8C9j9PPLwZCGLWqlEIXKZEoRvDvHBgkTRWa6BKYqs1ZKjOvydAnC83tXgR
hgaLKGQd35fn5o89ONCwBg2/nRfjrZ/b0ksi+Ufwyxzi2X99+wTUlHU+ENZYRKnw
/nPP+hsa0kZZmxjUE7Qdz2ArXw1UaiKGZpd640TGcryPhJz4cljquQGfZnOgaW4m
sf7fMSCGtL+iVKp8WSI7eHFJ+HO1IiclRAmZFIU/ZRFZDexO2kHHd5TY7u3WHshL
3fKPRgljqKluTGssOKCx/dnQ8YPB3x9ztXJpfLAFj2ixU0U7Q4ZQtS6abMowOQLz
uX2m8N43GhGAgqDIeJZIjWLAPJzuTj9+AFIKmVALTNo70PVlMsGTfqF54Tw9F+y3
5aci27/vVwTDAhuMqkYzt3UQmaTlMHcNMXxblFEZQDv+GInKeEVWSQ4A/Q9C25ut
LOGkyU2aN5v+KMfQxqfwrQds/zmtdTrLfA3dzxYWHkcWXv27gal5dkYh1FClRfbF
25TLoGnDCAwbL87PAvpPQuf+QADWwbwOWaTrXI78QNkhg+55T4b8Js3o3i1JjnsT
jGFm6fo9UfuacHOExumFVOzSrIisbEV3iRBOkPL5hRsitpLEwlaWFCzHGcwYWzOZ
T0/m64Km5xxmkqxYxqWoqa2mQV5oODAH38In0ydwXiySvKWHqQYUDnfLmnBOR0lW
nkIGZT1RzPht8suh2/OkgAf6iKeLo/Nv3sJQ7Lg90kjW9ZiWpFKFSzT7SCvc3nfG
1tEACccRKm9Lk+PjQ1M3u2OoVeH/F0vSvDpAylMmWmfOIP9cEvK3ycdmPkwxyYu2
SUk8/HqU2raeuFuUjkQ5u+Y+ZYZTZsv7yKQx/Qv6oMablLzhMo17EAZF3853C/z9
g2bGPynnOdqcarGFRlwnnYINrYzXVz6alF7g1rF/vmfY5Dp3xCLLvbzwqjwnBdRs
heaA0Pyfs3YWVnvPN64QO/AxdKq7znyUsYRw9ico9Uhz3Fs2Iw9JoTQBxqvMKDNN
uU53VwcWEU+Dz0Z/Hze3sho/2D06VY5x3IIOP44StBHHCAcvQQeT9J1g5RVAhkud
lQY+Vz+5qFIVC0aXkJQ09PPIdyUwNFLD7jQhrR0pXCvJXSvoFtwzx81jDX3aQfXU
Pw/LlpCqlhU4lpBCSHGqjknZM3gVzTPWyjcC/BPuiKHXr0bWwwVqzNeXhVS0Au+K
yA+LTykh5U9oqP52SVQ+D6v7FVZ+uh4wWwcJkcShev6bh7TTvwwFlpY4JjJN1rvq
swANWIpnxO/xVp1yNG/gHQqUz0J7V+helYHnAeOX9DL7i+jROwxJYhT7otFIWl9e
hDNQ7MEVxTEl/qt2eRcCYH7dZm5ske82YFLr5xHq1jO7lScagE9qBg70Rt+Cr52J
t9gYX1oDhX/rUBMg+Z9G6cCHlioJmuwKFoXS/zcLaHBCTXWKWJ9PlHh5oLe4sgpt
9m0kW0beUS+kELp/2nkrqUXpoNNMeilrNwzO3BLVSYXpnJ4AUme5ohFlJx2w8iPr
cVwzQsxS8rBFFHi7v7DgWWayoMNAdJVYWnquppky9VTwxQjTys8D06f+Fzc88bcZ
piRQ0HxFbIm49wcLbnZSC+C6sBnq1Rdy88lkDbr0wFUpDHcvrAJ0MXWdIQBKb8B4
S2v3Wl6axPjJc+Lbqa0KGxq6QvAxqjCUGYvIzwEgIPWmD2YK2F524yyDUkw3kV/b
dNL0BAlBA8si/l4vnVKmClP0vmcJGudhPs/kybc7U5SgGHWvfryer7Mbf7onxrvU
VGaRJY267yXP4nPOntJn0x33XiEelpP2eLDmF5Wilem261NauPhMv9GGJJ0tKoLX
4kIgw4PCbYLufD8tCEyIDds4LV7tuhWjpgajPq8DUrJunvNbLocRtV88UgLsTd6Z
fhAVUbHLWZMmbPNC1NnYgrRlU4VmYBChp2FextPSIoQmFE1x4dhwQffPFjs2oMQo
O0EjpyrxQhGZRu02ezcOjkvUYkCOZV1yoBOxcW6q4lQDWNoO2u5IqQpobgymObF+
6D0j1ES1TEFME2SuBBoaFcAyrdO6/tWib2kcfC+xKHThL6DQsnjoRSRi3Ci0feZY
OE6XeHQZhu1/IGMCSmJvTlsMfnmo0f3xITFehn8erPxI3PRjuTTDdPdYjYMfc9s/
B6q8KJF3IIv3i+PZ4+gGn4zCzN1qwxsW/PsmMaoUM88ApgXRGOoA09Z5qaw08Nea
O1quDTf8LeMIAHG/qzEKEnZenS7VdqL/EtPnZYUJSlSHf1546giOF4GNLSpPUCXC
96vcrninabGzJ5xB3eHLh3lj/FzZ6TgbgEw+Harhbl2tnOONY7nC0yQe1j0TgIWx
kbJGAUIPKSInkb0ii2cvVMczy0iIVMKTJlRuISzywWxaZNy159gSk8OgtQAzIobg
q9zcnuvQIS4KbUFk7apiS6MkxH93UmA8Cf2pXkoRe1tYHzMnliCOKHTD4b8AedL2
G+IPlsp7dAOYvbayqwvZ+jGTJUGv9Js8SBFTR0Ys8cVy1NZgwCRG3gV3jwM0zSm4
jvxoNqRprF98LZPUkfR3Vxo5JL7MZfQkKqp+c8+99ksvNyDQHAGcWLaUv3yqpB8D
LU1/nEhbbtlHY0szc1tnPaAWEJwwAzv09LR3TMD7HNGgdhFo2dxjVchpJN3xAOpb
culL6mqaqyR2ofQdNxdXmZG07DRWerJfW5OF8VRynaEmND5rhc6MIhIUavTcD5h+
mtpustjwcc2KpfwbcjB0lbLWR2L5wqWpAaXCLo+wVPA+45bTZw7JsqVMmoiMCy7p
/k5QdhlBdpezOz5tNGApeUFBHhDTQa/tF1z6eHNiH95s8KDKF1hGFUraj/6oUe4r
xPvdfN3ORf522q9/W05a0I6CAjgPLr092jBDzSb4VwsZSP/DJQrnu8oKAVjpQGyS
INm3zSYrR3ohr/nou7MGHLCDABNZzCWgqnZ3V+9ltZ/v9qm00CNeCaQ4ERyxgV+V
ZgksybPI9ypeZ1HKRj3aK1uYSUci2g9aajkwrvbAIV9T9T52zun1l1BweYLJLVsc
PQwn+4jOmsG/Tx+qrAp07AIePmzjI8Zp+TNAANQIIAzjF7fNbXS5BE15cRcCPr58
GohE/7qDul9yjmiaZGpufSfx1VvRm5hoVjRUo7m8VWTSdwm/U7uakoOURFbxHUMS
VOINWOxSF3RG0lDfru01u+j/+PJEUBLdpIatwhOGUyfnHIsJXCx5yX7l3KyNWWzW
xj/3CjVpqY6Eq5mrqDh/iQq+FUQXlnGe/l6dwJRjc8OdYIneG1NpxKn46BYqAW56
XV+ZBK73MNitChj1v4vYcp1PYqU2IvVfVTQ+MqB/p7z5q0NaxH1RM3IwVvxYCWRG
8eb6U6nIPsLpuvUe47aWnHX1Fmv5mWF0LUxul6+u/MrI79tDvln+SU+jB9SxD1t8
McRpl/h66vflAottz2WzB7ebMb6IxjELbz/su4qrXurplv+5mu9n7OGBGntsEs//
ljVmp7AHLsdaoGehHnWpb0EFaAwhY4UxE/NXHtnj7uu5pBd+Zx3oMycB8ge+tKce
5z/9wAGFG2G+eibXidapxRHAYu3+3x+sykjq37HNj/116l1GCfOe+SzxIq97Gy64
oLkUnuao+2Kua65SUPoG9mWFLFwdF20nTFl3JlNQi91wfBKvdzVivb/oqy7tPlp2
vvO59Ew5G7fDUWfEaptiKh+KiUKAgiqxsY/8dSATE5n9aOBl6haLtM7k6cpw5NSu
2S7YQkFiVwE7A4X5OqvKphqu7caZyX3ScM6e/9/lQz3X5EDHPEboFxqRAkkkUG5w
ZUEvktSu3L6HQCdQdEQUz6+JR4MZCjFlXgyuQUii1Efl374vJWwuq1Dx8ljNCGRt
Kjm+mSzV4u9YL2RFrVJpjGkD1FRpfXR7/H3cZCySkY/ylOB0jooVMtCIniXfGfkW
xqLbR6u1Rx43rUxjCVbwDpNeYNMJWIxeF1VN4YPFICeaHmaV+SEOQO5Jsjxy8TNS
O8JVz7XrlScrewsClz6YbVgMYlYJNeEC6BM60Lc/n+z8es5rfO2Ro9oHRcTHljwR
Q8djvMIAbpvn6FdpbAWIrn4slmQTpE99W518zjeY75qDypLmLf/XOtwdCv/S5te+
KP1urma6t9NcJtYMjki8aLwTJX/10Pdx5EyHqdZT0PBUgmeP1Bl/3usdpGW+vQ48
eFOSpL+W6FV1ACfpz9dHXNaVElt4lRBb+e88XYUiC+KleAz4E1L+DGE2e2RfyPiQ
UwpF1bFjxJfHclrC0erBmxtsU3A9JIOsY1oc2h0nCLaQzOcrJdMZFqsLOo+KwI7j
jyLByxLrnboT5YXql8cuB2lpqBH6nTfdB0klbNc0/owjkW+2gGeUcoXV2VLJtbGi
Zi4zazOWvs4+iXZXDgBqV8DrllLTbe946MHmH/Qjv8xuw/ZLW7wp6E6+W/7kO0IW
/pMyxR15V7sQCA4IJfD+28YKaucARRn0s6mQYhKr0OUQjcKQeVL3ArkBdXag2toS
phsMPlvmPR+HEt27mjIWac5PLU9rhgmwsAcpOkfFGa/zxiKP0kYDV5ZXUPlbZ3Ni
A3YIHG27j/y1OXuakFM/K/L/pkrppaCzysKxUCFZ7/GTVB5IAfB2hCPGtzf0uXNC
j66s8VWaP8g1P8ikCiff8fLVpRM4WNqWHYbYluqp8rBLYwwvVzyan9u/cUbNcN2v
cQM6CemY5fwl7gY4KsXiDYarX93rMVCl3jHfY7+W03ajlHJiQR+52ujzVsKz0pgF
JYubvgtodSkc4TKbH7QciljlY/ynULVhKTF/B2EJn4JRUHI2H6EpJGOKYdG4meMT
MITLUmOY92+h31MoZ5XXCx7uEVvDJPJzj6Tab+cX5HNynWMW2MzoCEUP1WWwbRdr
o9n6mzpFU+2/9RGmyEMMvmxUGrgPxHcmrjKBW/IENb7n8FFQSww0lLdU6vdgY6Au
H424CS4fnUMjspqLFdiaveiY1qJtHtmWTVk6Aj44uXOatcyL3VHDXAMbt//vC0qg
L35vz3cjqdOblwpOHySGapdYaIgji2I2yXEdAcq3tlHUCjBo0HpfLeqFMqGrR3Xh
MqPN4Nmii1wkGm2PQnfIW8ortKRgPUoUkt1XmEIE/qwK4StdnT3LBcCOYoza30TC
kQkPwGa9MC6durjZQpHOpV/DW2RmuzW4AU+EmUSxI8fRdZ1fLDIwAvKUw3IqES4I
tzD3Gwiehg/SOIYQ62hc/AAge0LJTyRum3q4pYcm0gfPbNFl5b50cjRnOSUHD+ah
61CmJPrJvaUaPt5CgiQHxOOC2Z2wXMycblAD1zPL3/W4IxYB6LfODlRGn/NKcD3l
4m5FiwbdS+AgSRjpwKTVi24CmOmvqWpQnriE0mTiCTx80CgWbbulzztD8B4Iq5FF
93Nvd1jlpkCnWdY4c5473C7v9zmrpTyl97ZdzXos8DDM7ALwdENIS1erowtDdDHm
2umqpccm+t10x5AQ6kMzd9BxyVwXCeMWBgT8YQp8UObSInum28eqkYbXOq3fjoRG
303+O0u8QHv21EpFM114++SSjt///SVJSlLCGfgsUxl1uLNHNwSSTsmZyVTu0zCS
/DTRT+MvyDv1WmbGvD5Alh69GwLc8aO90yuBa+HCkb84RRywUvqWYopLwAgab+N3
0HWbijp8J5Y222NsY4+NPrSDGpcL+jpi9jOnQCb0sl9rA/jguAfsg33pKtDqSe6w
Em2MM7pEeCyKFjUzD1+DHM48QWWrfBPi2uq/oFmHoJx4+s02XX7+osc2Pewwi+Nw
T57WAFkbfdhEzn266rS1751re1bxK4YmoK7aomyYnvR5cHZ5ikkX56PWZiGLzAv4
Xx3fG8+KQ7u46/gbVm1gx0k6uNoa9MfOhvOaRbZCLybC7xD+rjLdF+lSF8gQWPGK
HpNARZBAnFg2farG6y43IZZb6U3Z9xcOppThwUhovKIzXxRYldVgx/LViMJUoQgP
mR3ykamrhEzckz/RwAlYTL3FSCex4BrAOtG1yZAYNO0/7BKwaXSa4WeIEeyuiby4
aMaE20/CcgwuliIkl1DENKCqOqIQsE/IIEMwzSJM91sb859TmyPzU2XlGIf+51mR
e4T0KeFtmTVxMzG8NO0A9Sfj+Lzb5vycbuiQ0W5RUaSX/en+/+joPNsZM/5JaBPb
34sItFzMej14yBT2PxClnoaw0i2g51J/oBxwwZTn9SaPLpDDys8wCLNG33K/YaCS
axyPL4EFFOzzzjnEwJUst6K1bDesuMYbqcuUUO528HhEhgUyl2ELvuoDoPYXlQRp
6tXbRTjMluJT2+4DS9YR7apnbwXRg594YWp7sV/CJGxWTnjzNZwyHdrCuDxTZFSA
2+ExjTlLjqv1Bc+fk9CfFpxzGcc7jZMY/VUckntPHeaed9oPsBnecm+rNqluVRz7
LXPsuXxWW+I9LQoHL0bOhgNW2QTwWeFqsOwWSf64iHDlwjcTGSvta9zrL+rx9X43
E0/hxHIHRWNSzX6n53F8424iCvSCwDdzN63JZhO4XPqkrSx+CaMTdYnNOX052IEH
L46tLCNwtnX60EaKiir5S1thBNHGKyFOc54PWOKh+RxEcMIM9WO5T4jtbInEoP4e
LkB7exlYysP9daADFdXpd/8R2+GuoOCrFpbsqupFqzvt1FbxLn8HgQ8veplqmhLa
sLSA1gfZzG0vmDEENenho/J1x8SbOwVCxJK5ng/JDVMDwjOJv0xwbAOwxoz2F2YN
yGrDZ5Y/86H8HnUZOpVcrcfWKC3Zxab8rJVSEJMa5CDwsncafl3XgIIJlVCejmTD
j8qaualPBeINkndJoyfSWyCNYm5QyfsVENUAbd34cPTMWJP+qNQcae7HE1+DflDo
lTEleWII1XPcyLvkrxQ+cfC667cwKpFT6u9KGqeDW7nX/1b3h9WL4kG3C18XqeRj
hR3vpltvjZmKum+IvUjLNlwgrRPfYj0ENe9/K5f7l6AB+CFLv9dN7rFbGatqeeub
qC/BygQyRqPxMQIqgVQD50fpM1XNTzzPDXkVS7aC4Q4uoLScENZZBHCBagO7fMcw
ztKXJCKSQTWgJYdxrhKqbmWhn1birGk3Xu3yWobg05a/r7MxVOx/YJbys7FXpN3s
036Gpbvhn3GW2VUVFVTWJDx8kYZo0ugJ4XiJ6L9uwexg2U/RC50WNVzTuYmWok6g
jHmXIJYXsqF1a17uW3Dazdc3xrIlhU52BBbuSIcYXrKb0jhDqODTUVnn9OrlXeMd
WdF7tIAEoVfdyiOX9yxRbxpO5bT3QHE6lKoNVC2HQXPZygDDlWlbq7eSZsOYkmLl
jPCD9bFXkhuTxGsTu8G6m8RVOdgdUqXjZjAxJeS+to6eEBdwFp8bQQQxX7PakHeT
LRtOFlA6wd2qQyfYPBzz8eDr8rGLEfRn1v9VNeAju+7hKDTh0+vAq4k18ooxGA/3
HXqV5uujhMWV1X24xst5K8+6mKoQBJ78nWxL9InbRmBshTYcouLUug6vvXWbJlbS
nPTS8cyx4xcET9SjzTPlnT+dXDHsK9qfwJBuNynWANDw157vXo5rxEOCou9ulA3P
k6O0QRJTQ5cWUwDsPLVFvvsBIOhUPb5+EUZKPbDWL3qr+NUTB6ojYhQP+b7dY4OZ
zmL/3g0b/gXmeMoRxUsEpMRWrW3LnKOA/0Oioktiu1yrm0dshPrEONAtQkh5jq5A
VmlLrGY9RFPUMd2jNq4rBfHATOPSSAIvsuTmnsghYb0iKJTDvKOsZ2vRnI2xk5xC
IuIjzKjv3ZUqn9P7VuaiXlbPR+5V7HiNMyCodOFDUEYIIT0+09WoQ/aqobNQNIRo
5RktDf+Z+oK9rtJzuRhpDXeOA9lgA32GmTvxFiGJ5xECS9H6eam3+TQAylTbK71b
Sd3cespE367WYYTwucD2Xiyh/MaJ6Fk0li6Dhfqp1fI8lVJEUZdyW4fdUu6a/7yD
DLDW+Z1ZfAD5O2xVcr/Z0YRajSFm0kwR5re6xYLldOwsam2rXA5fdb9WsrjCNHkB
AnzmffvMTLeLn3S13P80j2gSLDfXqg5d2Vhug+Zp1EWfifr8oBpZ+ZlSEQjYj+fc
UGVzWAMPGHfBfvB/o5kete5ViX0e024I6U1PySn9SDOzd2Dtjh0XeoAohKPs4SOz
KtjiQGIodOCcl7hO0QgNMrOLH63l5TkcKrGf1ChPVhG7kvRypzAuWeq6H4bIL6c7
M6zpDYCjnfYVxjNl8jiIOGTpsJBcuf+hNhSokzJOJfT3Nqg6eKlmJZDMUCY6SLjq
4rt6o7nsY98TqpANTMuen+Y3ksl+T7U+sbBhsGaBznPGXSyXeEllFq0cwZdATDuM
x4NYaJIYe21RrPgs0FO5/gXom6QPWaJ0mJnVt4amfxxsCMFesWYKdVglGGaMwr4D
iwst902dOBJd6tdb66WkwBPJ/MC8WlAK1DXm6e+u9jgB3y+3wyrCYYToRqaJrrE3
lfnz/rUHVrK2sAwpjBkuLcwsr/2qKYt9yG87zypoSKxbdHllVBzP46aT7WTo6JDJ
Zk1qHI4FGSfQ94JlnaA0JT8WfZ5YI6qOivc6QRlR+bisLmO8+H//NNeO9rpwgROC
Nlp3PCm3fUh1kD+88wc0VM9hmYKjIL4QvCdlZXX1LkBgo30PkqOihXd+qpWGoM0s
k+FAtEdpyUvG4fL99U20BcTTWzK81M8F+IzqwYzjytm0u5w/CQOQxYBw8hp2L2QT
jDRG50xyqmrrnbAfpJ7GY/+W6C+Q8P56B2f1erracNl3w/Xkq8Wg1ouOHXexEeH7
3+WWj7ygfhf/1Ct+RPbcRTIIRK4Ql40Sk7JQhgNUQU6JRkPyd/gzCC8eAJrNEF0g
tujGKNfIQLtVtP2c1Ku+EcwpKim+rbQWNat3F8jt6C+v8l+DOP1XOdZ1nIgqyk7T
mkLMVj0ru+O/qBIStiLpUyR/ttWqVmkEVdnCyCNGdT+MXkLotGv5tJMpvwZBWc8Y
YyTzlHSzbRRcVjq9YQR8OoEdjNiUpAFhQDs3brMMDpwOEWFDSEC3LPhqACJUC8gM
5EZhoFlCInHpX4q86MiQaPT2a1MFrDyQNA7Px8jbJozh/ledY7lajj/Wl6JUvClS
t23tXAqdYDxsTc1BBRNUih2lLMnlpcpV2xTXNutBTiseBz0TFXLgwvpFKKL2GEkU
nmtszJ5CuIlBDu86FfqZw8jNzkqDsS61eUOrYs8tifLqGrr2KWVbBhRbhDDj8uii
A9mOlHj075/T5kL7Mu/xIcjl8dLTz0OW4j2HUuTBUwr17TMPdbqFEtksAhYZ8oCq
+7muYl/CfwpAkXLpI1ydoRUQuWpvutHqBhS4ZeJbKcwSR9O7cnvnIq9xkVRnW1c2
14Ytltlkiul4joKIkdkz/vr9J8woK730ACPqvwFQXMkORcONqVDVZYI0Qz73oxrg
dIqeGpTJYLAAOlj3sHzBmhWhRQ//xz/4UlDQbC8GPiovFTxK5YWzp2w6v8NWc1yI
LkbsxQ0kOyiB+SUux8RlN13zAIbNC3AlCtKl7bD23O+jmosP7L0RDTeR8+sWiwVe
Xhu7iSgHqX8l0nKEtQZIbadVBu/u530IbQJ7sMUdywy7kDeCgTWh3PTT2cYieJne
4+tvCNrheCuTi3uxxeg/Ml/KlqteyfmM/OOJGI7Zsp+w4cn0mLXd7iikiFH3DsYZ
uMuqpMPHCO8FeGBvodqaDdlc+3yXvBUUcEko3Y5goMoVLpSzKIX6UHr26oXZDidT
XQ7lS4iMn5LkqG8rORxuGkxTEzXA0i7oF8yoAGPzrWxSrxUMeNlnSH24rfA+yCF4
H+aYFV8u1DkphE3dN8Ewmooo/1AFjUyYiDk1vX3X4mOhPiUbciCqPdura5zqB7Uc
B6mkmIR9WyiDj44KyAsHsjU+SChDEislXRC16OEkbrgNJYHVcG++Un+2WyAsjqVO
UTNNmibmkQsMYRc45ANYOxRpqKXDKBRH31LAXzKIvKh6mRWfS/BrHA9+NY/vYUmX
r8ljfdhtBDJqjtcV+JlnasSbrR728VyN8g/CHsNKWh8nzPQ0/LoLhruMdBuMmbec
fgrvfLTQie+1hjLxuYBBQKZFPADjcdGMhLFdc+6WqDpDUPUejAPBV/dKtdHmN82C
2EcVeveeKkih2keBc+VXG1cu9nG/X+2ftlTKCBgaIK6gKjtETHMEdGjYNqdpLqLJ
EXsmJpz/QN4JxTNV3lLydkq4wmrtzZV0/lj3gBYCJTCvdJOYcZO7ePLatUxzz1cp
r7G40qgDF4GXLkZEw+qVEwxcrsqEdJ2MhC5t1DaidbRgnUlQlcb9IwE6Wc1iezrJ
y0lRgV8jPtczlfaZ20ZuNJopqNv83sSlBZO4sySYEQL6Zp2eW1MZArgSCcVMKB3h
sVwHMotj03Owh4oAqbE4hUOspwdufKzyllI0Ra6vaZEUAT80N48xlACqsCiYTvJU
FWde7DMRH+2HJbyVCCZw/y/PBoJzJE0GfcIcUecNQtAt9wFqJyXHGqYt6VFW/y6a
j2Y65XD7NZcEj45QXwUTYXpegKji2pAyEchiliraamNZe2r13RH+qs8bO0PoIrxi
lBOcmWFNYVj/9wqOgz/0ZPySUgIvLcm/qWrAk51erth9oSO4Q+/ddVyJuQkUCdmP
LJvubCUna0N4cJjv87C6gMmro2E4M6XwVzgKRWdBaSmgKg2Vv+Lsr5OqaEqDfGNj
oTIcxnnfH7hIhcAKaJ4fIKZ4F8RlOoLtiRgHuF5Y7avwwvEyejTdKLT3xoMbf6JV
R0Ko2PEZosCyWkhYSCY02OI1O6eR4sBxFFKTsQFalESKdsZS2yLONz8iovX6q5Ht
3wxLMKmyeDqBUZc0WtcFFFW2BDdAEdkqypmt4QA6YEZkYifCLDpgrxanXsXeGAZq
4tcltTek1XNhXyfis1wkKZLe5Ss2mrmoYN25bk0j6GFTggxuOaSL/v31gl/7ChAc
vmk11PVxP9pX4r+0E7nRxgXzeRngf2EAiKztSdWSnjqM4QObRSyLr24iqzTdkueF
VmELZBwQllOJ625MWlPelZzRN4elXwgdek/rtj8wPaVbjer7KvHp4pTXtCHVRxF3
yu6EBubFijgJHR8wRn+EMmbtMqksGwOIHIHHT6YAJaWJCRK0e99a+FoZVnSETZYj
c6+Z78nc8JWlAEjJhi2uIN2lqy9L37a0d6QlJtiZht8deorOyVqIAF4UKf+2Y6sR
U9z2/dxrhGiO/LQ73/0DZxjgz5rdhHXRRiqkxPDShWAMT0pt7fA5l8r7z6Z6CKOe
tHZCuoZ2OgCtmRSdFGNshOJh1djdG3/PJ9Ej8nPRsLUZevvEetoL311sH9ioc4WF
FeWg4YhzWxZsuBKbHP/4TVbALO3uSMIrY4OuZOiqiAun2OYqtkqgGQs9bi9Kt4Jf
Cz4Alxt8YQ0a2dd457gDxDfwALC0XQ1cVeZlHFaovsOXuSemmflEhaphU/P+BXJl
1Ylr0N3CPPJG0RkvUKYuxj6JkWM14YjJYBvvTynlxZNqd2d/Dg2MgxfIpEjIBjPg
KCGvruJZFJSWAjveT8R7N+d1eCu0hzmCa3Ci7CXQbOeolsNFOD0RI9sXMW1PgTG0
/tJMmKaxsnQxQL5Km0vtD1hJpY6y17po6QPLHYR/jFehamtYN/Hh6JEH3r7GxkQf
EEP7AQkC1d0sugQDSgAae7wHoeZ6AG1hf5xwJPGcZz9+jwJLfKzgkzyB0qEMyBPo
Gw0wwVFEL6rYkjaHpmnivvgVVQKG5d5MiQFno5qgHSejEyBLfmH67X9jEplwFGjg
4Ce4k2sV+U/JoCEA5F+CUoUoIgGwO5EVaOSx9eOaz11dcCUm+8/9oUUF2PoTicnw
/TkQ5EkWZcc0Y3iXKuK1cxi6WpP7+aDGn0nQFZ7saKS0/M6fmMKh1Lhob30V5/xj
/vQ/o1wD5WCzPZOueusUo19EqQ5/1X6MVjo5ee5tvFyUx+mHHP37FIJmGejqqBiT
WHi1A9N+T2xWdFhjwU5cCEpp8XoJRo/YhA0o5yZGINDRQi/8h/gXP+pU/NIclngk
MIGke7Rw9KW9wzNoP4W2R6Xu/CsJ4ornqeroo2AX1TXKWjzj2bLluRNruQG6znF6
RTmoy/PygXFALgXZSZ9Mk3rwz+Yy4VV9BIxgnO3DBohibu41ZsNzNCEvyijXaJ6W
74wgc1wyW+eyJOcyuHUPhfz/Fy/kAAPSeFCPQwIVnB9wE8Yd0Y1Mbu+lmpC7qsAa
amcPjv6RFrle2TQYMp9yXjx+p22lWwGUH1omeybO51oWkjiufspaKB6X33vqmXXW
qbZCWBF88KLE8Sy8Sz8CwNIkNIwVUjF7Z1RApOZiakTW/QoKWYbLvRyBiFQVdTDt
S2Bn/wbdIMwGF/JgLas5yJp14qirJdT868zdSSQ0oQcsHwfXEoOH0xj2YAiRACCN
LgV9KK+mOB5If6IOcvfX8+9i9uiIXaKd3VqQJ57VCTV6z7Kn6FETrIvFcfcVSW1e
usQLWauVYzuMhjQ+hsYJCkWTfDykPSvMrJn8VqcIey1G59f4eldY/A5+sulUTet/
c82BRlw5e3xD1L4SsPIlh1W1j09X+WqoKTSfad3sYl58XRBdwrQXHx4Jo17EEYPw
3j1M4NiYQ35SohjQ35srGcEDortIhlU2Yt4iNQcZ43pGZSBwARizXPFlOdVLrqby
pgjHBRMhoFSETdOapO+DZg+KpokqnRFzLGvUNEgbGaA6coMvAOweM6cEDAI/NNTt
V9pd6RN5cWRWf4mjeqsqmwdyHPBk6m/w5472TAeA1GsHVLmDgPXfmgsGjGb7sEDO
oADb8syDAd24Bh1+wh7+us9SV1c2OuDBigsXHsbPQsaFKt7DOI8G8OE7GqG//R86
U56/YXYkTUWJqt7RrxHJezZKZF+2QaEfcPf0qFEN1iKFLmEqBbo7Fn/w7VqCrjwE
tms1d3PnDJVjURR1Fi69TQZDSfDpc7zaPswB2ak4vS7kRyxlAjqnLQQlmb4K8IXm
ea8htD+hWg4zrnzvKTGjNQV/eEbiCyucYnYdJRESSW+aEEfi4QgC2TTHe2V4nPJr
nbqXjq9hBTLgQBOgCB6WWCjprTaBRPAEMM/xRTLVljgREVdDLK+NZKoJrECyZH0A
l40M8C8wkgBu57IkAdco3o+jy29OsZS29eTgLkzaM5A/pXzH144Zm8L0dzCmWa6L
vwYaM3AuFc6l6jghNDQhUDzGmVwgCrtgoTRCG6hadqDY7IRKV1PEcXYskj+WhBSF
Tv0mYsetvbdPjBya+nyZjFxoTYetBiK13iiER1E+9VcHBiGGmchmT9x77zN0qKOb
OFn1qVpXclXov4+rT+J+JJ2THYbiOFgy5pxBhpO9Px3F2qHRmpOrFaSBtzkmKi7u
hJpMsO6Seg4fj+TfaXIPz2cR0FlXzEv7wzVBBxNjgvhrC3kTLL1DKgqeDOA2u25T
eeZu7+9tYdBPe7+mrT+QotDFru8c/jJ82XZdl9x8Xlb3C1eOmHXS/IBKiPHaluP/
tDhzBkaRWGQo03mBZXVHxbM1zgqZJGs93EWzp2D1SZw2k+RRyvLgT+w23dFyzyWa
+92Zg7Zg6zJ5F0kNEXPul5pX+M8YTOysPPQN6Rzyivv68DrHatdM3Ii9EYTk9fvG
S3jApQFArgOogP9qC7frskaNv0brhylC9jzNkmW/5GtxqO7gwtSVWcW+T64q/CH+
ZOKxWh66GLIWhv3mud309UBeCh6Wa8hugx6IVlB4Ytxbg6d1V10kV9QsHgOd+xQi
V0wSsfuff8nr2QvUU9ZEfhDqvrXzC4i8mg5gq9fdgLe7EqTiLfxCN4cvC5fMe0a1
zdKZhrdCHFqHsHuESIWOYDvf5v42uyruG3dVqdlAhgTeSk2Ij4sZ+mPGS5IInpAt
e8Ec8JkNrrsi4WVk/IJGHxlidLW8coEgOz8wJCUWyPiECfH1kNuo9MfVIvCOCKQr
qiUDKnWqHpdu8S7mfEKSA1WriMj8FFQ0SiNVEIOUjW/Q52C8bNRoz6UJtVLqc2IH
6mZ+qpcMcr/DVZABV6BmyfyZTx6b2Nij930vWuIAExm+PGVQIuZZZLKKVH5YowO3
HGw6VxMR7n3pyZwZchb01DCyvzIbFe9Q1SgFAQSs9NZMPO0qDOJbJLxPyuMh/agG
eDiW8fnFobejnU9UdeNaCmy+ZWATbGjAQwD8jSkvIJl5pP2hvkp3f6Gmu/xgISm/
ca95CfljT3oDIIFYaoJqlOhxJwdMI4pCKQ4mTM+s09G/B/olumAIF+42cWy6yEDG
t/7QzBpSbBcxzZhxjgXcX78nfYs7fD6QHjg+UHMI+QyNNLvE+Xsv32/Bvv0bY0xR
r8GC3+uq7m3SNvM3KPHieXPZBzc0eDqXYSpzBD+4Worx/0Lc6mZ30hnw0Rg8NQmT
NpLpIIiK/cl7Q7RUMa+AJii/C0fCxPriHfTWW4z2G84PMczhpUUfqUrEB/lsflsm
3c/6RL0cqNjKDs/YRxE8CLjkDYI5uKkV42sB1UIvF9wGwSTqsfeyU6jpcpxuBmon
fydUmtRguN7VGJFtOJrv+cwRnEIMF7B8UbaIEIrBlYWTEaTnT8UNi9Sq/JIbyuko
WSMKNumsL8wa4ihtPe1dBOvo41wE7dbxe2pnK2ocunnV6T5Q5gNDkA47b4kWtZRD
tVOrVt0ypm66iqT5lEVOZVHPvTR6VDhs/CrE0+TrKxRYVx9ATdSYUsygR5qXO4WE
sXOYTTa+N8Gh1orH8O6dohoU/0HKcITcII0mZ3kDi4qUuKY1bFGD+Fw3IdKUPfB6
63f6YLWlicpLkoNN10nGJDwQXIdjT1SRE5e9u1P8C7eLunB2ykDjuG+C2jXDv0dd
iW8ScVTnFUOsDllMaz3r2LF1nWIx8zl0v9kFvg8CUqfkbFyoqcrMZhKsYte64Bdx
4BRGvij8EOwC9Ma8gRAqLjETpLBDJ3cGY6nrSzTffC1kyu9z87jBTKHCU+7rzXEa
fDTs2yjEaFbHNdYfQAzZ29pOyyDumN6L6cRaz56qh8gGkqAI9j15TKnVo2o2lsaU
ts4TKjWnt4kpl4juCEKZrAfJ1P4h+3GvzsHQzJ/YFqKFx91oWtGSRhwE28u19YqS
IRTZj38ge+a6doTZ8ZmOYWnNuGKw9VIRTjVPatosFYeZjsj/wchVZ5eHVttkflHy
GA8uA4ZW9OS8bfd1YC1fVf6pA/rxPwprjy8TsMELzrFb3SUYR04KsHysSJVJtkiB
o+FqtPHtNTMTirlltNVphEeXfIZxNmSMGEocRoKDfXb3RD1o+VACiYHey0reZU2A
9CMwU2PvAXD/UiT3Ipfg0mUfQSiMqwMzgg6eQGj/pqIs+SdDQ52jmRDRxMp69ttY
4IWyQeBRtqZ46IXQmcyQHUbuyJjWTCVfO5hQzGTW6NmZaadMI/v/uyRKaItxhdQq
ylXXLBLBx7jR0jqNBPtlvPozFoFjKf1WvL1qNbfSEA+CqzhAHIWbDWdG7hjeYWwH
q0LT20EJMRpgrRDbDV90+I/w8Jd8pm9HLXyC6yMjczTj9ORst3ufXAI6gnIXaFCb
cisb6t92QhJyZ1/9mdJw9/xKZG2wNXKbd3JUpnsHvZ8wkVQTeWNYGh3LJKNbkMJX
ksVEvis2f8e7hoT2semWzOTAMfbZzhLnEgMd+b3ZuKmCb3QmSZ+tUZc30obS+ELN
YG6SwPS1ql1WiDr/mxcOpUe6qtqO5NJhmHauMByUH9H0UbrVDXjPK1oT7gW1dRYH
jHqiaxmNv2xaBfquFTku9NtfYEMKSeLqFUtwdD/JUw6r+o/nF6J8K8Rw7/JMJnlv
IqqMgTRJgnEi7dXIg2KMyTYPwDzy0DKXu1h3eYcogsJy3W1SA7Pb+DvzkILm6sRd
CBqF12q/yMF49CvTM9XmYRH4tqopGaVBvV15hXBCfEaM4xlQ8wXxr2LWieGIrhWy
HMkk1AE1vUt1+IFNdw3blXSmzK8PAgHW2tD68WgiD2p9QHr2F00K4yKxUFVrfni+
N+WnvrNlidzzAaSsdC0NuFKjxK8YvZWWWlzucQW8hGloMcXwm7p0kUr5SS/PlUHS
WSKxaxxzbzW2v5L/DnAjn6xNyM9XaPiSeK+O94MgunGiWTWv68E3kKKxg6x/bfEd
MVQK10ZCKQnhHQuDhJROoTUOQN+aFFVauomBWoQnzKGOVjJKIJIPQ2cHF6jEaB12
OO6J3UF52fMrpUJbMnRpeKIkzphtYdZYSI+We697hymFAmVbfbwAN8dErHlpvHeW
2y2QinI+tl/GDKSegTw0orduUxhhYL/8zlymslR+b7c7eKkR7ueWwePtQG/dcCM3
SpNLO4/A20cmkZg3RtOq7L/OxS+0TrjybBD1/SsrzFeUBhofKPrkHeZ4AF4qhlln
LnqiGYgAfVUqjV62Tl1HVESVU3MuMvadOEmRpQPhGZyNZnG24GoMkb2ItFQvDAun
X5kSIA2kI393LuvP8eKw5UsNl7kV2V5KfNv/uMoGaHDeZtP2m16BJws3a57rfXqp
WPAOJm0yybMbKrtUfxWmiZ7oPLrizcS5EQMstAnkc8RGmMhXFth1hvrhdjQyTFSQ
0bn6EHtgQgntScH7JAAxXG6egq6zx5qTBlyxF4qswPyQ6hwHfHeTNIxphYo/Z7f9
s4RBr8hSuBKdH2hldEQ8ZYbW+8mK38F5aSLFYaXGyWVvpscQ3o+96/qQAf3oQP1y
INHsmG4fyi2GKKRfipYmmRxzZ0HMnjWS3lKBqdpd+qfso9BvyRfc2MWV+mcHq8Hv
i+s6GUV6muelAiBEMeef+SRHmrqm2amdUzFwQqYMgm4fDj47LSEgkPglntSUpvds
Lxf+LgwmzyiCd0kIWk5I/LyafxSAhcAvvVlF9DPJLD+P/AJsgv+MgdztfvxOe/zt
yIYHEQ4NI1ddfWwoe8ah23epF//hEZdm4OBJjEtLy6C+mlvMioIMBhEupUnINwJ4
PFcU0f3pAuo8YloPW5oGiywLXhfX5lhfPWK3HxyZuwlHG/vf8UdiaJ4xhe8d5c1g
ictDn89fqS/7aKDJELlCcokjj0emttZ7pxvGKVuOgz3rN1qa7nSY/Ym+xUQnjFJL
MQjBti2cvWQ8dpxGWGHCvDYADgs78zc8+0uHZT6rZNgvlQ8LfiONK7vK86g2RJ3D
VxddEf0/7RkgjwlFxu6r0AR90oDUqPagvhu2XG5eEQAScUkqGECsHkmLKodFO/ih
nhHRb1pSFH9QmwT8lyOVZzxv47wd/fWKTGf+Wk8+tGeEa1uS60fuTQa/eXp7wxYM
S3qgIMj/ZgVkMsuD/uE2cXMAh4mA/zKI+xxyLmeUkdtT+E0/XH6U4wCO5TN3XqZJ
8Aab8CnY2r1td+MwTJOfcBE3Yjs8gGhcDkFX7gHvM7X5MvFXuauhqgVzCbKYBGgn
JLkxHwLT2vvGPdnWUiBB4/u098XEMnqUsUEBr1WttjzTYATraru23zkDfVZ4n1EL
+U/FjBGy+bj8HhN0XzkNAxz1Coo2qR4KHKUhTHFzsapPZC7ynJlpxlTArIfnDbuA
188zlXn+fq9wvR5A0VC/nGvjJRdWCUkj1lL2V9vZCniVSk55cDv5OBK8fUabYMIY
Wv1Lg6SdFV/ipHTRp8lOWYTl92v3YbgFN+FNz2JP4R95Yt73DiFNUMcBv9P6uzBS
zwJOkt8Tg3a4r+Id0wx/Md45ju0LvhIrk4HqRWSqRrGzFnfJ+pVGkXVNzqyxZOny
/DAdnblcK+1T5r1ZgpT4uQ/IOb9PiSaahUerTLGFbRQPKd1zCZXeS8VPdRVz3GTk
EklirOZwta1Hfq7IgbCNs45/wWdNA8nHnOd9GAN+byPjFXveaFVbRZX//WKi307e
873Cw6uu1q8Iil8o1cOojcFTzfn9UYdXQVDSm2eP/7M8WKFgXTrvbIhfJb44HZau
ElgEIq+rFPAyKwJHqUuVOzqHifT1fKj+GoyYucQfO5lsS9CscyJdB0/bu2AXQ2TO
ZgA2ftCE8Rmn1XmYcuHklLHRoRVE1T95M0lnsaJxIcxHgVn+Taz2kV8bNd4nm/Je
TdexeTS/O7OyPRWtWuC5TWVzB18DZNnI6Q+/e8L3gO6KvEdZB9+bdHHE29k+afBz
Qgce1GJ+Wfe78/1GMd7oSHLL3KEWvhcF7gc6ex1mT5fhC/volHAUiqGTcjCwOhsz
trJdUXE4ZJHjXiVGdzR/K3mFUHMbQ05wmvvlGk3WhS3FsYwItNvhZAf53EViZWB0
K3f9Z/zvjjut/oq1IMr1+PDPYOPMd1iWzwBM2IcarRE21f34mTHQ4CFnUJ5sSWS8
wr+UxvCV6moKdHD8+GiUQ0GFz7cLFOkFaIumFLmTh5fi6JdgBSOIWq078lzOwdVW
+VfcC4BZtNysrc1bFLsuioct9nTvJHTSjx1cMnNFk8gaS3fI+JIJcLSZ2AXOwrL0
m/QDbS1NEOgP870L/TTtgymjLd7mmS55JGz37FQIoNbUkUJGwvrCdssEv/n7t/gC
zxLdKGXtwVD1VKmBjYgOhj72dXsFD/kUNcrH4YNc5Bxs0He/4HX8SmuERhOyxDmI
7EweRbBFx92lF8nPhuqL7UC4XomItoF4O/N6OMPPBY4aJI90aj9kZNdTBg/3ZZsp
MHg4uxF29YimR+OH2zmw9wiS49j5bfZbsWMFc6zfdgpa5eRNkbnId+BNXJeBbm5E
vOntyUqHqWufdrH1BVJN9uqACh5QaWGSYi0aVUyrNuOapG5OI+aJR6GWbr/TQxBz
WMZehFxvnYOdgwxCsxX7BTgUUMJwZnKV6CiTHrSdzOZvCFhgGcuXB852y9PBIfZL
eqZlyQP34nqjAz5zWKourefAWu+L803O6z2rJ7nsB4xQn5QuFg7qbCEIl2TsS73q
USQk2jN0XWVbsNJGjnrfN5uwgHb55t+xYGdoWUVr62CqT8+I2xZUSGnKqnvDg+Qb
NejfnOuGa4fYswzlGSp5171KY2pO7us2g4M5FK63FGyJRcIUF6R0+PWRKa0qaUxX
p46yW0ULCkgGM1PWigjRhczP5PHeHKYM6+dsfLmWbnK032gdUzTquPD1mObYmznk
ErO3eGd6WQKhhfFPCkg6DKqJJswKM1tgX/BeFiCPZ8RArXr9+zozrmJi7IJzZJVC
2vfdr7Rup4WioAGFzbQMx64UcDIG+TEsCqNdnR+JiudbQgzUFud3AK4I2n85RAgv
F5+fR3JoEGp8AeK+QU3bxCeFwzFnEhFTCpFr4a6bynZcUWJVK6ferSqaQ/Mt0I7v
nVCFutMtyEeY76C2DFG4Yt7aVaHolA2KzlmXUGSy3KNMk5WWmLv+dAAdFYoqfu9J
wU2pQhWQlv2unoL92lpZUbOjf/9ganmkVdR878IN1U93Aiy/S8t1MRiiNvW8Q7gw
b3wNxdWxVVdDhe5xm8F2ZAQpOQAjgyCR9UMirWiNZ9E5Veocyy8Unn7rKSgbn3FV
zP7ihzhONmd+vh7zCLGtv8XIoa+52+XjZ6pB95f4fUnMFd9qdWTh0vusGYMhCtIk
asHW0Di2r8ypXVUKj7yWX9F5KK2Khzuh/ab9PZOD0mhOsb5V1JmuUyjKKCvHqDH9
jeG3dOcpn3D39Ya9nVYh17Xsfy8MOpfv6+P6gSIdExo7EWxVI7nvLaySLqAYJXAt
ACrlALqADkcNl+ZfU5WST3EQyk5rwg9HnBatA0YcAvXnRnYsUaqVu4k+iXuO/+fF
DY4vzdMdnG4p8xkMJBWSIXoB0/PQ8fYvzrKP5edDY32+x+7jjp3hDDwj2RYuJPVw
ICf6QpaI/QAbOTJYsFdf7nnDrBppcGT7VrAKZcMw/9x4cmHfcKnfRZBV6wV1Q0O4
1KS6R4JKwGi3IOCtX7O+g/PHXb+lTAFp2FkA+Ni2fYOkBv5S6AEcWWlbJfgB9Gt6
eSo/sccitV9dRn00LBwGIhFRSq6q93KvMkZnWcKnS40mLem2kVM8FzqxrcOiShbp
G/ehfM1KBqUXj3NsYKGNJghvN/u/cbAhGCdLOK+JWnogKxbDjDh+LrPSLv7Xj7EG
0ismNpY2Uxpg0l7dkQv6nz/tkVx5hMY0Bi58llOhTosJdNz7/aVbwS2dfg+C5egU
Qvp1D+c6i+DtBiD6CVcikcAfB8rEa1cyJta2y7cii7JQvHPejyR/J29NOfCusHoa
V9SDYIFbrln3eBJgaqcpi8WXmA0HWu//2WXa5q5RjzGzYOcmUEHZZhq+FjbM/ey7
eCIsbD3gP3YCMGtRIWIX/xxU7JyVanpm6ZDBmu7z+rzh8Rq+vOOeb224LhDTzvRS
K+i8meZQWO4Q/8d+0V0s4B4LYDex9kS4X+ux+TU0IiaVVnNlA7KgybjDhUNpXrZv
1capWFF+u/d5wFQCjmpMcgPqPfzyv3BVgMxvJeWPmXxhQbm/b44YLK5NO0lkV/ih
8vnVhoHl1KIC2kwR9B5U7cPWt8X45zufLKFEv2WOoFrg88I2ASWv0+QIg6SYsA/5
v79pVqJL0lfxG3zyteIXhFH5ZvxLNAA6C6WemJELb9k03IhhIULwwzoDNv+1WIiE
Eg0mytXld/OMnIl0VctqkG2XkAPStBMi2Evx+owZ79G+1wqqmV7mEqZfrV3OLJXw
ZFUhn8/Qw4BcpsXwbtjDk6KeS+DdoC7Pqk0xW4PWDM9r1w3CbP5TXOnAA/+ZeQh9
61nLuzaNXSfqBeP3vu3h6kEteWmvdQe4XRoT6Gs9gQsoZe1GlN0IcUHGMzW8V1+P
Q1zGKiIJm0L0Ypp8NHSjM2xVQBm9BTyXFeiCvKbDsIKvc/B5HDvAlg4ucTTggOMb
RAdRBgD74ERS3CgjvjXHQ+1Ou8lwF8Ki2ArEdq26/PfAh3WyHJKVdcT/gws6ja0x
+nR2/4n+tLB5wJnwLcZWh6khWvrlkmTxRg0GBkS+fMsE1i7SyIoNzZRIB3mBgbS9
/J/tKRCTmvIUSyYBZIz1JY+DHm9R+FlQTu0r0+YHpuaBtQjvdnEUQD9Z1OGl5RZN
x34GmH2AQSLUR12aPv+C7IudjT/FC2/iLApdw3r0lZvEp30D5a2o7M/7JPlAsuFi
fecMvEdc/JxlgJ/VmKw9bcZzdvLxx8wjMXr8xDkRRZrUZc54WWLkfdXsIZDi2/zt
yhkAohBPIe8UsfeQSErbR3TGKlNR36c9GiZni7dicoiUZ05F0jrnyFIDQZOKUSfC
KAEQaycZzx302qf1la52wQ1SAzu3t5aDru3RJ4DRCfCi8HDk1kwkCc90wvifpr2I
+NaiAFLDQaV1tdapc6tvxS/iybeV7jGfIpUuAJ9i5GCMfR0y5TsyExjmfyhIn78v
tWOKJ8yJWI5E9Te10FNOufsA5vJJjee/3eimLmUY9RLV++ql8IWv10OoioHP8E4B
LiGSkj/zyumIv993KVh7+nz+1oYeTcyK6IML7OCBRLGuJouLuWoGcoGyfxJVdBeL
QZ9TtcWJlqsFX7EcjO0vXRQqzWzYchvcS/7ZiGZQLPnhCXpbSvqR619myC0dnjzA
X15m5dHSge/c3laeb8RyJ6gtnJ9oNxRmJMqQ3rydg9nhbMA9GIQYpzTr1HPKCe9j
+eQ3kegj3GwujUjrxJE22lkQO4UqD3f6NCOdStc/jAeiUs1t6DolZM809AhAxRAA
dVKadh8XXAnKkN23I/iHvmrxjtzdUpY0ejZEp/Azpr5w/PnT1dFlC8Lv7KJsEOBl
/21OeGS72AxnmydBuKphsD0FXBzRd2ptL2A6aSn1Mtw8NDbo/Gw351SBYrHWWhdj
uyGZ6CZIG8djV4jLIgr/XQhbhCwwY0/4HW1HX/93mbEz0lVGd4ATK5QWoWf500NO
ZpQQNG6JYFBNa8vcgIR/Lh02jwbYq9pvXJqdRRt2y9+AtwlgLKrACt1mCSKifIaz
leLPvHSEBiBumO2z44rqkmm7NhMzG1KqEbYjUNcz5ZsrDX9KInIW1csx5egc9sUi
LAhSy9nH7vNEynRf3Nd3XnnsrxnGwWRe3rRPAw+Hj/HvBD1unjzMCtov3kVe5VEJ
sPoGDi6KBtbV/0WMITS5bpW+lavcOTBgNiyzSUYwa+54UEVc/BRM/7+hSz53pKuw
s4zXOAH9vkm3HvEgOSVaF9UOFwahwAMEANnhIam03x5HwmGDu2Yi00El8Ns1Qbr+
TO+kfCYTWziPB2sAP600Q8LkBM9fOSa59nbDsHP6N7U/2tgzeW3WJupmiY3fLhAy
NrBakfTlaC5HonEYTHxq7RbvUm+yW+4KaQUOoGmfDC1Ck0uEacBwO8tr8+bfGDY/
s8DMijaPeHXb0QDnnah/2heJmah36Zdqa/O1R0Amu6EdyFDu875hP5txOhyzwovT
W7sQ5XWPdaaDO72xGCjlfycW79ag/ex6uFCLuYaS/DbjD4JIK6qs3ncoS8lqg0Gn
6Eavpi4mW40mduugP2frFtUYY+C0y+qtrr2yE1O1O/Avo5OA8xJucuik1Qo8Ix5O
sp2k8X2Z2Trsc74GZ8Tb4MdtfJ4Wcr64wOWZCTeZxNNm3SyFLrBoSNPJJQ314Cnz
DrdjTgA/f0XXoUXqMkclsfGqb5TfLMfLzWyza+wQPJ/f3uiwvN9ebni8+1JBNFF4
ndYjMVNDrD0OM+huhV+nY5w4JF7MBPVxCMbL+nffDYLg+qwRpZ2W56oU2rrNawI0
rwroq+J9OHNZbQI/WRrPiOb5nvdH6AzyR/rca9yRrjhkbt0llAKAvp9rx00odXcd
uTVSDqs3axyLxkJ5en1fVC4gdHEtjll2/Qaym6nFOTg6AAbsWl2S9xT36evFGJWj
L+/NHJNNNSCn7gSvO/GXDAgpeSX9YvryT8sBExJjT/CV0/0mxRnZuxlukGk5Vld/
Muto3UgI5hqAl4Oa5CinfN+Yie1TM1uJMmxePJHtAMAkM/bmIbYa1TZA41R9QGxc
BrVb6hpTGAg/Ju3Q/0TEHI7sCiCKqCZHss7Tkqs+n/tOpkPvh70Vv03Y32v+F3qV
NvFvOmVT2CmOqDkzvU1R6knqwZ/jIh0vYg0jSsKE0piFyrBfBxaYsXGA5ZaBIVM2
wJwBKakKpQL+CxObPaCZPGtTkg5KZVkLAATtGOVFDQ5eSntGms8Mh2IjB+qe790r
KPGq08kfC/USMR/HArO6QwCrf5k7BY1VwBm5vIwE5aJr4OKboNF6N0+YakinWCj4
Meps/9tVB6BZb9tUMZxfJhNFUZrD3WfCUbQtSoJVc1OLR/9H0gk2UJlr8w+wJiX4
eCmCzXcbE4ufZVv+4beqIJa44jl7R7HHwQmoOvaw/8D+uCZqC4TlkJmlIJrjgqm+
xhlid4u6RnF/31LjkHAKU1kgy/SDybuN4dA7yrJD4IVl/N8x/QnSB0atL8IAAR8w
78AohYl/Abys46ktkAXZq6Y7qiP+7qatHLGi979xbitDczZ74ai9IdH7jdcYvgC/
nK4bZ+TEgzmdQrZgXdeY+eDec6TelOdRDIfsUbwWadfYE4RwJsHRIM1jztgRhMaN
DH0gFBPOpFVZwEYtoQwzfzvZhOpf0M+0RqsBm4vsssC9qqIDYw3vfbPTwPc6aDzP
hBv2LslpO8IWBliggFGg1pT4oq8KauMAWoIY6p+GXg40U9DTLQi9eDPeyWfTPuBH
+nRHCOtSCYRMHyzoXUZvl6ELgX6kKq9Awu4nxSPPhnBg48Bk0VGbezXzXfUF9K6N
eHqQfrTNcoXOuxE3YZ8x0R4mWQ63xc7KxvOAumSFEFmyTi4lRCZMVTzmgql6qvOl
6oBjNF0fiQd84iZ7P3ZRjHixLtYC8MeH8EtAeEw10IYxBNl5xM5bnKC7L7CAJzKr
/j1BeGtlWho6IhV+/l4cdybiWoV1J03sSbHcNKhLPpA56oAwJ/ajYQ9CUlJg4ZgI
e5pQJHzr4vdE6NTCZIuEo7n6PDGR8ikTQEjkRtU92iR8Hvden6EbpOn4Q3f/oG2s
vid5DM+vy+seZ8C8VEgY9hFhxxghjgdJNS2QaWvqbN7oOQXPzlaAeGjhEDxMXb/e
QvkhlhSNxb8ozih0qzdpgZrseK1sbeIwqmAGX/EUiHeHsIgG3PLV4jqWp1wT/ILz
NLf9re4fRSTjH5/ay+NdtKmQHxmhEo4BWSlPzv80t5Fdnh/nq2yrnaxS4CUOGLqH
+pjZ/CBUs7sT1jdDj/A//wgLTfM+kFNrFcJqZcTdl2CE4xgptxdgiWpGWXvClCXl
4jxlHpthTX9RAdaHkn6Bk8RbWybog7vixBn5sFwJgsDpued1iFDAyx4QXTDFxyIQ
cS7qRkKIwapZBvIlWUJ2BXEVfSoAE6sLqgUjz4Wj8RWBn2pojw9eozyXWmzQeyim
A099cTFfAAV1zNBdI1J15Qx1Jv4XU71aExAjsZXuzAR4OM6EOYnlDFCOg2miN+ie
OmZCY7gQMOIDJZLoD8DkWj/3RgictKRg/n4LHWataW4nVwVZNdUFi1XdcSfpaexj
b+6eTA089uOuVzD5z73sJ/XaeqPxKG7COeX9ar8fsAtQykpkIdz0ukJrQPoMkLKd
YKqnpbjKs/a8jdYvv8RodS8d86DUSoS/ywTa/0ZTgeBbYKapMb1CDaTiq4/oltis
UWpImCDx8ib8kovN9cp7FeJByDFvuJ9GEL6xL4y/JmNLcVxyMopO6ODWVRZp6gS+
t4LQo6n2y1oH5WKn+DemvXhTSaicoRCO/ciBFOtn1BWEEjx5ydqTRDjdCX0Pf9G1
LoXGEBrFUz1xn3WuBFuezaIbs2JF+AIiHsNHoIvU3Iw/2J7yxoMe4rGieACefS7j
PbipvAdoPXb+F6PR8T3BC8bZO3gzSYeJcJsO9dc4Ioh4opuiq1ew11fSQXuJAAmZ
/BsP+HtvFKlyB1kYJzH0kDDu97xsY4ZxQ76hWEQfZiEKlOdSsXu5tg1OYxQW1/W9
NMx8KLemEj0tY5IPSeXIsR0NNaRHcdhSVYsZFMjG+orWa42pTC7ZX6tR1uw493kO
dm5b0bnKx+4LFhh9GAHRhy59dFwFr8mtSWfKxXzPx04HHFN6/nEeH72+Wjt9/IgE
X16AsQT8axl2dOEv/JnD/9gOxSth4xZLgBCOpklZ/yLXXZgTa9Itv/Ze9LId8N4K
5m002/9DN3oE1oaFNLNPgWXj4J2ATjfPbXYfwkxODc9Zpo4TQE559yegn7mA/bB1
YjBrEfTXe9avLuWMYmGZJlqSp7qHMwwmdXgXLRLHGYeZRUwFZQhyDkxCaKH1rTvb
8lckLPi8LGgc6KDdUNggkuMkPDVPUAaQgzPkbXEfPAefzahVn2sVKr0575GDuEll
asY1BkJPD722sLqR/fQ23fbSuok2umFs8oIbtzJY4+7E9c2jufp/fMwHrFsnE6Bs
N6g5rK59N9RTqa4m1nu+xVg5V8ohvMuQ4MNUiNgqE9yg4HTK9FJe/WDXMiyfD2Ai
ApV8YEcHHq5oooGvlmHkpR8Gue6BRuewL6r3IOzNiwmAHYx64dUkVT3K1YKvZdE2
1IJ3dIffAlI/MU6RYZgIAK4b3Mm/zbAeNuCPAZQtSPVxwfON0qX7UbsjHa3g3qBx
XQ7ovKsehITl1M2wGVZaqv2OijSVthAjbkVZmhIR2dv/zdylWHRQZDzNRx4rUQyC
2bpsmgbhBYMcI19npqdUPsQ5ibDSmM8SQuuGylwpvvs0zoGQL3ohaVpTPCCVdVII
XBN3mJDpXvfhjaIO6tZ4O+V7x9UcpuFZloqfLHlMFq7EhirPOZCP5gYvxU2pj3Cq
Rz+2CiItGUbEIF8Nms/xXwCQZmgvAQ1FlhPZNH3QYZMjeCoAWfiChphdSwBPGic5
P3vc+7rE7kRw1rToQYZYNIing74vTJp/rpd8pMrBxtT0FLS1Nr/CAqAGFFYUUNAb
9GlzFf6A4XYrCrso8QZ9Gzb/hG7/VSHLbTqsL2vL6bk/FEEfxKf2deBqp9DFdIdZ
FbuKWskZypwEJM0PJZRbBRytqb6emfHT5LhEsVk1JtyG38fchgpBw3w/LZGCqnJc
Q0+PRrVTfdPcxOUXUSSS6kBXl/BXwNb7c+NnAGiThkECLh2CvoyyQwdPrr4fkB20
7O3ZWXPAXyQQrZ0fZXYtfMNfB3AkD+EkAGJ8Rn8DUIXhSiohq00i3LkB2IpSDtOj
vFx1Z4nrQd5yWbPHTsI2Je1OREAKxrMoSMtOOizRpHo1Ajc3pfIAto21utt4Qto3
m0aOGBjIan7Zqzu6hoDU6ZQoE3mR2mj/PSFIcrTeh9OWYiuZ+FHGmhrC3UKF/+Bd
P3u0iGorg+KOrBm1NwhFkLMLBV+DKaCCCh0YY5hti4cx/Y5d1CU38Q7gP41ZN+GP
lZ2MnaBo8ppUh6NwF0DRt0LIF2aTQP0aN40Plh6+XBrEDnZxRj3DsyfMhEWAuteM
IMJ6rP0Ci6rsgqVY1nrehWy2VCKkR+dPg4Y5048I9Gj5in3jT/UfghXnHJO90mW3
S439ZLgi0QPmHIjWV7osP00+HtUcZU5tsVxAfMsCA114w2F7sjEK2ljfEwgUPeM2
zkt6iiQ5KW62mQTaDrvNZ95MToShjbBlX2WdMsgHKcznjhazxcDDRyiDQswzSyi/
Y9tOgNcEIUoKMjhr6Bqdf8xw0BFoXXdxlR5WW8uMbLfELi0eo+/THIWYNmOHIcf2
hC1imN19WmtbIQDm5rNW3m4sVprxbmxgOdMl5I5jrxjZZzob+SFyJasaTM3hobj0
LlDxNtmzQTNW/D0brzFGK2lL5AxQUalae9DwwE7cuPsE4MilGlcWolW3r3zP/ZFK
raYKm+Wge8rdzCE9S05RPGPmO/Ma/t/hPDkBelf02Om/Nf/7NOksBBBtr/Ckv7+/
LyphfoSCqq2kix/CPmh8NgTGYvq+Cin/CfOHvu32O9yx225zLAP9+s09JmQTN2r0
bB47bxHwqxst4bZ3HbLiaJgiRr7XzIXjyW9UN5VToiV/yJ86wql3EKGrjCdvpK6B
RkP0l6bwULGj+W4BRxtnVl/MA+Q1TYsZK1uTfxWptF2DEna3xJUQb3kaDFrrUrK8
L0FI69B33zjwlwyjGrp/ezzhCfWVjEci7jFFn88X4tyXt8iyA4XKP3bD4nLGzIOC
pjpKYa5xug7MCMPji8mlyd+F0DK42F9hfn3akJiw++jw7K2RY3r4CKgfwn434Nz5
WvwE4KJ2+kXuy84tfDdagjzeqfJbXxr70jJQBGVHcFzt+y4863p4FRDZPb4VUprr
SkySfzaXWW5tMo6gjtpDUS7C3V8hXCfCGC6+mMg1RISF8ptJCLrvr8NKCExuS6hL
qugqFkWgo9NFNlScqLzscfNKqy16rjsfg/hA0ASGDcr98VpyGnO00IZaeauLceR3
tzt5sGYFAPMCTJVjQb/SfrcrV/Sc46SbxZV0aK3zbljmlLPYJQuhUqmGySmjzMC7
CqdP1bd2vVR+Ir4Y3hhRNlbHcVUshg2lv33iNPTsp4hSwT3ujl9xldlab0arhz+D
CdnigsaYaqTJt8sP/gIDYLLDFSfQdOtvgBXdE8zvpgLCAsw220y6AWAf4gy/s1e/
QeWUCO/q39DPa4XVyePNSaCBRMXbl/e4ITQtxxmh8nNEPl8T5KTUSn+rs6vU1SQD
MlLGiaNQX4vt7HcjrDKlZGN5VTMj6ZzTCatprSjmyycd6n4kW39NR2P3DO6el2C/
ANmsQvUKzCevKni26EH3CyDpPQHtpEyFV9Kg31E+b1lCfZODpANj0E0ioq2cGG7O
KGhUAiOkhOhMLXx2lflkC8bnYgbLFyiyYds1R4JKGYK7GUl1im5Dv6EH/0tjHtXW
uW7F//1KKfuRatbMyHUBbamt8utxMZ3vqYVmze6NZnbJLDplt/mEbR412Cz8u1ID
zP0VyWyBajFUnxuZh2rAiNTUrNSixJMF8mLjrGAGGJkwVNVib71J3ArhsfsQub7N
dJYHXYE6zHB6Qxz3QNsIN5a0Gkq6RJ2ficegUw/flBrMOuCXkuXks1Z0vadxxhju
C5ikB/fBWLEJF6TxkecaHd27wkQ72Kxy04S32plg2pun+OiNlA0GLF1/j8mCtiFa
NKVQyfY2vCp9zEYVaiHOvZXiAdFUDtBdd0xSE6nRc5I54UFKF3aXAeITxSBeT3vm
KUszeXcPBpzojLKscocFTLzYO/0k354VMQ7fSdeFrbpBjj/S9o0so+8c4JujqsDu
Krfz5VdkhV5QCgVx5+bjjrvTpejMp34zX+LCPaIIeCGchHjv/AxvuvdLQ8th2B78
Mk0IdXDwvc5RTVFWHlKI7SfTGMumnwspCLyGlOXxYVnpfmTNggtpO4VmBRE8ej6J
p7I634PVNyt3z7RsxIFaGGzfkvXwpN2XZOiHVKuhkph1MmWcb4R0UHBILpb9D0Pu
zM8WIOfLgilCO0DwLW8lnZTrJ5mGkYyrFZCrxgFbG5kG1JfrVjsOWJkZ/BqrTlHa
s+gAtf0US5EmxFG1oEgZ2WQvrOTEM48s7xh7V+OqdrAuTwNFvN6W8gOppfXk0lLS
mSBHny4Idd5h5mgjE0OmhWI08VVx8AAQ4YKXNunh1lFQHWSzF2YMKctPqnCUdg1V
Inj4D1WQTqFBSMaPl8F1J8yEyNa7+gqnlWDXA6ejJ53nGr7pSpCLDJuuYn7lt5sf
2UUs2oGaYO/EU7DA3+W+nQU4oGVfW6upigfsM09XwHXLZODnvV1uERR+N5vLx09M
cQ13NhZCtukW4ApGu3IVL3ptUd3slTb96LXDadbZZhv5p5Lq/qrW4Xt6o7xb1XOO
hAgPPr1YNfWSTGjy2jbZIGwFB1bfhD5RmP19x/22gvlqX60az4RTEv0NWV9Av+aq
JprPlRX2vhoKHfjWbQLEX/prrp0UqODIScL8Kv+VSzNQdMROyqeIegwz6uUwKuk2
HHW8ASvRqwcpQUlrah0sIbluW9Nf8GyykguhKKqjIyT+Vn9n/eeCaGv4w8QiGAhv
3et6p9ZX74qDRXkQuFrtop+FX+aEgmiavux2N4lJUjCAvnCfbvLICjrmmKUNOltz
3e98xWHC26Lgm/zdU81YxhM1Fvrx7skrWlqQ8NPMIlSpKvx4GZXA586UKpW0cHYB
ykxr018D8UVo2kDkZniZwKYQHgj/UHjlqnWiPEX3M7IW8d1d+JPbhiMOVAuV2s1d
kLqGRTs3UrHm/YjXaTCUQLKhrsXHd7z4YOqRX5ySaFGXbsTbec9ZwrB8m50uYwvY
Tkw/iF29q+yEHe4IHUk/zOzFl3llrxHC39ocFEYbcv9UVlWxEyi5tdoXpD7je7kT
gw69PllArh+Uq1JbMGfp84A/aSQCIF6KD0Mn09ovsib340b6vYi/mVu2Jx1h4Rpj
sxwKooMuZyzEBNtd1Fb0lk1wa8PhPEetc+mMGEZVKEFWAp70kqlvPxSGNwledLfR
+sMTC5EnqKv90zdeUcFbZbiSZLvwarrcrcJWQejKA1WzkVGNkOrVvsUOycAJzQ9f
OZ0tD0NS9mAxAcILsX7nzzo1cAX4awLTzVzmBfIPpKXldlryid6Rz1UfQSnYE0Ku
aJJpSMrWvkpAd1m0k7AZvZobYdDfTiLCtDeRqOSs/+iy2NNwkSyceKXmFdVTlUTr
8svVQEQfZbh2Omd5CGs3zvWkK47ZV0s/u6XWBCMDrdIScZ87fDyK+WLZWH1ml2C9
anvTjkmih5va/C1QRey564Q1PvnBEuQ965+C8qOVs8qMQRu1FlI5G2s7ooNaIGp5
1Ytmc7SaRt1XWGKSgUaGbHdpqmbDjWmFFvLzifQalBAU6m/iB3/NW40M/BNhwdnQ
9xOazOeQ6CN0F53e7IZtA25zpxlqBnfbPZQ2Iy4Plmt+TgpEogiWNCPzsGP36EWR
xASND8yhXU6Doq7to57XQ4GOHmLCYg/oiTN2gvbCxICI21HH3v1+M9ZlnRsrAIV5
gNUBKQFlPlha15zeVdT01DHLqRjQly+ZgASRYzXsTpz6g2u4KJuMg/ZVzGpu9cRr
+jeeIv6mW80y98adDSPDv8O9bo2LrxqGd39lRZ6XbqQNfFbQBD1aBwC7AQJQeYrk
vrMgV2OMndNSh3aqrrb6SqYMkbMC8WcwHyiTY/+HA6s80UF+Crbc5OyGqG7fXK6P
5L7aIL9MpRT/iq0NcCSU6zXltU4M1hQf2p5jaLdfILWWDlYnbEkGP+UIld8MN13h
s7KjRl0lCuvhkLpiU/R8we559reXuyQ/y7Xuagg1fWzEBCYsTmKBhmkE3YTxH0Mt
mYYMlxWVvk4k6ZqcePdCsfNm/LtJWLr/QIlk5PNrakAE9eptRcsmgrpXLZm0Kiga
SYsjxxtcx0FdQbMpiwIwMFXO6YxuDsCyem6mg2Nm8F16NS+FW+tcqLGKd2gUqJ/+
lWED7CQXyBMFHlO8H4H0wDfHr+ypWY7vSISpNC5R59ogsut4AFgKuOHbgH6Xmj9/
nBSxsHl+w2HiU5YJ8s3jg9/1RJJsD9vuYkjidyYAYT/NsBT3jVcaUvTX+h/JuoF0
Zlr9ub7EPEQKN7a3yoW8FDC43mQEuFBJ9WGB3luigudbhRUrc3jhV7s/1C404Xwi
3obb4S5nhOuJD5hm/VKVp4ekYtcKWYbPrwB6JoaNFyVhGlJE6jb3GfD97BC2Y+7R
cJmuAS2l6zhXjEwiq3o/FVH6xo3fukOgEKxHGdG6oYNY2tlstFuOhOxYLvkbfMDo
qE3Wz1e7IMWK5QTlo/vYT5+vmb3pXpZc8G6q0v1JHwgzYT8GfgU4sOIRLLQZ0Q2R
wqqLWKnfZu84QtkwT0ZRUchTTHQh0qafjRkGvHqKV0tf2TkzUf4ze4AkDv5dGJLx
n16CXJoFGxZ0FbpomEWCAPlP1bKXSXh6374VB++X7xYYHgwSojvnw5eDEulDS0Iy
y2graaWwDmHtMHEADL2Lt0PVW/pBHguaDSaz8frFJMK+bbs9UdQGJTvQbRvEF4Z7
e/CZ/PSUlZiLfyoFlrMWjsK8mpMEWvqCWPQzl9Oova8WE3QQ7KsoVGKl6xc2s07d
m8nUaaSfj/MzJrP6yQyJhhLOOYHyG0ThY3OM6aCBts8PHi+4lQaQdAIBAVg67rqC
0rWiQ058QHvqHb4VAwVW1r8oCKo8oVN5FKBQwYoxaFrnj0i+B91xHUZkqmJd6b+e
lWeQux1y2vydy33D5s4/bEhXB+ErxH44QxI4szw5NSfAXSUISSugKSi9rdQYLy2K
mGFF47yRacRHcgl/4K+f3/WWNdCP4n5SOIGk5cB42KfefohTZpabzn25cQDucOK1
DjFXDKVnb8zI6O7sHmLvo6rm3WRigKm6j9bn5xWz9sNe5Jk9bC5b2H5tNlx+yWiw
+4FNNH3ZIJ+IlRyDcYXuWuN/ickxsXHVDajSKyGSaLSStXQjIkVBUD2fpEIuph9u
FXfXUdRexG8Nkl+eRaR+B0E0kbudxx2Hzo61gCeqP4q7/n9goiLNn1wY/45aiFaC
TDgRQ6MXSJjrYBmO/WU4awkTiwyQ+MVeG7nXRCm95v1eQR0dMFVGQvlCWA+DjlIz
BKGN3Y5N7V/sblEKayRAWwil9A7TuXeF7JWEfjZavlsXHUvda3/VNLWZn8bjF5Nl
iKliDYWCGWvS8MhNB7LQ9i3iBPFhI3ZNc7ZQqe/oAJjLVK1ux3AaIVvOEo64QtfZ
L48O84jov4vie8IWBl4WgBGyHEzE2v12Zu2RwD1IYmFeXBtd1i0lWU78rwYMeHLs
3cMsdfIvOA4+WHTROZj6vyHuZQZJXvvYlHA9ET/7UPbZz9jC3xzsvHRGZTHhuC6D
XxVDXpjxJM3iYcnG1KZK7tobnO9Phn0hUMM0Z//W6/sVGjLpP+BG6ru5EUOxqnJ2
CMD/3lTjAaR9/MK5bEjFW69nIlDIpB2onHBXJXFVqji0nelZV+S2UwxL697+KQpY
YrP++539eRrh2OEbtA9v4IzZ98Rew1sfWYoF3wvTyoa5XYrpFiWKx75yeMf40wYz
PxltVPDFEcM9RdTEkcfJYVZgglHAXbZkqBgTWJt60iYIGl4CuWKdusaJj6LIoBSY
PXpOCWCV2vz+9yQtbMqMcmfu8zD/CoCLRuQ4s6TmFHsFkQvAL+EehloLCvig2RcK
zXm38ek3biE7TaaDR6hWx9z7uf/ODL4YDsXx+FtceDF0V+Rj0l67qNtwHXhofU0W
f0qc6+RchchVvg//ltJA2aerKUBV+VQpzUE7clb1+v36u6eWDhcZBoBi4s5s7zH0
f6AjeQ+fgzSXVGHBYVrVpNXQo10ZP/Ik8keRmAxO4Uf8YDvbUCUmBEnKn7DgeARK
b/6iNEPN7hgAGHaYWykGP6xBeqBktBNzsOOCaexdX6iGDTPXcWKmo5BPpsFOQb79
gglrosM3+qGroxCCIu9uL0nRESAOFrv3UBDDc3gd/OkSveLbVN6SsLsdKg+VR++m
OdJqaXCLOhED9llcriqD1ho9onxE8qSNWSIz8x7WuhITVu2WeDdNNY6efbwt16xV
nWciYkYbmdUXPYhXWzAgH5t6pMkntHwz585tw+e4QYyx8bU/WwSmGVzWmQrh/ZEU
0XzPJnA3Dlnk8SskuCV6AfTR7qvgeJaw4wTCHPMXVGV3RsbVuOxcBGan5u4bCMqh
614HLbozzd+39I6U//RZZRm2Xt7yAgkCACXLyCdnVxuRoZ6lqLVdtFrfa4O2l2fS
WQCx/XtIh+7ZAb9ME20/7Hnsiu+U0DR+NDRtirpXc+03Q82YlEYd13VlVB2A3BNH
eNBvAFT0PF/jVyHUgpq8239Y6EW2fFHcB9Ql95jecf6MZ2O/HHGlx4Ze9A5+U4GA
Xd6VscYT/71B1x/L4LqZvR963A1hC1FSax0635Z3gN4K8LrDnQt9Q2oVsswbpD6F
vrQH9tL9PEUjumax6YQK5sy9ZniRNQx0jEDCKTd1HQAl7NEix49C5IOKF2lVpYSy
J/VHXM8R98/NloEE5GSyQgbPfVYlWinGCNWRMl7af9HFor/XlinXFAlpZR8+FU9K
DHC+hHLyyb98FTqL/2uXeMoNZGezk1rLlX9nbhFQE5NmI14d8SA+mhd47lf3zeVL
tFIkKRYedvYmz1loQAgFKbFNiVFWTLMBpEDm+I3CAXNawTBgBH4aWcI80buFFFN1
uuQwN8iyDOTA+TmrscskfsizI5TCjqo5eey7ShaLG8jwI8wKB0rvqOWOP9I2V4nN
bVzCKsCFPvU5a4G97ko9GEIfudZEK5PDra6ymFD0emTtXtCpwW9PgDT5JbrM1lHD
wwriFSxFuwA1fnGL9n4C7Oh+HRkF1CmZirHAblecjp2fWyAf3KrOlhm/LHvO4PKb
nrP8bl4Xdh+T4HaCCh6Tbb7nAM/vVpYrJs2aWkiS1n2EXt5jahm7Yd6rYKHeC2Ra
ARX941M8KtJhxGeYd/aRnplAGJMOF7tf1rRiMNjsQ+ICxHEd7SMsVfN133fXSHpG
PHpUfgXigMJ9XZhecJLvGWvYdI5UTDe7DSHW0m6MT1jAVqQAFXlj7k8/a1A4Fc8l
CIoB9Tlhc6ro/LKpsSj5Foe6ovz03L8Oc+A8Adk9OMdtbq9qiSPti7Ijd82SnVBG
EjoDexwXfPi4hMIsMTsjkaw7NBWEWsNY3nU57riAfxaZPYfOrESqlfUq41c1A35s
br1pFHPTb7GAMm4zDy7o0uhq6MnSyxkNcp1qsyYCuiygAzk+O3E8GrGD+cC6TkJN
IhI8fJvMbZGkdIDlwkarOZ/4tQYmCEvaWI2TF47Hp1bWfNMqIFI9qR3fmAL8+j5o
rfC6qnOqfA561kEBqmXb9t4HWan65Ig5/rtILU/0xf4scXydrsDCb0xMlSM+K9AD
ZK2nJNhdq2xaKfyRDxkiPbUHxiOSwWPWMrAU+/So9t6+WpTJeKdVU3soDGeRjuAf
ij++nt5vaw1J9BARZGGsPjx5zvYbemXG6byLkJdAWAaRKfY4oQZlw9bnRzu0jJV0
StNhfeAaRXzeb8eP8QRrsAe0QCgrnzvFEEZr8cTaqbGV/qG+Wh8DZYr0ZatUaKUX
sks5rLTbMS6ld/sJPN+BbvRwE6FSM9tQUUjOb6B1MQO+D0DQzDW88qoAiFDXh2I5
Iel7zXAw8N9Lz1o0TUMJNBCvs7aoujca5IIM6Twq1SqCuuaj2U5qGzGzSNnpKbl4
RLbjGrT1eFTRwHyIjhqvHBvY0HahG9FOWuJ3fmUr+pesMZDcJtwGopFHruNIIErc
pw8NuXgdxIgftY2iuRtSUHd5KRIBcnTtftJEVCYrLPBPMF5kEUQB/UxzgSVnclVN
MPYIEUlN7Kn1Vegq6nLF68EJ2jF54Quy3MKE7wH3DaPLU/wpEYrj/kMp+gaiEhuk
bzMF9mprP36RC54LAa3vGMRCa3TM/tpSkNUHQEhs4lAhmBY9nJgM9U19FtmgUrOa
0karh+7nlEqvgVIyvm2uigQJjDV5tVqXdZYpeiAeTijYiTNYiT0Lz53/dN1YxwEX
46Lv4uSdBXSu7sTQxQPJrGlIWi487jmgfZYfXmdE5hBEaWrp6NMjKjNNqRNssYhP
Kqc6/1gvGFoP/Zy8ixzLCoBsCkfGukbswa2m48lF22GlErILEHJ/V8FjFkVh3lNJ
OeWlL60do3ONET46iJjh3X7rq3n00ASIYhpjTIMw6l2QK8C8xNIf2B8jzYPKbsTu
xJ1XqNJbsMt0GaMjPYAGPeokC4+RCQu55H2F27KFtEFwcolFou7KtvmiFwAWXU0x
stk4U6B1uzkMzKa3+HdGNHwl/qhb0cirxodhnx105o/1VnFuBZJDMzgC+LFk0sL0
TBHxtVSm2RdGIYgJYR7kY0Yt8BdhJYADhWq/z4/gtFFC3vUFH8SEkQ/Jjflc/WhN
1exUuvQa8ATkwPmDW+xI8U9nTiFnEw/ckJMZx4ixkjYle7t6JKAoWh0LmvjnGxZC
CIJrLcPORBfUPrmCOlHUUKsCECmEgyBNBGjIn2gnBvyfxPKzwee61r08nLjgTFUA
LDacgnoeA7fyAHqsFCzPWkRnce/Q4m3fSOSP+PY2Q6ST2VF7+ggkhI+Azci21oqO
edwSPfJWMjZex+FyCwKXTeHzGqWVsc+xZGg/85o1EnJfk4nmnmSDCC6ay7cF269r
N8QmaygywS/Nn2IElJ3IwRaZ5l35ts57fszNgs3BIn2JTxJKxcyTPUsw19wPsKPd
ti7ZfAve5/VFkY/dW61kQjVvXXQu/zMTxw8XWxH5iW9S20tNHpbkPTjEoAx83Cmu
U0ivFY6AZHpIkWiQOToLYnSLqFd+6HA9RBYnHjxeQXYVAOo2fg1xwlbMboo6np8x
RvINvZ4vRMfNq/aFjEVYlQfG+wcG3Atl4DL6b7UoO0E9kN986SdfJXUXLQITtEaj
JQMlcYtyCcGTDfr2Li+txdTcaDFutFE52Za39SfORnibY/S23P1+Tid1utYg3ilF
0VVX+jDgJCjowk/yVT4zBDrmg5AKwCx/0QTBc7qOg1OkjEycPyKDPE0L8PFSJOTX
OVyK1b98DnPcWebw9swnNHwBqXyahWoFdmPKgxCm3VRxZG+saAwzhMd7HfErLDb5
Fn1WVpyZxbQ9YxBVqdzjenYApQxT3pIYyYS7849BkEPN+vPSGHbvzF5eCzBYUiEe
1SVflsgm6jXIZmKwUJbBLSsinDy4bKeE6jbEH7ocHhBqs7vYz/8h2qprsRxOxjQm
gh7hLafiToePWypjmQz4NET71nQZSpPSh91Rtvkfj4+exbUG9vuuNL/qSkKBinzK
jsomHugtIuHeU9fbBs0ZX17FolYrfYCY8vKwc8wtaWBEGJ3gjm0DCkyp3kj2CsCZ
kXwH5sU9mr808/n+d4yI/rrKzbbPW/P7yQG900XVdGM6DLcHJmF1J6VTQfAOfT5P
Gco5CT2+A23Z80XSvZLf+qdzVRUZvQy18PiRYnIH16UGdN8e55rOkvLvoR5VwZo8
P3rnxhxXsJ/nEV5iTU+dgToLLyHJyqU6BvdXrwFbDxK3v3P3O4I/O/yM+Wu9+ZHZ
nh3CvZOhxtwzizL64im3OQHgAz6/yvyMf4YB6NtagDqXcjoGYf370gbKphskV8ku
2BxBTPNzIncf3SjYSHQRYQv3hwnoTntj44qBySTghOBR0GKM5ddvdGB1zo+Bl7GT
JXzCtyDN08aPKpCz8boFe1WUieRAFMJ1oyFVqkC1/X47iOGHhvKzlj2w6z1ia1/p
iLWDbkSYKxsO0IDFNh2EwBnpjSB+IheVS3IJvk0vYoGoXuG8/HGhoawdRVf3lwwn
McwofSU42GeckFtOkl+RQD63X1hS3MXzGH6QHvgaY+W8TSc0YeC6Nx2LWz421Jlo
lNCZCaOZLrhc6oDKBLQaN5bGJuomhoC+NSAW3OZQGTGD7gYyzjHwsabwTA7WIigl
9p7HRfoHEcFlmO2wr8IaerlWTflZdLp18eV3haPdz0ofBsrRQXYyEyg49CXALj3Z
H1xw8E8Pq14BMWL1+FjhraHTidTIPtLci/BoHX0TRzycwvqE/e4CLLXdIlxyLJJ0
o/UuBJ9elFmxlV5L8QD5OGUfVcAK2JHUcb8i6LexRXa+9TRdo/3h4V+aY/rQB2Qf
v+ME9K8A/St+1awRQmldsMhqAoIeRLO3QbuBIoBCO0Z594lTgZ+k62DhEm9bLqpg
4A9ULDm8dqwKsw8mUrbbZHpNLlZmE1ZZzbLdsRXAeKEBYfoKTXzZEdjyPmCAoUEq
xq+kKe2cR9IFGd+ZsTjGIAB3VAboNs1tNj5/mjVrgXWZ/QyhKK3dI6QFo543DqJe
FfMxk4Y864KwUxdkJo6iXYECshdSAJX5d+W68wIy0A1W96vuGn/1lz9jtg2p1Vc5
/XLhtijCCi9ceectOsuPmKp8vYYEAVNAQJq19YLHLvT8mtg45rwhRrRbrrlvd9qa
WbS40IWEGVinCn9r/B8IPqnGvN7ZvcgTbf6pkqu6bMQT6KDIusLUqEuT9JjH3Q3X
oAoEx7BwadCa+vdRcXI86+61QgucmssdUCHMjZXXvzBPUV8mPGF0U865V5rhc7hl
xUMgVi32wq09xrr+Gdoeih8brp6/h4uIAJdptfyKID941qSzLSplen1FqEBtlvUs
aYfNseiUH1TXKJACmDGKb+U/61AmVziBLN7W+nWlSVMGVRJdsnWgWWcst33QmJPZ
h1pOKjWGsAykIPWetoRQ0EsQVjSQjCHRph/0lZjlCIFiPyR8DVIjSb2PLnVowny/
nMd7QmvP5dBXL2NWe0aBWM5JglT7LAkLuDQ0Xfd1Qb1RFYmsofeQyMa07FslipBu
NvfEjyO6ie9gV2Ui60VxvxfCAMwbutUGqJUMOpS8nGUfrHzxzqIT5KDRw+aq44yS
6DAt4zwLrdt9gDSrKsUIyoBIyKi6R3KPMix15wcAIKN81Q9285r4eUlEGuiJoZGP
UgVequ2gS8EytueqdduWVrKk+ECAxmrh9uOdnLyeJg4zIoMMwe8+u1TIYan83Jza
8TtMZH6HffEmiL3NYU8NVeM7H3CazpvA+9LU8+RS0Ff7J8gwa8l4Rj3WumgCiZr0
Fur1jAyVLb5Xlm1qzocS6mVVFV1R8rYXJ0a/ebgZ/u6WVaJCz3V+1kbJGeo6CfMO
dW4WV6HlAHdanVnmjEvnyy8qBwkSocp1CbfOPiwxCdCheUKwQziZ19qXlKFqZzgb
nBUtVK2/SHn7C1Mr4kbTK24iibEC2sx4NFaIGwOUHgjDkDtyxvl38/OMKNWuJXUi
Vdkh/R1CtosT5dgBVDhjgpwPcp6MpJtqYQYfcTCNtdrzo4HoE347XbGoJdAok1qB
weCj1HyCL0qxzA9qa3RMTST3CWfbsh2k1OVcrDnvt6PoM8du5lVelmVPSZaF8ZR7
Q332boYBsQLEO3FUqKaWuji+bsPi1LZjCVebMCQ5PrNhq/ozbGPMP5jvPzRbOXhA
7QjKngoAzh1rgdN5DqGXbelMSv2yNHuWhgs0/44fP5QQ37429I1yDQYovKoQn8YH
BfLyx9UAIjL9uoMfkuBDgFPGLbq0XT8KR9I0aOF2X5fQneUPUHtroSKD1Tt5tLw+
gc+WVQmzjvFAOfeCu4WG8w3NIdHME8voykPHbtrudcHKLwA15otHGBTn+7NVBC1U
BQHAaU9J+sEdPXKhmJvHZVMZ0xLLMv+o6I4dhBBoTatVSAMmJRkzyYcn8i61ncW2
mGSba3OZmUM2ensQudcEOf4/Of9v3mYc25R3TdyJsWzuBbw7AOzW9HHF0i21jbw3
K/uMgd3O1Ia+vBfkiUkrioeyW9C4s1h7JXQsb+OX0i0Kt72eDxqEXHNsIzLz7tVe
nnwK8c0LQ0zgDGuoEOUf3Uh/lADxwapaahkCt6jX0mV3+b5BViZgBW/75gHgf4Mg
p23Ae0Xe5Xiy6bV+saKfnCq844Wk0kB14RKS3mm+clkWd+sMC04Vrn9X1SRt7/B+
1Mudo6VK131h3yGC1vVdOh7yoZVj39/sqWZZzFoR5+3fenRKRVAeXJ4He8nrl89O
2fJH4oomnqMbflItWlKWbPQYZT45MSC1Raob6rwwiACKg+IjjZvTQx0Fg6MxDvZx
8i20kqUEJ1R+/wHDBOtLtDD3Nrs4a8wNKiAqoTm9eTMmwP0kAADjHM9NIcYZXGbD
pHKPFaSH0jZjUcs2QXFL7K/bhaSEftox7OSo+zInTJmYRIl0N8+/edFJR54eSBZv
M0xe2PZaj2RL7lC6Jl30rKw3qzcX0lr9D475kDJsNZpVlkfkgDdwmSNnWQA7s79z
IsU6lGQooD1WLyNEvZMqo3Sdw9O37dwFSiQyp1dS4Fe1YKJX1QNLvV63EqzWYAGm
Qmmostk4kJbHO13SVAH6ISCqXciVlAelO4IPJXNO84Tezw9/RdB1vbQLGdPnOVtw
8ThmaIHs6gc9vjaVSmeJhSDKvp0+ZHokTCB9XJoQzIwPaPJo5rRey1XcG/gFDgGS
8IEzoovzr3J+MWVZzaPPIOoJI7d7kJmSbl8ftOQSKVHeOK9qva22HOsFKbsP/tc4
WDzBZmJyIPGa/ulCetzuhCy5il26fIPyLFX46R6DNCT51Kw6m/Dws5CjWx8PpQRB
dWDN3u7Cu48fF8f30/n7KNMv824lQtqDZHEqZlcuUZ8gs7MDpCCqacZQSi91Xpvd
WyyknwShatDJ3HyggxnP8jpqHMW5xmmdmTgHJzUDbapMdJxZOhfJcMecRh8HtTNX
S48EGkksOrRwIHqSNOYmy63Ltsv+iX45/uoHRXomDkMHTtQYpb7Q/QJsAc0mHrez
G+Ag7KT3X+oGqABuqoEiAr2C8jbWQmZxqtJ84vr8uw0hEF+DLdSUqlkEqg3BxbmW
Dt3ow3FjW5mdsoKp15Q1Qu8UFNHr+Nx1QHTKxC5IDfCmRzpxAJZekVquU8X2Tk4d
vMxYb0B/EOniZFSV+C94pLOLw4CBacsjFTMRjKSpWcQ4txg4GFPY7hnczTxNTmuO
cH5Xn/+oP21hkLEcur+MIFsdfvE7oBhekHQjdX1P9ARCav+R1wlfyVRjcn95GH47
dXJejhkL9+OkqWT1Ef672E0jUpNMSMUwNfHVW88p20zNnf4DxvPJfGLCU7nXxLgl
TYuRUzgBvTXM9OyyAVpxA7aFAhOUgJPNjwgTa7MNAnVwiQlDm5BlUS8DxYsbdelW
QclEMS8SshBwa8im8wuwD71WmAgRMrGAt2GdiuXavQdN73wD7Ufkq3YBq3jFu3hh
YtmjcMk44VOYMAdP4gyk6xCXSHhgFc6tcphsiL8S6STaN9JAtUQ3+d+AluqvsGm6
sLUr5Ob5EaMdy+tfbOQQSf2SgvFv/Q3yn17YygffAiJvbsq2FiCAsKF47IUjNsiP
z7cfSfd8/ehXT3uEv2HkoheVf2xudb/iwGIQtDuAzUm5uUzL3+Yi47QivjGpRKsM
P3Zi/GEoWZ/S4Y7j6ifJ0y8aQDLoRdQWZwmb15rP+/vMLnwfKb4qnskCa+oy5Cgr
dAbv6IuKnG39G3ZjMkGNktBG96SLGfq9kQf1LMNa4orUe2bO+R0uLoIG5W2mzpbW
WhyiNo7g35erQ6sm9d6CxuauPIUxaROCaLmI9BgO67/3mcCA4nwpYe9ORoCmlwTP
Dy1Ic+e+kp4HKSlOLK7GfbP3h1tm6bahiBkyXySGnZ6mD9vesmSxrt7v9SFtzw/+
xc9401L8I+Q4LMKPOq9VWmQByaUG/4JUcx3wtGF1kEB1dtCKjRJKsGJ2NAoP7I0s
nw0kMHOOW3i1moWL++qoryK8Z0za1OtFqB7g37pM9TV/RpGtoNYM4khr74kcpdWO
W+VlTqxwMu42VaIcRTyRG5TqapHeK6kmficzJbnsX84xkHRNDPzBiL+hYKw7Wonn
VhQX0OyDXIXrq9GAqZGEtRCNVbcuTSwlXzv0NST9hYJOaayRH+2q03KkWxxai6Vq
Dh4QAXDysySZv+QidzgqF/MBGrDlUTcn63sj80qQoB1WsUgFZSkQINwAT5YwHfvE
9U/crjNBBQKjja36IByTUQKzK/Xk5V6n48glBmUVQ+yIT+yB2McTGG0EJ/T5dp6J
cXL+ThGXVDLlFXANalKjFM9DphgIuzv+cFrGV4I0TkD5/V0QpHLxq3MDKnZY5ovR
q6YbxyievQx0AJLYayTTKBUJHCITfIhb0WJHmgPmYk4O4xtzIiMrTprP+Ymn/QpY
P1u/2JGDDHm9GfNLZAZQSBG5KwfkNPb6q7+67bnYt/HfXUOumXlv+js5TbzK33v7
ex8eTGtUnUpUa6Zd/4eNXSg+Lo8W5srBXBEZkke5ln/OaJEP9ABFe+goQJNS+r61
D0JXVQem7AAu4Dm/Lz6oK4LZCcrCiDVYMfzOrWrdWYlzcE2Dl/Fd4YMf1TAL+lbx
09KNjDsfofN8EcgRsJ863jeVRqwtvbnFh6DLVFQ+z1510+zvCwZp52+mc0x5MNox
PXlY1tLNeXffctSgwtU7dut8o46rR9uJofQT3OGqFCLnkvMJ/Jrn1W35IscgoD9J
rW8AZ02VH10yqcucr1FNPf4S1piMkgMByNibq4n4Rfh/X+YPUnLI6P3OEw4jOY/6
bMtZHFZKaPAcfqMlJej5kqenp798rP8cDk9PCfg3Qmogbb8wy+uAiUQKFbRb+IVh
IoRO7RdemRlXBsd4AzQZwThoOrlO7KzUV5RMmGJV1aqCfS3PA+ifSdCzmiaXZ+oa
nBWmo+wFebQjeis48n77HZr+EL9do2wikpkrNyxg4YLLPk8nccs1t+GfusNzF0uq
/MXIoDOdaQBz4atGmGTosXrpkCJPjGF47rXuY/MNVRJz7nU5/FA45K+kjJwL7ef9
RelVH8S4WqBNZwQyqvnUnSk9vQEDk8qtu4RcOZHY07ddN+7Oyo3rnBxITE9fbHZ3
ByiC8MYb/cbXobUBrcxkmx8/vA1AozsMLWl4SsbiT/mT+h6wShg4sqCIohZq0L2e
uSp5WrG/s9+vaAh0saTZuT6BuY6+0q82ONtABLdrtS19TO+BtAL3b+PKOzMKMg3h
C4cgRpieIKoqM5oSEes6jZCBXWyAkuIv2jCRZJF0/gd+CkIAQ3MgZ2xDRlaaJjnP
yCXPESHhz884gp4Lv5f9+CnWc9WGh8OnHvw9geC6RTr2fqFYPyyKSUmZpB46IOcf
CvkY1n5wYMh/l3CDY2ioFbPSpFFZtiITFEL56j0COmIBFOPVIa+NuZVytpCHWq1b
3x/5XPJXAv8YECQRa+uvyMQioae2OSArpxbS2nV6TgbUJ93cUpxveOdOOW/FxKTm
rWF0uWQrz4e6qfgVPoBeA5tYbnRvUIbt6S/Eesz8E/Zq72WS7r48i91t7ZiUl9g6
3EuridFXntS0w33Ztwf1b2qzbwqXWzmI3lqgjxzxx+m1aNVOmQ3L090oGocfDdWF
Xd6s6Zj0crgovUv0b5mCcGX79o608+/gjgWFAeoFhUoqU9Wz5YEwR3Qjt85szMb1
bkALw3M2tZrGwBtjWL1Jb2yjtD7PVhyR8kBQCEW2vsJELRqwCEVKxJxVs7hPlRMV
ZxELJmac6Ii2WwDH5hE3iwn9TklCfLNzGsDlUH6w+m5kdDxOk8YT/TkMISRad4Fy
5cfcCn1k0PR1pVVwN4dI/irmiLdIc/3zp3Z7ljiRJbXfSaasq8IoB0l3B+yfAE3h
pNSXEOz5q3Zp69vqF3fTCIk+ACxFW5nF8vO/Oyea8yTuo0cJT2nyCA5JRzmOhJzu
/asunKXtqn+O4VOb5UvWfokFk/H+e6RZPtnfyeEPHjjRtR9908nDOQ+OL1RWa6BK
1PiksoXtYocuoGnpPcVreJPV81jxbACVAKGWqIb4KJVZCeUDtNVk9KEoy1syCwTs
4SWxEI2cxKtB8n3+EVV0se80SpiLCIsjAQv36LlQFt+0KiMq97n3vzOCBsLahUuy
BL3dBkUtvB5p3/+2AMaWt4uBLnM0GAi4uG6FLGlEjuu5iN12L9/jj75qQc0X76/H
r7lfjH+G2IfVs/jnSGw1/ARhPiwUmpvcOexMNrOQ/lGgqOYQmSBAAKrPmpjFbGxh
x18Q+VmDrHZe78B/iKj/Mu0Lr6iEl/5V4lMZnJLQOtKObvRLszVXFwUtvmqvfN6+
sZQw/P9RDN6RWMX8SVb+dTf1NjEH/IiSjcMRDNycEZ8kLyhaoPv/loxHzW2vGCfy
84HHVbJATzFO4CifoWmeL+HG9p6NJ2HR+1TyElA+TfEgch4hWVwLMk6JKF+nMcU6
l3XB3xKDlCnimzvuZJLRgkVq4Ul24QrG0SI92DjMLkMPMHOaeGr0cdbxe4jAOSOO
UIS3rh6oR7ddUICqaQqvqS0YpO4n96IBTBF6dKFK/Z4rQsJjkHL4fSMR/s3jJjoM
IIgah+6jjRQjxmhcr80dJUflq6zBseFD1T42FKA7cDaT37rKEa84bmeV20BnoXhb
/6y4NbJh7Ph9hyXz8CuUVlpkL/j1GDW51ImTXYghRMbB0tLBK7G+ZGLFphBSeL5y
UtZM+l0+1l5cUARS7pf27N1zWOCiuK6qB7k9vXRG8JQpzMHwFKyq82wMWyAqdMnv
9tKhs2tzDelZLLdybIvpiFJUj+TNqTh9U+JSIuCRW1tRhte7Gn4kYJ1cIXBsApV4
E4I3FG7dyLU7vHZLF1GYTsJITen41DinxlRKMOzrfQlSZG6Fz+FghseslidXdwHz
AIiwMxIllMDbWEN4k7Mx3evvw8EjkwUvLLDrY/MMO6XTIp4RUosVQhyNlAzbTNkL
7eDbzqTxEp2auM9datF+36jQbbRhjd05UikX8leC0lxeeoiQru3pGbAihqARd6EA
v4KJGpqRgRmyruCip+pegcTDfWloVX42UhNQBuClNNEEpNO4TePyJiRvwhXt+09p
AWAiD93EskAlQ7H8c+g2KPIAQ36GMJjH8jiG73nYj2YmYnFQUZVhRmOGjNCzX7mO
N4z9VqTcKTve25W2ha5la2sKPdGabZ7a8ybaXcUM7+YaqZ3pLN0NvRM5eHjBaZwy
/5iUy1wJ8+sxHwzWA0ghHfivlYpzJwo1dn8eQSSvaN4iCJptqYpH8Zjo7ADtGD/8
t+/Nou2amGeEgk647IVEbpp7Emi3aon4KB8vvgJ9mr0FPSAy3N74APZBS+6/9Ydv
T7Pdyhow1i6uV2Dz+z66xWCBqtyxdpLlvcR6ku6CJL3LtMDONHQEtZPFlgpey21y
hE5jRCJWMPZvGE4C6an0A1xJrw9kH8Ho/98TquVj6BOrwbuqnEVDrJnWWv1ipGS8
hFDYvAmYYwVGM3WQqFAmJduzRqV+zUAEmzYiyTT60+BG+JDEfFC1BcXvGOsOM62H
QkrbKcE6BLdLgprd2Qr62/r8+qtnpiKn8WvuCguML4oLvQL70X7uafk5YHHmGGgE
jGl25/BWQ2V1WDoo337zv8qQgdoNFNMBIKLTnu9omJkuAMWjjH8ptWEvk/HsgOXk
RsWPMhJN55vDm9bubGNcBZb4JenKilOF1l+2+bhyho1i9LndH65HJR9fruvrFTUU
WxX9ThC3c6s0fTDYqJa1VbipaaK6pslAPhorBlfAtuWY/GhkQ1UmNiR+P0dTAMVF
9MK3Aa0Uqe/U8oN33X1zmU6Ayjd//UBd0NYP+8mOMap+VXE7W5vSmy2PdL1dfEhu
F5bogYZbCfYktBPe3HuetelLsZLAU1NkUbuuOm/XlJcvT1YiFuqr2/s4O3Xvk5+e
Lhu3AD1FJJ+X0s7u3UQ1bktoIAfVl0JwwKOnAbbaRovVQoMZBQQ2bsKNWVCvVs9h
BJwn6oFOgIFgjUo1wZQTUEyG0A2T3k0GEEJCJWvrWwOR7lpnLHzR7nz1d3GMLIDR
6bX1JNVN+PKw7Qn+23YYn3xyQmuQc16z8voEghz9ZrBl1g3W+NI4LqqDuYuERuBq
s1rbbzlh+1dC1qNHrIdB/IZyxaGRXpDwiUNzdh/FDxr8xA9toDZwjjZBqvmyUFfW
Qd5hYQUw2d21/JAEo75ovc4doNOPXvHEjxQyNpWO/i4IBhjLO2sGz4mpWgeS4Lxz
MZ0IinJNhWvJtN41MRnyrXnwEOftA99+6uOSjoVqT0bJUMHQ1lLMScyLTrDUYfFs
ZyixCoPFV2FNjxMwVTeDIQwd/kuZvNzkgk6IXIwsdw6rHuxSZBDHhwK5aWCsGmyX
2FWt5tjwOhWU9Iq1YoN/zKPZ+mHEqFlngop1aSHDsACPM8SGYnVwmS0S3Aai/I+/
RsnjIKFlXxuQqy9fBTqsK45zoJaodxwFwwN48REDyba4nMXp0W5Z1kTk1mx60/GC
twY2wSG1M6kZ8OJQSi8tnjusVWXopgR5FiC3z4qKEDk0eeSE8q2z0yTNcbYGETLH
hb7rzo2ISS31e0g9aJapJHblarvHo0QWy1VSD+8AJ83TtiPBY1w8/hqia1GMbvjn
4JeUHMw35kn73gPltG4zkLC/6ReOg5EAUqGL/ugjkH06jzbvoBD/m6V2BVN0FZD2
xjmA8B/Oh5EDqfY+EeiPQCmYdGWNizjrsYr36QvVsjThMgVk4xdt7Hoqq3T1brmz
h2VUsGCWqzhRRmb3jeUi3LVI8JtIeLttTEsxoNm/gm4omRgN+o9MumcumtOZfc/F
0LTLwi34UgNn83Q/x64kmASIYPMKSBgrnMJ2NVmwBVDs/lJMtH8baWPDwtQQBI9n
vDbEukfF45T3TsRBbKbm1DkAyxRrcr1TPbUDU8HDZZv4jhE800mzcqyGyU/r2+rp
zXkHuKVhHrzUzS3xIYKmFDvNnK1XYlvqXyn09s4BBZOV4xxrN/HQeYxxelcnXzo4
B8MBqXeKLh+Am35zynSlkDIXMP6pXMPL3V+1vjTS330agmYu6cpHOZrA60OwzHig
Cjr3hCK2bk+4dpyqvenoGRFbHzAazXBj2of7sO8PzhDAFW9kBdjGegBzY9aHwPM8
ocCPsq/9F6PAfK3wi0pyrSbOLw+TtbWYdbikxrvp0Qk94Oaw1C88plgdJYMerVlb
8/TFeTkhG85e+hruU3q7G+FBc2iDDr2adpMZTmirHltFuwLWL4WB9lYXLSEZrMu3
UmCAvDaeRDm/TIoTKN6AdZHpJjWqty3BpO4uLOyy1zv8AOM5SDkzsb/Te+VdEPuQ
4/eSYd+f6YgLe9C6UBVt5XfOBFUk2hnbvKIWX5pOJHqQKQZPtkWewnKq7XnjxoMX
MrhFWpkKj8ylyx1hXLKgu0GoN9JfL3nGIL/WXm7SojTXuhCNn13cS5bDgqY2Gwz7
+Jq30IBu3YCnGmICrQUaU9xSxnPYwk+ZU0TrVe183wrMtK76yuguhE15GRgAIhrm
ktFm6cd/CVnX9zSQv4dvUBPZEj4LN80M7AsjbbmmK8ixlFE2yrm98YN43/S3BfUE
TvTcxcdXUs7a0WrqN9MqOUMfROac3WI43AfY932X+etHS9faZ9N6u529Yn5bVeMm
l+fLd1hm38UtZXjsM9uXyrURSttpfxxx5tyYpDwt439L0/qUG6oZ34N7+FIGORn1
eOA3NuRyapVdHpVRzzZ3HTPkY4vE2ZVoL29UwWgMW0a8Er3ljraLYEhFBCP4PuyS
IzD5qYeoZFkKnDSP4P1RZsagDQuE493MmQGkH54QyLOWX4YAHckWPWCyT0AbRQYw
doecJRrPe/euqr9gHOnfqguRJV537da3XcCyM/If7d5yqHk5nZRlyyTlduyn3pD0
oGwJZyTAVQYDIQsrO0aXjHLNi5R6nmytE4KeiHlg3bAvU9b5WAS0GKeLB1xaAMmz
ZjMInKiO2RU08e0OQpH8kDo9vZjSStuGTGasV10Z1r6BYtHohzbPS9BNQQmaFtOd
38aptRK0xVMpOM4pJJNp7VD8Bm44ZwRTgHNhbrBxclgMZUJhS8FMhKHFdJDuJC5g
yUV5YOHeWbq2+sAd6gu7PHCBpMY7dH0wiSRlmjYGGlfVuOcwc3cFKPC4L2W0rlrg
OvFKT0YP0dCH/ElL32FPMOGmitCteB+7BT5Wa52GoWl73vVyT1rQ8lYQf+5yo3J8
1gkWB+4KdLeT+DGsXWOSoa+K7pFb+hY/PhgFgrMuswLHtY2/1VzysbwShwAfhglZ
mtQ8w83tXyK/S926vlDGwYVZdDqNKywI3rsF18iWSdN7XhsPowY5g8di8LHbp622
agLuZytSSQISV9foQn+NNMIfkTI0lZnDpdXeLj0OvCieG+FpfbIKzI0+dNOefgja
+DYxI95e4RsJBsGiv/MXLIVylrpgv9iy695Ay0pXx+ghaWtODKP/QGCQgiJ3Gk9k
u8wlgh7JWhGhAahTrkc73ogNU9J4fW8XanDyOTuVdSnOQ4if6LDjpqApt0CqEpjx
QZY3XjGJVi6mvKrWpGW27viHUSIhOfwufMfMmIlF22FYYnBgoqIvv8AQHB9FIl+Z
EXzhgQ3cWUD7v0ofIfQ5i2FfnD4d8OZf9hElPK8v9kO8N1+nyL38F64YrJX4LjL8
fQ4IEe5ZSPAdDOuhj/KjujlsSz37PP6dGQ3z37NrFEb0c7l+1HcJFV9ZsF7w1T3O
rFlcjiKOWkEA6ARuTG2x9R27Q7m4580k5ZaraalbZVrVEcF7ubG7UspYzGl5EEKn
yhS6VH3osHVO/Hk0GqOOTyJhLTcViHk1tH8A9dsjYJaJjLgvLLkYqYoTl0C9BCdl
Xrv9wVJUOznips9Y++WKySsr0Y2uhkZgOBv8dOxTNHoRkKevQMe7zP9mBOZu98wz
Rn6+foiYYFhGvY1oEkuEaJDGg92jty5jV7eU4MtNJykOjc3fcgABv5lg5c0XlWuC
wLSCRVHAbAVBAGrDMTh0+7/Ij2MdAzTXtOAvjDPqIIFmY35syvWAhFmqvVe93bn7
GA2hZtjHdr1j3ilziB5MNlhXrhKWjD4Qi46DDilr461MFegOyONuXSk7XzYaxjwW
Z3jeZeXXODeFPpi0RSbru6xEJcn97tzto7gvkKBTfWt/5/Eh/cI4Mmg/18MeNPPe
QYCj8pKldC6PIZ+0p1a53oG8LercM+0h/4Hd2bDwbAcKFGlMOgEcNzpU6QQru+tf
Tyq4wial/XAb5bRYOiGeTXpoXVVGLe83jR3taTBdJkuaZ/v9tjKYhx7LgvUgqm0r
fl58JYw1rW+xxYCUkjOjL8SgAQOmEUFTm3Nu1ULg+ZJ7/OJKxUldxFZBhdAD3HRH
bJ/KhblkOtdR31ZpnH/yCQZAYenexNzMht9emojpQ7eHFfqMVQiubQ+Gc0qM9ZbH
uu70tio17jE3zGioAIzghDqNLegtj1ceh4FNLp966X9hBRVuW4674gWRze+hSV4q
V5AtbANmrz7mfcu6+RrjQ1OJMyNGhkHXpQd2Xq/M3lNwmpE3NydLtEpHpWdHwDrL
wtzBHGXFcKIM8mYojvpsao5LZerF8Dfeh/b3ZBGW+70fPp6mTGwycRKKcTmt4C8/
ZCCtNaUSBgV78W3gp6x46kM3ArFXNuNQlH9dk8dUXWX4OBZ7I305vpgSg20TIHjV
I5y5m0a0OP2seRfy+HIX+J25OGcDG9sFgDtupEfCaQsLstZnIjEO9ND2zRPj4CbH
txGyGDrghV8rOjBfMJjN/bDAZLbfETGCrdFF6Oy+Lv5j8o5Bfr7AUS8zIl13+Td0
dBZbV5x+nJwAWYaBaEKbO+3Vig+Qph9o+zi0m4TA+G5LDseaa0w2y908xu5Va98q
U3bXnao0QVPlQ2zSR5dF3SdbpGbBFFjTgNDKD2Te1aEx95bHjDBdB96muGQ7UUE+
mki5824GAboDzrnbfihqjmPlEeCJMMLnVYyoiG6QSudIb475AZcWLohs0+esCXUt
yxUjXf30q6WlAvhpzZNdR/fSO0kr6h5UrgZu+x0BOo+f5r/jmkMyRxxBJ7DynZjL
fLvxVDyGMdip8vfAK6rBd1rYHoEzNA5PhAJcQvWWZSELq4xWMYmdiju90NWV7VVh
LpGDu1TqSh0ObJtNZ1ZpXhjaxmQJq4VQD/Vrn4lddjMEi7OjbhkTYSP9+i663B90
LQPD+c1xqIbB/97ARIERINx5/ifiR2X/rzOSfSjjT6StDq/ZDP4jQuisYb4vRcDS
+Lh3wWqHd3lUn7l1OTHlcKAhn0RYHdIlspzLryVqKOwiDxxMHq72KOInDGBJUP20
xgDj0MYvjed+63AS4AUXMTz5TxN1B4AQFLi8Uij8lAUDzdkY2Pf0OTdwoFHpurlA
JzEyo0EKEsW/J411jeY+XV5s9cBlE3w2Mt6CD9RoLY4urDB2xCnP3E7+5FaIioeC
025g5vEgQTTFaYXLnrP0AJU3mcxNmLx7woVl1k+Ho4Gl8AgiGDUd2Q+BQpEs9R1H
AF2MQZ7HvcvTdhZoC0BO6ZIf7jn86gyPda5QkZVBezFJvVOeTKBn4Vh9DBI8PvLM
1aDtoQx3tlC/BlFzZ5q8MlrRc/wM2BG9Dak6kJBXqfCfFfgakwePe7EGC3MNE3LD
ZYie0hqHX9WvqDeap4XVEKkR5UnyLnCirffYkz7VWzX3r9mAd924evPk4mDJdj5C
W4ro5F//f2tlpw2R6dQE2cxElbMkytjpoO1XdhSVSFn4+v0f/qbZCUtUgorvwQ4b
SeFPPpTyVI52H0X/FnLXgdc47Uv67Zybj4mEa8hArtVgTdIb1sCzfF6Rf0Yx/hr3
0CdUCyQRKCY7KvYFFZs335reBUKIyc1JZEY2QDS+Vut4JeK8+xTteBKJjppGK4wk
OpMdRsXMoIz9B8AJL9T3fuSV2SEKK86CV6yUQC701GUlTGkdqp7QA/sDV0eCIENZ
wAcOEy30G9VfzYuVT3Q2wXZ57E9rJMIIl7vMdtpVKVUepfnnQ8I+i61qyXx9xZ6j
IDJV1W+NAsFwvcr3woI4BYwAzmyhxygnNtBP2vitvASGMOkiH4BZKd3QBKRIRVo8
IqhXG3/CtI3xqK2vs68cop4EC0Mzh5HAsQFgkwy+01zWL+XHI5oaU99xRG65sbBk
PsmOa3BCIdsj9AZHrbT5uZIG61p1/LisuWcvehpn1CuDuG5otf47x5ydPSy/lDu6
tdCF5bK4W4D/kAiH3x5Cec1zm2WwkZoatTra028XTehqJJEMIhVBiRUHKo6y/KRv
DmwbBGP+29Tl46BFRy9WPY4BbkHReE8wFa3g2BK8Hg/1ixClnk3k56qV9Vxoqy/0
Akc+ymhslEYz1f7cQneaLEPWWz3hx2ul9q7qUODQ4JSgOuoglqAQg9T1vpt+rzUY
WerKKmuRkyhA5r+O1ida0U/m+r4gRuWPN35mkUfOZ4JiCzgIzRzGbwe3kFRK3jXx
S/oE3jJ6AstSb62lyDtkCmha4Z7jBwHL50lFxmBfQHTYpgpej15KLiAkITkQfWdy
t1Go/jrUnntQ8v7vyLrLXIyyv6Fe9bneHsDHAXjluFu3j49gxcEQaN6Ogr/PVKcd
ieFraB7G/OGBhOAUB8fEjgmFm7AUqZEt+m7mg5zkH8w+eoBb0DqE9H29naZIUWlw
cqVK2mnIACUdEOBjz/gHwGIhGg9fvCpWO3cI/ci/tNgfU8XiRCZZm/FbXaQ1XAeF
/t7Jb5/MohmFW1yzsk6ZO94IvFvbphyObcv/ZSl2m2eopSGSMuj7Vgp09Avz/SDM
bt4SbVPiHqm+gPalbAWXA2Ew0OORzmhWpZMFwNd96a6GT+AIx6T+BzovciRHAmBO
3Z46mXrJDjlZ8oJ7lzbIUdQoWroE9kG7Dd4DD0rpyFWN5ZFtg3rYJNQtVuPVksvF
F58pvGpVUiN0NJK8aurN/BDLK3k8knjnJqj606km1T/oyOmgW/CDYDo0lv3fl6+9
y0CGwPhpJUQsddV99DLB2BGxfXvHuSQIl7oF5A9byBovL80BPkKgAy4ZIbLEK2C9
eY2SwMfetfdWaIGm5mCxAS77mSrfSaukMOcLA2cAZxxdzFlexx6UJptFcIt1m+YZ
SaBG0OCIhttVi+vFWzcRQpjvjBMdCVWHhi8rzXimN+8Wxf26k4ZhqEQhPqHIeTza
1nFEbAOjGbrfCr0A1XbJyjh4dlzCSXpRHNu+fCopez1F9a1+cJRPpHQXpZMTGk7h
X2/7FdKYGUAD9gDMg1OE7zQNoJTfvURW98qmd0vjUeovYZC5jZooETQHh2CnZ0aI
4qB9wEcPf80e9jd0V+1mkAQ3CLzj2PWONBAFcwzFfD0gmTksEkCXzljTeTpVnx2X
Mz62wfwe/2TSEnK0Y+mX6R5cUxBSu/PjimxgnOFy5FJaUJ4X/WFyuEArZtfs75fS
SBv5yvuM6Qwq8+EohSks0PgPKQNnas04D/IEqsEgwYrgIVqtA+GbDGzvqzslHGIg
1rWtWGCxDDPvHvzGSlwVS6V83tGal2JW36tsWlIkCz8fBFDrEXsz0l/fgN4gvFHV
rSI9FIjtIaIaGGsWimoA5q9LU3ZpF0tRfdTHa1PPV3EcTCew9exMXlh6GRUOdlPZ
a0ouJEi+AHtITEUWzUn/Tlb0lmVVAmdD0Gpo1h17awjgq7ITYoHgrW5WlCOqcZbY
kHBhGmWWkFWOZAQ9hYQcgltFCH+ZhnENJZzzB4NabvZdpmwL4I7RW5AE93nT4T8O
uUd0ijHGjit8+XMocIbc9auRiZs9fQUAYnYoqW6Zc7zQIP8KYKDOpBMpB+FE/6Ta
Umtr2ftjHPlhJVHObviuJPN/YrwG66QKgT7HksCYnL+5AonPfE9X33I5TlfufyRm
Qco765LvRDyq/H2FANI5jX7kACwoyDBoG2yBpzgFPjZeYHEXPULFPKN5Xg03BJTJ
TuzeJw6DyZEyHeCPHzhzmC1vWuiaY3GnQcYUoLl/JyKvmZpE/G79NOT2K0oUPgoO
VqkTgvomV3IQyPd1U1xXWkIAL6hFuI3Ab6qWFL9eNYs4p51kUB6tGRNByoiW1vAs
WVc5H3uil6APMhGuK29ZjZWdot6Op31UBLpdTYO43XkPExcApGM5ln3Rx5blSLma
9CS2ungfMvfX+HRzhChlNkBBohN/z7Ib85am2Bo+Ccji2Ci156TxrSiTbeTxwwmB
IQRbS0AvIUsUBg/vrvhFAE8vk15vR9fqTO6DYFoAjvQ9mAdgu1rkwTU+xNq5V2DY
Z57rOaFr2tajZj6fQXUWlu+q5TvrqH5mFAZY6gytwyQbOeKxb4/6U32hUZriUk1b
X3Yu04UFTcJOzuYR078+yWvPJs7bjAs5rVLGLNwTle+fqDEhiUH21Q5ToSv6MMar
jUpxGq/XG7u4NLgZwUiOBy4Mmp/sZcnoyUiPS6LPh3F0DKUhjNWMyYyrmK4CCyed
hbxFW11LG0qPu/VgyxTf7F622MtgYYTw2r5E2JlOUP7uHau4Vwfs7JjGK0u9XUuU
T2J/TbD4uW8wcxPulyOZG+2ldJPUzC7Y7etyScr/3yZlsZuyd7yvD9r3BTlTfUG0
3RIBBn0dvW7qTAHWHb/1v0jTj5WJlrRs8xQhpD3QNj7bo6BMuA+JiuZwYkhmpjcm
VDIvhUT8hnVbjRpBkN2Nj1+yv4XFRSKX2zs5uW3RY1isjKnN65iRQoM8y/4As08I
hF/5UKKfxedo8WQI/3RWD9P8Dfzt2MQZ5GIzpB8hnSoyNrkL/dYzw8XlvNkiua0+
KqLrGvAf3hSrY/oS7DynEC8NL0F1mwuWwxrIgN0hXOXjhJpJpTSbQ8vdl/f+Rt9r
96/JkRYdXnyVDfdT1uWnkDobrNchRG7Yyikf0qxwVlUeCCwBYds+2r2O6SYjatrj
AGw+OikXrAZo0EetYwR5sruH8SLA/sZcOtqQH8MLVBdUGaZUvTLj878uT1pOOnUx
Sh1ATm4mXpibzWtuwK0phHXDrnyo4jI5xay0YnL1U6XzQ1SpTGGq5Zvs6Zz55brG
IXi0w5lFPxB3HlIAg/uVP1cXHsTID2kYpd2qCqrFgZP/+k6rRU6F7HccYDSkcYvO
7qV21wzdmhL8i0AusVa4ix3sEss8OcYmScIkrMNHg+AVyd6kdAwotbTh4t/lfhQL
yowjusrKDf03Yf6coEVa01WPQblbiWHtjOAT6JaG4p/cxzEYsnCvV3cZt1PKI4SE
GooCkMRZlLwppmMdSpOVkHY+yAwHFLhRVlIe3Ux9Y+6bpe/ub9Aqs67jxWorcIDW
kvm68DLdv5LtB8Mtqlgj2oAB7YqA5ho54Rpsgk1bUYm8l3BxKvXzJ3+MBEH/cpD0
CD/mRygXQHiJjBKTBsyxmML9mMeMQjwxP4eLlm0kh2MFeDK+SGNST5MOZeDsmL+e
D6hJfh9R+0wnj06K6vHjymlt2NkGpK1wLHcxSbuJVfEK5eOfcLbwiWe+1MBSE4UB
AecUJLQ1XEmhk1s0zD6xXPkYWSx1SMpSY4WaLLM60P4wLoPw1kSZdV3dAoPRZAK1
8opljS3P0gGtacB9ikCcwLDNHRS6JVzrHkrpLt5HsChGue18YcH+a4nm0GbLOQec
SC0J/vYJAy1H/UVouwPtp5mgFrsCYh0G9CzBSKImqTomvEdbofAtlcoKTo2RGbEZ
yzI/MJLuVF7o7Iraof72158X1ud6zp58lFaJAnea1OwVdr0+QfuSGtS6gG7MFQ9X
BqC8FC8J/I7sEv43W+GjFDrdOmezRxekn4pcT6UtebfSsHBc5tjgl/ThqA+2dxUl
2TJ+INCx+on/wyiNai/8V5WnMV+Wsv576exIWdCM81aTWTGQHa/mYRFyEsX8nw5r
TP5GKIR7X6Oi6lSxfvMEZJMtEO2Fg6gx5s45Btp0C1tLJvM5xlMUbNqo7wHxUmMX
ckN+3kZwkkw7eCfhxLBB/ab3Mumg2aQkpZEJ7NLQgjXk1RWlUbg6ScLnCzeZAS+V
jY3j9Itcd+4nmLvJUhd8mlouHs3Lkfe3tPTjivNNN5oGy+bZJ7VZnxewu5np9Q3/
tuPBwLffqwjy7/ar+C4jpVZc+rA6GOlkWBgkHmo/KUUfcF3hohi3hHGu5vU3JFAj
xEZRdmmJt7xhq5Kt9qzz245xqLOV73xnjNS2rbVTjE3aw+DN8SOjtzQCUYspe9om
UB0yJs+CVy+Vg9oR/8267DnNfhWW6VuYvGftakWDeLP7XgRHPAJaZJYqy3PV4Ich
Tchj5+hvVoUsUolGDrDon2DL0YZvm+UFE//j1HHbhkm8CRirfvR1HtXF64RE5F0p
o5LIXEGclx0SmXV58xLxzyLUsBc+I8O5iscuiwCpiL0t7TGFJm0IzuwP5jyIDPez
EPmg+VGiWOY5ktPNGp9tnkGbS+X8E1PZhP/EXRv7EuIrx5HmwZSsnq7WEfgODPtj
/G++j0QR6/adqxV+DPby+beu0SkFTBWV4SduyMAdHcp/QWbDlkNwVjF6q8xe3AFp
wQ0n6eW6O55gBfyJfgAO2tdW5nrZpXvaDYTs0asaADdItCvsXNINseOuT5y17H8F
vT+GEaVTznWZ25kHK+sMi3fPQ6+S+sRqDbogUU9ZnAt1Qnz+b+7WCP9spAECmlPX
Kbb8B88SWeRs8okqT8kiyQS8DAg/LsgtLacQYNYwKZStfqFGy/sMBzLWsE62MtLA
7x4wjhuWcDXus0hjiO5LCQy5KRCz3k8wl4KiIQlFsnEWG81fjAHYDVQ/38IjjoSi
rn52/Fx1lAxtE5DXyFCT1JfRrTvg6Kd5vTj3bLfd5edWgRfFm0Hz8fy/IMTs9RvF
H+uE2LGOGueq7pGwUPrg+l/f5PRVH6v72DSkdsKKmImGFyIweMfAB09dxDvN84EW
bvAwsXbSUW6m81+4uTrAibi85yw4SZA7blqRm6meA/APuWje52wlHQYzNi1gom+z
qZyB5FXkzo/BZ1CZanpmPAR7yyc+fgBlNoMPau8g26Mb+BNLDn8O44XAgtee5O9n
Gn7Nf6iNEzOdZTSB4coFKYP5A/FpjM0XocP3nj3mfIBSGhq+vTJ+V7NXqP91OdmD
PYz1slBD+/F5pFmLe7MfWPt9CeYuagj55uf/h3+HlOriJKuou7TX0BeFZf8Ze+y3
0rpSBY5NcPscaN39fWGuwLhvKDNsULE5gEu5na8C1gErT6VKGrCvWAhfGTXKfl/e
Z7bQNtqgYc9aDPJXg834LZpnTzWQNWdcwG2HRHToO18slTknt+cdJv7MJqDe+kYd
l9v+FUQnBcycqB8DYKyj205mVtf58FW7PPKAcNhdOBTcCiZfmrkV2dZ9g2qM2/7k
PgzJzh+hgn3eDG1eanww6zxf9pvO25JD+dxdlAepMxdHjHG5YTki9tCgSQe8uQQb
9idyHnXxutl8/BH6zuaY6hVibG18yNG8K2mRwNgELuHiloXqnsf33pwmc2vh9bZo
ADvBiyVpYHzg4n7VgAxQZjXDCvrARVjOXf8orU8TEa1VQ3ONxnqWIM8UdOFhYxnP
rfZDlDkv4jGSTX8fDlGW3WxS/qOWY33jPgA+OUZ5rlPPWqDh40IitJ+XwKQE4PV4
fZP2zxvf7Y/UIgld+lGcSYRDrZagVril7i1AL2KEKkVZCmkCDy5gRlAae0fKYfBd
blqGzpdTCf7ZZuSUHXdODXG7mVEiXxSQNsRT2eAE0nqMFOfLmyK0s8Rx+dKD+kQr
qX6iRPH8Qs2ku8hBUPLugYw02hqI0o62wAhVzBOKPeL1UoeeHwlxu/WynAoVrAOS
yFjh93bt1rhO/2PL76ecRq3b3L3XuCp5fTh/iwahHoLL1jZ8s9e/4mnHb7/TImsg
WYtKDBvjtJmtSV9B45L9yVqzAn3tmAwrEAbZL/98IFSSv0ybBYjb2HYk1iLfe+ZV
sUzYx7U0uO2R9y/5yA9JINRUZqsvvSC9JAYYU4Id/PwW+6Q4IVV/6PBrWjj6Q/bn
zzLbuIe6yWSL+DmWMj01BdJw4wN8qSzFYLIElLNCxgnU28e6QE9IdTiZ669d/W8R
PlOIksbD7ghQmNrr4tk11rkDCgsaNJb14s+sIpsEFF8vaRozkRqYpN2QUZUmRGuY
4vfBufAjr+RBNGlSWc8NcBhxKas8jtGD22qezpnM9KYTvs62JMmg2zK35l4n5QY2
M4Axh8NFwA5H3dwAk5CCqxrmgsDK0Cq4qbygorGmX5H5Ob8VEzv57IuT5x/BX8C5
xT+zp5jyw4Ih8gTbBpnBaC/o2/+LVbNkSzajIQiXzGa0cu3DuHhsdTPX9cQG9QZn
N0peb6i4TsZgb1RkfEdQIam/9gsVW2SD0YvIEjyAWO2jGAipRziTn5eGl9JmpVPi
dy/nBEXDcFkGomA+FUMhvRI6WQS8Ruy8574kwRtYpAZhDlKgE1O+N8NDyPVt5845
xg6v6zsyiwNudJ3t1I7WeAxXbfrZw9jg8z0JelQDoXlUZBAuUCDrpZxOLKNIiyhA
Q8/Ei5Y23rPADohzmxXPaKwAcuydeRjRyYaqgoMwS3tgiugfvCntzJ+kU0troa4C
jh/pLayQY5kFHL/5EZVk7Yfx944nMqa6RmmlOSftmIodbTccGLh+7lJbaqLg3/jt
9sHLuglYJKoxyzsI+S+pdZt5h/BfSiemM/bwoBpoAbJE7SavOdqlFN5K2eo0qgDU
XV41/jp4SBmNDh2k1/LvwGGQ2bCOa02ihK8N6JwS4ndZsIsF/uHnylQlAmDVnefn
g6rshsZhvWDbh/OL0xmd6TSSLpBcTHjH4VkV+DZFBJ9usDLPYSxILpdAMpTtvL58
cuEpusl8oIsKr4eLubPp+lKoIxFh2ZbKUbuCH8qwP7WxeFQjhVrrtIqJLJ7ah5Hy
srhvWwdtO1nafNtpfsLYIEqrrhOJzsyi2W0zPDD8tTyj+Xsnr3ssmA4DwY8RF5HV
YUMXTOyithobdcOkslSbO2+HuiyqfiQtzwHS5q767OSZkxZZBEE1vdThRMgzbhER
U1t3SzFOs4CBc42H0wOzmvxrgxiNT8n3vWEynEph53ALHy0+PFckNkAegiU1/Tw6
u3FM2HDeZHIJKpVxXtx0Uw7OKbanentgOCOcvh1XoGoDdelilcrFrfJv+56dRVgd
2KDAMGtwzFqJI/iVy+8eaXU4VeOtbC4gG4YZaiGK7FNkEhZaPlID2TRUCJKRZZ32
M4QX23pXmMnSgZEVhDL9KnGHnf0jti+tzYZJt4hkzEj6IWhkzkqcv6dzRVJkr0Qe
b8J440+dRgWbZl1dL0+tHbbhJCRlTc60cNMaosKeUBpzJpCKdoRd2UzGHu1uwxUf
I+9z1Wdi84m8QudQj5RM4XUAyMnBdkFGEzNCHcuNXWd4Tg8yAj8UPSUfusU5n7yp
+TmH3LLUrNjZZtN1KpnoDit8cqKwoKduYQa7uzE+lCV+ZVe02wok69pBdymjGlkB
6XZ4Z4VBO0arVYWWFoN17QFl/bYeoeF9/Mv/UafdLllUd248WmGfWvMM7BFLfHku
PVj0aM5FbQ6sST2OLahQlns3/FCtAW1TQD/f5e7065s6bJS2AJwMcw2VY5mbpJA9
a9AZauiRkqhPH6giOZaRrKDePlYbfhrfhu+k7H+2frIi4ksXAUlgBG64YbkhU+/X
i2OOuMzPOPe/Za2dEGD97R8jUBd2p0phlSKSCIIT4SXCCTfvrq+13ZJdc9WOi5Qu
LhpzJbceZI4t4NTt2Bd8q916b93O5haMa7E7fOEk1ZG3QRNvsyrrlX/NNzfIXMvy
yIu8u0KYs+akDCasGiQec4KPBT0fmLF6LsfTw0P3h9KIU7MpNO1a5sSo3Pw6WrLe
Lu7WG/9lm7j4SdonC6AmLyfo+yGnTt+8ctPQu16Svrp+u6QkmQadb8AqeQTaa3F1
/9f2qTdl4lW6BjjhvZ4xq0vC2xmPtMPlEdQ311BQ1H3siIYx6i3YKe/PWUxuNN8c
SwwcBGsiRXSUs+zRH5Ur9kIYf6oogM9cINZ7WX6R1lEIkowYnG34hBIk8FQGMolD
Af7QkoqBhoGHMg9C0jqX9nIF5+UzWCh/Sd3uA/4QhvoFdBO63txHi19BE9hpafrQ
IWEZ0InmISqcEnw9ii5/zYxqtJVn0FtscRH7LuyH91+7aIL28TfatAAUTUowbXlK
I10mJ9i/fyQ/Q6PtFd+zOID/aPEtD1nNaVZ4zb5zNky7a4TXG994ntjb0KlWR/ju
G76vLkfj/IVFHl0tjN5RVxOHM0WOPHpObf98/wPjNttuQnxMoMBWwdz5miU0GB4w
Pb5lT5J/qPLr0QejFHxfhvi8uCDAQmpBwn9l6bpkwFMW8wcbhhztQoIpC6syywCj
V8/dmvlYLkcJyxdjUBq9C5X8QDvxuT1O4A46+81WcEz4vB3ANLn+ra/fFD3cqc22
Tsm4jQtTZKgMIGGYpMyT0nd0yEmGC9n0GwDvrLNWLhzey2ZHPoBvxdrklExNM4Xq
1PKW/FyB9dWh79Z2p+KWvX5HbZQ7iY8DXW3FRswXAgN8xx2+5q0FHpzX2VchDpGU
i4LUYe4cqIvLlztdOhWlURG3cenWLhtXAW9s9p4RFZCp4PzzMY6f194szp7OvAMh
BwtdKZJoZVn2og3CTJuPeZp43G71tnPbZa7wDkJnbL6Lr/PW4PBgeFZ/JDBtV63h
4adVnLSgArMm/K8bmqvq4iXWXCAJjdmxELe/+qlpgk6gItgCUkmCqhKnHMEtfWO9
W0yFaZ4zHX2vlZ2YgRZgVS9jghX4aqgVaXmBi3pHQfhor6z0871Nte3tuI3HvdFO
3KoqGyA+3Q1uw4dea/RBAbo75pXTArC+erEYmenv3g01o1NzdA9luECSXitpdlz1
ua5OZ2Uc+QCvWrM+1AL+AcmUXRA0S8O6R87ADQb+NkL3PwNQAtDvrCInRFJ1VLJO
KjmXoaGF38HQK1/jBwVCUzokxGD2j3JlwM/vWbgnKRyol/8T9lp2oxjcYFOZj093
i9p8tI43KroMUcDkOkirunImn8G2RLGRhgMgkK4MM/9G02fPzFKg8e4clnTAmLIk
pENaQiWLEDJmvV8DN/Um1hT0UUlCoTPERrFtdTqcMAmEQ5pP0lmtj0A9BGICA4rc
yDCboUTRaXoZnsPSnMScWqNxvMZ0mxFzG955ERJeeRPsXeWRqXica954k1X80nth
lHvHc69FPzEC/uTxIfmE+fDKWcRCiu+TzrAb86/M3ogAkc2wbRgrdQGB1OM51ZKl
KzlC330aXUrZpi9IGGn3KWA5DWul6R3QpL+as3J5qk0NugVCEUvlJHpsPsp0Fy/M
9/d7iV5M8BFAisfw/IDKgkKzg3jmW1cdCwozj0tXE/ikl9jxIQOlRDzSPuxZGIHt
hWTj+XyqfbZSGDjDImEJ3rCCBAhJCye6ZLBDn0bQmlHSUBQ5tnkZqvaVVeEyWDCk
EKegXtxa2JUz41C334yth/8bHoDagKvTr7lj3WcsEr0MwAtdbuF8ISvAcqJ6apm7
izBqudpoL/LkAxJIBBz2vh6bcHhwOVuETrq8xAbp6vKYcjgjeWlEmo71qvLzLzzs
rqnya2pEJhzRrujTtEezhZT5sn67zpT2DjQ/7u8ClEguNQWkSeeiIjpC4Wc3syJV
n7czkI49x79Y0k9Vn8bdAfsqz9wX9ZgyD5eE0zaICkmTqdklD7B4hf0mhmoNkIBP
cMZyShj/9mFXzZ8TqNHSn/UWuNXbzBWRMwiXdlnoRHmrV+1pYsyqiX4eoK/EPZiA
/pUo+rp+wEtM36UpCMze9WpPvIQkSrsbo1PYcTFmI4X/xFaFLREDAR1V0o0t0N9R
W45sWq/4h30EPRAJfDi489Yo1tFFhXV5lhlflIMACUDG7vhpTj5ykO8HWwrivpT7
Fx65PnDuC2TawAuY79zTkIRceCC+bWCUSxDv7WzsBUedO8+nFYWT18RS8nwVLekt
gL2QWMUdkRRq4chk25JCRORJdCE+qgtVYECowtzZF94F644B0mSAdxY20ixxv3OH
C3MJfd24Iy0g43b/TLq9Uc4ftF81Ip2Q5SWC1PxaHy5y2/MX5A62+em14tRHIe9z
3An1tnpkEgGBkTX+YX1+rvy0n3judu1nNGqlTo7iWdHPTJL1z6aXjYQtHVkggbj8
UGIHxxVh2NOBVXURtv/aKukBwF/f9txA8AJ4mb4Puy77gioTRqV8BmeHThhWkhNy
3r770WBRiWxOjDzDJKepHXsOaeypXT1nCz40bKRj814aSksGUtnFJrZze9/JDH9E
Y73pEekend8ybJPQc8NndGRMg+LSj99K1oynRwBHgG7aGwARWByjIS2Rse6fjVBT
tj1lNHCeGgw/CcEfR4FixEPUvOo7Ys+Zd8LkacZsnb/aLNr1EJKimmr3F1N5IBrK
KB2Ly682abwt9duTHJil6wUOnoGpUR+pBihtdpFbwvhg5JVCd2/FGV8LkErTlggx
bgbtwOOBBQSBgpWt38f8zp/lWJSxYtQ330cWyGTV2dDEZbnVYwHsNkKxusQ5m+le
ELulkIqVALwxtOyQIzvDgTG9gZbM6bK/GtIIefkPiKz22w9DJmoZycr54GIGRSNa
kT5zq6+VnW2GaiUK4/UcM49qGRtpol/iDmOjxX250nVEWN/XToU0pep1Si9lYRHr
W08J94bdW6IBIjpRJEd4YhT6DHFRltCH1wDmn9xN295FZmbESXZn/muBuphzx834
/pVCapvE66grLIFNJapAMwKj6SxRttEE6laEdzXEEgMx5VJAP/pxAcPBvmuJyPtY
PTZzUw6K810M01ESri0f2xWMoQumNiKSPGwNmmUZKWiCJ7PoEY4AECGFDCV9UK3A
g6bDB6qB0RvfWeJ8LZi3GlEItc+KoJi/8pokScjiyc2Vff77nc8YN7rOiph6/xs5
Z+c8p2WkbslMU0q3kYb0NmAk0jlWRHi/nG1t8iO8lZFoKrs9tm57WVhfaYCaAh9H
i67qPMTQ/9vngPD440em9CL9jw1tfpYNWpRYSOd5eLC4lwTYBN5vAS6L7i42WUb5
cNwtK6dhLoTmDP/a9OC7Vh+4hLZCwt6AnUr4VbwX5dInvzbktmP5pvZBL1tR82cF
bMg51vM2YnJK1grOZEpuGKCSXHKnoSwEIcDQdbHAZ97worNyccHJ/2E/awEqCnWy
+AR/hQgchnKPe4lZiMMiRil/hXNbrHrekYbPgR1ymKFBpvk00BxTbAzs1P8mN87/
mHLNg/Rw0MLHBgp+/eSb66vyGteIaewKbIfUtWGOVaT/tWiemTFYniPfeQZtSwUv
fHR3DtpERg8/q2j8D4g5Nognh9iMjuEDiDat3GWM4Akte0Dzoim61L0OOFidWDiP
4mDm0z1xIBtR6O8X6STU1Ylr9QwG+yn5QfyZajma6EDGx7I6ei1rORXcraG/EFUp
N7/7dwMe2uRTkiBtghyyQDFu7yte7Ws3gPmigqFHm/iauJp7cmOAhv7Z90E5a3Xz
RUEXDuj8pZ1vXbQQt8W+wG7f6y/iiNJrMCcUGzkdaz+2JqfxE3xpybfDtAcHXgsy
iRlvLgqCl90qL7hIUCvoEMRBd56mdtRI5y5J2B8kvFg+yerOtThcs5PUcLWRV2HJ
jQgWZi0t740UgG1PBahuHjw8l3IyB1WOQBn41VVyq+SRnL9RU8fIubBREbG1cL4a
M9mR8YsgMJD4ycWem6Hn/QIyc2ZYg8n+F/3wed6+lw55Olq5uDDMZvDLxcXc2TO9
o1NA3rSJfNwBWa80uDavISVP2FF5woQ9gyQK1ZOTQnF6ilhoPvgF/E6RR3eBwQT9
MzPb80AJfXcxA3t9iqC5yfZ77fj6HB+XvGq7m9ZvWMXPc3r1nMk3L8uJFQElkhKi
JocIKF2t7eFOgww+I/pN3LRxMKfOO4DngOFt1JvfgOD+VEWkRS9prPCMWk+RiDmK
u/UygHqm6WZGDVFwGhg7vSw+Idkq0BGA8OfXK47iw/r+B2C3Y5NmPZ579UFYtuRy
ZZdbbhs1I2m3N8XAAEVTN7V+spbZRoTHFgMs+/X5m5oh1fGng7svkXqBQ2FrOv5h
PudNGY/YwTTEIor5rt6fSc3FLkRnNfRlBBFJ1Gm6B/TF5xRt5jIsKjGcYFeRjdTi
daCa9F6pN5DVZPcl7m379Itr9lQ3/fQPPjN94XasPfJEFsZhs/MgOwg/8uMRCZ5U
y+Utds4WrdD4NaT+9cXwkIFjwHqYhV1B1w6dvQVZ1mvlvSLbMVqXkTieIdHRXG0M
u3sVCNRNiu+xDR2T57rf+4+iJPc4eiXWE8uVM/VnVab0T5ComjsXz5TZa48F+FLO
vVbNxdbt+yT2fYgEo3ZSr+Q9+XTid+RDjl3/pYCC8Sc2YWyXbKB+glloakNKGvLE
BqL9Bjeu5z6P7ZbWYJwKe1Tiv/5wxM/m7CO7no5Ho6gpXP1ca+D2UZHvZneIBcgG
tQfgGsjG90ZChBmKHwOVTdyjtnpTCTGzfeuSktnsLQVTO6zrmDELIGIRgnOvAK5j
xxizzikR0bRzlyTABg9f3pd0WrGC9h9jGVOZW893XleqDsHE1D/VbpklbkKDtkTB
arAJl1HjZbQx23BjUnl7IT4cjvZpUbyt7zkd1I8CvudgfBJZTE2CCs0wkgM5ns+B
Ma/bMAf+iHZu4jLiP9vQssJ8V6gHV/nCE0nWmQHNjhGhZk75sxS80th99GifN2vE
Y/aroGxsCv58+M+yCw50gAzq3ywMsv3C4T4hkVDI4zjeJLjgSmsV678SmMTTdWfq
yH6eqZkfPCm34agkbqYcdaYiYrQn3I4DsQ6yUz/t2w5kv2f3e4zvV9owusUXFu43
Xi5PEUuIlMhC/RDknLOpLDWm5N8FYEvFGnr+MqTPpOB7Gz17DuJe/MmAav0xm/hw
i2GyZoZdXUACL/OBa1SDaEE2IOSxejFYMmwh9zhyvldj75oPGKsFLEzY0gyEmSOv
lEkudJo13CArOGgn+8q8GQSZBRHQMvZdFjyEWpFqrwuGl0U6/DpkN5B7IZ5MpLmC
UALLPKYLSa7WQEBLVMvBh3H21vDwFM22BBnMtoRZL2e+o5cEZ7fz+TDlpsnxcEAT
+Ii4XFw/M2QCDyY26quRSOOYJ1PDxi2RquIgh+hSzjB4/BM1BWwRxDpZmFHXRozQ
v+iwYH9cGct5BmCq78vq3PGC05dTpmztORRJjO2JY4OhZ7PYrq3SEg7qsV7jjqGI
Ks/v8DoC+IhFTD56/0AMnsuwOgISyGJenu9ourESRbvq3bA57vnhP3a9puUz0uS8
tPjj26PvsUF7cXKzi4O6Y8VvNUDCD8PFD/RisytsK0qPCxVxXQce3OzH678A/WdR
ffYFbYWHrl/Hgp6Fp2bJ8/pX5rxru09vReCmvc3pySr/GaPGf9/fOp6c82ewdt+S
hCBWJpiU48Ldfec7yLVdhvU6DDCjEjtEAguQG+FK8XpSX+QnkhJebH+rHAKC8SOI
G2ZftG4pGRe+xHAcyrjA0R2itxjbLSINzudTfHvmXgQu2zWxjYcVKPmO9wWvJrD/
rshT1V/va0gLCUbXGE0gwayahEWQI2SilXPtPV+HZ33ozBDGOKw2z9WLwpRr+xNW
dR8YgYKmFsM++8RiLZXtw40u4uoU82woOarM7VRK9jA8E36D1QI4T4dT1NJruIgl
ireOEnRxuPLm4+66tXdL0wEYHfI7oSWOCUJ4wbn8LADIS7g/2cLS3DzTovbEDFWb
IIKCOvt6C/3vANa7ysHO4LetWpuUl2tip8xBU0RKghUdCbqU9QPIhSuFh0VmT0Da
1a+5ZpnhWl9IS3EZfoolEtx0iFfL1gXeu5+KDmyNoHWuRpvyKAz2q0PhF2pYtrfG
kqvVfBWKoeItqsH4oWVrQ2Bxxf6suXsnW+BtcGX9ZwCSejFvii/UTRyn4U9t4FoC
KZLjd4JOkhwYQnPWHY7muB+JEJexCj34TEzFv95H82ZnX4wMz4ZrEOof9UBmcJeA
+RjDFdOOXJ+IBKG0djGdxOgs/g2i7LR+aZDJEBT7BPHXdFU3lRcf4Oz4hxSqDXQu
YYiedMnAOUZAnu2m+hCYb/iRrj1litaHVQDczLSADNz8komo15FzGthXLjaPWlSU
wYaUuOOsWpKvyrEq0C6i2qma64DKHdO/Or3Y8vzsM2MH5CNMWzZABUl4l0Ts6Won
YEdstjIlDy0Ff6ydBQlSKPbSW6dr1YBAjcwkwxEPSHOX8g/S18fUsd1JKfDS8ZpI
TEb+Nu1Im8RM+3TQwAMDBLLsXeYciW7Bu9J6tsArudjxILgHKmwfxzNG2a2hjErQ
T9Zkm33cCfD4ipPqFp/u7fx9our4glqV+PEV8OqQIYaQo4+F43PMAsHQyAwkSWR6
JNyi14ecih8vWVmxrd2nhO3vgB9HkFaNhDyNbc1tyj0vteSmpzLwbuoSI+xqSXlB
FMSLs//5pfsp92UEtSylHwPCQ/PgMHNkTYvc4Dl552mP0AZlfuzc9Hy4T2ptz+wr
2LBCtVxR0nuuPmrBpwX0JCkQ0P5tAoZlwxg4JsRO7S66QYNrHTjjZ4pRWJn2d9SP
7whNas9mKLAoqeaIerHTU7LSndeFfzXyBZ2dmORGwF5Py4aQJs+Ra0hNPB95Frel
DqitVkI4G6mLycmzW85ll7mWZZaagcW7slyK/m0zXTcttyMp4CAEEdmMnwsW/r0m
F7VlncVczijM49gpSppUtBvrGyI6nYqpagOvOvztljA+QC3j8O8WZxv0BwCIvHg0
zWewGwSIGUqgDtUQfOLgH0YNuzAN0KRCFpn8vDl4YCkNA0aRI6Z8/HkiXWiwDNkT
gHdtTbmMMzwjR6JlDTH28lO0hcCHzLtNEciJaKh4PJ97BztZN6eXA9qSR5KqSX53
Q9YMBnTv8dNAQAFLfJ9ganT7fNBjbLip6VR9rWviVV3IF2dbVs9HwTq/RDv3L7FR
wXjJXAXefp5moOx/+MndYTmyCIkCVGFffb8JFBu/GIiuoYV2MKFIL9VKBJKnzF8e
ZooeXRoNl915topYna6Wms+fZbkLt6zmeIKTfNcAx36NrWNoaELv3yYWyWbqEFiY
65ZmIlZC9aGxXNm07+IzbxmPi5nUTVlS5yG1dLtx8beFfmgFO/RXqPxGgPvzR7qv
BgtpLppbdx4t66pT+DnO8kzmQwAUXtLhOX84NdM09d6BneshKc/+Suh4wvpew10t
HPOLZfKzghnVYFJeSYqgtvAtfWZ5qb1RHlazQj2Uh7W69nSQsSNvohX9iTO/NWca
midwjHsqUms5h9uUuBM5b+b2S+1BT8Xvh3e25xj6XQXH/iiXHnHpX3w6SXcKL4Cc
GXvXj6gA5oPheWeVrYLdHB0a9MO3ovJJkwlDSN80RTixUVRYG34iLMF2Hivxx6o5
XFPoHJNkeGe0BXoKnmZERD0lxORpq6Td8BPlemfxOODKuAaaTNPgG7roHpYS6LRt
iAwhAMxouNukuLJS6UqWiYic6hQmBiGaF+JkDUCHZl0Swpy2R5IGna+R1MLry6/v
SHHf/E/5mHf09wlKJbjH7uz+yrLjVuK6CqoY4099kyoz5Xlju5Akeio9NXXTCL1Q
cx1j7BC9IjnjrAJJkVL08xlDwe88J3N1fEIgrljWnVHZ3O1TkNOcjHNncL1aEf5b
imRDG7yIwLyBYOMHAtC0VCHbQsw/zodHLkNWQfKuAGZuEsL6gGBEHJ/TOs5ccUc/
l/fTwJOY480FP9ruFerCTiz1PDhf3RWMERbYIcyOYqund64oaPwaPY9UJ/xsAaa0
28Qp82OBX4hk9poEhZW8Wj+hYupCt7hZZSSGaXboCMUxsO0qlwUaKvs9JDTRBJ6O
F/pZ8x7bHdPlbfGRch/DlCuwsEU5g46vAzas2vqJ+9chCNjdbTsDEkvhwYCtbGGp
HLfEJTb6m13+QuZbZRkhLR+wDb8lYcNGQPIdox4oTd1c2RIzJv79WfHT1KRH7Gb+
/DBGVe8WgHtimunmuFuMDwxnKKGi80Nse7AqVOKOsknnWG4y3WLYrxgd69A4xt/C
f4iKCAOi3eWEGmTwOgt9O6PUfPmpxUBHAtulwBdN0d0RGoqoSHQh0opZRjL8y++y
A7l/grdn4bZ8GMuimU33TiKe2CaJGSIzDO4YdS7yoXuuxkXlarZNUuZ9Lt8SEZYl
6nFVZel0Clk7GDfRF4yNSxu9FotDpjQo5BxpPItJfwtHNX+hyCYYCQtkEHMW13/i
WbkKM6ubWMslS/E01c6lXa/xwvuse9bcTslg9xwSs7OjfKk+Asc2Aahr2mIHTHQB
yie9R/uB5wDvFaDZwZDLgPqcPk68UacvLpmBNejY7EGkcaAg3G9I9wZTm71lW1SM
Weat7TqmVV3b4Jr8uSsgC2b9xMMS56hEh4QvW3liZUWicXtMjLFAfqJUNau+MAtF
4v/tjXwI3rKeeF/nn9SYtJT0WAOveH9zUmkb1fxE7QsfOq31JJDFXJY6+FQ04zdU
c4clalTiRSEct/Dye1aK9R8PTfeTuC1YTlpsN5oHm6wHl9e7pCeoMHY3B3APw2t1
OcN4HNmd0e6Z8+cLWCMYTcOvYpy3xXhYWC2Kc7Z25OZsVusPr43EiS8kmlxWl0Hp
C5KNUSUyOMiAzP/TsokneGTB9T55SLWhnrbB/fGw2QFitvfWffOwYvMxs7Da44Iu
iFbO28PBbU2P06RVDRa3zrsmLV+TbRlsaeiU3ZC4dXVgy3KqGWWxDQomOyY0EJrV
lqtxTvhleK9Lu890w94Gn7Bbu6Ruo8HmEQn4XONjZAT5r7OPpA+RPkr6b5dX6NcX
USQvY7k34Z+s/gyq//L7SA0hXYlaRMYy/FjaPx5sfd5PKAnAnP8TtQaOH9/bEkV8
KD0B4ZfWU8W/tboaHjvFMWya7WHVPeah1cKLd1iqAqIlwTjSis4Dmd01VccsYcMy
L7IX97DKe2K1LMcoANXRkRst7CLLYh9EknuGK4pu7MTigHVc5hcAGygB0JsGkHOb
1KoRsfcoMCj7/zO6ozG78XtSH+lmnojsRMnQ1b854T2ctY0yreSPqeqT/ZtFWKnV
3w6dVrayqdplOzT3+6ic9zY1S/IqwIAc+Szx+8v8M/4ZihhQPZ/DZE+Ga42HRPa+
Lc0i6yDGL2HPJHeed9lF5Vn9MwqCFEzKqiEkCAFze5MhzA66khSmgA2xPrPcunVP
DXmDfANeXifhYJJ4mH+sqKPacpiEElQdonYd7hnj4DyzfezAUeBDCNS4nI6GJio6
ekel825zrEaXa0YhmUotaNt6p+MkM1mHa1RdU9yzX9+Jj/wWylpV2Yg3Mh/vY3rY
/bl0utRe/k1RovuxD8HkfGaltSTzn5jRKc+eWcH0ePGA6xgBTeqF4xpf8Dk5vve4
1xTUqGULn8tUgVzQN/BX+8RQSHsiJkziYc/9kwQ1svaIweUPoqDgYHA2p5kdshKp
QBD2tbrS+oTGkkAkDwmmbZSQSk2XxqIz7E64tDZcvbuwHLEdiDX+POe/OdGRLx2y
07XeAJNjEtbB29uUTzYylaawfhmW6c5eKz4beP4JT+geoooc7gVJhv6BdhzCpPfd
KnI+Ez9FzSX+ZwXmDVjIBkHheoSKa6bNMHXELlfx8M1q4HQYsueNOhuKpewuyIUK
U9l2hareQg3mRDdsWCzJSbg4taImX8nbYvFjyRNreMB7Vxfz8Slr7CtIwwmGJzTg
nTSnG8/HYrrtgfS0ncDRnAX158QB9Irj9pKPo2Eq7La9yeWAtI1Haz4x4U8r4t5C
ZyZ1JbCdVykhD2HeawhT2PBXSVhOm/FXt9gl+Glg2Tnz/qY5JvBeN/P5dFSJttjq
+OUIL1nxZMDrVUFlQbmt33KyPBSMY4iUuNnsnB49b0fyBX9U6fvgejsjCUDEp5Vu
jrshDoKjylXTXUVFFR/03Ek6qk+TPAg3ZTm2jdSJMsuMj592Bv84HbHeZfMWS3K7
bCyYJLgDbO4itT/bvVhPaMKb3xJBcEDJyJxNb62c2ssx7Bdp7atnu54B6RmXio7L
Z5lKKZCiMAipJBtagS7fcSf4P6g7VaftzEzX0pjyNbDqJ2khOX6nSgis5ndgF5uS
5Oc7hktab/Uw11KXl3rHrwrgPNdiakRFxSADlsgUEk0AEKrSFr96LoQgX4haTf51
0CNWAMAFY5llWYJo/1oCSQwb5GN8fXH7aakY0xBboV79RRRsl584zYqQFUIoU3yB
NpqUDI0ohl/tq/ry/Xbz9nL/IwmRsmuiqYM5R5F0g9ScjnqQbSg1e0+A72eAJH2b
PigSDIIQDyxzvU51gDFYS45vNK4vp0TZWt7BussINKPL3XaDwxn+RLLIqHVo1kHF
yjk914Bou0EhtSeifMkTiJiqAJsr8IPf0JmaRMgkFYrUhRlav+vGO+5BTbfphrdX
fC8dr8wy7/whRcSOVlMD3PaSqy+AHN2WCTVUK02Lt3J3uvjvKAOV9802hDOYTReN
olRPq4TJMu1tUGRa5tVZG7+3+9I04WsTICmGWpXzP717ND1j6ABdb2AVeorxnOso
BSEoFUChppu7+NYFZrVlmoqM9TD4XFWDkAv9k5MBUwD/iCsfOw3KTA8HINvq/IIM
ePAWEXKolKacKemu5/BAl5i3Sz4eUArUOm/vxhBlfM9QzZ9cYkjLTvV0p2FcG/GZ
BdQ1VjlGuiUbwXrEvARrM9wMV2vQ/L7+dugd54+KSxZefjdyMTxZvEfEXXLUjPc4
uiNXmaNcAVSWtUM5KousjNcSfFE/VVS17JWWV0jl56rSHN5y1VAMiRot/VNLtEf5
NpXcjm18JBjyEFaoApVlymEZgL7BhNcmYsbdnSnunjREAsR2DdltQHIEaj3X/rkY
WqYllve/Qar/dSZYbU9VzZTPgdXo9b6Le7+ZcOOMfRJ6KplxgGay8f2q/k8ng7Sa
Kb+ajifrnyQcHpSrnxMCaPj/YPfiN33CvanIHQy1OD926j8hn7m/QW2J8AaRT0Ae
kwQgGDQzzXHGMKnphIETh+WkL12CWkmsWy67+ZWhI+gvv/QsFNBSAuy8PPpTQ/nF
VaJXJbS1UDt4iEfQGV6RWCPchKblxcCpsbUv2mPs3+LGtuQc/VIx+76pBEE/ecVd
wHqY8ZAG/umgs7K+4TVlktqf0euG2qUNoUtVu+mb7JrMltxQE2D2VoCfgLEbSKbD
OCKNQQ9ZGO5vclIw3csGkCWU3juVSre9Q265iGmUuEh0zXgfWH4OA3AqnWLlijbr
lADA6EAoqWzj/HQIJk72L9usehFSv4ATJi6lKtH7FHfEIvNcd2RlvyfCsw91AZnD
7XLC/UshwKdzPAAt5ZIaafb3fkAxSiKUR3da8OPMbQ3fM4zE+zvzS+LTQoAyvThy
t2MAcAndudWRlsxza/vL4osYWVKCVtWMvt13x6U4jYkVqUA+rDEePyBWTZhlhkX4
/8TDfd1qB/yr36tTSmPMrlNf7QaiL3q1sI5aN243bfRL3zbhOcLrNNStxig5R2p/
/gFfP8DX90jnR8WIHp/0VSMFKWlmdjTVTdfMhiark1mQMhmVqApov6FI2GY8Ft8C
T5X6D0FIlr2wb8VuFteJ0ZUjYepr0lvswWRozaip2kLRBcwtLzO7HBwH7b58JHBR
hwZi5KP5CDHGwFSrEu4JdgmkE/qFqxVw5vsjD6KSMFm2YS9KMnemLMO51X8X74i7
KvMQ8X0QImuLuDggGdrXfbFDOl73e5De9jzTzXxbnz6AseNGLmO5vz+hcf46hE+m
lh7I7HKTGxK/Va5Dsdi30p8s3mr9tMaIApohiCecQ7l7UZAOq8Rtw+OTq978EDaC
EY28OnclFd3VWJYOlvWqzuyHcDm6yCw8yAEiULQjdlSciYIVwegzKTm3qrbtzAaT
kdpOU5rTumwGCS1GoTMSYjvSBiWsoayTyTp/wuhQ6QF8esXJaefW0LFol+A2ZLOm
U+oKH/ln7aZH0+yWg3IxfDlw/WRLvtUwf2u07YVXg6Bcqj2Iwl7xJAZf4PRYzIqu
JooGOXhxG33IoD17lz5PhYQ/GIFYiljmk8ekqtzsn+66FD+ZQ9gUucrgvlybWAgg
LNF/0hcD1+XcPiAx8dDIF1ik9cRg3J/hb6vQDSs69x8XYv+K3MbAIOEJwm+SEdau
mN3ZVMW1b7xoJ4wfifaPL321KDHxQE3v8iYaEXBYB0mBiejjHBwsKgZeYTyC5Wow
Tz/5Sn5wFA6j8hbqf55DfszWoEHONLFW+tVaQKADtcYMPMteD86YPIWeIPQqM0ZW
Wbef85WufYiPgVL6ZUhNwdXMMnlNXyhelV04diHpDWGpPGfUcCBZRSMpOX0/UZNF
CvGJW6vHsEUTVUZ/samVCx9kXBdeMG5sKapVBB0iWYSA/99ESQiDJz0j/SSgiC76
ttgAgOKnOJ0+wDNF+IUpu8K9/cvVBS7qdJ3dnOzWHUdL0KpuGScMjKVqgL9N2mlf
bLOiKmqc0s4gMIxTgXD4HJMDH1AjMbD2VCTKNpZKroggtGEtGzyHULb7c7NHleUy
Ai+SghoijCaaTYP4z3Wum5eTfCCwVyPWTBdydjKeoLrPgLkE7dsS6hjuXaSVL0fH
Ndtg6OQPalIFDDBP1qmz1r2qv+r9/8mILNY5uqqwLZfmIFNSSNEtm6/jNIj0Tn3L
hf1s4O6ohfgMbyZBFRuEY/a2P2pZl4cXrgiRsHD5FXVR3f4Sk1dOTZrhV97YbYh+
3+KYw7TXAww4KjXEHAHWfmMcOUXcRiC8Oi9YDA+1/HLaXa4VegAPSkemivEWNR/v
Jk+RD1XMcyK/2KK6ue4NYrOA8PnfS9TPLP0K7MAU9fV+SkmW/HTqnjeScH9O93tL
Ck639m18LMyIrRBUWLpa2ScvssiOFZYgAM3xum6vhiLAac+l6IBkT0+SdtKZ3rZ4
pGLS1aP111+crYoB3HHP2sa6VR8EI0IZDWDSGZZ3VAWjpw5upvRyWvFoHmd0dRFu
I3hbpPsxTE6s+j18R+av/EqmUVNQTXiwDOoSpDoH0eCWr2rTwthe6qpWRjAUf8a6
MpvyUaFPBoqOkMYBAdEgKfvTq9nAjj72I9ZJcgGoZpJpGuqdYJP6K24eIkQGN+VX
HbGcMH7JTPe+Ilwg6R7nvD6H94YQH8H1vt1liKy3F0Y4OeEAz2f7j1lfXC5fUop3
ieNX/cZTpt8Jga+7J0m78OrArKdk9EPiY8bPW60DmYLV96Ez2ENLQdceJwbAFcP+
GGd+pdx55HPIQYBkVIXp5ZtZ5OzUSp0Y/Ytgj1RHAYkxqgx/1B7IE+fO7lMFc3/e
0Hs8l+gz8HjccO+nu6W9PfWOs0itg9W2qf2Wuj8mpKDx8vgok1WslO6Dj014ttpZ
9PCQKYWpssdI2hP+aCFnr+PvG0EinwrVSuSTNWWHn42YsxZFYKCtSFs5CJSWYOBn
znBnw+UEJrBcSOQcOKqUCrQr6R8VpLPUXBsxa6lhBy0mfBZTmhunpw10r9TS2mfs
nTdtocxNmyv7wZ8MESTJqgLxswo6EN/Ib1mKULx64/SjkNkfUH1w53K7SWgB0uj6
ldU0F9ZYh/WnJg6k/hIGuhCdpBywikT5e/b0VFYbv6vnryOS0O7HlVawNmb7OvQr
SwvtSxWLMQfNx4klG4GRzOCWe/pUNVkgEq+D452ck2f/JPmQzZRwXq31/3/GJoY+
SFDVE+Bp+T+23a+Hk4yQDDSzt/2fjS89YgKtG9T1IETTpwgJUjNiITbciicC9WsW
vKthCxPp2jSUd5Y2FxtZ/JqIeisZv2U7FWirYdik3Tbv1UoQBavZKEkmLFdJ76SJ
VLHaOTbBoxO6f2STe9PCRTksBB7IbCZWzMw9qGF/8sbDTpfii+VkAenuXGf1SRc+
fdIqI2h9bbDJcJQlxfC6WQ8TQlFKcxIYSIn+OfY+a8mIdR7kWmVd+9am/eVm6Ftq
VNMT+Zctq8coCmsw9TnlRp8pko4iJYZljU1ia5zZaeghvxgSQsEdi3+OfSfTsdI3
XJ+vUUNumIN392N4/EU2PVbYYyL88wJdATlj0sps8zj4s/vNRQj/CW5rKSOyfhqS
GN/kkQ9dF1qoY6mE1+FnaTTs6WucUIXtHQN6IYlGs26tFVdzlJVN5Y02cxfMoFCr
7SIxDIz97SPs4yN7SWjnbvHf0JKex9DZqyGRHiQS5kDMe5vwx0aoXrHx4xRgVH5h
jo6zLmoETtAz6X6OGSB+fCNQJoJCOGfoniNRb/WDue1g9UEyJia42wJJL8ucTNEx
ySDKZ/QFDLR1IufmuCx+1fJkRpJ2DWihWh0ki5yglydWrrXRzIzZuZjHL+gRsjAj
hjR6ur6AkgWRdl9f6NasknNuwdCRmnzHriLK1wQ34Q5vbl0j2c9bI0ShR6C11mCs
c6H65oC6m8BR+Lf4qJmsoXg2Nd4oDHr/xWex0+8aR6o+5dGzvkfjMpdeyQZ07XlC
2Sxy2DTk4U8j+7JbsSy0LbxaXeCmoG6FG1UUSAG5w8+jCyQ/IaXo1P6jH3rkQBwl
xxSMIRONwq9IehP902K7J6Cfkj3NCmvIxQV0v1iK/YegSidwqJml7JYe7NByFpfN
ru7BXRZDu4B/pn+EQtH0xuMHOwCW+o7iWbLDamaHRAePH7VnPGPLjACmX/VeUaND
CLp5oqMFmH97B3BJEtIc8JQGQfbsaLfxXqbEx9Z+GWjBxOaluQMbt3aVekwEKcbW
4GztKSfF7Ry3Ev0yfca79QozREkujFaVsfM4r2J6VmaJg9Uz4QARygWaa8Z0dH7c
qNb1FRVKHbufWnpVPIGIvDe2omZAI8PGK37MJF2sKM84kEemrPDvowPu10RIL+dy
k/IGoqoLsFQyhmKE9zYhx7q56km8KiJu8ke0+9G4ET5fReoI26B/AYW5ss5AxvYP
9AbgVRxTEglGynautHzPZOnhlQ36RL+a67qEqcMRyAeLvv6mUePJLFQS8b5L1L7A
PpiIQbOv0DlsXAZbOvCzQt6Xdbhzj+d0jT/cdG1Rtef3glFY6ZcHxpkQ4QqFNVrH
bTaS353ARMC4cHiHVB/bUQty0t1eIlUQ2tHHMEA6pU0AR7crANTqsJlv8IsXipE8
u3+J7iMg4sNxoKp1YgIkf+L6vUXpb9AMhLEFywmc3/q6MRf5BXsj4iXIe4Satx2f
zoUO6rmoV8u2lb/2os8GBuz8E+NGAo1c/UNGjh9e8cuBPJ0yiE9rxKv5ExWEQfyt
YJ1HFB8oW10c51qr7cUYKhbSEEBVjqW4kHM0TcoJn55UyuzoHnb2/5MrWzTLsm08
6uPXeKTvPxDfrUA2pEGakaDTCqgjP95Ihocv2bVAvzRlIvts2li0bL8duhyDx9CF
T0kPC+ilOUw8MlC77SdVE+pXkzazv93hXFtHZKxTP0S37osn4TG+z3QBqmF5Z73o
osNiBI4N67ixKW/34pHYzHuS/8tURGVp6qYppyBmN8gaZXavBRW2hjiSDORmQguK
s7cQ8vc9eo6oHlSQDdRMLeBly1eX7wq2qVR6UBh0MYiEi9UCoElNG38KgXCnuZVp
vrX0Cy16TT3XVXhrfSXXFiPFe4ZuFJh1ag8hJUTGIgYyX8QsCeUZwRjBbcjXC1i5
fBwXrBGFRZGlf0XuQgc4T4y8YK3ukFSf63AqaseQZ0EfypZydBw9jabeeB11+3fx
t7yGKHoT4kwZ2jnkPtvf323dE88qFsawWBswgmPLHBlBX31YI5jyQXd6oQc1rzcY
Wel6USSoNJD4ai2VoAsmi2DwvpnCDy0DcPTOvzSsnHYA65W5zJW8aHpqT6U70PMr
KVJO7LUfiSsyuo8iJRP3X6m9mdBh8yoSUejobaJQdoctDq6GPW/2s1cySH5fwgdZ
3ZSWfIprLEXhIEfje3662eDgcrmBOH+/88nqDbnQvuYwYzn5rjcfWy2CGcpXPA1A
J7S1u++b/138kKQzizFt42MuSqBnaZ90MhPHIiccJO+TfwMTqdHO6pGlRwj8xP92
afdwTRUUJbwHzy8t36zrGBtLQOQTIYmFkAmw2W4g5AwMsVGbwbsQHYMBV66VIjg7
+fmLzLmSY4fy4t/TtMSPLHBnr8FmwmJkZwxvsPmFrZShTiLcwdBfb2r7e3sp/Lel
MWFr1sZMXYDAeQjoP/jidm351XLLZlKN8iJ6t5YL2fJae878AkncYdpis34LWyWr
cVC7siWKh266pwKNNQYuiVA0VF9gF38I4BDt/ii6pVBdTpHt6yXLZmEGhkAz9WS1
dq6yOqMprUGqts/fj8LB2bX5hCnrAqfwmMeb1TAxG3YxrRCKdXbgeM5KwJ1NmHKy
I7MKkWU30ngM3YU7LleWfo2wesGhmI0Mz3u3mi1o8zY5+sOk4luvBXXlpgEVMFX6
F5oq4Dlk7CA/7lDb3G60hoOX2F/yXXr6Uv8JUiadcuXEb7tWHG6jC3TrM8ozCNk4
u3GH6ol0CF73zmJ3/vHQgLol9MLYPJpUyJQVEFR983OVIizWYBaGEw6v73gD9mBi
vm4KDZuU3FUAcd7vLEjEW5BmLoJnnpEGoTkFa/teV8gkpR5OZ/fDq0Ul8fN4FqGW
sa/81L2xMkU5uvM1EdhsF3t/UUqGFDsWwGXecYafwZLGldvFKgUKegxsL/o+EsR9
vMOS6rl4vFLOBChMvAtekGyihjfCIDPC09uKKhablf+vPNBuDjhlA4JU6tIo9aIs
cV65l2RtgP/NXs5wTVP2/Nzq2bHElbcSTyvRJkCnNuyLUp6eWWB1n+i82pL7cHuP
QqcnkHrocvIHumslHnwZkVnHKh3WE9RZRTZ9AxMUA0ql7+jTAJZVNr2ld6WdAglG
XQcgZBsFu0dly2LmARz5Xjz76mYt71dl7S39hY6EyrTsaWhmKT0PymA5eGi9cUYS
a6GYPrfoIraBf+6LnZ15Nq/cMvi/oD3e12jTsrtpaMyPwLpDaXUEK7ZAKTsHKhrp
cDP0xzNK0YAultCU30xd071Tx/ZOcRt3u8c9zpSr8L0540Ut4w5waaaNz4duPfZ8
1ZYxJGUIRtakhwRTydL6qvGmxUwcHGiD6QII4YMqhkBXCjSnMquxp+BymV1jxNHu
YqwYXGs0YHfDfZdptx1pNWKznGV9I0zWva1eGrX8MupDmj4BseG8pKRRuCv4Mibh
PADYNO9h6eqG96I4s4ldV22lZTxFXxhZzP0NQpPWnnYVEPA2wqfPp0UfWQ8e8IQc
/ownZzUIznarRF/xDIpNfvL3f89QVP5q445+YCIu/ycLzDijPxVvbR6uMvIX1c3y
BkFMBLfZCpXZ4T91QXuCazEJzPlX5KX/LTyR35giRv0A6+nhEKMGaAAfS4xJUAnU
yDFxEyzK0+mo9LbJZGyorToQ+IUrP8jNAJRVjTbKVeNH0ELUZx3dGNDMm7gknNZh
z+UZQiU1wTWp1bKt62Tm77jNnrmPfM4HNea1dKbbC1MqTsbVg/NundssAZ32Fs6l
g1R9k7FHoj8P7r1zrnS2pBvNaSgZ+7W0Sio6sLwY9es26krF4ccdXNqtn5/oPbXP
0qN8IayBXQ9/iUNdq4R9yBcjAug1MnRmlwxHExaluKwhSIdMuzvYyPXhRIQMP2EK
8JIUTEPHQXkyn0+mcHM7tj9jZvDeSl2cduzqZm0ZsgsaqnmDc2cF6eiQsTdJ53Dh
5393DgWwvyXJLziabdkCUMF7xFeiuZZtGpIfZRWFW0U26+7wsTltHDb4Ry97ZNRf
1DzfNteQDUVLgbsIYs58xecj+IGnW4v/N/c0fo+WKNyPFmimaQ3YRLRTfqaI7TdN
6S/aia4GuMiQ99pWGecfrfT5PX/lkI4+g/yWzRN20EP9iYx4KeM6r3g4CaRVk9mW
Md27ukjWkGaUU8Xxj1X9V6Q5jqK3jzxqA/sHxITeLjUCEnP3mxLYmzeODiDgIxzt
0hQAIwp/wc4gAfqsQB9kVZOTi2+sG6nUJ8PjZiwUDGKG56AjrSvZSsG7sZUOaZVb
1mxK7xPaE5DJjPlN4pOXdczTVKTpaNcOgn7FFPmcd3l4I6WSg4G7Qw1iOJcT40yg
jXoSuepNGvXjvke0m+aMLUeHDxzI2vbXcnwqNXrMMZA6eq+HCumofAlj1Rj6nvxH
pjESg45BhqiMFn8Juaoi+51/qEfb6Ysn+T9Usp0aic7cc2bc2Oc8T43caLaHcTXR
MCF/l17oHr+H7AMzCUfT5KD35PtVRsDpKwY+8zp/Sc7bYo0wVIAtp7BMWc4/6PRE
5Z48w0CLLBRoF6bsDTo0pTp58eO2y0KDFS/SqHkXxECupG/Cau649HKeCW1xfY9j
ljgTfF5avzZJQMgOS7srueeKupnw0VQIg8YjT1Ilb5Otr2qOQw4XjdJYQT5UhMaW
X90pNZTd6ptuX8lSeeNNF40t5zyZhCrXEKZVzmMgJa9ewhTM0zaPicX3V8n+pUxO
EFnY+35EwO6a9/aYuz4EBOq7634hSu0zMgT+z+Pdm4iI4POvrxwph6qhpKffqsAH
m2rpuhgdOGE1CQcYxvzejh9DSJ8BDoHodlQnrTqyCAJ/oi75ItKsHIFgTaO7P/y9
VGKSFVPS6EKNLfiiVNYVs1RAAomVhqT5tc+PGN4RXCMDwAGS/yE/dmizSOSd19hv
4lQ38O0GjDv2KEZUZrAiO32TVzoqZGbytTw4bN7aBR9oEODi8Fi+6Vc3SRxX7oax
tZBHiK26z6RDVFzFL0r8fJgtpgwvDgoDYJ0uWvJrlRK5QZ/XVRxl5xxbBXS4naTu
UHtezc02z4raVMBHEkpQB45iHQU+DyUd41zZylkH6mqeOgH18LHe+48BX1hoiWJf
8U3SXgZMBGXbcxtkwFdhBHKVHcvtVRqFM9zd0PiYsj5f9rgpqMdS9vEmEu3HOlr4
wCINx4l3yVTFbnS3OMS3nxelKGsHeucmezRH/XiuLdXG0jFlQ765nBOamfZwZYWK
lG6WNeWbxVBmwl/um2ZFWiRubtSbQJnFzHtmrSPfDmTyWJ20IOMAOjDNW52a9Jhw
KNpAJTB/VROnXQt0cZUOXkKXOcKbWzkwnFNHvzOZkNMhRUj2lxOSIja+h/t91sz1
4QnleiM8rMcnbaROTu3GYqviwLs95D4G/BH1HTZvw/SHrnpb3bE7+BPgV7lAZHho
DkUPGazwgEtYwXriacFMXqOIVru7WWvb2z5qVF+uCGEybbWTV+dW6LLJnebytNTF
tPKfls1vuDvxn2dExVLTNZbOd00+GMdZqPzuTeK/6d+hTTLu6GhHmML2TvdvuEi8
RdeVaYsXjWF0YRKf4kANckl1FIzZuWBXpJtnHVaVO0ndlZIOC01Nrtxj9u9l2rUR
UnCuvlfHrJd+8rrGhNaHHEWVKT+3FsK67TLiR5dPQc0YNLczZOlwDfqU0rC7bTo+
/zFi2uJII7ehnxp73/8MZt9v/g2Z1GjlTw2mLBtJNWU06DRDxg54WOWImNv236lS
XGi+kngXvSYnQShr9A+sIuWQqZ3bpgXEG8T6x0cjJxe8F7N9koOYLqn4/R9KAkNf
9SddOcX8DO+7XAzu7HaOpqwpHJFcDAHrRW61KBVrnrzNjbglN4yFSdFZB/UR+4Yu
PFQvWPf5I4dOSdULA8Otok4pnddEMsXeYO2nPsRRODdHIghbj/Kc51G189nZTvQd
FkWGqArVfIfkhUnq8hML51L3XKiZSjeYx/I+5GYvIzbhWmSpD6wtS0l5XKGZ8giQ
JbSu+HaiIME8Vv7g5hMqIa3Kn+gJ/9Brs2smH60r0YazJjuQQq7odvvShr9edgWj
+I02uaYO4zz7T+jM3vINojzW8KBOgfPfjK7Bi9QzxRwFtc5a3a016Ja51h8X6Ikz
9h1knkRbt7zC4XYrJBa3u6pfHgLgttftusHlxq57S4labYw3tJu5G3wOMzcWbPC7
BJ4AaMUS7sYhdZzBdyWyYD2aBx4OTpqE2sEAAiO2UApoaCVw2Zbd0F5JBw1hCmaD
kIXkncmz4J7tmMcDhITixpsInPebo4b64pUr2si2EL5d4C/v2S52XHXyxAfom2sq
8d5BV4Vjnkj6YlDaso/Ie48DjpwoXG3RxF2yKBaYziuvrOBjOCi4/ertgDEHJded
X7wSkBkdQX6Oag9edlDM5TfglOm4odqXN5VnY9B1VT4CgwcR7AKl7XW8Ktei3QNF
7Rq2RQPRRee87nNEqr38zID1XS8IAjcf1eFu5OJubYF5ntBXpjM+3FTXlD01594d
n6aGWaLiLw0xgKQXa+DCCw2q+59xu9werCSLgn4tUrMFcuTg+WaaE6yLUbE+ucU+
5ie+2H6kfmZxWH7YsY+z0nBWft3UWghqfrNXTkhS3XD8EMnwhtfigr1JPUq7Ccry
rAH7bCytS1OiZpLLup3Zs51sHLwIy+VZmsJdx2MO6ddUsNrqgT7MYtL6IaAXVvt7
w3i83bt010LkxF2O4WVfieyENJmD6TAcxOuQtpa9RdXnsGTA+FvGPAZYeXxkuZ4b
LEnCdnr4oMeakEkQCBeszBvau26Uvc55jJp0jGkbsgm5Zx4S5qB1Ab5Ht0ks6qcY
XS3BF0qeDjGEvadqTWsmwvWVxXZmnUTzApe7HLG3b5pNwlTr0tu44AoRE9oMr9/7
9rp7UODwKq/uqnJ1VHByviDRQzfjl37iuolynTF9JXxReK8Vb87nytZtsjF5SVD0
PovHSw5qyPvqNVpbr7JVFjriifNFTH+sNnvw01h5W9EY8J3PdNu6T7usoveZnjP0
P8dkP57dgeojIKvglLyYXC/YLXhOlskXBJJehD9nC5HbliSLuoTlqN8FbPq+q7xj
ZkhswZCEEHab9aflwvmOYJrmE2CVCgwd2CSbTE+KMOxwbimEW44q7HWZ/XZ9+m3X
/S4FFLA25UwaFAKGJ9ovi8k1ZlWJkj51FAVB8DU03gqE2UafK83MTyhml7UGVb6t
E0Eould6D39RoFlPDo7BrTb1jsIGuaL1lHLhQrG8Y1vLbbkr1otCudVHSU0wob52
3RGjEATs2k2yXI0YS4NEDOhKjS9kCD2ahKuLv6OtbXm7Cm4s3Q3CLM2emdillGP8
kqR8SK2ORC7eJOB9QGW6mw7phsmWfCq2UjrkWWPPanjKOGNghlL+l6VmNYycaN1w
Op+nE5kixOZ4+QOvTVpf1yaFFJkuFBCPl5EsfrF4NZwZ/Q4kUthpXQS/p1u070n+
Zy1br64a2kQsYvNi2qFtzqrKrROWMDJEQuFm0CQub85FdbMH2QBB3JfTD6ogCdVn
xfsFusd5Z/k6Rp368TDI8Rei74biuXIW+cLJdhldMIITufdY9OGUME0lHw+cMj+h
Krvzw+owjYq8FL5ri8QWDzuFw3YWaH+kU372xHNoA6+0z73xbcBcY9MwKx908T7C
rhmkKOwfV8A2Oo1xbhU9HluDPAEdrxZYnvzQFXl/JPbdJLzdCKeK+szS9rnfprdD
wrbUkAPSVwhhuxEQVP81ZfLbdUpfq0GMKgpcFbqAjmvQtRVN4C5WhUZfRHD7JvBj
5X4G1F/wUUNFA/TBZjTGOv+VRwxgGSxG8zdvPWK4IYJeqllC5pokOuOkFTufIsjl
aiG5SNrw1M4w1PvFHC7YARDmQNgCZDgC7FMvs82O3I9drMs9N+tLSKf1G7v56/MJ
LiJjkGYB+bc1S0w01AXxCX7PVLASe8JpwImywHgtZXxQklsAlW6xkkQTMuwgsuQ/
DFjl3R+3Ayu450e5OFySwBCJCgVOPYsks87oHA0fuWuMBV6141KkhBXY4YJj9AQT
XvFqxxxZJJMK880QBr3GRgWIttowyiz/lsFHF+IVEfcQkBJ8TXBx1J3PpT03JjE+
tQdnthxbq3eqzix6NrzfWP/Y1UDzJ0Nojws7iNCPUurEHY4UuaLhP4SMgzvYhmZi
wGaa2Y1qJjutGMivEhkO+trKzTO/YjDnuLR1C4lTLf0j5UlRWY/pyrChz5wJ2rfB
EAZF6DvPOFwr39laAwxwizpn+9pj0GpnYQ2rGzFWJT18u0ATIF9nsY2Qm6uVPEa2
oVL0uWN7CbBEw5a6JPQ46af4efjca65lG6ae9RPQ5mvWapy9Jy2RHIsWOZyRbzWe
XU06G5lznN7UWOnY1OtP7651fxitYQYEyKlgy78KFvo8di+RVOhQdSa+iItxdQ/q
JoQnxTVakXfgfxLWsC98RhiKSl63Dnf5hqU5qwERnamnVz9mrDG03+lh7b5u1M6t
VoENIb/iPw8aDZ+2HDYs8/S3f0ddTv6oYxoYhIPFmchI3qvgSSG5oZDp+0gvwm0b
UBxRmCDFgRWsfSlueoCxGvV88Y8lncfU5fbdOFkc9O011uXhZR9vpwoBliXVjdFV
9QOnjvnOYDUh9bS1o9s4qZ6GCMDtrtVLT4i63Q60O1xRc3+ol9x5V6xItdtzc1A+
/x+Q4uG4BRozeMfrK+utgc95nVGJdbLY3YXZPJ/Lf6WV7jR6FMRWa6IIeKiwPd3g
ICWLfhyPdWWL4t0EApx2C6OapHWHMLBYeQrMBdvQV+fbzx5zeVkbSvUJ723QidSk
KHJtacTSj+YG3spGBorpT42TVxgbWNyDEuS9l2AjfcVRjJx8926z48eWWbx6smtx
8Lt3ZMUHRL6RtHz/LcF9eMlhuylADN5/9y2UyXle9q7gL9Jp3+ZbvwYGveQ8gFcr
Brh9Wr1BVwKUoacUcqXpqiejmoNwArbT47eX+ePwTRv5iFLP/KSbHIqv5ixK2+sb
Wo3Yv8yjMf80Mk27hJu/GUxcMa2KIpnystK1sR/nblfYttfZXs+gDN0EOa+gF0Bj
uBJNR1N76dUD1X0N2yz9Byzs5J6h9lB2+q8kx5qhy0QTZE3eMbhn9IbHxGBwsmvD
bBO0PTPnq+fWAfTJ3PwKJY5iX9s1lUbO7Zi5f3ejpKdKI4cbAZtHgHyfqQLsFYxY
fXhCXKW1HiPD5YKLCvFdpiS+qTVEJePHGOferLXFsi4glX9NX4A6PKTTN+mohi9k
PuEoGFAP2hUJMtLb7BoYQ5R05v/RoKjdL324S2G/V6FefmpZ+r4fb0oVQ/nn2rhe
rSzZFD4AExPbarflhYI3cDqqDTpKnwsv+9JZ8U9GiK+la1KtD9m3P1eV/I6AhzTD
yA6Cg+oVxqZtFOd56/UO9zspRokhRgW/ujSyO5Z7/xazcP+jk9t/IUgl+XihDNTD
NWKrIPo+TDREkEyeVJ1tGmuG2bcB4IgwQ3t7HIny19rb9aCWu8E4vAY58dV7pw8g
AXfxUpDiCi2HKIl1Hz2ZTb9Z+UbxV/x+lVrpjoizaENtJ4m52y5H1pxhVhbK/ion
esA6h9rI3U2hgTKokgPuUExWl83yCUAtcdlrdZj3KvOy+6J+QPTWcTqRNdUUAx37
BFETLmpcshkzk4g2NkVeewergDH9M/zptHXrL1B7Y61KPoYfkZJNOkFAPK4+LUsO
xW/VeSsILvqNI4iHUlgWX8f2nEIvzubxtgk48QkvZu0gs7b7lRtjXrsr3tf5W8U+
xEXyutPL9lRM44XdPm0J88NqOs6Ttbpb7bcZo0wVmgxqvcxJOZrdjt4PaP4zo8RC
qeYevjwNINr74ZUaZPoUO9rNMDutqKXJRy/kL8V1UC9QlSoGS9Fi9+v231OcBpbR
dMnfYKW1sws3+5rRWTdL2tTJS4j8vshUBg1j+X8vMqb1j4yed1U8DZaEPoyf1dEt
FKUCH38/vs4YlVH94dVx5FxaOBuivYO2gUri53geITjSxJlCMONWYUNb7E2eV5NC
RSdia699gq2lKfsaRY0K4Am00fe7i157VF9+uuFN20Ph/8pntQI/PbUM5fr5ElY/
qM8S0qj1GXgYqV0igD+//zxsN+7nYBBoCINQwHTlESoI+/AedHHfmEW8MYmdf0B0
nnYjLX6YTsFyNZKP9mXLOlRbrmC4mUxP46fGIGFAL/TxbQZVBN0AFFAsc9NJcSWs
Uuw3Rz5xc/7tqtGicl2ly1g+AvxtdCtK85Le3TQOWHdEovkb4j9pQaJ2FA/hAfS8
r3EW0RMQsIGUlz0kbjemIjzHx8QcOrXTBXVnrCbu9rBaGbo9tP42tZq+QzllUSZc
+kI07pAZV46/egVbcBuwZ1ULEnHcha6bcsjcPlkIUjFdICucaCU/b4esUGa4fqOS
IVUEGhe1/yaaFX3YPhjRc/4YZLxBe7wwHC0+M3v56Z+19OVUwbVm9Kgr98JWc4fB
oANXSvV021lTiOmo5qZnSzFwvhIp6zNFrvyLupqk9xlXhAD7MtarqqArZNpJgixj
BFfkOT9C4pUU1FujIMx8WKxrxE5cNAzpHsztU3micyhy13DEehGZsD5bwWv3Hvlq
nZQZYmnpcaL6LpsJgzMhWnDWQ5B2zymNArusz4TMAyLwF029apSUG+X7ix3IzMNJ
IY3nkhWC0+KLKawKrUb9qm20I08HumNzdJCClmkk6Kz7wgLqLV4COFUFajBvjQ4C
DpQDZyHE6jbC7bmadfEKvlvUOIikdGwnqQJlngRAi5TlbQGhU6EpVWRvOQGdhCDf
xNlqhVA+dFD+EdIW1QwG89BFGH+4sYj9i22gyPPf34ZdtietQEplZ03bD8ZiP3ng
HAGnU28erIlxwhSX3gBL95Mv1HuVn2zdhM+asr0XH9yyKKmKCRU5HgMZ06goL7bD
0Z71JydldGksQ2NsDrYPYugNHc0lQITtn/Vfy6q97srs9Ulr+vHjkvW27jJQeTAn
Q2RO+GhCMVyg/AFp8a9XbPKzQJPFAd6aFLhShpDLRBM2LqBJ3GGJFykyflgzU8kO
8kfDm5ZZplzy7PHWL6gPAWlo/GYGo2oqVt9fiY2QXN0DLwZkDHgUYyDtHM67kmBP
xO1LMUR8u9ULWcvknf+GLz9h+mu6iInwzAoAJ0k8hGS1kvjqT/sBlYLzhae8ARj4
75CL2bDeM3OGiZEIU7N6EIvsGR933QcsBz6plZ3H6Sb/UoOtYHeVpsQN8X8q+4tt
S1Wih8XIsTe4yVSF/10danzd3Xlbp4bBENTTxasKsN4y5UFYEfsy3f0vQ1vsZBIv
SYUWKHgMK9raxiEsN/XLL+3/SjYJQH3NeNW3I2tkfbrE8i3yjz6corjtpJu9Gi0u
iuNeMcCeqDX3/7AGBMvXSLKBuIyPHdVYzmLMPhYZt72M0xY79bPqGVIA2ds9QR9c
/aoGgDWyojvRdxUcDQw4h7uSg3ZKbX9f4GkPgF0o3R81jA16cV0GRvWt98KAukGq
j1RoEWBbiuhDHaEhC4AjivBlriCBbBfJqIzjanN7eR5lVFQoPdKD4QzNGiAyYzAv
aibA5sfcElOpFWPikVxYBwlq+3YKbNGL52RD+GDbVf5gZYkKwqs2Jg6LWPrXRiCe
k4saAkMVy9uOYLgLbeMVcXUUNxwImfspClOdPmoxYLa4I6yFCk8roeg70L1EcBNk
1eB4/8vfL+jRk/9jGJo6nqQHelqn6g4BCz2PpQZNIhjtsBXb2KaPuPBbkqarRDzo
KqlLLDJ8ttqzDL/6jB9hM+hG8Zf+CSOw+N4Vw/li2LtF0GeXHtKt/w1rrNIgRt0X
pg264xfNUpNylXfYhUEfhn7dh+JC1vGNSa6WH4jfwZtDxr3qvxecuyuAMmza2RHi
99oHo/RPOdvSrB7ey3TgHsO+j/l77rIm7UU6gh5dXNFPz2JcMOO9+NK3ESPU71xm
oBA2TqAge7oDMjE13De7JqIaEec5CbAGyaThbQo07HgnpIfZbO6CkKUB/+Z1eNiP
wSjwPmGhFu07KXj6RJNZkAPl2h7t2LBycrX+J0gSiGGjbUDLc6zTHRXLqDF8GmzJ
5nmQy7pOHiVzMZuRWrfV831EcuSz4QsaQbO9TQM9iy1B5Mc7CkJys6hrXP92gEUh
vciO4cJrsPUXJxfLHvky1vAQHvsFMPgapxGvUxxHz2QlY1EZxMYnJIwEoYhr/SqF
b3CR/6NzeHai3QDa58hyVN17dSc3M89bZ8TLGwsQPCSGzjCjp0Acksphc/JDqBBG
7y0CwLkdlT/Kqym+symbubpWDWBairtmEL3zj96UsqPhNn9y+ek0Xla00lhTxgbe
0wewwcc9atHqOu1VuXrSxAZaAwzD6mUWecC+f2x+K8pRhIckW6/nVsuEzr/6Rw6P
tYqXWz2AlNzqa9MCBTw59ROy1XR28KC2J5MCWXJYJ9OPUhYN23hMD6QmJYB7Oi+n
7wIfjUAdRpmwIGkkKK+O5tmhpP+P/LUrLyG6NdyEz70q3YLkAMH5VR4K7+Uo9VK3
lRGhE+xHst7I3FQzhNLyUhEU37GFgQje49CLjUGGBfRMylv2td8RblhTtdCcLmhg
dP5ueQ4EVZWLTl2P0dLHBxdz+Nu6Oa3XYJPDzZ08kEMO1ti/RiK3qJpqr1reCjUM
F31p0bHeoa5bMMK3MNB3HS6wi2z2i5K8SRi19ji6JOSoP/P/eecxu7K9wxVxq3n1
9J1LMzyoYF4bXbg6HS7d44RSag8LzBWIDC2izWQk9vqUCcMVpKfOC+CamFQRV1ef
IcM0ak+pvh1OZ1y8lOr25kH86v5vg7fNZ+iFDWhPG+yEZX7KyXpyBMlSrgPDxHdg
MTgk9ZtOpuu6mttk+svkni2mQDE0Ri5sbo01r60TjQpVZxgZe8BykhkfW5zDuNIK
ix/FcPLzs15KzwfOfhFH7oQs/3gnqPU916aWeTwSIbS9/Euwb5YcBTG20SNGA7/5
HRwA3aHhv3uRD6B3Sp2hIQSsAG8TvcZB0MtfE+0zNCmx53o+4NcK+TrM19Bltm27
mcW/tH50OGGdIEmw08Ac2uBjg70WSJzXSNH7gXm6djQVbh6B81lcAtPt2UyrAyQ6
ODgTbsf8LloKgudPdlcqGDGQGEXDwe0a742aQhjxpAexNfzhPfDa2krCNRJt8Adh
4J4k8ZuakiVl18AK/Fjvh5LrPVjJWncnbZ2vV13pZEkoovntFLoMQmOkOgFlzDQy
G9nUDNLN947oFgx11MbyXgNECtZUHSEvt05qOsjKAcNctiEx/K0P92EbVem/fhUU
LkmGjYdNaSg9DndDP0ZbRzIhssx1FEaqOFTysPi6vECeaDNXyEt4yn55WHMfKUIS
R7xKkZqsWGFULm5wRS87Gp48LxKcdjkv4scDbB9VTCH4+s21Qrfj58pWNrHWD1rg
0q7lzarJpnxSueD1wYGeOA9Uf0M8DPjwCm8JtQZewR6mWv9lunFkQogZuXg0/ISH
16A4LhSavhCPoKYp+1sYYso5vbbmuSR+EmlNyZPGhZkhMRpPwyZtZJ+lsGR2g9OH
nWH8BRI6r0QLgeuHweN8VP/lEhAfLd3pltg2hOfceDM9JB8o4A7B+SxaRjymuEKP
1NeIWGTi8sHeurFpSuHw3sQouy84mzT9scwVy6J2x6neE1Q+V+WE/HNzLBuwjn8X
kdLnKSXvmAaH+u0/5VFFa+SXnCFtlhveNy7s/cofnysoEdv+9ZxsYn9g/V9CTmAG
A3uofs2XF24An1CDYA6mTsFU3o09PMPr6wHI9piEJK3LQv/8mCL/CuvJIjRISZk+
gP/u6gdvL4ugQ/CiiE+ebOAER+USNPCDOBoNYsjMqt3bfIhkjLH2sQLPsVWhu9tq
fDGFb3AfTED2rNEikbl5vb6DnIoTLiTz2pRAHMSKwsCV3glMYTltKxhF14rEt6SR
sEvW94caJ5MnpA7AfUE2Tmu8KvEECCFde5EMXDhF4obhYwZ7rTXT37fiDGl03XT9
s4OWATiPFPAGMymfE1uYCP8/HVlcY4leXMHwOx4mxR57ySpDlSRhATLZwokUIji7
DPy63NXNme0+MhgTDhqIKxpDCf1eLXmMD+xMcYgN6qTgU/PIKaXmB+sTX6Tguiy2
qI+FUAGNJZgfLoKPAboiWUGAPS5IWUQ6ogERs7R2NLVD4su8pvz1EuPvqlRCBcvh
+Ls3z+xyCO9DZTT+7zZTY9whNtdh+7rfJb2qz76e4kAfytYJrgg+6UHvX4gq5S91
U55cHCRcz5NxPgFLxSWXtMNQX7uxlnojrek92of0jd+5CKurVS0qWOVq+V6JhCBb
AK++Z8OJmdDvb+ZFmbyqk8LBMWtbf4nEywenJHJsrhtAgG8tMLZ3LOB/38dhRMEN
2fPTrlNeuU/pcBhG9tl11bYLIMjRKxiQgZ1d6r9pi4zvdb4KEFqg9oBW3BPOM5ZB
kvSFZsAjgnVF1e+T/fmgzGN0VGch/+llKCEAOaGhJhTRz3rlZf3uW1GATZe7fNM3
uocRUYxyROSwHgCU1rgDwIxt8oY4qpPBLfU+eyqFreUg7UM5aDpqOdMQ6xrd7Lhe
APhWdpFk+DI9R5RekVj85z2zx9XLoi12UjqCsV+zq17zABMj3v8KoCBpE+Eoi3hq
+p0Th9xJxxYPNq3C0cmhtXJ7bhBJyDuDTWItVb7HfsOmbbcGTE27SpiG06iml6By
+dAaJt6T4jH0a7bOmYzgUqzLQ3sD+IF/Sp59y1PMEKgSeZXY/KLz89h58YGTzsds
RhwL2j2uLVF3V1uWfiviYHojrqUWEDa/326aEeKlFS/NZ9tSP0umaJorWVOLPcrE
CZXNCXdD0eGk6urlF4/aax8SGTNRa6jR4Vbwv2pSio8Orqvhg0K3XopAWs4NgdVf
cnq/jB5LlFk7GLe1EPpFtsDwzxjTn2MvHk37OD8X9zABkgYTpD+FiZ5fUUWL2QRH
OvFXytVgfSROgW5+qia5crgdQRmylM7QUhKpxExOti+UORup0Xw5nKKSN9Diu6gA
BOFDTYj7ynvLyK4v4UF62FNCjLK8o2olINAdIG3UW2LoNV6nNWffpIls6LymtaRp
lzZvnq4SuPcRWHep9ohonMrOAmyTRcsm5/q5izAnZFXuW1kyQYqUrPk/UV5DKG3o
br1bvgdu6IsINnZQWxzPzm1Pe/gqrDghrkzFkXHke1LFEl9u1KoemIblDo/DcppZ
6XZuEQWmcnk3mCTSs7J3UQHKDy6puX93ad7jnALqEVLCWMQ3C581g/mOQMy+iCrW
CsFeRzHfz7URDE3D86G1h/odvc0+vnL8BJ9ZS5rVRhjZ3EqwWSk4Sqg1kdhCbJXi
NBt2/DOVTLtt46U0MdkOnJSjB4i12/HZfyIsyNk38EGv/2oSF1TMvhYTQsYDaGmO
IiRWOPftdjftTrWH2pZoOIH/XIksJjOjnM/nSqsZmfsRVd4YhS29BU8k3ZkXB6UC
Pwu5oe7jLhrU8FgTOdyFJYcJ63D6SiI7JG5PH/pqcKkQn93/DFOHaxXskDOlMtI8
AhKd2Rk5rf3DowWRn9JteGjeawJtJY/MPq0pzCd4Wve/erUN/mWCIQ1x1GlDDmIR
0SdCkrQI+iVRYePl9JOKi/y55jedYtJlYKBut1GbDqKBQrhFa57K65eexKCrR/KY
/NVWMX60/iym12hrqU85TZWWoHkpmYtxwrg5RYykIcmfBaaIqaXP9TtXhYCKyFQM
Z+EJx9F0iX5OS6CFrhIHlAlmP36HNf9hh22vuTWTFc3W+2A9qLcJqxRYSmSX8atL
J5zz1VZhMKqDm/EOIVCUo3hP9xSC71/7XHl1YzYqiyocLAVfsbGjKXMSePjSAFBV
IC3iCPaE4BLxWkJelqLUTk6Qca2Od2uCIV1nZeJGnh8skY6L92+PUQsqI8X7zFEL
VPiNvkJeVtyDz1DkiVTqwkRaIRWd9dIMSpkzF5Mhy+82Et5gwqF4CUay1Or80Mej
rMM4fSnOI68GDZQTzdxwF3i9C/dRoqr8vK98xbtH9nabXTljFdYDpC0DIHp7XLep
dyvl8BF003fuxHDAwvj3I2FWCK9YnNHOjBog1yHc3oWOoO6Vv5j4dbbkB8iQtxLJ
8Plwzk0A/RpGzgL+wcxaIY7Eli8vjMiJ3LsGUcsSmepRQ+VMF9H1IvQJaBSjg7px
CqZm/2XUSNEPOm4VEB6Sig7JrToKbmxQOIt5yWxTqh14kPN3jjm0d/mTQcmI38eK
N0KsRjK0sDj3Ji1cewqoO/IDYK6iw9DC3mZUTq6LkliH0WU18auIl8L3zeUIUhGZ
iumMUeJ4pV2VgWbXfugasmgn4TACVOtlpdsBzHeTZznfcqCqvtfd470lhA2WfVMR
m612MjkuRvnqB0aAk8BVKuFlPb0WLA263N/iGnL7qsJsXMOvcGXySL2VeGULo67y
LQNUcjYTPBa+TEWWxtu6MQOV5jC3CB5Rk/5GcRr3rEq7zUj/LBMaT/irI86XUGsY
Ncvt3q3z6U7gFErDvl1bbwPQBG6WGQHQ+yGhwCK8n9fhcBJM60L0vEdrh84laJuH
GjPrBMNKyPFf7q6BX5iiFqBHSl1nJsFfvM7f8TiI3yhM6VOf7GtWoe++L3YKeX1L
MUrPstlM8Zp0kSjRE9E98y6YmPRu5R+95v9FGH6N5y1DCEGUZ+NJO0PpaklG5Eni
0Ts81qtFrsTINkN3lgj3Tjh9uQkGXQ/TQ3tQhzWDH/68rV2U2X/5bEVWoars1VlJ
pWYckAdM/tQpuZYsKWtCuvyoXpWWpMQ6ueqj/vRRX+Rlc3118bHd2fdGTY4o4dvL
K7peb/CvBCR/J6KFQtLujeIsN8Kogs2digTy8ammBJz44NBzumW8cKHqfuEi8nRb
HWuU9xUuwi6RmtfEPFMH/oNGwEoQJkBOrhFIVdahPxfMEh0fNMyL3Nxh5WL2Ocn8
vfO5/qdr0nu564fmmOf5w8QyN4gspdkgPuOML7gnY7bGMp6xyFkXnVnKhwIT5mZO
svGTMjFcxzVdQiLYRZRmAW1LNjScbGW/wfcuMJc0fyTAOikg/hb53V6apyh7BVuT
81hV3QuIsFH+VHXT9ryNZcC/VTJZPkJZWDbiyjZuB6P4qempo/8pxC4+vz2yzlrm
kgFzsz39AlpPpE98A95MlTPUdcNbDo0yT+vKauXpBUu2ef2Qq6GmoEntCC90rExM
qtbd88TDvfHnaxc8KyZ4dcbSqOcWRzJV0AQyq6nqPg8uSmyi1R5Ztk6vXwDow2jW
nPgRDShHl45P97Ab0lUr2HP/m5MTByRQSR4PWfis5qfVcSeA+yvyvoeH2jkks9Ig
KleMn00CjwQkUipCKq9lantxA/MFiF69ndZ3l8Xart3XedPBXvUjkbZaxMOxCPhb
0eUJkSRVqlrHbnGc+t0Gt9rZ9DkxzkOJtV41bQnzPr0vQ5D+YjSAGbMzoYuRWT+X
Tk/23bEjCgQjQQ74RtrZrB8/IurYqphS7fl8cxY7bvo+YwE4BtEUpouUx/9w614J
savaszFIggoviBIHVPXC1N5Jsq3EY+1N2u0ax9XPxngTSQYGfcSLF43m6OriZysh
A7ClH+euklNpjJMD+Vyc3uXhGU6gC8DD5uFidvvDR/PjLxgfcUi+Hkv624fuKWV7
q0WUOIjaEXuNDss2ffgovU5DDgrQ/1U1EFaIEiyAMdBCatdEsH+mw9rWoUkicAMo
n9NrieuBB0/mTJgWk+utQc5/3z+9+4PfguV4CRO25ufQsUHXyfRdUwuAf7f65b/s
aguQ70+aCYPc+8UTHFFWy+qx019+aKdhYb34BShVMcFyFJsv7rVHFYI9zE6e2sK0
Cva3d1Z+JVzAil+Ro6LkbaMgdBZTU5LlcXJTi5FDlrKO73n9KMFkMxP4iZvbdYHX
sQ7f8n1K0oAt2eorlPHzcuJgx8V28i8II/S4uzqfezYFJqP/1BMuBDlW5REjUGvx
fr//Ewe9YuJWsTlzBfOq9ad19FMDbX52W+U4AJKwjHAxCILp4OHjIreUsavNuyl9
3SSRYZMLw3ATHKCKX/0+U2281DLIUzXN0SSnDpX2OBC82AySjcrcTIy5d3wiymok
2sKyLVu8ztowkrTkYA/fFIJ9MF2pDYPNkYeRkmbzYq1QPBN4Qy0GbIJ3Z/lEwldr
G1amCqJhvyJ6+Unx7YJMzvHMrGD1rJMwWIuOfLewaBlcVlB+zg39RYb03bFbGgGC
FNDnRm7RJTFuDC3KkqSw+ObZJ0BHUxdW55vj8e3AXpnmKwShBW/UlQdcsvNyA5Pe
gszV9oxVCyQDyTIexQeRs3u6aQHMRABPFHBdSO0aSkwEsH5A9xbk0DmVccndao5B
l2S9j0wi2GLsB3z+gGKIhPgde/ZtjHqvRZRKBCIvgm48RjmoMAtc+sBtbKDk1a7c
vHBh1OpowLsl16PM8Dfgz6BfyNvBLRu5OX2Yxjc4tR61u1RBySHGxMiw9oCiONDm
XBY1kcZpEVftOqd4YtvKA2+pnV/eKhjfVSal837N2DvdWnvWVULEZpToVF3QYIPW
mAU7Y00m1q9t2KGPs2x9o6XvUk5nf/+U/c+fgyN463czajM40Qo/DQEGWWsm6k0s
5WyA4eBov3jzszQYQdq5k8ItvQWaiaWcqbjuGecEu+Yx6bqFVL+sZ18gF0+fLbuS
GUwlVt3io+mZvMrjORd5RTz+nZp7waATIhdd63WIscFAK0XsH8JzCn6Hp78fBH0r
6dPd+/Kv1zcwi6+8Fh9CqfCcIYeB0mcP7+0Id0mX4EvXdNznGuQiZornE1FNdN17
Q1qgtn0QxR4r2mT+a0DFz518dMU3M/9Ou0rO5knTZ9hrn1JThHIcwujt6+Pef8Oz
VnrC543MnpRPrEWC31BBeDoB1zQexC6OGMQxAtsZHu9qxPlbCTz2lu48XTYEdyf9
8eFQLjajA1JTJ4HtLKJ1clQPtI9NmR5fm9bN/owrPK4kSTeZcyq99f91pHAzANWW
v0t9bc9L0GhONQPsS0xGe/7gti6Zg6ldzJoAyCQEGUaf+3ji9lfOGsKiMJFUeLE4
s/Dq8gMU1d0yxDUhkRnFGj5Li4ayzPPFkBefMpkQcjEmoWbuzg2dt6o11U4A38zU
qxNxKNqfAtj0GyoOggGF50qY2hmab3zKgYi3HzhtPmyIeSb8yEgLN+OuZC4GgWl7
CL7gl7/1NvPfsbGMEU/6IZXOr2qIOUNME+vylJLKnBlgyglCy2NtRa7WaYpqkPl5
QWJJ3+X2Ywi1dXaKoRgYG45bdckL5UOelbdsLnJ8u1ECIGvQs3leAeBYtEAAJqkf
sP4nRdzvg9uwmUdy/Xjv2fUBoi3P71UiemOKMOsk/qZ23CiHEf8hYTLfZcH3I9Qh
2DE2eYsH5YTxRWdEy/SogwvLz9xFX7E2YZHc8a8nD4n5R3JMTYNzDIbSgFGUpr/P
CXvYi1ZQfj04n8I+gA4FlCDvs77WxWqPotNcSWLNGTcR2Lm3N/CZ2ukfE0gEOTTf
xhL/7618XOQGpb+tLIfhxLJ3THFLRVbVKYvm5kNaa3fQucMVCWsulKViBtCKh/XS
aas+5+kcaIheDxBKAJAtvfyXj0x2t9wregcYGjJnMnr4Lu2A7KIcGjIqMm0ezx8u
b1foY7ONMKs4f5mx0i1lnd3uO7cU9b+4i9XllgLgZiRyE8ddM+sDUQgaFHugslVM
djqNBN0DcuOCiUy48KHROw84ZgQkF2Iyr/RuUzcjtL4CZULLlO4Qg2/a9NJWNVT8
xHuDrNAWWhsxUdKmoIEcdqd7A/QzEN6aux1/cK0k6IPw5IFSSrYmyXqO0laKFH89
/WggN6uW2beeHZhEAXrdqWDU+zuSRyVV1qa5/YkaIQPVtNo2gYdIWe2hGnkB+D5e
sicwB1yVZ2C0dOjBEid1DQKjT615owG0NhOmZSnXRpO9QNgno92+9I2Jvv58HHSr
UopBj9aH2omK9eHYsycct+xzkLs6St5A6Ubvpizwf7BMOEHClnioU+Hh4juUdUUo
xGXrfkPot5x2vitkSLi/uEiD0E9RVQLr/6h5YpE6BJkvW94Ct/ArGikE8OC2Xz6n
MZzFVFEso9aQAJzITU6mB/nL7ym3bvXkfZPC8KqSDGE5YWRBmiqUwNAkmEhlrfcF
svoDLnKAPVGnj5jdTSSuKstINEazE7JpLNyJC8ZKGyCHj0EQ9PN9FJeOTaQTCeVN
u6DSLNK5KIE5zToT/IUzeiZNmHAVW53oiN5tUrPHD7Sgup31F1dd4wBAo7HT9/4U
f+J8sFL/6FshyI6yArjhyccp7epLnzqS1O9Zbka80adB+HG4ttLv5hII8zz0xrsi
kEeewno/TYxlQggcTDbZFut13My++NMgP2Mz9VG9d6sKuVoA1cCS0t61q1CON8LN
pnIY05CMnfLt4wiWhftUlvg0xWR9XO2HD9uEYhLXE9wqCSu2ICmHxqX3m2UyYONg
npc1atq5hgVBTsMcQjm90ptYqBJGw2EFS2/PQHctXMWfWG6yiOIba7eRqzV4HZj1
isX20XrBit3tcgMB2pGlXPFkoXJnErEfnWXmSLfzK/9e0laRRacbnHYQcU/mAjkT
selLbFIikTqPvUK1edXWmSieqwaNCZPE7hd2EW4TZLMaDWMcdGWaqcBQgR4Ex9Kn
DwIQO9DnGuLR6AmC2OZenuGFXo3OYsB2Kla3ImtfQRMHtDoAVgo95d/QziHQYsRE
Zzm+fMyxAlsyhxjP7Uh0DKkpyepMFTuwvXPh9EM320WczhVvtgAvqDdAf7o3wPW6
WACQxbvbt3H+fBfWR77owfEuRFMuXeBY6JiGz5iiYoaZbpg0twszP8vtUDRXcS6h
7XnZusSTPW2ntTfScFuTf7IyyaUoz/xFzv25T6ezvr0lJPo+U8H4T5DuGkEw/OLQ
RhpcduImrVEg+4u9/WPteEyiaXsXVyqbHIjEz+R91IVFd/WaeL9lxMW33PyVxtlQ
hA81MsQ6DXTKwm0fzGk7EZQnz3JbpzoQ0NlZE6lpScvz56vPPq3ASP+GFfwQnxXj
hPWlRFLvqJvd9yH0hczmiUCGY98Xz0ZDWpSXxDOyvWzYt4suIL7WtjlxjTbwNA3l
5oQnwlHmPoa9N5UZQNkjxqIg2nB+DxLVg7n67bj175k/yjLpYAMmB3R2PuYshRSM
96wiMFIc0x0G1LMxkQvjNMUQ/DcFj8xJzphTBMyLS3WVtx4y5LH/RwGqdc48LFtb
IAHGVhhhdQg6CXKojqFKDmvgaa1xcLEzvLje1yNXdkbmwok5M4JbuX4bVl9ZL2lr
8ZQZuydkVxk06v9DMjijO7k0BdPWiX5oQhl25IuVrkXRGWEfXdo06C5qu0EKen0y
uq3kUROYwgamJlxfYsorty0mwCMHqdLcZQLfFhEBudWWTt0VXmZijO+97YQpFr9o
lFLwSt8gngRwLIvxdn8CUQSXOZ4tXXZ2rBULyu4A2H9KifzHm3vGpargvhsDXsI/
SKFh0X6DiM4WrEUVKI7fJP3jyiXzAdE/tdIu5k14pyg1bBF1mM7tWg4f53IlIFe/
ya1JmJr9F4HqV6KDRKNUyA3gY0nZte4EmXTsA6BEH6Q2eNDXgxX5praej31JVigU
jlUXOtKH/E7miSz/z+YRzXraUNxDUKfcU0nSNJQeksVpOXKE66JHQDa6ERZ/9MVZ
BHGDqnGqVuKC53pFcjw9MXxq3JJmWgVwzRnswhY8E8of/Q8TnDSs4gfyP/C65+vP
mbSbOKkOUUK64/NdwnQ3PpXFcFVL+z9LVdtUJ2WNJTkbwj11CuZJgRWZtpoZAicH
UbF9INT/PTzNVNcA1MDHeaflla6K+xlB7mIV4MahOtQ6tLvSya1YIydOluQYNYyM
gtdhQvuV8h36EkjsYWe9CohUtGm5jWJBv1cKsPL+EZGvfz6lCxviCNo2y1R56ACb
4aJ6RAwJ8qj2wNxqx7rSj/msG3D58NsMEKKkuN5gZAi7apbWzQupCkTUJQ6LKL9+
1qgmmJxOYSEkSnxPu2lBIPUrrNT34ai+T2M7BN9myUQej+YzG33hQhOyGFJpuOvO
dh+u53sNqtSomUXrAiYLcNOIxdBAAFJZTN2xX8KRDPMVeyMQ1UOBnw4InmO0+npw
jsnaD2c74M1YSbVddI8Wj+79QytVmI3h4RgzXgSngz09RzkQm+SACqqNfaCgLg9b
oyoZjVXAuUEInnOcLWsTxsmCh7lnWKb7W+ZTYg7wSWnmQapqAQGbwZ8BM/R4tkvG
5+PZadZd0HmBq0RjXD9UT815eUIfUj0scXuiatmKiACktID3B6wNzFE5mMFC14lZ
NHij0OkIWHOwJUnbS752Khdi+lhMXDQcQBQ0o6xfYv/QOvsqeP9clj2ecFu9cQck
wU90ASsGyTNX3sWYluwZZQtC1TYJKgZX/qWTRxRwj9MkVUu7gOXRON00HQKrAEsG
Fzig4llAHlOJpANUowh84mElC/BNJ/kz1NnVjFPHcB4uEXoUWbY1br+VtfC8jZDc
XoZJ/pU4Wf3TsI01Q92XCCOiW9G8p46DwR7RPFYRR9vG6UEKoF3Jlt9ugzfRTqkW
KidPVrK+MMw79spgUjz5KonySK644bVHmsFIXNVG0dHElWywfu/IBAzycBhbhcbR
WCQme7+S5cLoINxMHpnO07RKSLJZDT5F9U49GdXT6hPERTU8zPV1JJSypBeuwb8J
zlYVLVUSjkFyKVSEmwa8LphNntof1EdM4PcICJp1Xjswj+2xmwl2Qxv37f4mB1Nx
+30AAmE78RoVe+IOccU81rkI8wAjve4EAl/GpoOJfOFecw0zb9Aqhoq8RTuY4gYz
t/xuM8+atIuEhHY9u6QJYM2IsBaFc+mkAXknr0z1JeuPSnJyY8tF2WqpDKybkHCa
XZVwolLGfEmEjMNvlYlL7qsIMFRhaLMLrz2tDO++tSB8KQnoFwOHTZtLUGp16vZ3
KZSMzzOEXwE6pUZhQVQXr7jHYqMK1YeM3Sgv8AokFsTTXvcHnR8XuYoqELppK280
9UnH2jZdKLl27uYW6U+p4M+C0K4/dsyHNCsuACCZZfDRXjiEILfx/qRBrBVjuJ3i
l+aF7NSYj8DaF415BxXIf1tOBGH5AX7KgEDcWJzFixeXw8m03cZn8bmTLWm1cy4R
T9XBKT2kPYC/W2blSMVTgtAfFmjjzv1dmkfYJNVBk1Fy9N+zM5IZE0gxVwaQogZN
YnKWMkFs464W7mzyFK9xd3iN76lbDlmcLo6LYV+AimR4HYE1wfTzMPnn75Z8V4OB
ZDwfIRMdtru8oFMC9eYj7NmM98aRUEUfFw7yHFb9EXXykjgaV7ktKIUCdjXIegGI
BNsExTteO/SAsc3wjjHy1OhF1eNteWu9JQGctb5Ov0AC52t3Bp//svELPz4WCJws
OIc3QT18Jc7AiLF02OwUJrpnW1lXS7rJbhWj3FvumSuwA9PlQufutNY+E2xWpqeA
1NSHItTO/kNsScetYkH27WsSgiXhBIMyQBZXXE4y0nmK9/FPrn0wYLLf12TDEUDa
CUPbr+W7b2b3Xf5AoAyFgP1BGKeI4NIsecxpVLONK3+OFi2l8rrvGK0j69/Zb2tJ
1qROQ5vNqbx9KnrbISNdK07hoeBa/OMZhzwWhgFIwOvbO3HEvCbEvzY2EWgNRgO9
c5ipkX7yH3VUU/km6FXMDgoiWKYTKtbtnJy9UrbAFw86lM9YTrXZLlzROT8TyEEE
WrEZtQYvBH9MKe0klBSsxw981wl4DWHJr7eozhxewqapauV7pBxACYWZcnROrAvt
7IjCg93wx04BWII72TkILm+VhiBhITYE3Nk+qGuUQfUSQIUSSKeShQEcdRU9O4at
B443srr4+tqecUkMByW9zw8EkOEGCUomtOg2Vkqb0peL5pgEnuos37zKapEZN0m+
rgg57d78EoyTaMfv2f2RfFUDl1/4GU43Cb3fXHld3+F4t1OoFLDY/abasb37h4Yz
WCIDArddfva41sCUAD93ayDpMDwa4KEE2j4PCnDA4VUhYtVtpW8bldw6o/srWgBp
+T2uoPFS2Muvfq8z3+ViaGkdwzMKZq2OovW4/alFuKvBfL85Gd+97M5lT++GfIZ0
zFjlCY7KCnCn78n7gtgHZkKYP8mxrUbfGaK/5ibWZAefSyRKK9sGctJ96uZyCAC0
TytLALBEFIe5OVzl4Vi1SQScrPl1Uno155p5v62KJLVyAS+Mr+g5aTNW7wCBEXx3
nx61LdcZfBYnKpPSWostkk4KRZdB6VgrP3blLw6JUqQyQZpKvNmsdEwCMWz7iHiV
yPAN0nvO5yw77dg2fqTBzPL7JquAFQ0ZS9185TJ21rMoAwL+PHYPX0fEk/HPBq4c
KmfHbrS4kRroPxOq5diYXzzePgtA7oN/5i1NsI91nHchwgLXPF/UqYAscBaxmihO
GxNx9X0q0sEfZyadd9NO5GMhRGPEriOloFJB56DjtI7JReXlq5Rm16iNXDt8Wsxa
T/C78IgjmSQAMKCJoo6FDdSL3rtqMWDt3YRqfmUD2m8FC2I+AIBmrR5+fy+lnc77
5hkFwFd9ieiDA9hmotF8kQb3tnIknITVAA0mmsbKyKl23coapQbN38TeVyyeSiO0
9+yVi3R8RRZsn3JV66g2ZZ6q1nmtlxOhSxX830LZCpSblIGbiLPQK+JHLqvLeG1f
vxLofAP4xIpHP2yX8FPk4tilqRGCjM2p+Xi+eSCVrdKsRz1CMVCCIotCIWVbGKzH
Ad3z56QdX1bmzbuvSizeow156WvzsP0BrZwZvzEm/ZIUl41UxWlpTKhNKg8hbLmy
0EJpYedF+amPNw78/UFPCNblku4NCkBPOjTT04srHtGwQmT9XGIt4W5rfDHPuahF
xHd9F8Cr3EZ3yIqxSoMr10Yw4PnhoDmdSkX2cPq5irE1gQ9tI/b4/NRKwdMpwkxA
7Fu+9UaoiG1d3GqhUao5W7N0uIjfHAYeezqT/kjesZvUw0Unt90FHudMqvay4joC
cdcM6VCYrQc5R6HDfSNjlb0BqWCyod033HMdQ1bfyonsulZbhlHWhutdqiT1mr0R
0MpYoLLs3+kR3hpW78gnvU2TEUNu/xBhUASGthl3xbXFgN9ZCRwz0v6SZglCInG2
2+rIIWOsVwscD3uFmIYzysOaOD5JPcB4yg2OKepAEK8CqWzaiGATBfDt2Peyza5V
B/P9Lkym+GtzLXlaOepa8MBqC6vTkRLBVZg1F03bMRR++o6RgOFnt2gGZWS0D/Jl
8oCPlkkDaS2gZexCxaBJYYqCiMepgCW/u0SPBm+a5Unu1+gPNRjh6qkzJOLssGbv
GZbNQ2E1+LiEhJRHNsPrhEh1ZA6HPs1iRIckM6YIYlDFsJP3BcV7xnH2WmGCWkCu
VVmoZNy0SVsYxWCuOOR2QlehM1Jm19T5WVkiLl+Liq97zMBwcJj81ZAHzKMpqglz
++S/UI1EstDprhyJes6c8O7/PQcrMcKTUa8oDOsPTt0ZT+niTmdnmyOzXDsUHgPu
iOMNw4i3hqzp0KXIU1K+Ds3XXS7oPvoRlyp7DitUA55xcYeocx56sLF0CDxnxsln
B0WbIEfIGhuP5m0xG/JkcI4RXZbZr16/Fhu/4tBxtgKGpUP9Jhip5YaF9DWYSxp/
ERU+Js5S5xhe2lw+bJjs8V0DaKo25ZOoCDS8Dtp8By2IQJPpaSDApYK9nD4VSpfl
KE0W2cPMCm2tJfTfktmPfPoIvKWBvMiylQSaJwS+t6su5hDIfqau1W4tzd0QF7ko
UXdYJxsEySiH3/17AZiWiB0k3BYorHIASUjqY5PwXD+5iXi50GeRv9X5NFnrNxUI
399/e8NGm2U/2MEgb1CKRQGK3R+uAvL3HQ3YyDotypP9ABdArpX5XevI0/iylgEY
XTSaKIq0dzdoxNkJ7VaudY4bYB+HtvAoPvLUpfcvvsCUNv+lpLBW7mgfCJEVd0gE
h0hjE8uDkJwhgohqTqWZetbYSA+K5yNF3Eh4fMYYc4Eg0Gl9HoBVXIuhuDA6Uxww
mn2qczM4ikrk3puiuzI/ODZwOSI30zAh9GCWaS02DphIp0+odQKGu/eo0CRQl0lw
01zSQaMEhs30OkXbFxIaWG6UGlU4KJfCWs2i0KnM+YlEToSzYBhk0ZAJEGUuXUGh
tnGuLN92PjaoJihoMdcyVVjFMuji/ppXVFn2wYc3YXpmctd1bUIobXLLnWSzb/+l
bNR1jF8RNeJHiN3dA43N65bxIAft129DG9eNw9MCM9x/kZfMIDXhDwTB2p7obx/U
EfqFVGDWf4FD3HN6LZyUb9l06lbkHthDZsQ+eUlgIdWipwlJHK6jQaQBTtGLIOWP
fTV7NwNZZpKGtTnlvl4QOyzogYlsJeNfwlTtCyD414tNtoKtRVWJdWycb98wMaa/
B5tNfK1SfbjCNtPaFOlUkAbbIMGdnE8UCi4qtl9XJnNJEfc9hAouiQZD4AANkBqt
i+9mPFFcF4LH2xA9V8bYYL7oAXo6F/20EP6i3KeaFQWazwnx+wIN5LzffcX+Qkpj
Fn+m2Wu9tOFCEmiJ1ChRepBvlxE6+SzWEcFw952p2haTWEEv9NYeI7Y4/358/vkb
4cvjPnrJOUTcy2osefXiP5AMMOQVkOGSL+513QLvqEZuhmABooJFmykHDGGpncwp
v76kua7/u4b/q2IL/rKEeYF9SykHlhv+WBvT9AzpZzqYPUA4qDZNVBgY7X0WYVUg
4YHuJb/R1LUCeYjjRJ6yZb+bfzdDBW6Y4OCohqm7J+uOqG0NHgV8J/BicQuQg5II
NYRDlNiADJ/oSRhVrlQoWmkgfBorHnWn1XjviP2fKeG5KqDytL7kXBVCVCAc/5UO
bkrrpbVZeYWYr+KSMPicUfYcb842qQRiISmaysDsm/JDj2KW81gn8A35vFBZXjl3
qrer/5PHK66X1xI6ZeXVtFZ1jW6l638iFcpFLmdYo4x0X9CGUQ5EgACtA1pr85Wy
ckQqveezRhzIThEYSoCC2nnx0Ikdbf54OpqQ4BUvZaWXLI/9PEcnY4Sb6thwNkl6
hu8ld2aDbkdOjCMeGGCOFuxjydVr9vStV0+HhAeaq8oFgVLv5+ACKWXEWS1ZynRK
oH/W/1KqkZ20+K7ggrFRtA4ZSSQVca+Y1k0o9UZYeUH2nsXazqjMNAVc8tt9MkU2
rogUbcTd5LbT8rxvM5Fk7pG/PJhd0SNMHHmsYFz0Caz7KUG293aymvSQFp06lZPb
BZsgR/cEA69tNbS/jTdzP7z1OWl6c9ApwCb97PZDFrE6tfFOkibhnedd4JP8wGRu
sS2kg3EU9muTTV8kgR0rGlF9CCYrJOTmPq2I5U8HctcktwCEE7eCIDH2Z42aIonV
dGZff7p/dFzZ6FEgK4rtSjF9kQXX1SxnGHwYJdVcBGI/nUCpX98b2DkMq43nW9K+
RRVLlE+l7Jc3M2Fm6W7NK3mkFNqwWpX8sU9OkdM4figiympOKx7pHNUUfgHFWeYO
YxTmae7y1C38+hxWSSzqOGAodesaFDdvY0EPzngb6ViLbrs4Hpix1V7/PrbvVSFf
evByrDDXAnETslMYcO/+mcDAs/rp0B66g7W/zBgH+tMDn7gt3xcqrJPGj+CYjnW/
7y6k67xTPGlbXg3csMpVALpHqhMpDE+1+24iEF1xuVqsBhMV/3Q3Ue1juygHuVfA
UQxZnS+tkqv4/eYUlTBuquS1TEvjJthDTqiLb6cEEVpADg4AVpDyQl0rWoRHIdEz
9AcIPd+2/vU0DmXhs5S9XLaS/utd0ZxAJP1N0endu+V/yt7xVyntvmvQAZdG+IjM
tA9vZO7y/LnBwBmaB+9YsWph3WN+lA38LjTXsL0xYDC5NHpi8of7M/AZIORNQmyg
4o07QEuy/YNNnsPaeuyxelatETbqawQVexxeBd0qMiuSmcevLJRDhGLvGQgMgHlq
8LV1ySAnZK9iGvsMJarAsexYAZv0mQoy08sSDaSS+Sjgz5jPf4H073IJctTXAi4T
EoZ5YdtEvPIFTvGW6LZsoLKGzJIi54j6x45LxcvBqW0S3LKO3+t7C3nHcUsM0Etl
9A16lmurjjqYmdDeon3wdzAkykPlX0w335SjvFTSiEqmOefKrIDbQPz1SUeiCp60
mnQKP2sd5QjIyuq5lebtSvj9UvmweF7Y+ziUvD+z/APfU9qrQwIuuDYIWswtmTn+
afDdx5135pFjxSAJ8lXkj191cByUdZksvw8a81vLoRxlk8Rq5igRphRCHAaHbEsG
4y69Y9jcPuB/cedcGH4NRIEzjC5VimLc9gYU0K66Fljv8KxBksIl3jw0v2YOjrmH
gQBVc49v+/txB3F98pGYLSzLPkR5Za3LdwaDd35HQS7HOe6tWhlU8bGXA5ZONj7x
PIq06dTPxit9MlHuW+rrQgq9Kn9s5FzUXSyNhZ38yxqEnpn7EkDSpDBThQiSLWyl
uHsRr33gGN+lHGIOTm2O8ZxxdQukH+5tsY2rcy9fr5de5+qQWNRu04Gds+Y6v8Ls
efzR2kzqsSAM2wzv3UGWKSf9uv8J82zqQCNNuc3VbRfZxu+611IgcQATzsxtlWOo
+3t3z+eiq2AOX6p1nFVoFV8p5bLwGY6rG3sYSW+JE48aoJ7RHy4iE4H5MD6KVcoi
x0paoGDymVhV+TQT9nvbxHX3op/IgkfBNSvERtT7EpIOGncKzLOEzFsxztVtL+1A
H+qShHZdclr6KYowb7xddGOqxolGzlEwfq2O5AVtYel3A2wZnyxG5nrAqLDXzf6H
yKCyUlYc0HyInbMgTS8NJ65QRLNIsLtwNZg7BVU+RdhDIu2c3cmUQS/khwvMW49v
UnnnlxutKHUoa2zrsH9vYS/gtPQN5COFY2VhpcfFK6Jw9wLM2L0wTu7lEp/SzMMw
Jvb042H351O2EdmDNkU5SXcUjesxXQcvDKHhZtEHQOTJPwrx6yJQdwy6GAak2tbY
bYXXGVv3HJ0T0ZZvV58aTmRjG9N672Mae+1YOp47o4yTZ21cfXJM6l5g8UrVdOb4
2lXTp20XUYphFW+uDlNKVZ817ncyEnxsElso4hEVlniGGvpm3VhuyxbolbCtmIpQ
Jb3DMGF+NAZtZ6iC3kzch7uGDp55MneJmipCYLtxexH1HVRiCsNyKLzvp3sFVYJK
aACmmXCtbN9jsI1xkKMxtUdmDtmvQToKbvM519S3aGKnrLRwKMmJL6gGP6K6Klrx
vzMUTmdkFALCYLd7Ai1qFaXiWohH55ymPJHfgCnJlqM593p9m7/IjGk34owiDh4k
MMoirvk1tffqt/uxjG/hxgTeaSN5K/Acq0Klm9PZr7ipn8kHX9HA2YUrp5fFelx9
SrKHuGZzOMa3XRRCDJgyEcaz+7v3xgmRQA+GbHSk3LNUTe5o1ervVeblKRdZaI7R
2SMxD3dipe0ypjIeuLd99jxkbK9UGmkPxMkLZ5IieJjkr/ed9RQ+MCN9sEUJ/IJv
Lm3cZJNX6lgwYFxhV0gHM6zjMi7ohEBNk8XkrogXbjq48NH0ADWg4H3dd2VGtT1D
2BWsk78ZoHd39RDBz5MEK4V/uTQZszw+K4sItC+iHEdE2NKl8t/Q3CsaoMxfkiVk
V+dBNSO9WWXI7x/krOA9aWBq/DJgxNsgUtJYiv6+IYbwbrpZri5aUvM3bNx7chVX
FStKF9X8KU7GQUI2h/d4YGiP3AjgU0ZKTl+hUlK/5hLjrjVYeBalo5sSfjrboAWg
ptMQwE4OkIWCLdzC1zvYj4GkWa9B8Ej3oguISEh0GFV1tRr53d+9qhm10F8STDyG
lIwNY4amaL9x7IhVPpCEzgmuzvHtcrqdBwfvslOD77vsfAMOlSEAO0TWqoV8PVdr
jJkYzxbSOPnEL4HH83y1v3Mqqx9g0IhywzKEf4mma362Ygd5kd255bp4fGFh6EpJ
9bhTexDhx8Q6w8baNLMHhcdcYJ8Ryt8laCc2mzyuB7xNXuqB9K8ZXZpMGhYacewA
LMOZY3wYGbLUsTik03fOQ/lwJsxZZbFZb+XOWJI9T+XTDIhU6bc3hsBHcHLO+vag
f1yhQwrRnXf48ZOX7VThW9vDsqTHNahzH76Nyio4cEa+6ulZKt55XEPBhHQ8ywSs
W7NqG21mNs2ymqDsF6GW3zVxrQiqdC/43r84eUOD5uMkT2yVEVgb4AQVQQ/q722f
gR9noy6J/U26OlTEMKgvNkBMa4P1b5lllaAxg8BWPZEfHJR5vhE+M3ij2HGcVsNq
MiCk6IKGguk42oOUzXcgWmtecR0JDs0q2UpI0M6heDJnDD5ViOax8DCCmBCfaQsW
zAPNBYzHMBY9qOVrhREDV6h6rcuiCxQktjSFHUbhU2hKndnPe9sLMDhx5CM8LfQc
51T4VXNykXz5tL0rBbbQvFAEjXrf9AKq7hcINtP7Jhg6PnlZPV4TCA0feXP95/+G
YqxzsyFmeTBiRCFNQBaD+mGiYIhkMOxYLKYFcCBDWU8LwMPgb68SGF9e6opvUqKy
jFQbc3FbF/3194dTQiouhlnsWPtP9tnGAI2pjziklqKfsh1drSFmEl87Zsu362AZ
arqTbdtLdWbOMiTOLRsa8MH03NoV3PkhVJaVRf23jno5wmxGXfZWxFnw7xz0FoJG
ZURdZYDKgA56iGDvXOBtSP1jnM933CXiYHPM4OCgVsfwrQi6qyAKp2s7CAZ9JlJj
rF2FB8IPKQmxo0X6GmFQC0g5nuq8h+PpSRSQvl3WDxaxj8kDxL8nqM0hnzY/uAwf
gxDde9vLBS5uxkq+qkEpSNpGTNZPGOB/eH7hmhjBY1km1WcwxDVcEDO/RYGUO2n8
jylKSK+Wb7Gq1hVNaeKUA5RU5sDxEYzo1gjFATTUR7nQeqGEOe24OtIx5hkiLbeB
iGxHH5FDItlE6TJ6oabdTfBznQiE6fPtcAYJVVYsoFoznHgjsQigIGfXm0OksDdu
F2LiPH1yIl+MqylfBzUWFnRDVsLDMAyQQyBVgePnNaUqluV5XXDtEXN20pf3KW8u
XWTi/eegcYSQWoxF8uYhVSbDYfljAyqJgy/lraTK71WPnlR3OmeBsg5uEjHtaO3r
Un4mz4yi8tJzXell1dBrYs9xvlej1ps5LAM8jmhdcktzc2P1Um4qeQoFWRI4cxn2
CHlpB60NKAT4H0/EgDKzHAVVSKVY52JsL9KfaI9FdmG8wK8XoS9St4j6tJ9uDnu2
WNsMaSG0Ee2XwcSQJvavm/U36GgKjrEFkUgl0E1nXZFAD4a4Lu+N2dKuL2ElMhkh
r6bbEdDolnY3bEn9syVHGnzKkpAklNMJXecdleXu46ARnwQZJsTTXfN/mlY24kHH
3/HVWvUd2A76pUHjdTmgvCJJrj0wg2cZLUktyau17yps6qWddR7h0ATVkaP2N/4b
qNYm4UcPfNDtj6T1O8lfCw/gomm80DY/nKspX8Y6OU6XY4p0r7YZdDvhjDL8xNXD
eiLQaLKL1TAHSxBLjZRnaAh34Zm8PWsy/AniLhKMQC4WlgoVWfPCPisKS1zkygig
NpS86gw4bXIA4yGbhbGDaJFODoqYNTqdaL/q1cqc1OcRp2VsdInWDVavSjFZ/tOG
FWDkhqMqLykSxiga8S49KUjeONK3vN8fC6uOcDHXRlENH9nBxqpz8wYWKuN45aGp
GY3vVMNJeueICevU8je996s31zopo+EEAdEUjdt+NbKDZ/bF/ikZh8ik/MW3ACmk
mg+hR+3yOfhsUGX5GGwdSwu37U6Tgk8RiM+m4TxFsF6hOMEmdfAfdPGEXHND2scB
1nfAGmslDtLBFzT9HEJh114emlzv9Qfc9njFFnYw5C4BTXAXMLx/pmoj/ReKJzie
NQtTgkee2kE2rSus/CG0UM0nOTKlxGLsNM8RjMAyqd1/2GGD8fZa824qDqzCHvGk
3mqdKHrMpEb1hhWDZB/hmj6cLP4Af9nAsLQezqzF4KgBYsZglufwlHIT4qQvy69e
7jSlRCkWH/DsjlA7Jiw3nLtKSAridu5vl/kflKMrIbCnb2T8XIsAYxA9jXcerh7+
4b8cvcATuHY9vEZo5x/2/Ky+T2inDzi6JkUM/hPdQUVSFgOMRVZ8185NwnBCkBKV
/Z4oSn8FnNKcsNlNMESDec0EOunMEWiqpGvB67h4kh6QL65dBu6otCDaNt5ftyqA
u08T6mxRy45rn3HGyVo2bFGfeBwpV+2KUm0cDIBUkTEprNBCsreTeWtNjZVtdW10
ywRYssIupygy5WuOCz5sdlp+Q7xA3fdLkCizmcyoOJuVGsbXBjE934CK6kVwSrSZ
vnnehH6MxfZ5e4GQL8YiSGVv49oUB+/fOhgcn30pZs23Y47AVluqqb4sL5Jf5fGT
0rEBkUgJ2LI/BLfx47i6PQr2nuXfxxFjzTrTRESYWT4hMpRb9eKimBpXQ42SMDNS
+CnVBjsocB6BOa+92vS07w12ERba5L50BH6MerAX2K5zHLsSKPBSg+Gp159NdM3W
ydCUe7BRgp4c2KJzjbuPLxz21/rCuLo8hOAOv8hMivC7ZVWEkIg0CDsTmmwwV12K
K9hjgvbhOBAUlB54oaqQ61BxpIo2ISJnVUqugHRosU/gkWVrLCR9rPWQFJMoITYR
ub67qakTJ8w2xigHBvvnBSEQmqO097odbfiK71bGOgjfnKBVHDuKOyP0O6WaNd+x
MFzKV4z5dDMctNay5eH70GW9jhT1mGLDvtJYvKUyADNq1EZ9YmFbQWnX8/gQADth
6bgsLbLfjq7qzsxEjhmE2BRocZXGd9kma7y6j2Z2qVuQlzp4OSSByAmpQg/1zuGw
X2he7bu4FhtVvm4VQbef4DhVuCAXFRqcEPAV2pmaF5vKhv2Hrl0V47NEbyXJNFc1
1LDCUEhoVYHdToODR36jIFYK/1snB4/FuTNM/txdnYP5zWmf7OkuIM3+rinnHPY6
L516Yc158SghLhcL99JsAs78omp6IWiRHrTLWCbTEMb7rHJkmgh2Vc62k+r07MiZ
a0dZ/JQEGlpfia1jCQ4NkFFKDQnToOYWiWqzGSd33XGZ7FL1nu1ieRw2X4XSjmim
OSx5hF7iVZl+AnqJRYaiGX7M3Y5UfBxCxkJB7yZwer3UtRoaFFZDd6v5PPxH51s6
znhBuieB2izqR1ZMsCbpi6kwZ8VRdD+V5RtKF9bPUveTAOxYTotmD4yFDqQElgbq
plGqHs2Y9TgxWCqw4eEoKd/T0P6y0ZfxTv0ysxVCuaPDEbYshTAWBg1W+khSd6Un
zO+27CyDZZ1HxQ7b8yyOs3z4uyqwhFJ+usVPyNpwqIsjufDiTNALio0BT/Sm3+/f
OT1HJKJwUqJVXT8N3rvvsndYLluo4aCN3jWhQpXy/bj9YxWZP0+5FefShgTr8emn
yyhvnKGkjwVPywrxX7fOBSoCF+MaOoplWb82KySUb837Y67r6TdYEwurbCgxsw6A
IJPn+NUgX0l8K6+Tzba/Q/qwjhOztPZ8KKZ+1qKFIBWoH0XPuwF74dbNe3MPg9k/
prp5mF0qSVsAA4hmGkgGEABk/EuF17G3kg2MMM76bS3Uhc6mx6OHKhBBeQecRw8D
VZUAT+d2AFc+IA/2vO3aJDp09NfElr8JOAGeNIG9Q27zbNvp2FsoO+/RFicHGIdk
VK0diz/K80xOgu18N6yrUEa/Bz+kfSRhINgx9ZHVnMefTY4rmsvprhpqPcFmN4lF
NT1PN6fwQNwFuCQkZtv4veEaNhgHlm0pxIx/wbz50bse6wki1ueiFD2vdajuOISm
qCtykrEUnK9lhK3ao822XJ4ESTcoQLjj/XcyuuOoskxSE/e7GWY5PLHGEMvM9Ae8
H4x2LEmr1kvUnoXq03cbbdPX6I3lEp6lV2BA6dFQSgQAr5ZDu0V1SMX9oMch4LZs
g+lNvmZ0OrtekSuCGapvqmMS5v3l1Z+OGPtXgPkUOiGUqqQBADR81ivQa8xO9vMK
e9gV74nNiyfXRPSJh50un1+POtkr312D88co0B9MoVFjp3YIQ4D1SscrKURBRx/2
XENO70bBYFNcxWvbMnAYgq/qXv53uQUZ2V7I0b5gvjOJQnHFYl8Y2Z6qR5NyEIIJ
JVheCf1XyOVA2/nQcDOIIGQ7qbyeopBoDY4jgQi670Qkcqqy0v8VFXFa1XZ6t3Ys
9gDfuJppgnLP0p7g7qzyXRcAVuRg0eIky9bF9y9uBySWSqtuISLDmfusQ+JqFE98
7gtGwCDJzj1XHVAU7oJvoaE62ucrU30PLHUucdg43dsb/Eju4WtF0N4NeItR8w65
f9j7xlv0Rj7ngQmkjvCqRxAo7t0SaHkRK9Cxx0hCzsPOHhAocNzEpfnNZ3/UjDhs
lX9OqnxJo0XUNxL8YEQ91eLTQZx24xOWYQRGuPezp3kVDw/B7E8roMSiIW8dFIIw
jk9B/ETQ5rUEyfEqODThwJd3sNZS+QTZ6y9YE9aqiVE6EfBT3w0MoNkxyOVu5Nxn
7w/dhAMM1W/4nXBQJrBPTc3DJy1kTvnABrhuy5ew2ZjLOWqF8F81opPzPZ/Ti6TC
q3Z9wR9PsqFIK7riL4WOJInAz+gomF4uzCvkIAGUEO4LGc52pLVAIdVkzdMIxpbg
KuHxMhg1wxWkMgap4NBm4ywJS5IZ6hQyq3ssXaYzoHEX7/GGM3dE8jUMv8/yG0i7
v6t3tVlPiThu10aEGyWtHsqMAiEJRp4oscOwa8NazqpOZuwfdyWvW81mX4ZkQRJH
AHyLuKfd0rcCWGXvMZBv9skX3lU68WZwHekbjnB/JEebJaqIKW7F5K2mwwNS28EV
OR7mLLakKo5996s0xDQAZHhH5VH4eQRoEWilWFOnKHdsdsc3zE+NdoU1Qd/BELzA
Sc0Ly8rYllkJ9nzayKxZlWLRMIJMZAIB2yE57evYrbdX4EaddF29zgx91FKdJynb
nmFl7rsekDgMd62z1zngFNE6DWw7JEi2ev/qmoTe2M4IjoD6025qeRRFh0AJGyKo
7j7a5Twg4it4yIcRt8lEXjs/BiXOIl7Wc7WG5pr4BWNIMPreDs/OvOi5jEhUH+pp
NIb8S0rYHPYBWnZH7Yq2ZonJzQreArq025J5hJGNtNcDJIT7KD5hOOVoQ5N1AnNk
6kz4wPtn2HKlleZHaNvixjP1KSVQkrSadzVmTlLe8PjD/Dk4gVMYDhjolUmmKR1W
ia5EZl23BPbsWgnFyXI+06jF8dLFwRnAv422onfvuucN0uWt/iSUE8SLyWLLspws
BU2ylcrKL8eflj6lSKsAE8Z18jzc3mQ/bOKLIgComjPgK0IjGrd8yB1FX1NktwfA
jC/86dVOGHyUI0D1wSzbbQMpqKKUsoVlyk/jR3qy2/4uvn9lHYtuMlZnz3W+zG5o
dg85n+DPLi6CYqXqCnos6ZujoBeEqnThBU4v9yZsV43Iszyn9qVmJ50govFeVjSb
rzxgUGxYt5vhVmBfAUeClmb4lx81WYD0OmVsCTV5c5pFXMlg/EnC3O3dDvv1H7Um
vwbs+8XC5Ppt3wDDAOCCR8oBztVmjNW5c8O2mfTww0x9suI4axmbBLQtVq1oyWEs
+Vqb3CcB6ViO+entetqE6wVcG6sMLS5zDkR4lI6Axb2DdMeFAPTqdR7vvQ2UGlV6
lpKlF31oCEL0FC/iCFPVvO4ukWhkd7Qu32xrOl6bsN8es7Pw8/Q9Dm+9Pz0+BRCA
zB5IDKyFAP8vsBlnBnSpOIz4PENCNFveLktgUFgcH80KQKWs+3/NLuS/ZsSFvMHR
Y+rAVMkO5UCxJ8DEZ6GwTuInkCDSrRJaGzSFVLU6FPNRqcTxz+YXkDYyXusf2snV
QAA0HIb2LzHiGaTd2AV14/NNvJ4j/O6rWwynGrE+SFSu+dbaH8pbY6PDQmeDx2HO
5jetCk6s1udS150SYYx+W0nZwwU7+A2QPUa8zksGy7/VrnvXALJqLSnsp+1uIzhK
/LcFiAluUO9E2/twntL9YHwTzUE1AbmybNNiaA4DYMxY90tB7Ar6Vn7tPWElQej2
Rv5AtpjxGJuHXWlyliqfXq6LnNDyZ5p7U/f7XBoNmZdnQ8GPM9iIXCZD6C78shdK
pg64RYjrOTrubej+PO+3jfU8MrMkWbXF5XM9svTjkfs7Cm6z9AOV6q0A2QoxEDgk
Ys9SdxvwYsbJe9KM3SxTZUCEbm5IbIYiqzAJD3TWO80YlxdPeFJCw2GuTIHQPD3E
WdHFWIO2kgbt5hrMSLn511LzcfhOpjXEWRbzUEgByunGzkV8rs+eSDmlo6JgiXYP
8DfqGixyfK2pzAUIqs0mPGtv44eXX4bxh+4qnBs+eZAyGJE+3QmNGGNdxIAAykWH
GsyobrF+LZoHJvwHhsZ+lFdocASKMDtFLw1kTjwFUKc1Dp9AvmXZEQ9yoc2Q5KaL
GOV+roitupJV1K/r+nuFJY7QxGdpm8UEf0RtaOOnsgRLdDOZvorndfg/ZTGoJM87
Ukbz6xuK5AOtbhkhBSGKEuR0j3tmPQI11x6xfzT0psPCSFLYpav7zIEXx7yJP7rq
rw/q4MHbvGpg2wAwjKbrrhZ3jhrZFLGcJjkZPLBEl2zgKNnlWPYPhR79N9PVEcTH
rLqI5ghqbcfbvAKD7OLon5eP5vU4nQQe268fvtjJd6604Fi0H8R0hSZ6SjhT5tqr
BP1cXNyhtS9qj26gK/M64LcB/STB8Dp3hVewb+f/R07QL4wOqrbcA3lRwhZPwCN6
EigHr0ouPeqLwDf60a/Y6hKnll413zrLC6Wv9+02y/ObWLbCX/7ujbQA0z/kzAe1
rNxNMgGssmAA7YXD4dFZvwNYqdN8Oi9NMW7XGCSjBHFrc75lByT0qFPr0FVqNNGh
E7U+t7OcJj7YuUqccC11pdmlTDhFyTi+vHNomn92zzOigSR6bkj4QJXo6uHs83oh
Se/PGAe8iBAIyJU0za3IJCmX/BUR7d/dlXsTHBvuNW5HdVUKUCPlq9GMtg7LfB7n
rUC77fa0O6QxOJjCiKjzLElwGRA+odW/JOtjGlLJuLIvFK53DRk0lvYcFExlEiTB
0MTGcjyHYiZJQgkF7jgExG/M05ug0XScvBjoKwGcCISPhVbRas+mMBXaY749TL44
cW59Cs4R62AOC6090Kn/4EdrBHMw/ExoqC0UDLdIanD3ZoD2kt+RlaKUe/030uAM
e2FbbIyy7fPtUOvV//m6cbqa+VTgvroYeRwoz/VZj07WwlaeIVwHwBplJX6Q6Wue
n5flwxa6ODI4Rb3r2BPOIPAFtWSIxV5XaS8onNBRQD4IDzph554EJh2EyR58iCPv
bkd0YLq7xOV5PKS5hHzUNNv8sm7aujUdNOarsnVE9kUC/lhzxddDFiy7XH3wOSjI
8Vf8rtaj90h86ARrXp0JFIGt9mk+KNE3yE/BbdKf3bv70ZsY4IGufmGz3MwoCp8J
j71k5zJoIHgLxAyV3ZJblSkxRF6OpRWunPuvnZnqNMwqIzQBCiJq0ztPZUdq8bgO
gIX+FnPBnT4nnbgk9UwpDODYnvYdeoWs3N1J2m7uYS+JqF5AlkSEw+4ekBmSHulQ
O4rkWWDBj+1SC0SsIpmPr49oMQlUnqsBQ9I/B/anZNFGO3QWlKdqfext3p99gYRz
czmMzfloUgIVdRWC/H6c3gxp5iLR4TBFj5SiGOmXKm7q58TsRxzwdrXvM5p9teUT
jm1Ub0mcYQ8dV7NPAjLXwrxtnx+blXUxzRg3N6NJmjqWOJLU62rujJHmINpxgoTN
MuZQWm+kv5gkmfipMRbOmIeS7I5rM753x059exnyH2h5UqrTMt/MHMOsiia7/14k
o9PDCw8awEWmS1gc0UV5J0HIcuQZG1g427WKoykmTHL1lCHjYG77LcX6L6k3+2ti
I7UeFcgFhBeoZaT6P9sdIEYdvl+1GFDh02MwwbdeByZ2m1pj3JegYIlcSEACJxa/
gpI1aZ2W3pJzpBV+emKc2197b7Lmg2zTcjFe88TaXyiWcPF2KQ588ldMoBrIZ4zt
QGM0s/eG544Iuv0n4f/9YKNvXZ3KAv1vHjAQmq5kJ6S9SFerAG6XdqoSL+5vF+8M
AnprqzVRICJJKDI8G9W74k5pS1eOEFs9g5vgEZcL82D8xoee/vtoga03sYvOO8Zu
HZDtz4E1LH8rb6Bciawcjl8D/FEhO3+dvZa7IF/tK4DyN/m25SelEUyPsLhL0RN2
NO6Jp2scsF8yjhM2ba/P+EG/UncLRisiiEABs+tnHru8nxRjgUoFYk9b1maye5nw
qCFkh5c9vWOvE+DSQnZQMaZAyP37LiEaRdMCnGW4myo2iNhBYahJGDMhLXLeKKHb
hPWkTRrGCw/H70icJPApDFRuGTNCxrKtDK3ePiqALPoTzrGeeaC7xb6qdimwTk+V
J69kpOwjnjBrOA5sgjS9947xAjOnQkbkmmYLrjwWSKxRwYDGnUxSBjoDn1j304kF
GwDTbRxl/f6qHcbAKaP5bbCPVPE87WupSipENiKtpaqCvFQWAY9itf7MdPco8muE
tM9dLii0bxZGEF6Okr9i4xXUbmOEgDGhKkYE5D0E0Y4m6p+lP/HkCnYmEFab3xzx
jqrxM3jHYabAVDaijtC3Xpy3P44XR7/SEiefM94G0y3TFuB/DNmyUyh6CNmkfWrB
IjBjUgfyz5uHF/mJUPESYYmd+wcX5h5QXmxmK0RcjOAGZ/X4wSGZwkBtMY2TGPF/
1Wi1sQQgSi6J+exM2kpHQ8Hj/NGoyFVZWd+TMDzJGtlNXiRXqOkiRxjcctMMSswg
oKozV94hv0bnHyxaY4VYTZno91jfzatyArXY5mIWan2BsE10eEyaNha1xFOQVlQf
Op1eVmbPPtQU3FWVkcFiBGMmmpjoNMsnIXmzTHDedw9NjGrd+VpD+RNC6AeBFOuk
zZ3LJaY0mExL6JnR6fIVlEfpVtAAmwVc8Ro91V2NzxLWZCK7OTlq6KRBrlslIgXt
Syelt0DnXwOyeeBwiTIh5tPiKtDzjjSf0fG2ztcfLiHsP/l4liYVSdkkE3761iGC
iQRcQCXRt3kT4bFbeway9YKjtUGd6EZTkTmSM8Z9Fa0/v4ZmRblQqxDxn2EcJ0/e
h7GOIKjVbq2uwahgx85bzcfZD4c2kJ1iWI4Tzvy8mjp0d2pyz29FRmVwsTd6mU2L
unod0cSQk7lojClL16IUv+XC2RNFEmp0804KN07xOTMGcJ5YXAtZDZagwJ4r4wnW
U1jrJQqXOhsR2Qgs7qIzc4+S5+r3X4SDMoqNVR3OM+cBtH9YCjUU2I3Rc89uWoqg
WPDjvrymkFrWNgvlE10UFb3wGaKGF8TXiy+vKvI+7i/Qsi9c2Sn9ZB1uLCmmmVwk
PnZrUNAW6Hj7rT1ZVcD3KNJOQL6RNsLiH0dvvP7T+kNW8p4F/hTSffK7ZX7S9y6H
ACg0mMIOwwoSw1ivKW/iRYd/waIjFLJTy4MnXWDVhVmTBG35JuV0FIN7Q4z3JaMD
KmxsNKwlu/J2agktfV5DkE2UPmfEpiozdKKjJvThs1FL/3fq8ReFM5W5eJlm2IUT
wMTKcxTVLjJfZWLEi3QZ9r2g/3GdZ9au3/RuP/kJzgJhDYbBVg0M5uUljrkVkORw
GnxW3Gkl1V8FrtBk0C/QdbJVooCHQY71+d8XpuZvfAm/0q7t98ni3Nw1AAqzd50x
pb0O+Y9kkuxA2oF5iepipslPM6pyOYedskScT4FnNn+C9E1BWMdeZhSDTt379Bot
65IfR8X7zKM1s5Mk1yG9uQgTLkxuhSOh9tt30osZ8J9rg+2pF8aDr8MKU9AbmUj0
PztsuJI5KGsREfbp1VEkMdTrDS7fU6K//LAkuUFgKcdTQ+/G93TpYnKS/4j5bKhs
czXVBs6QXnz2d1g4zyQMFUfdHCienadEGLJMEOZkmDZY16DyIR3imsesUQQeElFM
0eE/YqPFyubJNN4iYzpQXK1RDuH4H+DHvLS0q+M0aRswcwaM8PAW5L/29gNn44uF
q8Cwt/ZIL06CXd67fCa/E2vkSnaLgt4ugiCsJAMjRm8Hg77wD19DbBz6Q47+deJB
gb2PDtbQOU6UO1ETrs++425LFxhSS/QHmJB6BDEvwUUGllBoR9tG6LOeXC5UWYJG
3liUCSFnOhCzeque2x4Lhrvg+JCwgyuKH3FvFmrQ84qmBVXbpXoMyV970z2TBoso
0RHylqXwCSwSnHA5M5pkNnfZ8rELOL67zFYHnqfl3jIJNc2oUBDc4pr7zPA8c9sq
VC/qmS9HT6azK63mpym+OoMC3DHib2p1o4ManDiJwTUgZGIKBGjJET5fKxpqENwW
NOQTLWrZAbsoXmVt4L1iz5Ur/YrK88Qbgxky6DESBxPCc3Xm9FYVTUCZW/J+gPc7
i9yzDDlOSlaFymOgp+TXutc+XDshe+C+qxDCDCUNDI27dEoMcF3JcmLPCiLy9fsp
s9BgMPpA7xeNkkxbdg7VxZ6M5ueoGr5vZy4iruH2jR2uQXMh3ztaxuInQlNTcs0p
nb+Rf+1uG59HtiJb/aU1D8kV+ez4lVMlXplgCreuoc//2Jf+Vsz4oYD8bdo6Yovw
Ao14nalTWKxQmT86MNF1X+/vA4UZ3uq5tGNqLs71eDnsTsOY+R0mcfNjOPi9JGXb
C5PzNTBxkiJYY46E6rbb7c1TNeTQ9fADlEgSm5IM7varIlKwbB3klKWefFRsg+LE
d4hKGNYp3dMYH53igf1fdaiYXhz87LWBtafrZxRIOkhwIa/KhWyA5Cfyu1iqbJCU
LXK0pdZFg0wrJOWdf+DGr1s0w5l7zLKSFRwVdzqhLQGDic3pymO4uAD85z4Ef8hU
pctwDAm1rKYZest5HX1LL6Wz7UhehuJazUk7OLg1DFzb14oIWzWdLW+2VyuXw4tD
JzA9e87CofTDxBI4CYpMhoV95csLcBkFmcIjUpWwSXUevKkBU+prt8tM9DrFcVPb
CTD/XFzw8M5Bc6bMFHk3KJoRE0gX9uCIjq0fYtIGUZVxn+XajvLgU+ySowrWQD9Z
X+rlxZ5KAoovptr8+D+05J9SzOYnzzeLxL4aM74cuN6DwOGe2jcGDh8z9+KsmoV6
sWBWveM3XGxjneBPTBV96/s0JsahKn4f7h/SP4sVsJMvFAScL9r/+QV03Wf3ZpXe
/j12opoeMFC1w9AQrFipcNruddozUwj8Na5tOUIEtvs5qlud7TuW8iJ5WL0riqCP
xO+roTBnPQl0pzkkGCyocXL8TODgCoZiGq9jhDdTF2e9PQCuPqmWhRuyobeEYy6M
nmIJuCivHPv/ncbHEphjKTRbM/8ajcyLsaI8XRVYH5YwJ4HFfOZDij0WLEfU8X8u
CLniu/IiV5fIpFGLHF1KwNEtvg2IteqjNhWdN5E3vvz9vEGSpgtGzbcO+qy+Kli1
me0j9PK7NKM91jWwl1iRmRrhZ2kR3iud1j2TqRPvwXDI6WBHWmD4i9gcYi6Kh8xS
czVcqabNeHVvCt36NA6UQub8aA+MKXw1gZn7IJLHQe9t8jEdDELNHIwOL8fsp4S2
/gaDEnYsPi+XD0iPa2IROBwtxxt9ZpveKfYvhoreJUPfkAxlIyaOGsXU1CnmSQgp
JZKqaSP8xtlONFpR7HH0+YK5+saNpeu3JJ6QdUNpQdxPB+On58wOATJ6pvOLUBgx
k8dZ3XfBniGHtLGaR5ChlIt3/0X/Hm3FhF1T7DKUXVOguVKHi7XwwAhN3PeHy1/L
02tjSjZnmJixS/8hXSrrlVPNRUBVGBMB0PMbL4yAC+g2PShcH0OJaIr62cQveUbq
ErtbtBvQ9nIqWwflgQNhG57Od7p8twkByRbUWaZsK35bpzoBh/y9YLBPPeXMEOXE
LsowUnXOTu5fB8IVhXRwJkJQ8OM5LZ45/0v1s0ERvXO7ioCMVFfj8yAzmV4j/22x
HI7JfIVWZd4rbwMLqxL09p9QMmVNt6vucpqJ3cXQKNuqs1pRxNXRf9qQBo08303o
pKDgFKcsqoERG5GtK4KdUEyQ82TPLfaFV3PqEqfaXVLVegeS57h2V3gM6xFjfGrT
S8kNEqHKmSa1splc1E62W/b1UMI3HQlFfMnqcGxzFYYtw7ysV4JXtDGgEdko3i12
BzZSPoy4Mv+s+Dhpn/yBw1FteF+/px/7b4hWngRKT5h5/oOKBlnazFxSJ4k7tpG0
eq3Bem5Vl3gG4lWgYE/NXuCk1frU4SXhihJoNkhnnVphLo4YlaYDJCRIBwJAQm5i
ifCb6+i0RTgTFVhUTwKYRcNmat7jHDOvVcHHBjjjsj/0GguEOHKJO7+ArEvfUcvS
GGjxNVLBccQgsy3e7hTxynaYbepSK/FLcWAib+b0+y/lp6DIVIflxyJKn3rW8SWy
B8IKoizn6XLM15b3uycOfAoNWJ/ygkh5WORwc5FTW2TDWgsn+Kg0ew0yb8nVTRcb
denT6zwwW4MKn5e2VmqQLRYwIk0wOSRRANuAp9k+9xkMkZwshIYFzQl6H6Mkbkep
PVqPgPfL2t1MvFGKeKZNs0SuIBqRqrCZFrP1Xtlqj1mcU+wFEGu4SKwVfT7w/u+v
dZJqSGuFc2aUuKu1g5TTV5nJwoz1ooVuLkFIh+u7gCPuK5dGVt27t54y/oDpMq9f
YNv0wX8c6tOGl4O/8uEZPlUacr7ME72ms0ZUXU0yTHYiGrG0DQWvoxc2bzmbDmZ+
PLRZtbD7+LxI3WuxTHNRgzSLSdkjlxhJv53DtdNta3nWSZaIqW1HTWL/zkmM1UrU
uhN3n2Dhp8EEW/C14Z34nvVItpiw8uknCbGcErofAdIgrlghnJ8J0vleMkYEmoBr
k1LXBFSUqaLiiMVCAyt8G+Wl85QepYPkw5gz8wFpVOkSdQNYg7oQUN0bOhnwZHFx
cUsEz+LVN5WdA50NgGVZGqtLOT5yF1//RREcOlOLHnoun7lCBEmq45yaSOZypedC
+i3cBQDgJkg3F44mA2L6zUDCkRQ5MZswJ9FzlAIty2QpaIPPwYYWgD+2PiihG9y9
rFkrspJHgqPBEWml4Wy67wl0LIeiE5P9lmkVdpwAgikznJvCr31IQ/6u5rQcqinS
hz+qeuzBRIansSu7rGkFjM5HeaCANSRskWv++5lkGnfU2a+5mdGk4txwFCkCC5W6
gkhyR3rVoRmFd5NIiP+dfz5RJkt7EsPq495WwXW56HVfcputG8AHuEpNzO6wlt2M
p3GKlE0mUb5ro95svK/RQ8xYkyxykIettPFN1neXhZP7N/wYIF10L407rJzR3hVF
YlBdlThNrl7Ka96K7a5sjLNnBTebi08cGQjUBY1oFUA221Fek1PuTMWmqXwK8+7j
VA8rEpAp3lrBgtFvZpTm3qp+vm2LGPL/yytgCxhNDXqvF7/yVERQyphFxV/fE/dF
tCmTV7MVfeSC3eNDhi+JmLiQ2aFFWwf53YRd+s8URqHftDteoqcdjoAl0l1c/vzb
ouz8VGznqTSnpT+WGH+5U66/TAk13hGr9N8B3ryjMMOHoLvu05d2P6d0YN/y4x+N
Hkf6Y4DPH8oCJk89KJv4HmZrvEMz7lAPp9Z96LYeleWEb9o1Bi+t5FoWFmqga1Ve
Oqzf6eM1qHaAxN4FEyH6kU+G7itRQ3WyyswWUOUWFVJ2B4oNMMUL1s6yNuSUzVQ8
Bf1v3hGcnwoYPPUORMyL2tVmQN5y/m8D0LFr/Awui4GrOyL24jqjaL17ms9FRpTJ
bgaJQYvJgx524E5VjM2JALn1+nrtIXgeWRutItg/m+ZsZnD8koE8N0x80E6NmvZ3
UcT7C3mkId3m3BZ8teYeE9w3E8Eau01/SmxazJxgoTigex4959IxYFkMVi/FvVjI
BZngOt8I2aEMlB3QC2vpcmpRWNrPzD/l2nsxsGg2vuMUBnkXw46SgLA5M4YKmltu
CUwjyjZ6BVo8CpsGsSErzwj5wGp/XPYAxfl03+IffFPAoPnb7tUhG5hatMmEZhrb
WHlh5C4Pust3sL8jXTf+XvjsyVvyS6usAXZWImnjCfMW75HQbUDDUqrkblvooaQs
9d7iJsLfCO6Vl3jTQi2cubhgNM7lEdF+AH6etgNQqmE96OeklirvtjThfc/JHnzo
u/aFpCtMpgKPrEedKFY1ze+tVTxWXkQDDX700JVqL+zqdcdS5L+5RFgVhwLtQh+M
7zlZaB9MoGV+DnqYyjE+/8Qkug8iFqVMgSM/wmGJ7UCnt0S1v1PdBDrdoGJVD9kH
0rgs/bfKeUWYGK7ES1g7pGVDuMpod9U1dh9eKlH8aeOxjuSg6MIzK+z6qsLoi4Hg
ZyfKlKwyoordYKO7DCqt+Jy+ZvadguJYjo6OXE+ZBQe/iGOdeo0JsbIvhz63ZZ6B
lzyihY4dJdWt1jPa3wIsT1hMSvZKDlVSM5nsd3c/PbuR3ZuNUe+mVC30t3/lAHKz
3c4KphjOpTNRRwD427bfZy2v3kLonft4zYwpNoLKUcUyR2Ru3x5PO3ZCWyMurjdt
EFCv9Z8o3StOVy+5s7e2wYC1fpFFdEKqwR0uB0fh4TvejRRnoWN6vF9DEPvNTxlS
D2fCZr4ePn4W8TV+XT/UfJ91/FgZ7ftqh1M41+SWAjSyhvWj83qCAyH9iUunW8ob
XYObfo0nf5uYlkpdVO6S2WL/BY4AnGiPL5nQ11qcYfbLVcNvJXPZBvp+5yexhrXF
cfKxsZ9r7RYEZrcXXivIMDtlhgfsd3Wb7iMrbSxcj6ZoJPtP5PufWNJchY2j4DPf
fn3v6irGphWhI/WWhiy3c3jkkb0c/Z/AyWp34eIm2T3E284ywfGcFG6AfzJp+gIf
UU5RUOhv9U/JBuU951xk9Z+oZi32m60fsy51qe9/QYGqH1giNMyiDIMxICXfqOuv
jXLVqm1LZrE9WF5+7fOgFjoDU7vJVLIMDX/jKplqcN1xU6SUKacqVCWZxuhAhWJt
e8eStZN40MkGNXiQGWZuJ6RbBVtvVPKvfDvgDwNWQysSSWRDbFWjlfQx1c9PL5gA
Qdf+mEv/wUq58tbKPxNuiuMSAXytd86LSqGWIipSamGjxaaw7GHX23RO8iIi+9YA
nyaK5NSDbCtoxUbsh5Y4458GlK0RFmtPCpnMV46TkiLi+QTI2Y+WfVsVx+xGyyqw
GrtlXJfO7p2EBzmMz+juuWgglZ5ZH8tD6rMZzvvxNFJcCih6M3YyFjXumjyl8Eok
ZzSwo6zaQa9fr1ILEZ0p/Yx2l/mjGkpUp4WWU+UPekt/oWL0aMN+Wi1P60edU/ii
bpAqrjNOZ0Gqd2TPUcHNREblHM0ztGvo6BqVxZXftz2RTBeuW5u3+4h5NdblgQ7Q
GvjGAJ28dtIgHQhXjMWIXUbC3AltPhYfQNxh/OgJorye/7Mlm0RCcXVlV80sNTqo
Nz9+EtJwNcFc/AFoA/DRqmbqJ+ofqJ0D9eTAdBiNsX9fBFiMXElrNrvMQmhio2ND
FDEgMT23yHHTSKsC5qFlsBwRMIoJ7uRv+LAuNH2Z7kKICidyypvTbgZSyG4ZWI6e
0PAs4wZKscR+2x3U6F6zazbxMbNGskqvBUU/lVGJuCWNm+wyUlinQV3eNbUtWf7z
l99erQo0SW5knQwLmCw/V+hdR7c8h8Lntc2z+I6GYdidx+eKBIc1oe5UF/KAKDb0
cG9cmxz9cCRo9if2nQN7V56ZAjn4pH7BtVX3+rTw9o6WaXs2msZrTqECO3pJYf5r
185w8KC3qTRuydBvz/dof5yUTm8uXAxuVvXEg/yXU9bVfa7k5v2tBeaDlce6C7Xx
nSA5bUFsZl/ozE7mH9cWhBCJCRx0cZyyl2nCtLlxPmyx+PW5IK5V32OfDFMq+3VS
u+9H06Him5OPd+JNmgaDkVsMeENgpz25xsIBNCazkNud4b/Mxf4V+Df177m8WnjD
W+g/FNtnliuvnGIxpUn4Lqnl1BG0s54KMnx8/vwhy5qc25H9jezxbGii6zjlhTAC
igSBB9DDd5uTcyhkbQvj80g68veXl/m+hLYB6CPSC3OVPieaOr5RXEXHwrcGZwLa
uKznhnG/ohJLUMoWVdXMT3ufQoBumMmPVB07JMCeSVjW3NEuS8wwHbBsP6LCjiGp
rmyeTdkQGgKHLXtH43XH44Ki0x6CU+0dNqESic1k/B/JuKkjXVigYKeVFA28voYA
J9JWXXMcy5trP6P32kVRzvBRaz8oFJjfvwcLvPjpIJIHI7DBgLs6O6YbJWBt9EWl
5ZEHucFbTDeFuXO8xWVdjjTBPIQHm8MppNiRqnWkSVa+drL0+qugE70c4KXhtt/4
8nMYT6pIR8haoDrUiTFnK0La1naP6TuDkX+1JI3WQqnr0gxVe/EX+rnhg5Bx+2+C
WSaXsLrStyCSuSymAbor+y3qJCS1l5AXtqO0fZGCxlKItWLK0yE8Fu+5wSFb1jXn
1LtEFWmm4WWdRWWhTo9Wcp+bbLshSHGZN1LR/QGY+jX+9zDWVRcZCd84latZG1HY
3KMRJWeuA/jUvFATCWOPreE1aKK820dli43T+WGKnngXVQIanRfTkAPQTG3Wn4O6
+D7kVGkhNRKvlRwXu9KQWjUuW5uhUb14w+mqeBh0SLik4mTrBHM3qyBp43qXZmsZ
GYv/NNMxgMV5aIW6MiWIHneZ5SlUZn7wdAnyyRZY4RNGzxHFpLYWTZPHSn0saZWo
NKu/FlMqbVe4+yY0I9Gb7gN6o8DzqjdWW7adVpPk+ltmkT9po2Ct1JbegEDuHR5k
NgrZ5+J1GCfw61xQaSUjeTb4AmNn1eTLbrRXhddTwqWyQeVjFh9yB/6vcNuD9cZY
X2tL5XhiS5f77hJeOLa8PqaB1+n3zGuxhXELT5dVKRhfeN5tJJMseJ6JOtHi+gId
Lygu/ah+YQgOT5tYKoVYQpIp8ZYlHCVyiFzO+6PxHUShDJKq1zQvEcu45XTNfRpJ
SM75vhKQiS6d5TUI00rzdImjS0skAP2d/14q/Um+hZtumDmV0Y5gdZ90oEMGSx4M
7G6jATOdjT3QRSl+uWlYFj+7k0+YSuVpUykUfapZghsNFwK9T//wBJnjAwCbIV/z
MQnE/L+hwoZ+FWCf4IB/ckGrMU0b9xRe5HOigxJCpUSX2yoxiUd7PkMI7LdxSzQT
Sg0J2kobpa7cYmpGGhjx4+uHUQkaTAyzeFN5voLRS5a9TwFeFlP7QvVO2xTiEdzY
50Vn/Ar1oP4HxfETcZz41R+4cSA8xhFpgYgt6jU1Xvro0iNwjk6caeJSn3idtfom
Jrl/nXNssvjZnmRwdUWVHG4jGrAogRwoIPmfSkV8nKgiPbtegVymCfdkQ/2ofjpB
zU9+qsLpVDLRwqUR5KPNuh2RELUpEzSjwjSlNoHmcUTD7KIbN65cyFzRX9dWyWRI
mS8CWCuPJDjdaPgPXzBf7F9qoV461w6cUghD8Jjt4AWTyONJM3ZybjoLi1MI/Xsa
bJogHh9WaUSi1yNAlDqYRH929YkzdjUEBjv9mB51nRs2xwJ16ba4Lrt/i2uMj+Ro
oN/IY7BYRBVXFWG9IzfPn1/ScPfFY8k/KI6pgmBoEqKIXdubQ1lueWhvos9fP5n/
ZP8crDEm3OpRJ4R4fgVl7icqC9bR+lYVsoKG9hSTwBmryyGkYKah9VT8Kryp/pwC
fOjZU5BK4ciHP4YftwLmuKdnkBeMmIoHQGlCyQrlSMJWnc0B7iEunXe2Ttk2+7fd
TXSrmH59fAO6sGmyGLag8rmnYDTXVDz62p1WZq9he19yYuy9XnGenmLNIJruhujz
+xuKs4wJopAzn/sBxAv/A2ZcNXqr6abMyvL62A3BcSV0ALipHxLI8YDPr+BmKlmp
MrTwmSlAzfGBMVZcxXudDeAFK9m59EG6c2HeTz6s9HO339jhRjhXPv9kCsHDSEB+
XZ+qLo6imXoP3xHDn9cf905LzahncbZLey71eb7+xMLVA4qrRfP7n1es22438Agi
CHR2hP5Zx9xLehFzOGjX3axeoVum3/K+iiqTrecj9NZ6PptmSP+tTe5ootRuiBqZ
K/lK7nmuGY1fJfFtN/NlB6OWZIgEH3aHDxFtGdEmECeLRKuCxXmSm5+sjPxaqd3m
X2h8O3zNUflrhMkAGb9zdrGNVZ53Fv2f4exltSN5nheZPIxRNfVX+m8DmgdmExRk
EiVVaZnFJ32DkBYlwSJv493AibH1s3t9gFy3rrH2pJTKGtmGi3bYAWieH5+ud8/4
U9Q4C1/zkRITKZeRhRKTzK1HMQn1KSmJsHfUBge1jl7Pad/PBwLTtNurLwiscgYr
wZahTQx4JqG3/Poe6i1dNk6p/H6Lku7leai/ezI+H2EhPu8b17hsTgc1Tihxr4r/
2jRhN+raNJG38piUrTFWjlYILQVWDyn0m9ANUIOChw2GEQiRBS3PcmAO2zPag/xN
49Ptj7BxRtE7/AaeatdeEVAGXl9VjT5BYpsRGDo8A8LryHDODLxdZtqwtwJ+hHxp
kv9b0nhI8DmcjkNje957WaBOTtkU+us5nTJykUYb7KhTMgVHBRViaAumQai6Yz+z
0BXfuCTRudendLQmeBbUvqT6PzTRlVEjQGNRRCWpFnUk4jtbMRzxOmraGkTYpYz1
ZaVWZs5WSAPlgMiEbOJhX+atvGLC4niT97y3rqpBFfGSTLdLWS+gj31dy81MqBHM
SSXQP0B/rylgxz9yQOCYW1qQ4kE8YsLOulYAobOSNS/4tq2pwOpH+IvO+i5aWCPu
JjU2kl6sl/mtsojNU9GOKY+x+S4tvEQpYHCQgkqzmQhJ+Mb2gS8A2erg1rFGbwXH
4q8QS1ttARmdY/1p2ipx63L5R/tFOTGbQHy/gfHYqDsPDFFc2iFAG6qCCXktUQfl
eoiJXzIM1sd/lD5kasuwF/WsLOnbnPIObJzZH0lIBRTIQLO+fPxE0LqlQXRxDO63
TZXqqmhXKWAN4yamiyp4lXYECfFmjdYBXQyXDgjhf/7PIgLIDbLQfr9NyVedEc+e
hbzwS/DDn+0cSwTGNWDJoUU3YIf7TEuu6TAd9JGMBNXZ4xjEwa7F07M0IUwPgyeQ
2PR4W1sPMdXd+zbSNwEUQ3Cke64fSxs2R+ERhfSb3xiW1SvNGUleJGvK0v48YBQp
+uLU6MSUKDqGpO7fA/7bRPXG6V/2GE+k4yKmGTpDaZk19SPWMOx8RRwGHLc1Fa09
cUZZspNwH2jP1c5CKEd78JljaASbtGAZf1FFdIEShDZhQC0WZR32ybeR4amz0aBI
5XFhZX8OgYBtYfpLuB28tYC/N2Msgqf3Gp6uNv0Iqtbrwm7ZmEEDca/gt3RtqEhf
CEq46l+mdXNzf4u1quywaNTiuFvDsaEbz38JC2DrFwlWOmsJ0LFm5liMX4EPclqZ
wComg0qlHiZsmZfFVBGNoApmJ1DyHkWRdV2S8GoGTKJwD8GmiY4A2jzmyagB5f+N
1F3c6OU3eUWkKnK0EaK4E+lR+BgsFXnI1luXwlLjwXwF0+75qvzhz1AthAhfHuda
g1Gh5Petsb7dCjj8rxWYjWyllIvJ01XpUUIvtktyas/kJMbL0MEDUmoHbArfOysR
PCIIcMfLQgn2EnOuhUzJIjmY6RLRE+HmtJVBu8oURJcp3NESCqQ9d0bUXBaUHBmH
a3KgNVMghe05wPKV3exzyoeJ/+GWb+k9p/EuqxlzPKNG8/htwFwZMKc6B1YibD8V
PYLihp8NyPt3yT/mMy4GRqLsqVl8E4RSgt6CuERjGwq5Yc/BubtzlUtQibuINCxO
Eo3yx4uuzWkIN4LlnV6Ncp7Ktu0obPdTfb771yi9/m5kLJvzJ0OWZNyW7ViWMCxJ
YRGyhY9yXv37L9bSUDBTJwFWPJnOFPCf3CxMfbtp1XkS6CXvjU+fklLUEGkexRDD
G8lkiywBOkad+tr3g2HhJt1vK9U8w5fEaCyM3HJxaoSdnFtei5NgGoy44sYCJfGP
/7UkUwUA30bOW7jBuATdYgwHXdOTUbuwgm1YzOBvve0624NJHIbX96Qbi4tS5CTm
XubUTj9gUv2gJn06f6sln8MTWnLQBHP7Ke02nsY83smVK8TMl20gNSbLrbOjN1wH
p4baigzessSVLo8TbgcNw0M1sEPTrgz7/wvxi+gq7mL4aoottvisSUaSl6W6UwQo
lTL43sLIHhKtzEEfBvZcF7A3zGgMyv/jxzwsb0pEVeCn2nbSsE4V9YnAynEr7Apg
ETw/g1T9PLxUx9hICxptuFHyruuYAur6fJ3RXdifS/Dcwm9Y4j6Bn5Yg0kYPhBuc
6UFjjPa571SsDrGMuy1nJlEKd+rePDDLeBLYq8Rjo4Wjda+i0hsK/WzEWDDiXVP4
zc2rbeNVqN6NW/XIWj1U9jmHoQtUfqCzILl1oy3XT2/3Lsmm+ytBeQ7HttvKb7HD
w1aYM8SXUDv7ekmQQUL8CTduawKwA+TgMhRdmsSOZrcoU7/lN3/Kd+0zrjq9WarZ
bgTeOaE5hUtkQgd1SAV6EVPDNxfpfmSz4WfEBNuf4wqLyjiXAGTvOmbhsUX045w7
JkURKp6mbQ/GnVNYKY9RK29V1BEiMUmF0XCwTcE5G/kfbqpfQC/3V5UnCrIKXKv7
oxUNul1QT3suQt+Fy7rki7eRX7mOkQTBCu8fqNxEc3IBQArXcfpY9cP1837npESl
tlmDsbkt8c4EQbG/hxWngLeC5l+QSWiUyXQaONcJvnB+OQAxsKi/l7dVesWPwuJh
tg0NYxd3BqW0Hq/NHqVRwFoaQbSMNTJDDBPdxTF7wh0b82Uv74ZQs8IDgw3ZYsiR
IBHQ9Zkum7+MAbwOslzsCUFDVCjjTY8fbZWBqOa9EOgl8Wc2fbU426KYE9EF/1iX
YdjH6drgoVmNzWa8yELea1jp/HwwQe9KfiFnM0EG/5217M3oHaXlg9tMvr48knXs
2GvYg80W3Nwsw/kCnDiHGvWA/g750kNbm+LlOFMXG/YcuuQqYSyYOLyYr7It/chU
WquDLGpv1BaaB0xZI9O4vBv+ATL4fsU2SP438xex1SR1+1oHyIPsjr3mEPJ9mujl
Okv5yA0u0tqLiqRRN8pONIPYBgcUspc9i0yAs5I+jdvJiaQ80MNlOkQXSjBcvj80
W1xxLqmo/PJEz0ziCFdmPoqPn0himNkzSg/vDGnQZhzK2oOi1NZ/wX0qRMRsIpoi
T8kJHA/sQ9wcqr6ogIL9d06XLzEiGmZdGQipPCcywjFOzv6Vabkt6iZwNMQROeIV
nR3Na5R/fHPKV3jKb3Y8iWMvl6DWnMUgugjntz3C6AB4j1WADo8fO2xHpkV5Zzif
qxcNtR1x9CUHNRJiqK56NH7BD0D1ny51jR2xFDT+URYNpToXWiRVKmZfAEbb/T6l
nTb+N3VOL8a2afusKIEMyR1uWhoI81gSq24CO651q0HlAwm9dVhJF9jCqvxafSas
jznvDhffTVgrXD0CA0+FxkCJazfmOjsjmxydCNUiX4M77jaD69XFW14Ofu9DuoWT
fBY/7FL0oC1WOxWSUrkDhPNKNqCC54l/BeIi/XsnJQwE44lyZSmMXgXkMlnwz+hb
6t9bTdg6ata+mFqkJP1nrisJWsZRDbmPfa/3zfs6f5TW29vFg30+f1NRyTutJ9vK
LU0R/5YLVKCtzV4nCKdQ0TmqU7tY9bOP/fpXYUdzJkyiqZ8dhkvf5jBXlHMYnosP
t0bzqSJENl+qFFYe5VlsRSnla2+mMZdbbVJFpUEqxSd8FFjKab7n2QLF2+lmHglS
eZQvqv8wQ4Eu7g3xA0GesNRnzoOWv/z876tGbYbRimOb4BAWsx+7qy82QhVWz5uK
5qpbfBRwyLeXomgTzHsC1V2WvPw7DxGebFBm12AHWP2HadpoV5eKDoB/ut/b4WIz
cpq8gtWoVb85QVq2o16522bztaNjH6eeFZHvc56AdG579BE4XF0c+d16RePhJpfF
VEa61714EyWnPwNIUuyi53bmZAu06ht1PwQ2WtuxpzDZOw9JRdw3rwkEETJxTcLL
kaTJ+YAaTYguOUqYki15u6PhWE2280SuB1FW6lV6IpAR7y49w5yDPk+D4awEDpyE
YotV8cGQ2SLaayYVvwcVkqrQZYw/972bIVww3dAEAOkIZtI/jqCq19k0U9VdJfh3
RmAi4Q+uf3z37VT5uoWTIlUBe1K0gBJLKYJbLZKt5ahg9ZDXsxsx20bSTYSE66eX
UNw2PUU89awElcdu4MQ55dpyvyTLflfO6DDDpvV8ksW04uXQet4EciaieW1l2fZm
lrbvbDwuZfnp9BtAg8ZO+WOuoiWYHpFQqgppSwDHTAdh+aQbP3ryMikSlmvvuvno
BiaUhFRAXO2CDLd/AM97/J5jx8pid9ZZX+W6eemyb3mEejJWCqnFmHUSUrpzNcyp
TpZk8ynef1tQsAEq8EJEOFw6TJ4fVDsZHFQXa+eQJi0zLY+K3+CIPSXd6mvotlJ8
VV/msIy/vCBCTpJFiZBq9+hy9wRKYM7I6jZg3b6CYgAe9cRin7bdcxE6cf3UtaG8
oLIJrA0Lp4IPymvAruPW7o3jtTU19HK4HSZZwEHrLecsfjtZW5AXpBy7UKMOAgcR
/d94lUzNPoyeDBtvZLNV0Ihm9wj7BhYG4S7dgg2K8TsWBXVqejg09pOcXsgcPBGy
jQO8c+E1sZS8wIxAI8+X2M+Hs2HVkFHDlCRz1f6pD/cvbgHMou6DKSpWY3TQl/Fa
e/LIhUIbjshJzHSkaqv4ex5zknPm+6dWHGFj80LjvEwWGLssCUU3+Ryj68T9zYFl
WVmZOtCVWGPYG5VanC51CdcM2gXqNncnrRLpyafCm1NjyaSNK5kD7vjavY/Hi400
buR1+FSQUvp9zpqnB3UXwaIOdAe/jUXgd9Nio9jcy/dXN5p9TJiaRIQAXWUQQ/zy
byt+iqSGrBUpDUF41+PvofLLavMx32rLdSXkZH/5JDpznLNpa/fsIgSwW5hRL7l/
Y9eU/pbzmoVDmrYJeshYq7NlsKsw/2Kw3fmpGJbFKuuY6BKoToWBAN8luKdfTugN
qFwGb6KMoqK38nK5Nc8LFBdpqgjmjtXAQ2U1FlOZ3G3WmAuYV7pDV4jR5ep0FVKn
UHAzjDOuv9AFGxtrhe8EivIpnSr1RWFtMOYP4X9r5a17AtltbV/rF/Ny7OW7DsC4
UgRj56XApwWCb/qv/Q+siDeh75WC10jXB7JMiUcXx2kKcCl3iGqbx5OVoDyTdcSI
EuuKqlMUoqoqc6CYW60zCiUenLuDpGln0TZwvMUBCt0qeCvWjQuJLsmY/BN5DavP
bQvP/RNt7ztl9HtSQDMehZCBCAMDxN6wkznBdXimi/7jz2LiVVt22nRRVfEAamDE
lIGP9YFI3HG+MinE0ClkOg43AwQtb6k3psD4ER0Qf8cACeC36zPnu/xMpW5bbq9q
eHkcR2Fy65mpmLS4ZIfe18jxamSkVaGq+KNSUqiCUDm09IRtSACngnYPXo+CPuMZ
LwK4+FaD52jUWg7sqLrjCibAh0ZwnA3SOX0m2cTwJmnBfnt5bNnHolo5GFW5MjiZ
wE2ETUW1hQg1Ab465TRZVsMdBYp6oNca/fnYQawUBiKt0xfLCZDnfIwPTvHB6WsI
bcEEV/CUy6GuvwykhnaZMA8c9193H8diy8Uyp92y3kMnJ92abpJ52nqHVBuOeXVm
8A7xbzn9uWHB73k42jUAgLNvkrNyOcg2hVoBQ8cVK36rLHMDG45LST8DKkWns2OO
kuxGI0IrerP5qy3Qv+uOUkfNMFRuVazQEYdXifn733QIN5IlCsMuL9/Josuv4IeB
jZMyLO7hIjcVEX14PssOpfJDjheWDdquVCT69D82kXH54mH46bPD379WmA+zyOeB
wYtXzVheh8M53XoiFMneTothPpBfTSbhdPLh3QD5UTLMkUfItd2+AXF3bh5fGs3c
0kNdKi84eoDZi+bvfU1VmJg3b7jBaEfoMBJlxsPx3XFMRyVSOLhYNjOHo2+MgC01
xBh4Tn9FqaqkBv+e8AmAPMm6tUCNUPltP6xgZz194x7d+4N8cRMhzihhwJflNnrH
4QEFVE0zaJq6qkw37l5d0MX78NzEYB9md5GnLmp/h9+LmUFB9Ylnuv8CX0LofB05
zWR9Qbes1IS4wSX5pYWQrbjQXzRcjNYMoGMblhq1zYTIROqsp06ixwqwUfw2Uflr
gciWykGOjFnHE1SIzSG3wrdv8WoM8vo8mI0FZ2tdh7jSr0YJw2hkykxmAr5DRBmt
z/jEPvTp2123UJBtXZW0CpwbHPzrUu6G30FzZJtztFFL27iKugaPKHdWq1ojW/qo
MFomsAwxvJF6WBWi6Mo8Dl8rjeLcD4gKjfWuokalUxJfWqg9daGgR8EHX6XLlLUS
fjKxiqvgWC/GiHMd99N856BRI7xXWf1AOSBSeI7jBSVhczLlvyo+16BMecpcvCOV
bIUsUK3DpDoq8ZKG+GU8MzuIB6KaZre6YvmBPobiGnonhABEYtWSQm+OH0w5WOY2
16Byil0kPIOWRyysZ5pMxBSHfFbDxxDw6F7Sc1kfqoLZ7xkn0QQ5lEmJE1eCsK6y
X9uhCC0OuH6/OpvWnKagr4yGgO9SdaJKOU7/Wum5un0ETTO2YmbSS/GR/qC16tYb
ljRiKoYTjXWSv+Oqlu0NUc58GBvyaSMYc0jdgWKTsDsn+qwgunPZx585oflFjygz
JaS9gW09NzH91TXMdG364rhMVwLx5poKAvpmJXCtMAMyp50Vsop4mZr4LL+hQ8Rs
JXXx33yLE2E/MLFEhU8q7YS6nMoGWQv9RnSvNt1Z5XzxUTcLiaLD1cd72Ps55soL
+EYssoG33ZKqcMLIJMqqrRk+NSvCKUJnV6Ts/zqo4bRSI0xThLVHAf/YLIz8+2uw
/wpLUXHEt0af9DCHcoqHGxEp0VWX98HoOfYhru/UT38WqFlBz7sA4309GrG3nPhw
yOb0TgqRwqRo/eoRSjtynpTr5zHqYZuMiJ1zTKcZ78o+ygQrqzkFwuk5pqASgRCb
3MeKtzz+8O+itE/HZ6p7RZRtDMlKZjJiBNI7j0/GXKnBzeb23EoqXER0H6TGTUGC
mpSzr25Z64bqRW5crHwfvd2V1CeFXbVfDbtLl41yvbX7A2yt+S1QScP5fLRsoBV/
XdaOcac/PxF1VweUMWg1yPwgqdUMBQNUYtpsPKiWNDSd0n51K27eFoag0rWbbHFZ
ETfTfah0v0ES8oRjbIN9SDMuESjaCfWck8+SZtmPfaRVo4iK8k5hgNGBfqEjYeco
/lOQKLFkY9fuRJ0q03soOsFM3V1GmcLav3vbeGP0JFWB/APQF80V7kTdppBBd4wf
Z5xDk8J/WyAl2dr3+OaR0LQY0ptO/eqFG9tpmRP7LZeuSV3hNOFUYDXuzFwjOx6W
xtLpzc5G6GXXhRc9uuQ4hwEkXDLkOYyHJEzf9QY7aNKXpUmd+iY6y8DDpWaiCPtQ
vg1obfSEIDBwsH+D37QXrk6xG/oP5svudfjL2ns3tJLKzqpDevdPD6W0TsVldmcZ
I9x0K8X1jFm+RACqeEXyMPgVtWpuNJc4awd8s/aqjA1TAf2oYAVX1fMoN1vBVzth
7T0l8UIu709b1DIwlY4vQSh99BsktNKz/I3D5x3E5cXgI9TlGrc5pLIVsbX1p34D
p6kVFPknu9cvWoc2gAlMfVupE8TZlq0bgcebte0QkFHGCx1o0XgRCWaee4b1HWDd
0ctn6GeQwApKAxZLuB5Oqumbh/5uyrsZ/UuKxWCaN8knC+93HO+FHhv+VaeWGI+x
8bS0BNnfkvoWptBg74u2Qcrvx/Ht6UfUsDLaBt1fg7eCkMxkdcRxQPTpnBnJC5FK
LguI4BdE6+sp67ygNWbttp5pytQ2KqE+mW4B7zuMw06S35DgzWmbCKaGCuxYwQdx
r1l0Y9iumDEkI93TBOMjRo3kkB0qfcP75tylt7hjPCXLWbf1AS+As0UBnFQPXEj9
pjhFCNuljL/XcWlNpl9HL4g4cHOq6Dhh2NOWK5P/iMXClr7HgrDUW3Y9F2CI++d5
v3HDZg19kE3XcgwDwV+mCCkxuHrpEaQWXJxUd7KuhqcIpvQEKANGce/tXuBO6IQi
DSM5B5IKuONUdjknXyva5GpZVcOuoKxfIELUn1yZIzNs/7VIYrIQrUAdGGuJOyk/
aekdvtp0g9lM3QALiewg1PJ6uyeh1SkVcKNAM71GzONAl2T/GINsPEv4WFSK1xzz
vIB7JOtui/B3P17HsaFsXCrHauJI5NmpPpPVAXvNVZ+JwnJTUOnouipOl56Rcdl9
uZ3z15/b+dfQsIREKlHPyOcHJQclj+X3GcQrClGLrkL9DAyKZTOU1JlYlJYMVei4
LkPn+VxHwW7rQ4gvQVX1W1qENt7sTQmwwN3vPm45qrX4HFhspFoXt74gTxr5QKu8
uCP5QOaxVkWEJa6Y2rVXeA+dQv/JZlyFoKaSyEMFn3+L3E7A3fogjmDUhb9lzE+1
Me2zrOq20ZGM4pIQUN84xJ0Nyv7F6WAli0PosTiHVIoBYKytH70icjW4dkUNld0v
mrfoTjnE/ggG8IFS6t3vMvrWl2kcwcLV0zT+SyrfMrlaXOx7evQa6PwXr9wrH02D
ogeIGk3g0HpSvk6X6IBVboa8dzU2d+sBMZG6EFpfu24SQ4Xj2fxGN1GhzTCoDacN
uaNxYe+CiR5iRWZiPR4VTSInUaZAijpfhmBcOgW0I531Dx+qdgF09vI4o/EMGwZb
ADb2ZgIRY+Vr0B5xG2cirJrPhy8EHLnVEK/54Vprs+6PqxpQ97MQ/Xjj+ygzQ/e5
Z+mIU+TYHtOpooo5waR5DTNsj/WwUUK6MadFCK5Li/RjjgkaeYfXupy394nJnqQL
Iqcg1yqGR36vHdnj+SJkhkRU4HE7vEudTtRU6t0hCRIlSw2VcnpCQkHnKwTVaykm
dnPT6IoV8T0hg10kZku1kjvQ6yUCk3W8dfgjS/+yBUh6Jl13bOtQdmZPqAGuOCcu
Uabe2CSICP6hPpXKZXqw+HVp5GmDqT7bho2LtQA4cOMrNmTdd2qtjAcIIE1VDAWe
95imO8iKtY74yQ/Bs2isGDedQpxds6fivQeZE4Zoa/i61hK3/297w2hUV6rq37Sl
L8LF7r577VqCl8/zdcWeOsT72s1XFfSNabZ5jGkgBlNJ2J4HuYG+3IG9p+hA6hWz
gxyA6iZgsUyrRsdDKqTWPGtjGRw7AYmhGHab4lVLbp3sVG3VXy0A2RUT1h89zl/s
aaRPJkOrLO0bk5BKhCu1HOZaAoCJhNiEkf2hpS/kofZLCCUVrS4s0xmlxyi0lZaa
9EoaUZViUOX5yzVNV1mEj2EsCIJoFy1nTTr0uPgNbFOLwR/1pMa8gvDoSPSfHb6P
lv3K0Bc/FhZf4vntNzB+99vmZEmzYUyXrLXOv8rxTikJlY0vmM/kYL386woIlwsO
rr1vIdgKluT0lw5Ai3IFV+XmH9VVNZjTcpOe8pJw/5uBxZu9yhZiF+JdVS0dLKh8
cKayJbflvOkIm4UEX4a2CShXknxRonba4v+YcjfpwQxrImS/RYxhKut5u6xysPEx
71uz/EmzoJmQ9gAPHHSKrZa7e0rnCxte1llvEIVn3Vs9wO5hwEuVJuFYenvx1Uzk
2EGGZBXXA8B++x//dxoYsdz5rcZW9O4DjQtWG8ZGfKf1F6JdB2HfCnqXmgikWvue
/JMNOzBRHG7zf7zDMwle796COnoy/a94xm0FCnw7jIaupFMWccBmcBF7vzWrAiBH
geNWlQ6jWFPXxcA22Uyz3lxt+T084DUuyjI2WTCCqWqsPZ/L7NFUI+byWyq87Lsb
7qQHwg4LtAugH/X3KFxlon1i45L6ebQ6WttgYIL0C4KB0Amsg+IuVsIvivRyeA3m
FxREUwwfJ+MGCITJVhEpq2eO9IKS4MyAGRkPdrtwNRYM8ghj0S5lIgVuseuHSrmh
ARkIRBYzvPXHSEQGPCg0Xulhd10ei+DQyu5vKMyky6QtmNxu4888K5FtCllDyXKH
tFFY2mFmhpDgwZQbRrH5z6sQj6ERJyDrtzUrHHRf8WKVm2tULiajd7ddd2DVEq49
YJJR9CTJ4sx3bP4/T4nL21chKTENmWvQUpPTkCzpiNloeweIgd4nLAoBMI2ishdQ
1HryBWRMc8CpPYfYb/MZpWzDpmWEaKVFbsiZe1bLn5r3KXnrvIM/lRWkSYlhymFz
bCsQoWKhMGMsT51OC73LomLSfPLhlu3s/D8whO2H4PcbqTD7ZGEq+B4brK2HZsK2
nriFAkHtfELP2KlOaV6I5C6XHVgjsJuLFiHUJ+UyR8OWsaYc1hKMIIwJX1pXyp9I
c0JwcXFp8kaeTNvXv6ERp+SbwevS9c3QL2HVVXjdA+4FHCYGj/1nrowUuIPX2HKM
Hy7O5EgB1y/iUwAQCF5iLKLxGqYpBzg/4XTtZDmNiNuHThUvokoFcoFsABLX97fP
+ZZm/iiUqvVV0bYlwGUgmPlo+WETer0zKh7DxWhfI9x86uBVPHo6Znime3q9blV2
Gt5fqM3Eg0fPH3wucEalJHJwIIMd1kyYs2xeYKKuwZzsAd0MkMr48Jdbj3cKesXQ
+2/mooBZsx5BWskcqwOKfXpz1SoWJuvFEB3sEKFNNdaeLZ1JyV4wi58EQuSom7fy
gXicSv937n5F5nkn9NrEBZyD613WZtDAm75PDfL4YLEsst877mOHJypndBKBP/Ow
nY+EwuX+lhmqa7uCv2eaRq7NOaePDPPKuJ0Frb89LRcunxTVPfklWZFr08K2oaDG
uhH7dAOzpJeNVuvX/6qJjk6jpyCgQbPx3dco/YHl6dYEv4zbOEguJ5pz4+e2+jGw
297dLyL9wq+z+S+ilp25q8YiklNLAeSYE6ZmdDbow1BX6xvX75XhI0DxnuD0wQQg
Cy96pQtLPAsgjWiD2dUfMk96yqqrq683tbwQ+4DAV2ScdClvXzvdx/vwlXowHk68
ovtsy01FUNpRGtNEuHI1lVx0UhsiwbefkoMYEszacl2c6RVymsMhprDczGRFBqE8
QBgxsHgPbMzdh9G/9FeF6Ms/rDd+FDylSifp0D05VbzOmvTBFLScnGXP07Z2LUhv
Soo1siGlHIg6uzXREZQlNUKOhWmcxZ4oQ6dmsHrUNmKffmkIALGIu5gOMjvk4riq
cSEP6Vi5MhhRTdEUhtbR6/dYzlzcX0ugSaDH8geKpmm0KqZxTOauAw4GBJtX+Ozl
OGYO8+YxThtfbgunHpe6Bjhj2aeB1H3Vz2ryFDm7kDxZg+43CQx9hE7nWOs4kN/s
buLkcOWC09Z9Muhcp55trIOWbDNS1ilW1mZJEZ0S8pu9rJzOL6mBQsX9V2tA1yhy
rUKNLq+Mm1n2YbqzKFnqyffAXOkzdHv/M2GDS/wvDYwreuQeQ1o0yjIss48PvHD4
1XX37WK6P2Mnl4sRiM8WBVbgxfdVsL9pNPiYCQd+eQEoKvn7o6UIBy8uBA+lXdZn
XjaSSBB5Lck4KVfiSvpnkhWjoZAcHX8g/I/fL6s4E7AdaukIxcWL3GRFvsdIdQq6
7XqkeMxSPpEncf2nlhE1StT/Ik/odam+qt99F/6NXCqJw4L8LrJNyzv0ykwWATBV
H/H61KM1WWWG4779/jd2FGp5mJj8d7bax+s05wuWNTBnfTKCuWdm5mnyYxuxBDo/
SX43dY61Fe9JdV/9i6uoKqg/cK/X0Kxi/kgFufDR8zMYVu8TuaFjMe2ktdZ/kJIa
8cpVJUmgGnrlkPY3nxxvIrIHyNiqblrmtIxmqv+od7jQKRmRi/7s9xNLkL5zLb2G
kXPmgODUEWEO5TDn+gp4ukayNCimiAUpOJA8GS/UD9wQyTcYtbLDHGLJfQH2tKmh
Ik/21vUWUrT8Jre1l279UaOQxoBkozjPBXJTRQ/6HQpA4sOP6WV7CXjdVXVwQ6OA
zHFJ3gCrnRtyeHNbZLpwMCEh9iLEzWOUx3ByI/ifeGAZK6kOUPMBxr94muVP26cQ
oBGDZdwoWZKxct5FpoPgrm/XnXPCDKDE5q3ANojwsCZP/N+vqb9aJHtgnuK2ecXx
tSv2WNMlqb7axwNzp3qUFFbOZebgcCq5vMxRG6SCwlwnnnmCdh+jcCYkm9G1is7j
kVDeAQFcJr+KD+0mO4v9BK1tex6OvoQzUAPLGjI4YlDE0KgLetQv3KxWqqpk6BA2
64yO0BvqCE9bdx+qChHFmX4BI93PvLzNBL2Lked7a5hOtR7tAyzDUmR9bnEj5H+X
vLyVmtG6CvQEpfZRzXV6Wy1YSdHf1BNDfmOC9ZJr3uefC+yOV6RedD7dyWn7PHAz
BDF/EKbLcC81mY1WW63onR+cDqPkW32ba0sKshwpiRqBjetTxsqpTwtX+iGjBiFn
O5twJCpdjm3C0nBIhWde4Dei7ddEyzz9aNrTJEWkwvImNBSXjvST5WEW9Kbwhfca
P+40SkP53kRmsbZFGdu3Cz+koNMWc8l+D0UyEYJh4/FNxnjOSduZaIDA5qwmwfUj
QomiBzTTtdG0/tmmNj1ymcsFQAZtstn64hUsBMx7C2FmZUh+ZeUXrK8wipFSFWTE
/Z9qZF1S7/9mDciY8In+TW/JT199kI4pJG/9z6prQqVy7kgHRDbV1TLsGZy9PP2e
F9+rmoumT9HPFXto+u8MHn/0QRoj4sLvz9P5fKnODg5sHbbjSDHdvhMEwmwJJ2QJ
npgPHUq+05yw81iccL77NqjnC+aCw16e9bZ5zR//rZrXtvIrxbau0Vo/Nx3KHC2R
32kZLQP/pl1SAOfjNlukvq8vWLfNlDK7tT+GF9ZLOSO36ygTValvYythgM3/KHok
8YHO88vEq35XCwP/Ht60VpKXLVqKFXQPPN/Qg4qyBMVQZmudpRyO8wYYUxrlG0aR
YT0NT7grEcpoSEoDR7NZnfXqf57IlXXUPUErTuYmeO8XNmwGobi+Argur+oqR1mo
GyAqQw4uo6gZCJz8khrkgsAE69DS6dfXPayIUo8BqHV9LL60+SWsIHQE03JNSoXV
YY3gmFo07rKJvP7f/BD+aMCCvuQOgFy0fD3nUC6jwlxTLgUtS+UlvEZrLUfm2m04
5+4K3rgS9TpqinrlwPAPcyCoiCRQj4p3HRIaNm3Xl7cAOx4QnBpg6PlrAmQphdNG
8SHdI0Qizg7fJV5v0z6cvWNQP8PJA/fM6zTyesjKPl86EnPPUV5APPAkM7u0vWKz
jeJ8Ue7uGUv3b3BVfDAb7uEvABKzchLOVak9mxwdPLqbmEvIjW/+2Vsu7Xiofpcu
8xtktsR7/5qdaMo4C8V58Mm5JSx7TQHnAHu2uoFYVoGpi8Ak/mVXjqodBSRPnUuY
G3xaqUJt0Rr2bNMLIU1gZUQDXbr7vU7yOCqRdFaFKPAaDpKA9cYj6xOPSiCsnYU0
CIG5vhqzWMwVGQYEwW4YcImfpAzC6+ySEH6ddqzAsLBsiO7jbVsPDi0w9h6OxJC4
eMMO6cIVTvsrC3G61ML7cM7R3Rh+FcsOBW5KHozttNHeKfGTjvhrRkJuBgOjnz97
RN1sCki3f2NBYlTojLuN2Y76ifGTbm5BmNpkAYkeOJcx7nKtGKsvSRq7J8XhqGfK
QNeZMQhTovGpStuKf6a73BuDWO8LnUfx+y+/JeoKc06/ldMWZM3NQLd+LH5KUrEN
i6NAfRwPOWVRFw7O7P39QtoC/U4J9mdC+Br+CxaIE/t5FuqL8elJs4EcFszu3Rlz
OcrtrOYYi6q3tMKASDjhcSgmQbX9+mjpwYGLEL0F0+TdHJIqNWSP6Qh98xFpbVa7
v70X4lOVdyVN8qiA0W8oBUy5Fps3mdcCg6zTQzp6l65hrszBNFz5rdkYdPJJ+0rD
rPK1ZiGi58hDycXip1pHLY2lM3R6r0Q7FR+7iiNL9CrQGDEBloSKBGfq9HLoZjhB
nH+A0szvgrBQ/tIrk0PMYDMAT6gYPvAXFgTkPHYssLiRQg1rTSomV18cUoRHBXlv
tpQ3K+PCnUTD/Kgb3nouBE5ocIH1rJK/GH/8O8+0FE+Jhh3f/jdBpBEhFGTTVEBy
CFZV+SON2NIkdIVJTKoZGwSRT3U5f2u9p3LnkLJwtShJih6AsT0hVQrd27R+gj35
QvP9P9wZQfy9u1lSWG/LmRz3rNa0/VIRee0RTiLf4oECX6wD78qD22Gt9/M0zCKV
eb/FpE5kLe+peoyJ5fMcyX9lb8aPfcZbIW1u04+KtG47K+UczhYpwWrbJmLUpJTK
oqQ3vnhlS25t7w0B3JO6ciQC8abwJrQ32Kgx9HyqLt6p61mqc7BhNnAGX4uQcfhS
psqAznbsxeg3UH9iPQC9QlhJwbIor1lH2IN/RrR0fAKR0Q4Py2A+qz3JTmLgBCwD
j5/xPh7mMUB+h0SfWGX+B1Ep6EHdVSwSU3LiYMjNt4wwUWm8ZpXHoz9hR+VB8cgg
iRe7siFSDGvx5NtMGGxrmFSxhGMCBleU7AVFRdmPJxyN+30YwcX3j+Y8vsXK9Mzb
c8bqRcx3ivr3wzUyrQ4iZ4agnPtls6F+ZPYmwtNkOHDa9TbA3m9pVFHbKhfWdLSF
GUUawYbh8gkSHXmsG5Rz7aM6QxJHtI8bHPljC1eelrj4gtZAU1w4Pr45DPT6qIjq
NO4h5ejMIlCUBskpu+e2VKnvsK9EfENWK8YqmuDGoEnl74ZrocDRR5Lf5208iC1a
BeCGBNRsz0l+B/SpuR4RKqHcQgBYdET0K+El5mLE81P356tN2zYWd40VNOGrJ1Dv
CVh3eK6BAVqNu0laLwNeL864FOtYhJyHzvf5npZGTmn7gFuOrzP2m7MeF8LO1jty
wYL0eT+VEypbab+BfWglhmywxw83BLB2oViHXU7fcMoGnDWBWZn5lYy0TWIAqQMI
qU6Leu7ZQ0itXm/NbsUz9pc3ulhzIw7PO8KOA90UxUESOiKMZQmFa9NvvE6cXAV0
TgEn1+kG40FxK170YZN8eDcw+mC5J5uzp0XZH6/yW6/13jzZyR61YEdtqE1awzek
07iOcf1H2wmeCUiWcTTBPti8qWwEYx8PExpp/e4iWy38m6OIFQ7FwMDyGUOOKavD
rWRGHM9JpUs3uHsUbUIT7Sv1GNq3i6H6ssRONKjMg7xiMZ4VWKjK5HEqgkvcjrDJ
o0gnI/ZWQ47Jn5VQKMJ4drsRRybLVguzCJIRJOfAn512NWHLXZQoa+lHWLCnh/aY
E94/+vzgC9kv7A699ewnFzP+NCiwLjxPoVmyJmZ4zhddMBAaplsZ+aRHb3B4dqG4
AVt/61SrHdGDCB6pyc1jwuobOrfmQH5faH37szDSWuPs50Z4D8inR0tQibQTrTuA
W+T82GJ5+7P95272mEQYO7fZ9swyJ2sU2eioP+o8StZKPyF67RZ6gCwnQtxubx9X
CxANBWcSiV2iwi6rMRSIuKpwSm15v35IHVuPQdYcQ+AnnYZ6CTgwlK+tLu5LKDZh
nylu9saVFISKgK0mZLB27jiNUycCLX6L9pBFJ4Yc5mMLYqB/7WZskUEM1OuTFeoo
DsLfQpfz70OG7ZwmH038NYA/5BP1zTd/ByqPG5ioflqYpnja/0Lo5e8Y6tqGLpSj
rywDXoogVNLLHLoppyJCKjFMRkM7xsbIsj4k37uyCsm6qLaEK63wBqwn0m+emfVl
SJ1i+Azfn+0OXrl4JkBNczyIjaEgfS/DO8yMgRmYIL9zGUWourDopagg+hmg/Hdk
fNA5SmdRjOYCeEX3sNmJM+iRUSTWvMpYg5aQ6Apv4QuR7tYBXrGJUa/n7UjcLEwL
86s23G1SDMEzIJhS8eU5lSp3QeYvmG/NLsOw3Mh4Bn5wlcDlX8tSwj7U4QVXIM7z
gYjoQiHmvK26WqOTimunWXlDbalARRuuV1VnGXmmZThPt3Fxz1GQPVt31BHQ6CNd
yITyiT5psM3tfztf1AiJ2rVshYoIyzqqkxtMbkAAXNduCPZc48cej6801RM8QBoS
4cBT7ZUyN6nzhuo0Dw8nBjPCX/LaUuW1x15726R8RnXI4j6QSTbtnRqVKPcoheYx
7fzzsLHAHskZrYQztFtJVaAL/qcvVFX4cV3uP0ZS09h7njO3ObB2VskcybnkmVVG
q5kfUuPshGyFwsTWrlpCSE+XZgkULBMygkZi+txgVEHji3U7mogbYGUn1jsQ6Lpm
OOAtUV1Llk1vvBB+fWqVJ4ZfU0BldchFFGAraPr6Kl/xbvlT8phZhVJ25uykH5qm
NYGtguiEgpZ1tATfzIKr3Qvm4wjy4sETTQHLX7KxvsGuEtzvje+TIPf0g30/sPsm
HnTf1TFxcreB9b9cgMMiG3d1nBy0sYPnASyJT4/GKfnTQoPvNE8TNXt06RCN9veL
279yjy2sY5JmyR/aZ1McaI9V6u2Bo1e5+BTo8RKINFJWPxVapmLpQ164daHzL8bx
n3FAQL/Zj+OhnZAph/0+h0wPZtts53EjtXd96CkZZE6L3MqlL+HPG9sEmJs8kZCH
ZX9hoAJxTsvkBoyKr4pKaNWGGzlMviqv5+kQqmYO32RZvyIk3JcqE2T5IJ7RAltu
fL+XfCxbonI4NF2MPQfvbsn+xpjOZJyfuuAvH4dsqL4JtZv9359IU3+ooxemNz8K
d5YBc5pZkC+qKXHIPXVLT0POioOANU98kPTLHYc5T8tA9UcEHHd1ZxyoMGQ1hk7+
iLwy0hdMVfWzhWMuGfo5kR1aKT0IB/seyeOSQBo6RF00SIVjpsuRDscJGfvzEIBW
7wdalfrfxNGVs9tTeO16GhnLMD043y2X3CAvGjcU7l3cAODi/Z6sWIFNOlVqaT3f
WsvZiD1pS1dbJgxIxlGcOD5prITaGHUIkvWDVtHuGLTI1JK4UmwZ8eEc6GvWe53z
MzhBjBuO7Hy1tmhml43q10yKxx84VN4sBDgJJpKO39zqUrOOO7hlzRUsDgiUA6Tj
gEX617LmMUhfBKJSU8F11RkCmwGO+sBMumR5gUj//MSFVc/5XvUVtjM/MOCL51BJ
jaS3W6wNDoTjFauf57DMJd6CpfaPygBa+YljWhgx4YeyQUgAIutHpiyNkM/gceX0
Tcjpmlp4Nk83cTtya2JjibP16jnIT9uuZuWolJ09IoCGJy3y3X266LpoRJsJzjRx
zqFe7ZZ/2QxeEnxvCWypG1pwNlvdq/Li7TaY2HgPod58++SvhNPs06pi7DL2iFqp
h6eAkWAP2sIBD1oP2Ky45Y1O5dwF93mXj/6IbVQ6pH/uVkPK01WwapOziY7qT+n7
ZTPLEgDHIlxdWCItO+QvtuIjrcbHEIxyViiwyNEWvNskDUj6dB7yK8129F5zgqfO
tRg7VaU2W4l8o1tKMwFunYgnxOAhLb8jKPpebLXEH4VCyZqeM1Tc/NaG0UdPZDu+
8B1EvUBeHmbFmeN5jzMz/loNS5ry1kumKmRWbwLvaRG6AYXEAglYRAITjEbTWS3s
RNjisoZyfF/yU6fwSVLTyfr9cNg2tkh2gQwC6YqfnrI8oqNbOShQJ9GUuyr3WEyX
kZ3Ob6LzU6k1DZiTYxjGTpNfMNKUQIvEpwyoVtpzHC8uOKoUMxlvbrKXg/lexL/P
BECcXsLBjO/nu8NV5XSQibiWW8wbOlfB208IRw2Y+rfodgkJep/LYOd9aTN4nHtL
gWGZK3MZtFvYke/F2Z0NwjJHKzOTskXmvuLGhkZ0/bTEnOdUk8EFuEnBJ8Z3voRL
WKMTn+7T+T6OFE8RICI0/QFH+lxoqiqMJvBTsgIqMs8HirujU1oab9HhqA0XW45l
Ihqbh5xZJFFogsc07Z0QZK2uoY3L/KD+I8RQMu/WdgDxMZuj+L2myS/qxFzh47mn
aeeyOvoAJGwJ6lIfAQjWi3XZjUZgIXZapc0MayY56DtPXhoFwwoNL2VxtX5oxDUR
2ErDeC24BNShvF0b02q8ETDzhL35Ar/Hiec2uizoJXe0sQx1i6o+ST8KF7zzs79C
v0XBrmrocbz3jt+cGPpvFu8n8x0KVghCowRX6ppELQWnmQKIiUIkxa0e8PvhCXMh
9t7gITE7asYTrykGKsFfMJcVridpqO67idd11OlpQ6TrJpd0QzuHB00uY2RMfgNm
3efF/+WnkeI6ZVGoXGk5UY7KLRXx14nbvJJ3nMd9vOWfOcelKfxcgbVpvyU6Yiv8
jV3LQf9hcjaCxMl/mPPL4oBTLMOg0KFD6IQy8rXq7I68oYDUge4Fx1aNhPE+Oh6+
fzj2jGmsHDF5X69EahOpNg7+rshCE2xNXjaIuaxF/ZnhbDQ6FfsgWWgaiF1APkwo
CfOoPPYwb6kAe78Mj5mIycfsfd9xVwZXUleWDiYWYknZgB7ArdJijwD2kAimN5yW
GZFb+Mp3MTX4eiZD9fpiJJ4Ouq4Q1e+FL4gp8tX6MLKw9ADlFDhOSjdcVk5w3nsp
blIXTMYtcRgsSIwN7YAcwQYcowNvUlDBKg3amuY53IoNYIL+oh8GwyWIPKTLBRGE
u2K31z3omIJl7voQMM215rV7E5cf/OpHMxr9HDFwNMNrkjiAb2SB8nUFsIWQex+A
2wHfOeIyqh+gM5ZRuCczUbUp3oTYagrTAbuNPb94O05yMna5L7RXKqVJDwYGB8Cg
rkp7y2b9cku0rZ729TGn3QeTfgUxL50o3vy15Un+QplmFEcSfiMka2BsfamtpDAY
wfvxlY4J1Mo4N3Ckcwv3a53Sh35iB5k+gAC/au3aeZiUsbCwHLPw1MowiEz3kVh9
2WvZQAzkQEHDmycpATe0ydyTU0nkkPl9KDP2Lnk8BBfvT5bi/S52lvQpf/2cMhPe
ROFzsa7RwowTzYXPQizGxasPIT+zpmuCXIOaEUJl4n8f5oQyNn7kqSNtXUJKyjRL
y0DlHemh+IVVbyIRF7CC/6BK3fWqU1oeeNEaXXN7H3lHy85HAUZ/+ZxhhVqcq6Jl
Xzgj0hS1PT5d8HuR9jcVhGc+1l2OmHDvohQPQ1Ak4PPO3PgPi9Ha18ECndRkfWlH
f/Df7KXzh3xucX5uTddqbfo/ZUxTtUwwmYyLFumc570E5qMRS9zrMvb2BcH1o6bB
aLTMEZG2RRPsE7zhq7L9CaXjKCZJaN2rNc//ffy8vf0H9SskNDKA2qnuDIt/dP52
g5kgZvMV+vg42tQtCPM5KHQDWkQvJV/rMlzUl0jwanBC+ucPOuIY5bJk7bAyVT6V
+kwcU0vBOB0z0D/uMT285sYP6Es1MRtg2nhvC7fRhBAFGRSCRa5KEBPQSVrCEeuw
+O3HuveJULbJegaP7DesU8hZp/lvtTkAilG2fQDk9i7ljY8Ue3/B+SAnUyAr/FGY
jNpBqYdcxk9YUSFqbxWl55gSqM+gMsO8hlLcrQozE5P5biBEWb5TWYClMd99Xpv4
CinZ1QhPEmFWKP1GOaKDwBhrTyeDSx696Tb83E25wb2r5h50aCNazPqTWl7PQwET
TTYemVWHe41honLJ+ovPTzrTei5J5Qi7ZaZV3kqaYwcgrgrMOu4ar+7Nb6Ii2B8Q
+LbWqYbTtFeGmSL8H5T6qaMbJqVEoiTViUSPE26ca4SpT3a79qoZCcj6ll6A7iJJ
G88wkh/23rwoyM8qMh3fPIfptlnOvN/MrKljoVwZlSFvrXvzMl4agf+pYlvVXdyq
3VgvApXJyKCEPESufIFcYIpyyl1RsXrIPtms1U62rA/GTlugZ7MYVfSNA+wShl66
NLEQrRqW7q/7AhrRuCB37CZomp78JW33BIByeqA4Kcu0XrAYmvIXeunOSMslhOFW
8TSvh1EBUw/n5A29yV9q+ebwfPpuzRThel9TQ9QnSTbaiq5LivBwOLV0YTbMcxfk
HMWJNWMEE2ErTHB+ya2ohGGtdpchJFWnIGaSXSgJHCAsFncdYeWBYY9DuQJom+Gv
OS257iObERCMfDIO5j4MhHXAvernCslm44Unei+RGkVSRtV8r7OLVUcACEjwcgyz
iApKnibMVTaccLAOP87EMC/lDyz9br+Z+x9unC0PpPHuFkmXPTK84/oAtXZGo6El
hHl5AXdjTAW4cWpHdUG5XLR1Kefi470wotqLWVp5kLrVECBrftuhVCFje4yvG3g5
sbLaq1VjS9RI1JosA/+6sFMlf5+CJFZ1g5a9Atc6yzIUE6e8XZJSaNHIr39Zi05P
amTISJG933QIcOl0g44/TlMFZIQehQcroK2iDg3+LC0eDPDWEpqSVnTT3MPrR3Ix
x9fX6pks4fmddE+U4XzUYnaKEdpGATAPfvOtrhsAjwEZrLUFFa1GtjhTwfGQj65F
QHSJ8RdQxUiQR8OogvO/6rvrMcdqroaHMUwoiR5iD2g02G+GtwOuoEN7CK7l8ICw
dNBLDOyyWViNtTclCKJajSncZT2VixDcVySdFV4V342m9+7Km1V+Ze8D6ntdse+m
eLJJdRGWC2l7goUTdhUH59yFaCw/30K1LOkU62tu1D40zI0DG/MRY3JDLSNGb1pV
OjpWva60lEmKRYZ/5UHIeb+BbrFwy+GPtQf16Da748HQQ/UMFpD8zWG73SVTFU9D
As71uqNxS+i9avmaiXN3t39gz1kn6adVUX5LukneBwdLiIHDfoDPGhbZhQDeAb5Y
uIqdACKvN/J9Mp4oTMp5q1y18RJjjgMP52MmRhWj5aVR2ocbxuotcPs2h7MWve3s
mBEdNav1RlLE0PqjXZNhQ0+otMu+ifladL2eLbaqhUZBpCjbev8SGuMYuUrHNY/a
U3aYmMZrw+DAJbDmmj+vf89G7/efIHAIzK/NTqIGsX8BvMy5p/yYbX5ItgEkY+7l
Y10PxEb/7q9sYPTF2vDZVs9ePifNAdVavDayxbvZutweXcaQWAdmQjpJMU6SciZf
RkjUj/WWmc+GSr2F0ClWDY4dJEFZvo2fisc5daxp5x7V8NHgfPxvLPdNpTvRI+6Z
N08YCmQvJq8xiKJOFs3AkX7OCs7Ya6EDbatk6kRwbFVQJaCQrvRnpkG7I/2hybDQ
YzW7owl417lpiuSnWsMkhM8fyUfFk/LZdOXZoyWYeDv6aHrgdgYGBT7apu6908+H
G7ue3noPrkmXu8IbwZjNYGuf4UoPI8mbY1oW0+XK6+TPKyUPLO34sDqlLGNXw07J
dn4DX/JG9U/NwHMsLHJJ9CNlkD/WAl+lZq/3zv4RORZLKwej9+VAvi5dwyGyJyJI
begQXSVm/3ym/2v+okf2z94TUyIjlrs7dwHIsLX/WSiQxDwx7stWezuvjsiKBda5
WEpZJ+W7c8+rpyP8E/PPVWIMsDxVzHjTVE/H7LWrr3Xkg7Aepd9PyykHD+ebZLB7
ueqvwJ6hYFizdxGdSB4yGu7Fto3W1LfuLpImFueqLggXlFOCe2sOF+NO0DZz3j1H
QSm8qZbDGpUYv0UV7Lw8FharYGCrFmAwepAT1y1FHH9DhRjKCslCa/qLavyWDm84
dEVHZU/3cbMRdrOBH6uhuTyY7SUWpw8DfiT3ci3x/DylqDIXyzmtSUrS8kbegj5+
rp1HrM5naC/XJW5FKIwb7xYUA//8V1I8xd+XwiL0Gi4RhgJvb3SJdyKMDBaPqGwa
NaZiHzQp3Mb5fZek0ABxcjNs8t3F3SuQJ5NBBywPyH12lQt9idw5o1pJH/PzttGL
je8yypcOgfwJNd+PLmIprZ/LXELhmzNKAKPa/oExoefsB+Nm7DiW7mooSW6X8Z1P
gzA83WepJv9P0T9c+JAm00Z8AW36rRkdNrY2XI+JgwrN8PlnWY1UBV2JI9vr6j6w
lbHK+NxmAnovoFmV7k5mmXr2qktoRI9Snp+f7EMO/FIGOnwBbRaG7L9h58fMTpkv
PEV9pW+SXVqTHr6qkuBzZwhO6jcpIFCt8cx7wJ4q/KAzMRs6vWfMv5DH7GfJ2M96
11O/Fq2HEDiAqXQjds+0rLNPCa2osw0ezxN7wKkIM7sQSAK7hmGA8KWPud4x/cYQ
qKkcgOCNg5stHvCaLTDHb9+K2mYFQJHd3XG9+yYZ/92rndXTh+J6g3zVa74xhR33
GwKwkHiA09XSMDl3vAGq8PwEoDe8EGWxDMRHSbszmJpKG7hA4ykTWPLXmX3bO/Nq
PvkVeH5DVfxOekpHiQIY9bfIJZ6JfL0SB3E+6pReOHnYnQjhgvLVPg5wvGdceqZD
b3GcDwpr2TwsNZECVL5gCyT2fcO6BhxMm+5YIoS76Yk2zPGIn/1pWUXFUqtG9lE9
e67EyxPo4rqvI9AZjymn2KM9ljBKy0nZ9rjUEA0AXEPNWqYUJuFWIXW+utV7TJn6
d+XVcwmuT8UQosOL5Q0kPEwwtqur4LT/jYjHZiw1tmNKJqKS7GhIKftFufpS8T2A
Ml9EJKn/xSZI5oRjWLgOirZm2iWxZYIBj/JFlvsXrqXPFyb+zwNu9/iLVoJqsUu0
uq8q4mOvieRXUWAMt38LLClhEBIdaFCT32Ocht1nhzw/sf46djzG5/6QRN7vg9Sj
I13vitE1bS5MVZ4otOerhhR8GYuVNjoQSZKN+jkYiYZ4jdFVUi1yhBZaeTXDI4G/
0QF7P9lTuBMpkbFBXUage6etXGNatY6IZwa4x9VpOdwo7bSjUtdU75kGUsR7AYMJ
JSn0peEndo3eQ2R4RwUx2sQrxiQp5iXyGta7RZ6DX08AuU81a0b0ag9RHIMwYFny
BEmeNi0ji/cj70nCDwTAB89mkI/ONG0prbVloR8edFFsNkPLOPgKNtFjGCmP40bG
JrKK9C2f5N06ItV3DAae8D0gnkps+MIGKdEqYBHfpi2PzsbU0PfVJmGwLtypNeUf
sYqUpIV0ukD4xoHJ+fJmnBPgQ+en9ia5GSCsdoaM/XPbhdttMs8ZRfXeui/C1sFY
qDXmagwnuj2uO7Q5iEQYBtSxTJ7zWzetVF6hhuSDS+y9dH1WMHk0mRtCQL2v/EnE
NAFw7qLXMSVmpDRCvkhvb5Y3moHHl4QVUUb23AwLzqw0b7rneeQtCUjpTJvU0bcM
BZeEDo/b+1cPw99vTcBRtTlViHpkC+QbYORurMSNOaYyzgpdiQRzviv/Ocw3M1tF
A9S7H1s3n6cZX056upncWO/Xw0ZCT/D+mqJ+McO+qdvJiJ19aVt4x5v/hu/d6BMK
+X/E9Z61mM2SoITP6VRKLTYCu8/FtmLFIuPMnhs7l5OeHy6QeL1vHuEWdLFw7rcz
ZivwI0YE23Qv8VFGELJcgCYNtf69YVJ+dnmMIaQJEnBoIIjgRT3l9bXd6ERNpkHJ
p8mKAr2H6wo8j1DhrkE4Rp5AfAi8PnkinIh5/TxdCSpdid2uVIFNgVzC0kuJCOeB
GxHIrkKjZfnaRgXXZmwQiaqL+nkTJxKMlUBGErADWPRFBkfI0SNjLQf6blMx6TqY
lB1LxPqZ993a7/Ke9+YXCNUcW7aSmipuIpLFFO1IZIkedeI35Vhlp/Kl8gWEINi/
28JiCfYhCa2lak7v/jvPCEnVJCzbwHAlwyMuU1O4/TjlhAyOZjGtgjS38YMaXnPV
bn6fIlzh8FaVyVAhNfeWq2ENiSYQiItyBnSiLlG303wwXngVPOQ/VdhZuqZr6Adx
4nG6GVaVm2xAvDPWvyWxbfU6xAeCuci9zYma/r/gYUFywRQOIdBh4DpHNvExRuRX
GwD/EDt7BNalBCcfCmF/kQFaSFzhhNbU4TvkuJo7rUg6ZP5lz5bjZ6cXeR8wDmtn
Ua7WoT1BS0dFrz85mGEOsxJEX5eKNOlFJsVAZqzD9D1ZnDqVS7hUgd9wh1i/kGVS
brZqoMntUdrZOZejYXGwwe7RiloxBs2pBEHgG+w/P0j1eBSHVxzAT880HbeAqFCR
E2VsCHzvIk28kkG9ck7aZaQxzvgmPy52cApkbsYuIDICGMtNsu/gtJ4kEFjYoHpu
5KSkPisNma2qlXtfw7euAMqQfbvLktghwsJB/a3pNxcvtn9utpL8PDcE3CghFP8W
q64JlrhBMLZf3NvK2Tdrxx9p84DjD434q+RxtHQ7dyCRua4uYeC5C/m8pbmzV3Yg
2s6YBzBB/eexFXYEOB3OtTUxG11d/XoOLW1AEQY2U7rr2Zm7gK1R6JT/KgjkjlYw
cWO78frD206QAiOt2gOhcLpSr/3DxSvkMC2bS1/RULL2jkYZ/xFo8lJSNCXuEb0U
6Hn80GF1jWf4Zj8vBToN6Zrdd5D9AYNhSCWMEu4AqMx9/qtq8TjDk5fS7qKMJ1Qi
UsQPP31zmPJCTTVS+5Sm350Bof9FLOXOGLyRteW0OMse7ZO3AccWU2iJwTE+MOYs
dWg4dP6v1Hz/T42iWJRuriYbYwQ62jFzsbjUAEFWwwWMTmbDfyuBioi6V8kOXMS/
jUewT5VX3vx/bc9nOqL6F+YYrMYFDw5YaQVkaIZveGNya77qzwl8ZKOe7JrB+GCh
qEDzhmMs5bxeHa3a5f1NDElOntLpeTjtwP89Hr27mvxKToWc91JJRmmgKIGGMAQH
kqQFRhk4EoWsgfdx+5h0gjPbfSs9zzDXYXOVSmU4KCO1qR3P6vrWJp/oqVV+j8Md
bJ8FgvL77EcpT/V8b7VN/vzchqmCqOEGd1qXSwyO9Z3TTYjZw9AsDYOSygCFWY5x
dBo0EhFuOiVuTscJkYg3qwpHMl01l1K0wlLSWxz95K4+YDmPlXWzA0CWugadcu7h
IXQxkO8Am9HxpRFTpjfioc3xgsL4yan3BBXMbAdLmBvahy68ozD5/7cXT+LFoMmD
EXG8VDeYlAdwZlQ/PIfjO4fgf39doDEe4PTjy2yQ8/5+ixkg/nyuDVKOTSL7TvW+
AFKhiIPs9yMMJC/6zs87AiZNMdHQIltscKs+eQPiw+2FFdFi5GQgMaZDPrMQHXVs
xQcRrvSURGsJRH8oihfCVsWHiSHh553sMIiGdiMtWRamXPyZ3rF2URAzRgmJhB+j
L4iNoX3TEvCTO0z8qmSmmALy/+cVp058FLjgIAwK+VpAM3eglrgy8EN54XdpJSo+
TPnmYD0vREbR3aVx2DTdoucUjALqeDzacvsxFE3uXs1YzzRO3Gcf/royATerZsby
wz2Kfn8OKurToFUCSqyUQs9C7DyJLl6vpbeE/eEZTu3dp1qrKqEl3t3Nvhd5edkE
f0CMfvhPNrj4htQPOdqBB738ZXQ2xm567UFj0kHhn2jq2smKTBw3JI++epCASqWT
0bb3SqgOa2nGcMNgXbZzdihBDUyBNdanmBDGnzZgErzwfI3W0IHteYGLfqDG29iD
aLTGuHQm4wbJMlm0Sln9qaAj0+UtiZTw653CqRtLcTHN0q/Oo57pSrSUWoCvvzUP
+DoguMH4dtI3/dWP+WN2xn9kT0DihffTuKtT9Qocb4+4kABEL79IK9p1OTULS4Un
ILSJpkidhzOo7z0Aa5NkK1ETqJLlFhuSaYkVbrbspSAkqR5DUsjr9nBpXA0ztErd
DcC7Ku51UuOS3+eDrEh2d5yb46C0D0ayaf/hXfppu5jXhIATpHLnTlvb5aJbZ+NM
WwXKMFl4vqwOvHndPBSIAL/C5kqipD4xIA5TTVivNcAJMKpcTBv2GYr+yqz7XE1w
cfFJ4+d4Qb6439vrTZ8JjBZE0Ha9Mvh/J7bj8eOAPe79uEJibF0xn19z1gIClzkg
resTvNWYHJGIVl+1F8NBbRPJP6Mnytwm+j9ps6G/0Yw/R+yKfIw1eUndIh8WjOis
K/yVuEdFDGhg+2FIpNXkZIzJwmHLUNuKMcWx5aNJfSbjOt/+z598Bh5DcP5iZxTS
CRCSuKwXW3d1HncGW+eIyIR4CwOY2FOjuyyIlgfYoEqCvRkIWPj4BcPa624Bxjgg
fbkeQRLuREg/dvFW273L8ftGJ0oWJPUUaIPUQbSOvFr0E06dr4u3sqGe/3pBJCLX
wfcllGknvoQ0mceztHA17uDUdDX1RrP91ZmpagYxjHWKs1PnvBe+MeVRBOOZ3oWU
ns+0icnPwzZYTrhAz5yg/eDyjLhK4kTE4HdARJnwm2KaQpNL6tYEI7+E2ALQVHry
IVHcJn3HUOs8c5CEjVr5uhg7pDwXkeLW/f+Lu5ProAOQNTGFy4hKbzp1er0/mAO8
n2BBKv4oSbw+jbFDAmFB3ZS4njjuTOTv/JygBAmLmk2JOjfbZd5Fi7vHgw2Pk4gK
RtMmsJiq66f6ngTRDQhkplm3ns+j8o6No+OZc/GbTJKQkApwikay4LPtUt6AoyrP
6Ow9FTGA0lOL9NHR8/2zk7afrOW4fI3XJXPJW0YcxyNclJDcRQaSRPAJuC1LSY23
slDt2QArENsgmUh3IHr5II+TCHLQixTzxaL2pC6/T5VtAT2nMEi+zdtvuA1bc4tx
AoyMtFb7Rza+es+nYRBJXIgIvT50IVIo/pAFvVAjVoy/iYfOqsSkK2Rt1pW0rMny
IYyRKYT1/6b8kIU6qvHyH6MYOUSGWaCtcY8kbS29yUIt9ZlILP+f1Ze72Xp+EyNz
QD1Y/dnCifbALKuSnCkdIYshS1a5UdqTYU1467EZt3mtD7ZsoYyrnXrqhjhrdZOo
J/00xcFYsiK1d8RL17pAUIhJ9QmkVZQ6QCxfvENTagzJoR4igDf9nJdtHeJh2R8w
0nMFQx9yaXCRmjWdHi0aGckPImaycXlyKLqljx6+udL8uXJda06b46yu2tHauoE+
mHfyWNfZVnHub4/rNG0OSAHk/DG1mzET/SRap5n0sifT/mWmw7ErHvf0YFijV08z
Kqc4briE6EcPFbfXcqY9oE/0L3RIxNSKb/6GP+VQ8q9kqogEAbiZPCQbl8vHSM0o
bWP1hr6q5j/mzyXSLvhsiFsfiLDPF/IJQPa4UCqGJa/nTmnwkkuzNNz8l0B6h4xa
teT/4j275Z2qopmfMUOtyEut2pb4SjHWXTY85i12w4UvZ1EWqWs1YYkcB31eenAq
ySqCe599CgJZWgenCpMSVFr0nKMKkpUO80u8mztpUZtKUs2eIJQPWMDBu9BLLN5X
nLkEfvc5tDfh23vNgSxKjTKyq2YrZjsDjZjM3XqhwfLpZ2IYzN94Jih54hpeC8UF
QBvoswM7oT+INiUkZA2wgC2quIZa0oM3mCP7SKNxeI/PacdecVz5JudvB8TKUCpQ
cf4qlekcaLqXO8lTk67MIC5WkWveMVkffUJ7LyIuXwJ5NK9tSJfapoiBjmxKaFh/
ypAA9A9IcqmkW6zJsjxYFjl7VP3MgLqHbvsC1l83AMJ6BD7AoShuJOMEvs6XsVSK
/p9bW1eFrBga7UqJpJtcBBMLaTHpnkHu8T2HNqo/pFep4R/K4J6Ye27E+kuVG0cm
vnaCako0kJsbktNbHD6A4KcxdKFw+rYdllhBqtH6WVitKdg4xIubffOjNKcZIolV
HEEbXxz0QcW7XevGlrZKdNv0ayTFNpTDS0JXNyB8YXzFA04xgIFvlcn33EJaLkmx
LluCNH+fTy8gsnoEw5Lgj7JFdLGWzq5nyXxHWaod4334IJxMj6PbJmb8W8I4tQQY
K08mvzl2bnXV5whNAqDlh60ZLPuZQcBH27D+m7oSheQIiLPRX9/nSBP3Oj57ptlJ
S8WSCTOkdTJyj8/3aJqeMX5r/ScfcGVsQGnnM8Yvh2f3TbMJe5T9NcYbufrnHmah
2fTYFaPQmDwylRKhOICB4+DTfP+grmYy9v/18odYraEmy0M7r+1tDF2CbecMxhNM
9eLER5tzuhnyXF+jYx6v18B+LYuPr9Dv6DD5NwW5Gsi86cdr2dDXQw/Pr1gpxaO9
DuPMX1u84ID3Ytxg9TwcAKvDSg8xWY8Yn6z3RFkmlkgcAHJuZE0lh/qmTPiEpjmX
jY8sm4GWviKEe5/tpwuI7AwzSIuo7wV4nX4MIsnY7elfcpZGbTMOGEcDR2slXQ69
IA330MYvaUbiqWkf9wusRdzz4VAuhU4EybdQ07LYiI3T8QZeZ6rXBBuug3XHHavB
KQDKPurYWhNcDEl5mcdSid4oquZ70CsfFfOiE034crfnknxfGkQK40EXGh8kdwL+
JAnNyj4MHHhzwklST7xRKl8ZhQumYggtszxS+/5TcCd/BXE0So5vWvwAmECFDDNH
5dYEYC1EyFWRl84qFe3EkCVC4qy5sdAgBQAnjxoo2LcWGvBGy8W169/IjnmGjP/x
L4L0lYNguqwxT3GAtLBUgro6gMLjwS/dvKafj4t1l1+wN2CWuOy2UY/WFPtb6Vju
TA9k/FQzwhbq1jAERV763UqDPRHA0CUJhem3y3Q4vOVOa6dGDqyNuOmPpiQLRnbZ
a8Yr+P4PgztS0OFfM0IxJIx4eVFj3ea4jrZbtGzcz+xV2dnrmripGEpLQ6vbiha0
kF9W78ln6BKHF58wo0ta+OenMPzCLZVhOtqrg/B9dC1fqcVDs5Qi+2AoO+uQBxIM
460ga9cqUmVPJvPPfV2rtih97Qh49EAs37ntiIg/76onG6OZBzUxQE/c4mELn0Oq
wBXCB4Dij9J5JM1E6P/nfBlra742uzcVVydeqExYVjvJZvovoBXfa5R/U3NuYPDb
jsHw/laO4GALxPgWxutmt9dfq9qn+u68OWylOsy65sCGWlos674Xk7yg9UdJTadv
rK/BG6/pW8vRgXEST0SAvW2TWzpQTKIWkitfWyqlCznRi0lbl6YFz6unOqqnN42T
zaUAX1kGNAmtIJ1+s88ffn6P1FOgIm1qujMBKbXT+oE38cK8Nc8LJ8ON6EpahgcD
qR3+6Zl0a2b1ImszaVAsBG1wSJQ7C08drF809NLVcdD35hyuidJ55AsXqZ4wZUv5
wcNWMXn+hQ4wZCDYfVl+I1QKMWvutYOmSPDfmziI9h6Rdm+6bmdULeONSBJAiNlC
aIbTHj2UsOdaUeGWiJ/kcrz1I36PCUS/BjlwoTRgwvKFGjq6iP7CFXOCjE2fsQqv
CRFXYCYt4B6VgK3o4TXjM5dDJj67wSLWOlsmGgPVu6FZRH7ntx9vmo+AHgkSzqP7
VTLE7YZicO6GSfd8seSr084Gyakv/qkJ1lBVkbInVZA70gFSJ3Dgz2yV3R0Ifxtb
Jrl7PGC+4NicZd+SVzy+TKYixdGB+pKG6wNYB99VVS1BmtQZ3C8fBlppEXOLezek
blf6D+jOPHqWeCTtTJ5pPH8ek64fh9t8wZ8voBMy4qQ/QRkBHSa+AgKowFgEUTiT
J9SgEJOs6wh13K4roqMmccY7JiV6ZN7+I+QslvznRTh/abAx5B1+D1q0PJExNMZL
9/6vVrY2Ma6+gLrrJeDcrg2Ehm0Yo1OuHBwvUJe5UdASc6F/BHqxwhODkZIg7VZe
7jhhjZ+/jNCV4jxK2shUaDY5XtFyg/7qpRZj6mQGatAcmo47gI+WjsylQXf3gePR
0Tn+imLTUTu2OJZeGRBjBvVBXk76TqXT2XexzCEluGRYIqbg1Q1U2RZ88QxGHRq+
H+qnDvxXuLriSVkni3dJJ9/yCghH7Yknk9s7MvfEeYrfSWV/MO1f7qgspNcHhqZp
HUkwYSYVXE6P5YDu64qUEV9ODFCuLCkG8Qp8g9Y3sjhJz0fX7YD0o5zSmWqe1/1T
8fEhsydH0XqyZ94O6LSyCXm9RGi/eBvQGDi42pIvPeS3dLF0iwhgUblxD5h10fkm
P9vN/QDzxmBVcdTOKDhJCqpjVpAiIcM6TXnq07FEJ5qYW9HyyEg5a1Uk/pUZ9URJ
a3ji0Sq8rln9xtIQ3xiAWxc6IQqaHqoQ62blK9veWYJ9c0UNsDY57VoTV2eyEEZ9
bzT8fNXRSXIFciEoWs+4P3tY2DRP9PgtMnKP9Qg9CSbtY2OVSkvkPEL/R/3LYIhG
uh16ne2PX1izt0QzdbaQWbQwtBXsQkPi7n86MCAOsAUt8YVBgGV58SoizUNQBX9w
ja/dECCSDE5cuc5Pz753TjyOwSge6Vjb43W2YHetQZzjg4Hfjq70hZrjX0y1qZ2p
FjkPs+/oSQ7ryoLtbfYFeNdhMv3YkThoXDPhggmGxup9qeNjXka05j8qDrDm4UzI
wVrIoOHAhdiDTNVJgzrGAmD0uPts2iK6YKul7sBUjmDHyaGYkHdzAXlp/CeugD5K
BRnqTeUV5QXgBh9MC6/qy6wDP8ej/CNJXahzA+h5/B5u6J7FD4+9RrdprVy2FdE8
6e8GGJUwguUnfb0rOfqJZGrmt/k8PHFJDPdKBd/q7WqfMfaj3rZBdXLdIiJ7rkPA
GnYZ+2ofT1tzHPWQzLtWwTESmYZYxnl2GM4sm3oHvJsbmQnwpbVHES0X1NGfZxwX
56i3T0Ka/xhRdJq7PwTvEvLPmPy/OrRazpgFl15KCMq/5wf8e1zvPc2/fAzQUjWq
glo+uVXh4bpqt03LrazWTmG3J6YySKgyWo6At3+BAf4xkmJOfFFqfmuWIk/ZCyla
RIw8B7WxkDaNk9stVEaYYE3FIkuNLHZhA95cv6N4MVm8J3+oVpTsrweD4F3WjAx9
7zKQNcf5Vcsjz1H+oluIrFXYVH6RU4TavyxLPjQ/CsFLi/bAdhoowqzGbHA20omJ
NKFwHBW8H0+9CrgW3rulnpaUtbZVl6nZxFm06NaHaTvqbj1ywcSaqvYgz8Qd/+5F
2Iu1AyT8g/Tkog/ov9NnyDlBBdPQjZXf8yyogg4umXMLZt+VMiggjap9fzqgOQgv
0A6f87pT4s40VLvAqp9IXSPS3xhwDjYOAW2AWc8ukgVAiw8TnMEGbDA8IaRQ1hUy
fbyXTh9OhKYPINmBWIEYS493+k339nQmhwU8bkWtBfbgU+uPiiXtoj6xgiCr+uqy
y+gcJXdJXCfTLsJ2J5FYLQFphDPHb1aqLCvBhWhl56jqkwOZA7t48QraRRmB8ohM
3q7BPO3AImP42/d5G+s3jM+ctKiGMwoCaSxCxHsMij4pU7PmqEl7rgy6RQk/BIRO
Cf0rza5RRRoFCNJLktR8g+rB1pp8tHGcFFanstYaGiv9LFH1xmYZyU3dOglWACFi
w1Nd6FpzZ4dX+YDsMPAdmgpp7c5XYMLXWxTFI926WqCv66EtlCukoFxq0LZo6bYG
x47MLcy5msh49ljgQxJ4uKZMJ0dggvLkNykwgBGn5QvBD4BaB3JmyrK/VSEjhwsA
bWB+7EXuk2cRDl33E9VD9H99xVow1VXcsOWBp5dGOgQZWnDIdAYpyr6GpgpEEk6v
VI40JdUuLY80lwR1V00h3bnAf2r35QjPjLMk3p/8oMJW+EVAxIvzbKyJbW7FGE2d
QO2khxaGGqrfinrqegsKnQvc53RVLdwLYH3bb2bXybgQtEbkJENmz3v1wZD4m8sf
YKfUhMMmLDOSCfPYxrBKPlegGKLKrNpHyzFtXniMdtCb6+8wI9hulkye+rKKljO/
zXboDpWWWHBLuZf4T/BElwPKzU1vyj3x50qE4aSlpEwdhzKoPLmZAXvRWWh1l43A
jix0c2atHFXqZL+vHbwOES+ezapTjy4Qspv1MSmAdcV4eNYrH673uSrQO9fnzK1o
E3NXSkUJ0wM4obI4E8gKnevHu6dvEir1aAUoHKQy4olVEXb8jIIKIp6Jg6KfpmpK
Qp8glF5WISljbcb7DwOIMXr9c2GST7+miLb49MN1tz/maqhN8hh5Mn6w2fpoP4rx
c1mcUuz25RPk7f3StsS0/TyAHNrWGlDU4LM/v8/xr1i8B6ZCkffIRKZ44264/rVd
2wF8UsCLJV4OTmbhpgEMkHPeF4M/OtgBit7OIbeCv3wCLRxHRjT2ThFtNRtrapeF
HwDJ3JLQffD763JJwTbZpT7noi6z4XmgMFOrYGRdiXz6NiM1SQeS/91msM6iCjS9
HVGly/crBnuQ8DtoBc1hKWYKJqGHGoPsQSPkm7jbFG6scpMgOepKI5r5xG503QlO
/vXeqbsQRY3q3f/gtZF1o1M4pEuTLluOxjAEJ0DYCmatsjWIBqsWhQPe51g3oclb
9F5LUVFFkHxx0rhIlFRfRWphp5mEbp4aZorl83OfbUa9zVxjEJo11UdpDjLNcalS
OCveZqFlpUEmVHFI+w5P7y85DOKGtTKmHdu6twF2/e8OGtlDZ8CQCOcYnsXi9J9q
/LCjXJB6KFxZj+t9QqyMNfagEUwWTpPgSA5pE5n6Ke6ZRFF2Ii+c7lR8iaDsUade
SDrwRQse4bvNiHLbVYCXpelEYAkv6T3QKwndYf9JUm6nDfu/2yUGLox2DeBn+GSA
e8vKewzGg62zU4GZ8zveCZTS+T4Le+WCaDzFh2xDXB4hKlI8FVdw9QS0tNq0W3wD
g87ToRhE0dsEkpXxwSNIrYPH+QLrSWI36q1FhM6OgCISuJ7IQ0HkwOPvpQEHQRjD
sSNbRKdIoXuPiTH5xaTvkRLXidAa9obLqAQke5FunK+V5gl0PUuByotLY8Ce7R0i
vU4o3nezu3ZuYBlNgcSs1nvMfWSgTcuv1ud1HyIHhSFr6Qzj1R0ST0ezIIEPWDlx
5UqDuM+Ad4rFp45t9wumWumReVqMui0/fQHSwl7eUdfsjEN6IFifsnch6A6PBwJ6
tZA5HaXKKtaNbqj+98YkwDFF52bJ5QGM77FegnMPr6hnD8xh7e9cCjiJ7Hp6LUiR
EYdmXpAdRGLqpKE+SeA/LJe1v+ArjX5oZy57I7YS5mSCpqqgTBgUENBR69dZTocf
trPOcqRX5050EgB4CTOidYR/6kTjo+BMcdTzKvp0alWecc5DcXaY39JFn7O9491z
OoFz5z+78pvsltqqv/kJ7eS7tyiRAN8hTxzIBS6yYJL3/vT2ZNhjwSUQZiCZixxa
ENaKHHpKcith/PUu3GoHGdeztGtH+Z+IM4vy/9wgjJvvRQVE0f4l3ocJMo1CL6db
5L9jcm0fQDcNUQ6NfHYmX+ngoL6vqY6lJmO31V4o4KNUWl25s0+72mdGuppzR3Lq
NUyU11YNRYqakoLHyQ4uT54IUsgDC2klZh5siGZlI88I5AJnQGcWnxNciefmC5pK
qubw+S5oSl0TA51AYHiQkxtDnfn2ZUj6OUfmOaJ9NAKQOGuW2lXN+m+OuzjZQbqK
tOGWHnMKgklXesOtCOm2/3+/7+vb4LEX4lCWWuTNqFfgZAptXX9S3mkseLIdYQpb
WfALGOR2kOenVryUQqjvIgXE8elaWd5Oso3j5Ch2g52AmN6Mwyd0u9pPToU6Fgn3
xSE2ih56koflfHKVk39yi5jRoTZ2ciWZ5tblKufHtSgbuThImv2zfos588QOUl60
tDP1JzGl7f6dUA0nCstWjWCbNqyru92H2Y01xMh4fiMHyxqhs0Ft3vo8fNCzcgSC
i+fHXy2JI2rCNffh9rqx7clZqF1Tf77FOkrRigfYpgFkq5PDyaJ43sB/9rjHajwW
Twhes/eagUg2hECwCEJhh4ZbpLUdsrQ3oeKIVBFtcK6zdNEOtvGU2gPDz9necGrR
YnSGU7HR/8DKx8ovC7TjOtLiGvJ8g84mhQIuEWNp2h+rolUewnxrVU80NKM13feo
IsXa/nJSNZ0/mH+qJjCV5jrW/yQrddASEV889j4dMPb5LyvSpM2WgCW2x4gJfj43
GyIP1j0I5q4QJ0DUN4IARvDOiq7e+YTHgUfWW0X7U83HEjvtj8KCvjBscS0GQVj4
MuyB5YK5GtXAC2YIiEP5ldKqyqj1wxKnJ+5U2PV7og3IS7z4+Nn+J73O7r8QypxE
RYg/orMd9VvZx3qRccpuDbeIyBy9wlHn3WdeqssuE5qk+egDKftCn/EO9az26UDn
1Df5e5HjLwSkcXmgxNvI8eoigqdcI5bS3vm4Gnwpf1OAwvSDvavyTEL9EMiY5yGq
sg+bFsbpYWX3UAgGudxrxORhPcRNx7e5rb//nrkw3EBFdivAY6D/KAsHlNr1PiPH
2JZj4oSbyRlmZNIqBOABzjdkwMA15TEDMyo1nJrb5dUcJEXe45MT/fRqrEjiE8I1
k2sFrDHPDQePNXEanMhVTmCu9wv1Aqa+CKmwhccp0hudDgZhW0c7G5q/6xHnstZ0
aU59YCD9ZoNuxi5Snrvy9M7mUPM4ybv+xI8RuG6gX8VL5v/bp6qYphrfpA5UBZ9I
EBD9LlPnq4Z23pAkYBQwx5X1VXtnlunI+8JbVV/a3NaEsqUyoORPUJfWKm+/MJAD
Va46+XbZWqvtdQfe3uPCKchAIvE3vyoYqx4Ta1w6SMzNCp495t1b+anbpgEJ4MzF
A84WZhZejVbvtM6YOvet2LH2eveq92iiYWqQlyL+C3d4fi/YEQc63hCsScoXQ8Q+
mXU3w6I/af6ZkB+3Q698a8A3Gxm9KbSFM6RjpSVf1PE/DfUnLBRr73ksPNtWyzJ/
IBHG8WaHko3jwOm2q+PMYzHcRct21d3MkdlkWkuVk5PaNmWbk2HAdDzO8Md4XxIK
x+hQ+/OV9ALMzADrL8zaJ4Er/eBPU+ARkfKT5Owb/BATo5p4SdFz2/b/UDJH3RwX
PuWkJMDPIeBFwzvxxME4faqJmHENfiqhyOfzOuW4WpPeJiRS9Wgwmy8RN0cTQX6T
KuCj0rsQlBJbaem6NSXp+PDIYDCn7ZuayC9DhWV++F7hcg9pfPwCcODHPzdCYMQP
h93+56p0Wiz5WjLhPZ499ys4FnlC/e1NQ0xdMO9eGvbfxYcXC4wHcfIjFCbwUMp2
8/lc6V5FxwyKFhWgAHxsrPRT08BWo0bbW4p3N9FXQB1OdGvY/+tODweAHiJEU1pT
E7M3yyt7tIy+8g1cPDo0W7KK2tBHnW7Cp49X0YxV0LifwFSSXvsYT585hezP4ome
Zx74dGuonJ+YFGcaT/ixYskKWRNIXCGvUw5VbmkIHhS+wZbKfgLy3Ekzy23xmupC
H8uSS0HlLoxdD6B5cQJD3Ope66/DGWMOXcTSYkevydOCCQugnhLbgazFNlV2u8cW
L0mMAfJZeh+gJyyQ2Gr5e9fhvSRNBxnyKWxqIzrFbriid5or/mHB/sMDBnskaraL
jFQak8trjvLUhh0cVhz0LduY0HL5rS1RUvkpB0uOOIyFQcEv/gJYJYBMENsmrzQ9
lONZ5e1fHXcri7cvzIxzKBm4jpvCxQB5agOLBcifhWvVmx6GvBXC7FROw8i3tRIi
t6Udy5XLwhP39+TJImCgeJXmBL3a3E0dQ3GCZndfMI3Yt0fLMVGp4O53xgiZNJxY
69eoNpSTDcx3I9c4WM2CUxITFZnxbjVgzk7OUEuYbY038jEj3+l5FL7mx7rn8Hqt
6GlIev03yR84AzS+/nHcFJF0Bb0pgrBFoYOv12K+R8kNf7fTcGERi13pGlU83mOy
0aGGEAzhgqXJCpMWG3WREt86bz+HZGLFy37+XXYoqvBsNBLAt1Gokn/8tIIcEhR9
14uM6ai1mT4eR7BUDY+rVihcXdPGrSoDt7iavvVc2n07beFjM3MuxraidnEFrIH7
MYbr+ZJ3hTVKUSQX/G33H/+/jG9DXuDC+b6VAa4MDjd6Vik18TEGSzeVUip5Sbii
j7aWV/x+1wHwEZGw5H1W+gRfoH/E8MUq+REiVQ6ydFQUwpwi+t2KwsT03Z7GBEQO
B1GAwUQLQcCkL0GjiTc2TDiLB+O/NHUkAb8wJe+LyFRScy5sJdjv4ocDE+9lvxJ1
ojeCZMyK/9AL7WiX3rYSrqtFIv5pxlZRhuSu/mdb2PAd2WNGjFmZumXhgd0wYwdO
Rlccq/PJBAtIae87+W9nfMAD/HCC9lrh7vqKSFUQEMn/fi5iXa8cjDhzqZ1p5Yex
1uz+oET4hwuhCrPfjOD3/iTWo5RymoqdM1htC9S3+IaIpgTI/hLTWxv60OhYhR/n
K6yeiGTIeLb8vRnYDj1ltJdEjq5PnvC302HoHROql+aWIutktkXGRu/o4dIryEpD
Kau6tXFLbkg6sGt44NVHBFMufWllsunBB1MvrlnHNeQ89GRhZ2lxc35WJ3j7398+
CC35XcZGdTy8oV1VXyYjOfhRy1OQDfgUa2uU5SlpZTGXYOHkwuvDmQJKHGOKe3xi
BWjB6+aPoTiC/VE0OCckA02ifLaG8IHPt5IQnlRGVeHvM0Bk1EmAPN333VniA3Mv
CxD46j1hSg59J89x8CTdL6SE1VG6RyRpwpOt0AXU+T8Ap9Wg8HdRqNQ9Qgli2O0Q
sLBtpAstVHRBfum8D4IEkbgz4cugiEGMvlBs7sfmZJrxcXvVWX9DGXGHMt4/NQa/
rXKkG/Q14TuP2jO2OdEoeSeJGMbI/e8peJTQPl0nBV0F7d9RR6fW+LLWJr5SaDM2
QxONBZcoWMlXlGKbGiQEHKfKxBigULmupt/auQXblHmnP6iRT9o35D1/yO+YJVyr
6vtGPEXVOY8bBMLWOcfnAChgI8Obr3rj5ETj522aj+zoA06BV8NntcAUosEEy3Iq
pYOYn3vN9yX8eaUG7EeRBqsax65wxCDDaOYuQqXK2gflhABQG6B72AZ+fRwHuq8Z
PrJ72R2Pe1poktXK6u5i27TTRweTt6uDP3YSWisMjFG9tEIW2CvAHOcqT/RU9aXh
arM36zkAqNuma0qUDxuHMjgxF007PuUCQ+yvCHAp96e71Ytin6R7BX1KfgvOT4pl
eao85Q8lx5lLgRaiYt1/YMa6wv7ogIgNc1EU1cpUjCcp/OXbQR711YOz9mkdsMHS
F0Vur/+gry4WnHgx8ceXsZDYjmPTg+7P5653ERqr1cdattfVcAJtrPipuU6ORJoJ
dGuyh9mIAV9/vDs0U6zM/39ICmYypxw8MjM1HnvVVlvd6M7dKZWfaqfTaa3RHXLp
EFRTvLcwqktqPgiwGhyyaVz7b9zK0QSFEtQQBfYro+qnNW7YbIVWLH9kw3FnNlXr
qXvzqkHHOZVVwOIWJPkCVONYofRLjil3KEY4gxwyGwbBdDuhnd7iVB6G09AU6/1Z
CArOTfq/qq4kNshO6BViIx6QemGO+auTFv3tMZ3W3fN3p7Q08/P2jpQA1b9qNXR1
xLwF9dl1/m11J2lNse3abAsOySGWhQuqS92cnugHgR8/kFqqijFYyPtfy/2a2S9D
tFGNv8Sxmv4L8YEmqePBG54QoT1ayXF3OQjRhc0gXX4XNqAVfxwYSdWWoF1Lq4S3
SflkRJ+S3tdEdZl1E3IKyfPYx8ekD90RxU/bz01WCO22U4XkwAMNz0d4ufJIu+Ln
gLpaJsuhy+uApAVllD/dTOyL77vTNYh46oa/BQijUpgudD5NQZAQvpirXxvl9PRT
VRKzXxxihBC3apA53gEWg+eSftEvMDo4DDTRWRXMIwuMU2BtVIPwMy7kr7b/KVCo
5p+vvuPFhMpecxA7GE0RkXAy4qtVOXEb5dLErWb/GK/5v8dfW1/6db1O0vL3AzpT
rXlLbI0bKGfH7L/tWBV1/ecbaXZ/vHnwCbWmNnI5k4tdhn0JJr0/CCItDINIRgus
oAEA2uyJHkBd/a3UwiLCrEl2miH7nu0tulFIGD5z/P79ONpybGyQUaBQg21eRmuX
wBGIfXUU4md0+Ap31EgjcAwX+pZtDWJFiMuqjQWDbuNcnw2o7EyTZD0Jk/Z/5OvN
SsXbghpOSJK1zR4QMjAOjZWqto/8ZDJrWnM8ZP8c2u43u6E60dBl4IDTsvAN0JPh
9sPTTF9LdCvaCMI/pBKFL+yuL0LboIswPA23WpI7/MQkDFQI+mYXK8ZGI7RiUHi6
Msj+4DwTvoes+IzF40ZVJAqsJ+p0+gUrXQwhj/D4AeurqQdg9ZTpEWzbuM7c22F8
BEQvrQrbObFlj4RH3BmRtsOoOiu4y/qtCqp1rQLGBeiaERbiI9HWlGOW8cishZml
hwzBYDXzWnkMxVdsOT3+THmsVc4Cz5iUPoh+6xAFdZeLull4m/8CVY4QFR5SJW/t
1VtMbQKX+0RivK4WYkaNiJQatIhZh8UcnKFuvNg3aNecIzF45xg/bNxEOI7vCa8R
4NZpGMGFMR+SzdwmYm6XJ9scjwu6jIx01PYr5DkHGs+VCEUMZjeJyCKgZ54jJ89w
fPEjNQdAvYB/8losnJi5HgqfW/ih4O/R80kz8Vl69AyIwLNPWhD4CbIo+j+PH/o2
hDRInyReETsTHJ2V7R7ObMDD3n3CE09tHXqg/H+3buqXckfQR2oqj0qvreB/yfLt
8sNSIPjLIOSW9DQosPESkMjBO2lnOUNJUyvIcGOGs0uGu5mDyDTl8K2rdHU3ymh3
pV90gNGIUcxrVijTuNx1SJ5VgINee5Y/+ZHKZBR0oGRv8Ml0aGcOiT28wmKOZcas
wCv3RYa3MtmTw5k8JPFFmYN4T+8bAL9cmtsAZZVmu2VILafkIrfgbfrlvg7nP9GQ
iYoysnbgpCYaHqngrFbpFdObjlmcKwDolTBxnjdJlkegwvaT1i24pfH4ncdZMlJ0
5/TZZMLB84nCJdy50MBW6MEsbMGlPCniKG8eqvMTZnO0oGf4jlk94HuivpmK1ne+
Ptzokt3GWzEq2naQWusNgTUbcCOwVdDUSQj0QGLie65eqxjVwlxBXs9uHlpOZIbI
v7USD783Kn0Y1lAe+zVTZMYkIV45IVUX6tfQhP0BXrPYnrXcIec2nBrYxIRQ2oaP
7pEGaTRXBySdUrXJiYRv9hTxOf+4CVHxw0HH7zbanIvTtgKveBuika5UodOSDHbb
oTlDLXesFhBV2TuhQXeOLv6OF+0v620QjqsYHlTJMLHRs9hKCJBl7rzoO/5asUEK
rewNd8/IzwW251BjgPKcv39OEzalXRbQYU+LxIGtJ6nfqQDnOmYDWdUg/22KA9lB
kP+Frhg4W0RQPY1RcKvcUvfqE+ZJT1oYIntKkXSe41e35bhnC5K+WWzK4B6xzp8i
Rou9Rcpu/uLgYUKhj88FJ+Mk5x1IxquFs5LsUlO39BQ7QatAE3kpVcPenPBSK5fP
BB9GY9wCj0qk1zl3/eGkO9lYB835U2li/krhy9rVF6iBsojY3uLSLLNm32AYgNS3
AUpOj4wQYkampPMiTF3RH6bMsZofrLYM8TXkPj1zFyzPcRrzEdYuLs0cIyUWv66U
z8yNSUjSpVAQbCMOAbgD35CU1arM/yiloyijqlhyHdmv3tx1+4TJ+SUjl/V0oEgI
yYAh7vR5O7kci0JNsRP51WI2WTqbv+zKcjbCWn7Z7ZTAw3gXJpD6JlnxsBRG4R4s
zrdipp8ilWYtiP/7/AVT2lmhGy3YvivSbxXCbV34/mjQr4f0HvIYFuwNobNBq7ne
tbErVPdzKtUBhyFjR2AebVQoQcRf+uQJJP3odLJ3zQ0aTm1+7u6oxQfbPvTJV31g
BDMZzR1BThExdB+UTOgFeRMQFWUxeyosah6ln9LUlTuZ4HvIrQ0BQJdewZGWwQCS
5YDOtgnum0ejnmwyDE6JRxx7UE1BaWhflB8hHMMyjC/MM6M8wdPv+syAp+8Fkktx
y4WL1+tMNaIZWis45L3ITpcdR6MqmMkTxbchVOa/mVkKN83tY09KRMCgsBWzBDGV
KTPwJSr+XdZ7GNUHSeMhvQ4mfKQzpmrBk3q0qex2TePmEQ7FAgSWndk/Skz+rtsJ
Y3eL4E+pNsqxNa8PXki/31uGiZoKUtPvzkRmA1Lya854+TSVEOeasRsDobvMxrky
yaVEp6WFBzwVjhEM5ft/B0zBYZpl4P3eCEask8yuj5HxTgNUqLPZqmP8ONdcXRnw
NhZik0yh5nmix+2kRwM6AHvPcZQ1QImyYi+o+QzBGtLyi1g+1ksQFjb4wXVvlxE3
xtDDNOCbO9Z+MV89rMdz8aDuizUoIPHJbKTF5vfuxCweptnx+Rw+SPf6MGdj81ZJ
dYU9wCC1pNl6LkQbRTcsXIhR01LSeXzVs190QEv4SZnKEEVnODbrq3gFx2DrPYvq
Q62poAGIAVg5l8DiDzzyj93kpKENuHmx4Qu6ELqM+FeXwbsmHuobb0hCj1FU1gsu
7Nva8ILTqneGsKLpNwuJJXz+eaOPAgzDY/A8O/XiWFsv/JQO5rgBJfULWrJsgICD
WhT01f6/fVEo1TDg6j8kIY9BIRJLz3dxp/abfuW8kIAWX4RRS3YxJopDTlXB6MTe
Nnhd/UPuUFZSNBuPFI0VdxP5R7hAAKiLtn+R7xr/eu06tuwmQStEU94o0+rfMnpc
YKdiZwxN6CRbSMcCa3lToTGfVsC/b9LGLHGEHsMOpI8D/5qBRud3kNPJtIY0kL5g
wWBKiJwUatkOA2lqiK9jbvEqeym3HiDWzyvrP2Hi0JqXd4LqrYxxj1KJp2xDKuLz
LG9DKPXJwAN6DXEUpx0W4tgzyAq56VgsBAI6mLUp+7Uj+l+YUy2juSq8b1ozE0NK
vhtkKIyU9OK5MJY8QI/1xhuht3iC/Fzeq+fGM2FBFUJX2amNGMEWfxQl67emfNGu
daULT1wewjnd4vIV8Lq0+mVgE/LyOGZAIUL4hBTS/7OApshrbZnC3MGroO9OPSxe
Ith+HGnPCGQXtA70in1Dd+HhnhQTv6fhdGN4D/ISOAHSk0r2mcbANZM/eZSEEfts
QRbjUb0cg0L2xB7iGTcRp6tBCyKbbnTV2H2nM2cnYQqJ0WUH/akcJiW0Z/xS+aLl
0a6s1oKandYxuZVrCtR5K/i+ouGAnj+oDZyJSOt2Swrxbfw7r0s6Wq0vIFC6UH0T
+SOnQd47or8mWa8OxB43YhVvyOQaL0YXi4DwXd9sxOivq3Gc8oaiyrmsy/nLrmyo
TtgMRd3RzQjGqOF6uiGCZb0+wV5qvaD9sxHbDmE07U4NA177v7rA0YAHlka01LIi
brGQGxSyVjxM0S1MrkMq5M2RCakdyFj4AHQ7Z5+9FwiLTQtloI7VjOnHL1xBuCBl
wwiNp2YYSOYhdFAz5Oy8oRqqRN5jewTBt4sO2e4l2u7UplnLdgFT/JQpdNIaIFmA
gzZ4rsPBb3hAZroT7e6d0FZGAk7+tOsnGstSuqDsbv06I/jR/yeBZ0IxrhmiVQpB
L8Oqzfm7n0wssXLqFzmAOmuwq35KNpx1p8Z0Kvvz5MGuuLOjJbR51oYxVN0vWgwT
hbrQx/5r2l4RHu0Ai4NcdPx1ZeQKSlpPHAmM8fKTm5a4MVoKVR8QLKfL/LcMN6Lb
pdQk5klaJwfZT/AKj4IaQ3vGFgFDGLJogZbr3tniFHaNncyDkr5No/etM0dr9Spk
pWyuHXxsgf3CrjhYnOAE88Vx0zacbXKVns4YKPXqAoBEY4XrcecG0Fbep9QwHCnh
8Coxj56iqHQLY6iim9CpAcfjMZOEyeGmd7Cy1eCq/MMAquAMrnGPN+nrnoJX++7e
28Jtsv9IwIy9Wzazeocpe0R037f9W3VZt82nYzYbhGl7+d5ISLRV1sQVw+mex4So
44ubQCUapvnRmKbaoSHfGY7qetkEfi0fnF7KclS9qD5psOFsyay04VwjRbRwHGrB
BQU5LhKbNIvCYzfHbTDNRSf3wK3QdrVryyKn+ylzjABpibhoKdrcKXs5yGtKGtGZ
YERTETzSB9DTVy/+NIqrcpv79VehO9iryJbwvTwdnJPg7sFj1/OsPne4o5mAT4uF
JCP4pd1lGdzyh3G5FhsIRWP7BgHFdnN9OkZSKloHjw/11OTx1MOErQX74vULj/tX
5XpXsCXwuQjUN8Oe7MfSPpNM+HEN9j89SCRqOV+Xngw7NjZclmdxF4V0dNQsIZXv
T+5BXFedYtmg6NSnMuBmjdf433xWGxIsVHmtMcNxiXvdMBIOtC8MX5oXb7NOrXWQ
W54MSCSPticyuWO7RkG+ADxr9JFe5uySB+8mkDg6eDvQz+nGFWz3BzkCS4iWc3OW
dkVaHCvS5kmobS2k0/cvnFOYZCy734zwWHFGrtbz6hp0UfVHxjPUMaMqsdb3dg/T
sU5RlMy5HW/Tc+EILQ5WCizuUeuWv9w7JnxqrnRpBwYkeoiwBe8uI65rvitn8Hfi
9V3aZs5sC9FYEMbFoYT6VZ03oMYsKLHmt0RdETOu4wII/GBcZVUZ7CGhBTixQiVY
sZtLqzQ8QPEgKRICN2b7IsfFC4r1vfYO/FlR0OI4sICIwEkNYNu06tSlw2YBM9Tv
ujyzcFuOKrkcjKXH4RjMvUdYnpTJgT84DINQOII/Vlm6y/y5zNc1g+3bXcWoIGBF
gPnTh21zZcWmY/1Kb6Uhq1ow7B6gs0g7+1y7ThCLvJ3UMMMjVSH5keCX2mofPg7h
peudZpZdFkzoIBMuckZBCrE+c9IkNkNXT+gOYstoxZNFMlulbLY5ywemJ4fK5oDX
nk4Rmx/Gvpb2Ji3XYoNtf/rk5vdaFMfHMO0OKBOT0UNogtyqzLQOegVTqJO4emmE
G3WlzL6mr24mn8Mn8S5Rzak7LoGLVspSStkGibeJePHEznfjJ7EyRQrhF93gTmEd
aU5xXYsmLnfoxITFW38i3RWwFxfBaTAbvBIx99yvgMrl3x7rO8Glzh/u7ouC38TS
d+65qelC4lkU8vgndKmO/UccfE4IQimMgtQQznrBl1IhxJ8Ai85EmI5ZWx58j3no
wVANNbjwveBNkhRkt6HzeCY0D7MDhhHKy+7HRfB9c8PS8qnREdHUNXP2lQa5hHb/
64OqLzxxY+evMmUtqzRGAWM5Zv8tZYSREC4/xzN6B/FmJhtsd9vivnwGO3MXJqWT
KwnNoeoqeCI+F7FM+79mW8GRufDNRv7Hiit2JPPLBKca/xt/YXAonA9C5ZWcfYfs
6xzv7JS0KPE1AUpQ/BRGvhAcCWhRdaiwIAlme/eFiAq40DYnezuk8fw8DHrLZcsN
eybdx4DWD7n7DAEtvJUdReg2EMjbPDB5NeYV4VJq4wIDESQiMVY39DyMgmF1zfvS
McrIPOGv47tIxxnnaWzsGNhCTfHt5WHVG2dw+Qni1WNQyjWpU/SkwoeeNbb+p+Ay
JqRjo4Hh0T5VIJ6Me5hQdNi1WLEK6ubCD29Jkj50G6hAhQ2glATq7kTDQfhkVfWy
ztZb3EHQh64C4D35/JcD4PJgAEEZ+wOwWTmvn2pLwIHshm18e1EkU3rU1E9XHz7R
6AThbJ2z+5TNAXbQB2pvAYseTaRmahJomo7HjdUhK80BdxqdhIsZ1S6jyyiQA+ln
MekYKFkWPUA07Z+kCDuUl38evTtAUSQW5lRx1K58ghFqWebT6qBc6DDsg5icP8dp
2/3QsvPCvsS9MfaWiAgF9PWmHQ8trYs+s2nLrUD9FjgI8Grn5PI5cma4y+5EzmbI
fjAzN3GU+9eAIZhWInO2JVZKNiVgtYwmIAgRXnnppUEQl9MunynfPNMEVeADNafT
1HmiEGJWfVHGLZrs0r2XvwP42abNFSPDCaT9kAOqgTpNBZP4mgvB8hB/nDQjCxxZ
ruLZdGj5t3hi0Jfe4xDTDDYOmxB05cCJuAXi3/Uin2/4U3v0kFG9DyAQtX+BWLkz
Gh6jugCsr5afldHJjVkzXaSSM48qOFaU/MxjDdDamF/9pV5XEHHM4HNaEbrvQ5Xx
wZO/DKs8CNTr9SSLvIqhb2k7L/RKxUg6w+k+crSx99gcoAWG9C8tZ23J4RYs1hVD
WaEegkmDSIS/FCV0ugwFU6MzsiTRNwHxEIMad+SeX1PSPGwsRNJMpiOuTEmsUbn0
7cSkhyD9DVA0QRN5ZfT5r2kXIuK7o11EU5xHN+hJV/TXAWSf0yoKiCZBPMIwAnmu
D1fukTDDkDhrhK8NrvfHK3xcq6K9gvsdVY+ayFXvGpupM4BWbVr56ivOGpYGFs2+
NakEVjew2PwQqnt1w3JYHe+Y86ZoPZ1JlRrXr1uzqRZsO0KFnY8Q6Sa7NHqLpDSr
1MB0gc1T0oYobOOoLcYFr8XiINUTaJAYHoJ+3jrr3rYLfYQcoLlzTiMw+s8fXBH0
MR45sl3nfa+DeFjGpEMwIHvrm+rkg06mJDzBt5X5AhKY4fkvPdIbBsG0yiB/3I5j
Hlailqu2MoDmwSL4w9rJotsVC/YW3ksE1mK4oOd83Xtd3wojYDCksvR2g+mXHHrb
yLCcIiouksuNkrYmsJek+b9CLiJEG7X+5nX3ADUwgB25ckJtJR3SpSHqZfhvND8X
Ra5fIX+RpH+kpQonEE0/SYFPvUx7OrP4sLJXEx4ZRncV0bfGmE+9d/xrLTBthtsm
upp20XKDafEA1MyY6wNt1W4R+Q98hI8a1qXXnBrc6KJH6IKmzugNou1zgj4Eo+zP
IE8t9mjWj+xJh0FNXSiprMbaLx/zrNXesoVvEtx0zN/4AcdbCmVOu9Koi+fJR7HO
ZSEa+rNZigGR8SrUFKgVA6vXnu92F+PfWJFkFAACdrlYoWna2Z/YXlq4MdPO6RMz
Kat5tVy2n5uCu979M5QI9NecHfJzBOuPnB8QCsb+lqwryQXIhzmBwZdTxCZy0bOQ
qcCokYqb/kfQFq/A7zuapZsb8zHn62BdOKzF6Q9QVObQvyLZw7Fy4AY3jr7R6o8I
MDovHMCowyPHnL5Pq33lX+yWkd51ZFxs4usqsHRqK+8amktUknwxA4OYnFXKMV4v
Kf0ixL9oVUsEpp+MvbCxe1XrrtGtEIM6HIWFa6TzxsYGHCAEA48DFph6gU6JXcH2
zeEbmcNMLhIvGZQUPTNXVqufW+NyKChKgOfZUawDIO5bxDcriJCD8daHEFlFidzW
wpDWFlWu63o+JbirCaWC7qcdMhTX/kfAmNzDEZmpgT6wnV5wwdv/1egM18rtgXvm
YmCOB/NQLidIbJZO3LuMOeEWpYG/XTNMVKm0kKf03eYKjAGhIGao+5Diirc9mZTl
lzgUA/U/+FWjmvC7Xx0sWTFQQ3p40U3Oc9UpqKJhoXh9hFC8pUueXLqMKof5Vnm+
J3S/QqCM7jKoKbbmYK+jC2oiwAww/QUx8jcMGR+AZaTSlr3mtglQO4L/T2NreNSb
AKiPkWD3ZK0LL48/cyL9Yopshhq27l+9dRfKVU7nBPS7LFfXS30JHlfrjRFtgI4w
9+KTc0FDqI/+D289J7Xy46e9tsjeu/pfxzMFSuSSDUwXNuFrXKwEE+VQ5z2kDnpl
T5HFyiuY0r47cNEcZrNNMPeDMdRCz1FaTAUa7nqvCDjjKz3u1QzyEOgktmBUGiTq
PNMeVrtzz1ne/4oYLm8PH5Prqg1824qKS4vwC9OqTz6zWGWFkF/ETylrDT9gdUuN
oRuzwIWvja50VxO4+hyY+uAL6JZN4BuxFZVDiXLcsGQlqOng8PQSFjb/Aw4cELbt
rD1wzaB/aatzGedecmxDmqgmvjZ8WxDZ6hlMJmGtW9Z3jbToN/ssrjWOn+ILlck/
KTjOvWLlVI4wVY/ICSBNbGykjSKb3qfKm+GfKV3USbOGXf0EdL8/nFjoeZyOhtt4
/O0UKQ0U5kY7HO4bqxo0QKx8WjTSSwegdCf/fWhhAqGqmYoDalIN+WCQnVMfWAh/
XEK6/13KUgDhHvUTFs4AxEOYT54GhAsQ/MinOxJI4q4hWby5xBYPOUPSezSQXlg/
RPdVge7JezOcoG5NLNPr2NPTpu9r396AI2h9SwQZSAl3FWYlf3ky4IMXEu6MB7Dn
teC2rPNr/wTP6MrzTiQlqjXp0z4AKD9i+uYIn2v3HiaxiTPQ6HUytyidjHliT0ez
8Ns4CSIyLBUIn/hxFVSllxgYGitm2Sa3NGNnazW1uihI9AlBtvRBIynU+t5IoGYg
krOh0aA619q0+eJUEsXwMdFmtaTKkqvAi2mHtI7HFFUfRLEUo4ocPCCdbTmsi2O7
2I5Aup+WGe8hct3qyOJZtrZ7AGo/ndbtZDJoZSuZIBTBSp50T1H49hCD7vtgMAql
W8V0YFaDAKRoD8toycGcZrWSumgmwhMhiYwr99J+pidZnSISIoNYnJgAudO4IMmF
H6uKSBoam8XfHCAF2VxnQyIMcDqMLk/WTBUhQBpZO9O1Nhq4R2n/8/xEeqdNYIzc
35mDhKniaAXnQXJGrsHcJof8zjYpN43Sqy+dqYcGvHv0ABsr4bSmxk5JGfX/JRiQ
oDA5zLC/yFUqAXiIq0VYc/hldZyjXma6JaWhauG6Shu/e+N3OJP7bWBGDfkzuf2d
55xJj7YjJrzhIrRrYcOzaehUMSqDBgUVgRI2zsIJUvWe3h+r2GcjXlfbPClF7zSB
fgmxcEa5BpvkXFzvhYHcj5IOG8nO6OZExEivqoiyEKPguVrLxUiw3lh9GxH+B9KS
no4jne3Fbew+sXM6CSzZW1K+ODn+bU4GNlslpsqUTWfJu9kRa/xJjAJ0dQmpreSC
pdYbxpbjlMzM/F01xFZJ9nRcO7R94njjs3i6a6WMZzOOrj/+qnw6xWGVUjURD8D6
FIhXsnPHlMbuMckcs/J36MPhOEWJML96QvXFRAEFj2q7lCC9ZsV+nPj7Me9NuGsP
l6bXCAUaOcX3iwhSksMlUK8/vOXtphTb7cbND2j+7qSlddHqmMvt2JRggPKgBE/L
QMQ+z7q9abwBCBRf8zesjVAobl6WqNbxb0fqQduZBjCeNgNMb47SEDI+5y3o9pq4
J8isCdZUmDXMg8tNHv5eaiHJJsENwfEC1Hpb7svZLzANRHPAydiBnnlpPSBdrqLP
JZx1W6M9ajbT9g2AtgpLiQjQOksIdUA5lfnHkyYOd/3JWKt/Qa91Bm1FSh5IZK5e
Y+0PK5A12xKJdgVgXNlcx5C03z0x/cThmOC9w+4J5iw3VWQ1rdLXi/MK+nQCQzM+
AUeuBXclNXMZO0qDkH7tEDou9LkpjxOkUsIgWLCJ2SB1NsTyboE5nu0O8/8ek3QV
romPyd1/UyiAtj9gae/HH71P8uuwNnVM1QQT5LryUr4jTyCYH1YincAsFihYvd57
b67GSt7+3VU+1grNuLa6uqeneANgMAgkKBU1FZC7t/b00cVAPBnjA+qsAXQQx/Aj
4CBQyqfO54VYgWwHySKgld1AMVmuZAYO4NXICy8bYlI+oSypyTgo5zJkV6Q8elOV
n3h5+EZ2PKYJQO3tTrWq3dzn4VQeZDPHQr44RjQa5494YmMLIMPabUpXgUWcf++S
9cdwCu0MzFw3GzMtZOQ4+mGJUtRec/fZyHohJ6/F5hWCREkdDjIoF/ID4OhagBmX
UREWlvJFDz3HxSxUten6SUFmwLnrY4M39KhTG5f8b1dp8BaZChBtRwZ+2EyaOCKC
lToH69VtKMhus68XrusJEOr4b8YcSr0uLMvQogpl2dU3NJ52QzsaGoTbl534Iw/E
JsDHxDAYA2WwRlaiQPCCCvMhPTAm2r/KjH+hcP2HPRPN+w8GZ4ylbuPKkEwH3/k+
C4aqz2WDbvkOnRhZN/ZgDtjj9zuU0DvRE7UyLLyqcdSWGfWyEdgnndRGz60527HE
47AetfVU/2XoQuQYPLx+f66EinOZK8k1u8OqxKCvaxdR6wfajKkYzGiJdxmW+uH4
vkkC02+jfIBIESUfug44OLl+idzvtiCo+VviWHLcPZTnl7f4HYpzln71Rn6frlJK
CVflD4H50h+6iEQhlfd3pkiALfHGL/ao77TF0vYh5JyeaTYWWI+MvSiD2/18/f4K
tiW0VcDOlSJEGqACxdg5P9JVvr8a/ZOu5wU5mb+QEnHMeOSsXEe49YNxG6lnOaT1
oHDSxkN3cgu8tggRTWNvTb+EoBYXQHMOXXeAJfpEdm90mS3lVdtkI/feeTHpTByY
tW5lAn7jA1paQoUlNwJrV3kkxeqpk1Q48LTdS86QZ7a4JHApkyKQ5fMz3PqXXfK4
8QnT/zdr9rtmngynhkk8mSfgSjb9832OYWC/T06wp00v+h4yQ2PRorv6r1tIQkSk
YPuFYxLdO7KVw9KqSWfk+Re9HLCEXXd1B8v0fdakyqSEvsg/o6AgG0EIH+Rkpn0m
XxR2NBMAcTeBphTabQpSD05MZpD+FzVpHCZ8/zC4bYixsYUOyR8FxfCegfoeOaXq
5qGkkCpKFXH54DtILEd89d/TVYX8Si2x6WfZc48rBOrTRRZqdzqF37N0fxrefCNB
uXj3A8G702fYjJXrbsIQpfIwiKZZ8BuDAuINPwoTlTKsLr5KlyP5LFISN3pOVvab
TkK5kvIh5ZNPsqIlrH+fluiaIZOVrSadvS8Ji1fLTM4L3e56dew71L25aXcN53QQ
Jca8q+wtyI99hvuQF7XbAlUlPFIJ3ng6QZC3dSvVuofMVtqvkbYFhod4toPwYhOk
pbtkTWZUwfq9V6tDq2zxRFzHsG/C35TPqmKR8dDZm8rf67+QjDT9J59Vwfsrx2Eg
h4AMDhfVG2eTM8TURtzeBiJn884qstlLqR3yfhFS4GynucqrNQAMaC7cCejsHdnQ
4SQs/qYOgZPjx4bGbULYnnVRb7LF3v9S84NLLtJCzCfwjp46Pvw6/bI3JYz2y6rw
t3KcJ9Ao3RDTTj1VJ/LxQiwCw5yG9o3mLJvU6WE83R3iJmuJhcGDy8YYwr8IzsTM
DFmsr5N5AXJzNXugClGELmvyUOR3voj2GyWM/dGHWS1y3pOwnLE80IURWfF3KWWG
30NvKuCfLSRjmPax40laqC7DvGuhHiaJ3s85lr7oGkMXj/1F04sacGb6FrQtPBya
6tfBj+RcQibEV31GSTVD2meIyuOGyAzC5Pf89vgd7+d1EgKaGFoVoApn0ACzQZmS
5LEHm1tydBAFXQMWvcv8HuNu++3qWUWqPkWG6F463+jh8Uq+uhBH+p6DZuimEbhy
LYP8+chOBg/OkKfoam3VIqJENyssoAcn2EBEX+bos1LXUr3av9BOnB2Y+ZW6MyXl
kKRmJL4IY0Oul3YG7w3znVfoNIYPkepONd6MRbTpS94xuumfl/Y/gR6HULSwxb6v
Wk37XJZYBCKaju+KrZI0n5M0rBGxZ6GkBYE2quU6U9x/iIm7KQx6NG7N95zrFJxV
swEedGywrpksRsW5zkR81YuXY2D98t4pquNcIm4jELekilyo8or44kzfqRBeQgQd
85wtePTV4bKhZOGiDZQpPimr9A77liO6ELb+f5UrJwoFLAxHsTxAEpn40sOTcORL
b7fM9mhsU+VBBqODd7iNWZeasHg/F4bfy4XxoLEketK5feMqzmDIqFQvjh7PxZ2d
Yl5jSlOU013aFk/Y8pNAQm5ORldL15TyXMeSLex5bedAFXW8bX09zocY3t5Nbjmy
/HUyh3t5M1dXaRaMWpK9veSqBe87VPFZrktY1R4qr9fp1Y3z7sJ1ETn9FtQIt0rF
3ay1UOhv+CfvhOFGhlJQrPU6xOBWnrEMteimAZ9DyqnEgpobr6wEIKdyY8ixyuuP
kRnIgJOvndEzo6KbLELufvC4MoDGx+ZTsNeWlVGFCRbfzsXvola+XfJrF7PgaUbc
Wri4MQxrsc+vEhg12liouquSlnI1sukQN1f3PJXXWIauH7CSjdBZshEHpC7GhnpB
CowRCKf4WihwSopAu7A/+B+/AobSTHiYGPRBADYn9IazQ3YY/IglTJ/eg3pGLD/A
aH9tg6duO1ZlCznxC0S02yzM3kI6wwxCzZepo6lrq7HV6obbcyJik9KvXdNW0Cup
ucr52R7b7b5r14So9/X/R9CIuMaMR7yOyPxrbk6BTAg1xeJ7T85hGta93Gdm+vYg
P/CEbd3VbfVj1VaYKTjPoazlTc1kDnRUXZWNfMpYu5OH1eZLz0zbWLqdgp6ZgYB9
afgvM+VbEKgOSxUPoI5BOe19zXBDdE8WmfhLxC2AbfL4QEuO5tz7ndsbkQHE9rEu
A8gfR5MEJIGy/lqhUsZiTIsHwamu15HIhHX8Ft+TN9ETCTT3wwD+fx7zbKAeP7Zl
ucJtByTVh07Ln+YGAm2C7bXNhvbYdFh35YLZqpz9hrdPuzNWG/dKWnkXRHmBdg6g
N5wr1IqqXQ0/SWeZ5nRkkERw0+zJsWBh4PHHCWn+56s/lpgHjkMxGEalCYdzSEAd
mv7w1HYf9rKC7EgSB0geZy2GESyZ8tc0Ru8uWph3J0DqWHtCxlj0DfCboyZg8Sv8
1PYzMzMQLyoU1vZq6goLPTvCvmlDkp5D3pz9KU6wk+5THuwgTRp3YvjPP/ZI7dMQ
/rb3Sr1U01g8q4cPo26Uc6sPK501mx2hjaKwKZYDmMpmbZQCaY4N6JNY636Nqyn7
jkYOShHfa5dELr1ccWTp8IzN43KrJ1Zr7NAikITLfh1+lAzYAt7SfvFCqMzzRmb4
HeAfBO5xL7ZGVCY794ICiDtkeCZJvobnAor4DUprRxs25pOuh8lPnsl3GTanAMA8
UQWc+/UhFskwXdIFeIgxA2zX1YI/UW8mn14LNeL8yADbKJPKQ+yFQ83dDAYhp2md
uUldHNeleMxOGOL+tj55IDMEVZl0jAK1WpEB7GOg0Q5dDQ0RorREDDEcFlP40WvD
cXSHWOP/wRvDHoBupbOKj5AE2qZnLPsC7UqKUEKIAYPyI1DSaJF++BHerwDcFDp3
sRr+p0vHTY/IsKwTSfh7tswk8Et/kDncin+zHZ1r8eJs2vPMt4l7mdwlB+dbYJD1
+r3+TH822yTCIZ1O/yt+5Pfif5+ar0zHOQWLlJ2Ohu8/jtG87AcJwrvLjmUrnhbW
pF8VAMFJyOvjsqu/HUqz7UIgtuekNe8wmn9j5X7bskTFR9WglSZEZqoRqNBXaeTF
YMvB50AznwLAPgHPlCPUKlDc3Xsx4+nt/9OV9c++wXljiOCtH26RbmI9Xf36uKoJ
1CNoIVnm0S9JIepa0k1XvKBAXCl0dJO4XaRTdw4b/59+VbaGbzJuiODAoxvMWBqM
+1u59KBttRA12A3nUq7GBbSNT02QQctJTdEsW/EsXdsG320lXLqX6dCLUQVZkFBI
INfsj3u8MQsbv7pmOpMQL22SDwGqb4tPlKgPcn8nVCjRJ8GikrXHxm2mB9RMjY9i
r6HsKCNNE1GkHqCJVxWp/MdA+vlqAS70YHChD4VDVYYa0wsabfYgJeFn0gzhj+NM
t0AUKl7hruP1HXyTF9CFeXbUCRnrpMHSVmnH6Cz1Jk85bE9XMISGiIlJtq4tDHK/
JmPTzGTqWpXVesDYbpyl60F1li7aZmhiwGIWT/ce0e6UvjRRJ2m/8phgWtDqwkbM
+avgmMMw9iyh1keOOrpoJQPUJamvgdEsF9ETFoiq2sAmc3hf8o+v89IZUXg7BTXz
t+m58qWKdjX3omQ5Z2QnV3xhwl6v7znADCnqGIhUExLl2inBEP0PSeX8vJ+d4y54
16L1/MTvM727OlCgzd5h9kfvkFGuQoOhQntNaJXxWK+dTOBc6qR/XSPoNZF1kKEv
P5RyIDEgdELmiSb3NAy0yLgtMqsVyywOoLHteW5amaLaqxy2FI7kT3ibXxI/3JsD
CX7RApD60MKjHSIQscg3+GuyIzpnwJ0uF6EGJCquHfSi3f2n09AxHVo05wY265TT
GEoTMABPf3V0eHX50EJTZDS7iOTZ6VQZuXTGLJ7Mlz0MmvPAPDE1Z943ELJtSySd
j7U9EKu2AENeV5ELwGi6hmlKPiwvL2ollWa312UQZJmw+xBQ11HgpSkEVoeZm7CY
qqFXn8Wbt9G1A2bsDV8N1zqd1WUX5wq0MAREBoZl0a2c11UBbZyatGZtsP7uT8Xh
gGdT/1wjQUywRcutw8tvF/hgD5rxzBbXdRVuQox7JgMFVeUxSS0bbPo8xdgWuv97
WOhBudUxEeb/uFeHz/wUnt7aUORDm1TBXFl/G1fbZbzgXFscgwfIafJWrk55QVQk
fvT4kDK08ttBSoRMqkOo+PuDvOykI+kjJ8QgMiH3pmym8y5Hoi+kDiv8dWkfYXic
0uDY9eTlGJ8zBSC5odw32ZGmHznHWOtN4/Xi/1fnniNYfypP6HXTBrdWUQ86c5io
ndAr9FMCPKeuYitdTetUxooRjbWEWe45N4o0ym4saewP4YbOPtAsnlnbsCJKa1Wp
8hNRQn1xvqoX9nqkw7mItqJ09m1FHRUjUrOla0RakvshHlZ+27p7sBzJfGa46Pg4
O09GEqRHfEvVzewVg5BSJmsPJ7ulOwCs3uN+113iBbNFlmPKYN25cUuAXdh1OmVN
g2QuaKPKo6yNLgmIxFi7hrhN6nPbdZerh2rB57rglzP5HaQqJkc3tt7N/7ztRCMq
8Uzu3PlNfR+pYIOuxU5bKgcARdxKyZViMUwG0xhdoNApVSlj6V5EoLHFUn8sCtRi
X4EdqOuf0MF3Zyn3uvnC2gvghqkNAcE0SdO3PpisazVTO3WF8DiyunlknaarB6Of
PcxT+5uWCFrBcfyjlXFU64rKw3Lz5K7VLcpiWsO1c26+lj3CtUXw8Rs54MzWqOQQ
yshYts9kXlywF8pyEWnkf1Ztb9q3isoEn9f/RHDLoQTVVdH6yq5Wxf+Uap48atue
eiMrUiaWYHTIcWEDXGU+ZJIHSGSL2zw/q1AeN8vqU8PpyP7BwiaT5RQElY/JT4hw
h5mb073R9yI0dfGvMVQrKgQg8854XNGQ3xjVG8KkEPdGBynTQgiQsmE40EqSLycd
62VyYJMyJ7mwFmlnoAPcxNbgbzoCgBHqCbrFs9dzW/kCZIujC0DI8qVh1qMIycy6
X65jReMH8109xGzRzZKQ9AR7oKbjQdYbl/aM4kGSh1DBEuyXpRsceLDkxaP13p5a
vWj6F8Fu+eithc7MbxU/vymCJ7kshWBqobDUIVjesAoU3/HgULAfV2+DkBK+RlLO
I0FS+1n4jDz45riT3454avjXf9aFb2OvCoBL2TMT9mFDLmHmdugXeOOFBzTU6Jpx
4kKr4Vlc+VKOqlxgMX1m+0afB/0ucyI5W4wbpI+BFWxf4trxOUb5XJeG+lGGEQWL
8QZIcUYHA/VlhbfMTbQiPPD6TlE7d2IbkbUMapB+yGjSNfLuswhL7Y+wO/XsCJrM
TkaIlrqL9FoLKmFyMu6Fx1yBW6AvLfiWoAS4sIuRIopflZJUMez992tu+Lozayns
2b3zqnBD7W/KJQJmHPtSoLODV6IGKpMkVRuf5IWSpAk7drhhZV4mripvPHE91ljf
flhg9DZmGajumPPBNwRHfYIH6S0H8CMfYRmVOmk8aH+7kncUNE9H57sPqAxjqBml
JrqHQ7/q9Zsu8SrLQbQXVL/5ODbV+mWif/8+Bwkpdb8xwzNAQ+KGjSw2/za+uMZe
WFCelr4kBLHKsrrfiJmedrCY/2qSjrDQzslyCAUecKQgrgfijZCK+KpSToT4rPCZ
nx2aBUv3qCqr8wnLICZ7IuarWSPOcqgUehM3j9ov4KL1V0FtEGcU7cSyd9GM+Ujz
+LK9rFdB9DFnPw0KgdeLRS5H1lfxM40FgG83ZECVrqGq18y0CeU6ySXClgQDmdc8
HszgPmuWTzHxTq0jzjBuat4foFtDRvFDAMFJG3iautSBSEG60etqTzyL4LxVKgQv
1Baq2pyw0zaUli3xGZLiw3qzUANaxVEvRavM2p5U0svdYCTNhzVg5pG/F/OkB2st
G/kby6fYTVFxltcuaZpBIj+vrD1+JL94+twr6RFWR221uInSx24T6Fh6A7FrB6vb
5STOynYtqAUSUKXOYhgz4klfX1h3JxAnmbfokWlL7QjUwdi9U6uWIojz/YpmYzWj
ieCzSqN2aXBzrVRFQH7wKhq6zoIW7HNCW2wyQZ5A4Mf0doIOdFfrX6m06rfiwMPW
9CWU1x6oPpDOVL4bceBKBS8UOL5SF2lVkzyKKNd8agjbDW71sWvdoMC0HSmcT8HX
6OiZZ7Eqww0iwuOtUiXRXeSmSJm4A8j//jBB028jCIq1SkhiL3/FTv1gh3Flpznu
PF0xgKaNzx5eHyRz7I4huck9GJlUWs5+5oAIuLSO5aYb9EvxphwUyVSWeQypXFWc
LQej3BkuzXXAZHnqpnQR+farcHL/Q901Yi285cRJLyPwLcBPqsTx438Ua4jTY1Iz
HnrIVhohu9ei9Noy+ZjICgEoTVsNeOZxTnwW072k8yTqaTj9NuKhECswdRHgl6t7
iS8g1szuRI3IR9/KgYGWghpNMjv6qXyY91OX20S55U99hSx+X105ADJfR832gIKS
BJTkPTvdG4nutXGOUDMUPdS9+b/oRmZsuNR+wxzZWgOvNQJWe931kjT4L5YDOAN+
hOqdL+qXMOOyPTNwoqKhRKsNw16oHG7I04XHjTPXcNuv4Dj2Fm1md0CqzNnrL5sh
/Lit1whFvf7RDgNJHogMcYchH/UIL/RzPOSspuGTpCSErBtIDriKplj44Kp5W8II
xjtup7YzappFCM6ed9h4S4fYfJvKe4POaaBq3ZO0oi2YUH+5g8Gm3EqLckt4QK8H
Wz0TfKneA8dCCdajGH8j1Ue5YmMzm0lz9NB93vL1Oy2IlC/kb5xS5ojYTtqteYZn
B/V3WsVF1nXKnQrvh44jCTq+7E/1Qx/M6HdZFg4wqfapk8A77Q6ISM1TQjb9YS9k
TmRmI3J8RvM6EcyJuDtRUNk8Isb7k0me8ggmLxbX3Pr2vcoasvzpZuAYOxrLP1v5
d4fqC4gvjGDJ3NLfIhlqs3vSjIawYt/W1QyB+durTwD2LikbrFiCONsMABEHE5lx
0AGfSu6Kwlm/91YPcP80it4UoiGE4z0cwvS77Tg8SRw2tACWAzMA7qJFSqvSopLA
402DWEu4/lI2hhTnPtRTsS8y4HylAQgrV/n098u5cDngubuWB2UVkWjK9ZZjSdgu
N7g0hr65/dgM5SQ+No1+LlTPoHZl7s372BxbqBqAH8AcJICsWA3QNyPCUNZ3jLfX
Cw9Fw4n07uzxpLaFv+hoaNDLjmnmVdzSlctvOIIwSsLPUzM4vU7JdFhtuGDyzdxQ
ye+8fKCKo7xroo1AK6uOdu4YyIBPjWUkn364TD8MFPwV+t5OWB7jiPQG/ixTyt74
9ESf0koCyzyrymCaEPn5QmOwluto2+VU3heMsmtbKUWuCg8JmaI1fWUvPKYKVDPF
BvGbhuQdFLKbXZPcp4ax9gDSLBqCDEj2bhqu9vglLNuG3Hn3Ve2yoQc/xB+B+wsW
cDiD0QX2dZv6GyEB0YlZN2NFJlf+5+BATGo0oujoenmDnWwx+zhbnilU/GXeZvDC
Z+2aJtrfYgo9IbOS8o80nn4T4wkAiBdO1cwCx3XdiCNkwF/LUP50DnDZYJe0kIpy
rXjLPmciVpMIzJFR77xgUzST6T43ZrwBveIihX7BrBUnrl9RbkEuDoASaaRLt1lB
QraPquGicK3ipW44Twjeuy95nitowaJQ6YQEumGfYOuoj4t2FGFRtp+KN++6WXgA
oxf9SjLNgU6cAhie0gq/w2GuZvWWht5P2c6JGKmFmUJRAOc1P60XQUDmPpiZCt/Y
Zd735ecTsiBFZAeiQ1dKa1dEuTpDw6T/oCHEu2Xgc5UtGcdOIVExcwimeQxFPnR3
jZGWnXqxn8v8VDNBT9wpS69t/ZwBeriiS59fr3S4PX2ogKakJdF5TbPgNdQ/R+NR
05GqBndRxQkHr3iFI/a2DzkYMfmoZK/lx/zoxY25NojQr1kwTlpg55WroCW3I2uE
8kj7QgvwBWcf+sYpg33kgjm/sKZG+fTnWK7KKv1FlafO1RAI0I3HglKVHHEsbmvc
9JrPXQKQq/IS0ybzCwdkKgk4buAR+9oFuRKQZTxQXT7VfaUgX+Gi3SojNpULtTvQ
A2nIHTYW6uSxwXYDGTxxqHIyB0PPnfwNy7L7d03lIbZJOj5mzREDTAClVWLjQU29
CLxO2CF0t/t8GJl5Hpf05AjRVh7md0p5N1QZQkXhs+TfHPdFDAxIudR08PANP9Yi
0Kae3HCNtQj49q4/8a0bGECfz5nmZzcHYIf4nrD5UZkPOtkhtxGHG6T3GQYGEM6H
sMldqMzzFoF2ll7LTF7BrUy4BJl5UwakBkSXvxmF9X8A8jxs52VAwhKK6iXCEncA
AZrb6LsiLp5QtEoly9SBeXwHIRhS9gryTadJVAXdLqS+iM+Z4iwMaLF5O9OmMjNI
y5hUny3quWtSOWdEZebew0B8W1E2c1tORVyBruMngd4oUMV3LRIg+TKIAdQQQfWb
ev8I6byQR/bBag1u/pGzYkRG/2MML4LMiyY4Fj1oOn58nH99y1gi9NxCfmtz2XLB
LDpPML4O0hZsOhasc/VH8Enb4UJP5BcvDIn/2S6aUfwvzVjnzyVFgNrtA9ClS610
PUedwJLyLR70wZYjq88o8HM9LBfsmW0qFPRep+Cgz5psb6g3dk7ciyqwLftMEPf/
ZCvWBEWKksBQiQS8sUReJJe8ps/HRQIsle12tx8PEuSkzq6wFXvG6AsmjhbSGJyK
XpjUZgN+DdntqVxb9Kjpk2+GQJ/FYj0rS9UpGM7NRAxmIbrWINeDy4P2IfH/KwQB
1LeaujV4KiLmi24N1wwDw8aZs1EKR+QXHdCyfjU64STBlWVrL2TwbK4oUY5NbDfL
JLGN7mvElNgii1/IP/AQB2UiWf+jjBR2Tl3LoozBqtYXQXcbO3iB88u3d+cHwBdx
q4pO28cVYH6U4z1J2KTNwMcQMQOfAd+oA+0UKjwEQaA5J+eoyfGpGcTITZ5ZyXy3
XjGDohjbz+eLnaQgqDGqPlclZxyFlimnh/G1JHOD3zCNDFh8J/v2MDLQbXSySmEk
As5jh7vMVosAa2HhmeMszTRtt6RHv/OtVnlPRiaop+ZdmdI/Lr8nWtX+IDtjnF0i
m1F/tM2z4UumNB9YICij2+ioFb69uX2zX70Ub9sX0ZrQuCpJGsDO8JzOwm6YbaDm
AzD8q9SdU0nqJ5tk9wU4h+omU/KjOV39f+Lt+Obfrti4FSNN7S1u2nf6CdcdDY4v
TVwLqnjIkkihCIls/EbAqNfFHv7i5VHBEg7j+RqMfQojfxJYyHZZlJDjM3UAVGdM
BB0+DQW3wFcyFTjATBhOttRHW6vCOWRjUCS8THzun1sLocS3v3LDGJXWqPe9iUU5
vUbcsZ2EtoL9/RQCqCj9mw4s15h4h4x4GQ16mbQ/3or+GqUetqBfUlBkNZr0SPW3
VvUSsh038ybYgaeEGrB/AYntIgwTxLF6N6cS8zQpHM08eH7xb1JXMuogjsRMSXIW
d+yvwnwi+AGj/SJbxJpzieq3aM5T3iAh93W3bVid32ixzzvpdTQi8lXFTQMqYA4k
PLz9ty+l2zbaRpNV2HTYVkDDGvBsYYajGklj6jb8oF8QK8goXYcxuCqF6JjQNwCV
bWUPRtniL2Qap9NCcjxCinxWXkF587VFaIixbgX9k142cpkoA6w9xiUVnzDtrGH2
0S8wruq8kdYyNOvYEhkuMgLgTMHtasALqWK2EB8U9/ecg76dmyTHcZ8xnzvipP2N
cCWjcMdLgL+DOLHXqK0bxkU0fS/TlHDU9SV1UoZtqFk9zmeba8bK1vZe561+ZGxi
+0LMy8QeRI9+sWxQaAGRsoD9KOQDFzrYd7R60bw0QIduC+3Fxd8DkWT0LwM6CYqt
A0Kcu6IUSyvbOItn3a+ExxSm9xpxwHGgVRi/uS0cKT9Z3xaQ3k/ccEJ8ZyNGrWhA
pXZaqOlM8gf3lAFJr8XMs498JaGsv1dnTLY2HfQGl0fSoWFttb6SxP7PsUec4M6B
p+qHwy6+UxbR6hdzmEFyKYFiGtKjT4l3VPp927ZkWOU6Yk2tsJKdREFAXwvrz5Uf
dnEpz7lW2aOwGRXeADOZdXQtKwo5hXXQwDQOtkuhRm3WTQDNkQChwM0/+CvSydAq
MheoHcR6C3/R7QWS6NReVOzu2pHwqp6lAig73LqSxsu3jHTnI9iHJ/8Xa89pZIuX
aC4H79tIssCoKiSkgaE+tVgwEjWtvDgosYtfocIVtZnCXjKWX0GtUkLvoiX44a/o
pQHxm0yUcoKhHuKbh/E0+iB07ZoHPKGkmPuoizeofUIgfzSAR7JIz+6sn5SoledG
jDB87BxA1w0so2LSg/hJl1GDjVkZG4y7LDdlzJtnmc0+WBDP/zpRxtlrsDNxz8Sj
6fXCRUhMoRsY9mlLrK6+ehd8O9J6trUzHfduxw+n1fDEe/scA9++hFJ6md8rl28h
aPkdGCJaFwubaZnb9JygPWTACUdkHk7NtUkqGLqlbDlraynW4skE+IGVz10u/vKr
wDAxGkoJ45h6ZOlHnZz6xb2ykFVxSgnLPSUnIJ5mKQobRwR8ktd1EmCymY2CRNc/
1i7X43iMthSFOQega9r57sB6A7pFW7+bf2G0GF4ya7oecdGUFQvtdPFhy9gMPVGI
5zYvPbevP9TfTlsImt/74wTGFZmvhzeGeR7suLva/63zEvzj1W1FpZ2ssOLAkRTe
O2ibNTqvl3+mvGM7O+Umg5Oa375BzC4zyLnbbd5s1jKDTF5xvG7LMtPfS89iBf/y
dschWjYrRKl74QFwgeHiegUDJfLmVMQMNgMba54SI0LW8fdxkrGm5PcNoq5Gf4KQ
RGuwYFjedwmRepieAWbAhOYX1BkJmhe8PrfVTXMdI084TUkEGiDc10mA4TXy3GKW
ElhKD1BmKzRaqNI/jWcveWbK3hnPioidxwAGz71W1MwItUq2roPfPuMzvA+Rpmh9
77Ks5bhmihIoHlHmpHsGUAt+EI/O8pavVd/jYsMa4eGmkwMJVi6GB70ZQ8rqbfQr
hCgbos3A4f9bZ7Fap5wu87tcKhqrN2SE1zpYLWLWiTOTN5eXSEjjm31MXTJzLaIS
4kA8vxZTgW0MPTnKFmEFy8B7pc28C/BrNqcyDh3yP1fk5mmJmDu/LF+FmWLZgPFx
UaLcxjJE+f1H437ZcagWJtG1fuzoW1XAbV2EaRexz8AJ+jeEYT0k33ccRdbvIA5Y
duy3wKMRAOe9eeEusW7R4DS2wys7BF9yuiNLiMPKonwVBrSPc0QIJh9MF6y5MAsl
TDTkLM3SCU+A1ZZPRyoGimxzipFoutdVkzUGFxWwdg6Zji+DtU4xAX4TxMhAu6ct
HPZMj0cAlPpKhF6ReeOuh83gAjeT5JoJwtPBRI15xuRzRX4YHIt4cEvvrR0wZ9T3
9cvL6n+AlIhSqSkgGpsmfBPLq2dM8ci7QujK1/d1gBMXDv1CNMoXuP1NpbhsVORr
5IbdocCK2G/jjCWhf7doZixLMeP8vvsexBlJBTyBteZfB07bX0ApdI/ptI8rtrd6
IBOT5ULyXMiyDaJZDeA0gsRUOmF/vmfQ4F9DHck2fH/IqMZg36YHI52md6FDwodk
eT5mpRBVB9rFRgE6NlrH2dR69Az+17KXDftIgVGhy/DsU1U4duDFETpPrSdO6jxg
cT0VO7uCFIPhBHF7Lyx/FPm7UaE/dsVa0D0mm9C3YDQna4yF6pfqAOHnF+S1gsRD
LOPuzdv8U+R+0IqGpNxXD8u1vZxD3DKlkS8vB7/XiyDsUkR4As3kCV3F0uWqFoLf
//ihgL7c1Ud8m//zS73yYo5wtIPmXZKSEvg/U0QI1kZGfDvPDaubTBiFlVrCWl9w
/y2gIwBVJS3w8tv9IuTAhQztyzAOpGtlwuoPRZjwYXKah/xmeQkns6/7QoXZ93av
Xtd1kGpBhr6KLozxXP3LvhhhH4mWo9vTuvYuOO+Hn5lXdlBZ1xvYghDyK+Y9MK+p
ZlfdcThOFCq5r6sPXJtYo7FEkwCRvfkSsVgJ12J+ek+WPSCQFZBe1rqEdXjQP0UW
CDvYWuGaRFNVLLzvTktq9VZy3Rr6pWLd8FbJSxTKAkpSSRiwWO33m7Deb/STwc5Z
xiTRAEhvvqDry4jn9Ib6TZgfK3D1/3ark7aZ8hXi3N08prn+HF8NlXPV3WqQk/Xv
6KJFg1lya3LpYAnYno18aqXehaD29aW1q2jrbjUieW1bU06jTLXo+ETp20SOMlrv
/1fUKtNCtPJZLDxe96vDMGLKKKE1HbNf4qMNm/NqX7Xhl1V0SFDnT9w42t1NiRwS
6D4EHj8qvuxjMkh+5dQEbu+WHdVPHVKzzSk7shTIR8E2SPu0smJ1+7ld77AQyeT+
Wc53NCaAGMpsydxIyd8PQ8FzhIMsF4Ozhst/MsUJDcxg06/IkCpvxfm3rpXL0kgV
Doyts5lNtisXlU86recuNwRGbUNCB7fWaoYXsiG+1E1mNJpcv0/8sFOR0sVoWzb/
1GmZ3j9rAVGE6NT78agj311RxVoLSSm7E0iN7jCE1avP7wXd39E0sMv8kZU5qFuK
uT9Y4vl8MDOjj+tEd5L3TwOs7ApkE5u+/cuKEQXCZhWqjbzjb3HqEV+PLVc6Deog
mWRoRC3H+/zCH1HIfGjkrJWP1JACtbzqdb/ZkkrivsLCdQKmoc/RaYnOsu3hJNlB
bnATYV8d7rpThj5Nrc1AavU5sRAHRNABvAwuzsk6ca+fXqgtj4Nge4Dj/thoJfCn
uJwAbCeKkaTThC62ssTkXjNCp2GVJmuJYoiGVosykqyzG/Ns4OOnGhQOyVWtEYrK
wALEmiCvbVJLxn5BtH3CcvDj9jC/4oxxx/KTF78E1nvUV53WDCMZTgsxTPng47mm
C3ZohkmLDfvXSZkYM31bjjT13IgvK378hAyfP04umjxqG1OKsWtGwFjLJs5GESSt
e43AkxA25J+IqVactB4u6nJDpHXJ/4P1c+Eqtq/Gj/dt2ITlRtZGdmauw0NwswIE
rW8KKztuNwyTH5cRCVe4Q/Y1dgiYyzQzXXeib097UoBASZkKgBa33EB1P5zdYmml
k03ylUOUl9TIgA/UtHonMaVebwFOVwZmVh9HF6cwAkNoPW9n9z0Ne+c33UrV+nx+
A8ggIYKyWB4MsqwkyIMUJUlVQtwnwf23Jiiqi4LFuqB1xdHx4T/BFkl+5LxzZQJn
9Lk+aDWBUubbXFxo/LKJiKT6sHxblD8CIhIPeGLNA63XS21Yf8wQHhMxP82P00Zq
oxqanSfm4jwq8AzUJhuyknTmFdU2TYnBVv8Af2odjRdSRKcpxwgsxXlVYyz11lgW
zoT0wGdJqYkXLk7VtqK9FhRv7EUU4REkh1NJwRBXJjHDWgEAYbL3my8OpvXnkblf
tyaRIBeZLRklv6byLr9lscWlqMdHWq68nvxMWxJp96KxVbQR7mKnudUQhuKkXFpD
5PLLbA10Cdd+wN3IaUn3W0TidXyMqEl83KHp6cBU1Z5yhcB8StmL3RW+z0Zoytkd
ilwe5FbeRtS2U2oWp+e+q40UrGNrlG+EC8Ys48gxXnLAH2XXGGG9TcaBoi7uklU9
o/AlpoL4MX2y6IukguwUyYZThh+uujqrjWa3PjX9AQMRXTF4/TxNHsscqwUatYPq
u8Z5Nsj6ERdjWhYEIlTgcNNrMrqg0RyBuf/jHXg6Ms6gWL2ir6pdfSehZAnP3c2S
w+x+PGaBiTLqgv9pJP9p083pyYikLm3gMISHDWX7le/4stiVwCSq7nSrIvqI18ep
GL1B/qrvk9ibTbOXBFt7JBX4vKZqvjyS6QOJARd0OPhJfFfmAc8edfBzKFbpreKy
LTxJy+W1E4cP0rL0ECGEACx7LbY/dBEFd2wPfLa2rigB+yh8AymrJMKjYr7bIQMX
9sflw2tWP+wmAVSfHZdiYhJvbhYMbCiJVIny9+YRkhwFCk2s56v4iB8+qbBlJiq/
eqlRlCO44qiQZHuA0AQk8HFgU2vhYHD1+HAo8ILe/O7Q6fVg53LKUHfZlH+sjSK2
6kzC4SzIyyHrmlgBbXQSHXAUfkrrL6PIs2802p6gssXB8R+a+RLp3kpcWPKzno2d
HRxjUukg5MtYnqX/l3i28tU67ig/EjfGDVQecX0Mbx8PX+k+fr1CVLsqqPE6ao8+
SlhvCzdKDV/ZRaY3adNgDgkVgMPLhMKYAsugNMs4Ajjmc49SCAD17nYXM667MiAl
eS0rxAh5nIvud3dm9KGfs1R87uqvDaCVAYI7hHK3B7kJ1mqHE0H/WWyiFUkDNOhu
sP7L081b4dif53fu0nCPBXsGwuCMJFZssUOwVoMlpG70Z5YUYVO8W0JAF+EF7FXD
M2S/9BOwDQy1N5Tsk3D0ahJF5VUnlZjqtjtVY1oMcNppb+JX3pfmjUrXpuejJm3d
Y1ccH9qEZufv2ot8x0a/OXraJSRQZEmpDsKd8zc9YHnMT+XPnhSzxoZgvZta1umX
vkZmnjrN5vakEaD7zcJkn80FvRQcloTV7Ry3PYKm/owv6d5WrNeRMT2KuCmJ/qoP
DbpNssRjmohM7I3XSaPMRgTFOAG/dVXmAzGcFFEBWTq6WWk+lcGGBF8W5NpzLTJu
TPiJmbK5YNIQyGHh1dc7wj4XT3yBDrV0D7XRovhjtxpIPakRD+2F4JTf+kZYd3wB
LAZ4Vfgnet2SOFfDacHzt33qE2xLkx9UsdDJ5jpAJOTkxUxGm2y0nGildvHgeFvS
2KMLnHzW9r2kNi3ACcvciCIIaQ4GKS5p2VpI3N3pDovxySBVE2DyLPMl6UgZpVB4
jaX5ouNBNwrsxaZDHqUaqbPoOKZQeoj0uhFC6Qu4qb2i/41illgyU2BgFKfwy96I
DHzlQbevkCgYFFRf0ZqKekF2ioFAwCleM89UDyzc51XcGF7HbVyOaYrw1WayuVLC
qc25ebO/mBRlHf3h6/myfzCZHNzg2b43XDOcpqwfXNaaUK8nCDZukQKax29GVWsn
BUnFiFxu17Lw1T+FuFM76/dcN0pjpyopVSNCnm4c4fGOYIhscDX+eVAH7i0OBkNq
LxO9zNjlmk6MQNWVbIZ11M2tDpRfjscQjrn9FgDK7ycRQbhVD9RpG1gHYj4FiKQF
H+4vqDkf2XJhHkAB6OhKyMDuBDs99i6mljvXS/jwV9WTSnVBr/DXlAapw+t4sWTs
sSPcYttqrA1wsg3LA5LoMYT9paJRtafS2ZUuwGT2MrtFUG8zVV2PrEo3GCPy3t3f
OphdmzEqhjVpe8Vo8crrkYlnynKZMqdubWEHCgkC0enNAfG4/nGvxE8lt9Drwnnw
kO4Iw+/jBizYiUKd+VPlM4tTrj0dLA8u3Tvoq++BMcw7/6tRyddKkRGdV9J5CH5W
ACqM5os9O3h8lahxck8x7BsOC7YIRYo9cwXRoy7oJ9BfgvcSu7zDs6gBpHCeLNNA
sZnideyK4sfgFnkQlEqrjtB/dd1WXOYX/ReHlgMneA/a7SWPyay+XBSm6pjtxgLd
Hjm3Es9Vp1pnxZ538PufrdaD3YTYfxZmafqRpkGUa692p6bNDsRFo7P5+RlnmOzN
fjEOPc6fzaW6F2kWYwVRiEZ6g8xbEorA6HoxAv/l4eyCUinwQgLYT8rTUha59rii
twERd5o1R6S1qes/SVJnasHWQy4xYEE02luISXqhzqCSIQwoBe3wdG3RWAssici1
rxEIFGSH3ZGittc6AqmqzBTnieZAXYcN0zmfUb0puge/GDxwP7+EutHkl3hDv8dV
Rhq/3oJOLCPsVw2zz/3JezT7eXbP0Gb/1+zoKLziWhMfViAOOP2t//F2fjCyqjzV
k4+ejOi2hp3ImwpIN9lPgc7H6MreaJBtwnHkyJhRvFQ+FPpdjZvg4FKX8zWBIaSK
FZbVWm0UwkWLMxfmsCl8DJteH0QCDjdMB9X9ekJi0PP7H0aXSwjZFIFKO3wsGJNi
canex67Y6oAjqL1+LayHp4a3zNzfyFxgxkInkFT1y2PR5+e17heacgXcmZHtvxsg
Xn5NmemSk/FHCR0UnXGeyoUJP8xU525orYXJX9RRKavJkQyn5FKINt4fuHZDrqTT
cxm3n1ldXfcgYw94EMdPtInENxAqLv6ENbDHnuFc+bJNg8Rnt66WeEg6lU87fhTc
26z/97YZ4JJKuziNTNhFTzXa2Hu4ztH6iDEL27nYhwG3rdOd+iRxg9wofpPGsKPi
1Dhg/31Pqi38a89PpLaPfnpsxbmn5p72cZG/yoHRBkXLeIK13MHHt95yq+33iHj6
8YhTyu3GCF7ij5WsmPlI9Vqm4qKSnPGky4IWux1LI1WJLB1asMkapl9JJa3j7h91
UPol392/WtzAz2WC0qHyEYspUOAgJWfZ1JqA5a6nSg3vosPoFSkCL6AqX12TBRDt
xP1ljMJrc46pvzH4TSKqUcJD9HrOsekw/1wBFzl0x8sEhP+6DF6G81OE/iML6hRa
0JQqqAkLpjfmFefd3FeiA7nLU9lSPsiH4Iz8JXfA8iat5b5pSJDhsiRNSJX2RCdd
f5CiS8yyaJHQXf2E0RIYTaaj4KGKt3apBNk8gwGC6XT3KCgw/cA7bjY66lB0nrB0
CPk/AqONAwuIvlwNFI32solePH5z0UmOkZMPnEYQ2i1qEhzAguQsMViLaW8mwHmq
ZGsNvsU4Xe25fWpozs2vmlkJqLx9AIxR484eVCp8rDUA+/aga+x6keIgn07e4e/3
5eZUX/sCCsVPlm85f1pkl0l/agED421xNajio8ZsWRtn6mnVZFw8WS9E9yMkk6Sq
TIrli2mBroGnTY9j+B/GrwAVVfWWS5jKIKRMbQLs5Iu/glIOUI42HYGMFJYi9mYb
KXy7Qfvlxb8BU5l/54sc1LuiCv6w/ImNtUnaQy466NsGYe7tms23eMwCKgB9IO0S
U6TXChxpATm237TsaZxX6KZgiUeLfJg+AcKNshF/oJMgIDGsKpMfLxd+1NIy4Q/4
qThkMzfmdZzclnDoZL/DFgne5eq1A69bWOqskCJtHKaCSKmtKeaAoAEYMzI1+SAA
edmmlwBvO9dV9eeOEha7r+maeIrn196tyigyr/GNwelxp2W4vU3cXIpi9ODIxYWd
C+HvKBsYE/h/5L/lSj8RlQT/IYPQxW8LYbHkm5YhQ8R62GKWMfXdTt3sovVxsTGT
EzMhYlWf/A4ReshrCg0sNmme3M+SDnS3rZJFcwMdVTDvi6iBxR8kQOSDk1ScyFWC
Csvv8i5HpUogV9dpIdoH6kHE8TvVoFxvIF2SUkx5ljAu0X06hdSVFeJibj/E1pha
LYmzjpXAJDH69ZzG0U+TRTDlBiXp9vQKUlZ+RlFTytBG1cKonzkEuknSLyIf22Du
ebhyyF667xB6et8GDCO9i0c1ldov7elMiqED4lKukAbRlN39O2zzLLKE9/Ih4wZx
d36OnHXJ0V3spWJ9jnnBi3IhewfWhn7ujJpOgrJ5sUm4K89G/yxuD+MKC0wnMx59
Gry2p1yXf4M/1SJdlfJ1haHGSkgoLpwvl4xXooyZ7EkGOFpvVm/xfV0l1oxC9YE4
0Zrmy7Zl7x3teMhTLlclCIxRoimNyhMzEcilZsmFQIbtVAFtlXFMztRQvvq7RTrV
1kwdMpkn1LXIXgUnnDTqv0le1BwIcExBaV9I0+UyDKlZ5NEG1ssHHNHLZu7/ZzVh
TzZXTawkpMvphG0Bw+FEaSLKrxAoZ9KopytgtJWIQe12hggKIjrNBWq90CuMtfFu
gbNlSaOd5BidTd3wHPUPkCUzzdziV3Jr2kikbKZv+i8KQxiHIn/o7XpTspOU6/MY
BHlyBKf6UrvJAVuRj3uCv+CkDRNH0xlaxICl/uE/GztdciJ5F7nKWsdmpz6DpVRv
oaNGxHHmlPMySxeHLYawX5FPSdFQyWjgpUkezAb6m0+7IujRhvndWcCXwKLlZ+41
VzAKLU/5MEXEeuNfDkVcQKfbPfI1Pm/d+A058nqKGCJnrN6XVBAhY4sPWwtlFW95
1NfZaNPh72UYYyXF8D7gEbKiH39lT+3QEJs9enOBuK+E/BmBF+J/jDnlfq8solkI
ARwhNtaT7Y/wkSO9oT6ORCBL5D6UUH+dqsgPntUdmUOpNafKx1QQ7orXkBP46BFK
IUJA79ny2FzVg/wW+T4Q3+vMRDKR7XtXjua4Ln5OPM4pSGobl5lz+UZ1d5ZpUOeY
fb16pPO7DrmrJyq4rMNQPAku1ERAnQDn2w//s/X4MMhKYbXGLde3Wy0fY0PlsrVf
evv80wbJOdXhIp8hDOgyx62FFiO7oMhxLXJrCJcn4eJGTCFk8JQ5wqK6JB7bhs0a
8FOlOeIHr1B4AobntS70O+SXvY+w6Zt3ptBhtb7uT8s+7WPqyy4YN4vUJG+tFsEJ
LArqHWLg8WkjwtPtF7b4R4zvySyvlNxsn8l783Rx0bsWA8iSRwLDMbwauHycFkPk
X4Y3qukig/Z5tIxx3OQbIyQS5tce8SC1BTR4jF9R+vrXwqbfNyGU2L9EedNwQ2GJ
BfD3Clu7WnLmVJ7PzFSJv52n/Y6PZkufsZSK+juAbSJ6ig+Yc+V4M3jGQDUz4Y9j
MaUTY/dqimMN+fOgRs0CV3JLc7jJCTBqjbgEY/wrrX2bu+xAAVe8tZxp0p55UlvL
hICptA14ePXarf4HeUD93wiW7Eb0X5pJGbFisQMJLEcFYWQnbP1SFXeMK2iDPz6S
pEqH9JlTc/ljcAn/9tq6I02Z3JbsEIIixdYcbINs6S+gZuEnYp8b9Me0vZUv6tnl
9OdcxMi0bLxkc4FbyKlchtpXi+EX/6DvS9JAWPgcEs/tjojNDuBj6EEMDNhxyDZ8
RYepUMdChZswSgQLZH7H204FkeGr2yVHfR1LvxPhRi0p+raBxBA5XC/3cPlQyz/W
kjKiXy4fiFi5tqnpovZuadZfnTeyshwgWpIQTdYeY1WUo6sMfvkbf/8hwe8gajg2
F1w2FUYOQweJhEglDxGQEeLCV+ZRkwgK/Wmn1hk6gRMKvviLRTRYfvT5+F2cFoFU
GDUmYn74Rg8bOjSbiNHH7v/fPA8DT3ajCo15d5ukiwia5eFR7VkHIfi+rJ+HcQTp
HtvHG+cmsvOBdJg9V//mW/SfK3tMQoos4l9KF1owSlB37gVjZlJURoSgt/jpwN0k
HuhpjFkbsPNnZDP1g1MD+/nRs6rr/nqD7OYXTOCyECXlAAaUOz7onfQeOvU7RLVF
odckNmKFN2SsQr7+lCcV9iI3vbsXsFbMG7lwJQi0khAnsNrPONs2uncODFCN9pix
kNUWQ63DAKxtD/NaumJWp89+6eb2amVNhhSSEsXEepki+Kpl0am7CUPQguu/mNN7
dQB5pZ/HLlBZJSkkdRrc8YN9nJdb8SUgfNztveg5RXobQGz3h3LHAlKhWcrdrCDd
LsRnOEFZ6PShp2iYl5M6mjyY+gX3rrcr2nHpap1py78z43ud7Z/0xeQTBUiFKiJ6
yOL23qzrt0x1uMf5Ovlgjngq6vm+WaWh3iynWunONGZcgP5SMuldXR8TpD0fVnqz
8/jidqjHdzakaHjFXSo1sF3i6lxmehefEzffq8u5YcDkKaXiFE/dgH3Mnfxc1Rii
CATe512RK1aEYDgka09k9IJaadxFjjaA4mxcMo+lv4jIh0fppDW7N8Vu1+lySrca
UYR1n7zK0dBZsq/PNYKuoRqHJgHhTgl+SbGEVmhbe9s6IDeRmHYWD2Mk10q9eM26
ERZZIQ+CShnQcesjaykUnBRh+w/rnWKyWDls3vzjEi0LtK0Ie0ndYGJtZhNtW3rS
jS5PxHcgOtprWdVQWv8jTzQeacvA991+f+FzdbHh0FIZ+VWmXC/9htvK9IEtFMv1
twaHlxXg8DKb02vEy8Vl2C+cdzGV6HEMWOGVS4QazQTY2a6IL0ZcJQXA6FIF+LsY
3ajQVha4SQiGhlPVtpYqSLgLU6iG49advXRVx22m7WXd1BemipB+hSgupyS2JLo9
pvstmdmhNag4k/QTk7Mr9hR6PlvdsEccXxo4D1OL1TIpJkhj6ywWtuvAPH8ToCxV
tPBhdCIWKAD829lVCZ/FcI2Z86nDC0TIguA3gXYmxoOii4ra1k5KDwzxgcTmH4Vl
2cCYE7W8NTB4v63+dxTeZOt2wHZ7DZ33V1lNlcw07ZdCFfqnh8hsW2FLnrqaK9j5
4hxwMvp2wYV22Am5nk5l8AqJeda7yApWvUmlrc+nOkc6VdjnASV0DUnDdimTPT2h
6Xek5E1qXBdatJ08EfADFYYz7YWnBEyGci1ZGAuYB7GI/JU8BkSTWiwFU+egEjcX
ZtXcvwdwL6z1uKklVrW9vhKuOBAPE3RRTfKdPM2LDQr3iWCPnKzgUKt34TZIyj2W
6StK9MekjrvAd7JthpozqhNTkp8W/8T1hCsYBXA1SxRHiGFYO4Aq85NI1DoTuJOY
ljk1OxjlsgGKnfYXcnPy3rz6+2QZs/HcaKlW+1uRnD7cn915OcbMMF0iJ8kr9Lg5
l7J9ztyqOjJMT1Zg+2PBoOfXQ9WIZFzc6InnoFRExps10L8EuM8He5mxCNUYgAFc
mu2pNxyDCxKX6au8b+gARUJkmPWrMnE0q/Ovf8dJewcRYIvJ3WsRviBqW/qUaR8U
ibv9H7u1Pa7U5oc1hRfPxjn5RNwGlcHPnGD8uihFy6/JnWoUXB1mTtuOYZKgEulX
MVdOahIKbfIiEtk69iRbDdE6z4rkuJFIAUbDbMpugWmX8oywYJB/E8DiIR7j4MHD
yoTFg6r2flnvM+vjRZTAvekXNZpl2/6AimaMToQXf783V4BTdndm1iHB8nV1aK0P
PpDAa8x/KfVjsA6FW5Vp6to2zr1b7IgOvvFJFIVjmKCaw1Am/CI31VihPoIB0soo
BckJiu/3Cs8GaFF2nlsY4oSAcS8eNTcIa3fVV5fFbwB/8EoSqFjIZokD/774cm93
2sTiEdU85JY4UoaQB3b2N0LKNH6QZ4Q7yiS47o3qUFgCR6vRM44mFCG1xHWUMFNt
YgrdnodYB9O3nDrl9/6I0vwj2KvYCWoDrOTyJAKm6lQWcGcYX4THjkaKylxb1cCB
+acUBuU636wNYiskGYBhxxOV1b1o7nep/CUC9eQ/wysXupG7vKj97nR8UJcY6jPF
5cnAOmFBwGKxf+4AcuKkE07i0X/wbl/TCk0S+IOOkRDNjFL6iSi35Nf2RW2a1kgn
LZEfEXg6SuGaMNxN3qDzqyppFTovwg7grNLuoI0oaSz5trBOrK9kWuiMMGs4Z+Uw
HWdBgvWLVhhBAc7seAa04Vimp7cR9GOJt9jK96Xln9BzGr2fj+AvUh4doSqT/gjc
OcaweUqGwQIlE/jXAXwC1aC6i49r5Z/QksJhCbCG5Vd02dZ9jtxhQrHLye1lzCXA
ZqVJuG5Hmdy329hAHShwWsdiZYDAGeXRCe+18VjWpwpzFPE5JU8jg0qIsHr2Gjxg
H+xV9DFX9F2O/HHcb8N0S0DOCLH6MiHbZXxADhnhaZE0HEJ2g0BiK5BL/Erkb/pV
OjAhe5cooLdiqT7dKwgJDBFqj5NsRPZ1qAsRVQc1M+zEv5mn5qNVTP5OJfQ0UPrK
YAS0aJ7jA9GYqCZhOHak0IkiWe/E+927OLTki/unpdRMzDM4ZtSdCsNJCCD1jAMN
OXcqM/PFUh4IN5+QdJA4pBgZEPnS7td1KdBvcBpRLyhBRkxXRY3UdPKn1MBI/kPz
XTKaGIbA9VNa+SmbGAwQ4pfszhXDWkgofY1uRXOXhf4nOcEsvsPz/EScREhHbqmj
OL2M2WE5pKGQjCbd3G37TXR7ikPl1adWeMX1oqJf7+5FR0C98LB/73BqfchZEySf
Pvp32bYYM2i4p0o1mKOrfO1IbgA9dC3Eusi75vXdIRoX449pU5BbOKc27c9s8mE8
Wq/JL7q17TpjjdS78wMdGsvKKRtmu0Aifsr0zbANVj76fEEyKjwT4gg4Cu5ZDCt7
CQgdK7TWHALnFApWmKxtYA7Cvw0VXI84COclqSQR9NKICp/s1yLTWHWmAUEb/ON4
r391zhZKYeBLR4GH1sAuwkveLV/ASoKvCgUsZmwM764UKg7ElJXLsn13uGBfz/P8
vP3ucbpb2wbI3Ooe1E6r1pDUNpZ6cxrrcRYGyv6cxup4z9VPFDMSXHxBFU2FwRG6
3vdto1EpbEYr6f55VA21DSyy2zY863rI3rjuBs/jlBVAwkGGmPwlN7c8Bc+WT8jD
HymYkFkyNFhd/hyqivo9gr/z6mkb3wqPhKfRwuY0ICdsR2QcjLm0SDv/ZN9A0OWu
bIwbpgufAKD0WP4rCmt/LK+RjQpnQosOHykOuFxdu9ALn51hNMCA3x67q/Ijy77g
SjUR4ScS47b+ZCAE2LvfYLAzc+btmwfDkQEL6oqaCJvDLfr5CAte3pvvtd9PSMto
jbnziSJDrSUNE+pXrTrD5RA9Aq08+ER8nLBtHugOlKkjoDXNqlVyyUml0Npfkpsd
aKgbYEwKFtHrzdCdSJzbYw3Ftq/Y0X9h4UeXNBLL/NzVaBaznDZULFTaj6qYnTCP
IeYwulxnqTTn/wxTeBu7ZnV1FZQBoKTpZxvzwa2aZwZHzajWxILwahEuq+nX2dGo
V5FksQTULO2Adrd0KTSeo3zhBOFpEdvEkYIq1tBzVYcHHgZP8f60N1wgrj3aYckg
p/U53h3eD5D4HL4H60eViRqFYl9CBFNaR+t2miu/UbJdmQ8nAR0OywRogS49cI2Y
Ms8chUzT/wATRVG9xyEETLcLkxDT/7dxW5yr0JngnvN70rXCQDyIXyPay1WeU4ty
HUYQ3Ik5AIV9qjDjOAtJfXAY+f4m61DoDAW0CTNRtXA3Oxq5wYg7PEuqQyMMW6me
PlFHfTT4RAHrQ8pPlZljLsStytlOL89nh5aHn/gR5zsJGWYjq/HbdRqVE4718Ze9
curppzspwJ22V7X94I/4Y4Ht15bI7+VW4oCkTaN8HkWfo+IN4sY1D0jEPObfpamD
SOOfUQI7d9WA4YaAhM96Vp+IL+RzH5qRLQa4cxwet4idKFTKV2UKDG0Tb3e6Pl66
lhc5eRToch+MgtCLuxLsP5EdCEhWGrgCgzZJK71ZM7iDUDMyohHGP93CskE76Ssy
4/KVh6G4KxS/N6wVK/VylSTHNY8ReIph/8qZfk1oqb8xx81a1fmFubDSeqNzugfP
1ogxr27AXuo7n+PyhnQ7PxVoIVEqc9jEpQSyx4AqQ9O8iVC7nhn/xAJJD++QkN3t
1eEEXlxuqu7oHNGPlPnmGAC17SdEgepm2PNrAeKZJUCDiyuUOwZ7FEuF1sn+ct8L
o4SvWj+UK3U+hRNvebB2X42I8E7e87k4OGaHFc9UEFyRz0CRtvP1zLTrDtZ4iXon
TiypGGyvLDGGhkUeMxkP4CGh1apGZVNZ/CSLEzRnD2+U4LAa/MalrlM/QKKSBqWU
7a+gO47CA7eC9ZmS6P58R0sJCM9/QVLGMHTf+l5uzgBOo7o1JuMWYLHgb2qX7tWm
FWx5//RSKVIugwHAaQj8Ux+8j5Ot09H8d4PGTvJVPIX5TfSM1lanHA75VXJKBlE9
bg3L7pezT6sVyMdOVvLF+Rq6szU/5xE9TFXOw2tI0S+bJgTTsm1xwT8X97GxnEAj
dZQZGo7rzsNohJ13NyfqeOhmewN0cHmhZiCRQLAXx3R3NMVmfu3pCJQJ7zKT52cS
PS1crIoSFJ9pGGO+TAKhNbg3SRbigNAdSnA7UvBRMi+QIuh5LMZvMLr+Y0IkOnHH
p6gafH4H9ON1qQAzWvR36xmIUnMSo6414HCYiXag2pVpM901EG6J2b47kfitDbtw
ZAzdYER8IpL9xu2pvmZrgPtQbCvqZmoqjwlZNdJ3cKloDmTQcxHbIPRxe5Im9diQ
CPFpoTM5oYE3pk2wBAPWS5gg8TPqbxuWAtnJaDMd2fb7hZsPUiCfZ/eQ9gHIjdjf
el5MYM81LHASFIRD/MLL3WDNxnVPMTrBy4woJlHb4qHrr8ohLe0ypv64OBC+pPfX
gfW2117VIEacW88l3Kn+HW7HxTMOQQy9xTgcI2+LY9mzxnsyGvhpPdpUUlcsTmeY
89Fv86gF0APvDs0UmIgkcPrZlOkdaS21LXa6uoIPNvq/Agbrj9GXvOGeHMkF53Eo
MJ/c1uJvbQqZaKWTAShK1gDfxpEUl9QtDGgZggRSareFzNVtFDoKiipDmYaqVuw4
0QC/60+6ujafw1aVejZg0LtZskguXOMKeKJAx+icRRNvj0m7mKYBxz1Nlgw+cs1E
E0FI+vDR051GSdzt+4LZWVwyR5o5otz9fUxRr/uxM0sdIibVnbW6Rlvohf6tpQM3
A8MWel5ysQFC96YrjKnkCM0GKN/TuFLOelniOjazNCf4iXM4UYby90OdhjppkVaI
2SI7j0erhq64p5ETWY/5/P0UrfhyrbhTzUDw3ZcbakzuBn4OFYSa0grXMX0AtwJQ
LhsZD0+ilSi+7hu6umiJEGamZOeIDQjLrYsO1j/kOvmvEcYiLFPH+oFQzkekc/HC
MO4b66Jp+XGCBY7vmT0x9KiJixdY5WapeCkMqub02oXCevMOlVW1eIv/JnXeM6Ws
GRc1FBuYtBrz/QE7m9vm2HhYNQ7O15G8pZgpHIZYw3mb07jp7uWC1BewL9jv2DuL
RkNGDOb/cSCqQH9pgiL0gEFuhcd4quwnMs2J5WjMOTBYJMjB1KsqN66x03SliwxU
ppDer54o8ROKPB0GdhHwvx+4LMM4wXfyL6ejhG0yjtuJArtEyU8ZC2PKNgWep9qX
kgcN4Vwy9puT8WX/4+yYAfrD6VGHXKfAMuQ0GH+gd6UVlNYf1awhk1eOEwMiN5uJ
w8Pcut+y2mAPUKF/sctwG/ae5uw9Sh0Rm5HkBQOPuy8nOJGKfh3zpkCPaYa1mZkC
DgmvIvHG7of+TjMVSI3PQhbY1d1xJBd44hQRNjoKmYhx3nRcD8M8ttqf3XS/YAYd
eSeUgB/FYyZWW6mY4NCNjCC3TQTxGxE5FLo3D46Iroz7OD1MRfKfMIgNzPWHVJQe
0FnK4airzNIze6ez8VtcLKdTP00yZut2BTK/YupI/2YeyYPXbpIOID/v0fSF1oLL
bCPf/GeYuDrdie1JHQoykA/h3CgWnHh0WUd0P+8w5BkQ6Br/4Sj3mK5dHXIJbINj
4ERFlzhNvx/GWx/hQWTM8EBl8yARenE9JTVDnt7UhaTmH/skStBJCTj4uexYrwyZ
mBCa72FcTJDK87SZYApNZfnwFQE02Vi2Y7Q9PO/tRChTj8nUwpgr918eUg75q0gM
Jl2GRRi0IjpcL1oyEN3vgZZo1XCGEpccijtHaleYGjWDLq+FJwg8BecqgljDCDqj
y+Y+Ut95Ojwo5XGUH+3djAiKMQl6HR9xg1E0CxetPro7wPdn3TOjQnRvzoW+HBV3
VpEkqX0Bl4Pan0MlKWTMZyobDL424ywOhAYnVzXp3U7F0JNwQQdOjW+0SMDXxKIh
RoFHKFrAOsYBVHrN6T02em5vASXQt9yCNj7npzW4elZBo0prJ1g2PA+CEG/JHEk1
d5WpamZbf1sktMtstZ69bp7dNtal8+U2k6D6n55DkjW2CjtBLlFTYWe968II7lNM
FSDzIRS3XpYmPOVLJvmkgIwISKgN5ZJszdwQmHrjZzIdJslDGsBPLI8ifO7k+vTn
EnGdea3BsaHfBnfPQBGjJJ9PG98A+sAVX33TIVtS65+Mze+Rr76urJuOPhURbIHw
RrujWTXgNyLXD7NH43awIFhOdhbvF9qbl9HKCamqhUkBY9gb0IZrsnkTe31zPIUE
D8OfiTb7CUxkMS/a2DbwmlE6p3+RSKlWJfBQQxyMVpyab9nuLT/ABApxuwe2iaSk
yZdIHvZxBrLEuzOwWBg7cD7uzx6nAabQj1sc0XOi0aWnOKmet805NLpD2Dnepwh9
sgn/tcrO8h2FAZxsL5FrW98LYw7u26FtEYzpftFswOJ9KWfoqgO26uBd2b80Mtdy
UtQvnUFyOxTEomZLMq1fqyUW9F3W1SxjPuZe6nGPBUyaYpBff70mhtyJt4OUxwbU
P6O62ymoHPeRsndH744+8YX9Hw2D7EgKpwt1kRmC54dwKLErqpJWANQoTJnOYYPM
Ja/bnnYcDrKjKPXXdaE93IP3ugJRniO1p6yMzIQboGzAF+nyOY7Hp2x0/2ZAoeoH
2pXQ7IP7CNCm5dGM2V8od7QoQ/aRaJOl875nKGlhM9nBEATGI48/51upspsU/Orb
JXAolcFuwgcQotFsrm5AShpfChCssTTzY+eYiRUUQpEKtKm5jr51pfqGEcCiN4K+
RJlw1Y0NwzccmYqOzo9WuD1v+uSY7p4h4Jz0Xr4A5/cLnB4zerwrgTZmx0nwEeo9
HKr/MsmxTi+s7Yhx7nyZrivGidnMs3gPSI0kPkrwOP3kdvrBxI5DgXk6RTm/TGYV
2FwZ66B1+/ru5vz4l2ZKJDaoo+zHRmEyUQPDnjW0Nm63zZfgxTFyVi0ShIIKv/yS
2zn2Z4ubTkgRqhMXJfTahrZBVmiGoAhEIPiXEpJrwnWhrGIqowrNDHdTkrocqyH5
Eev1phnT2ByRNL9jul4jkN57ss1mnA7FLmXxge32eQSfyYip+2BceT+y6wkvR/fI
vOWfTW1r6ErSX25A6ccbhcY5xfF92juzbTc6Iw1EAqJyZr02+XlPbVxGx6wCODKf
7CaOfXxcPVUudBWlnwCTQU4Fgo8lpxXr8e1uPIhYXZgvwoS0+UhCH2xNamjttWtG
xLhppY+520rZUL9ppc5pXydBVZt0spMXjZii8XtRjvR6T3Tm/lDF58BmAuFUZn6K
5DfvR8g4Xk4ulx08XwNz7DNas0do3d28iY5kk3XEEZH/HocEiRQ6nyJK9pZ7mMC7
jlf6PcM1SJRokQMYl/3eUdgAkVEV31dD2Hs1iygei6Gm9ZbHpFMhCRKoMz7nKpLp
Ot9jdPsxC6imiYgbk5wmPPc6CVpjlwbY9i5aAvoy26rQwnlzLD9FaYJeYDYa72ND
5qp7Ihhe6QRhseCZbim159LfX+9XCgEUsTeAxp1nIwfKmcuAopUlqa0kqkrR7q6c
ayNOmFRh7VIIRgR85S+vaWu60L/3ovY2YACuQIyX8DoL00/1mPmXyUrttixlGaT1
rklVAuA8q/465CSUUfeD07lbqL9Te7jx+5xxC45Jg8c8UtmUTZ5EWMxs9/5Mca7K
kmUd3oNal/qg3LyX29IIK12GB/AxnPbwApU5uPhwkldv35pruDKA1po/cT1s4C4J
BFcGHyf3dhx4EHXRnd1FSkZe7P/xmYWjHWJrEjIPxxOu3jTmVhPVne5nAKyzmEgt
O1PKMH5fbjdxyYH4hSdNUuBM/9+6HmrzYAeWuJ35cvY1taP+C5AIBYoXywKogzj7
7WKF5StLQQ8oPU4mE5rZrOPVnfYlYNkQPdVXnT2dQ3Lm1EO4rOj86exzkY9CJkaZ
Rj13mJAQrnOfLoiQmj4NWYTvji612pX67ggbvBTrZCj+eCyxLRra7Up/o4auKC2H
5UFiTXbP3W/JRk9K1/tHVTH/wqMZAGFhlML5N4aeT75fXgF/gRh57Ryhl6FXQAoS
OrcxQm3bIxYXnGQnCwGkfqahfk1b95VlYfu/BtreQo6e9iC80olGDuxpkTJ0Elru
/ojXpK+DytUgvTuakPjTsvQUJdHTaTC6SUReZKWrdtIHFolX8fKloi5V2mWMVi6H
S2ojdG8/pcGFZnFhYpwSnqFqU3LLPHebvPitdCKscq+UwPtduTnrojV3WL1J/eS2
VIBltY2TgmWbr1Q6ddTF84mTyRgiypYqo32l5c522T83I71NUaPw+1s943ZA95iY
1yXppqBpXCISj2y0ZI26VTgHaGrZbaipYISXGP6AVFWa4nr0rX7nQoHsgH4Iapmo
bLVljwpZLuCuWG2/PNbmSHLGnsd0SyfbwoLx3orK6O7nCwERw42UrbN3yDQ7lVZ5
cRq7L57oDbhdaQaBoD74fSx//pZIPeB92nVb0mfo7koCuX615Umc9CIPpyogETZM
ALrOXRlkIu/X2pNp9fZ47K5LBHbqnpe8wASWy2xuPGoJP8Pqc8/mfyeRkVtQCXqJ
0Go9RZ1QUQ9IScpgocwEnIELI6h824u3I1bBub290bmbbX8WnY8/D4SE/19p5fOX
ZqVmEO7W2bNDlgPpak7N4r/qd08+EA3p7dP1Bmpwj2fyIPb/cwPpQ6nFC5XLjFxw
lwCFlFhP5RCGgKqLK1lYeCX7rfI4U1UPVnqaiCcHLqZDtyLFXDIkgsgif46aXGyh
8o28rUVLRneW/Tv1yR8WyqpRoWcaQ4d21f2c09+aK4r0RN/AVq5DpTjU195hJN6u
hluSQNHwaTJP5a4gORIO0yuGFRURHoxQi/GrOe675qMLoA04EBd/05U72II4Dv30
A++We9xNkwcbD7KrPtXc7Esu700oyibeyoW9UGxW3ctrZONRnt/RItBnT7Cv761H
HmX07Bx0lgwJxTuhADl8dLIgCpq9GgQ2BPgKSWPSBJgn9oYAXykxy0pyJwOKG+dX
GCQ8fLO/E0Y2+eSnJEm6CU8s0cZu2zjfq8fRYrMCwlaTvdbR27y3LSGGIfL9NjPN
norMPPK0N5sSaT9SlOG1eegfc2+KQi8yeFGsxOlBrt8YvdXb8F5Yjrm3V4C6+Zd4
O6jAfGtKXTSIVlOnfxnlcMMjItr93RbBxnzGuwKXSHS2ZX/+bgCiZhx7XpeQYFGH
D94jRT0prbRia2d8Hz51JKC+oWx/lfXtaR4uLqMI0/B7stX2EsW2N2VIgipOa0Nr
HWoyH51emubxAaBVqUUk23nT2PIpvRap3HnsyvnS5SZQ0D5Y7AM+HkWJhYvxfRXM
u8E5oYmfJyo2hyR2NSodevQkmY88nYwTV7yL0h7dbhoJSko4D0gTWveYffgyK3KL
PfanlCoZdgAOivUCVJEt1uRtJ4wOYQUsOBySDRzA2NkVeE60q7/BYL+Lr98/u076
/QejEhmWEUL+D2NT9Hkk5wlZoBLfsLJX4lPwpj8B+QGoTpRMtebZYNx7xtbvJqfD
sL/nk8R8sKf6Rqb8BwdMfJPSfGNs089OqSPyz5rspHKnLCjdQtBE4Ay8LicGbmdo
8tQ8hYAjd2A2rjhxGULfJGz4z9yKwWvVH2eplXbLmo7Mpz7wgDePytHQCA6mzTfu
Hx+QztPtOA3pKq8eH2y3+VnUULwMV+Qx16H44A2qxaeY8bpe0WtaCDvaQurX8mSk
fZ0GV9xRm4AewRSqrIKQ4aXBQ9+mInUW9YcSIxyUH99GLafRN082iGxVrIXQmDoL
beK0Br+Xuwhd9mBg+BmV1bfCOuMkEQg0B9CmtpLgiR+DMNqXGmHG+vnS3KNszMzo
0WDMaaL2NhHQP5pWXgyXmclsduxQM2JvC5eI9S9baNFv/OSX65nvS5Kuitb09K2P
oj/TEPS0j4cC5qD4tTJXsRAWM1q8OcN49/JhzUuZ7le6vMgXXTHWQLNNVOXJJ15C
eD5gC4BICRuM4Ig4vazRXwETvfa6tiKdcI0dDMP8zTtL+8AbIGaN6mbR3SfLgh78
hV8DEO/FznUm0DwckhKmxEsnR5Nr8Cc/W+4olqaSvRWM/XH8Cd5J5VUYm8Fg4dVa
EvmLkyL17C7mJt/jvVyXR7Y0XYb5BTLrxv8IMz3Z7F0Yuu4DJW1JcIpMXMJVWjCq
2f4dYEG/e/uZ5NxmxB7YgO6wFUh8A6+BSf0/71VzukROd9egMrF/RbA4/rIaJlb/
Eb7geVTJzYJqfF3TsWccff5dg9qNUTEf1ii8BF+T5tx0ABkXQ4aekjVJtPMaYlHF
GWs6k4PODUM3YkantGSOQvsLXZ3nXo1uzhFjNOVGO5gxVTF6AmVMDFOVl6Vgv7aV
13ItIpxI2u4M9v73LXmuBUPxIYPp1yVZ/FTJg4BKh0MOquhAOAJTYGW6z2WteeB6
cgOIPdH0dNwNq3pcnSl0wyi+hPKxcAQJ5ii3WgXhzCZhXHK9sFMUxxqGayfX3eXd
zB8qHqQseXbF6t5bKdyz0Wo5hgreJJBNth83miMrKoG+6Ay/mxQjxzTgdfeg6fF6
En+xx7LfGUUWJ8j63rVbdzpvoswf3j+KYefVVl7Z/LDD2+GhD/VI2kFQEQheYLC5
1hUIhZxhZ2lxbmLZamDcAOOB2mQxOYdxGsSR6TysUe3LWxJjrQ0nl4ZqIfxuDHF5
oYyX5xQpQ2t9IFqYIkQ4XUv/XkNxm30i/MJqCXTQ3vOAeM5bvtArXgMyWTbysvUQ
eM6X39aHGq9EHupLh/ZJdMcaHAQ6lw2mK0Sb7zWLwY6LPnc4u2yO0VZ0rKMZl0Qk
N06d+ZoptFr3/5Cs26r2ztRAu/P2y5+9tnUmDnrAlBrcfG9dJKgeMkBi5td4nYm6
unVJ5879XLgKe3nrga1WeZBObjVPvvcx29DkTacI24oOrD1j8zSx/e58OfxawCRU
KsECAiYUyIF784koQtKILR/1Zf7SDYwyDf/EyZJjDTphUBRXiOUGapXZpKpwAdMB
Euyf9HqHYWTxrpiLB8z4UzrjSd2CULT67OTJwIM6dGhs2botYLeotbL78EX06YJa
KltmLloh3jI0nivJPaaA17oHighfdX6cWhGv67AFT/DqRn3qNhe1WRlRXut4/6JX
+qbeY8QAjBhG7x3DEs5YkfMQh/A5WDd7Q8FbMKNz+m5aTGzNBscfEzfVAG6VYtWt
qRH8fT8alLDJ9B0G+A5hIwOaCSkwX2Pc3C1kM5V3T2+q0W2TyZpotlnhnK4xY60w
uurOkAbai+7I/Cp0z+BDZbYACfUrm02XwL5vESWmFd+079AisQR7VT/024RzD/Zn
9gFfb8+skJwOUx6ftyiEg7t3w30XSwzdQmA8A+RtDW985idZCHgmvk0LktelhJGR
dEK6XbZLXji2rR+F3S6lHDXUBpjtskhyayC62t6hLQatNawF0RdZpRJKilwozyJ/
KvsK7UufKMKGBI4pSy0hzpTbUCvpa6JGuzf8lDtKdMgzOxb7cQJIq5fpBHg+c5fU
OH6wdDLKsv1qBQqeV8ubBXN8rVI4ZuTUuBWBHvI+u6T3az3IHQk4OMwzP/fgLSY7
RivcgocOwPHXlJeHDTpbrEROoD5pxDVwJyAlpFgrApWHpyKMORY3BnF/yXS3jiFb
wmiKYQkutTnr8bziPM47Y/t3dhOzcE7FLAul/Y7G+EmX+a1MJxQ3zD7U14HIG79E
+PG9UCZP8kQ+vNp2juScTxA+fK4UM0hqQEQPyngpb2BTzbamImcgvHHqY/Ho3R0m
KNb+HYvh+p1S4VK1Ytr3AajQbvPaqYtIjxc1ozM9kcliZ/JJKxFys7qTMA3axK3v
l2XvboR09uRyzdJKi6tCxTOie+eJCNaAZvy1GMUe0DCHmJbewhs5u/o/Aa5cVSdR
wo6ZT+EXDJ6xZ4TMkg9dS5YiwUPaPaTCrDmldWULAz4xoFYQg/Q4tGLW2MQj6K+p
fIpoOqq9Ci7GXsuLaoNrWGggMZ+gNMB1F11eXnZB+t0osJlDrqj+S0gh0h4dwrcz
wvc/f28CKd5/h2rO80FXnPDl6qyfmpVayjLZxEsrJfHHKkVpSCbxTEuyLMQSjTJi
lo5PgANVMc3PVTqV3KmBfyxiLx6ZJmA9fW6ctzAqgYboKMJnq3r/HEv7VMP/3co8
mha0gcqQRdBWH98qaZL3jOdJeJAUxzp9unfLpJphj0MouiQmGVX4DSgtvgJoVB+m
S1SRUAL+x5A3e7mV4QPpIwApHhvUxV8wRWk1SUyGehdHVwLSiupbLHXL01teCnyt
p6XFz9s4wRUpbUIlkIHKrpVNaHLt9H8MT+hFx941DshfNRedH/LhRU4UrumY0Rtg
vbY2WbaNS5e/2elN0WXsQMru0v7nJePT3vVSBL2LZjpqCrRjLj3iCHM651MeLHq+
5NeBXBQKqJ5d05pCYWhPgrjtMwTg8voEQLVBqa+8wJYpozROCtNaq+F3VuMPYSpf
5cOi8RMrk9sixK4LNV+DWGZIrYK/JhJzdsawcZYf0r5zzg1GzhTYdgv28AEq+3rj
sLruyv7y2bvMbx3tvRJSdVrqAa7ML4NDiNO/TEisHL7MA5fcxT2srLg5pU2+mPlW
Z4N8KZIPuLj4D1iw/QX0BmjmQ85HioGjgSvJWXX5V2A4HDZRPMVSk6WRiHpKDtNc
fffNHgzBL7LNR3f7Qz3Cq2+P68PnDXMcNaol/PP0nU1DgfWhpV2qfj4Q+m19LoO9
HyK53nLpOC57ajeKHXizSVr1sU98c/EOkSSNKTapD7Sdq5aBG2bN7XklsoeUDfdZ
xQIZbyyzOIcUJup1f7feTUI2+8DKKCktbdzgDG8gINCD8NxOBSWJgBGaGVA2GHkH
N1fdLqtU7JBs9AgrupkYpaJ5JxEE2wliQCaVXpIWR3yYVJcyOLzKfwEn4DCad2A8
tcD4pOiVpbzs1zUg/6Oii+ZiJPFoFjCFIZ/gVvQ+SkknMkRUYsj3HLfw4REVxaOb
DChDqYhN3KpSwn2BLZH6yObVaYF3QUMYO/0VbQw+K1GHnU/bd5fSy/yyvorEoMlR
DrdkwzPBocOjRHgqt/wHR1Oh2l9tfgwTrqzOVn00TGUBG9jeKdNn02TJKOZ+tU8f
XEyycxcC8n2YC1sVnpRsNgMR37OyI5h3lph8vMN349UJ6Bl11J2aAHYobDRoQ16m
czk+FtBN5tPqZGmu7u4Cn7Cxdx09Hx2CBKi9L85MYAeTKmecnBiUO0d6pi8YRx99
s7+w1uX9qvBTaKT5rP2YOHhVmuTi3Vt/zVk5ABSvVJfTxR7VoqSsBBsS+rW02HrA
cLro0S3+SGRb715yiL9sqty7VXpNqXIwxDkcWgSuK8cPqDEVcRM9EV9u7W5YtGmj
7F6CFOZYL5X0XwLWeLkbOE/2bQPnLaKB2zZnIOEZfmthcfZ5Ls9uFr2LiJUEL8ZY
lXQ/t8LI5kHpY9WCwXRRF2vyOdJLkJJcvZpcs82NHKBMKyMyQuDqCHZM6lxApvpa
FZhmW3T6rM8hN6VHLRng69ALZ3uuQ1uGYkm2FVrGGNLOl0vWpe4MzWUMbF4U4CS4
Sj+MIRFHagjHw9q23xUHoT1fxZNdrfi06cnpRCVlADqwOe0Ab4xW9kdnqUUvMlW9
Qk/ClMJ3J7vT+R4GQz4EWXDowHHOZr4AbEYMakqc5/vdOT8YOvgESilEVgxeaLtA
z7d+WXd/KzEaUsWvfA3Tcwm7QfwP/4seADfaawl+cxf4UtCeK9HX9fddmYvb8MqR
61iY1wDVUKMga1umHT9KND38WSL7pE6u2SYT6SniAbpiVDe/oEteQWe8J+NtoFZ/
gZ11bo5w0lsC7ePnhMaw2Ay0P+1vaOmlEvsJEiKYPNO5hcFL2rRvOaia9eS3fYBK
i7TIHStKdsSGWqjxYmLQaQrcXM7wC0qkjz1Mt44ifxvI2bPzlwgfudmu/ZrJTMay
Tuau//XJOgXjoVUb56Rz/6sGKA47tup7H0sBs2f0sXCTE0mUvqhzhzpciIJnkXjs
K1QaoVsczR4wW1H2/84X1YZ1dSmDhN3nZ5tQylex0NefCOeN7aXGPewUC7xhxC70
7AVqJvkJDozOt9EFpam0xAsphhlKlCVdsJSNBnOQ3mGwsxPwJeEgPxperjncKQ0q
NR6g5EFqWYzWTlQNxzY2n5+swvpHjs1dQSY3aK4/NxQ1Bs81peErq8ISUNjDwzk4
N4nhjHYJk1RjIcGpZpGq3ebV2tM//OFyo75ssq615z1NItOzpRa9ir01Tf1fTlsR
lVIc/w9Dhyby0fMGgl5chip5a4x69HbOyY0M3YgSVbWsgMSX/AJMRf8yG57B4T8F
p9OafH0q3s/VkYXB5IECeVH0OBF1i5dcImmFviXasIB4P45dWFMH26eIKr0jV5zz
An8uU99c6aQqeOnnwuHLGfF5aEFizjYjzDg4ysF/qDQTfZN3LFkXFIY1w6/x0vJN
InOtpgDHjls+R+JH2tIA8MK8V09SWUcgvbsWuUXdNu7evFuQkIYF3DM09Qdw7I4/
mbkxfi52/7eRsmJOH5VZIo1sajVvo6SIQa6mbTn1dyx9pC2D6wUgIe0xeA+EtpXy
d7wsGOSe0HW2djlfd8wbl+S1yJD4DBW1jHRm9OOamDaeXbzg7HLVd/TcEDQlAwUX
0J3w87dL7IQrXyy5C4m/7vnG608yYnT6qoRyL72Jgf/gVrdNaVp/Vl5KgB2xMZ9v
KHmYuy2EnUyaA2cvVK95Hw7K9HrLNvZiUID6Yg7vNfIBHn6NTcytS4QVNtWVzTwY
1ZYsXVq8pHqcLssiTdNgi2TxxGNt9QUdmpWLIZPwIUb8hIDsglcLme+5cyLFNMW3
bAbZnS+pml9/qUsD20A+PSvL3s6B0FKAuh1L/f8b0XP/Y+gwzAUuvh00dLmECB5T
MkqEB8wtGyaQxAzTuGaMCpgcqfVhEzDsUCjMmZT2ypzNJCWM64sHydVPr1JAuBCa
KkIBwvedzjtEGjlbtmCLAl/j01A5KCdtsOzSLeeEHZpq8xIxXzzsD/DzUCh3GLEP
XY6OtHu+HASWoDclp5GJKo9HLWiCVFN1ZQpnJr+CeUxomXNT6KoYIpsjyiSl/LKN
M54M4EyTHodpROhHnS2B+0RLhzcqBaqq6s6gVzpl4Nib5FI7W31GsgvbgQ21mqJc
LIXd1cPe4xs1b4Di6oVlWpSpHmIJZ7ezr4sbTAeigWCYIEtGnKT8NQ7tOWomR4Q/
NdMdzYprPa1jDefEPBQWhqjyzYbaK8Nh/37L+tjP2mBLJF8mjosiCZLV045OJPXq
RtFI20JqMB0xK19NNGnlkdVU+Zq7aJH5XCDGjt4670HMdeqIoYiqKnX2uZ7D2IRo
vDnnS9Vf8qmA4ki9nhcvd+nuVkSewg4Fagx/6R2WcqJCrQzLLmedorNzHji1GhFh
jjYs/QN8wyIgZ7jJTYqfL1mUAVSbsWzHPg3CHr+ujdn2AByk9xfjQsVtAJJvL3q5
1jfy0Ltkn73QdXttd2WL8GML0ooNm5CTvRKEs2PGLC+6f423lqaNg7WYggly6Yjq
V8cLSgUrfABbAtF5uHY8jiA0w4SbK4Q7XeM0XMvl03EB7QZ5Dg91GYVl9nJeTb/o
wSMbH0/eIqFFfif5j93saIg3WUrQ6B3gKOZ6PNJBDFJ9V+sow5ktPJgVW7jb+7z0
RDGQUf42nmgR9TyG3fzQ6p8BRtPvQa9PvhOkJAJNruKks1qlCTdiw3J3wfW0y0wi
Ax8NwrBvAmYEgLlELywpmKIqH2SQNt15PIjs7zOoWZOjz9/PQgOaI9l67pjITtLd
GIwWqmuqorDAoDpji55A2/9q+BhkJMNus0A2MHkxD0fmRQy+GVrA2ygxUxVEdLAg
G6GDQPRNWEIxwe89H9SQmqMroGPxyi5ggBXBFwvPVHb3S/toDFpsGqvfyxEPHIzS
WtEfeCryiNSXDSEccHy5mAmTfdLCKLkd6rsaHAMgdSG5iIYOGavYwB2FYxshlZeD
qQRo7Y+G9/tz5/01mONDdPSYJImjDl5pnTWF3+HThReE0edFAcSh5BJrjJ3wZaL8
3zgJJzwDpq48DcPCkzOo0mEMTfjJvaYF1/bWFFq8H4+9e+ZdhloM+NBkNwwYzZ7s
nFoPPfICyIqRkv3Q7ecj64ZvffGaPsXQ8G18rZC6RkL7rSaA8OhgCfL7IJXukzjh
/byM9/IRb4JAefi/1det21pcvdlf7DGfPnqTW9pMpXY/TQwAonxnfotYrDJQN1a7
JvCArwYEbn1jY6jeZB9fcV4I48nFBJY/yXxI4uHyB7NonhKIRerUW4cSqVU7QgJU
MW8lImvQvZf1QD69EozNxysuYOZ4mK/kWkCHwMq0/g5BYWdRN3IfWuJwYEoUbpwR
J4wtsdMeC+p1tBDkhl3fks4DkmOB0F9gkRLDL58Kb8B0+3oVqKw0Wg7JETi6npX+
P4ZHIkoUVot6x+Benhlv3W6V8lSiLXS40TECq8OjVDlJFWq6l7zQfjRMwBS5oS8M
IvDT2iUZkhU3wDofLsetHt/FsxcVWJuZ9IN29Ye5dvCrcc+DiX06KW34bHTxtpP3
h7K3jJocphxZdWz+W2s1TWPsoRNVIfIHvxwfmmmb31z+ggcuL5fzxOlxVlwPNC3g
ra5DbdsLegMk6P/zBKPoL2buTZC9RVBQzoG1xI0HNNwj8yafDzLxplqYFxDL/4h1
4Wle4PLTMWObb8FehB7jHkSnCQDSJaTMNaO1c0kLUvcP2O+w1F70zQfQ4khZPMHs
byBI7ItMcvaehs9QAMroMZgX0KSi8RbuWsZWeWtdxlkTqDAD0CnbSf70cFmwh6Lv
w1cGdEurCwFI5cPpUY9XpXHuFl4V2W/6o077SruBPTS4/gnFY+O1IDOGQEmHPMfD
2ylkRtAaJtU/vhqeg9Bdb3OUVNcd7/QdR+zO+nR2XM8oHJ/CYxSIKj6yLN3ozZvn
9O0T83EDbfhT0ZQygdMmvnj1dmAtoip1cMP8axw7VDVb2ikar89vhAojz2JHr9AT
Ogt5ud1jjPX3w5RVQPYzkJZXuGOBUzKR0tbg/k6+lUPNgSKJ+xZom3Upm9+r4ms0
U8XqkuWMsPkHm35wnBgvnqjtBqPrSn/MM1IBxl6cfL04KgUWOOUlYKgzsO8dPu9Z
v3Yw5573mxGvtzBdMCQvET5LmFgLZMrQk31HGIc/To1EOF3dGpSP/lQKe/bjjnJN
240ZVM8XVsIZwHHD64Q1S6dADqecf/L9yHUgi0tVZi4CRiN/V4U9i0B73XxNBarJ
M0lLgApSRfyuxFKE90NXs5G1UIJd3BMhC6t4WZq/rlBRGMsbUQYUg+JZd9OIx6q3
UoZEm/YuWbb0wsGe70jvkvv7yjKHde47oZ4wA6T5L3sILa34Y0Urm9maHKCBjbmp
c7THM3mD+5MLhUdBaJE3ZOIHuQP0xWTyAfy/TgIOtKCTDvy758IV8EyHl99jUn54
9xNtEAohqQNFTTRMHt6EMVm6usx1iT7hpQcA98hiUcqZwUpjx0ALBQ8yYcTy1n8q
vBc96vsQRpNuhwioTmFXK+/xUiv+ZHguVZHoqOLAtpe2wSfxUMtRyGsdXvVIn9FW
XaHD1EhvxeHO0/vxLg7CpJbEloA/K8N9uy/8+x+LceuLI6FMM/z9D+1rdm+aq4qc
6GogMWKfcN5A7n0dAqZDxMRaQSlXhCu59CxOOUtziYTDjpWfuH5MRfF/T098/WR8
Umcs+Jm3Wk+dfXkZbaFAdoLyIUKoeFGNuloI2BzzRNqEY+qPtEwZLUXbsIppBtgi
CxGcYj8sictuYkhrwhmaaebXGAnrrwgIoPxcz5aBkIVkYarorEHSKcZBHxPSi9V+
4ELVbWuo23O6HxiZF85zyUddfQWX9T9BcbLUWWJ+2xOu1fQ+qGzd925iBIsMQM4i
TQFzduHAeyoxe68hJCWHSX3S4GYubvTLMyHr1YgiWsBAE2Zw3DmUnG6sHNb9e0CW
got5mc5Xl/k7DkX9OXRUzsfmHUG9H9D4o/DVpGSSz8WQZjQxg9TPFBUBTvmFOg+q
D3ft/lf0ng0t0BRs4fSP/iSxOz9qN39jJBszNjzm8knNYXwpu7sHWVess6IWEHy0
HHSoEq9rD+oikQfrNOjqba5C8vkN1qnhy9T5QBDT4ufrFxsmuOOV0neAfGYAEYGu
ALZtcUP08gAwZ8i+SgXTUWN3XoiQhiLGzmbSH/FS3cut/Ce17P9qYdsxbPRF8xX0
95DfQI/04u9UyF94zxnnrNqPM4uevXaYKEO+ksrPfcalAFACsRi1llrah6bJghRw
cAUpCwr/gteR8DCkf3vTv6Zh5XRlt5Y4rxsoidRdGucKZitZX6H8BqK5kv8j/RYH
jwaQgeDwG9u1zZ3FkhoV/NF5RohLHB3XUxZhsQlWddOdJhESqtXUgwLnFMLbwBTj
AeWD01EZFIfURRAnEDEnsTtBE8l5iHDP4uNUjSlT/suelFF9V8fFmfEAb0pd+9iI
R0LuIfp0MvS5Ngx678lhR/BvZoni/TG3cduLIi3/J/aVgTQzk7l6idGc5NVL53DP
FLagw6jVXSgFhoE/pL/sakb0tp4nEqD/vTjSbTuYaLilwTHfRw2qBjpUVPz8fXg8
p3PvNczQZbAWM7pB/ghiMLh5iNPLiJ12337gFpm0DeKwNY6PRi9iTK17yMMrQLEf
/KAF/hsrMrmBtcLyzBvVBFLJarcTAa8u4BZZJVKuFrAlXpDgM/Zyvwywp/pS+lua
3snkBxx9unvO/Cek01SwV8aZ4UU4gu3GXxOb3M1x5dj4krIX4aJuqJ5w5UvFrhWN
MoZ9j6y6nyk3ZWVcRHYF3Jkq6aCM7CWkYiXmJDaceTgafZugU3Izrb8vffgL6f9m
bGHMuUUrQ3B/hq6GkxjFg6lQbb2BKzZlnQqKu96MRW54pDw7A63zewqC1USouakr
VkDBf0aOm/mTpLIGQYVhVgdh6TeLRw5MeQ+BnEUh4fUE/Nwmb6cisiGVnNOtq3Ur
xe2X1Is989UOYWEhvqIMEkL7WyQskbAv7SATjFQZD4H9TGuZ6Jw2bqaUuIARDLMe
MrBvZr5r1WjXhg0+KPFCudAAtXfaFQq6m87qfxeZz0RGcQRbuai0Au82sjPp7O/U
nMq2KtD17hBuf9QKhpRAxJ6JZ6n1Pv4WeB+p4KZJ0tgzvPC2BomZJaST1cI/IO7E
s5TczI1rWJdVx30ynD1giIoBXdKxR49JhogesBpJ5xM06yFiatmEx7TRF6RkHZTX
3myHkG63o8Z0gBXuqklQhlJyApPQhQZaWArCm9DmOFEpTqIjCDKdaCwt63NUbmBo
S0Ev3qdEo91vVaca7ZMe2nIDyHUoy1XzBXn0UdXBHXf/8XRBp7wm4RaLjh4vyLPq
I0GzF0cicGbw/XRU9yI5FgiJBD4+DWYhuwlqdwuIdfOHrJQGsRcB8t8VPH0J8C6d
8/ODzFmLJd/ar53PxOpI2Z9PEWDvJfSDLw5XaaTqq0xFFRd3s15FV1aNBsQ5sU+C
cFIWH7Mlb6iG1zds89ESTMF0iWhVMvYBR3YnjcBHHLYH83UJ02klZOFeEwwRkU5P
crIFbJieqMmlCVaSNFx+4bLsI3CQwGxySRlSNQZoascsF407KWwq/FUUv6oFJCYi
4tFmQBGoqrFqyA4XxtjDBecfimYVu9RVfQ/5uX2jRfWGfrUwgQa3A5sLxLwA00m0
uvHPVpVAzW/OH4n6dWvdgo44i88P+NK2T2jB0qwMoarvH042zDsy5PPOUpKHC2j7
hsWkC5wkYPPJu8JKGqTJdoAgzBNGfSqgpq/OneLpXF491tIuBQ+bTrGEIfdBvyDu
LIjqTU0SWYkFOZuhRBfhn/u15If+dCQ5kTLtvW9K2OZEPknhy7Qn89OhwTawS9eP
fUU2+QQuMHiSxv8ZW95JhTKVl/0SPTvPY+JsSvAf09M6eyX5aEDvbZnFuQowzc3W
H0GdnBkRTk/hnSjCYnKd8LAkmADwZsKCA9iMhv2R7k0qjjoQIpa10Z6pADJG+dw3
JBGULjdBqpgYWeL4k551Lw82Gf66pBNxgsgjnfUwr4aTvvM51mvr/f3++0IQRc+2
ATeF3+XMUn1lP2Kq/9F2oGmjs/7O9TNhjd6LOQTHAfqfydBpxAhELYnaBEVMUtF0
kqkgkZHhLuFwSFf0Yyq/ynS2V14DiiaTZ05wNiaE5H/egzVoSpMgs8eSTfRKzPfh
sW4SBbdMeGfQNhV36KNvHha9Nko/xOdb8eCXOXD7JAotickYbvcp/pSZrN2DS5pw
bNyY36YJodyx1BgbwHLGrw6t2DxdEVe6l64ObZrIg8d402DsQpyL2IKrViHse8HT
lGUdpJu1slQs11ZrNV1sfQ1YO1yvuE37kHjggmIqW5gdqXwfgbuNwMiYflg7/hVB
yKnWJg96R33CxKed1IVjilx5Xxdbzy92r+3usxyYSQQt15WgA2u+1GmuTe4iVVqk
jgQ3e1LCUaVK4BWCE7Y7G/FjfmvlkBO8zXMF/50LRZWYLNsymVpPA2OaDZxFbUQF
tPJezy+2wQX5kAfwGz3gqEVe581PMI1TadW/+28frx+q2J/0lBqK3C1Hji0LYZ3o
nAkRuXb60vgigUXVMiArk1Ki+qEwC7CB9DbDa95mm5jP0GpCueqni4K9xuFb++oP
sqBvw5/Okwax2KMAMJjjWFNcVqp25elNeQtRvifmN33ncaUK2aMLt69gdiIa5v2D
Iea3kfq3Ty0Xb+iyReUXtEB3LG3YB8sewlJmHW9TKrGVAFMc5kbp//5jInPoHpY5
d9KiDd+RoWcX6/6kTJAGyI9YTMcljmn32OoJwCBTOg3FaZW2lw9rJ87b2huIjgsF
3NGNGC3Qk5oOpZ3NJf77X+wQtQfxNfkWolCPw4mcI5Z17cESvkD+KILP7z4n/ZSp
Uxj47Q8K/qR6wDyXbQ8F+rDbia0PVV/xTmbhF/Fwxuea/QYBGKuL1XdP9i47iIqG
qhcoWUFXxGa+t1ATaw77urwU+mOU0mdhDDy59wC+nOXY0+r5PNXvaVCPmBDKLqpO
amoLmJUpZokHxhtqa+ltZnNDkCu2ta37G8XYFtT37i10R+w93xp725efJQPm6p40
Gx7kg6EXrxdY45myc3i6Vr+L6P4zSopU9OtD9Sm0Uz9Y5j3upE8GWm+alPIkJb3z
tDktFG2TYzh10guyhbBBpgtteqvA2aQLp1A7DGoyUD5tH5v3PTs0OTs6m5VifJpx
oDV46IoBy5iNCmIaKb9bu1do/DTtAEgeyta+ASaVf5RIeWyQRarAxv1YC13EkxN6
QTPIdh0FC43lhHxhnpwyIErbe2aBPFW34IfDoECPxFDF6DAMTYvF27XV6Ps56a12
Bxhke2eGMvgIZpvLMmV0/ClkAJdcJHS7VzK45br3tIS0ITR7b1LIYn2ZnVuP9nkt
9gkfD09dOtSDkd8M7mJ0GdURwkw/6XCQLPzF5dFyGjjaxlk4xQolfWdoVzZB02xF
s8n0dtggVhkbOc/TiqJxBASQVCBi7WC+r86zDyHcIgR/ZVaJuDPb4WtvAWh7GVQT
CdFD20F9RClAVUZw11nbEhF27PNw1XcjJqMva19s/OPDuFpydlUQ293WT+nv3kPP
7/XzF7vzNWTlZonFa1X3zmP6EQdEiKoGESngrC5QvDwdnx6EoX1HNtntqBkYJBHj
HHtn1RHyjBwg0guC+IPCI69vCQe5gozmBn+VVOWOxqmGGTfQyyQf3+mIqOf883zT
PoET9YOmXDeeI5VgP93/OaZQi7ddLEbct9qqGKjc67yNKmDUHwSlPdiY0HjYZvkY
BXf2pKBuwiy1JSO7w+sb/aH0Frzho4lbgL6gcELWc5Z4weNfYxQ2256KsNqI5GwX
PpVXwyJnbSZwKLwfeMBJL3SxHe+nDN1gD11+NrajX0Mk6QnaHNS/lo/VpADRqGO+
xxZMphL/HYUzG1K/wGezZyABf5Rkn98jTYYWLji35WcxURhj3uOFS59Q3ndCSppD
khAd5boUN1oEqGLi31NEcMhxDFrrdeyV1FZLhFxNdVM3sPCaUmBZpE3qKmPG09NG
ySqDpBwLtoGw3KlSXCPwpD5kbSkK64juDkKhJBNqIdnBl09JZstYPxnRgjvnGaO3
rMENCYlKoItIa/gTRMvdLC8Pvh0IOMia9el1mnlKao7OAlbjfu9L9+6QuIYBnNyE
2YKmf+ppSebTlOys6Oa30l7hX52a+x0uHQrRftdh8HlSGswxjZoDPFc6se0jkMDM
PGEB92w6o6MB+CPckIcsQCOjj6yxQ1z/IvZAhwNFKikAhsmDX5TwzApKG7Xt0tdP
3nMH7wWEJASJNMDxfWUxZfyi3vWmefkSFdWKVuf4ZrWdLt+9AKb4Qd5kO+oH53W3
fTW3TK0hpIUFXemRExcK3M3yAQ2wQz6TCnBY5Zu0DoRnmDz+hrwQRiXSqsIAYbAa
HhGBNSZLMxGFilcYtJ474SiIpL2F4aDYwHCsku6RXkZBG7PROLHi29H8ufQ6NCly
yKBJlF22wk0+JtQc4BAcphPgXAhkd90fbrqI2Xy7bkUJJhMSkqXrOY41eSjz4GVG
if4NOt+mwQcslPAbDy6YQj6U57cFd6SZEB6zaz0Kr6RIYP9bgKq1X0C2k7nzjtr6
kgYZPeVl20JSOeP/LvHr6DWZXpAFI6ZK0m/dpv+25MB/NgCPt3iyTCN+3a46FwvJ
PQG2H2DS+3pmsW2CeoEF3k6QNRaU8h59/gx/YOZU2d0w2WxEQg8deOEW1xbTkGdu
wZ7M+xkTCd944DgOt0U4epcnwXmg1cnsv2KXOfFflhz6EwKj0rXM+6jvgckNpadC
nHG49YbdsWUTxM4NowoCnLe2pGPhnOtgMqiVIwuErrJl1ZB5i2RCAGDq4ZvL8T2f
EaFp38gVCIW5ebyNXSSJFqTFV1KRckJRInYrq/9TJsWmEKxFCwD1A8R6ApSRxw8g
og7+ZL2gzo/YPQMtw8fgAiBIyopAo6XV/WJd3vNmkOFUADLUrZiWI6/1Uo/FTvpi
Qeiiu3Yinh74mnu1pVHsnmrfrXDS9IM0e5Gr06gNqoZgOwyEpwrTjdqO+mBDW0Ke
87WCNZTzVYubF3kHaI4buINsKYDFKOhjFXkTKojNmJXKGdm72PLaiK1q7OQq7zes
jnIfymukQsxTlByiny4u7OWjhwqGOhD1lqblMduD1cGKAUXbkBU6xs4lg0UwMklz
e0/cRK1VqhKJdIW1XeJEqQTR+mVjazVvYwwSyhR7yVCmZFWqEtLp1rNKHsMSOn1Z
fDMvpPkegcK5+DckwdDIBNRs9tL3/qGFwaOoQdSbJzrb4T/BHi4rOjpmw6VzZ57n
0ZaaSuYtOn/UgTgI2YU7L9o9nG/BDVQrVsQ2hh1S1lQdT7YqUptz6Lvyq3XUWpCn
RHMAl0ndXw3/w7mMj/xPYIHGLn1TBPuC0rwn91t4d8zKE21Wp790x9JgX+90HB7o
5B0lVE/ffXJUmlXSrv7s5scPO2VgKL39nsTSrGR5ixqWZQZut2MwwivF2UbiH+bA
GAqxMNaRY2Rf68uzIocsjtKVVdEvX+uqrCkx+6iimUiL6a7LXvkKsKNnr21YUgUj
+aGHxhVvwb/JRidaB9HZA0AAWgTSoC3spUnupuFuFhdry+ugYOF1lzHllTWoklJn
GSy35lNruhWCmZ92FI7O/u3NRtWQwNp0GUgUvCoFH6lA4BSWtgOgTjlqkwsm9YaC
WUaAGPZdZy96aggtsjbA28MzbUSfyx4Y49y4caKQb37uFLGFWebF2n9MGZzXHZg2
UjZzrDFRSxjHSBdYixylmTbysV+pfUJL6xlTiWpUFTTX3A4yE6Z3rRvorwt647Qk
N5KU7T2j0aln9f4gIYRdR11wakLj6lw0GCrobX5QJ4l7shvtWMCQFQs5MSzPc6QR
OSA8QQjOqCy3h8iqxEJaczsC1tL1qKY6nKZ/8iqxka1vAepaIgarHO9sZ77Su010
tQTxxmuZIAUBwNOke1JST6zbrWV7r81vkdvtJxgpfy/cUVWU0kELLsNNN6LuJtO5
3ZPqoq05XvDxIku3gqZCa4dvBH+AiGiFaLiNUKbda17t0dxLE30n75IpJqMf5Ug+
v+N2sCV5xQubuwdYCdyIjrzH/QCUi9qqpla7G3vgCvita8FaLM+7L6QiV9d9jn8L
LBpIuyVzb9saIWl48NS0a/HJO6HalmRDc5tbA214VQlVHcq6ML9OEPCFNsjr7wMt
ccAfJzZwHazVxeX6eQ/bqAVhb7IQ+fLIRQQ5vdsjwqRTqk7QVLyMyeT9Un66QJkb
R8GVHrv5qlwkxlU23RzqgwpMLTqN5tDor9iN9BWyd0jU0Ip8HrzR8VM0glVi2Etz
G6BFb2wm8ctkVpIQYlhpVhnEDbUpXa7DkYV1UfH+Sskwco4MNBWmH6oWL5slXeo3
Q0Gg3cS8Zp1lxfjOPHrcCe3GtiqLYSmjIj/jvnX1ueuwJ41HBGgVBOSTYP/T27VH
nAVPXL3RjPdf68lkF349cAZxpjmMcJtroDYzmfgM2Kk36UQt22y0bmXlYvYZXfGX
/vmZCdRDFc5syKUZzqiOOGtOS6uR5zuRlFAFwDAiXGnegBYQ8meR+6LGfRZsZRKX
MowweKksZDweISWE9akRmEOXzmqSYqneJnWeV0ms2N+MkcLK4m+UESK7x+vA3eWa
4mH0v3n6EyDM+XA6PJC1eoUXT5FIc48j0iWrFxUsEj6bZu35Ot18TzIkoFvHfWez
nBn//bCqUwBXqnsJGYukQf7Axqc+8KWaYt8Kk2uH2AqcuzR3bdy1i3old1LMGBSY
UyG5QA6dmUuwB67wfbHVNcWaZMa87MwB+XSF/fUJ6px/qGZXf3AhOXhT4jGeBnVl
rn8woRx33+6r8BVGmCw15UQRpr+11rrbqEfEOQaUI/4QCsklKMTrn5jG4dKAznBU
zQ9oY1E3e6EJnAoouPYSiAVcQDqZ9sgnIzpu2+yfdEMbFLWSYaHulLxqelhxbXdp
JuY/aWthLUaf8XE8T1ERrmzWs5pgTbXUsvSmN+343BkYLUMgb6khf9SqiTTwxiFs
UvXsIhHaITIj6NxeBbHZ4ucoxBkfPiB8VaQ+nRueA0rxOpe2BPWVF35/Ns6OBPXT
TmgV7WmR4oAA0IU9I63oii8A/sDLJE0i3L28Z1P+2O88qUTniQ3Cuwy74d5UKZUW
665kU81lVg4G76Ncgmqb8GX9B1ywThfVnAXy6iCJhATkR3pVBHeiK7K0hjzjGDeQ
oQ77hLLuWfPGI9KhKWOXPEfv6O/KxP961mwf4jjiOlQ+SfIoJ0WbiEKrdUSJfo59
BXG3/doXHE4qiY2yqh8W8q19ITVsjRTftj+rwdRFNEoJnHgckGuL5UCSTtMAegVv
N/rfzZV7Dj/WvdrIn4M7Ztu8gXpBerAZV91XcCyV0fjhkwhgt2ALORbXWGyFE7VW
MLpNPGAtDb/hy7+dLjaJWb/S9UDPHKg+F118gMzHgn6st7HuJHSeIfE/NxYGpufA
3uHsJN6IKCVsObE+SFaBRety05xjn+CXlqUBuhplWjj48c4Y+k21lYgUVx12Xt1h
zeWVvcIgnyy1P5Ot0jjBItYx0kkO4n74lknXmpNZOnwDqrhxUykVdfgIv7IrwFmS
4+/otDjAhKjOw1rgMJKlECFpLcVadndmO3Mjv0WbbkuYdHiPVzd/bZKTd9oqIjOB
x/9TR0ZFvZE/87D9emef5bCc7ZvrsZJxma0oYJGvj7vhx0yfZEuU71Hv+WI8j7Mf
e6fcWD7gThOT6okKm46GPoLZReCo2rcqKLHAdWC5/g8dkhXB8US/gi0PsvQxYEs9
0Oa8GcP35yCPOL57GwmLjXYfyn/tvd120ZwyLJd9xV2gN15Gkr15VsXygsBV/iCC
f3IuXPTuAdcCnfjOerlRY7MkknkY6TDRQDtioVVRYxo3VTjTTc4cr930heGb6Me7
LhmhZWV11EskOO+JZcHOLZ80M+aaEZGa04ti6nWREVodVA8ai2pMbvqzUgzsrLDj
PmG8uUx7IjOaChVY2uQKWHHq/vO5ijH6I8qV4kbyg6z1pZCSDRd6fHt2S/aNgJEU
8pvpmqxSwHXO0olKBJgBMOyY3ClUE0Q57/kUaMcmidxX8MA8Zil2Gt1iDZiRYGld
6XJR3zTeYmkHdLlTfvgsUwQvgdTsIQDw89+dlx4ZQ0m/vhPogiqo1cz4yvW055u6
bEXEdl4E8ZcFd5nY3TuXjWPlTFLejWMkMKg3Z7xis4Ueef5DPrAS55D970DsG3xT
GVTN3/IS79upE+IsMckwGOb5PNs3fRPWcfzYfXb74TXe1IkESc2Pm5EyMZ+VZFuz
ql4iiOk+Rgsx06z4h4ArINnApEg/3eHLy2rGz9m1o8ADUy7+SdtIvAKwZx7vUhI9
ps+Tm/RuIVjEMI3N6lpAjgoVEFbgODWKv1sFwOcxH7O0PbTGC0lZMfqMl10yH6PP
r3Xk+xpWjK/wp3/1RO9Sg0AM+pmIWmjzR7lOavzDadmuR6EGHVLq2yceBPPiWO0x
MQZLN7pfGbeRe5xNnjQW6mYW6bF+oGd9tBAvg7etQkcimwk4/YWkNlkgXatV7wt0
IyPibuTlAPmCDEhtpJwkq35GKbb5Xst/0Z0jg6Y4DlLfNTwe2jIMLAlsBiyz2Wee
hRaE+Fnr+Ux1fDym5QetHVuzOXm6NNEN71UO92ioINN/+ss9gTLWcqh275BgVEpE
TAfebdENA33VSMztskPCexKX+mWk9gtNVfXO749r/OgiVSTUUcv2nnXqeLgAf99L
yQH35XCI6IWnEbYz633to7X80vg3tGhDbr1ABVv24dkKrXa9ipL8m1ehDCIjAF9l
tO4IyjWyBp/KyzmMF3E0GPCi7rNX+RCbKnifeOhuA2LzudD3dZaVhNmahCapDIsV
ZmidGnAMPkAjHtV4shuevt04ggSf9t4LetlYu7aW0bskaQjoXZw+iYMf/cgRbw1E
o7ejHd2rZFpTgXuzd05sJ+BtaLFnpS8dlf1zBfc8i7L3piWMGoML7Dcg5JrofI6C
43KbcN5WsNjFUxCECTQMVM1y8YjhOF9OwRUW40WAiPxDp+1yuDkpjqEixjxq6kms
agLBB1ZJWCrlmh2jjA5/LhKtyFAqyQl+8dABdxHx1SERU9wSX15jH7FH2IvOaFXX
rPraiIQWXBUTxNuVObj0zuQEaQe9/fwV319xFfG0qDaQc390HbWvhCWsQ+hGkfhU
xeaK/U0jMP7oGp3u7ED8RiOJKGHg2jeS2eyjvNe7UtQuDS0xeLzYfbZTAmORl2e5
4HBk12KduOQoIgQv+I56LSR73dxp6FRhi/DiT8uZCp0qG0iBnw54M8Nav+c8xpzn
5dXt8uz/MPBH/l9o2E50ydhkGAJVu3WnRBIQqY+aKZhP8oZxE84jGYk7NRW8FtME
taxgCQCqxF/O9WlBEFOQwiIY4B5lPudUmp0LB9S13/bduwBSTupJp6aPq1U5tTQm
cyovmr8mGMA7ra0MCtay9UO/oQCu0HNyKdXG3i1TnNIR5fZgvyB0AN8POR+vfcBF
lw1X3TXXlDneVaQlogNHmDIbgaa8A0sgqoU2pfqZl4Mx/Z98XJ9gn1ztwMnOyz4a
7+tWmLdsLXTM1g591rAzYfP/W1DaoihdO1QbpPq9mVWnMv7bgnquyJ4f+IgweDVO
ag8Sz7pbFcvIh8SjZYD3BwJ6tJfdyQy4YEvq6u+NKspiwBhg7qBczMahk2CiXXA+
KqcJc9nnLj1rB6YF4AySARB64wN0Gw8PRTZ98Rkh3wI5/wKKbuPgwmGgOQNO6Uja
oXbYojMq2drFj2/qV3xgq8aUzdgfHYVRkJqatjEBuBW7E2oSAqgQ10EYKtpX+nHB
XyMDkd36X/q//hVjb8204t458Z19vuqwRxjaN0QOMD+y3/6Y5mRJ5K1jec+TtRGq
E443leesKptihVhWKQHjzizyFETA2HbW1jNxL4T4yifkjR0EGVIdNQjZZOvLuQ4c
hpgu3GUy07F1EojJ969ZrcspptfmBZLyAu1KBzmeughv521OaUcPutdMcYRGGGPL
MPPIeW7ZP07+HDwHuerYQ0RKWnm1OYJjbbRSSFMMRTBPnggHmOUWu6B7kIiUDw+x
U0AuB/dm1Frq55eqBfCXHxhafFu1HZ+jd0xowl7dc7/2EHiedMkhlgzStrkGKdge
VZpQjtEXlKA19d1tSGmlmIZjqa5jrRJ3YQN5VoBILrVQu5ihuC3XASrfbOVvYlHP
W3qSeFgrsBwxCzbalTS2UvIA+fDPKm0Q242KoPeyG0SYcR8FitRPG4NyxaG4m5gk
T4mdYGGG6EBPlGwL41uqPzRCvpO6A7rTdSw5esgmOp59ATpJ7rwJVEmnwrDc9LXJ
XGWaLcUWjzuC0vpvygAkSPgMQAsHlrwK3uCyfqmu3x24RhUUB8Rhq0KLbbnsAek6
8RJ1oxEd8U0mOSBKmrCekvG4xp/9D+JYzS1YYuI23oJnOgu7r4hLeIr2hxEDQTeS
Q3n/Y0sk91leBLn5bQOzhY2pE4NVCv517rXmmwrU+TkNNdAvyV80QuPxxk+6EL6I
ykrnOlg8sN9dKVk4CWHZOdG7ku4iuDdtV1yoQp8KiU8sPFtcz9r2ujrpacd6ijJg
idAweBhydWR5btPE+rZ0SIss2H2T6P0yIKZWapjjDMDYowtIMQOZ7t6rXV593HhD
qVQzS94bmoW/VQ6uq15miKFUVPINhHEd9zJ9tdZKZgPxDwetCs9CmxSBpotiJjAQ
4nKmzvcfMwA75GdPO214ehgfr1uU2ZQX7slu/2l7nuIlKFShtX/YsTmMJMs3S0kH
4L0y3UjEgJowmEJDe+9vp9aKD5I7rKBvYAH7VylUrTfjLLx4K1mdz4xlrnqzQF3j
wfWSHaJ6iuuqYPgYsneCuilSPmq5zQkvkndIMUICqQa+0Na5wZSdxikwhGCSSsG5
6rwZXMVbgURX4MkzWoZ9YF9bQY2c+0TxNSUaAxSANrr9OGKprjG9EfcRr37QE1iu
O4UPFzAuUWv6F/MObTyV3XUC7Tq+Ov/+2Zhhs1TNKGEpCEi17u1tvZaB6vW1WaxE
G+AiWXV29R7iEa60jOJUP7ndp69d3AlbdjexfCtVKbCmuyI8upXJxE0LRDgZ8D+C
HHy7srObrdttpyMsE1LA4tURc9JYV+833G45hf8tlvbGptvgo/mEQZLP7xvR74u6
W9Nz66fJqKujs4jdWXoiIQ+bAKjmOCsKfD1z6ORyIam22NxXbW3aWmDyXvunGZ/j
U6VXxBuTcZk1MhNc3idgG395EJR0iY4o7yoYz9qKdZZWwZ+hXdllgQMWkT0Rrggr
tdMgyUbFlMunH0Zxo6oEKX+xjM2y4XfiegqI/gDhsjNpCeuUEk7lNd2oCJ2dSkHm
5McOwdGgyLypvBvtKacCgScpLwgXeSSOwHhxUFAK/JCfbuM601v+Ot4ifOJzMiEI
/gMDBIREyj2w29ytAHYUqWQzC+8XIJP34pa4zEdgUeT/YhwzHiXSUa+eWMrTc7Nl
38V/GxVesqlGipSbLczn1mf7oD78z99LqDO1HvNVqizMwtDofZpN/kei24tKCTA+
CjoqEMYfK8iQVAkK6UDyKXBt+nz+MDYB/gEDTkcRGLjMdeHSS6Rk0+hTTVksId+i
uKGGbnIoI/a4Bgv6U0etypBWVCUozsLm2l6XijZVpeuKG3ToxNYYGQc65f+U+dEt
cAMx0VXZHve/xiaCF750lujm2HR1vLCRwb9s/BHIhwKQCJKcz4hZzTnHgKkwICj1
mMFQwzL79DC+uX7WLUoyedy1U2EBjyi6gS3y/8nhGKiJ+1B6/ZTY3ywV97EvIgh3
EfJs4sIz228QVKNAxQqTmIhfOFrlAeQgPK+JaKv9C1ad0f2zynwd0kU+yJyDOWGh
Qo2geZGjHScYFm//4kekErdvn5nMtyjSvNvXSK6l/X3dZSj+xGoQWHYMgk2BFX0r
320lRo1QRbSkzSgrszxYTZmqeXRuHRwnFTzzA05/cL+FF+nSzcRZlapTHrP+jaRh
KzfVxOtQMcSyNMYnlabY7pO6hb6Yh22ZiIJeSyMRH1M6uEydKK00LPpbnIq+9TXo
6qzey++X6rB0aoKSWAWvOq08q8UevA1B3UBVhe8L8aiM1bBqrGNZ5KYwrXBiiCfm
Jdiv8U7761imkGuqaw6/il2FrbK1Zpba/k+83P7GdOakTTrjz0VWY+0S/wWQnHPb
tzr7UEE9IScPAzJzV3IEZIPMR2+5j7a0xan45tc6KKqR7pywNy0NIss6MHuRT5yw
We5i66htCT9GqeG6EpLsRiIAFpKlCXc5MRtIbTqCiJ5Vz02yJtVTRbKx40DuZJyK
XabFKrIt0yAW/6e1xJ5x3kY2mJIlzFB05DUG9k/7UDSGL9EYv/kZyL7MOiksq4oM
CFL75HZ2hZuWBwk8AykfyJMPXRp4wmoahm+C+yX1X3KZKNUJLn3EOQBkZBh80ozd
4qWLwJ93eZg139Do37mWS5ZLR8w7EGsHUIZof+7ftO/ng8L+bFEhQ492JNqgcXFm
mv9IWi/o7/VnfO/zKv2X35mbwEKnTH3Ubb6+BoE3RvD1RtoRDyxujdC+PE5M9z1j
+v/uucGOd8nzdqbfrQgyyWv/CBxdsiX2lWUBFD5JCMoGX0sZdxIsPycBEJJQuh2J
mOFEnVDIDJrEGVuZyz5jC0bOggtpJvjS0TkBdBpx6mEY24aKhdg/bZ+4GzPQ66Hf
4mV/YXqh4v8GpCdmhwVmnUUr3IAR8bejzd0jSl/lSSrW/dM/dvJexefEgNkeVvGX
v1oHkwAVAaoV635/c59adC73xl1tfVUecCMwy1knazFJwmx3VCzuHmFenMp3WwGc
RCXeVjZJV2iQ0jhhC7WhtJfIyt3z7H4wS8mjgxjkG/52saVGgx+1dJ/zxu+KF93N
OTahsKtjp7Av4C/ZFWfOHIhd8AB1W6m4NkErN6A/yEm16anGgv5hITJ7JI790nIR
dilgqjtfQtFk0fZpExguiA7IRg+batMqTy2gA35k1LYR3yrbW7juPnmkxsD9rilA
gmAKrXu0ElWi48LVlrAJHTRsy+0tvY8eRFwOAH9zqak9k8T3OgUSHzcWM+YKO7N7
f9dfz0flDQ3pssGcOOJ/ZByf21Ahwh460pE24/MuweJ6wt6ubxwLdI0ONGik2e4g
NJSWX2s1hKV440l8VIJ1UJCrYVd4X78iTC9h4XZ/AxALFG+IZweI94QFxjn173VE
KHkl/G6IzpQrsfnz584WDb3cmcwqGeB0gTf3aXIVdsUtK+Mei0M84equFF1QOKIN
6hJ3v1h8keStS8H9kPtVIz1JK6nOM36Fi48k4O6fZ/Zz6A2iE91xK2XNq+G2Kxth
45HZM5ku9mBwT/LYnZEO0w/UbN7vtXj9JSjtl0sbz49afxRVLlf3M+Ugc3G7ypBk
iSCFomY1IjPSeGCfjA+Un5n86NBFPFtDTpBFLW+uPaTx09HYCnOKuwM32VxoBpzG
1UgNl7KKv8IYpRjJhXZZ7bzA1USJZsfFF2tm5WkVgiC5lKsQWhqaa7IVrwO5J3qP
kGeWFcgPTJwcsrDEJrkKIQau3qW1IoVqpSkkFLlae74BnSQnHZlWTIpfXojdYFt+
2hySLVs2wwdsjOlh1NtwueE6K63ZCiIJo3ad6xkeaDuepxxOUMXvcm+hcRVM75m1
JNXSfysFZGuJ5ft/NQ02Uho3v8enPihEAZ8TXRJdyjQgioL9r5q3D828u2b0GQEI
GXIuzTXmFJ0nQMSvi/1RtUiFuWSrTY5c5k3boeo0NWf8DLQKTCHFUWbyV8zlI7Fj
dWi8IuIlIVu8a72RZUlwKzjLGSpA/zhGUS1Nb6wR8aDVr/Nc9bA9/DNw2kgCG9pb
iYU0P6h66YQD6/kE0niqhOcv4A2xKAbv6M5GGkmUegGuRv82+zFZPnJeAO3zDbWq
0C0o1Rjjj4oddJ65TtZlgHuHNS5QD+SaUyv3prCcSkQ5T1wVVQakizNINld/22gt
tB8tI+qkX48C4ZQiN9kLVrvwM25pjB7FSQe++EGx0ZADsEP3CpsS/F/yheUk+leF
qYUM/JmIUUD1BzRpYoyERqbKGwyCTIE5+18XlZ1Bv9/Nk8SKTrGg3SRlJkGChElS
l28Qs051DTC0du7UecHZOpI8VFYyPIVtpQwY984hY7HfT1amxZgRrTC7j1DjWOfg
mQCbQvAbZFT1UhZaS01Ugz4MCBjkE3IiUVJT9td6X9wI1l+L8NuWo0WyqOolo+ot
vCfK/4eRrdA3kbzDisomTzN0PBLoH9SDqdjnnHQkLbHufzRReEx+arSsuDtmwocg
2S7R7BSUwMDblkNkFEB7mnYBqBe14CPT9wAeitb5FlisgA6dkAAuRegNPTSFEi2k
5C4JdQOObJIK2KSTHl2vhLV0F6hNnzGOFklX8cR78ZJa6VDUF3TWQ8/5bXYnTulY
lDZ61pOmo9oP1KEfVV5e0Qld6N/w1+awtHuBNjOK88RcR2gFkxi+po7zdqeVufVX
expT4ENpNU5swCVzIsiuSafYLryZmi4+sRnc165N/0eqhBp8vF3VfooNr40uRbXO
BP7+e51O/bwK2ZzzpFG6fp6WS2C4MV2yjGAWDIiO7sCfvHDkV5zZprmhHlp2Ez16
1i/4B39NjQPIquXdvs1vPVAHM9Vaj6Gv+yoWmYdEXPzYJTByXm9l4GGYspzMBw8+
eFgHm1kAfkMhxMAr7U4QPtdf5Uqg9BvZwqURfkUxWcMDVNyVlEvNO6Ur2Do2ruDl
p69eOj9C8rZAlO50EtW3HKeOkg3BxeGH0yUeY14XmYkaT9skxB1i8svh5xkVXPXZ
ts6irxURz0SmBFbIObujLnvyaO1CAGCsZQgD4d1bp/Ma37VQbIZgRhAipNoTtPqq
T44T6mCCsa8AMA74ZyEMbqOVMCtrXu9XTnNAqYRHq6eITXPrejLjgU2Eh0YRab6B
6+Jip5eeDlcCK7bUTSx9bYpm+yX6W/cLtKY5sLxGoE/wyee4dQeCa8Q3nnJVvQgd
qOngxidzlKQNveobjSrDf53dV8tRO5YLM6vSXVgrHtWHWD2bee2Qpy/L6w8prxsj
NmsZr4iY0myfEWBYtVsam6uS70q9Vp3sSQZApZ1Y4HMGGIW4+39Mv2qwO6lTB3AO
FaljYcK9u5r3lUFs5+p1BSBv6Tp7UhNYkF7nqHIv1cWnRyRa/2OzSy+p+uuyXp7x
p4I5ciKtTXxT1N0RMjrSIS+s8ucbp+MenWlyDgrv7bPsE4TMSjV8zarzjdQ353R6
gKZRzIUbVJzQs2fjvfOrfxyNoGkfblPUQ13JlgU7qHP7B3CHbwW3Jc6nY3xB6lKS
tdCk/iWB362Pe88wptnOZgsS5UQR3iUAbIm+/l0dtLtIYFTfnn/jqveI2IKgOlWt
wjuxOsT0gWeWPrZx6jchv4yArUDjK/nF18XpYh32NMZRCmiNsUn4GP/TVOiETXLB
Ewn7NwZy0vSZbPNVDZZJjyfrUJv7TvdFfcfxkttuu3ffLBvvCg2uOqximHnydIIK
/NK/zvnViGyp7IDHdQUszcM2IdkRNRJawRhdm10bBe+12j7a5+LAGsr0mZztUsfa
JlMIXC+KVwZlyKUEsnBf7zEUUuf7AbWRk2cL3Yj+kZJo79CTqqBrv8x0l8ILR7uZ
+7lKqL61VqxeNhz+PKxawrLRfsQKwIhYWnGIdwItUSQuEYzvPzfPjaTEnye1iNVr
miwe80wcFs4qSZkQeSxUX5+VoCCs97VHNyIomYB/JXDcnxpTD4OO9qfv/DhUZxKl
ZSdmyf2YGAoJ9AEsvsm8v6huQKV948FgmWwQ5esz0DhgqOstioCsU6EuKWRjR5nd
na/ANyhWnM2eq7eRt5cmEC60YfGewLTQZnsM6rpkKSm3NSv3+U/M9zlj42/anPPx
y01Q+q3aMZ3iFzTdHWgw1jZ1yERdA2YmE3bmHjwmyJII5jkIvxVaYbH0AlgCzjCH
fgO5UfIBqpav9BHvsUz2HSMH57cb1X4m3m750s5gayYAKnS2GVJizvXg2zbf/doE
Y+hIyBgFNla+3qZ1M84uJjia+7CHrfU3/wQiTr6R4GFiDFwJR5wE34wYVWUf9MFH
vWck7WMUWF7adUsN3zBasxl6j4lldf+jmA+SB67XLbUXO/75nnirUssLmB2o9++2
JnPO2G1P/5yaxeHbbhhqKsJDdc6GbaunK0i4XCeqkC4ZgK3tWfkdd/TgnX3eSU/k
d6HeuTHER5PcCk0QUv+QOozXR98Ud41KyG7BTXuRwBkl/QpaVsJqnuma6HiivViA
oTKMadplj55OJoQ/RgnYUUy407t/y0pw/O5a/5eKplqv8ccMoeVU0SCEcT6r3FBh
Xs/gHqrNAJ4YWKX0ji4XTvvdBjtY5kPe6nMsyyY0jOEWGXt07Ns9EUJSfroOHlff
xWawmbWCXQPorBvxAf2CfB6kcNJp1n3lEfYqbYPLDKrI12cN16YQbJcdK7KQ6aFC
zK6nLGb2pj5jaCMYTXzGhVA2y/l5OMSy4YQk0MMQHkd8P4j5Q5/9yLEqP94COPa8
dh9kYchznTCVXf3CHNHVr4ur15OAXRc7WXfDlGYGptpYrUjAzCHUz2Z0Wk9OWIg3
Pisr0SqWjRXmeeE7HqcOlZDs8Aa7P8a8z+X1na8stolKa/RBPD6LvPlsYYvR1Cm4
47m9iwoPZfBqpm8vD2ODUlURC2JwV47DdaAmBUA/8kCUy0DbXdZae6OuYV2EtW7M
5HwD8ZyvzY9bVFeHGSXdS5YXCvTqoiZnfP4yC7zVCUCmhD6gx4tXIviX7L1fnuNg
5GE1bA25uIUQl3F8EreheQQtndhfz8ZBV65BA4RDbuRgZxi0zSTrQxKf4v3UNdha
VOOoK1wOQROgPsy66H7MVOs0jEztvmQbDEVloqsFBzbEZFQahm8aMvUCqEQiWuxl
G0akNpwt+K7wp10bqWnV+MHoBm5n5GC6CctHxVRj09vofo+lmD58nJ+GJHHFqc7Z
lmQ1t4J8FfFEH7nfImVPAgMLyre0S68MQ+u9xVCqHm7WG5oRXcT4v+HQ0p4xvOqO
AqS5OnckIh2LYq9g6g4K8om+Bgc3GMtZpC1O+cW08BkQWMfucfeS/T7T6iQ+nr34
wBWcJ8V4ypGZjT1oJf+OUpopjk/wMk/m+mepVBG8QZ6XcgySHa982x5MApIYw/F1
37r18480WxOvwOUZnBvyMPFUKQFHVVThx0/P6X3EY/tIQagZIwtWbAeRapMS3cG/
GE2Y1EVcXc/ouVpZuiZjDtBSSXnhtBTzzx5UfzuaIB90wFdNBAmUgLbmcHDzLrOF
ajw0JjU5YzSG8rdMRZ7xem4d91kMebDaBKJymEiJopxJsM11DLA5ex1p25Z2Shgp
TJScaXZ4Y7UR0CN5PQPa+Ufm+26EISXwC4qvxp3LMgRH9oicctkX0Q26/dHeFKdd
sR50+KglLBTwTyT29GTFz1uH+42huJkt942wrfYxFeRZJKQF8m36mghFcSpaN4RD
WWZDUpmGUdGpMepQhnBb8ZmFz4/5a1WFfwgzvnfN9zcubSmq3pRN7zRSfr17MvvY
Uqd/h9boTthwpulXNarWJUINbYoTCv8umSucEp/Z2fy4R5o64wG3H8rqKFps/zqr
iwz5MKsqjRyDIvHVw9xFg/tJELaBo1Zed3ZvVtA1kb1EAbGsjguz0nF2hF1W1Dvm
NUqichydQDfuTUltZ1+fm/jPF0rZAkFc0rN3Z75hOizQH1VEPAzHDqS3mo3e1uV7
+dK2OaUkiHfnde1kc5aqIhGWh97rzSnOIso5GY9qJSGS6uTg+VcEVUgPp/5jmtO2
uVeaxsbWExtP7vSNlCa6NqG9mpGcZeDttkBsOqvJx4rF7vpoM+QjX7BxAz7FAngN
N5w24XZ70/UR9kSBgo4BnHdPs2QudwnszQ/IO4ce5rsyP6BCMldSGxlXLnMd2s72
pW0b4DOsAa1DCnxf4CLOBBuwoRaYSdhtHBn3UFlJ6zaCzCGC+N9dkdabIcx8cfZF
uF4tJLRE5QZNVNXGCMjvtWolHnOTBwpg5Nei3llMCVhcILEdny/VIVaeueXrVtvQ
duDaJ0myCmrfAv63bspzpnraCydePGMCQKxIpybmpic5KwmCr2dLnVwU308pfPqg
HKdUWO56IyRLSTsn33TMqYODUmU+FiSZLjae7JjAV5DInOLe+9KpEcyTyr9/PCFz
bFIjE7VI8pL9yRlS66L5Gcnwh1mqPwkeVqZ+/vtEsX5Zfd30u3zY59Sw+uxfq9jM
iLL6EIa6OPKsg9Q2695KOBr1PFkEwZAo/v7UZPcBpDGc2jHzDTe4yVp/frv4tYWB
mIke5rMfUmwKDqagyBRLqxRyjNnxHpaHCnkvMOTdXAICRVCmx/wk6IH+gF+Wgsfb
EuyXKg/ErgLdBiz7kcxh8T0bk7k/iZwXN88Pot6HSKnaIJHIdBZu6a66zjP8JDRy
bRRgVQuVoXU5WZJP6wizdgiuJ0PiFlyM+xbAn8r5sUBipMMIa7K2PIaf3dePhdpG
/MkuKEpDCVwsSbbn6r0oNlYXpr9Jsk/omWs0uFa94H+wFPrJZ7FLQe2XsdfakgiG
hB030k/H2SATDwZJu1EREZwQ9pwDPivE4xsj4BNEaD3a8xa+cv/bUD3c+/oq7+mu
ollxP6w4EEfyrmnKunTuvTvCHWk6BXIZRjICHaaSY60JKK/6KVzEh1MaUS8IRg6N
s57BPazNR5ppilWP50pLLD4AM2QAhTEmX4yRL27GjKupC3H7v5Fci+iRPbPShO6p
29vF9O/IXeqsIYk70FNWx7Qp8Wlq7YtTp5XUPZ/SONvTIOp/pUVqaxrmQSvcnVbE
DZM9s6KRc6rQWPuLbn+zomkVz42Pe1wTlfrTiEk/+XC79FqDXPLQK04A1tJn7yud
xbBuT357AR6evOQCgBJZh+AyM1ckHPz/ATUrOxoQqub8nWhVY4Hzp5ClccEfL7FJ
vhWlc49GxIvMrPfCTYWaNko9RyigEtXlXJIlQ4mgf0qDlvFw7eFMljjweitsqVqt
C1Q3fCfkgjV4O2g9aBzfT085vRrgbdkvuWxMxrE7RrJ9mS8NwqjXylL9uNzSzpmx
cVEymxbLePDCQY8/7MouGpqRP/nr8C/UNW9LZpesZw16dTKVqbGhGT9HFjQJJ1ob
nHEodHYnIAgMyPDaXtPHw2BVY+A71sEPMicqfUkome9weMeZzPwicqH/MirSuuwS
bOHUvxkGYsiziHC6LnFelgm+u50+2gR51/wu+NNMQ0+rrjKv+r9MZ2mr1ZYw9jUq
XeBrZHNU8GIV6df0jNZYa3FbT4YIh8P1nn7tYbP6Rea5BDNv2EtrD2Ms8ou2Jmvj
yvCHDSiDmOJ9fn3LubQY0mnngUVn3ed+4/fo9fP+6DtUyFg0iExmA/D8cRn0UHYk
xMJ24xm6zyxr2VqEMJ7+ge7B2ORg5KvGDBuDh19tezkp0JFR5UVYu1Qnwb8g+UxM
QzEMbSXx2Ht47Iw+mWQUO80BbCwfIbym85P+LOliH9nael4Hg7t2sMgN3KGyRFNk
V2/R1HLo490+Q4PTuRiIA7Y3ViQzHDYkzbkZLe8WsVCaSjRJB6aaI+EloxGT5Lqe
h2Q6LTmBUGBlkwOs+BjlUg2a2mV82lypldkS7RugRTyR0tTHtiMv0o70qcc6xqIx
pwlzdsdSD3+xszlS2XtHF6Nkux9abmKUalrk6TbJDKF9oDwpMVzx5ZgHLzmWV2oR
kMJX+nMmdfvJMLOAC4VvANR4k+AUGMLSfKozmWOmnUUCNWvBaOztz4jmK5UeHZJN
IcwbcUqvXGkd17DjqCFOYUiO3kDL3iFYYBR0SIHc9N2spKyCzHARYTdds/xTKYB0
bH+qkZVMOY94yL+/PDMLLX6eHNIDYEboogFlqCvM3Y22AP/PwI+n8WtMP63ARmJU
tpGDtAn/EHJr3pbvijL/v3IZtEDUw3xBB7Z9Swx9+i1DV39iyi7xGqCvxunw5OpK
QBwprcSFoiXCX1W9Umo/c/0GrtaiEkIrBGIdnh8Jxp0HX9l0UEr1R5Knl1FL/Z7x
5fHdqSEWIzo/eMI4BB5z72O1oPKWaDuJD3928QPa9LKGWoqFGx9pDMJdO2pcSj78
RVQfBkXT2P4yPGIu16WcdFHwiONNDnS1bG67XJbijMmSFhbhLXgx2Nl/OrkrGuS/
K4ncA4h1AORlvZMSSa65nNM21lm5CLvkfvauOi7cGpntYAH2VvIpf1fZHf2PtXyn
EuiPnfgv/hbcAmZQHSji2MtImA3dhxUhgM5pzd8hbVtqpaagyZ+3nYXO8JdYZSq6
2/83+F2ZwG5/U0B/gNZwxY+TFa/o+nAUtoj1fx07OuzpUjB2JzGSpkolkP8LVA78
XwrStLuS1kSH5Z28ltX2ys1TAZ2DTQITmDBH9Dta2XcIND+WO6vIzVFrqX8T+1I9
LWY0rYzx0yKjIPEeAuxFbPa7ing2B44qis5TZMgq4nZhEo+UF9dhM7hgIpKS82sS
3HWSQq0CKo/axes1u8QD5PKSrSKJpwqmjQZ625oE73yRZkfa4oTY8UOYEMIW9glB
Kttak7wDrXQvqj3Pi573YrqLtP65I1frFUbpO6kBbeqc67G91we8JndLwTDLue3o
e2V9AiBu8E85ZekNCM2Y1P07UP0OKzU52Oa1TCEmw1WCP96QmkpVzd+CLy1c6eYk
D16x3+/9zdR6Fj67YPW7y/qFdLki8mTfWpHJ5PFOJwntGVL1zrdAfBNHOkeAow9L
EV8ChgaKpKCzbtCDk3FotvHracOHZHtLCLABQjfjEZoH6JwlvkmVzRUkAFZb25pt
bomoef0YuRhi9g0yJ0OjzrePSg9FMtLNbOznDJD/vcjk65pDnVIzmdwIhQyk3/k2
eDAzXXnGLPTWsSeO4nGPUgrnKUdgFV/HWABgG9VxeS7Xas/T1wiJuxi3CgnmqOlO
qyNe8lr++QghL9z3qcQa2D8saesUsV0fau4UeZwIDZQgS4Ac0HuThDq3C6lLnbhW
dr3DxMziULKso5jrlhni2I4hn0PRIjdMWQkho+shTXmUxtU/1174rqCAvweiWDRE
6vZ+kAZkA3ObW40DvzThsS9VXptQs2OGOhM8FEuNYGkAeIteLSQnk1znQreC+HQr
e3J7oKG3IwW6S2tU8Yd2R4r7KD/ktPgxwV8lc9xsEeYxq9FImsV9nT+4hcwl5G68
MlLERz8WdqU0c7Y3fmx9ZLTTSK+zUwxmNTpHTbT7HgJ+C35cye+az7Z0h0k+Dsm4
jJ7fzxKUbVQEzkRMJzAw/j/uToL4XseB23zBCPKofGnXgavoPe6m6OXJYwh41VDW
j952h54OAgdJgIW409hNjWaZqnRsOe7To69g2r4+yhC3bc5QeE+uyPi0RUP8A07l
a7y+GOKJ/fGnp0GxrkL3zyVOrPWin+mXFKqFJP+7BGGqLQvR55zvUBS0kakq9cap
Mc4QbXLYxgi3R7P1JNmTIFpag4YRtlBTYPE9KEtQzof3eTtAnn+UX5mnkz+TlY1U
QMEFe6Cr4eOGvCcw4xBjDGOSRhvrNo8XxmVdYCGq0bVJp0rKfasw186e7Hyss5t+
+pAW/WL1VLvWYnWYVgwfczTSluehqV2i7qB3Sn4BFduBeUYL/21XRK8Ni82XGtDo
tsltwgcv0QVDvZSOzTLF00AmhTE2/AODNmtktMgw0X62BaftkFv0ttfa2gWu7yP9
casftw/nkpqFZT0VxuYqlJL0cDoaH15dy91k0OBTZHYdbbYtmm9hDjwk56WfMYvg
6C0mHYl2hmm21c8MBry66emqeEXDpxHx5jowd2JK1XuKoJ54hJqFrE/cmS4re6Lh
mCVkWSVn77BmmOp5rVWdVTKxBfHTyzrRMCz7Vs40HJCUt3+Qd1syQdRzVufhp3M+
pK50SSUYubb9LeZ2w2uQ7/nor2pQRIZGcoyKhz7d6U6l4GSt+t4PrbGqgUerdUa3
c5CpYNhRCzCqwTFeF+12718kH4aM6qDkbb80aUl8e+QTyZsv0na8oJz/SUy4k8u8
GVV6oNo1xrW4U0EtHwZlhMsi9rXOsX45lXpDepxMo4nPS0Id54PHCxneTNP04V/L
nYdeE7Ce1CwFESpxHD8IIdCBGusEQmtp2+wllpVEudaj3RAmmjZQ/pR9iXhlctGu
LQJAGkcictMJyW38/oAchowehJfZaD9LoiNHhanLnoSTwdGmUJM779iIFmpJHMAB
YpFMzpXA51DfQl18njOUw5ymb7w7BECptQtcEjiDUSwx+DR9ijR+32UMjr0aqEMQ
yqTEu7+T7Z1RJleQuT4nej21QNtBXZ+ipUrXX1aOpvmMazy+ce3eLNVg/g7rNBPL
u4UAc/kUiwXgVfzjLv4fJonbfV8mIWprpsz3JZUr+VZ5CguRh6V5mZhfn9BQJM6t
CfzrhMEgmsQaieJA6vbkSbh6s7BRDUjUsYN9yTHlpxdtqBtGlBiId07Q8tK9zgav
/GaPL0lJ/ngVYje4JUiRAYi/qx8+4SPo29UmUscMksT6jAv7Ggy4CnTIS63kzQwj
+PTPRdcfQCvcsrQt4u6ljtCudnwBRqPbCoqsGPSVFhAbxP2W2AUCa6HEAN9MDtAR
K0lWoTjf2VKpHC1aRp7hGU8GjFIa8NJyC8xrEqKGetuAaHbmNfptKHesjkbMpIVP
Bm8UGhTNt4OJyUQKEmbbYjOaChagxrnegIMTvfmqDPoxdCkcf7kM4rzAnXrbffob
FZlIQVUNAdeJ5BAtZa3PDoY3J6z7HKzdKcZxMXL6jHCSgDF+36PPT+R5TlcTr+9H
QkkLR1Rim8OGP3a2oi5Ora4n+1birQShiXYO8p/JwU5pwAl11zMpX2FYUh/STpOF
Linpy9DR8jp4Tjfnf4KwPjTsTtX5nuAtFhRu8ibBh8PWemkPT1IejxtzCOzfDmwi
p81RfSqNhEE4zsUaDwbYKLsJup7KqJMzHXZjx6XtojbWkGx/4gXJAIvukljFxIgW
xOAmynK4PW9gEFR+ep/esEr9TdtnZM6oxK4GdwOzeCR+RlySQCDPZ0bqDrn1o7F1
Y8a+dMcWodQZ77eaKBlzbmsx7D0klS8Yx75feVqr7J4GeBOh6FLiC4YcgdY2JuDi
/fltDjLM8n/qohOcd3goBZe8TueTECSwFtYAe8zf1kvKs1LmWcHZMuTALEWlWGZy
9kYVDL6LHTKv/ZJJXwCSandcOubRrFH3Xk8a/kvVM+KMQ5ly1EX3+gvY3uMJ3BIP
PJXoytrJRtnLe1NQXIbUwjXNMsnhZY4AYs/hW0Kl0NLADyPLUuI//zQuICTs0UhQ
E1Ph9Of8CQRpMk+F9mP5WFRoJPmGJ3OwzfMoxgr7ygPVGwkCEjk29Q4UDza6RTbu
rEUQKEJ9XcOTNfJGEVkZiac0z4dZt7nabbR6z7AWQo0+FuZ+c0iSFViHuYFrX1eo
ApXB+Xk0aj1fU4lnmUTwxsdCL+Wn0C1HadNoWZIMlx/v8gBZyc58qoAwTdKFjL70
rL+qSSD7B11mBKjFmqon5qbfxye42cFlhUizf1X9OeE0Ba+if/0TNplPt3+CfBRA
JukITFYP3Grwml/xv1Sk6Gj9zQYzY/rz227pKYG7q8GJlgtkc1MnPmOhCPGmLoy6
Z6TtB+vrXwDpwRoR5ErivkNUBlsomMWwPmLyjLpj3BIsWkwhr3hHDt15KOeSTUuB
FqviUg48XEToiOTbqK6gcvt3oZk3Ok9HNHLYCAImsm0bHpHgqhZBuS7gXcN5mFbI
6mERwmza+FpKStvGmoF/JR6nG8hO/7BUC168JJ2pBy9TVJH6zb79UXLRfWho0a8d
1W49MPGWjbKlyE1iR1C/XeZqXoIDHwkYtlUUt9dI9BeVCFrWKPEBjZM1t8Cx6GWR
lt7BjStAdXFZcbbFnTupaafRuZbwnjw3boRbeUW79dbQ7jDYkZlgLYmglK52D70o
0gdK7OIW3/AgwkURZwk8vRFAlFnZcrhTrGbz74SiGlsElH803KM+7HC889+MRQ0o
v/F//mbLz9tb4Bbm8KyP6AaeLv+TdBOLPTNN4E0hNrVleigg66U5TwxTrHKya2Hh
tIciSY4dHbhhm/+1fOkD+stmSAZc3YOMXXwwENsFjX4zLH3smQZGukj7cuJF81lT
eas/kTishX2ktH3UAs6fHzlPfoQTEwYh+jMqGRE04ufyywH1OLprqeGzN0ynltkY
/3IqHcv4XwG2ou+rNbFOmLNH1bUJ6Kcr8eg3JfbkBJUY/YKe2exll9/RCthkTFkQ
A+fItjihs/UlbH39oCGCHB4aArimsNCKz6UxHZ+eeXis0dk0uZYcaYeAiz9iHzdP
J7TAHR2lYoTq1Z9zv82Xl/eh7tL6ZJYC7bFsWa/jbAnrCwFCLEK1GRybXgw5a35z
l082lI9tviQ0g65BwDrv97MfzkqR6SVAuTS1FvSq1wrUXvNhoiX89S3le1HoK8Cp
X0G9W11DFKR4s/qqWmzswRxxqqMFfqqsimJQvIhVTVScY8oiu0DHUPuxhLcN79cG
7cabWYUgO6joAwTbXCG+tJ1u4vm8KiX0btOo7en5IRT1yAhTPD7znka6nTxGYrgw
pZBvmagOKb1+nWlLsUQwUkwQrdBkxWUUBEXVEIZf37boSWGIVZW9mOqHhAJvoa+g
ixfSOwkPGbbILpZ4rBm2n2FLqYU5edgerASn/NkwTvmXLbWxXqzdb1XSnch7VV5L
KpIfAoZJXfGzE5obEe+Wflh/zSwcz5UDGOCKAiKGuoM0uy2CnN7PTc2seas/YMPf
0e1P4bCYPNGWplVV/M/BbnTIs8mK9c2Xj4KYanok+x6ix8FMDToWH5wdcF61mt8q
HAgLa+vZwQ03gdA5icbj780LipVlKPq5RNp0snaAFldY2bY67R1bZ1beSHzRpHUH
EHDc3K6eIIoRTAwoOOeTh4pzRyjroSCBpTFFE1gf+OmO7rw5s3t47QsWJOOBSthO
O19yPLL6HW/Tm1aOuezS+U2+RqBU61yY1f8HnDDL5YUhkpRKoa4yZkW9MeVresvC
bELdftPaSuBOBSCcxpvQZg4NZsCX5DLGYca8XcxEGpcC+O2Q6KzVV/mP6r7s09Hb
NwFJk9xQnuolzR4iQR0d9SbGnHTFOaeORvx6o1YK6YzZbXGJM9VkzPzSTwmDhaDY
Zm/btTvsRbAKI0x1b5qTUZaOJx924red6KIwpd8EQP/crSyiQKY6vMDstQPkKdlR
8fzM8XSjpkCZVxMpwLtrwpslsCNEpJ4a1J8FF1Ko2/bWVfwCUdSR1XpKA9l3xIeL
URETtX+4iSh/xIUpHw/m7/UrDPPUBdbe7nerkXz4EWnDIdOg3E0PG2mMZj0GCJUO
jb25O7ishvdCl28L+0yw93pDYFK4I41y1onCMoe7P7GQRAd9dS+wIOKQTH4s/1wN
baDLlAdT7q6Y66J67wItUrUD8KjfpAjod3bL8GJgea+cD2rcZkV+zUwk72fKzZSH
z+lvbcs6w5UGEBPXXLC7dAkta0X0vFzxToxyKbYi0fwNLr314O9R5Up/N0abyhsX
PrLJCyJxNsUJgX8plPFdvK3vQEY1kuZ0gTWsOXfL0DPL8Ge7u++1baLfplbStj5e
yuzC1lC9r93Ryh1xhaKtfJr4UV63f6llMT03Qt0Lnv7E/XvfbmOEvBEht1HasxFH
ur+JKRx+nAE5Wl7SJFw/BglzpHWjNAqNcNqZav/KyZcMSfhsVGVK+HP9YWZU0v54
zQFTtvJKLmUej924y4ezY3Bkw0+mYqyJzoRL3nMGhv8qyM94CXiYmlxTcsq9chkc
/Jx6FKPfX7SSng18LONEpGz8ZvOl6hUJqrNiTaxhRashoS/GIuDBZhxhOnWPcfXS
yNiJLsfD5Dq1mH6aAe137p6wvdihFb4vMxbQB5Ih5wYLirDmPmHsaddBzxlgnJFB
8aA2tmxLPtKr9+mpTPDI2JAyguOm6VYCHzkMKKToQ5htNdkIcxAViksRW9IWZxQV
FmHdsrOGV9W1qL+qKRGkq6+TWtbfjVPRVzTTo6iU7FTKRgRMZRwRzHpwiw2+xwMn
tDb7K4x/pJdc3b8lAt4mqAQ+t8ewthYtDZ1UwIfXhMhnKvOlewB4tt11H7WlEgRo
5LFVqaXgvBKiHsEZMoLTHSND/Z3dUpIu+IowJx22aOEBpVg0b/eGtgQHOO81tQZn
bs7MSyuvcnMCBD06WJUJ6a4dQe4sIhrqn9WK4B4qrxupQFrB+XHeQlzsOjIqcTTo
rRBQWknjrC0suh63/0GRDbf5hc4Bgzq2D9Qe8Da0USkIKLumTj/l3A31bn9nOhgt
rme9U5pnmvu+EkKzwLyjPeisHuJW0pgIctSOh5Xf2jKj/DqIoHaUQ5UbZzieFTDE
XW1VEbuS+YwhNSenW7ij0kPK4avJRljqiXUdo/Rdbe52Uc1fWO66kJzPo+K4jfxH
9Vx3xjyxsKpftyMA7ZYDzvbgSiAhnjudYf7P9wugkp6OhFvpwDhYzhEc7SWetesO
JhIkj8AM8ZKLa+KyuCsMOwHKmH7JCY7OfZKKC3/Cv0vZyHK/tOwm4K4D9ZMYgu0b
5L0FpGfd39D8GDXkI7uF4YX4Oz8sY96LEcm4l7WXDi551W7yFah1Vh65mfmQYuP9
x20sCHTOGcKkTp5yO3jtex8DVNVGUZo/3poMNz3+JZtivGTryEC3gUo4QsA51xud
7lhEDQrDAUzPFHqLMQZzh1bFqwrjKpEazgtvzsnGnThNYDjzlFvZoNrAbWXwSP/c
DUanolqo1eUUQa6mo/6P91pTfcOQrCQguTsyWftntC9Cudzhtdpo4RmZVP2wT3RC
iYNVP34BU+qZ0b3VLV8nn32QSvQoy5KuNty9/U50vb7EGVdz4Uqt2oUuJicbwAzj
stOH8tQRMxMZaY64NrciJkjY1pA2KBFTySq2jdNFdX+XdQ30CcSF6KAlVgJI451X
mFmPXG7a59SDYDvGcGZCgDQ1zbSbJ/wi2Juo1Zn7GUb6cVJLhNH10J//mJuhXz07
9ICumEhh2XQ3t0UmXYjipA4qvpbLxulpMCpvtLFVjjeUD0qMxS3KZdqC9w0Fnz3K
HNs34uMWEHAA6nkk8RhF303ChgYFXrVYL2Q37be0S+tjPlAuK5dnnjC3iTOqZnwz
XpDg0KEr2phyjSg2HT1Ypkr0d/RvbZjndyYDLP3/nuy0mX8oa3FjzNTiZcCDVIka
Mo/WpbnxTxTjR8khKgS4zhOIr3K70M6dJVGDkI5Am/GFI1veLBwXu3jiwSFn9i/j
5amJ4xvrSbuXDQ931aAGwr18k+OCJ35SM/0J2TqV8GYU3jnhMVe4z9OI8FWB022G
WSjCofMEM7ogsfTCKHRabQ9XrE713UmLQU/pWpHHwNeZFvetIYru8p7vL30dnDx1
6oFpU9wjZIl7zeVVG3ACmDC3v2ewwP94tgkBj9wIpSDs/MbvIrmTYGLvG+DTCvT7
Nm8onRpO99LKLhgW/AUlbaJfg3Puzw7UK6Rawy6FfrApViveyWg76gWFONq97RgJ
DYcbKloXnl2sFja7A6gcep4a+s5Mb9MZZJfP70UUsG2FmZEOE3iF5Mf0VBrdP8k4
iynpECzSYtb6Oe5zqp2zN6l270sq/W/mjX98atK4luyu//DN+BiyS9dab3fY/Mfk
lPh4hAinQvSyR0Ksjx38WHP/EbLpbj/L9Zq41Fp+d18FTsGyewC3GbxI0IvALnf0
iWKHc+3hSvvcD6UvqB6nT5o2cDHX9HMIL/iAtOUZcnlBjSnVeQbJ9OERxiLm4Oh+
mfYPeLzpPnsUUfdREzjJWRHSvoGvoDlikkxt2pqb/1q3OT/SSEadwIFnkLlXGoqc
XoJCR/80jYptYwEJSE6qrHD/NV5icEV4odz7jDrn9z9KyJ8hc2YTIxpBXN1LiUn3
kWawmLyxY0dwSL57oHcByXIKzly33u1Nt50JJjnbswAnK44gtttl9Q8R1qQK6+vp
CTwOB40QlXaIWqZHzgO0jQz53hfMnZPMB7/szDiDcWcKZfG5K4CESn+HWqDC+E/9
c5Q8ANenST7cpX7yf1UglU1L3zlIJS0sXaLL1j1MAOfPGSHt2bBH3vcFu/ov4CqX
ULMZegi1sLuTlJKnZsZbkHn17ElspWTnA6GzAUc4XnEq5LLZG/v28i7+hsoU2qQM
TkQZQLN6Djs1L9/SkNhjTN2l14ZYQxvY24tmDtqQdQEJeUaNwMQzrqzkfBvLO0EG
vbs3BirEgaznGTTw8ToAX8sIKW9QediHT8xA1nY4W4drCSWxYSVn6H5vauvidOuq
Jet6ChgTH0vy+i3/fLbPDfoMDpmCMcYGf9OmCpGBjUt26pixYJhZ4ah4sJR4ZzWL
SySXKAYGbuGAMGwVpMLjqlPkYQ23uI1pknUEUnNtU0BWEApag0BZhWm+ZoQ8O5M7
IWG/zksA7LQile1F5POfF+Hl0Y/aNrSZAS0XsnwfXo4P1b+HrWH/UWD7EoilLYdG
bB6EWcxBxqQjz5lu8CS5GOsPCmZMrPcVSBobxQlp6/BZvw6dWTj+uVoAn0qsKaET
PXmfkzOP8AbLMupbKp/TnG9nn2oJqPbyQUiULhDyXZ+oUbcB0a5Iq/KnOFaAkARi
7BviP+aUGan+4s/C6LLEIVltsc3BN3ZRvQoQ1gW5PCz3dymCDOYTdaOCsVCmlnO+
NONSawlqh/6+ZXYUVKh9dqWfEttp4QukYDwAV6WBjSSmj2tsFaqYOeZ95Ml1x/Lf
RO9HcGHyiZ9t0Xo/VvOe9mssN7OZnWO3JeSPjq6kmVEbAHSM0sWiOjMkqoKhvCBd
QRL7DTVXeOmTVEC94PxzvDtBcbZm8AG9yZ+uyNwBJsGYK7yes5D6VVzyaqg8MUub
iPxmCStHv5D/QYyUvNsqLsW7b0KCrozQ0xY1LP6bT4yiI+u9shgHeby3E3v2SS78
NaTt2wgPa1FQF4g80KAiR6fYjsESKBR1wSIh+cPL3hRnQa2+cB4+/SLpHsAxUlg7
dCFxg5gr2dTsIxyJKPWvGLZT1fMHOKbFotNW0aEXG2FfN+dWbLbR7q/QFdED84YU
WxqN16MRvUfmGgAZGSWlgl82hY6akB2yHeiZC0wX6qABSNe6sqRcS+bjHIK2pIo9
lX3V9d1UBubgk4LGwTkq6oqWjk7SbcZJ5RfBGkDS//H7lYDvv8uhbM54EIhV216V
Np2KEmbKBxaFd8Bcj2PRRyjJaaqoOHfnjnN7GicJTn3fxUIL2/TyULPU4XSC7K5a
0YIyoOtlZaCyJ0AgE30sTyEzQHrx/PoO6FDXqxpey8sAfV0UqSuStDbDRKXQ5m0E
sumr9wNlfuyS4rTOIaQAjyXKEVMNiJke3YhNQIq1x2UrRt4V6p2mdczvtrKAp6d9
mXNt0wphw47m6Z1a1PP77H/88StS+7YOfYMd1OQZxnBG6iuft9Kfl0ZzT1HQxzbP
SRzcv6Ep8O1fCXshWxe85uSBoU+HtdRPESSg9QmcMBftfEoJ34i1kSiNkQKXIyjT
XDzBY4T/Kl4Un8+zIPfbu7HUZUyA9ijUOeK+I74X/l6pPSf+r2WljKoIP4WdJ8o8
tczrWBl8EEHpY/Nvwvr/fyQwfwePdo71SrIx+4oLzdnTM8nmVCGHuoDL/4GQsEYO
liC2qOCQm0y9ugS7WdpEnkNcbq1TVyi0I57kXjF0RuhlH8e2L1Hevl6yhHlcanKb
DBCj6m7EJN4Ipr536zp0r/TJbQCWuUO408gTz7Py23XAKfaoPVMZj+sJh8zyVyAs
E3Pk0EzWzkbUOnm2qwQfMKiUlpAmps+uD15HhOvUZFuceZddW6P4oeZWm8FZmffr
LgWuxEKD3B81HmvI9Ww8Slg0wl/wPTImbKM5W40CSxTEHKfvoKJxm3xWzAGeqby8
KfvyZ93nDyEaw1Xe5eQUAOe1Vg27/2uv63k+oS1EIVUWLRy9yy7vqb4pIN1RqcVU
gOhXT5ExrydUjGgbge9WR5EoyvXghTD2lQuk6WkUA0XMdMmhrfSWunC0TTG81d2e
2hBmjzhVVXhAXTMSguESW/ghkiH77cVRmOelacS7jMPw+qUm8+PTSMpwXFZFXX2A
psZJhAZS1zP81r7gxWDu67Kx3X9PSKC60NWf0j45py46pBo6uYQPxzyNnFs/AwjP
k7Rjov1nNwRa+RnLrIZQnGcbAqJ46QIDZWT9nvD+Udq+GSzZV9yxamHjurTSRgW3
3tz/Hg+zioQwu/W8Gdx4wFazVehCk6ej0EDKlxFjLPoZmIPdb3cHRNvzeqPBbSyb
yoOYqZN/xdY0gyZY3ibUfRoJRw1nguBsyfVEYoZXhHoDQiHTPa2fqTv2Z0Nz+O0l
ZbPc7H/ogA5KgDM83NqzKzhJs8OIcc9o5+AFy0bpNr0bS3eOf0rcGkCdB7HeACHW
aQ09VnXg1xort9ftaR2fwMTuEUWZEv1C8FX7mvf/2N1B6WzpNZxXb+J93g/KNbAf
naxoDQ2FX0Z76bB2+Lde0Y/Aa+RzDf+IuA4DuK9kEwpH0YJ76xAsSLFZv19W2VeJ
uBv6jMWJvPFJDpMn3Ek5D9fLDJ8NeBFRB+I0ng+5sEtqpKpDHdcUzG/T3RBhXkPo
a7oiyje3EkvCY5MR9Ixlv7NIoxMh6EivRPwqZpMfqL866Cyn5u9NY1BgqFgZrVPw
zGHCrUfdU88G8qaL1tdrL0vZK6qbqseAUExlakynrv4imWiPxRYhogEvYBDyTRA4
F1gjpzBsLY+8k80v0YDkuDTKZu2CEX0hiNMqP1Uioc+wYzfOd73eolfFOykj9FxJ
jIxAKrhaJ04IsZ8nFR4SC5fZvCfpOFn9QdYuelwrAqMbh9s07RrRc5SyCd3s5KY8
q9XDu0tEIcMNLbhZerjzjtX/Uy2BXtvhBqwqTeZNb87ekmAsFjMDc9IUy43a2g96
8eoUDzh+mNAKrP73thw23f63QeCnbPMIcr3qjvpPOR1x1zSsTpsnTsbT9G6Z98yE
bbzzNK69dq4RGMu4S3Eid6TyD/n8cSZzTzxYAT2iW2vUEagIT2M1UUtQgSsdgprG
zXC91uStmvFPGh06cd3UtgyEza2T+q2jaKN8ZHfwZdxue2Yd8rIkDaWOhywzh+FK
bjoqxo/nBaY/4ORQIPlWQsH6JsmuickJUnGTgG0kbD47cSag44NJUG1vzMm8OMYK
0v+guOIanK80if7mB6JfcIgjdlfQ3sWfr/83Q6qnthVWuHFaUxp2HeT/FVBero0e
0fKDNjArO4Vv6nL/R30grS+XvLvf3tspIb/Txskmm+qQpzA4X8j70JpULqT+WNv1
sIiU7Tibg+IXwsffPSXaWsnMxH01JiblbhKEyseYBvmPk5ACsQuuvo7VNQxsu2/H
uWfQQyOJblTOd300uLh7HXFfy/oBZovHNZ7FxURGYlRW+5KnIJG9nmMMM/uWzl40
aGm92b4fQRhBINwGj8XR5IHS9yWNJE7ZMGY048tvMQffItdDJX1Wi43KD+rFEr6l
OmUTFONxmcCJkW6cJaG6sM4NI5Zgtv4QEWYnOBPjCOQjQAxK2UgvXNFQI6L47XKy
8Jh8I32iRJPWPFPVh05HrBY+MGrS1eiaRQN7Lr9b+NVeBJ8ptTPnoOOLgXVKguzD
98I6TbKx+KUABsVNgne3TjYfgptHXJ886YWPgQw1r8tAPQ9Ft1LbMfIUJylu2EWj
VaTd9GcJJ0rmJWWdXOZ+3QzYXvKZHTHtGBbvgXoX8z4NkNTBjXBFJx+h085DmxMZ
tHyTK2xpt8y8sdhX08k/7vreVaRE634IrPVD2GOjq/EVjtd1rLJu+jkJKFzBzEeA
oD81qfT3HAiOpJrecEUko/rb5OwYKNHD1k9kzQtqf2RMOcPaitOoSNMlwKxi+6Dx
FfKm+DFDGg+myD72xQw+DFoBH7ABBLtEc5on9KUTOMI2TaCHCZicX1NpAA31OJ3f
b1QK6/uFs8ZGh1G0PMli3VgbDQ1cmIaeZn19QLEwqsQXxttS7muH6uVHyq4vsVmd
ANiYDu4ekO9NCEFXBqee3YNJBY2eTCzAX0AA6Ljxh4C4nVQrfGw9q3u9+3AkdCI+
XRcad0aaaqtsi+kINWBdje/sShmA8kt9dBm8al/pS04QAEXu1szPlx1gpBGBFXr6
5Cyb079UyZVMHvVAt1DkBgvTP4gx74z61BUpnbM5HgRXJj261/UmRu1FHI/aNBAY
jaqIgSC9MpNoaSyXL0KZ4ETCcOAF0tmAOHOt2cqWBIeu3ftdpx/WB+g1aeSbQ0PB
K9lizNN/me17wrDZ4CUhKIb4I6UYW7WrSh09Bav1HcSwvEOWUojQawYiL+j7Qxid
K6Qg+adyRhEmc6mhI5ugJI7qr8kqVEdKDPSx/pyKXQGo+igIRFl6njncz61VJSdt
NWGQL3+iKZ2eZkmj90LIFqxgTL2feMdNwtNAyS0EqIegULypUp3WMdwmtgnGwUnJ
k3MEXrjGk4k43IHmvaKv+/DV93Lvk/dbhj4zW5WpRscf3JUXR6SWncvU8WBLatWY
Ks6QuAvrrsdLKQ/dWcHkQSMYVCrcj+i+qG5n5sV8ujRrpGNeaHtBCrf8hoI+mZVl
ov8yVaWi6Fnxqy3D+qbW7nZQgfkGAZbdoBeNew/mU2KnvyPY/vw/jstoBImBI/gM
GORkhAqICwkGc+sTPFSJsN2QcQV6h1Q2xCX3OV1igctnvACb6MWsycOxb6unxi14
qqnJabVzCkbwawAoCoYE08XYXLdv7VNQDMAhK6rF2BQPruHJFz7GAtUcVw4632gh
8Mr2m3rlsykcP1OleikCWTHEuDXnXpjI0LnbgzRqSdw6c49NKrSdiEE4Vpg3UqmA
JeN99OygyFYG9oJ95uT/KfyetjIwadICt/eP0PjNXVo+7H42vX5uYl9F6TENoAap
I4Z9RYsS1YyRgsdGXxXpRZTTE/MZf/eRNlzvT3dDxCqR/fOK1yKyPLvszCwQg3aw
Vd8KzMuz5inhJ7cTSnqCwWyRTpRAVovPc2TlReNGmceY7evWcy+7qsLoAVwAzTXk
uV0dJehGg9Cl2JyMz8m83XErR4zPGEY3tgEUmJvsir00F6LqYdw3zm7DJJfkQgXE
hJVStAwJ3BViJueAZTQdWmor6qNEeZg3GtxFShfQWo5pazzU1qJkxPPHvDXan+Xj
eDixKIHwgYiE+UHF73/9LGSrUA89DjG5I1KLoGNaXmPO1SBd1ypRia8nKNbkEjx3
lH+ZtBG7vgGTa83fgsqpl4u3HmMBWhN7MqwekF3azs9s6XO6cg2JnJfOdHZbpdIq
wjjpWSCv33mP8wHYNXT2A0XsOUZO9p03Vjf4Blef31Xx9It5T3VP4LtfsbdqAp8O
0Yfix3WKXv9d+KGrZ2F1i9bOqRk9EmJRuTUsIcD/riEpIY5ofz+r1Idw2XlyVWU3
2aiGNvRhk7ztv+coYrUc5hBOxeqSf9JBAgX6jJSFqyKjIa9zLQC7tiVu18oAU0v4
3IQ9zpydJj4Tcxj81ORuqSkBoi/ejrEDcN341E1VkCAOQp7NGQpXzU6fscDmc6hA
Vs/XngEao3jIADQT6XQgCL2Nk6OpJ3OCXI++NF+9DwhG8NC1AJVg0v8SkBr0pQej
OL0piHlpR9rulUww3Wp+TRnUMWAiYMBSmXnSVr/Ttk6ZBoT99CpZsBEUrKK5j/fy
+vFC10ktFnKl4dViC2UlFmCJIBH/RvMMB+RjH9/nVl6UJipgurZdkrWVKcfUSvvb
Kom0ScwpwyKF1x8IbFmlUSMCuVvG3XMenUU9QxkNsbQYzJrIcmAZ/xjPbnG8+0tU
Dr9SG3CeaoifpbfuSnEnJf+MEgETJSuoUWgIjZyyFzSpuluUKlE5dZiuWg84Idt/
cAF3eadtKEXnIO/k3tw6J4/FpDZu2LxbWwI5me37LKsjM8ZXzyN98HKP23tsDPNt
w3sQcygi9J3zTy+kEy3t6A5s0otiMkwxTeGVd3q8JJlNleSOLAztuIDEuVSQE8ar
hU2vH362iPj/xnAk1qcqA3eBQUGONGjMgiv0xIdtAUBiwtnjiTHZf5rEIzmYRm3U
xqqsDDmORVOEX5llNSTYbbkTTc7TpQSClr1GCPDXxxgoW7BNVen3OWbmx6LHnUpW
NN2Tu9qPm4MLVMLixCWLU38qvSAy/9lvVMW0pRW2dOgO13ot01WJZuijNIA3AiqU
PBYE1y7lt7yPHbjQmSvnKeZ2oyo2lcwB8/xMSRmamZZhL5asfirxwxaQmfwKQuKt
0/K/2pr81z6cD5FdgRbNJYfGNCbzlknnv67VgDRU64o2Z5pGTEhvNRHGPAZefP+l
M5QZpYwacQvocYYN0tRSP9IE4hhRA7vRUAHLuGN/GmUqE7q5haXx8lHbRhJbOoAI
M4qT4qern4QNqK+Ya20M4lGarrbhqiGMbBvSiuvBxabTcKV1hnsFOkTQ790SOoVl
8EUXVKPlgig8CutBfCHVJcWFn1niBETJIPdXxYWTbdVRmM6lx6YytT6ASw2YXC82
rpYV9n0Nb1VWbHqLhr84odfKWcu3d1Vs5u36gOknweG6xAEPKZllOagOa+DW/yHG
sjYIkVIgcLeMjVr/NBELau1Leey3EixvkqB3lRzT8x8nqtRWfibD+QHaL2jOWx8/
h0l5n4Dyzm09FzpzeVScDN6MjbDbuUfHv37CoRAzevi60oIkBqsKHe6xymA6zqvz
M4859Q7s7Rb73ovzTvEBUw2L+/IhgKZEf+G1axI0uD1Rn/i8y2bHFYiZbPqW7Ozz
OLU6u5m47eLgp2POB39HLfK2SOB+TVaOxh6AA0Lv5BmVRNqQ9mimE2e48ZtCS7M6
Aj0GtK/y2tFPUZb1meDGPbLRdV08oo00EykmvT8zQnRbBXen5c2E4y9yikW4/y5F
2GUMQEHPch/TuvdbYEODA5YTspHq1322NZt5DVlx1KBaTcaPtMHPZQtUVqf/B2N5
4aGfYI2WZx4jcrCgFFBH6sbhBhMUgyuVTJHmlttQuBJ4W2V8VGyHeq6Ule7SJ+iD
VCM/en5CU1CclQLaGeC9mkDtptS05n9bf13CYSI/gOXIvhsAaUtk/byvrpxnulE6
EVBH8OmHwO+XHIuOzjKjaOCUU0gC36Dt3Wiyajyrh4PplNWtH2M4PdP3Tc3xg40o
xqJV3pqMWU74T/QvtixHJ74rCt1KOgTaztUYDcKCwc9StkZIzF75Uyc6ogHCy4Gl
6Tj8Fvh1frTLpsFBwXUI7iE8gNppWKtDz11V6qS+D+j0lr9b/k55RAJmz0soiEz3
NvhKOJJ3n13BJLhh/s6QhdSoLC9GN6naU0u3lq88JQbJL9uPvpH+06X2ZgmDKcu7
xw2ifHv5VWOOQsNXxzxaeAfCeuHT+bngZc1otMXfCSbeop/U/Ug8nFwKaWDz90JK
OfIdza4ej1Cl7iGMBQPSwtGrr/vYC1Li0tyC+//3CQE8o4lidjd9EHUsnGE6oxVJ
FAs3o26TAy9OZt/dJpouRdyLMQvexA5/jQk0wMTDgl+tiJzeNSi7dYc1t3h9DDfT
3qVFjyCaAKw7qQgvncB8yWnjsjMKcvaAwA3zrUpI9z8VWzR7nS2wM34wBsCuy45r
4x8Nfsx/Siz50jXYrm1NFXbZUx0fPyAT6+Fg3LpXdUI43HRP2ktxc7BeGH8olGXO
4xddM4MutmwMX0nn/+ESgwqQGQB0svI7HMS1l34iTheQ+smkddvdbLgM91rY0PmD
yNXxCKJRGQd/lbKABhXb3Ae3aXlrcJ5VNZcgU+QB6G1byoCQlz+I47l/3bB50ZRY
uiYu2/8BaP8ye20+eS7Hy5IMgdAOFXgI7EC/kV5I/HQFXjdLKnm8zGgEarHj15Si
rDrLJhEzagjFq9jHSbP085dg8JllCqbx62Mh3ryj2zx6O4DATsH8D0q+y9ll/uSD
rMliQa16Ajf2OvgRuWv/Hv6717mIxwevMneWrLBxVCAf9p/wnVJQ3dXd0hN0088d
D3bIN7j0u+Epo2J80y4ZLNd+mxVeTufOsUCxfCD/hrD6ewkJL0xqK7dixRmY2wt3
VV7hprDijYJjTODC9Wx2j+CqbJZ5E2fGy7ipEu3JUupPpNhSn6kWdQ1rK+NY+2pk
m8yOCRVLRWcAzXWtSEEBbF/IR/SFYu9YPd9QYpW4e2RbBI82ekNgpDBPN3Tva3FF
pmieQMFyi6ooZL5LZbtjtfXZswOzKot+c4sxkHl8XanCKEuwevUlJkdv9zw5cO53
5TNGsf1R8FhA9lzQcnKTxOGbYFu3PC0aYsk1aKfHP6WjNKvDoiL/nIuhK8YYJTP9
ziJLFzPDoPaY6gbf3Fp3kZCHKbjJy5CBCs6QqmdFnQCLrNBS5p7Mj59Df021cjZJ
Isvxqyl3EPeuLFu9agTFXPo50ROsGmwz8CCD3i6l1qNGjpGAe6dL0U1QZRtMgBTn
QVePmfwY3iu8XxXDV8cmXI82dEDVZS1aP9W1CLN0hiSfig7t5Bm9IF0XvaJ2ALNo
6iCpibmVi6noKgngfWDUd0exwkCVDrT854bjW1Wv/xOrVgyNR4Bcs4wFcivxbrty
rSfJKwlLOTXrzP5qwjPOYfw/xFbut1nsMTry7/uV/o1mr1p7iVMH+kpRLZsz4gWH
SUFjKV0bI1JoGVrf4Ok0enRqq/DQvOiXUaOzI0YPzSjlHSiyVJ4pPlX+AkN5f0cY
zEYU5/NuAiV9VhSYGsyi2bRKqkMIZPG+1dffDOCqm3DmJFX1MBx/7yaYG0jgCd9O
+UVZ7+tnfjbiD6tLHDNKPNDN0puO4clVoCusR6ranwEUzx0BtkjR6DsIqOZcXkMp
RPXczqbFYziEnxP/ydehvUshIFSSZvLoh3CXtS1llvSJdkQSejgzg1QbpyefAhVs
Er7RanQAyCdQKSNUZtpgLBlGgjm0HwPnxw922b/hpSCHCHJpkM0XIqngzH4ipAlr
NnSlyhwHvbvav0oQENIquvBgv8sRDn3SW+7J22HGALcF4cDvHiOWX1S61SlXqCNa
8nt0CzHe2jHpLAEWbp3gSv7uZh/xToA4JyIDGUv2q8U5+Qryl5MkBUWOu3s2Grra
hybzpvGCVqsTCA1hLvVxuwLE/BQJ3LeedGI9EToO0lp0KZlgqCVAIsR+gpJKXD8n
x1BY4lDH4QcO3kQZXMaEJSzvgNZt442t7qm5URUNDTCN1g1grYkb59Qllagmv6I7
iF+1aTC/T2vGAD5nzQF7IIC6a1igzmmp2Bhqug5DTKHHhKy+2U1APGcrf5D9K1Cx
aF0eZU8tXe1eMkIOoiFonBZ/RroqpslJBsRR4olgu4/evyus8eiaqAh1E2AjZDZY
ILFOJRzZ2rZFmRNUaz2UJPf9C86liRbtKm/3YqGnnAXYkox5CGWIjzVkqIwVtMi5
+cU+zB3EIaKMzzvOlUnyjNMICmjcBAChN3dbGZm4dbBHKDdZPvjUha1xB/ac4C+e
aGq8/T7P6jqFPk8vI0CKOwNISHqlYvNQL6/UK1Ox7an9zb/m3mgSiXryQoNFkPxk
Q6tUC3oRdw/P5RxyJsPvruhl9gGVw1dnzUvqy1Nso0cdm/cZRuuLnMIj1oxeuOXo
PhGwfAzn78QHtmyvwyx9dYz6c1DddNpeIyLNNz9536FaVtIjoyw7UX/w1d1uMOXz
gURzUeLKNI9AiI8Ty2dSU6QqBHj5ZdrhfxHQNdERetR07vbwhigTIz9A06O9t4dB
MiBfSDsd/EyNpg8dmfN04A8Z1XVZ/6ldfw6pM3553VSTXpi8rLXl0OuDVQ+mMYCi
rjReVdeRP0aKMo7Phkdy1hQ9ql+MC8zBAGGnmjy8FhlWV+0hdXsbjyslb9jLmDty
q31IljMJ1okHI/jWyiMnyML5VefT4LKnVWZo/sstDisULVqOWV9WAcZypElQj5MW
PrWq3EMLWSaoqkxn5xN6mlxTbRbgptLD9KQDB6jfx9Z19EDPh12o+YvjXjxQTtdH
A6RHP3qs1HkJli2NCHysDA8d+aBCeRRvY2To0fz3S0oRpQvJLo/tfb16hxPs0IL8
+gxzgKh8zizzKgyiM3eQV/v0xoM3TpaFQIZFpQrppl83it/YbO+6mkf3c6igWk0U
aAXgxtN/8ThwaGBI6U8TNl+pN+dyj8q281xzqoj9xbjYevBdZjcATaLYxksxJDju
k28xgRyeq5iZjOGAi6IzdP7Bv37qXIWFqUCVk+sxFLKvpqcnHc8LT5VPLu4TglbC
ZKgch0fQm4RnCP36s4G5Oz6fXtVqVfHg2cWep5mYrjiS0o1oNB6eiBWmlKaZn7FJ
ZVfSNuUBEJ3uLJk97ZW+yvLgcaSvZEPPLALn+jC/IQkoxs+7fP1YwKbzqy26FGuP
ICmPO/f/CHkZUjNDzx0p2OqJHA93U3UTaKQYhrwSGUl6Q+7r2M3IMcSBIjtCH5sM
jpXFA4ZCUVyWEdsONz3xkQHej+R4ULacQ2nntrU8Bp4Yq2RvnJjDpWE4P8LAfISD
dV1HhzSYELWIFLJXoL95WIHc3Ta+ivGs6KUd1AUAyZMgKhEHg7O8KuHZMcXwlMwp
mtqhSroe7iUsaIjQaWunV0WafUlslID0NlnUjQhrXT9kS306tRzXjyTSFeN5FCef
JCPyudgJQLniuUz+bdghQXj1KKCEeXoFqo73OMcWx/nQrs9U/Q0Nz7UT7kXxz/Cs
3a14l8QGxlyxmg4tzlwWy+8xl4jaC5Y0mMkHOuRIB19oCy/7i4zr5WrmrfuKYLio
ruyvkX3aO6cJ6zwh0fqQCWH0Y2PwYKru17kK5RgNmkPsj5b61cXY8RlSsxt1Q0tl
BhEINvKoRlqeJ30/Th+7KcEi4k/JhEAzxkUjammoJwdaQV/JTD3LeBaK/E2Y/Sf5
Sj1zAkXNQMvaw5C7A4MgUm5GfRuXMdftOzrx2M5Yl8bV1kEih2+n8WtHUhilarv0
ibpc08+0PWVETd2ZfPsrLyMULR9LCgcsNi3dVHEajL8I4iIomlLisa1AHVcNUzks
a61Tc74uIulmq32OFNbNyXRw2+IMThJngm+DQZy/a6wqgead3YRAVaDdC6HU8ozv
jwaqKoS/MTe5PQEbCcYx5DQ9vGYeluIR/hB3kQj3LuL0Lq4QRnAZNzvmjmBrxR4i
weFrO6aPPmyhRNP24nU2+nLBeaAO6+5SlU8GCg4natTNH/7oBJGCbMbF/VCo6KOD
q0xjD/eTWAn/IKDnt0EMbUbC9/I7/XD02pcbBoRmtBp1V5vKXOijsFXPtQGHDR1K
+kvDB6vwsMtwzf25p+ygMg0Xbc56CUPdO93+UwsWMog8ccMpxokZX+pxbIDG/qX2
vOEqFHSQ8acL/ORMLC5JVG96jOHUVNZwN8i2qpNzN1sObp2A3J20Y50UtbxjpPUO
xuQ9/ltcfzq6sNBoEFOYaqTQI73r31pjdA3iz9B2760cFEctyXYTCt/Tj7BGEF8z
oZ8EoqizXOGafElolWvugz5j/7YcTMtuHqjz5UQbxC2w9bv+cZyU17+W9YxatVkw
XUjzMOPnUOtbr4Berjd2NrE0C1TigQbBbuX9p5+r/J7nnVJp2ijAJ9vz+cRsgFsA
r969uwePqPWrTMpVyoXC9OtkDow+BNAcRH5as7+AhHHAP/JDskXLjmMJQC13ViHJ
lUER7RnlyfiJhRFpfE5FiEcrOj1FHBi8waAX6+ysG42oFnTyePmJPXD56WFTuYSs
O+NGiJzLB+n7/xe/4xEpDil8rZCVfNgyKpP8Xbwhsck5Me0Maf4+pt3YwjPnNqKi
Sv+yGQYxPlCEafUCyHiulCzVpk/Tk03fI50u08VoZ9J/kRztbL7IsUXkd/Cvgnzl
TpwzFHAw4ahG1rSs/5cHigZVkHtFT9ydN8VIlvXJDWjkloOSyZYSNedrDakacWY/
dc0k29nNSbhLF+EA1CmS8bsZYqqNzXgCGZKMDDLKt769bM9X6I2uk2fCcF6WqNox
ldKwvg5ZSToDAhT8h5ygZuxb3LWZEA9+szKYvzuHtELEHC/8UAwIY3LgHBcPWOxC
g21QYMzYm50ayUL87JhUOmIA+29VGWpx01viDUDDMbyn8icQhBDMLyQafQE6CUOc
nIK1Ttcu34H87f9563jmu6Xj5kd+9wJIFHlJUfGS+Z3vbRZ1/sewr4kXL4lrS40a
02CqIWGBdH3Ax+assI6PboTbuKVkwIVZ9zKkO7y2UyWU5jEj7gJS/P2Vnlp2RA8R
fjmmThPWv0cBntOmrsVCs+uJ15rP7eCHbsrLViWXHhQf/Np3TO7vBMIqUOtPzFe6
YF+WQGSR9N3j5KoqTTYjzqCN0y1WBSr9aZaNx13DrOcQN96mSmhjpVBHk/Rhiywz
aZuY7Zpw81N6NZDNPYshYpQ9AvA1trf4a4RbXnypdFXhj0Pi4MiXGdmJb9itlIKs
rEB/FrrtyA5XvxSn16g2CntBoryXB/lMnphlxnr3D8qDkYvilxRtZu44GMxfaYEz
k3XfBUePtI32QEgDrKBjhzsgkaXKWS9/+nqH5tt04lM3NICfN8akPj1yVdiuAhOz
7zQTUnOBawqomxvSPqDJxuXq+146NMmZUQOTP4d42yHtu43iBS5mSYbS8cp4k2WU
8Xs8YBRxgUPhM56EkWm0cOzzPyWaJxolX8AlypJbKPs72jY1ghb6nbZaAKkP7bAM
OfDcHSmrKmtXw3WH0R+cN3w657NHiwJbVf0zludsYxlCr8fVnmGQrSFcfSiLc/Xo
PrwgQCF1atN5tdDhr5nd4ol5RWYONKrWbg0DACWWpwnw24Abcg7ykzjQg0Z3cmnQ
6JCIua13/0rw/I3Pe0pDJRKu4Pqm/hNHkCk0KHZQgp+F9rvC/ddytRaw2W1uEn46
L/lJoTyHsKpiUO+v71Pe544qJCq5LqmnVkSAN5A0U6XBbGjVXm16cbyB+iWtJhWJ
TLdKds9jQpyJBz112syplp/tcn+/DLkaMB+NSIy1dZlenpRpXqjHbqXyf81wTZp0
lVLOlFaHl5wxrhtcyv6jlzpIAqqtTes2X+FIAju/11BPFwomzgthSvLLU4JgJvyq
BhEw4cY5UXTZNZRA8w+YovSY3+LmDYTi0U2jTWqI2AOj0xM/ld8JKELDdPFU3VOl
d/ISdmzJDD6yXtUhMSwQ4jKziYhEd0o0Y92qT55xYeUI81wsVAoZqTXla+PGfSPJ
SlAijuT928lyoiOT9WpdPieEyWFPzTpz35Q12M32d4S2a1M7F+5BzzeYd1V+tJH9
JqefFt7xJIibqTr30QnNcirosnxhp+pBfP64bdrkc94OiIIzcElhPrKkyQG2AGFW
IxgiLl2ajo7JLk6HIWXUinfIsgLxJqbu8oVaF78NFKOVE95Yf/h1/EDnSnOtamzA
RCfHwBInWM3aDM/37nzKvRwCyDRlDVAl4H6NGWCzu4QRdDvQOOmLt4lXtSvwCZzV
PBSX5LkumyRGCcAGY+jxANKvKHqJ65I2LrqoXglLBMetJBHXf1sMi/2WJmKrITN3
oZqbw8VgFWVvbPMRIl7FauiVo3RQmeiuWwVG5ARlIoys1nsY2NkJoHh4xe/RJWsV
tPXMpAMqL89gO/eFzb4Kp50ddJCj6+XP7DR8MO7gKUHZsp4m2fJjMpTvt/vYrFOg
DcsTma9m4Kp9DA9kddgUi57+xZPGS6GJz+sttyEQWXTaEdFUP0bzjb+Le5KwGKHO
meIZjHYbkqhZXvK097xYvAAruLXU1NVngJBbi9BKkgsDWwG/+YsBks94UqdP6JL3
1TVG1sAy34EpKu36bKf07Fl1Txv5PqjEp/JHQ3eK8pHhQBHO58AQH6ztYV8uCLpZ
tW5BfMgdMYwEHreuHjYzzrSeEX6fjKnIIoFC5ITgnTX/2kK1lQ6/DFf7cKaK1BAi
IpOWqdLKwXGZOHUYgT4l2RC/FNwE55J88Av7jkXRxNKUYuQF8mpS3Pz03Osv122O
VQ8OOsYzRuVDskwTCu+/2/6o74EgOQxTnH1CrkY4Sk4XphK2r6jHeEi+bzRhP1ZR
L/fcIeorLNU4wu2BY/oo8nnJyM/2beTOFMpI/PoNrmU9ndx9nPg99PdCbKZpk6fs
ni1mtDp8qP7RjTxO/IznxVD0JHwUo7HkAhbkWmpurpWM9yVfvieIeZQpG0DF4XxA
bi+DzrwmZW3ljsfdcTniRcIi+rjg9dVCj/SGrjx7nO/Ek1XocmIIaZJks4YsRn7C
1m8xhZBVMX/UB+kM/s7UNvh/RDZOnPNuPJJ3r2oGDKw9tXVd33uCKKQBfuLx4qQg
Vj4ClENAcUUop/iefMqdoX7hnidBScQMr0Ij+6p6p6S+29b+67KAaYM2mrTrXbym
t6a1ekTwEEdidQmXBwU3lFDKVXH8nE44Uyal5kR6t+GRgrHs6D7WwaLxPrr+Ozwz
Qexn+5rjn4AqDuh1IV/ADNzWZNnIpjvUbRktMcE1nMd+gL1hcoA4YfvDfSagQhbd
BTcBAPgKGUPxhB7We+cNLB3xXgq+rwPy9vjWX8ReMNXu1JYN7xzqkZkzVBsIFszF
G29voJoj/Lf4BcIhXw+RibtSXLheej1IEZlf6oZ+oKot8c0Wbxbn7cM3q8+mgHP2
NKUMXsQ/r+TwZhGXO+n9ezhNYz12qN701++3s8Nn/ZVtoyv3Lmuksin/W9QFZSIJ
aT9dMjXEgcFSMG0LEpF2NR88LRN5FYZgoHk1F0Ran+g+4EyLGfLn12YHIfWo/q0v
YfuP+56ItbC/K2BsBvDAiXaKph+5WKqNWafKB8BvoQpZMlE/gDapeG2rmAqpjT6d
yVZqKtFdhyZzNcZ2MUAkagm+JEfnVeNCgUd/qF9UkfbdEK1tUS0NB8IlNlc3EyyY
wbtD5CLKF92oUbQ85zGk/XIpc850LMEXM/b99g77vdPQTqHJoRdsf7ZGiKfL+YCX
xB9yGMfrWqhUzxRzJoUeVGSi4cKRExj/YETFRcoSBj3fwgyKWLbJEyKdkyvjFGUv
UqObHj7BaGUkc70mhom2qtYagp6nH+8fxd/REf/br55nG3HJq6MexUS5vQ+jMT9a
wem2XRFUJLDg2wURW+ORKQz3kpdTGFJFJCTHMyueOSgfk8WpaYyJkLc4+ysLN9XG
znQHUFxjKIA9qNicYg8BfLgBDny8uxFDEPq1lAd224lJLT8zRi4EMiGLKPXURBGg
gF6XX9FWU647FZ+1hahVaVvrfjxPhN2dzhjD530KuZkRZ5ZByboudOy067HdDQRU
RF9RS45tjdLPQUd343cJ9gw8FWOpJU4R05+ERXHMU9t/f1/HxWqUeNEm5hdj5nCA
pTOgnCOmNBKYDp3YMIaYMCI3qliEqLCSRyhkgnpYruvIT7rmNToKOIiRGNfgW+h1
YLaMsD4FUgG/Bm/ek0OCeHRSRt8o7Q0GZ3K1OhfeddfHL3pzluSJ6OZDEVY8zQcc
KMwNDZCxj8AYlHVbLli6ItaHs+w6S/IWt0j2kphHMjJmTsTDyxLFdX7LDW2nTVIO
kO8VN1zDAgW2D/KFwOHDRD1oqTW/fzSD6dSyIdg2AlyVa4nwKBVFM67TRZpYQw77
p+Vz94vgkIzRTVHkmTDyTW8UHz3zFxfY8r+y8MsWciDIRiH0vtMC4Fpae1htMkDE
gAU46aPx7OAgukHurfkPuemCEp7lyhEcbIkLIOFPCrvcwo0dKMLi6L+Jt5dWzoOv
wquBbEDozXEkVHH00eMEJowvzS/Xb8uMFdy48Nkify6ZPK98T+NA7nDbsyp7dAYG
5aFBPdVpXRCwunPHBkwbIZ1bDAJc9ZNgNZWGXo5jdR8NKELB1CACPA6OSIjvejF9
sFnTdyb56Iea/L3l6aG7SrpsfBIsf5gC4po3HW2EEvtJWbCSpoAxbBpTLVbv0ut2
L3415Q4blig+gPFqsUi+ny0Ycv4rCxMJTENjRi4C5XFfUke7F25R1EpmqjLvjYV6
EmvoKSiXVElgXkd/8AHtvApbbdpdprMUTRG2bd51fKs5OfyOJkZM0BrTWEoZm+7F
ZAHt2VeM54zdMc/3tAz5TiEhhdAAqYWHRGqwJeplCvXY/pxKij4a+grZM7/y9LxZ
i9Dgt5PZS+ld4IoeP85reWtdgWS7fYvDNUS+MgtjlJd1BwGeTNV8zHxl+jMbdPhs
pDmXom29BHqViEG6ittmNWx+i2YeVBt/dx7BksvPkrmvp+PiG5zi4OS7CWXU4vJQ
AJ0PyXF5PRUeMkrfvTMrhTn9u7dmKu+fDufBPXetqFTfR0MKS2JD4DoUe/WM1mzC
Gifb334YKJqB4m80bJT42YTtN/8iaVxbDflI1VfX7CCJyaBnS9Q0XQszI1TlSsDU
kK1q+spIoeyNPv3ff4xm1Ui4K2180mPVOYi/qWHHIaNSs1vql6siRLMzxKDBIWeO
LuojGUyaj/sIt5kIoK+Ylrm0NpwSlbuBC2sza3CsPp40+uTEN0BidQVvHZrrr4Od
3nmYTF2S5F9zVeTRJ7+bzsX2y4V3DlwtTMFiH/mlAsG8ZQpmfI6KC17kN04pG3PQ
mwHAOZ/ZjVNT61xNRDbTCAzddeUABXfOCuv09E7+wfV+TAH5xM/iKRMQWbuQ16YP
Xs9etAa5znl045nkqOQnBMmQBGfqvWkvgt++49TkVffmsbmRMRuQ/CgTN9dI1E3H
2Y4oEw4h6CufAullnw3dK5LWkAIeVEYRmN+C3DSGROcewP0vRWmH0hsP6Ruj4zKg
RiJnve9HmjRBRSmPVKj1DSTeG/inu5cDHs3p/1b2Thxug39epxua+qYccLXrpS4p
1b4frfHHHpkWbFlN8O5WnPC/b7+36dGc41MP8w7khoxBi9e00/xo1bMOTL1bmCNi
p1mEbk8+PcSV7oPgevHh/cW8yx1JYuXBbKil9KtunYBLvrRjMLoLdhnU0K8ozXgp
SYvuZmY6wtZBDpaIfbLBB12lIB0xcqPa7RdBBcimiJ2ZaEH8WawD/KMbGTbVWnHt
w3a7WfTlzVBcmOQFRN83oqU8OORBJ6/LHqhkJGtTZotacNupoRmlz8/CRPaLr5PN
4R/utKgQpqGjCnr3jluYXPOU+2yASOK2e1BbkcdB1zpup206QIpO1E5okXmzbJCc
Rw90hFFdzcc9Y5/a2XlTQpgEVCXeQGX0/knmaHRsLUmeW11Mdwd4AW8kevJFh0qA
oNYERyH54k+scWFj8cTc+6TwRq/nxD7unQyeCnlj+cJy63QOWWKvSAAwWc2q5DCv
SjvFyXsuNDnvr3BW5D1VPbaKh54E13GTFJga6clSAa3WGnsFWE0RJAaOjpmq6tYZ
wUO8WzboPXtFTVIhT9Lr5FcAgnmsF4PviN61bakm2qHNG2rHMBDo69U6LILwP/gd
9OHn7TdwaDVp75B1ZjjeQo7tiWY1BbD84JuHUyDPQ9ktyZqFekKp4sUOGLkqjOJa
uqMMtPiEMAkrc26NwjeatQ5WFhk4qRVMVLfxTDoH2SW/W7Pj/IycuYO6n4C7yAN8
1IzGGv7gkoTQokpnrRyZHRgP/f1H3bJ/h4cwnrMnlMLTFCmbxsjRImPyTN9YDifT
PBYvaKMnvxzlS9iqlPFM1by9Nx1lLN4DHF4ESmLG5ZRJ3wH3BgoBLFEgoEBw7Z+i
xm9a3rT9kTigUS4EDN+zhS9bRu1xNTXU57/BWvfkUBy/e3wurHQdVWWF0x4QOch5
OU7G2HbfbWj+RrPzkQsm6mQ8mtsnayBHLoElu6obddmgnKcJnm2GiW1fHr1lO+Pk
KPwepjbbOSmuaEXwaQlpD2cdCF7IgVAEWrB+RES4UsCwYuC79eE5IBBnShcgu075
L2S8DGaA1yCslNh0fT8sLb7+AG/4mshmc9nZzme0Tv2mBKIqtS9oJQNAJkApp8m+
pxYmqT5adWdhAxOHSGuZbwgRHg+RAyLFyqTqJ++NIispeQIxeMHD2E5iIYuVgO1m
2N4fUht9/9TzHPivFz6alGgmLdTBtxVlvk3FRsk1x3POLjnR1zLr3Rk+Tg0q+UI0
XamAvnwaLq/q39BQ6iWwK1r7DN6srKeEnFUl1EJ5MBjnGdn1MM+yT893MvLhLx1J
X9kj9p28DP33VjplFzLOVV/zT0O3i/BdQXlvekz47zzePxZXidnCauxcvOSudlQZ
mk+m+T8BNO33nf13q+YRWOpnHVpejWjqJ5z+9fGg5jj661FU+MP1oXsNAKhW4kNV
F+cPBtQMU4QScev7v5vPrNezjeTGK7dxM7oe6UkEgUkJHT2pg5+jiFqvRL42imdJ
bf7+196d6r1Gnufuw9wQcX39ncGHv+XuVR2vjKgL5HiNhJXOHe+uRpCUSvIjUlOz
zKJZ1bcS/nSl7O0EJYeS9RwYY4mxUcWqwvXAR+4WNsGAlWmH1Wc9DVZ6uK1yy0jC
2Kg6uNU4kpbb1BhAPlmLelhIVpoUP+9R+o10RnbJlnBDxJ0hUsTCZgnIsdEDwa7I
B/nAm4WtN+TwFV56dATbIGiY6Nm10GIE6FQS/pgdZJaRcsayYE2sEaIy/gWf7205
7a00Yq8989LnDt+6goP4I3syyz+J/WLTb9B5Ge0YBoX+o246N45FiU/tc94Rz7IC
Bl0rmfIP0kdu2EiygsvO8vpJHikM7uliX/XXyaYqq//6p5bGrkKsHNeuUS+SSMTN
C7Bg93J2x4zJPW41bo/7PtZMuMZN0TCkraW00KR+yd+JJqBy4J6AaJCDSzCo3tIT
/2FDSg1CAPCm8pbs+guVi+BpHZ8OJZypz5TeCEWT7+d3sj7izDtatRFBxxs9bOnh
BR7PGi+md/e1BeVPoWnfCEL/onoyYOaU9RUCRkj0mkC/6JBVeAKDxs1g/YbsVsym
AUS4vukxZMvEbgbZFUjk13DFhgbNgzABmFdauSZVXFYLR/1KGgGxKe6tc3W5v1aK
y+wZL762ilBFgKZMld0mm5nKdESE/KbJvpLr0kXxRM31ZFBarl+MQ6uPpOetZeoN
mrfK9PX5w5tIQtMD7rr9jYvVrPubo5oUD232mE0WJrK9ElRYQ4WmVRRMLwrd1MVt
YbN7lw8EVrsXDRRfhyV5GmbgcxuGDyy3HEBBzKp/hhMyGGowqTTqpQqte1cM8cSB
j+gnEXddCLOe5HxFkmvMU/Fc3D7PueNRVVKIzDPConvcT3PoINO66i3Oxs3Oprp5
lqIlIq1v7k3bPrzFM+sIDfqydflbZ5ecj4YqYMNLBZmf9p+LoB0Qx6lETsEISoKn
+5Ig4qrr2OZsOsbx3oNgP7vRKQzIYtzTR+O5yF0IQELCxWYpwUVCF37c2c2SEAy4
JHtwzB8XjLJ8pBEvxfV3bpIMMAJLyl9iE8CEq9n3YSwrHfvlIl4laUXAiOaHSGcb
WEciiSmVwLy+swQyZ+op8q7HDOQCawZVuwzhl8Ly/PC8cww1rdGskfE6iNup0TUg
bqnfX8PoohOux05M8uScs7oKsMZU4r1Jfhe7z2JSSJWZw08wlpa9thoQXLWDmRPA
3nmTRwgEh3T0g3AxLxVi0NqSaqmGTEe1Fim5/AvhvKMMmI8Gpf3bZDkFsB05gUjt
ZwTA00Gv9LcdqZ84IzixbStiYydKhJH5TsDiAtJ1kexP/OAnK+sm7kW+mtZnOk5I
zW1HCI47nuklOg2trblyeGYBtrn+6qYAa4o3/NZ7teAT3ZCWUUfGptXny6T5DiVD
loKJ9X6QZGyXEE2JmlHJRwcFb0advwMSUZTtp2az+tAEkgEQVv3CiRSRBlrPXcP6
kUqkESmZXwwkQjxWpQwFVvsFm9QVtK0SDdKg1nsAC3+ezMC6UHLjSPjmpabzZMNY
eeI1J9dA0WkdEjkV7PerETR6aYtNIiizhk3l+E6OKo4xCMp2zZtEb06emb2B6uUL
69ZmB4sPMv/aUcJyvl997UR4qop51eFeC7hzVa9FFa5FraUeQJ5aWAOoYndXB+Og
sqt8N2DndMTi8XIyFsGZDtdVxD5jSfsruKfjOJwzUF5AXkLAOjrNA8hs9JC1ipsC
CgMDnesbFU/WmBXqlp4wjS3tmidid02dbA3BG8bshlCg7EHUEYg3odkEiN2Xrjqo
FZVWfGvuBkvxTr6+O5PejzxTNDEfLbFAgPnkYK7V871v1L9GPF99BUULssPe5vqC
wctgjc27AMVkx0dhUVpFDdtMj7VGr0bZDjs2Hygqr31/LYmIHqgTkJn9js60uRcV
z5yKQSSK71RueQH1smO/wHnxhDi3hxX+CLkVnQ7W/LiqNgGvlotOR7wBkDPdG+9H
ainhex1Pr+kogWmudHffw9SD7FF7HWLxvNWZsRSkKemA1LsSlv0XD7YiS0/fGFJl
orTrxjKJgX8tBKbtlKe+mr6r6pv5WenzVgcU3Z6s0AE7dHisoI59fZiU38vViiI0
6KWMXFaCpR1luzWEUsWrxtzf4/JoktFxuUuYuBOM5D5e/ElZqsgf+Tix9ta43b5N
76dgdw8wkbHuwyYYlm2mPbe0hVTM1XSDer0MgQGNXsidBu1Mp2rj5rAGRcB6+Qs8
gUnVL310ZNtHEnuo8ad7qYpEnUQyGYWMi2YF0V3WYpoT7rfO2Cg6m+kt6ePJmUug
dBKj/YfOpPvcMDdRNAoDFnmWPdSKgRN9qSn8zr2sJXHhJu/WU1/m7gDaDeXYWTH5
tOnOdMFDWYdi3Um2E2PUWht2+CPkg3KjNnpL2MqX3wsc34liyBYfJ3PRMeaLEf1B
Amnq3d2vJ9ypbTHNRlHHzNbJT24GfTLgww5dYqdqlCxtk66oHHJ9kUFE+F5s/HRM
XSkykXYUWgYrISg6h9yej2h5cJoXLePZ9Po/BGV8mgs0nt66pdHyQpy9wadfVdXE
s39ZV3G/F+CBlL/trbdlQacF6D9pqKbhf0icOyOEe5astYk3gJUe4x0cP31/wRXe
K7DvzsEeEVEOybuz/kuob3Jb5y52VsjNJCq6NThiJru9UiT+569an5f3dFEeoC/P
w7EC0sJagpneu4Ohl/AXU0BB3di9QQOCKegE6tfz2bX5MA/BjoMuyCAkrqY9cr9Y
JQQDkCfi64wk+NCceCP9HUKsQyvINWgzJiaWe6E7fGHMPQnn2w43A+oO9UDiUwvI
h3BBogwVHkLvmpAhBjlA5soFT1CBDYOLojRcxU9NdO5UwZ1fYr15lNA772em7lPw
gx62OzXQD8Xf1aS6i9S2W2TgpiRw7O4md9GK3YnPOrQbsQabq4HrnAiK50DWnPmR
ohYEmHaJuUJGQrWwpk1LffDsb5BAsDelvu3C6/BBKpWYN89Nrvhqteib3tC3VHwU
M3GdcCbWux2Gat2tyzuHE2GGlLUBis2jZ4wKfg3LrNdzmjOPm0ezMuzva9VRfsj+
jksH0GWw82CW3t4f7Vfd23OqGtyCutcpiq3eIaWM8vMPjT17e0bU/mhHeY9oK7eX
us8ea8zCdIbHlHpwMLSgdDymE5EIUKXc/dBGbgfeONRoFaggu9cpilxqL+sPan0X
2x7+bfdkftGyixuciaXJqM5j020h7GNbFeZDKcfz2/V4s42G5VHBnr/K5T5Q+6A6
v7vBBt/MDi0Yxeceubi6jRucUFb4OMilvqvt7sccSPeEFD281/OSCLZDz0kyejLs
hd/ANFj8EU1uINBcsKIscRby9kIrN26B9VdvV/Ysw4XrPgnsrMiDwl1DT0ANFTz6
Zq9LYONC5fEUi37SJ+lyfjgVdFXlgI9AxZVcS6H6dT3cmWNmETOdUvSDDEUsvo48
XfAzERzDVOpHxenYAMzq0b9pFASbxKdzjpW7yzmlJi1jtyjMZ54pIPDVSBobIJ3E
wCTWtiRqkqKkx9ofS1TFaIF+wjyv+ib7JXnFZdQenYn1+2pyQCpDSw9sqxM0zUTG
XTaklgChHMKjoisTGM1bwk6WVfTc1R7Qu5YrXVFsEHiCoOE3wIMg7c/32vlUOQZW
CBl4xspMCC7Uk0kyESccsicyabdYpiQoKYJ/1oKMCAC9ril7zC7EfybazQSK7qrI
kdLY5It22JTSvot4JCH4AtJMr9WE2cY5cr1daEMUYkKlGPYWnVaXl4ceV2+iTdNO
XD8B/xj30vPvq9JQPRBjn/bu3+RXpcKD4yftxiByKqX9esUVwyTKf12HWGr+VNET
l1z+CZ2r8miuPQzliqvI5D10+6lM8ZZymjjYBClrrDhH9Brdx3PZRwe6cQFuXlL9
4lvsm8/JLRiYYLO9kPzza2GD121Fyd+oqIcfS8Wj0QA6e8gX7EnHaPa3nGnLQPsH
p+4H8URKAkaIh5S1dw/WP2Kl30H5RFXdOMAOSPJ6upWxiRYwzTW7PAJS8N+iqTXN
4S2YasKo75tOR+cJ2iTgIerhUlSHp/SQafBCxuKgMgx50yAII8ZFP4vTNrTcXPVN
ANnL15hLyz0Xcl3BcTpgnJTTP2hTvZzssu/pFvuLmcjSNjrQp69vJ9BpiKQJe0IO
mRoTcWossie2YTomH7BzTzqVeBzIU1itYhPzplnfKenYZjqdBPcFc3OF6Hrz0Evx
M4eH4pUfINld+IgljvrUos+BsbZ1L9AcUu63DebFMo6P8F95EbYDDFN4U1G4qB0W
BvdgRjZX7ds0UiTvYVRYGCNfZvuNHDZiZG7PBv+CKo3dFC67z8I5fcnDK/DY4T1d
k1wMLXvBt1um3X1FLziCHD0phFzGx4oieA+389VeRGYQebSQ/ngQat7J1FXrZfP5
6hkYpTbAvm1EP8K1PYGGabHKFCWavzo8MVr+sN1OBsh9YyidvYk1PGMzgJOqSjHu
Iaz/DVNMx+v3nbj3MYnvQnfTE1u7aXYf9tgyEIQnMNNDC6aS7vgMS5u0xbYQr67t
F/siRRpnP2kwhElkPLtxBMHMEMuFge//6mmMU4z6x0cIesm+cZ1G+O9T8mJh1v5S
w1uB6lb4B3QZJR56lMKZFd42CFBAJsZ8wZBH/xciReCisYN+2uJ2YSKlGtMbj8du
XY/YWiYCA0IDg+M3Ukdq0erp8o+3OWIaGEWszciYbOp22ICatA9QQ0x9WDzdrfuX
aUQ0NncNud0/8I7WkYXjJxh8laRNN2KxGabWSfzJFzlLyPAXLvB7Gff+tW2vgHyX
MUQd5RxR/KhYX6ZMqp1zE8ABlWSXqfmRS1qV05tp1954bgWbS/uxazQwE1t7LM9b
ExQtwytwmPSp0YvlFRi4Fn4+vcdSMjFyVX4v3nAUj89CV66Jv/npKlRJ9oco6Xo4
8nxd1qPjZvzae1gGL6mFOys/O6EfvvrywGkoJQ0mbFM96+pWVYNoS/FGPjaVM654
i5Y2JBS6Ez6h3P5p191zcG2gOpx5gAUG0mOEUkiUDVYJpvTJrafxy2r8f+FBa38e
+3/jbKCkhCnjJHYEvUZf6bu/oFMUKdKPeqrJZQy5aCFu0lntwnCzq2Kl31XzNesS
LmPJc2sGjuaDmdaABsPn2CY8Cp+W0ezsaz3sK/y9KXhJtz3rUWIH/zeQGeAS+kv+
qP7l2Ykebe2tlvLUspcyYHnoJ3c6yiIpEt0zB/oyW4K1pyJ0dKml71yl2fKADtVZ
7ceWDIwgv3rF6E7JpuS1rYkUkznOo/jaWBulC9rfFdj/rwM/sw88ptXS2FDGXln1
UbmNFuKf1QDr/QIlMOLh7YcqtTIvTBaEJswZ6SNSK/COU/0/52j7wKiY03AqT6Je
D4zW1qi80oX1GmGlswMLPjBetDhAeDVJ7yts5aaYLTXnfibfT+1userUbh8gRqrV
vcP3d9QXBhhWZRNOlXcRMUyqa5j9WP0ZY4IHnjMx344GoyE8VqnZsBsQ5Kh4GOkZ
8QVBQCmFJbPBVOn3MclILVEzJ1HpuVMCa3Q9iNjtuiqHP3P/rFu5EJoVWunJCUtB
64IYgSzbKh/e4g6a9H7/nBCQBskqx3zqSMfAah2rul9Wmh9H3qXTPL6H8p2l+5rA
tWGIRCe08DBcRs7e9Rrnd4HZKYlS/1S/RT0RLwHJWGRLZAA9moDLZC8l6DwMhwFB
VDOK5NSKybhIgFPnENoxp8KBvzWYYu7o8c0IfNOtZg/YJ8BSTrUjqy8kMrf/hNAh
Xz689RNY5X0HpE/Y7XzrKNY5N7orJl7CQH5cpB4BqkxFI3WnioKdiNoelI6fDoaX
XLU8q8NNzM35hyOEvIWqDUx9IRXhZKaL6ISu0+vfwso0Qajyotsj1ypJ5TuRctyg
Bh9RumSAPbjcs2xe1IlaiZxSpPS/au8iPWnYzzQB+0h+TpnBvrFePlUkHpkBfg6Q
NKidcD6XbshWLx+liM0qA0g2cXuL+Q9zODpGBSm5iboZUURsZb6z8MLYZuY2PLAS
QMXwTjJg2Uf1NducX+XwCmVEBK9GMhZazsDlCrCEJ3GtgAnPT77TGIEUTJhhVb0z
0c2j0/ltHg2Hlz3pXCNpdqGQqOwdSm/3aIAY2sbbpSZCJyG7qZ0yqdfh7vsmJMTf
ugQBRMzyBEKPsOSZ6k1pVDUKmyY/vMx6MWTD8zl9irdCeCkcJUlNaN0wNW02vErN
WeMLgRYJT/rH5vXzGxjhzLSKXE3g2NEzWtIJD8+gglT6APV4zX+OtKh/QJNFKbhn
8u3Tp/ssZDq1vWoS3kbhF0mt6S205SynC7ftqSrjygwB06Az3804LLKXaq7Vl+w+
X2/Wd2zNM9+5Ja793NpLi6DC2/S5J40tO0AgCvt0PJZy14wv459A48s97X3hCDWv
y7+xUgLnECcQFQOq0kUrHAnWLufIICalH1UMO38EzQQn/lHVURQD2agkFLTi0NDN
cwzjU3jxNmZeWPsHOD7fXeRdkOz//SUFZC9BHqd18x1WufwkzxHvOA0VeWbV7qps
hjVUitrnB5wn9OEJ9wcC2tlq1o3gohECgL1qgWisfkleNc3ImCpubyWqCJ0t1H4H
PHlWUyA+Ab1hIRxQ4pNPxZGmN2I5VK00QUi0CVv1xkTMKf4DRrNwqgGjpHVdIvYc
GHmeRIv21gsFzWp1Bgk8xYCEeBAJLGcb0Om4vYSXsRSQ5qIW3Ck0Meq9PjasVJin
ho07Zo0hd+vIcnXFW1JuUVE1me97MF0MzmXnQT/g8v1siaoyeY2kfkJnSsyo1v8F
OcUiCSpv+q2NJeaMvF+kzOxk1QrABmAA0eAaWb7Q/exWf5K0HLdB/ugd2y4bYjNc
S9mdK+FxYOrAGaZMWjqk6rZU+QhhXKMHanhznr7zZSV/Ep4obKPU3sWiA0yWDBz1
nX2keUaguUKFn1IlgNCqremJ0/h8TEa9WEBBb5kXkhnot0MAmnDlEmq/6xmycdc8
muRbG3UA+uTxxv8ULCZjqVOvjFxFQhEX7UTefh1V/PSID7UKvDYNnr4X6v/jPM+J
ElJi9Ia0IzpV3ilJGNy2rUVQ0EmJysJuzpgbAz2MpIW+bUbAa4cB/k0nnn1CT5FP
yhWNH0gRleHD7bmYA3Kq9iMwHD6aOC+8Z89L8GpjHxTqJv0/E9WMYL9mhSmJteCq
q/H0u6tDfAAyAfi72rhFgmE48Smdt5Ebwkl5JxMPlskPbPtssgpNBzOrK/yAgyg+
5fBz2Pf5ugDaG4R6JY8SN5uFrDPeX1aWW15GsOvYptajXGVMvg4K1tZadM60vtbL
UZ8pszhYeOGjb3268qPIgfbyQfzjkpZk+29iGybxfLbZ8U1SGka+hyBM0etdlxhz
bixoW27mbAmUwaDTntGiNOLORPcji+9XSLJqN+wfCY9ZB4K8A2WJq58s1aC6vkD0
oSpI83UWBtZ49daOgjGbYIv7L15nkrwPd/j5pgRNtpLsveFiQx0YuUGLTrmD+Tzf
TwgOZl7Jsv8JHUi751dFepgGZ1ucgtD/kfLpXKne60srm58y+KvVPj2X0kH8aX0J
dhKyeRUZwSdoEKttiKTRbtRdojIxLodoeqGDGKISdESabnX1r38D+WVEiu7s2EjN
72JSufyd+fEaV5htB4RCgVPGOPRgt77FljkoWXy3hcmF+tCBttGjAtSZVROhrnJ3
Ssh992eekZ5c3nEkPgcJKNoh0TjfTecj5y3AMKXJPznBGtgAU+G3+WCt8xwk4xQE
gCBC7I9bNKUbfYlZukA0D8hUw1zvOkRtLnCpbHiKQgAiNcRWCp44SKfNg/2uHENn
kFxISqU1Qjktt05ztCzgYhgT/FauQbJZ6cWvzkpjzWz2rAcwFGEU3J+4xyL6v7jO
O/sc+2Lx8YpSQpQogVvB0L/J8ao4g53zsdxg7Ga2m586yfonVwwCxRLUmraf9jHO
fWni2Eedz6v2oBu9x+Ne1LrsIuRXlMGS18hN5F6ia2BCmFtKXvGWXGhMyJn0DIGK
wltDBBGnht5khKquo4K1F8ZkZY/KAcy9QvOezvfYI7xi8Oyc640JWgUS2xzdF2qU
3S4bo/CajelA8kYImelreW4bBEt5LuSSxrz7ZMLdxUx+npDo5GoZHSpekGEw2V9Q
CVbGUF2hl9l/xTRCSr9EsIdKy/PalwoA1yQpvqyCvCHIIN37hnvNzZWdqKWhoolO
E5VIIN3g++EU7vi3+HKjJVZWAip4nLUVGvwzggQ21j2k98FeqynD6ByDt1lVHcf2
t7kQRbOAlOhsUAKoH43sGLWT7dSc7jWRONnJ555EVO5C2Gk/g839W9h7dGBNt/yR
MJ4NzFMuobX9bzMInqUi/c1SyK7pCr6Dc78njF0opYGNeVCMir2ApqhweZOh1DgX
xn6sBbtSD1H2tGJ65oLl2AL0Jd1TmdMfwBxzlbRClJfrfrq1n78EfB2YfmU4FbUG
3JSAfGvnoCdf9ipyIiggkZwSeCWgwUGtXjWYYwRiR80rlP9leoimBgXMBnuRZgZv
iEVm5gZXEK7WAIkpRsaM83ZXaCre2iEUO6T87+0VRbvLyF/P9nIs/UEKpUh2v/SB
XeD/Zy74DVVkqtuRMfrgqxW9GLKnqq8RGUMkHWmapZ9diestFwKTQT/hXpTNDXpg
GBmMoiSEVa1UlJ/CgNlVsm5Nuk+r5hyWpdr2TQ27KHWV4aW8og+0Ka67SRPRReJO
giwOAedCgMSlBK09piiXfBsDhcvXuWgcnHrOFZ5PywGxyTEhODf9M9LiIYvKXSkz
p/pv/12FWIL0aAYsD1KxmDbUf+ddosMFBhCa+3M+VjxZfP6zqiZmlrKggRS67g+q
wmDrOSXkgCmJjZaTBUB4x5TR9PEdAYNtqUzSLb5e9kofbc4etDSnre92e9/SzEah
ngq6lBb7ur2XuSkLZpUYK+JJIR9ZwH+v0Nml/LHuyu1Wfl+vHkfViRfFpyEvOoaX
Nto1n9PGqMbs0JUTAP6vDTbC6oX6YfWZszXjxKMvIMGvlVL7uc9Nih/TM14ubFHt
YMZ0c6fjxtEt9B5dUXVgfep42xa9EvhUeSxwK3HIB7BzNnyZOyo1I7GAQZP+ERxW
TMXHv2V/mR9zpdCj+uA6k471WB/T84Ensq+bmnO31pB52pgHrFTzvQNHFPM8ldJd
GTJ2cg/2KxFON4iyghw/fto5oILca0bjZssn1QuZtxncdvTba46LZL+zk+t+UWAt
UkZIW4cTR/gzDgxCJjykgcSqps+qdGbLScz7QWF0sog2l8sn7Rwwpd+y12BP2t8k
lMCh6TvkLxuU6cUI7dcC3A+0tfspwbHMf4WdXc0zQ6Pk/ufl4hseHOjNbZStOAnk
2FcwEPgw0X7eMx4MVfLga0atmmFpexypd0zOvvKRxrQuhv5/VHV0MqDlCa3pDO+O
t4GcIemvrZ8YC7EVbSsIfB8J4uArhP/C/Mgd9dRhH/GbzZ1fimEiA8JOeefY0BY+
6Sg1iV9l0WspBS8M+jPTs6l+KyAP+BETXnY6r1P/jV8a8MyAO1fHBs+hRVnldeQF
fuixBOwtRt6ulS2RCZug+xwGeNOr1t7b5mQ9BEmlZ2fhDmfaAUqYo+WQGUMlXGXu
uxpKOioQOqmta9jcKLO+v1K5bN0IkpKShONIbsLuFBrfGFpsXq3mHnlTcyu8bVN1
ZY10kQbl0Aq7BiUoEyVSTh9hQzrD1bph5tiK5Y1vXJy7XIhySWkhLPM4wiZaPfm4
azJgXxqZZb4iMpV2LfeKLXBsr24MMghWe1X/19XqTWBwPE5bQnRH3bKAtekAZjDt
1THbxid+6+DthBKIFIMTc/eNZD8SwAlThtd5ha9BfWfDXwyu5TJysn0j1OnBN9Mm
2NKEsyKkp1MQInj5Ugt1DA7QK8IGZUiIeCfKrHmWrM6yVcb3UqB2V0M82ksWbea6
pCffploE5A1rDUnadUWhsTR3CVW3rsrCVw7qAUz+0buRs2Yo+ROIvkq6jEHcq8Ue
TTjKl38q5QqEAL+XlCJirKtT7ix8w85SG8jEjswXXzM58yQfHL2ojJlcUZea9vOt
jqM/VIzw6VA3UGLlNelVK+wpqzraPHn0ykovcOMqY6vCJgJ0LpUzeQsPRE2rGg5M
DrWijlJOqkBcl//Z4CK+iV8A3VEr+0YKMWSXqsaBRfG71COdY78ExYRKnP/cYcKK
cDhldKcj5r2dH6XuakPOsv8avfGQY5X/OJlRkRoiO0cqGwBehgyCqa0xIFXU5REq
nfj79Y1kh3FW96dCi5ZN/qm0MNU+rZv4j72wI8kuVfpS1MwS5GTsJSBIysrBhiGI
AjicZh9lRJ1ePdJ5rSYrXzcIfYuHJjnhZmCZ6/dttWWD/ZkHwz/0271lACudBkaS
abOzRqez7m+Rlqw5Ctce827wn/zwOGKERZmYy1OJA94QLj23Q9zj5yTCkBlMUZl7
m0OLIWLEzrjdxcpFcjxbxVwp1Ukij0metNDaY93cmwwUGDhH3iX8Iehkpboxh9Zm
A5l9rFp8VUXqt2v8VuOSLbi39+jEPvPfW362gIkFKb42fiXZuLNGYv+Wvg0zZMPd
WVbuKzom1WtKBmEmqndjsWzULV4BC43eS4S18m2StxbE5uVL1rvDQYSm7E81KrSx
2fT1EJeR0FL6s6ByyLxGCtW7ua8Sp8EV/OkV5JEUGMdP1Ctez/B6VEsXiwOsObXe
5i3cZL0oveACnz4/PaapS2K/Ye2RXvM+aO79dfn+PnvO8WxqLVFGCZd4wqpQnjaV
13w9ZAg3C14iBRpgthXVLQjaopScUq0L3mEBUUuP4dgFQ5tFZTJ8AHDc5HK6tMnS
Npj/3poRi3wtHfjbQRAJeY4oqn5Q/wyyhQ5N9cHmPXkogSGjqMvJIXclTXzg+s58
xnSaLWTg/o55CdwXUYFuzoZUfOx/7PODuQQWMfXGPfN26tBSPsXKIQlu7g8G3l+f
9QiYKKaSsVb0GegoRXKxGhqkIZ8ONTJAyIXlh7wzVPl0TkQ+K3ID111m50v+1wuk
5ktAArcf1WJqkuYrzPYt1GgXzFLUykqHJsdTEaNLS/afIvvtf3hak4jhkrfM+1V0
y0kgXY8EG49f5EzKUPjFMRrj3rYypKZ56epnB2+uxxZXzYnGslWBksVtFg0SurkQ
kzKQk9jYJV0Wo7CPhOhLi3KLqHjg0y67lX3VTYYJ+1wSKK9IWboL3s55CVVXgjjj
/KuaRG9D25OYR2LX8m2xbo64u2OJ2c5LOE8wHs3wnnhG5HNKOztrpmjbUpyDNrlg
Jv9/DE+YpH9IQE2ZL/WGqDJCBg2lkbKeg5JbJakHQaFDhcKHDkZrWcE5TZFypQJ0
oUvNG4v0faH242+XXyJAGMMMOCwCavxUHWNCrAXBhEiza4FGLtRA6I53lK+Ihh9P
ImNxrGJgrAyqZMEl2yovAmQ1QWBLVzNiZf4Xm/EUScfaZl7GxVGZ3qEhv8LNkwJ0
qcqFUA8Iyikg+rXw3iUIur7C1ETavppLP8EIT1Jw0omOGmywlIixIXbcpMuOj2DE
f9JwGYmKwchkUyoh7dY/vpaCPS7+6hlsoTCYcnNzXs5EKlHJJ7+/UGmTw3nIrzhK
oNWlUE/vgzom3X7+AiLTCI8TWyVaaAD4Bk/o4W8XxN/Q0yP8hVvSI6mCA+Hhd0PI
l1PNky+4jzd67Ha0+M7eVdy6OVqoGeoEr+tp3lCJX3i/qnIFMiOG2+FMYpHk/uFf
HZwXRYO5JdXmHd7zJKAY8/XYE9uCLwtv3JivmRhxWIeb+hYrgLBsr6vMJzWEtg9K
9MzXBgLa2+sNwRGlEJG8Boxv677R18jQATtQ5ZcBYM1s8AUV2dUv9a3PfWSUbWcP
teWmBCV8wZEJnaHA+6IaidV+VX2MmDeD52vxtU0FQfUbYt37XByEtYQSe+urSgfj
cublIjMcPI4q6d2tyTgfhwsUOUwAtFYcTJ29Vfk7rXFO1MKlGovEEF7K+44+3jZt
1DvPytatjS18MHMAmbcHlJ2KgtKKmm3C79Zj/UWg86ynutIbVVJOwGIuNg9uID5w
RX5pHVTfmLzedGV2h6BDO0Bw76fDhuKVkLIFomnKfXOSV/wOtDmeSTYsOGCFj+lz
PfftL0lUHizTEJgzKRVqaIcs3cgBQ4RrCjilAtocX5NgCm1EASb70sxsySUheD25
0blQ24WMlkuIsjRmCkSocptSxiMFKOEOGztmpkZS6qgaFN/vS7LlmbKjKiSW1Csx
62r1fN2GrUAg7ESDW+416FUJmm3qsRmQicBm6YDQiZfiPbzy8kDzG3R0YwSOXJ4R
qSBiZBV936bBvXQKnLQJuB8Oge2tFeWJRp7Jt8tPzfMTX/EbMOInIYeuQ0tt2ITm
SQIiD19iOv+nPxnmZZkKOQRW/a8QHKeDjDVO8pj+Itg5py2Yj0a99xJcAtVW6eaM
xDfillpMmKOvj0fVh6cEhjxiHJMcm0xUid/apav5tXLqUYi6hnY14gOxaWrQ8/RT
CT80rnGdN6/mwvnJ1orGbHKBXyf6f6+cQzflm11m3YaVxG+M65vuaxL4rYaPgcjL
X34WRMShrKrK4zkmereaoF7lXkUNkHjpeNXgrJBB1bmDsIFPkQkrTbtIHHJEEv29
/uN1jWxrEz3PtpUBOGn/uTv+DxFmm6Ysk9WtsdmwqQOXyu2NdF57OyOrqlxf1DSl
cNDncyF31gbBD/z8uomrJd4BRcQqtoS1BH3aE7CELp0XQgBS8N90NWLtzyKfhlft
0cG3WL/46Ihr1kNrbQSDyLNKY4DpnaeB3A9PsuVk4sYvHkK9s5x0zidlxuR4hN4m
M7buU5gOxmbxwtJZoNErrg3pu9wjHmFRA5xWLZJ1R9MWy54R9/u+UhtLn7j7rmWu
UVj3XgQDMLb4szH4jD4UBvx1LxJwL8xvXWLzVcNDjtp7QwvUWW5TJR6OSylJiLxi
h7QorFpEy+N4F/0Gvi4Q+fpQ+p79cWlKvKRRNDpHtWWZ2uBQZhmVgoHrhX3rrNVX
0kHpuxVzHm5HZEwYvwi3VPNyYJRpKfY6Aa9H5Sf53xTegvsu/9B9MHTzFxBxaYBy
e7HzPe+75yKXlAQrGJ481r1NnUGGzgUSoHSHrBteKyltAg40YYkRimbemxow/la7
czhbADvy5wUCNorARRC2aOty9q0Bc0V0pj532syyuNp/F7kXaJbauUQOFOP3tsQm
WLNWGUkPnSa2IxlAXr3CNrkguajz59puxybbY+gDkBQog56mntMkmAkP9QDjThHu
3CrlK2h/6OgZR81XbnNjuy+EqRNmO07Us8XISAXgDRY4z8mOFHlHsTFqv3eYhW4s
H06iE2nS5omaqZcN6KQLzUuxGcEpDsSAd5vZuS1QOtd6Q7sQc4mVEitpK9kEI3tG
30rPeBkCTGUBGlnqu3APwiTpXyRN7Ikn/0bCIHhZUGAfE0LZtq9CZQvPNSA1VJj/
JRM7GakvItdWiAAGV5o7r2qgwHPfdes1ExPf+UgLbTDSfMIlbvatedW7jzEzzazO
UTg51dVEyTuCwcGcu34VMF0GHYnP4iB1ezpBLD1fzLoQtkLx5JFcRpvl2kfZFZiY
tglWTUt77Xa+fgLziXRNx/JcBEdOKkwy+Z7WiwJDeLEhSSMa3Q2qO/+U+CDKzySV
vbZrPrZcm7niECFo+qeZAeq8pcyk0b+JkWEEQAs1tYIzXTMB7OOZmFYzezRU79eF
bZ6ZEgT+L74+4h75whPg44tAUEwPJvvWPXF6zLpU04NnIVxRTNMtZNm5KMEDWVKG
SW2g0u5dcIubyYNYfVcr7W1e+lzQlpuiJE3vzQgPcgP23Fnmpwga56VsCRhfZuEp
pNCpMwSooXjxQWSSpFW3ueN6OzkQ6wn+gLI4s+CdvYGGktf7yepSQ7dhhw6ZCUkG
Ziua70zOYnQusH9X2siQBMuYMDx3vM1uIel7oXubP3PeYmagh440V5C/tyTvgY6U
BFkJ6FcX+pa07lGM2CL0hHll2i7EI+hP0+18SYY5eAmqms6Un1/hW8+FL7gav0tI
X32Nwj28Zq/VcJY2HIv9GQihD3EHerIvQ7ifEMnDEl9e1sAb8BcHOVz7pdjSwUMg
4d+WpMuy24wbtU5jVtrZ2H6Qbmxpi6HQ7ywrHPE8w/8ap85OODY9WegL7xwcUnxR
y0gmtNypdreRRzFTGj63Ein5MbMMGq5mNvRuTLs7uDwzT93p0ECtQHiPqtR0HvcK
0TtIWOiap4yKGflKC7O8lsugrnBQfdBTPh7CwqbeXqgfRZK/q2TomksKXtjuXm5R
7k4V1ZrU+g01c3nAPoIYSUuNmXo74Oxnor1jPGo2RRq7k6jrdqXPsmSqEXvF1KNV
ThKmtkvQA/Hd8VNXF/2Sz8JIDwrokNeiE6I0GL5y/2rVTlc1l2TuxkrS8evOUinJ
VKkI1O7K0siJ9y8ZvtEcgCgcpLR+QLEbjUEK377xwS6m03KwbcBsvRG9xhWVo94T
L+wOvagbGUIObiS0NX3UqLmUyk3Nyy1prhwyw1dn4gpvwC2DUZmabqFZ1K/pgkay
pukEQLErwr5uDBVtBCsRNISFuBrVJjuH4gwKZsgnlE4bEFjnLl7D+DhXkIdE18tT
xLSWR+967ka6JAKXLUyLdCFxjMal+AXJOGEue5CMzbLBfFeyUhj12BcBi/mInGB1
c/x7nzlQ6dvrwJ7lzLTUE5uW0/JNELyEZLMWisELmsZ3xAjZ2TdnmUOOlnKqdDsc
3Ak7yjvzTTcPEogHZfc+WrjtH1UD2MFRaZ8g2QD0fWDzRMG3IHyhoaCCbKIaV2FP
5HR4yukOpU7qalY+QdNoPK+EgRgcirWAxZX+Kl+ualkzN2VWUuGkHuGb/ZD3MJHn
OGjA2ZLpvAuQv3rhaeOZiJyV6q5VcgW5i3weOd0dNOlFeovr1sxGjZxDwb9GY6dT
Jyj5mv3dMAuIZRPmfadZN+ELmoSSIWnyfTEWZ8nKb1X4QEMYSiRtGyslWG+X8hDp
r1H3QdmUIzCvWqOAcBr2557NdfbMmCVg5tIp04B/Bv+S+pJJFcLToJFEyfnN8IBG
BR9pCaaIH8+2gkfWNv1E9hZKjgWNfS9y0yDycavH+g8r9qII2P1u8Zc5DumRHjCV
xTUs6NkJjvmXmjqddQGqMum/yj/0HX1Q3UhO89BJWYUr9z5Rlrs3zdyYRv5JbQxu
F0wwbhZgiyNE6gd1fuj5iw4h5nUJAZdUDLgRb/XNOxKWbYzGxSPXtmHX+WCig8I4
BdlwjxPK1cC6fJZGMN5w9Qyj67EdOyq/CiUfCzSfJA33V492GzNIvA/Ht8PuQQWH
KUAi/GEKjkImsbIA20uJl6qSpCe3PWejznq2S7jQFONHeS95qnvrFivAywEaFA9L
wDRxLdgXrkSOUp1GbZAkDB5NWhDYOTkjwX1dTcKeanszHtBcWhRniaxnaQyswvej
nZX5Ahx4pWnagpQerwnFkRHhrC1Oz6NjETIXLX7aCoQ90eOIdbATBNVEf9QoUnVM
0nKX8kf0n1fevM65mvcLbz/AP5kZgfwgUh8GlPlO10PTOZB+tVCobEBGzVqyp8hm
sqmJeCTv3HknjfdztOfw88a5sI0uWnFzVDhpvyl/7J8AuyVr63EzZtMfCN4E+rc/
1NZSM5VIKoEhbXP8Gel8cqbi9BC1G7mtwaNjce6tqwJZMIm8Qn3FvM0h+0I3ORD2
LMcjxeHcFlf2piOiv/TVDZGe5HvCDWVcw0+4ORkccW1y8jXCWi7eNtuEgWOVJX92
Zw638J7DnQp1cInFMYqDGpUldycO1lztVpMXcwlx3niVATdHUkcWPsWlLSGIdQe9
zjQXZg0U/rHh8tPM6ojltXNEAX/H7psm0K2lbXTbtqlQDZk6GGMVaL2QBATCXPeh
CMkSQKNwOscbrXR4bNjBHtzglvQIlz5OcaJQRKJZ7jqp8EaO7QTL5uZubC/6r80J
2ytFQ85s905STD+uJO7ti+2MnyPY0cMDiUg68TdY2cW/9g8c2Qdb9jeBe0mpBTk8
WYcSfN2G2kRalz0N1UOAjmOm/oaQ7OujOA6qW6vxt7g47myJdbQgCwewQNyA/fu+
FmBGCIR+oeWDlWXHMK3pO450uEpnPFBcoER+yRA8a14ogQVhKhl/mHw13Z2Ezka2
Zo1qsfzMW4drXtNNh5GxoGkFmk+JdpHuD25TYlG2a0JQg/pN03yKZlPWwBWMtdBp
MIiyjMsAJAjWrXlB4OZ6PETEnsCYGSbNu2ESe8Z5LaUjm/NTqFhqOh49mY/F97oV
jZUTjHmdzvIOuAfwaLKwjH1vXSqtXGukyDzO8NyTuVhhQw4LkEzhE6b4XTZCgVfj
nb5HHa3kyf/Exa8KxMXcjRZs1qEZQzaGMDTg0s76ArWPW8Uz32Hxu4IHKuRDAwrG
1XntC2Tmv5P4ZTHb86hQp5IKcFvIO7uUUFpzVVLevXqPOU/waqv4CCVtAeS6kqFZ
8UX/QHHTBRLoCiX1k4Y2bJFpqKb5L7b8CEI+ec3nw+X4yVUatmOLWBarEAa2E7td
AtpG6bkyK/aHlw0VnB6neTWq/kfaIP4rkMHkrogvS/KevfrK5zW8LJUMPgbW3I+D
XZR2/5MTXm2fTcA7cY4sREjV1fkDQGZG7caHdS/za17iVGdL9nhShIWwFL0KwpJ3
Dgm7+X7f0ZVHQBhc07GG5/amolCVjn3HfJP3nhiHi1WIAlokC98xILFHcgIPiJak
SOp9dmR6eqN6NYZ95N8flUDIx64DswrdVZrCoCr1mr2K0Zvf1i3WkV0MSO2E0fNm
Skds1g+MuJ0u4xVOP28Ag1XNhqvOr1OZb0rzt1WJ0Z7r4XDgGaYB75jRw29LcQt7
5TMBfdKhTjLKffAR/wOs+O0ke/HaGOrvbAQJ/APt1kqflGToE0kh54ojbE3tne+A
MXeALIAwmPHzH8NcE6HTpWWmtUyHa+vHylhOTCb1qA50yug23USdFnPNg9rWC9IZ
UOovCo7lTO4k9PqbbkGgUAirtbBJmyF/qgijytHcb72wWlBRbl2Y4utHgX30uUwt
aCFPBEXdRQId1NumE2bMDUcqyzM8xoTOcuL5+4HFxfepUJvFGzb3xU/4Xc4o+U3G
ZEPUbr1QJFp8SBArtUss8njFYNv0/hnLtdbhqLlIx/mSlcunI562/3jMO7Advrgl
4xotXcI/R7j4KT3sakuEKmfNYBnUkuEQIzt2+Tt+qXZnSj/y+UFppO+CAKOLzDXG
tGDfP1qlepd7cYiPJ/JDON4aLN8rekWjljCB52y54mija32SEmrg007tanF6LTtK
Ss+m5mlRs6QWe3TkOo9JyMvxoMRBBEonN1mlMyZ6OeTkgFUhnCpsYyJr6NT/3Ky0
gW+tdoYejw6IOi8wgHmLCqokTPPihkhYL2DvRdYHX1XII1B9awkTBFaXr3smwH5H
o1HfUT62W3MMm5lCenvPNrWJAO186sdl/UVnoRu9S4Ins7ZL7NoTobQnyfhKq6vB
xWFZ16HEN2fko3ACVdX1t5Z1t0YlYBQPjd3Sce2GBYwAm/HaiYHGOglMvBU+07Rr
r76J71gElNnnkJT3fzK0JvV1JeT5g5vxytRCIIpbjVbf3e5gAm3ffrUFyKKBkEcc
oaj1PhghYOua0aKL3eB6EN+9+XrWJ2GOu8tb1Dq1UXbXxjVQX/qTxL9a4jY6JY38
y8aEi+U5Bq7b5guCNhRTpH2kNQr4G+MDv41mqvdqCe/UYrUHr9usMeOOiwRxsv//
nxAANCTQsaXZvbIkS4cW/Ws7Yltkg5aua694X/OPWF5rNuQA4/48PBIXf7mznzpV
V5yfyX6ocBq2HIu+Qm9Tp2ayyRgAiIAAQxcw4NOhD68rz36kL04Tt7nl+N/rF2mi
Uqn8oEfAyFKr8I5yia0b1p+gCiDFA/5FbFs51StipZCl12wUJ2ZLXlZPqFsJGQuw
KRdAvoJOLtcW3bBZrhobPsLcnCOZPpBPGVh2oeCOeorLPrb8iamRUKoHIcENCjrm
9sTpKa3OKCDWFEIROFHuyghmMffsJjiLQcPs3ZE/6eaKB4zZ/X3WAMsX/dWHUYDm
Xd+7GFkC+8et0fdcwkq3dzljwKL2oS6gzL86jYYVp/1DhJyzE6QH07CnUSz2YF1a
9LIeSeWaOQ4j3l5tkp+UDZFXUsh8f3K6CGvlO1UM3PGUV2WRoh1oJ9FhKBV5pG1a
JO1p/cUFu0wWgcKwmVd5Sey5DFvNIDMzS6ShiBen1EZSmcc0NWHXL8I0Ea4oKHD9
HFNb/vWmEeIcxYxIbN1p473qNqMJ29dPYxlyEgkD715MG/swiAjh8uqD6yy9mOLG
Cnji4uUchWUMh0l6fZNo/xitBjRe/RajKiLCFBuIUWnwfV/eu+5H3X6p4RaYs2iJ
94rqV3+7WqxiVuz5EzE2OlqBrbwNQ71AvnVDsGfm2LQp76Pg9WdFNdXi4Li7ioLW
7gossCx4O+V6x9LYS7YU1aQi+MigQGoEgGzs4ztu5CHzfktFLEt7Pzi0asBhZiPz
IAy5MmqCm8D3qSwCrgHyG3jxb73s4GxpkVX8y9HEweFDgOX0+TIC/vcJH6qhDipn
7vdMyd2JARQM7D/UoycMP+XFwF8O+ciZwYZbBuV8RhoEnLzum2h9/plLxs1Ggm04
dEwi9C+2Z+25qPyte8TNDRYYI1eRbUJMjY5U+nJYXKwMm+UXuVdifFOriAZB/ysz
ie2arSglxHZ66YdTWo2+R2LKf78zS3w0F2bo9/PK5iEn0thiNhmIuAKQ4Pr8X9jm
bXC1NWwvcRJdrIuNz5gqxrHbCYBlNUPnkrXGMY8iNPP5aDtZrr9GL9P/6abFYAn4
/KCyLw6O1TL9fqtO+39GeIdSk9cLJqVzbI38xjwYdr86tP9r6KF0s5BzO4xDNyLh
bWgR21yBY3Uu67k36E1SXzRLTwOoaOhD5Nss/mU56BCSyBKOyq/L+v4uRkLaAf7u
MdMLCAWUCG6zXm+YGtFQ9rF7cVs3F+N+xuHDfEdymCQE41YqbTnCLQI8wErTBZef
CM96lefUXBnxdGvPVUnMUxLWp7x6S/mOh7d9GYss1sR4YnriBi9tfzzY/kYJEade
Ju2KnVm94rlMoTmY2rgjUfNwHDjIhkx3fucEl8fgkfFQQYMzty9mfZkQHdev6RsT
pY2oT91TGsHlJbuo1W446qkBO/Wa3S8jctgeHP2M19NKbi41aleWtfEL1x9WUcBe
r8s3nEIOaRSneQFt/yqRYG4fBHDBh04J8VyUWMkDo8zqv2hssV0aXsxoiBTwVAnW
z4x7rxJ5OZguExolo/AKC8bfqYD1R6JonejYbbXUtuNjh8/PKih7RXSWFNNNssLm
HzyDA6Jx3bDxb3qjPUbnUHp8TnIwhThIz1p63TzeDWGU0Hi+RdfF+m0RtGRcW2zO
naVnCwqYr564s5VeY+hl8cpsl8CHBKqes2B+e3+jYsErMNziSDATArki2jnC983g
raoFwtxj0ntA4rP3v03CQmmqfjxhmcz+u8EEekMUbw6s+TREJWu5WDxZO2JcKGsA
3+jFjlxZ2Y0BwfZy4FlQo/MSCPipA+R7P8m5pAUUiSyT2JgMIih7qnOZbJmm2Cgq
EcL3byfpruccTPq0CCPupTWdX0jzSZUNtHaPnq4hK/rDzCPPDFmhcpROwmOWvbq0
Y6VlbhWiToMXIvehv1acxgsk89p/4gqT4NfeNMU7i/kXV/2YdB2h98YKHlpStUR/
6xDFPS63TW18IvF4B6d0iD9ebj4mgAHIenAD1tdmDl5GZ3ZSGKiwKoF8J4gpbeEx
C0IJcrLimYb3SfKU/Wny++Kndw99ODuTQJ3VVJdcgtCU8PpIPjDEsg5TON6FngoF
C9lmnKYgbiDAud4gnFHs5YYFNQz4rzhpq4IgWNd1IaksFnncvDrzi6KdoTd8KLSz
vcABdITRMr4knP5O2VuW0l8sXToLrO2w/ValDjXIdERHYNdhChoPaow4pFeTP7wt
bmccVO8yIld8cegN8ik82/mfD+0FiMjUXCRiLuNHmAUGa1twzJPi7KpZA0mHd/nC
nyTbKl+IOHVnZIyTWHH3gRvaJRhoNAW4FLTX5VoYj4TkF+qgKbO2RcwucwtgWew/
y8sHLAZiwHGQ+ZDg88oQbBL+O1qP6FaWIGFYDNTrzCbHkrqS+ISe2xVBp+MkUlOa
SE+zscUAFXz5371I7Sf6x+VcqaArR3k9owqswDUHetmdvGWYbLLf1flkRjba9UXC
twnthOfIlkF1fp3vRZ0atbLiYOJ8xvDJBsL2JFwjCES/93AV18XMsRN/3ZrcVNZG
cAMAxYm4DY9sG6EQQ61VafD/rgglBhEXmbyZgXz1fgCjC4UNjBVco1VrXOnuzggB
SHIW/s9SdijeuL4N6KJihbXJayLF9c03j+vDgR2ocVunVIVuH4hYiaqNRjVcYclo
n3hGMvz8k30n1e3GipAnbWKDJc4VPWnDE2mbIcO4RSWqGIP6w3g5N6qnoCwFYqtr
sco/VyfCZhnOrfIdrrP1Hk2z9CVZK0S1Jre1Io9g/nHI3mqbIUaABTqM/nXeOjiB
behHxht8yLOsj7AGP0rFgSG+eIB4Ahpcn02t8ijYXNgFlHnFCISWhFQ11xFt9R8X
uJIpAYcxL42+5a/xOR5vHgcCsjMIgL+2kBD0nDSibLL9TUX+25TJy+y7iGmaRhCY
2sODZDTnMrbrvgHX5JUWo1EospdiltMPcd6SOoulM5/zllweD4N/N1w+9N0HRI61
V2IxgCJb1o1mPQyda3MdQbF/TBe9/eVlEu9JOXUA2vIbbtU+Bs5Bm/47dLD1LQQ8
5w4FRoD/2HHyn0tR7ktDiVHnSJHFOPIQrwZZzqham9R688Q8eqGgJOgNCKGaR+FF
MGYoY8b8zyCQKEeCkLI8MWm1FcJd5B92gAa5t1sQoz+7/AsFN6eDtiDfulXuogmL
bhKbgA+LRWCxCe3YNZYY9mkerkxc4vgrD9qgL+VLQrMtaKgvFJuvwL0ViihZXvv5
IlaSrBsPHlB74IONCln5Ee2fRR8yULHGknwEIU1bHJHjdHRquLBnlXnBh95xtKxg
MN1BnZGfN6ObIVkBFmAwsaP1fodSRlMyJKvf8dY6sqMQ+svUyFI6BftIcJ4V9rmB
cOlgKW4uUTOM9pLKCVC16QjJ95YATNqOSmeRdGCVw90pFmxnbt2s+7XmsZzU4oDa
Kywh8vke/pwpMv9o00qO2Em5XFUa49X4abpsM6AXJpq3gB0uK3/ELodsmFqF+gQ1
J3wVIHHbkCIYRHfc8w4y5pRzWnEZAw2j/azI0tHjLMRcF8SUNXrSel8Ld9sJpXTi
RlAkZkO34zfpPh6/KFk0yrImeM5oq6OUHgr8MCtI5CGTaraUkDYgoR3PJwSnUd/l
7Pz8ai61qlNXToERlCkC3fEPQFYFA5N49E868aZJbY4p53R+WCvyGe3zYjtjgR5w
Fm1Tw7JJD1gGep3WIrDIEL2NI7ZiGIIemUy2mbkD2+A4Gm+5jjZ0iqCEdKJk9FH9
69MZFSYztmBULmUWJp1rbZKFFqNEDVYGKHT43TKBv+M87pSVFc1fK1RVydw6KgIl
884E+C/k86/lrEcqdhEA1ezTiebpaxXPXzF4AEFzayPE4PzggjNYQneoJJeK5z0N
4uSm9yrXIoj40E+wa/mWIoASiCdHCz8wm5bcf7OyZ260GY0FO03wak33NMQSeyrb
RFIEU/gpceA2QHrPwW7pmjPyojyNAuwzCZO7hENhJRkCybOYx5nlAArq0FKI2n3F
dZOU3QkSwTAqCsk320m2ZlOnyXPSLmc0XKoYTR9YuVZeKUrnwzQQmG5CrZ4+t90r
Y4H8qgX16AarJQ0y1zJbr6QeCSwYUtg7jVNa9uDrMXqSv8YjNiOuVdEjxB14EmH/
le0soa86RwJOGxn28GN7KfvZl/ZA7O0jWoCcW3BR4W7j25lfQpoa+gRhkAxC2Ms1
R2oLj0YRcSGOC1CtxzS7OCyree9QEVJZ6ZIxDLbMHGK7uFJ1xqPDeSWaq3V0PLxW
HmZ34+dnPjYQLFGyfRk7PvI1VGzZ6t0YxdAP7+CznldQ0651pU0mG3npdMmEIh5f
iSKzeUQhne+RR7lZQha2xWrHg18T/pHLAhjUJls+5pf95YNz0CreRaXFUiHLeDVa
gZN0L/R2bWruk4k4JDEnoKczH8BTCcTYcQzqw3hUi17Wu8tNsN93byi12G4+ZwHA
zgOvqDTHgDY9Wr0kUHiBSx2wZT7acgOhSWU5p3HoIgIwJr/tkKXgu8Afp92OFK9m
FiDSoXtNk4YRM0WmQDpr1ndjfGXA0b/Ynoqmu7/vyRc75xSR+wH/2EELWxyjR2lc
boIb2TWKm5WbExvnvyTULbPn3sCH6I207mAeW4jtZxIhFZQGgvx4C7EKp70YhnJm
wHf2ui3u7E7GEirEnZMEJkLGTSls7fjWgagVTFcKV3TlHWoKRszTiBXduKL8Ao7X
+PM1cWZgAoLIkJgFbY8GcwyR/pwb4CBI+U5esnC5w6pjYPzYUSike6IjFyfWjCcH
WB6ngSgw2EovODJzQqHEck3wdpbaFSjoUdEKGZydz6r4dpr41GsLhfT72ey2AbiM
29InWMy5ubQHcFBQGm4uHg7cXxgxdA5ptU3eyPCxba4jD1U6t27wZbU9XBDs8mpp
rHdnHwXMFaDIGBBnV0F6U07ijQgm/UsKTTan0FefI2Z2JWjQ0dAFgNh0leJM3FUW
E5l7jQ2MhPRj6a9wrZXOYz0T8xbKVLAjan20a/7vZkgFzUYIyBvw2jYRsrVYs4Od
Y1s69XmgPzHmPV8BHEOvPQ3jn/g3Nr807cjofp5KuTUR8lw8fi7lN/8euzpbgSXO
2wZpdEUB2PWVne56xbvwTAHYKpWDZ/1p4UKGMOSvDjuHUgGE8ouG6PRb7eH+y7zM
CNtbuqqFTyqTOmiO6jmuaO4Crc9QPubkSEWBrEM5YFEM52ea0Yeu/jYXLjmW084D
GM37TroVD0TDWLi0ae9Q382L+ShNxjqlpD/3x8mKB0Ey0tjJI9BWLDquRa+kuEgX
pU8725cHtdkfwxq3f+ZH5gwamCHi7vDWKCATvyEMtHf3ft1iECma5iUIywzcNPlv
M6EdfFY9uxKcOup+z5aKNR1fD2GAz4PxFqosWgEWxLNqcJOyd2Ebcl6GKFesntH2
Qmw6n0MjRi1agsecqdVNxGpFBWUW+xsSuePT9vyGpJhYEeBKPQWFY7eShUHqODFD
QXzKW9STEJddzR/3UaHEdMJFcp+77zLUYdL1UrCehf7TugxQwYdnThhoW891GND+
MBaLJrdWTldO9+8HzuI7sGSWly5EyFM0l4V7hkaT7jVO7DDbUw13Jrk3zhehte5/
MpXJmLvX/TLsmGHcS2u9QihzGQddcao/eJN93/bUasanqGYZNGHoGLmkKjhDPAXH
HYukGDEu+slrIVxrog4Iyw+guO01NB3de6cqH7NYtQ1qgmEKGIwU2BEpRr7O48/h
oZuCHeveF7JfyT12HyMEGFpTjJ/o8w7l+QrnIYrKScOtTyozSaRqUeZniEWVwIt2
8UOh1K1YC5Jk9UscOzpB959HiZAPvPPJHVUJzqkPAaQnXfuyNFgz/4FdSlU5nc27
vd85lTBG7o4solvt9v/MS8O0cMJaFNhf8r5m/XdTJ4WVWH2ot0mzHM7yGxOu0QH2
2koqP3HpEirApU9U3UmS7foFEEIioHFsDc5Y4M10CVVqirAx1zLwReW9gL7HGnWg
83Y2uJdXmDuX/xVokUt1CwvoXyj3CPGnut582FeUqwmVtZQoV7tHoaRskbjDv2+o
q5pOY+0hfZmKo4SWgqvPOkP4jxqXjD9ypPShZe3JXQih1KHfUa2oeLb/dw4sWPc+
3VqVpNqgSJLLjxAG1epTEyk+Z2TYCts2R9D5w3a7lzJU8BkGL/l8+No/gWPaTmIs
xsY0016ZmY03Hqnsk0m3rVZYQnVGxdps+HsMA5jP1fvnVz32Oz3W2sNxrAVP3oy/
O3ZvOAmLsWN4JudJ0jOk6MwEN3K3jDM4ERDRf+D7ul0S6V8NOHrfj/u3gMK5BZXn
OlvoGeFSb/to0b6C7XZIgt8Q7YDFDSi0G7s5Yvneg50C3UlLXycbF75LrYrrvkyo
ijKzAve/6c+rZjTwLX+sK7isUDq/wsBJcPg+JCxZY93ggD4LQHCLWlcoyEEj/A+R
nmVIJ/Z+dGXtwNogaWBWPPa1F2956YsKq00qoLz5HM31H7tD7ElFDjV/IPsCqvfl
WrFwoVx7lKKf5lFFrYbYci7nmckkQeOVBSpnOE+1r+79E3rGl7YD7HBPLrnvXhiY
fKa7DGAV3MaJ7a7ExdgJYYzf+svZ/UweiiRyUMZxRo3jh0upEnoVSf1UECP6xD6o
rdi8jzKQiNn3OfvyILp9nM5Shs1e+rHbd/k/up2qprNPdhIGdOMI+5RyvZZCjnDA
n2PHcdaIjhrA36oO9YFZoFWpJ1DvjSGkWJglw8Ho5czipFzo11cuNTa0OHHvrpD4
2rWGqQmNyqah/ZuSOteH0l3yeG4vuz6tsWRraFtcg2X0DufjLxUmQb+SDqrCJNs2
+0AdMsBCxKh4cSf3eqZt7vYyndUQ915Nb87eMAAwrJUlOENdLCmQQZoY+kBShpkP
LEqOVhDau4lZ3Z30DVatxxwEr4ifz4hqDvZ+S1O9xG+s2SVLYblkLvoQ8/1g8Hr/
CBoyJdHR+iuuh1f/G0PIxJ2tWcS/d87XZdLXHWAJNCfv3/nRDyRM3rT3oIextUW3
adRE5YsWa2rhky2oCAvGolOH+uDei2YPnqjVN9UhxgMe6YelO+JP70p/he93lmzx
Z3QnrDJBGFT7ohWQBnQ8HZV7ggDhmsfM2/3mr63MYyZ6LdiRam4TxaGQY8e0jT5Q
dndhNpkI3vkiC1/hmdwAX9PaSV18tJq6Oitj5nSLPxOCOviJckLWsXt4Lm69OYAX
vAx411em3TxT+b7Z9UIrp6Y0SbfRe7NS3Gr+qUjhu3+mtCADzp4T6uGXu4v5HaIE
Q6humxtp+23dwomgmd2CCrbcDFoD+aaHGHcg8yjbg3ooczeklmgTckWXePxde2tV
6ALUZMqDFUm5Gh1KfbnXWrjzJOfp31TlOWXfAD6CG7FgqHJOJINL0gP5iVBJ/H58
m9yt0VQm9UYy3iHhRLrIsXkdEUZJZy0lMhWaUW8raYQdYCrcwoXazIIXDgdO+r6V
fuPD+5Owx1X6BiMoVz9uY2Pym1X5WAEYBbde6SSUmISu77ZXwaEuWICGzAExWzRI
lD1EmJgKOludCEnUZMWgNXp75xgRlLnGxYabbqpcM4h0pLDslOHdd7nwQGQ7mCuf
aRZAdyyLoKd8UCHpt4SkXrIbPEqxUWRedyONq03EYK1WWaWqyssPVJ9bRr972WV9
bckkomZiOJHC7vAUgosVTh8/wjXLoFzQY7ediGNXdwwqjc9M8uJAl8ZBwEFK361s
1iFmM4a84ofRRaLVagN56moAOm05GvK9xLPVUrXYgTA6B56mnxP3ogdaDazjraLb
o/VPnsFAwhTKe8fmBe0X6ciEAvOalgXU2HwY3qo/gp+/CINzB4KXLGfnhAx4OtEn
FlJA6/yMpmYLNXeFWdgcCM1lb9X6Qx56aBip3uPEr7OytrITu1VM6sNIyQO6hlFE
D9IamDajdLjLFdHlbtYTP0WCKJsYYy3OxV0smF0QIgEhJMi4ia1Og3BKq/tLOLyA
wO+zts56Rd8n2oNWUrsVBK3iiRYPooaJIzl7hsYLEScj+v0LfUoXhMW3+T7jzmL5
GMGFYmSYz+jvYWlznK9+CsDymk1V1cTQ4eT0nwIRUPxxYYicNd2N3T5X8sOVKlBl
EiP+ELSqAyKi+Kz6Q98jOCFcHRSI1iAGw6XcR4qGxHr3LjIHdCRPCNdMTwu8rlh2
n5cW2DLbtS5XXOIgcLbe1fd7rQh8AJWaN241fF3ctKrh92MKu8Unk2EtL1K+Jmji
46paNixG2odiRiRlFXzzWkQ6DIn9dpmSiuQU46ZZeT07GBVEyE6rkUYUIDX4F3Sw
LrRA00M/TN2T7SVfkN/eMLuvnOzW+S3s4JmKZf2gdTqdQrfsrjdYXQp2+5qnzTvW
K1ZN2t2fVZgSCwWOChdNn7r8JXKXqn8l8x57JgXugUBZwSE2EeZvW9iqPlQ++DWt
Z0ZGac1TFldC15nDVLf31IS+/6eamHxYlgwwfEwR5DbcH74kqwqU3qEUyIxGrF4g
uFXFuvOms84EBl9AwvYWBF5Jd5B9LamL7kDFyutslADapu2JcmE2aJLD1mprXqkR
hwwrMTv82pyDYAN80Ib2Yz5FANHZFx7mO/oRr5Jg/jSA/DBAIyJgfSCT4wVdMITx
GUYZUPZrFk/4akb6i3cmZY3IBc48WFb7j3dtb8S1WiO9okgTdbSgq57BodX1s2Uo
UjRT2PNK1pe+oe3rhpR9jGeJvLWty3b14ZdCNlKlwYeZbhvu8VuH6JyffTrR2w7g
FSPHnC+Y74Dw5JaR3VfepveSuq+FwPg0KbfhNWPLMBeyo2OwKwvDgISMFMmQ0j61
bJ1QLg71tmG1xnfNKJT3fLEcNZlSPwMFc3TdH6SGEvDlt71yEubEKV+3WQ9EQW1K
ratl/ejOaZ+dUNtwAdJ+3P5GZ1XIWKcFGTw6Ky/ev2A9u+I0/hJtUJD0FHf/lvTH
GZcDOb4C4vuySsidExtJzT86Wzv9QzVXI3vEFJ/jxF3JXu4WInShNZshk3M+kKl8
dQp1sfRlghOJZA3o8kkL1dsUVPX3/1FrdxiUVrsSuusXds7jioYxEiW4r0Wo5jbJ
zQYstyIHci32kVtXWqBCZhIkjqeKIRKF7+RNgctMekPlGHllH4ykpvJNDqWEQ/6r
/ZW+2ZmEPhlVDkeiN9zOZW+zHUH35GBNYlw/NkEKYjNOa74yKGmukTnBiDPoC8yt
K7i6QQQ23V1XX7rkdgnaM0JmAeZohUE6eIREObVq1qkdQpbMZ0FhmpnoX6s+8heu
e9S7p4Nbl3p+e4kcvBSJEXBDWgdUeSW3uFr7bqKTEuTeUgb3TDQF3LUlUVeLTBu6
e3AY/32ViDJu5wkEuS5BDvEKNYJf5wdKEcqL4Q+0lWD9nfmA+/t3054ue3IcnQEW
+1fg7HJPvYfCK1jE9yOjeg0myXBfhiQqkQCaIjbl89uKNocKE+qwHWQeHLzWDgMb
uHZByblVZaeXNNEckVh6vmoXkvQKcVpDjtZO9EUQQnamiqlLLUkkaFv+yya9HxZq
Pfrik0w0yJ0F38GEnCcAnxEP8fRPFV17i1oT/3omxetgm1YNmLJUypT47e3JDeUk
I+idXibe3gT1JQoiJbPKVuyophF83YeXegdghvh+ONuJdlSxSEwTavMemAo4qYkG
/BsMPFrVr5NMAwQrbhNdnZDg9+uzP/i7OLs6pZVloIF7rAj3WLYBecCRanU2mo6s
HncFa35PWlZSQX14CQjqNp9HjUGAWLEIMZNoOE63K6U13EKkHVQ14CcIoKSfKhIM
T9hc4e4fFxFX676Ikr9NekRDsZDNdNFFT+CPRUZ9BFofBUBtPgHGEZDmELsBbVTj
+HMP2S4s9zaFId5P61cch+qJLe1LV104WXMYIYgyKXnm4KyZQmL8BMA6y6QQ5ewF
bT6ZKglkpMUEhjJ4dY52swMH/DvWBPm4ungQyPx9NkDucnlytYSBZeP4vOW8qL8H
4osaG9tPOg0Lxxjh9JxlQjwqhAnw5gCNGPhEp1hAv9mo5vSPyeb7PEZ7hj0OQLWc
FgNkAV/ZprLKPTDph3wEEZ91UZNE4y2xI8D0bgzdwrYpS5vZ0NGMecXMMLfwTX4p
o9z/wPXUO0X/LvOhYA0YSUsZMRCUOlMEzK9Ec3uRmtbQCQ60U6FviSMwf61ya2Vw
1/9pn0RVPWAfSO+BDMiShHyBlsiPpfOOHTAoB0wd3rFIJK9r7bSeRcbIA350rlyK
DucWBneYmkO/YIgkGiMbbCVY6hIbMwJMpbQ38fBU/lqYIdPMa5YodNQvS85kP+6B
vR201MmJaK96L4GMHMTFHVMCNc6571w+VqeQDAhJGMUC0PZ3XTSwPqtnXidXL8+F
d8jMMky0C6n+x4P0DgNfQY3r/A3p95Syw3kEASCswu8Uh5ibDYNPeTGzzdgGOW3q
TvB4ZjqkB+TfO5zKULeLbAtWAhIaJJlzSt6mlcNzXv9575vMDFMRcip4cgtYHJpG
hE/Pa19lPAwEyHsAUZYyW+f8VsTFxxWmY+1tyzeWeURLSgrIoV8FtczuSAMCzyui
UzBl4V0ALAsvFviRzTqzqQ2X2DM4h686Pll5UpSAWUhl7Eu0RtJhCWKEr9MJpQT4
GOGbUTOvO4UwSlWtwpRhTwqT1jBERe4GtjJQa6soRVDCzbsm3QimS7HrsFdBX5Hg
2VG6el/Sg7MKx6tGC2SRXE6c906FIRSykzZJcJHAApYYGqi//VR/ZaX+3tMOxuUE
2+9wv3w+DBYLM2wAlNYQLUSWAMYSCJrwL2O/kkFHoGOJBRTMKm0ezDVdyY349t4U
8qLDY2/rTn7jflM+BRzRER9jsuvACyaaO5U3dvptUVmqaRpLT2TUEo6xy03/jE0r
AvQ4ggzh61OiOr89l4wAAE9zzzxmHY/Eg8thTBxpcV2PILc8uXdH9bSS3M3RErnT
WkEyqHx0ZVb2zd5ncLgpGGjhx81gqSR0Jgot5LuxZkZEthCo54prsvSPGLh3RZTG
kLsDKEyWbWE7CvOFL07v70tKSgYvpa2p8zezB6XZUQQklx2tpyDB2BahjPJLUlJw
lGqo1OMXxFuNRAPVXTnXM8RxXz4ho4IINDRIjaGmi5FheDjlrRD/s2SIprHTWBg6
o3O76B9DACRabqW3b6DUXCRYQSa693+WQXYNS5SvsvwuMazV0rP2+EW1ykwEp+5I
jydKqFd6i+GbtVQI39mxgvVAvTbx78/BQfU2oQ8fE/Nvm+qCUuWSSsqb3IDeRKce
T1YTq9FGFapZrMM6Xo6Invjo+Gl4X9f1UO25daDr4jNdNBZowmGhMKOtnq90W8cc
y+q+NBGUNKaQxdw42oUiBQv60PaMbeo3NeAr4lq8v5kaFnac6XEureqmUHyii6nB
8jgYC/n+GfH5vBCOY2z0E8AtcdfOQa6rbcztaz4sDJscYST8WH6c1y04ktPKYijO
c7wbI4+JhF5UMzPlRGCqUgInskhV6QXpMe8KxSp1aD2OSQb7rXGtehmsJwzo/7Q4
/5S7Jqwlap3QZ0ulo+hm3RTRDHpP9NENuM6DE3tW/iu4yFtDOoOQssr1nZcnMiZo
gho5BBcaLFUiEdKa1NBpqjOS4i4AVGT9HNcJ/ebaMtjwEiivCrJrSI2VnD3nCJsj
rcUFv04w7mAq2lEDzgNZuxQ/LV4Wzj6mPZA8ceRQ0+gHbfoLSma2vANM5fFaA/yL
/eIc/I6KWKMA+R0HS6vmHQRaS0UPed5JRXu2+vt7FD2AcwSYN9N7W8pdpKwR8EK7
7o7q3ol0fN9SzlKRK5gLtHe90JQ1k7Bao5qjajQXZ5BRoAfWPbVV5OwPXSAgD1jv
mmJQ6Hoq83NnbzStyWSeSMvEFzjP7oKrd+jgTvl296Lnp2gB3N121jOgpPTggDuh
8aeJs3PWNaHbOrNbUJuiUzYdHR8aftROSsYi/Y2oL5TsWXnWS5fox3s8mg472XXA
0/7kJ410XTcGg4lClouikgg7N14EVPBYcEjaUTygZDfxvGgFFHkWlMTts/nYdyKu
u3ZJ/LFBYENucDUR1E+v64eTcR5+SyoGbrzqnAjklgLTYP9I+48FUTLWN1qzStBC
idu3Mmk5Ck2dEXhoKWudEvrg0QndphOL31G1a02fjQIG474Asl7AehgONUTpF6io
lvL0GbiKDoDxEGZoj6h/n/amQAsIX64112yBJDJqE+tl47XhFjCtlujaerpFqs4d
QsqBKQiW/LEsd2YSGVNZbIQn3O6FwVbmFtBe4r5jzS4quFRWbNujEKUUZnIRM3NL
w31KOw0GndctqmIC13IQQUv7qi8hr8iOTyKws5t3b78WPLK0yI9Qdeug71boZhUR
J193ik7ifub/fMiHEPN+Amunx49nzZnJXUxJPGPmGY0rjpYrayGS1QRgbpSBja8C
mDuMz83uuGE8tES2BDn+0wrnI6n3NAyvwEvrKFoIGjePuhTXEvyFV/Iku+xCpLIO
irzhLn7FCDYeX5wwBWOnD1+b7rAjkHdSE5xhvOnC65Mu08KtAc1q7WkgEZ0qFExJ
ArLrfSRwa9bkuE3anp9rI3QewQ2SV0zvQ3VT2+P81Lo1uaaODTzOyny5AgupYauC
Q+FGXkydeZqgLELggNosT3nxzRHarv93T8MI3SdiILZej+JkYpgSpkQ0DRoo/AgP
wdVaLYO5Wj5qXSsx3R1RjbT51IJGqEcVCj0HH6VRUDDOc3JAYd0DgKjU1OcTRZQ5
fOdlvYm6Bm8lMkb6NK+HwGxVa3TOIi3BNzK6NYaYk/OdxsEcUa0NY6ZymrrAoUcu
r1zplbfIlsAolqsGQmwVVX1nMzlf/ut+TVovxWVyByl+pTIk0KjNUx4ttj9+Wnoy
jHtsW1KmJTx86P+YUC0S/fGnTmrQtA0ocpOGktMYLxDl62dekU4ikSX9JBXE12p9
KP7NyJcmil3qc39S4vt1RWsErFFKruXvyEwuCCQFQ5tXZRPU00CRtj3GJhIBgfPt
Cr5Cs2JpUF+ccoID4k/rIzcKXkq01CN+vMbcGadRopaUFJZvIKcAZzOfRhe41xU3
wdE44w8kP/zVWRfuDs99WBrcSfqEzsSq+B/UJIdVu/er2+PIwgE2W6NUOobPV6aN
taeahOKZOJrOE3sMs7GQUi2MMbzsigZ0E5FP5wcYfA/PwwSsL6IwW9rQLFFpr7kx
f+2BuVnXbyyplf2PbxCQ1e5EdaIjdeuxT0EMY0KAOArGeEPMwXPTOhe64YKl45TA
ki9VaQNbU0/01lKiESveakDw4ULi8Kn/9FifapLhc75CcOFHTob2HWuHflgdgNXY
54AndGh7HCcl5xouOPPV/UnqVRvHSFpRYVjOTUZYCz1UZKV+aRtqPxF9UqUl1Krt
4iYHHYGYB05t2jpzLgLvKtXjhNnechBhgbPHd9x73FsAhbCe7yhh9O2d0e3dIZBz
cql8RfUKT71G6WRSu2CuSivKfQMwEQH63XzZYno7A1VJtcTupq9trLv5Ap5uf/lb
MJenTWXgVovRg5d/jLx70qAtH0bZjBl3pLq6fzTp/2xl63APyqvPs9BIgI/gSHHU
DUYuH9e5M0TssK3MMtAMYBCk842qfHNh3qFR9HwAxd9WvddBFE/g33JwH9Cr7Z/B
gIXLgMmSG4SrXNvxImvHvmGoGBgaTOKGVINOovzxGToBR3EqhIKtiFhkgO80HGW9
cfeBsgW5BwlQovCVPV5UQegGKrB1KVv8F0fGKJBHsFWt1dAY9zP50jZcbRVY35Vl
xeyb/5UJTPGrGsKIWPjvcfzCgd3M3H8S4MQJQjIHPV/K7IlaSL4NP2s4OdALsA8y
xWwzpA9LqkrGtjBKUUDe19pK1j2LKy4CmHoRKF7hdSk6zyuPFwCe3cQPXSdFl8OA
dIRQlLDBZ8gjMaNyW3FlX7wL9cyvVY3ThPFbtsy7Ek7UNBx1K25uXkQGGP3lWj2V
EwT1frbx5C5wR+uzyalsQ+QP1BGVtwwLhEFd/zawxO/CpMp/W9XvC1t1V570IDc9
Uh5fvw0JAqFdiaISoIh8rhm0frpUcTEjuYn3bgBKIHZ8RTEoMQ2x44a4LGpBSjD2
Q7GotD4tKZ0iF30jmzytXd4w/egDOM48vMthIVrY0eieUK4GUTm0kAYi0yblKY1L
0Aax2R/fQliGIuwdSi/aiP+/mG1ABatns7SszKgE5P+dZC6vu8kXtbW4yN7zWJkr
ugowe7YtAsOvmgE0v2KSnSiwsoQGw2vrMdomcA+VBnQu4vVryySm949NaQgIjd3l
sIXjqSc6L0rStwhTE0EPl9zY8AYJuwwGHOKDd+5IO+EGaXrXUl19XCaNj/9l0uNa
UhqHVtOW3lSocEnpAhIULQQ4TiMflhnjzEwZWcNeInj/vVxnvyXKNUmjfN7q2X8p
S+WLCrVriT2Zvy7+/c2SmB0gO8AWlmL0obcATVfclDJEk0IO5gRrkkvrlLAg14SA
mU01BFFshjsaN1j2wxGzW4lvDXrv0zewKlZ0YtYFpMpn3k15hYlPvkbOqZJiJx3Q
mZQJK59ErpfWIJW69e3H463IQC65e7Rz4240aH5CyieDGD3sqvZp9KHJogmGvbzX
RBnjMtRDK7CU6UblOguTHRWSye26++jAlcj3MR76wyrygULurgG3Rlwfgnm2Mam6
T4Nts0i+U+Of4Fz6xHTJHuAt3Sb9/dRh7RO2xi4773SrqWoT8bl5oFGaKp739hSi
LYIYDMjiPpbYxrl3nj+4CBQp5j4sbmx9fOaJAOEaKOno1gW66o/pmZDOngfq2JHT
srTM4rp6CVvFZJgw6u1aVKTpbjF0H2DT7riAutKCtmy2u5sJ4IKgtTqeJFAFwYIL
RnsmB4XRlkcxJbDPU57C43LkY4sg+FBSTjwDfME964Hui8e0dz50nWTrXkMYUp64
ixdVE5DMCrKZEhkZ0JDlXgFZ9ZOHUhBbib1aa2oCenwPIXHdQ2KvbzcyccKHnneN
7aeg8hNhorwqJb282Nh7CnVtZLeMSVBtHeSNlacEui2JGVrT6EaLJr/+6eL80W9Q
jbRFcaL1rI43qX1EuIA5AmRibAVn2GoFLIfRTPkuZhSuPjeXEx9zitr3EiW16u8A
JmlAObBsAcJsk/vBVX7bLRKZLQC8HX6sj4yZa0Ter0UZx4xO8aDBMV6A6m+Su8Ib
1MInp1LuKZoz3F/+PWccwn4rSnmxSQAjjXj9+jwnDX/Od9Hlse8wveauXCTiGf4Y
FFHWqUmi+2QQ8SnMDgR7hh8r0nI1yOaN4K3Ohuo9yJlmOmc5wYZ4s75GbovDOKlq
ZqPXr/AM/XuHdHgzgk53905kYe3YthLnyEIaVKHHGMMML9uW4ZVRlBqOg92SPm/Q
mQ4rDlDreXfLf6Aia6geGITU7hTqoMBCvtt186/ZC4r15MkuQNOd2EpDkcsF2v5f
gZtclbWYq6t+jilomcgP9iWryQa1Rd/Kf6chv9mhGzPKH8ZVjeIqNIeKxwR8Q4CZ
d6+v3yngFzyAhlCWn3BmyktavLMoBewS22HbdDIVwt+0u4IS0k6s2+XLgbL43Qya
c/gYCloYvKOwe0sDtMju8uQIlhiFemx+PCSqHrcq/mYc03sac6OQUy8gU0QveaAx
pXmojrNvo9sgPSY1EWSD6Qm+WpEvElCpGlnGGmHoaU4FwUzSvkeB0glmGxoB3Vqb
/ys3/1ySsoi9PYjE2HI0akN3AcOSd+ETro0YTl2jtQI2ZBPt3o32J0ygL5hdDZs4
zcGvsID610YoG+imh1OdeIfb2sB1Tn9HI3EM6zSyonjigxvcnxBGPSSf0OLqvccz
LWDzoeLMAr//J73RLl6mbpIs4SEmF+h97U2KagU0mC7DKIMDbLQYStHxNRLtpNgE
rqbfJk4ikE9ZCAG5pgsvR7hevbbcrv+no2JJR9cReNK6ErrIijfYV1tIMWcbTxfa
BA2Xlg3+ibASXxdjqW8Sqr0V7Ds59T/uGTQggWNjqbDICmD8zf1ILp/muNaZLATx
VAlmYxKM3ClNbwHo5oaVt2Fqan2ahNwZkFSCyDlH7IoM0qpjT6/yi2J8zPCITEVh
FYhJ8SDekDaOexgq1TamLARjkpSFwfWzCXk6p7llvATOwhqdlXqU01a4kGPnm59W
5jBIG5XtIUG8IsmAr0T1q7hWT030R55KDrdSiLoRLztzdhbOp+MkN6WTKtMGMwir
Gq2gS3UwD/DuDGh74bXfYjMPkHmx4irI4YGBhfA1E2X+2mjlCJNEFNY0bPasLBy3
3sTyrwfSfIq9VqJLfOg5zyWztQNFI5nRYKwAWcEH+CesvK8NiYU2fE8Wd7ja8esT
ksGAcGoF+UkmVNKIrJMimI3J+BS8Kd9+F/jyGxQ02jywu5Sj+L9WouOXRaxsQkXZ
H+4XH3T0+DJ4N6NsS2UJbHg8YLhUK+UMwXX0lX5V978F+hKp7MjWZ+x9x6Rh+whP
/CLZXmAMzledOCPlqDY78K9NHFVaZTTSy6ctv2hcUy8UpjaAOt+FFj1u6lhI0hWr
a7ueDg3KH3H6MNXoVlal2EpmMQLpTUOKG3H2i2NiQAwRpKJtOyarKBvoYvZ4GA0r
FxTxPs16JgLMRnhl4q8oIkXlbYeTSkekxBRnw7w4BrSwOaS8mjo7nWRbOI8w4NzS
2zdjj/EnBgF+feer+zjy0h8d0hERdwXrGNS+qAcYRfc+hV1bmjyp1kqLJ90gEMOY
8xIA9c8et8SUSA0aJYXpT9O5/i/ZGunGGFXjS6JrkiDt5LGlps+44ocJYK5OzckW
yAoQNOKUNY9r2wCJMQMxJHwIIapwpDz7zbUzWetTubMUsbastJHHgzS2tPIN5eXO
Bu+msIbCjtBENuD4Yjwudg3eop6Lc9Wwpts4wWA1Mpghz4ODQHKbWhw0D/uw+C+9
MCeY39auHvA5z+mjT0VhmnuBg0g3AlHnlppYpmcaomDi7lzzzGMtd9E4WLwx1+Xp
PLMhSx/LQEtCi6TrIE47au0ODcnwt0Mj0Tl/ydhIXy+efkiimoUBBY//SUoVpv49
lT8L3C9Y+XolaUgN0jucX7+zeEz9GoYHK8kru0JMR3uuzdMImrEItstKzkJK9VHd
scDE/l7lrVx0S4a7B4Hl4k3vbBxge8cP1QXnOeGCPoBeMPmkETOsaqWX9onnucwK
LAl1Oz6gEJWybHVWNfpesTH1F+8LflOvbelJjwDTlCDTFo2+0/7x70l3V7hkT1KH
Bsh6zjYDQmTJNPErryKTlm6GBC9objUeNPB8KSXCnSprHNl6K6ph1hosxX2yQLCE
oIuo3oP039qzImlhT6vgLVL5Xjn+EG776CO6fmWvyVSoFL842+ot2hZWCg34QMzF
ULduhKz1D9JtYIRJk496OLBFzpKIiQo5SVSscN6D0ck2En6doFiAXYUVwmA/cItN
+099ZARcBWdhezUineeBY00taytZITJ536bu4Q8+qnEDVX1RBVP6s0CHZXZBS5Gz
EH+Bk9wz5YK1rg28R3mfw+fT57F8OVFj+PLt/6z412iE4l2SdpKBcsPeOsvm1mxS
/2phE5xlCnaEUzgFKnWlorDxETiV+OE10LPhuKag7qc47W9a8PAeSfphRqVqy6Jr
m3oxQBNEH0UBoJ/s9ZTYeT+mxDxf1v7Wtx6tbjxUtOdQW41sScTFFmzjVKBfcSAS
LxZGvWdYnxRyf/zKqKDtM8cENWJaOmNQ/Y2oVI+m3EBr6wYFUG7eZzVwGCb5qkQk
ZEB01Uzfgq0iPCbPT/cLZi5QpME7Ab3BWPNMn4e6d01lghHR69QraO5Wa7JKg1X3
oHgOELelmlcvmv/0ldnnodARoOPqNV4hDfV8ANGFW1lplz5T02g9UrOIjkFWyLmi
ExHOC/loxejfsbDKpDAhOxzTXGurxVgcLFTlMWWyolJxHVnUp2icHiD7Lux9ytBP
6SRJQg+JnXphoAO5eFmJfCRqAhXYDJAmEnFHwqXJCZ5uTaTliWefdxnbwiuBOuR7
faQ9cO6J2Ls7cwXIdPs9LAmIqZx1qwVB11XwfyNMSOm0WxuZQ/FnD8B7x5RjRXPq
IfauFPACb34hxx0ktzD5VICglwL0KksB+vlUqYeTyDcAVOhB/1Oya4pDdzx4B26z
LMcmy28/aPhkrJse5A+wf8hbU0t2ACIYy3uYBRqNuHIQaX6GzYAI3niHoeN3kWwT
yGj+GN67TB6uvuGNtJ5eZ7vwTZodAte/SkN6Acw76UYs6Xa89Wpw6Pbma1UqIAI+
WXhjwHhwY6FxkNohrU9aT28Ntt8to8SjgKWbTz0aEJ7nhLYzlbQi9oc+EzfQT3BT
LVfpVsL1envslqfESvA90n/9UQ2Wu9x+62uek3tLlDydvyxfpu8RJxP4DhiDhu2w
w/vcQ756pYKY2k6WlIXnCJexIIhniIfMOfhrmcLQJAyr4raGJ2pndo1FRUfO432F
SA3LKslEMQzzwQP/31qePUPmH/pHS5wP8CJijQVVJxftss6vqd/QFvlmJRzD2S/K
TvF5yFskQ2QL2bxAXzqWmKUFdSrjFlJH4c2VP079RktiTl1Hy8J+jjnmwm9O0Jtb
hdr2LHiNZf+mOOIawNNLggRZxPMs0kx0xt8VDf42cHOmG700eQT3U63Ei4bX172W
l1KwibvUBpT1L0TMKLedEQs/5LlJmVFJqe2LDWQyjZhnbBoin43qivaSiljYywWI
tuTPt/0Ptc45znCYrEsvsCX2rcYlna3Zkkmi6/hp178cXkqil4vzwScEVrs5vdzR
cFvukB5kBHYT4aWx9ZMKriRT6TAy8HWgf0x8n9/+zU6rASOvV2Kheom8j0jdZyuf
MO1vz4Jpj+sGKCB6F0QOQpuhEgJg9C1lZ1+lmwWibCjMhZ//vaOK1x/W8uJjE2Fy
B5BV4cSds3CsWY5MCY8vR7U9VhCjV0gyDTlQq8GThqoeU3WjE698xBiQP1iG/j5C
ASumesq1fCd5hz/ucSJrvJJruM1AMUSRCKQxSdMw0jbdY5rwUGT0roUFtc9GXysW
9OMEFsKwkkTpSQMe+NMUKhos6k/I4b250NQB1tXDQgd0KtMD9lXYJ3LdYUIjjH+z
4INHgpfsBmxyaa2/3YxQxebPHSYD9FBB6jqlc78AwYCbQ6TfVxt7IeJ8f2tHkr1f
0+ZelMj/5CM61w3zphJWXF3YARBRhX7B9axijbNEa0ozdHn3wxbMEEqMZfvAwuOO
AT4amy2a/Zp9QHPQzNV9AVgKMFTeqZw+FEjWJ8lM3oDceQW9jA2OYmJ7WOSx8Ntz
wjJ6m4Smb0mFIyDzSfHAo3VQNjeSVeX7cBKKFlVa5rhxlWGVAfCutWNBstE15f4G
IbYLaeFnuse+j1Zlk+ltnaytGz7PlFxSFwgoOuxtaFkhK1ileDD/arx+BVdMOLVp
OMm1iOXboPNoKXpgjCyJB3SL5uTpklhWuZeXyv+32yJzHfuBogpYPLlYq9PphrZ9
jkucfHR2Wj8NgYX2nelt27D/vgxrxRKXIbC6GxUbZAj5pLlUaihWPT0Q7V6a00ho
nZLMgT75rvb1LXO1EbUJJWkSmw20USUpO9LFCl/JGtVPMmkYF5nNCA4GIbaeZ8lu
zqH2MqRlC9YNuK/7dUhOmmAYoiBCyg1U86cjUL4iF7oWLjmS75SRKkEf7irL3V7S
R2UlFPl0YXb5HKs3QlFWOS1TtWLyT9hCJ8jQHmI+7noOVXPzQtK5ODLzKj6Tvyc6
jsnp7cnPWU2RQeyV/fhwt8HjSO51hfT3bS6mEioTB0QL0ot5HO2o6hP49ozvnmNp
MJYw0Ipsq5S+5RyFw+V3ZOPHLK13YkZsUGBAj3kiRrY1tZQoTQZeDUdgqFQBpHfr
IUQ6LEhW7acuDAflfBKn5ckke6iK9WmCfePMHH5e7LaNaBU89ZkNk0NohewzRTUn
STLYDQSuEzrotptjAuZ5qbg70PQP4vjp8pboxGRt0xx5idzm/juRtUbUEhAtnidg
I/825LKaZwOIJ/75vFTMV+qZwWVH28tcE2asMRZRxs/hPm+W4y8HAlAZ5P+COgI7
jRGrMRWopL7xyLQvXOmaFQaqSXxQaHHaU6gIpCxf/mAhshkKTLpgHpnh1CVHUgiU
Etfzn8VNRm46UAbDQStyeT/GfIkhADRdgluEoXjyliOYjX71aKWfhuGvkxr3qQnr
+4BQPRtNdNaFoUnWjxKstGd+2jrWbvPo8O+6UG2etdLK9iAbt8RT9GVdxdcPTNqj
KImcSacCVTnyCtRLE11rswKq5TyUzuhFdCB6T1oFj7sipweAcoTsN5IZjVwSztl7
pfm4KbxYKTtmrqoQ5ZsLTFyq8P2EbTtVC123uzXZHgyeMHQ7Dl/Prb4YO9P+n9xn
MMxatKdABXkB7yS0UGDcY2/tQerTMOTf7+Hx9tAWoJH6OWAEtra7yNj4dI4Tvs8m
DMjniRD1yRfRtNIFTO2W5dmrya7yT/ytrDqXaQEDaCsR8lwDrEO8yabzNVNQoEHu
e/qo2s6uWUks3FC+0BxwbO5gyvCZBui2wIvSRH5q3hmcGkp9JfKqW0KOiXiKeVwn
kNchMowBGvLULixptylZW5Wwh8+s91XTIyrq0M673/uc9DqZW1gbjsg8ELeh68Jw
iFnEPam9IhlJZc0VU0GhvXKPhFTLeXATpLmuP4kWAYa4DtgkMa7Rg8GthVQ2Zvsa
J/+ASzPm40hClOqWJle1t31gwsT+52+9sqPbcIQvJTwLWyH0fus2e1J1hQuCb9Xb
V3on+1uTb7HNStT5v0ClLLJGlHRCYmQCuiF2aHXWjYsTQBFYAC+51M3kXtT8M7hw
0MfFsFxlN34GWf/6Ytpl87IzTLVZnxLXEMd3imuF9G5cTY49J3MvXhVmtUZ0D5wv
V5WMBq2Gbfgrlbc4NlWqHygkUI+SE5Vcj/jnyl8fNVIfZW4Z78xzse+lVAZQc2Dv
W83/tPxZPoSQ4+BcOGD39vqDBeZ78krkAWziBGYVz+9oVcAT+QN2umTR3yPZ/pc5
i4Y46aZdxYahNKUwZsnAa/noJvzqbH4SQcwSbdEfESNTR3FyrmI/7FTwJ669tQVE
Ky9DgN+PB01OxoU5FDEQPuuPaS6yqTdds5UsMcz3ViuEGJuxh4zz57906zYZH7g6
J/4InYem2sJg0/b/UpZCvxWgTH1CPfP+fvEyaIb5VV0+mC99X3LC9Pno/xo8BPdb
ZiEfwYFPoVX0IS1DmRuWJS2vXv3jiLbLH89mbb1ADt2mJP1vkBkxqnNECK5MH0aX
kcCA91N8J662QgKwYfZFWppPn8kt80veRfLth1fdyP9Ucg8Kqw0igOqJoX6dJGe+
1JiJlO0PmBFX4TL9JZ0JZwM9mhVt8XKtfdq1LGb3Tny0Lky2I/C/JE22Our1XyiV
1D6RRG6v8RUcCdNCJykhWzc/d2gvW5nF/f+ALacU092Ru9j3SExisf1Hu2mC22ME
F5F5ozEywuaFiETprNU5+m2KsUTdC6Dj0yhsXbyPiUBoLZdLxXljitSYyiRaj224
/Sd2dXgB5cJoRjE0KQTC1+q6F6zJ5A8KI9GbbVFPOacoiQxiuCe+8Q3aB72bFvCI
GdFdMGDPB+ebdUoMX9upgJBFJFNl+fgoYiffbEnl+bz+4T5ouBUZy0WNNYwpgHsv
tav9TkC4OT6eau5y7LYE1waLUsiy71TZsfW//Iz69fwdAZmlz2KDrZO1AtuqUViV
TxhZBjAnhHMjbeO8C9M3h47P3vjoHV8zIE3helvZmMumOZwN6oGCc6xolurBKRDU
4aTNk5wdr4w55NpPccSxT3ql4ZPGBqoMh3DiNHguowhOdK2upwFITwTQzdLKwdxD
N3Q+v4DCfQjxsS6MePTazRcwisWCqjJcSrqd4Ty1QD7PhR3wUhJz/cvB00eYDvNV
6+3DERoDA4vNPkTV6cuwm3u4Q51uvzoDOreiMDzDARwI7CW+A2mRG0zU9k1r8Vcr
nqjMhDkz6kqoSR8VJH2v3o7tyhPOC+cHKewQJS+0vd18W02FVGbEya87RABY9U9E
+kqSGfem0ezjhBQfgWF5hyLIkojwDa/l8jTf/gcm4MclfGOynM9jtRWo0ZgIqUVl
+6nCBtjy5vY20hpUIYCSOYXFOJiV7I161EMVaE68QF6aEweu3AHN4noAJlagG7Ow
mISijVfYiO+pqZeNmLxyqZEetDR86ehN8Mw3zp3aMv6SD0ZPuPsHBB0PdZ8AcXXd
Vv9kd9AnSanvKWZ4ELqRvx//HSEK7IThmrlhB0dNOLjzSu5ObiLC+ygZkzdhSKfe
CzxG2dwZYYClsMjjDw35lFFizTLYTVI5NOcy8YqCnoteDANjC+/WrjNVXIQOo98j
2/m4gaO+GLP59ZbvHX9rznCwAer6Q7gASf59M7UevhvFztKRbmgvOqd1eQL3ll+/
Ihe9OYXGK+YizLEXnO+1EOZ0MHy+DCT9RB4IKqDknvOx3p0l8JMCWaAgWUrt4Bwb
gKXSWwF61nf77Qez2GfRirr+pvNc1zODU9p0WgIGsUMfVEsgjphCxvH+Qf1xeEos
mdPhdS98Ilz+Xa1QQ92pQ5JZjtbp7WvsMAFhhc4E1Ox+wKJUh6RutvAyXEwqn9Z/
LR9tl8pOkB6ZwH2gYhQm0uN2CoYV/seo+XSWcLVDeawDDFpd1QWWq0/60kYAZlun
NHoOISWxQJ3pOUQbshlEUe6x3xh1Cdhb66igTPTtn1y+Yhq59g+LFnpNz3sMEJ9i
kVDeqquXtn15ypbwGmyytjIQN9G3Mw4bl+BWaVYFpFNXR8iar3ab+A5+uDDlY7Vi
qmAazos5sfdwvah1KdjdzsL9Q6iwHpnLQbBfhYIIaERT2FKjqTa4n3/5utPjB25A
kFuJc1RffRWKAnGsfERAgn41hOIlDC69ZlpsliBWgZY0PuVLkQ2TrLzyojF+ktVB
cOehFT9YdUXctGyG8GpE4gkw6JGNHtFmUNGfWzct+jYOOY+kQHxmXJ8Q7u+TqyOQ
4O7rFZhjIldPEuGqf1gEuUGwTRx6O1kG3sXYuONNpkLhpFMv12h+C0N025WZGclK
sGTO0299pMObus0DchArv8GN8RqNG5oJgoEzy9JwviCbERHzHrlCOTq+8yLHg9ze
O1Hi1nlJ7GyIFHxviOcJ1QHV8frLDHyPggoJ6tFq7N+5NGO/vwjckY7dXzMMlFjl
/yn5ZxqBdcLX7HGjSl+vwsXqxCmI7Gy5KtWSHdver8N/q924lDOV7dfVNp1YNXRX
6yCNXUhV2WK2hXQ4IofJpsKJ7JdK5iWyOpaQ6PvZ9CdM1hSUg1IifyVG4SaT6ZM8
EqDrWJEWE+sqn0UaY8ANZMHtG22Tec3wWn4WRP7EXOSj2Fiz8tgqoyw/NFclYOBn
uevQMJkmsLfTUZQYe5Gr+hH5hC3zYRk/ljyF96JSNJLdNHVJ2SCpzR4/flFM+Tel
YDvBC/Pa94BcLnI4LXBb7Uj1uWHjHfbvj7NlCaf6myeuvTUbdd9sEU6DJv3/ttA7
4qECjM/CVDuhWA8pfp9XbK4DFMkv88OqHfJwbu2WKrgOqZjdU1cFSugSRaXtv8A7
GmQT9QVt9lqd26TAzrbAGj3YivtCv/hICVtfyRqheubKDVpSoWUhVl9nAoU59DZb
XQ38HIRumduShWDDKwKmLiZRJN8YpOdILMEJs/DR+NdzJRUatPgz1BBxGn5H63Jf
Ttv8RMGOurhOl/ZyTU4pvdssnxwUNRtBDT0Ra2zw/R0D+cP4bChXlSt8i4P71CJW
+KIIISM2iXldXfK5ps2S44cmJsOVCKJr/a+ajEGIvqDgi46/WfQiro5iwS86Xr/B
5+jUewZyd8zXoVc28jfCXW+p9S/ffMymo1vaFXuHsnachwKwGYzz0BwZOW1i6t9T
b9vD4y6DnTJnMnAz0tyA0EWKLj0/ZdgfqImW3reV++YRhm5GjN1YsVqqafCijyFR
pUgE98zwhaqbE+aUnf37Mm2xZI3H3DTE6ps3NG2vvZGkAr1SvpM4rXFiQpL3JqGq
n8qOu7xSJEr8h3bOwLBUs/NsnDGbcIAonr0PySJbWTdzPmxegUvuIs8Z7bX8UhS7
rJthL58POWpNSYi6miAN6j+8jXsa69QrbOuqXwQYHpnc7fuJowJcxatl+joj/EIp
mH5si7N0vDaNwuqfu0IzZlOBGY8+996uIlzVryd0N46b2byhhMQS9/F57Zr8cUs6
vK7fx5AK6RobyyrqH0pRvr4oY3KKlL3xYAX0VMESYWFpj5Fae5V4LVjSdyVgqET5
N9HA9CUpSW2n/Kn5gaCENDz5bPot9yplrPUc1kGtnd16oC3v90Fzg0xnvgaLxLI3
+lbim1YHIFDZep4QbYj43p1/8Eqfq3vpP7QMpuFW+Nr7pn8SO3WYUtH9FlJemLw0
DsX22tqZhHVwtXhrcAzXt5u5IE+CdVNqOcABr0c/qHBIHWb/e9Rl0RgjLxq1LBZK
eJxwpuV0lCHXAgWbMi2AU7MVKKJkElkjMRSqAplBZDw6UgiCsM4TWnzMV50ldLD3
2keZuK2XaijsMAt3GRIOjb5RiskF6k37B4qN1l7OQIERvWeYR79OM7rCyQ9dxMPI
yUbZLco+0/bkfrN31hih0pTqYgMzgo9QQbXHUEMfpLVFOk+fuPBTldlcP1iCrKlK
fpEwpHmrmzROIokrLN3zKFKcfIddSIhujvRjxiXDbLXkBvsPJJQYB4I6bCDgwHWW
xTpHTyPyw0lMtM4elyniqHZl/7mFRTpH7yp5d39ggrwbf2AueB8vZrCN3Ff6MxI1
Xz1ccuDhV+/SxwHEvE+KSaSg0zJZ9kJl95y9aD+hN4HQnLNBFM8i7n/haNAZJyNc
nppBvZ9FPvF6F7VSVSCbap9dD5ZG3Mpa4DnRq9qtZEJF2ZnSRaQGO3FmAECqrWxq
hTdQWTrzzoIHX/cdaUI4mezQEyTFCWi4/DafQfuuKHbqLAwK8ncd/p+QykE4e6n2
QUUjkx17QY7U0YPc/2yMZW0GlCxeCPwAmpUj6ZcUhsDXYAjYEjkAtX/f8DKQ4ufv
b8p9HKfXmZOIgw75DceoFyotyBU5gNNXkixTf6T19e8ZmaStqgI6tHQEW952rQ1E
bZSnemAOm8k1VjHx8W06xZySfcnv4/ZGhtMgwgQd9Qsa267uCXsjfK2vG+hXBNjn
UkTsCEAzB0q1nzNc47t/a6YvW0iZ72zY5JW49dbuRGzc5wL4SVHUMSqXRzC6rGl+
HHw1PT2STILwlndVKnsqKeKpR3Ge+TeSv8kiCtEHKQcV49Mmrj7CYp+5pijDwzgM
6ojAhbnuz2QCCsmrc2eJDH6YHg+dSrE3ATW+8CkODQY9/C/mvMJhTBk0bSiO32Wa
paCN7g80VMo3VLwcK6G7eup/5TgrRrwBuBHLYAGsjAY8Y0ylAbUjPMB+69Oc/vOG
J3/kdrtQ1SRzScMIS/A6qQ5wpQOOD+64k+VZJ+c12JeT2DpdvQ57GqVY/XgwBeV6
tKDDoGQHBMkApJDn+3ii8iYKDtf7BULgNwvJE9iH7vQxyMXTdWaFcBghCG1HYZLv
q4snhwxGTmREmN68KpY/nzdUeFsWWZEuUOdUwWkIFRNIbQ0zCRBmeQ5I4HPXtJkw
zfnIO6fT9otSinPcVaEi0TmIt0rWeKgEqtOry6IjdivXyUDoRXn/LafC70MwbWJT
w2JQmzhDjY9DlsVpxqK6iwdbQZv6VKoiRWCB+O5WF5XOqxAqm+3Jfgx0utHLdhkd
sMgCxgczQo5nDBQmsfEZ5bVAVu7SzVf9ZqHwdpQBnwNitSHh5MYttraF622FMI1c
ArGlzA6s+/ErX/OLhhM8H9+mJibsrPdaKhC7EbWlfcBQpqo9zfhIG5mODWr6hVhs
v0mEaQbQYQYaZLCO5/FSrRhAHy6ZP1tbYVWnq8T1LfTmWacQMEu5q1492/MdTQgu
4pI23txCkHtFoPQcy8KaxmunKpEDZ8hwWky5v7k+nbNbkfV5ICzrHzqEDHA1mEkr
qcsMSe8ZzwGufXkg2IpuEoPTKF7JvJThk/R7holmT0CxPXIvPfp38cgFxr3CpwIK
F0s56mwtfddz42urKfJNL0AU/yq2rm0TCwE+k8qG8YHSX4BcGPCUWUH/U+2BJfpe
LLlWhU+Xksj9icDSMxTleGsPC/2+22iR3YuIE5SrIqQHcNVRXfHgGBzh5EoUTb0R
cEcinJfT1W1qDeGpQ9PdV9iFGLE4iHDjeW6eShOjbV96g7sa+cliOJhdOgyEEapc
Wez71rCY5XnPUS+s7devN9AbOIvWegqLIEM34PuSfJjXjOSfuqZ7vwvSe8091UUr
68LmqkJbSISnwo+gYfTVIf/hkop6XKO1qE5UawT7JW05F/NlizO/QUaVprtRVyp2
IyGqTarvrHIa4E+Af1Gs+YRg6bUkFPqDiORuQ5ZvRhGIlAgT8RxQERage6iTPIBf
E9BLFFXunli/RvPoU08d4cTVRanfUxx0wzziTOy6G+4foxHseX3I5ev7fvnSaXKH
WcbsHtcsyGonf4JtiQXuRGPjCJ/0LqZTyz2CCpMZuWUUGq2LxLteMfv68goweCVe
gwwon/wNi8dN8tVa+ztZngPxNkTB11CL5NuCg9bpeZ/i4TlRjI1ReCsED51DMJfo
5uz/MsgJTK7qKnasK6DugB2xafJm8OzZGooy0DX1c85x0bwpjOiucWFv+SEk9GM8
91r8PILOnFAyHYz6w1CJiFLWcTGHFLz7/tim3CbTD58yNPUIk5Lgp7NodySN95QY
ot6ptqC6QxBqYUgid996aGdF2uLob+2ul0tPPtoHgfqF8QWFttAkKDjuzfugnjlO
nfVxhdorJydjwjc7KPMPr/ET40POuBTCjwbFcjNq+iP8oEjjs2/sbWjcF5fQL1uw
WXpTVqfRXNaxL64q3wY8TgCicEb5QKgHSO9MHlBsayeFPEgr1Pi1cBNuDlqzT4Nl
zdvSLjusgIxyOcG/vBkUEqCV26LfI3nvoD2TVYHIQ8zdSb+0o+x3P9ctFbeMOkBp
iHOwOkR2FQn+MFBmf2hoOG7kEIjZ/n0FbNk0EQnD7LfcoUnFwhMtmMV6DjdqgsZi
6kIC7Mffu9HT6uiNhjIMu+hdzrhE7VJ+CSNc15hQDpYauuasIXidpPksUeE3aN/r
8HJon3ZDYZJBImMk13byFxfFd99It2SEO5+gzsn50t3Xp0i98fskagFjiZnTGPFr
WpxvzAaS1mqtn5oi0aCNMSr4wl0k4CMqepq/nMox/8PyO9ia0HxRxur5kqLYgIvE
mOroI7Mm9R02Gpmk6e6TNGrv3PO/RZNUJdJnTbPXEGIBVEb8RaZX6gt8rf8rJQJD
KcwFprmzxuDFORhWhDBQDOSulvmzhh5I7nGLFZeu1WcPvKKvNx0XmSaKAR3iM3wq
b8FQkkNm9n/C3SylNbHwqUMj8Iu+GTADDed0OasBZZt59btDb2TY5W90ny9tucRP
N5vM5wiosZyN12toNBkaLb6qCuo1wQ+iOvjTTxmW0oyUXU9NfNRMErRVcZHs2uHH
OoGpCuzb6nFXXJsyvS2+FWpeGhTSDatG81ZepjcuxoHnWSH2YUE/L3AN1o1c7vso
u7AljaV/F50jTFhFunG5xKCZYstejGJ87H45V6IgKlN/ogh3GT86ZAKnslo5lLCV
/E9Q1YK1jhbff4Ejg9+iWP+BYju4mKNjrDQttv7X0LzGYRtX7TqZHwdJbNCpLqkr
W2KWwu/znx7xnjCXTEwmHkbtTTitvJhTeeGtN/FUovUDS13L4t5R/q+jl1l+hGJR
yKecXAh4H5XtOBSryUI0V6601TokNoppdLOqnZMpeZ9YiXirSlPuf4XCn23L9IRu
OXiyLrvOMLRHe2Yo8sfT4k83fXXdOz9c+q/oXRQC14nDaIadZviKyICyzqMay1Fj
Dst4k7IslVpWFq/3gTKZwyW+l4REUSZb1eTQrVFmoH0yDqvZfOZwsZtJADNf+PuO
Mb1UII+ILQ58oipnfrISY43R1DQWbkuzWMo7ueMIbv5r/QCdLTQE9ArbzPBjJShr
JJOAtOT7o78gpnfb9m7iIUS1+w6uFyjlhVbxS1HCQ0kW/D32Jn8CjEflnnILOG2y
yW8zRAjYIb8IOsD1x9HOtjr2FhFlkcjQa7bHw/cwbruu0RKIi557RUgoaPdjEehZ
lkSvz03PBapg83QIQO1BLK165t7t4kGMqD003Ya/jWIb/OtvNKREKDvMTlZbHfFu
z8S3H6Xy3cLKp+716IwYhXAYUGBCiALtkrYG9JCG9PP1hgI3+Xl975KWidTzwVch
V78GQdgE8PhGj1Aw0qHTGQXn0EQG2fUKtosB2pmob9bdPV4m8bxGvHtX195TQzEP
kQFyNm6ZFp+VNL6smeb3rwoRtR9o1wM2Hs1+1N9SLnFTH70zD2yj3cQyG6/ZoE2m
Xoi5l2ni5bUH0jCEbnjScdTCD1s4oyRMA1EntdX8ktzw00w5eXv34Aalel8iVDLT
yEQ+jGha/LSG+cEDBIFj6zFtIgw1qmzAiV5jrXrHMgQjIjORCBYQj9gfVtvonn2R
RPDg5nAgurByqIVZYVjgLNCGSd67x8ccQ8o5G3nEIJl979xpoROIgaNv0mJW4CW7
20D8hoJyc/NKLDWww1KoFUe0JenbEUflRSGAcVFhENKS/90fyXJiSDLuTd6lA+T1
eWJOZLfr1o7Ha5muzYNeVUgcsDJpXJWLyXkwLQv+SB/XaUGmkArKwTk1iPJafnCa
OIMphJvMmbwGlPKbdLa5tEcbpPOaFQN+rQc5BtgWhwO7cssrr5YV0DE1cqwkW7Wz
7HcTVk9z1SqIw5Re/Ohb+Z0ZZ7aoFs+Ii0FvBBQzN1AqGTJGqoJy/jJ/Um5Tnqkr
04sXiCKpjyQxzBkkP7jfOBPN/CL32PNV/paS6eW3IvrhYYX7oQYf91f/95lsPyP6
JnON/8b/cJU0pma+E+knoyVfUcyG/NCcl1mlQHcCELl2nGlgEaVcorqhwr4AynW0
eCEdofSawl7bqiXP+9cCV5lQrFgkhCAxSBXSms9xCMxQ1HH+/mEqImee3726VZCi
k1v6TkiEB529HEAwsL81LEEPySrGfSdX/27xUZGpAI5H9hO1n+t7Y0WbX0Kk0wZO
/0z7Ui8GYpHg/O0cf+jOb5GcLc2Y8LUb8uj9D840o6IPxHIerNsSx8HMm2ABHDPc
KGx3TwpTJNETqHUzE3Dz6+AftaRb3xFpCp/GO7TKE5Gicki1Sd+T6PF9yPTOmxvj
KrIPoKWKRIn19z84oRjRx0L9NRVFTSOUH2FNj1BviiZ60neb8H8xA8PttJCRfGLS
/cRUWuFDJoVbFgRnHFaiMG7WgrQX4hqPWo4ANQXCwJOnzu71e4NI2YohqaQhkRkR
849ejq+lROiIBrJCDu8lNUMjW+BoIQSkBd1i7DbNE0jsH7rkKoJvK49WtSpmEqdS
qB6tmAczLMUO5A0ZoiWGXbTp7mTf8BhA8Icii1jNTCxEYL7iG5yMwojmmwbuplFj
6UGc1oSIpyoIJemsfLAcm6b38FUfa9y21ryqxrJLNr5SFJH+aDMN5CqnokMpl/Uu
NKjMsc8SZUfSWFoo9la8vVbTqAOplfmb+fHc0YZtbsodAlvnxdFTQNtsz8csY/GA
vL0WUB8+QhnhFI900LwjPPVQ9GF5EdDqQkPmYakcuPawFalfFIGKoRc+7VPcbNEI
vmm8+iJLltcYETMg5Ph7mxPBs4ddK0OL3qjsOd2r85LsUQMePT6VHSRm/JnKci7S
k5+Lzk4tmCEveV0TBnqEtvW2/+0xCFoUO+MBhvUZDjKL6/LD2tWNcTc2sCaGya+8
RN+1cQbxDQ2L4OT3nddu6mEN/5iqGk1HWKaxZq4w+gxh3//Y55o+c+QDdp8O9KGQ
9QWW34CGJ+zwPTPzfcsB44x9RcsV5xJlt7b1v0AygcqGoKVZKGhuK+NzSAQfoQje
UbQJmiyIJMNo8GAfG3/6EzCfCUdAlsxHizRg+q81pVnJIr2AcFOigygaZ//O2tra
TOrfcK4fXsYigwny9SX0UtBOlnG80E58/DucCo2WycGuB/m1MNV9+jq3QkBNDuB2
hH71UIA/qGOGV5ZLmcP2/2mlQtMuYGhOiq4h/FLOHRTfy+20AS6Ol5QVw7M1Oc8Z
s3RFEJzxcff/XN4/Ig2xwPkg0Dy5Wv2CgsVc41D5JPouLTeHhRSIOhlEjPaPgycS
v6XO3AADjf9uC9OmigQQu4wEN+0FGG45XVoX/9+LBBbuWPI90HofOoNc+aYnBngN
N5OGnfqf8biPoEXF9/cPzzYLOgfXVJF+e70vi3oJEJ6s1d1Ua3eEFJSVwczIDUP/
1PHOKmkJmW6zjGNXRis95Vx8fnbKMgRVwRS9WRYuWp+ih4og+O1b48YQraOa6M1h
uPVF9Al1xstDigcm+jW/6qw7alcDEjaXXLcbOJtCROc9XDh7+r3Jy5V2kzD9lXzs
HnOYDP2XXCWFtYK6VCQBnRHLo6hw9c5Po6H9gOeHGl0/UjwTdT1vIEqe3A3TEzMY
lchAHaLOIl1z/awFBALhQM/lgQ32ch/9gv2fiX9EYhmk1zDweLFPUZi6GS+EeonJ
P1+Ie9cwUKoiHLsuzXQtX28AP9NRu5TkGTca3zGTECXGs70Lv9lL0Adfv0o+es88
AR1pU1dTXcKHJJ8bG1JnRQVzXIQSzi/81ukWM1gYSRf6pMpoAGsMjf0IFuzEUHag
hC80W3Kvsf0PCiugq3JISlrWZdOesMoSpEE1OchMHSNsq2BpoFn8h3mGKZc2Cn4j
eb0lAjC4lvKcr+uJDvyh9rconTqAvsECluPpUsY3qV0as734Ynz1B0aAn6C7DXhw
GMurC5b5Mc4+hmI1leVHROUoNpe07/+OkN1misxSWfVeEZxfcffoHt6pmmD3uyqr
rloo3TRzacEljrmK0pWR8SGptam0DiLlbvvbqXZn2WTPvUqN+nSbaJAsvWwDzEGJ
HSwcpKKvHAQorEwMMT1dl5TE2VDkT2cqiNFgFC/0Tpk+N7wsmgxJz4z3JuG9rs8G
FDG7IyTYMuP1OXX8qef23bm1Y/iIiPznF9v2ZXG1a1vz3rmHQ91kd+OgfTzjr1o+
8JezWGMoYJ3gc6eBLnBXyB875+va/nFY+JVMXFTDGhZWLqnLPMCzHlR9ygOqD7vX
sxhnh+XdI33fW4Mgu3IMHAg68eSbgi3WYxRLuHeeokAn3Of1o8oFpvs6IMHFpTu3
b/xvJd/p0U8lJpatUllh48hdRbauUqwkhwfbraXim3rHDK1qwx/hfqn2UtXfe/kb
xrt0E9BjwDpug1rZ5ANX8+UPsHqfgliCGA51FgKx34d7cGw0tio/qydYCx3l+2tJ
KtjJyvOauwn+cD4ibDwn93yq1pA7FhgW/H0j0ecFJD+rnh9CpVggnrymO3efjsBQ
jPLb1N6meagRYdB6KYJQcfwYMH3GpzT1KTQDCcNw7HIwu8Sfp/ievbzPwCTM/pH1
vxovo7C1r/haFeemBiUBWfW448rgLXDJO/w4YVZOvpWfzlOcCgZTu6XD4UjIaKeT
AtPGo0GZwpoPB4p5RElVlP7dbmtWolOYHMy2DXW0zaXCkzxgIVyfbERGK1kA7kes
cZ8Jq9a1s/fl/qwUH2AptgGdWjkAloFsAaMbc1U0LRgbtipWyO1PWszqBxY7c68g
DrfGP420NJePa9XSGxcBJKftRBXOgVrYiu3b6EURTT9eoTVzrs0XLXo6xxGkaBOq
QkAvexIyQlU9DecOobXvdoWgkV1e4t+qIz6Vx1Gs4hZujG7zunQgmRKxbu1UC+gf
kGk4C0+7w8yQL2S1/Lj0NvrYIYdOhssvvKEvtECKaOUPi1QcASph7fXaXQMbL9Zz
OBD6BwcxiXMH6uthZUQe1NdR7jryfBikV7KRgsRyHzZmIvV9uIUDjAg4c6Uv+0cw
/om9i7JXvC6kZfBk9eN+TnJ8ijKvelleh5fPMWPK9KE/1eHW4QxMEnGPC2VZYDmz
mgcP9GE6MFHMmFn6CQNOPsqedLBwWoMu2whIUIZmtaB5DpEmvI0oAh59gfViJDcw
t5gGBCD2zLQ4Xv2t9Onolq0CFndoFwKxL8mg4cH6KBNyRRg7yWbjclAsSF4O807W
nyTNsXAGVALcMpgWbSD5dzNH58W45KImbBLBT/q3IWomkrhpUSWbxIYxr0rwko+J
HXxC4tMzUwpM54RFXAz+QpU5fZwlpwvJTf0E+o0i3iDNFsgGZURV/w0UZxDW0rW4
aG1v4NwlrBmCLi3g5hf1f1R/cVGVC+/IhzbCFpOioxBsNijLN+uQrJoyNF3Z3/qt
NWy2Fbgyzv2OvEY9zKmU/9kX6PJP11Afve7fzwAKaKWwZXLe3QB9J3Gst914We5o
uHMsGsK9nf7DMlSrz9TZVFh7tSquFvylwL2WqL/h9mdTT6u10+NoTgp/E4qMxywm
e4eEnYHMMDyqV0rObxeLNM2b7P3TequW6qRW96kEUDOjUnwBB7ug5Cvq3Q+Ar5y/
Aw/0UR9ufiuq1qhh5n8acbDqoIO+rAfCb4Bg61v69EJqDs4qkj4nRY+va+i55jA3
PeKuvFw/5Ku1ptd+sKTwbSY+ItlJmPoVdGYz6GVM/UI3hSJkVEhc+b5aAOIlMQtT
2N49KcZKIA6J5LF3N+mXKVL+3HtBSxrpCxao3gdM8IEfy+h0z20BVUsDR9Ga7khj
6F1pgTJQo54lFGKYS5/9bkd6S0ta8M2hCcGAMDPUuqM4Dlw2/U5m5pWbFfpd+UkT
UMBaYv0T5XsgmGm9v1lK6O2N56jTae2fcK9S4Qy6X7NQfsxgLKR3QHqWvMvnFHOH
06AhmJRF+5OCw9Y23HkTmZpl8FmLmvPI8OVpxUSrhbruiqt0GG21qmHL/WMfebdE
sDoVoqPbYhscs13gymr/aHUZa97zu75qwx8vLHhajJ7TxHWae8S4+PfvlEr4bbnY
E1KFO3QA/0MOBR3BIhffgsH83YCOevjvCHTc1pDpH232W6npq/3YRSVaZDMYzscl
1gh/b1lav1R6rRGYdlIQVn+VyS6vGSYpSsB1rVx0kjhaXu9G9N/qUcmSFKdbhukO
xLj9NfRejI7zF8b2egCtMHyEx5ETGQMhMAaYk4BdPymQcogPcbZM48XL67va/fnR
1JIkbLGNV3MedThorzDVtYEsYzMr/GmnWQUy0nVOyEIwZ02LLp04AKo1wC0EbfT6
izq5UOYmq2oh4GdDFE+WwSiPZw6nL+mzCfECz4Hcji7KiZ8zG5WNEC015g6o9mmC
sdzykhP8oKUrMn6GAhbBrNrjtXfLZHlw6DtueKAISJcIUvsuUHCHpubhxlR/Nb9s
7xo/Fti1d4BnlLkt19wHTarQ8XKfBOUJuHAHzd3zBWG/QUGosfxF5b4K6kKns7cQ
LgDq8BdVSEjNq7WHMktYsEKK+ZNfMOVkSxP5nCi7nlkM+1OR0Lk7BoAd7IcrXbFm
PUhxTJSK374cchioaK3QFf6hNaIYJIO9ytq3xZbZeVfLLO76JAUDxoLVDIEJmxRI
t1JlBHbAfEGnE+gmIcWFBdFS/WIYl+T21WHm7ZacqABGoiI55PrY1BSp4H5TiYUe
RLj8Mali6DDacIfWfHDZ167QHmBLBSy+ma7GVBH+C5dO3IWLhFfqnLq+Wsv08861
Cj7I7b7lXKdYHpPQ5V4MCb3iruF713AIpI2vTYoov7pOZotr5wzLaYzk6zsEcDwE
xqUKOW/KKM9wXzJOzBqbKpvMWco1bE4kJboyr59LRarOEnrstgmHgOHJ0qwfNNix
CPygqyQ7uHXInSJV1yAz9Fc8BL/au4CtaBle3yQvMUQQOoc/KVXFaNX2WfrxVohq
tzc8SUMprXRCzvB9XAYGMMw/ExnKTbOqueffGg4BlnboV6zLx/FubQBN7gwHyWGa
dDR8fXr6Lth/8IqhnuUSrX5BXvfzJAJxagGbDn8z9halboKn8FXVRJ/qgYyitlvw
YZFiPNlVocURfFMmeBTxUIQXke/nrf2KiB4ZiPVh4A2JosrIBkyLeqtjC6yRYLeM
rOIsYZKB9E8DyWB+t5quTEKmlP70hE5rOTMxh4sRHWFoCHX9un6BgEWAz6EJi6kG
NrA3XvYpalwR1Mhg9RIVM4q9jilOFcZL27TFj0YUlW8X1A0wpolC43/9NI/pVuuS
PcgyIbX3Cz5UVP+u5aHuD8cJx7zTD9TgWjL+3e3+ObCtjFwFodlHGZlosrtpzmfZ
fPAfvtgBDc4WuSlUiNsmXatLFI3TbT7jWeYQb0520NAt2VfuCW1ovr/9W4JeKhKQ
GW9sUwxBdR4OcLegl6QqpGrLvQfMRyYQLqOW1ZjCSBfp1g2uwH7Si3VEiPDzZ4hx
eVLLI7HAqgLegs9a7PLV+07um7p27jhNfaelb+uxtThL8k5m9eQZDVcbI6LVtw+e
fpJqw2+HAXkVvT8TZdFVKSFlszMaBNumHfvwWpSwVjAmXaxXNqQPYdN38S76637E
sXoQJ4c9rsJovFQcmFDUq95rIEPY/oQ2hcD7aB/B/73yK5+iNFCRXAqbUYukiOhp
wpksXfW4gqNq383rW5cChXCz/t2E7raJT/+011W/SoXB9rLM9u36gV8ysyVkW9nF
fWsjI+pLVjJJ5jMCJFf0VlLKH78ZUKTRpRJ2Br/K6PhDR5YOp8MoAA2SZXtPQJsj
2BZmuhGdZ/9NKovfWL7+WgFwKiSQZni5t3WSjZmkVgT1cJpz8JIns2Kh3t9NDc2C
lOVFu34X2hlSDmfjtzN8KkdsQL9MgjTGLq30Zz0YvOSaheFNnOyFxpC8298mj/1G
UB7kCk1doCExVZ/+BcYHGn42m7sFob3lVw4ldtHX9ILqH4XkGKm7GscByRAIL0ZE
gJp4J0qErgOxeisa4Sgso2rg8h7WrEsfYfKnhPtgwEy6imbRZlUDrnLSPx/ToPkg
osXdYxE/3G1mACWR3D0TznAVuI/CFDsa0fpaaGTGCYbca85b9TIi4k+m/XA33wpY
4v+K34ePwOh/qNXpNnmghNd7RJJcAffDNWYX9qJJH6Cbkl6RijBm7hZtn9u6dvtJ
Ahc9A1c8mlCx20ZCCd8Ux8Rv6L8adZrvLQY3Dbivve0VKXtP99h1Ot/qzm5hMAty
3kAHjzJ+gAAi48aqn/EuS9CQopszqQT5btX5jroF1BwDipV1ggTQnQ8rGrz3ADZB
qjDkoBRKMUvt2o+Bwl3kt4bmKjCVrVcC4qZdW9PZMxEPCzkG+mmmKLVzREBKa1Dk
wpuBsLDRI89iMRt1PGQN/02Eq6yoFtloK156TkA0B4FBssCYijIB5Bra0PhgCMAX
O46ePuAHpsxvExraxTQdbMtvggKrgoHa3E163B42WGfPnluWl/URglF6eFb1wM53
jm6noUmvPZVK9AY6DeSLL7zvn3Run/b291j9gqsKdDsfuMscR4+IaUzdtPVjLyWy
Zvvm3acKrzgkSOJo1lJw09wnHI4RYnVSKmnEFd2QtEC5ru3LvJR/BvBTDP4uLzc+
cgCcJG4WIWsHIFSdwDoGBJUBkv58RIPfOmFLwGIR8wijvz1ZwHCNzw4fu5BqacgW
w/gpvBZFMJ/mIZioWL2ecq+oWSanR1255iUuDNldbnRmI5MMvkptOvNZWj7PjiOY
t92DSB5oTRs6Qzmbf0i45/Hl/IehOqlUz9BOEmyQDbFUXFDBLeD/h3pzA6loQB+p
v+6e9j2kHWEVbdOsEwAFfh6S6vP4oP0Y4M3/Samr4VOuvCrXmelradLU8HQZ+zc7
d+9lixi6JE4ZD38DvY0oE3P/b7TTd/xDgTw0LfY3jSnH94udnuZXaJvxtrmQaAzR
HHYx7PNA/zZbtSE/CUocQDxN8RBBapDpEJZSpYhE1mgi97nt1DuyKDvlbBrHQ9El
Yi+lNP8BUhTqOmHFfqdnsAQrA/CYKyfkSbTR8Y05FSucaBoveHyu4d41o3GVhGbs
+tPCHyCgQXmbV0zRzDUPwaYqFlEpoM+8PDo42IHXXMg6Tjxi4goekPrKPLRdd3qK
j4DcaniDpXczURPOFM5gAE+/nvtmE+KiUXj0WeYlpGew+hgnkSednXA+CfPsldCO
mQIJkvhpykSjhyBj+2ehfp13tKX6+szigOpwS3Gz+7bPdbEq2HzEqefyxTkilTs+
+3XPIhviY7ejw5MDye+xyJIlwz14bZa2uBf1r7EzuVb81Ga3q6GL5G+AFwcw27GF
JO0+/yri3niI2mXoX1mpeccsxVolciYs44wWd26BoaPT6zRl/VneHeOnpoFUgi76
yI0gspLxyZk4whJcscmkSntkz+bti9/pTb2sUhbcfzRY8K964zaRuU3V1Ew6lIIQ
lysPp7AdEWIoX+R3bZtrVJlI2G2FzzZZecdhEdPHy5UlO7g8cdYvY2UlaooDUiqy
V3nWREylGqH0eubDcdSj6wIURPe6gHePP+zhateflxwmSAPGfoVwoGo6XYeSUFqn
4z2uIlhuF485MBsZXedgWyH7Y/e5TIly9WIC2L9U266+2Eo43Y2KLikVNo6iHidw
pkwMY28yN4DX6vcQaKNDpMkJ/eFFhb8jMVcsnhieWN9kVqQ8ffssn9IaarwXFedA
h0hUc/W7TPH9ovbIA+EFFZnTzBQdisJrW5PF6pprMIeYzYBbPBL/NM6c52shWGtJ
0G+jcGWJF9Yxg3c0n1WDvU6vD+wcXSd3+381dneWf+aNCEfzu0cZoInbVRctgrSS
LLt+qPiZgDUfa0Nl0NxjrBHlIR1lCVEgqmmgFa7l1NfZKWUXxKSRBr6VPiJ452SY
4p527a05TUSGzztM/JqYSnjikTp60VQ1HGczVFZ6Qm2Ex/dL892R+5ObuHLg6UGO
nD3ew3fTK/vE9Vw19zU4kdfPxNotg/qgAJ14nj6XXOdgrnAHRyu4mTbkkyK3d8Qg
jtzJosJ1gvk3QXQRmKvs0NYjxEtbNmjuv9ypYpeea9kgyb6j3RgzR6GxeAC+YbYb
isyfaubNq9AodhARstHmMCk5NNKVZfxxyCMgjGzN/Jen2Z+YzfdkBco+p62ZdaoA
nrAR2oh2Fuk5LaxtwJHkIYSv6iM8js5yQL4fYFjcyyLppGFH2Me4NAL5XgiIJ5ye
ndJX/4svT1RKoa47aDzdRJ9qMuZLNYYh3p/PBLbmwHfvuVZkcyqwsOZFIk2p59y7
b5kog6FTpWDknnc2iZG6SkJqOTYGtA4FjcuytQ5UTC0G2vTLHS2CIAcF/IYmxir1
Tv4sygTFkF1PKD7vlGVlceIiFfYgzcdzypV2SPtT5+NhqetwsgxJKX7WdXbu7H5J
/ESaFQXrxbE7f3v+V8ZI62TQ3eUfTqb9tbelp53hZAuZ7vSQXpjIlERvUmki75gt
wzPTlskBdbiWJzk/4eqTYNy5au7APYX5wMmuyThY/s9+lnAK7bCCckawG3seI55h
Wib3Hf340F/HFbR2q+gToeLyMW5cwb9UWvzalrdAvao6oubOezrBBcHfzJYaXASP
tkYialN/X48mXMy0mL7q45tpVyd7Rhn/a27iAm7q6Cpd0buXUjAlF0lcaRV/djJI
bSjiZIAWGN5f01POyac+usI19Re5W8sk5cVdJ6VZ1FKmxUeOYOtB8a6vGsQD1FIO
fQ9EfpxsP3a7LnslPb5JVXYAZYyEZdqd7jXr0WmS0uFCPAfBZfHCUMwuBbgZr7LE
hbFPTyBbJ9/+QPuWYLdZsxzS+Vh7DfFQqBXDMSPko8VGpND6TRUDHkvSTKa08Olk
bkPEJtS0WUzlJ7kCcYW2XdOkVqU/uQOrh6J0ZKzkXgQLZOs9K6Yokx8QMgY+1y0O
wJsTacy5Q+vGoZIKYhAIKGxSjsr7UZXqFNqgZ3KS1jX3QSTv21w+YqjlNnup9dJb
LtLw7dNWOi1x3j1j6/xTUj1BS1pKg6c9UO3eiEaplFww3LHaRtWP9rl5m+mEwTju
wFP67PUHuKadxirhfLIHC3MDGU8lI5BOj5da5ug1WujqadP4aiHVHSEYHPniEWUU
ygEGrggv1uOhAz+ATo+3SpJvKf2znMCE4r7WwXDfrKir2uui79ynZ7vL2Hjb9TRw
fMZPP45sgRpzGpFTr4S1/Uv1n++YRM2/9bq2LhL5cDKDnFRJ3cXRCW28x43Bi2fp
LYrGX910VPI8kse39b7EQgJxP47Xtu1NiUXMvmxaFFpQ9dc9QYyimDcRzJx7Rdh9
vw/69nxDLmNJg4eR/T6Uq7XYez0XdYMvmVLK/PzGqVuJ3GlbQxORENFFIkcGVGg6
VjCVw20vA8h+wGdW1cFnmk9ZgBRUIpPMQBviiODJtmhUrKSziKQIIDMp1YlmYx4P
uWW6jb06z6SeyNLMi7MRcwTgnymZc3/USI6PIUSQd0FYBCWg7virzAKjRCULedus
8DIDAb+Ta6kVgXfT1w61B57RI/Zv884RhwU5A4jJz4Zc1OReOim4BBWIataQsMCo
zs8wSqHHo+kx1GfTkDhjhPwsZ+MudVnM/g0GzszBZQ1F219e1esVCqcA4Kh2rHpo
Kzl7ccMSMyLEcvbo6gSyM0mUQ916O2sogRQHlzG0zR4vkgChMxTusxXvg4+Qm9hv
MXUvLin/oHpkx4IcUEaNuU693eqXNGbHVs4f7ytFK2FTULsUFtoAmQ4GmPDHhCwO
TaHttBDnM9J0oKE4Kj4VL8kF7SXJ6Fj9ZnKI4g4+3XI7SEsgN+bXDS7dXrpuAiQ1
hRcjJZFaTeelddu9VmPVQm6nzwBzPQi2s16fqYas5Y9OGl2c3ZKUFEZHkn2Z99j2
3JjM/djFYUo/1Mryrs3hl9M6klgJQMI/LvYmb6LWICpMFU3yceqIOOg0RSJv+oMk
T3x63S8YXIrDLmsxPTPXFngTQi7LTBauanqL2vvnfQogTmhqqldHBSG4g6dq0MgI
Itohjxa8cl6TEiFnw5rJUioFI0n7DJCPo8WJM0vtrV8LAec3hykd64XYors5l53X
GeQGakKicis5jtTOx4NiJ/Zt5Fwfz3RiXegjPnCn9GkUiE+IvlAXARf/iJplrZOp
kXtYpVF9gK0Wa5NhIFYEMCrb4xjl1zb8No1RT8oJ89CDTQEVYzUJuvNpWZmdHxed
/kSXApNhETqScY4grv99WZI6S6mNSWYuNBdTnlopdiEz3Shgle4hC7pKoy212ONb
IfjIxRcuE7QEh91ds7YRoqIUY0RuwTPNee2apicOeN+60hubJmJAugILb1kOUCo5
2z0lLdhtdKvt9nEXSIWRTRtydvZa6z1rGOmvtWIrukD3EdaJMUpM6x3vxwPZy4iR
QV30xYkbxu5Px5VCE3q36kyQmp74E1Kejr6WT2yO4K1SLYa5abo9euYZz3QCtCFj
yKSMI86lJe3e2fO7C2POwCxqZ5U37J5DOMqC4gPgLB7cqdG3Y1/dXAoc14eCc89Z
BVM4eykdxx6PotsAMlmqGNVcp/o7GHmmCfNlama8CeSHRjgO+dQPphAgQoems25Z
5n2Ayq3R8mSd9a1I03sAEEorCfLB+qzbcQ81/dm102L4LC8yKHeYblwcg3hohNKd
elT5OsKgnmhP3hKoIHRde6o6lt43+LwxgWGL60jNlrF5N9tIiJa8QekG3IMYIWKv
GTYCx9tACshluGcVh+NJ+pTnqnDrDH84jsum2MA9HOl1uNrRPx7NiDM9QbqHluAv
fjEv5SxTdfec6XvXRCVXFjljclHEqMToGCB5NZDxAgm7f7RcqbdeGEVcYNnJ73N/
r5QCtC4odwCuLncgHp58blsryVMfaFfVNnDDEo1VydkITWo7jnciVew9HITuhI8U
AhavayN46bVUVlUAymkyim7yLb0Ef1B3nz5GUUvHhXenKPgcMUKgJWU1aglzVoAR
KWhvr/rjx3g0UzipQwU3WFPhOBBGKgLiInuoR+v6CqT3G83cHnjBicdnImkljLJs
AQTy0KzX+vMymJ0tLnBo13J6bhQI6v9eD2IZEPjZy2EwUFgwDTrshGjwh3baRNQf
YKsfpXSP6M3DBCPOhvssSwQhq43oHqMSW3vnpWFBEV71N6l9Ukuh22i2G7pRH19A
om9FW8lqPAED04r0um2bhRLJ7DV/6r2Y1ex42WCjAHyrkBzFfB+3fz+JTXmk671C
VoUP48qecRSJ8VDw0pRH2oZakJ0o8y6q/+7Ahg8w9ijEIv20zCPLcu5pRB2LPuFB
VeEOHU5CccARvwlhvqxIAVf9JtttYrgRR7DCNo9cm767fbvbGNwI8kdCt77Go0F0
alHcT1AtQ/St7JtE+k9bKI8pWeZTfzftrnYllJALVUMt7kbP7RqaaZ4IehdDxNd5
OKnduBI9EAzeVZymb0nf5QbO1IK3wYP6V8suWD6aURa4uVPuQRQbdwFW/eLJc3qb
LKhJ4bSGYuffp1pgNzyaAdofK47/cNHr6LzRlVgibEzqrVKtGh9iMXrhmttNjwb3
7G90AV/RrNS31TWKdad4ayc1zwK7l2dEVr/K+RGX3D89c9utv4l4qfdOeV/4LIrH
5J4Z15JWEzQo1+wRtQfC20HfZv+nZq0OCIOdnfoNA1p8yZIbDk6EblXtchDjK3Q0
+FVj6PtNRPzLYUyKe7y0Y79N8iHzwLORn1opqGgIOSnwLJGD/akjLqLVfmbtQTCB
nZoUYl4XlNxcw9i5T+pAjt5DagPAg6Oc8sAo6Qs+R1GO90O+DluvCeRDZp1g7wKj
C31gxw/feATxt9X+tgr2h9c6xohm/1uEvZW/ixXPF8HdFtekinv+1S/NueOpDW/h
lu9IJtxtVANT74aZLfQZTWiSoc3iAQIhM8kcf7GvwpSoO1CdOylCv8ig3hKbzxsx
0vjM4/lPwfkZIkocEjImQODW+aayo21UAW4BgUEvWlk0OmNS7c8C291KLjDfWBL6
cCzkiqdS3y3RBJWx17meutrwKzaDHkRlskA1+qsw/M2sk4H+MtOxV6uHQtIvbgfD
yESaZcbqAF56o4svtOKny8YgiRswdcj2Hqk2Gw00oEDLy9e7sOkFB+OGXVVpBh/T
Y4VYRfv36VjGBQRWsVkU3J5mecOHSav0PpNCxRKx4bUb63lf59mqcII4fHiC7Slo
hDuNJtN7hJFgFQuWroWOa9qE9Hm10438Qqcf7TTjPMCAS9Czp6+GE22XgnXxZE26
bf0RBxSSPLBHhJEaBZ4p7M7/rh+DLDgu+SFLpFn4g63/BeYqZ9T2vxexgSL+bcCV
9H5uVimr3M78sWW+MzI5XClCZXUXtX8YH4uS0IV4bxt0bzWu8nIqs3UKFNerP/F+
COC4Im2uqn5zlJppio+5XiLSkjQMRgPGP2Vp241dWrzLfTqgz2J4nS0Y9nCFkJFL
ODKQKq+nSAS2Xtno4Vq7TFPM0ntny+INMjbHuWcjL54hD4yMA0XjySlGpxUvCcyj
jCfZDsyvfTmsVTQUWJ7ofZy/TPCERtd4AqVI+fzdeElJRAZzvtsXI2myWSeONc6q
Wpu/g+XJnpObPB0N5KTyfef0IbbAky/X1hctYUxKea/FOIZ3SyJ1fJG5pS44X9jh
ZDEflXvTykkrdiDgznmczsvTzWJxjqf9sgFxYuUwRRA1/bqvpW4Ht3AQK22XxUfZ
H8PAeqrpp0IZZneHQBeRdC/y0BISbs5pXJdrZoAWAfPeICq8KaIP98evKO6EYnTa
+hA7F4iN2GulBX30GjJ4v9QTE9/fCrnbbL7tk+XgAuzEUa9hu+gjtZUS4Xcjop32
+dGoihYeteRSKc8hwFQBgXOyJBC9aoymF7sDsaMk6Ph8d+c9qhk6qzgeEJ34ZShO
56UUPoRddegJ5pwfg4HuaRsjgt2nu748vx9TSF/STVcJLped+fu+YYVLWcw1hSeV
94O02f32rk47oYDdzFc0Vb/xjAbXwFBlDkZ8tzeOxdu5yS2sXjtTUSeGOi44J/sx
j/KLPiD8bHquw0eL7p7yWnC13E8Ep4QEqN9HF2jM7NoZU1FPKyHU768nMooQqZKl
t3Zs1PW1C1/sMRvlarYbstOsXCu0SfJCIByYZddbhceEdkIRRqej8qonw/YHGyHE
kKT2/1r+jtV1Uztly0KRtY76vXXEA++10expSDG6GYd/Cp11ZJlbg1u/OyM5Mx5A
jONpUq8or7rOEYfbP7zZUxI1Lf/CNgwPHOuEGf53o/h/qfm2vIvVK5WCh2/Tyto5
lNyWNL5avL5FSWaA58yN86inUoEDk1Hbccppld6h8JQxweKnAmm9rnFQ1l37UsYt
dHahoZ+XsAPtOfBKCMWZHTMAMyp/Jf92TjKB1UIb+YengrUnZxIVzMSP4mh5wURY
T3Ei7ROLm5YkuQN1V7Q+rGKdbKJCY2kSsGSjKVW5yXYKgwA1O0pQMtP8UbYiFtid
P+TvlW2lij7hGM5bUP2WpJuOKdD6hjLdH6XyZrDjzL7lHnyrEGwdq4LHl/A6DDMn
kEyx8RrdB0REValERh+LcWkL6dz6aS6GWDyjFabasuqn37q4XUX+GhI2GdozsalP
VHkt5TIOIHYsItbgig3XtWg40Qo0+zy9G5wqiO6M9Rit8WAHsx8KnPPip/whAfQ8
ZCCWyTRcX8LwjKDynfIB5WVyl5Oak9ZXYekLwSWraADHXfP8R+EOXV2J5JXLERWd
SSapQJAIDI8FNLBLxogcnrg5Uh/ZFi039w2ieTTOul3P4SeBRZBpXmMw8EEh7+iG
Ct7d8TjmEbsmYvi20jAs+Sdls+xwFN0gPkWUFZNXsL0Hb2/1sGt91wILu5Z5pYdt
eeiIHP8IhP0BWTZmGfUZlCXQGryPMRpRXOy5b/3bphlQIYbj4WSVFXNTBVtTw8+K
1wrmI9MhNJ9mJCbKoLfM2hmR/d9YgZsFisRsV1atpFq1yymxKCMzPHpdoVIQDMAx
nJugZIEzzeNwG/Gmuo3P+J0DYZuzUdNzccU5AGlj+ZAzPNizcIIJ+33HzJF/NWcb
qbZK7x7gd6lrkYzB5RZ4W7jyv3ILmqwEJ+rcOv/Tf+BqYjI5vEVmSFWRfOUM0+JM
2Zzt9oYWv5y02wvRvO8T4qUenrVg5FnwGP4rwbi2uN65elK7CUGJwEUrMhUOUpfZ
KCT4BsD7K1DnPrdvlrys4BI4n/27/HOnp8O7Yhsz0lIPt3ru+8j1sBpmPJa9vj6W
RsuFam410jzsnS6S4dQT5OQmOcehpKxOVeY0Uezb1oTkuckbAP4g5/hzBvfWkEQn
XNSRdSntuj9Qpqh+8XpuYkyt4HU/djC5+h3oNj3+narzjAP6/113q7mgwq67/Haw
SuRfa0VkAdw2FL6laAE89rDeeJmaN01MWfYsX1U782W394OfFb3whGZfkGuFFS3R
xL1ps4LAeiEP9AomDlsO5huih5tO16fb3hbl4ily4X9ni7fnW6lcEfYTVdRcs5De
dbFAqLGScsk7SghgMgPl90E4EoPVhMMQRFhUHZdVqoBFBoSB0FcjeMZphAv5zkc+
4pEnjaWkv62RbrTFMqnzoD7M/4b27qS5hioIfsLw+SnnK4oEhJGkQFuqfO/HG2C8
YBV4Gm5xHt0UWb4D/ftwShV2qkm5HSoVwUBz8iMz3PQdKUZSQ0oOTX/5Ubl/5Z4c
S/Jw10fLz2RQKjUVEbF8e2mUazFTl4ljR1dfGHezldukYN5hsPoIbJ8i7vfAn7Vi
hB/qbUx1Bb2BCsR0WfHUy55cq5Zk82FzcP86LIWFTmqAC+mVzB9kebZK86G8dot3
chtkAdgue3csvm0azsHoBpu6jtFgjIVuUnaJyrDnXQhdoEqnmRiHgLz39kKDsNmT
UX8DbZ9B8d2/+yowOX9BXSptxiNTWkfRYxH5gjOEo2FLqhtNo0DJd3Tse6pcIBD0
nWdbJb3NLKoT/En1M7tmoBcYO7lDJJ1Rq2DLXwHdQZ2NjYcuZtVYsot+Qug4jZhK
J/X2+lmxplGCG1EcSGVPs+5Jg+2W3bYifjD6D6NRt+0Vr4zOVhzxCM7beFmuyjoZ
k4FKtietJlZxbEgd67koQqhWsPtl0qH2HwZHOuNJjN16GA+X3or4gkgPQi3v3zbM
xl/3fdqdPFHMiWNwe2tVjoY0aVlsdoy5YRBOl3cmnH89R1VzQhQJToPnP7l16ukS
hSF9OwSqW3JPU1vfYSAvW7PntSHrTOhXWh2IbIL9adBh8qh0v0zxcdqM8OusndYO
oRnBFL9QWEJ6I+SHtAzqfIFHwnmH2LK3AJuOkcV4ek9jpqMI63YrL5HLofaTBLZ7
15BRoUbHfQzA9aMl6w4+g2gvotPGYLhAQjc2Ds7RBbCdbZZVHBAXyS1j75FxNBP1
B29lE8X2sZf4XJuTJGhRJ6yMGze7ofnagnWO18yOdEbT/rFx773pNFKSgWJZchK5
UqsKAZ60SlrWN1qQW99/cDjHLMrwbhhbs2G4huEDlhXRm6tqX2CL9oP0x6GnpBa/
Cy4N7kmvbbeL5AP04de9eE3QzWJ1e6RBrsXIUIeic1DaVVmhOPnzA1JB6/G2/X+o
YxFBcSOw4d/paOpFfyBqCWWvawSunXIuPHeNhG0i3TRPk1/A4SSUcrM6WCNcPLpo
fxFRGb5bCcJj97XENh1+nDHQkiOCC/PCwgYxPtwEvcIAg7KOLeG7q0bHK5AWiIVI
wPkKsx95wPrUQ69XblaJlYfRFScdfTkk1RAEV/L+dRbMNJEML0AaHx/7OwXJBBPg
D1zaP4qPLE1EjOZsnIP/9nw3MVyXaIz/3psV/PbsRFTOsxm1/8ZxIv2192aJ01h4
jC/4BtztkY/7fiKcvvGepZJOiCeTVo8QZBBfHHRz/DUSAunGmFvcuDvtcPHmi+QE
kL4klDy/FDOGghAN0bIvWEUj2pJqkjVfncjM0Fw8u/SxU+udPtLrdAMfV/xe3yMd
5i05sqJx6E51pECyT5vzECgPYDHnmjFB93B5jxCYM1ZRGmflYVwdlQeQydXtqxPi
KOLOfYL9apbYYp2/xIF9Vkzhw7SyO56DXrs+r60FIn3jVnkK/Lm5J0OsAXR+VCse
fyCNDnqmNu7BWu3ymrvhIlaZwB16hotXEbd6aNURuo+Pob0T+1x2upHjcb8XeMtM
NYf5ddU2bq09thNQ7D50wSJkNiZRf7xrDi8uEtVy6sK0YdVTsb/F0ARbHzVqBf6F
btR5PWTeUySlLzytkXDytorA6NwYFr0LfhVonMVmT7IBglQtOZDUxQvWKZfYok/j
6ZtdpNKaI2J7UYcs+ANEnUMDG6Gmj3Ls9349+mbgCn3fX1QX1yUqUMYGwdV7n6Yq
v3+6FsPRKsp0FoqR+TLrRPCUBq2JVGDQ3GN91BDkp5hq5WiG1X9vasMZlocI24Pf
c7lem6tIDNaiQ/jdHKTBosL+MaMIsDHy+q19l9VROOFkOVq1rb0xUzU6I0h/gIc7
8YcTWfFNj/zB+7u7Hm+CgWmJHCDq3R2NYVupSAFzs50LKGv0ODyOg832k/GmDdVX
yq0hvWiuu7pygL4/nZkLi1wVtCmLfTdrFfDlkbQZbLHOxdGJjLGLg9AhI6CUOmFQ
uYeOHNUX8qYf9IdHogZcmKUFk1exG/K13h6YUOSYtNscXXGfTm39HbCWtiB8dmaG
5OjGM+8GAsQYsdmfNucn9H3Qo3kv5GH3ZwWWu46VPsZbLGMo/YxMMQO7LAcJ0cBV
8QoGPA/BPtOnYG+e/eZ2/L2zogYaAFRTL1JeHZPF4n42dRrc6wAfIH8YGsCr7IMg
wsrHHlqd7MqRk/XbdQ7pY1sQk1ZcDUxbS8Xr6GYVMz56o2QrMBZn0m5GJBurDZ4/
LLZgoId/khlTk4zIUL2uFJR+sbz3p7CX49M+yixBAD5wRrivgV9CI+/zTV6B0Kc4
GaKEGX8ev65oAz8QTzUvIWdw87w2XhtR5UCM8HaDwwrHJmEPnep/6eWu4LedZAwE
QW8u5PknsuyUvBwiR368IOC0mJR/3C98NEulIstA14D4Mw3hlwTMdFMezGG8vj05
NjgeyECuTIzLESRvYvYwNJwm0ONlYiwM4TGu+j1XosbA8YZ7fqOtbgiIeu+SBnfk
62q5Pfi+aC7R01cGMw9ijm5g/HqrIMfaEPGBovuCv9fEWba+Dw70MXOG6EPsoqQg
+LMGV6PmmjLS+PqwlPx1174obhTIwJ56oV2/sDjn7W3PqAivEYP4/575Lb08CQ4R
KHp7+iAtqLXYBWmDofDOvzLMJtYGCoKAQlrJwMxq2VP+bxguRDGNwkOgY0JoShWi
3u2D0/Rfrsm5gAosTHqC2+3MorzNwdzf5c/dsY3yZZitvVCsYDReKpstQXCphNGt
p8071IHr2n8rb6N8xBmT9u++MYqfST+Q4rcRVQSRuEZI5cKC79us+/NhBk9BMPHu
nN8ECW0l5xINIEGtkUrIRoUp0i7jAAdNqZX3LZnmGFXQNdSGWaSnRnCw/aDmnbgQ
jpGYLKgOtOoDA2RNK8siF7MlmkAh6SNe3EFVvJxt1uXmWqWrERsACjZJDQEPWYGW
Fui0YlVVw0e2VvPWB2Ht5g2tavXzo4aPfHt5G0s7T7o6lh+eRGYi7OsUAYb9OplM
s7WsYoLx2lrXiaOICnzKKrsg4sEsDc377kZiawjvVfsYqdCXz73Wyq9J9HCrB7Bx
tDaMs9GjSUI4VEtl7gb8w28Fq1jp37bw8XBk9fsQ/eIsdbnzEnFJDeDvHPZtD9wp
x7/SSoeblUvY/s7jatfrtD+8joEYrn3u+lI6NDg6OYtO83LFS1lhKpqhQhFZv7du
2wxfIC2U094xYbIP5M2XjlSoPikcuYXb7fftSetrmTeifXpeP0YNW9dYRbcpCb2r
iQCPd1g/rLfZem52c3Ek4f9TMgaQNFUY2weCSmPuq445PTDeR6rUagrxPe7H8kOQ
lUXxOHZtlRCedg6xyJXeEZQp/GS8LyUQjUzL0hA+Jn5VLjxuxjt2+iIljKwYZEIk
RndZiKUumSOK+UD6uf1D8ffzQsSfa/KEQsWm9sAvSziT5RQGDLlCU3jz/w2FM7FZ
YGt5rg89gcdKVpEfZrEfW+OyBEf4hqtB61rzsfgyXUZDRMJEbuFNdCa9tYA2FNgw
JSn3fYvXpKOdgKhzn+nTJxBhSzgzy/LQZVa7rLShWvReMWPy0SFuuGlFH95QMI3V
7eKXy6Iy+VuiPHUf/i0wKQhLSrLqpD4CWiJJKpqsNq6k5ISvf9YKr1j9cZsKLgcr
zLS6Dm/4ZC2EnmYxehZH3BHQQmKsmNfbtlqwSTAdPnZs2woaHs4+VmEGx5zsLZkA
4vlS9dTD/CZSvQoMnneqgoOTHMJII5r+xwwTsObWqkfP297658PQHGAv+vWtbIsa
4Ns69Hfs39P1TYBSOCTAQwMYP2/0mzFC6CHi/LusUEpmMrFoyb27Q3DG/V2Af/ae
oW28KdRZGVcfktjzaCQh7vJ4QU/0BupGOeyWU/Ryn8L40/vXpX+HA2gi8FbZDIlI
VDanb5oSpRv2xJ0iDZXDXbhDEnRJDJV7xwgHB6qkujArKkgpTugHHgrPvTfd2zI5
smFCVYzY0w0+iQq/ImApqLIlckOIAhkloP0WYWH80/pFaaabD4brTCLqMtVKcCgU
TU4Q1sZjRIapURIkmj27Pe34bSQQzW0I2PZmuLzRtBNiPwE28DibLoT4KN5AQVJC
r5WqYOuDaG1xyEYtK/NlsJ0NEZ9Hj2w8Iybb0mHca0qTPtAcplmKNWidicHyzSVv
K7noTlAsv33xdpKsj++FKIASC0OYMKmRqx1R1kWasQyr8k1soS35eDDaAGkDdXd9
70avNfdy12xoeAqSDTjdwxSeSnHCoLj/jxynspfcAOdhV530qJXcpXlDdkOob1+s
8FghYZiZJlKM+XKAdM27efL0yY+3Pd8A3kI18e52fSQYLvXez2XXn9xpWOyZtEox
mbuaeUJgzGfbF6sKkDXdp7wuJCw1Cb+XXWDFJCyhAIDvrAaaCzFUJKrd7k+7Y1Al
qnbgiLR9zQKeGpLLMoqIYOwlCwknqMzTG3vAud+yRbz3tFHGvSqZdMKrrUvSrLpX
sTT9fU/5VsylczPMjLs0ev6chhkpqZYHg2WvsXJ2nMHOjW18IGUJsfy7JoB/jBQw
Qxu3jY30V8SgxFis1zYbp5SLy7lpCFAOoZQmCbllLgIdytAprGKN4ScUS6ieOSf+
5mqiqZ+c1kTamcuI8bfuYeiFbVDO3RpxbrnpdpQxtjQbSLPxHT8bkan5drtx3wQ0
06b+NyANvIkl1WCSkglerCqudYMmxEEkDglYwCQuuyHryX20xAPEKFGGThZrd8+s
4xfNi5LnQiDrhxDLPeJozsqATFp1H92Q/RvVHMQOjMb+1uwiABE9q/tClP5A8+7a
ioztNsoZaw/nL7ea1AQX7bRIFUUtDYkxccYMFwvkbYMlPcDl2WN7i6xxq/0CcZcM
t/B3cFnoLcsEu4wSYjXQfB2vxC7N5K1R89JIkc9ygkz2rNW5ocDNyJ0hybGQj6of
z1hVa0eiabY2ZRjvzYUzaf06pzZbzshn0srXu/itrfyQ6YA44HBRxMRhn7aHxUmn
ESIwhB+9d/7qh+GxLpKbYEx/43Li0J8LmEQ+xu8pRDL6plCPkGzrHiEX3YZoxwz0
zLAQhgLM/BDrYfNqi96UjtA7b1O/CVlMNtOpx4LHhP/f9C73jsVAOroh43vhiyFN
Elz+kBsPaNzSN0eMU3GZqF8n69o6uk7Q7VNcPVlDU3JPy2yLL/AzIP08xqheca5v
YtvC5yCWa3V9pvCwdEfdEOWnxPttYcppCfPErbG03KLPg2njGCmvqgvAGLsMiSl/
PsjLNu6Ruk0bE25V+aZtI5gkDac9lFPwzciBB03UaXYNkKmoRB3+ZNvPip7rxBbY
1HiWhwsZVJKgp9rV8Gs5eBJliuFk/lXTzqRRURybq4DwSvBr5a2T2W2ousPXWDod
As9qhBxk+/4XG9saNMFDttYgeWXFiROvF594Vr5Bwo4QoLA//B0IBeTxvln4td6e
bvrh9x1CbL6Iq6ImEQhb5eI+B0RZ/ZzCTPzdZTFTmew4UxoLBwY98UFpyUDovUMZ
5zPC3YnKbyWaBpjNCBVeTQ3R2UIaWUEST6o3BabdB63kg/85qs6nAZjqmW6Phxsr
0bwdgBWyoNOPrZwxnUnsT7LNxxtBqfcK86i1HcSugSPFDM/9pPamto40bjzogrbl
4BAU1dCnykuLWJ+/4ahkd6TOKi/JsWsRg11c0AXBroExU3s4p1Ir+WGUldfQAESk
2QG3O/P8uw+fsjHyvgSHABhzbVbE7hLCq+RkgMxsdBWTXacg7bXHV4X6ToMvfid5
pbD+6x0b1XhKdacjmEycyq1/Gzn4G6dEpTJv29/2Ty2IT4w2OF4pOfRDKGVF3kCI
lMyammZu4riGzjz0SeqCm9GWAU9Rc2ZbXD9if9cSewzixSQ0kf+BAR/6sUZBpACk
2qHznilwIGaQpM48hz5qQdCT4+eSZJ33hQNHOY5VQAJ6POwB28cuYDnS7ad+RNZN
6bTO6LXyAgM7eLl3P7s6hnN/blsG3MCAF7OUTgL+B9SpgOoF/XHdjAKZRKXmhA2J
aaiG+AQ5dpiUeKshkkq7Q8qgJ/X5c4CEFMl3GPwAKVTxtAWcN7oIsVxyRSFcwGJQ
/1VYRT42k6kcZPqWjvBu17TuWsE0rpsfFqvoVOD3uPIjr1ANnOD/ns8PWU3rs2zn
cvpy6Eoe/QF+4iGkBlqrsSbXGrsAwXYurJETGCU7jghuNYeQTQUeBIgcaOtggOcq
wdA75g7EhUhjPgGLxRCB/oMOCnf03Q9O+La+zjD2XvcgkwZSfH1H8j4Knb4ljeOg
RBKX1KfGFwviTr3RhWx5ZjZnnFx0LyovRjYeGCcAR9kHHDKlsUx6aWvacCM8TZFl
jp4Np9/uXi6J+6ig5aMvJdPcZXfle40Tcy85m58oI+OSlECzgAOKbfCLFCfBsR8M
7txVhttLTiZQNAKzFKyD5hczjYlwOs/ImkRm/qg/DhnS/6HMwwH0455hn7ZHRBcV
UBwI3ai8H4ZoG5A4T9OaNeK6Ei9aEtd8CFClyMGTFAteA09+G/BXhUtk/niey6t6
D8hzAHLb0K40Tlp4LUb+TjwJKzoLYB/4CYk81LRovyK9r6FZmsVj32vk4bu6xYfh
ffymOCIRJQL4zMgtMKAoUMztP/rieixLtSTUGJzCd7aeio3Xzc94mAokBELLaYoA
ZLGHMpFWj4qGJt5IlwdxcGecXT0EC8qQYcwrKcuIQwTkkg6ggDEKay0etBvkQ48F
FwvAclM72THazAEamaeq+tgr8r1Uv1mT4S3fdJ5G5qFRLAKhe1Yg8IMu7Jaj3wWm
xo0re0et+nEfYi9vgMgqoOsGEskmN8ldHdyJXqx6xkxWa3XFMxEcRMO4RFJEUWy0
N0hVXgw7dFquQEdoduZuTfMKt3jpumUzwnMwQs/hozNLWj6QSLUtzcQkG6usSqSp
FjMQMCK7nOLD5QC/zzYrjFRiRGm+JRvX6YgKpeJl3+snJDbfnGOC30ey6ei5iCt0
x7HLsYcxh1QR76hmeKBmPdL1plbgZCQe0S1fbuVJOCHlNa/a2YaNfiHe3xOqW/iJ
n5mNY0xhbbpVz1vMUQz0AoHvcqyT0PxX4qHblTCahYUeC01SEgvvAVPDwHWOi1P8
LrKDSLQQTBfldCQijbpAZAF44ripBmylhggEQ+qobt22jkyz6iTy9KfMsSis95no
9MuhES1U5v27oiXo5EYqbxu5OR83ZjtwIl3ixqGZh+XZ/q3DN4yUs002+ipY1TPT
Pm3GAbjkGGHdZdBPdOpS6HL1MCYs/R0vXzk9KnnFqBH4hlHO1iP4fL/SRW+n3Tba
kajhq51taqJBZSaYv4bkIPONgkf3b3DK/hz1dAnaaY3kzT4dzREeaU46vbpFixAu
h33QZvCDvKTCZB5t1TnYVO38j9FaC0QloqrDm3nsM/U1KlYJhOO0B+HwpTtAtO//
NZLEhNqArhRNmqYkLs4Y9Y49YbdrzOt6PE2AxYGbJaG4R2LgwliPGtKy4s7wVpbC
qrQShFKcxlSCGme80pKe9SXL8gT6PlIcznPuoRWhDKyXbqZvgwqBMSXuKgermklX
w0P44aAOoOU7JbCw9BDCcmGoKAzj2uyjM6aoOkGmmexIBhVN47rBFA6tpAZV1TpN
iyT8kV8zFbG4v2LjcNmL+6WtTg9J7Fw77HMXcBZW9Eg1AlymeoEPKH1FqaGSNYF4
n4EApuugL590nQgjT9fe1u8G9T/6Kbi1FehBqvGTWDEPJCZ4EpBiFolv0ffdYLqv
NqdyaRklKWeMo1DiTBXC0UuHSo7x1Az1pQN6oQ9HmoLrSstycgh6phB9Pl4it6h7
WyJXkJkv14M8sLpno/5zB8Fc5mwy4/YytBNSgLUjvJzpir1SaAb2mvUs3RkI5cju
M2Gc3Abw1hrfx+mxgAzPR2TPenzUXQgI14vjathhCeY6tjE0ea4WwGd5bSP9Bsld
0xtvVyAoBMGJgy7cR896UR4OaEY52wc+b9b3NZcHzWMrQxu5eumM79czgTii9Asb
qn56+jnpckxhCMM+ynshWNB4rBY2eScu34YtqagxInKHz46CXEKRQU5s/mepCSkq
2/KgilmF7hBetaxnOd9LHuTNseWJjCvVqqM+ChML5FSnBrIJmuJ2ob91swsBk7QN
pQuqtl5nNeIi/l/syiHv9EOUx9l/+QoUZItbc2RuWVOIRRFZIqkyVvoMDvROdOGo
750igofRgBqvk91lnl6UeZYk//puS3IsmjmKKgsNbB3uEtMP13tvsfWlWdX8dOss
Qw57tCGBrD1tlN6wgaTfmFIujP7hngzsL8hceUKuLfF8MELm7iao2LkOrAJTYBw+
nZzWdH7c8FXysj4KiDc2SDRcvq2yksL6hXts8YzX9Wps1LVDcdoezs2L3eC3S9jI
66o6g6KZujfz4o67Li4KnYbn5SXTR/j8semTGm5/BgoEL/exMRekpyikWZzO6NNF
U9Nc2v8deJw4riMHflAF9aRXg5rVPYC0Ou97wOPeC6DMIoLJk/6iRDcJbdmjhAx/
5cgrcoKiIB7TgIa6p3qVP5CNu8GqxKCZKhYETU990t+FBvLgXXu4M/aTHK0l+rdB
U7bkd4SAXWU6DoWeJT938QhM+gC22LCwUf6iYuWP+IcDGhjYO/PmSF9qO0tl02LS
V9QLTZo7EyE4inOteRAd/t3gBnxKbFCjLf8EJVrfA2AdKG2jDYHbU3iH04QWzmYp
YVPSJJf5yBTNw+m+RPWeZLK21Yvl0K0QD8o9r3W2xUymOPmS4FoMt3oKY2GvDQpB
12WMevWXJVFozUDqjqb/ezrvYV/L3UwlF2kWXm+sqAtCj8MyKy/frRmbCfp8/iLO
QZ5F5MKHxONj+YIMZ0/Tma+kZQyZLSNd+yQ0kxnnQaI+BSvR0cnLUUCLt6ieEjFn
2KjoFxay+XV95YkFvTYWOeIlYl4QxizLjtYWevlyr0O9cvrvFHjTf8x2KR3f1uxQ
ToRz/RzF3/l8FmZuL6wf+YE65SPgrx4u0d9AzhDetarS+zGisgvwRaQ3MHmPOxhd
/c+CTocugA8YHBsXlFMQNAmSD/jng6HVyvEYpmDfX7EVoC3qDCl1AfztGzvkvf8Q
LZGluOI6kvfHH/u0luqBffm8T5Ys0Wf8JGRuL0fReRnoC9/et5lm4Aqu0SOEo8Kw
tTqJEny6Fnh+N/taxn+LDc4n5xqD0aMojuPTpssmiLA+uqtmkUiBnRSXKuEb4Aby
SaimZ+MgC3jtsl1lblW8TDHM0lQl9erF4N6tOMkEM5/i3XKJvTiRhGLQG0yta/ER
jKAF09lrWphJe82GKOgjtWOMKmcfYyKlqrkrEGG0gpqhOWszDDnFMmpkLkBaWbGP
j2umIxJkXMBaOnQjN8zfDUqiXJKDlrp1k2XLV1PR/3vQj0oFenztC2smYUq/u8QJ
aagw65zOa8dmaIQH94ASA7/2JROUf5mk+QusdOw7g4jDSkn+Utdy61opNZzlh+eO
pXcUOG94BGixP7xerxaVC/h2HRXV1F3cLtKM63quZ5qQf6Cxue/dqojgk1Re/AjV
rAD/bHxJ3VdrTbpTDwHOC9oyYMF1qSQPd5Etu/VAepGcC+Es7xotcNWEaPJIlO83
DUtESXVyuTIhoZiTogVgUtbiWzPDI47R2eo6wkLCqSQjDRlJB35gQDZcfZIRPfe8
2P38KDi7pb2nEn5CDteKVba/8QOTkl9M+4wfFLvBkHoEKHT+fCkpgxPnhZRdiVzX
B9KhWxHSdA3AcAk2D07QwJZPXEGq6bDO5Md3gF5Ry5NThh6bD1vsmNp9WUolqP6e
3bkyGyh8EnOlq3DlvvM/d3WQKVW1CNAW44ib8/RiCSkP1meGg/9txeNmdHmYUcSX
sD5RgNs5ToXD6B1mckN2+JF43rnCW7cuEXSboCm2M8Bzh/5dcoXGo6comLD0xTRa
zYQk6JQ4AV0gwpiQ+Co2yos3FE5OOFZC6pWm+6mqpmzyvQclkULRLHpN74/EVY97
OZsOVQB2BdLdyzs/e67Nu5eNwmezyA0x7E0rOjT8mHsOjfCILOWg41ddbt0zK+0z
4IHuGFiYlwhEj4vQwxuack8w/94+ykrxVplqsxiJyThYWSLBpdG9VJBb8nxdI1Ra
s98JCU+WsLZ0OjR25i6rLSieErq0p3udFbOwUy1TB0sIUXLuz1dHnsdl5LDjGNZ0
JcajwwdsdiUJAU/xGM0+3cWPYT6T63AYPXOFMQm0RWfj2ixw1zCpQPhpCGefI+MI
YyFU61Kix/kxSvg2MSlMv5R+wR7Uf3IzkozXcCOU05CvEWCYPgNr8YqHEsueb1ao
iDPGZmEmrcHSZwudXI9zup4ppYrcqYOjGgPIHQ9PLm+gpIV0ZjYMOwA6z35pTYcl
0pQXrkObNkjyS/pqdp5ylMXbquwU7zBhti0BxCM8aYPoHV7twfpHdHZvJxVjQ8hh
7LuZ3PDFPLc7rBUCLtry+I1u8Fg7/StHsBxsVYKp3rs3yvTxmtyo1XP1l+rC1OQI
AwzbrKuBKdQbY8LcuUXtYKymhuMpRXLlt+DEW4QG4ijs2aTG6thhmhae3+SuvDr+
OZd5Yqismn243OviVuwM0Ke6enT+emBwVeseMueOrzohj986YFr8BXwEWICWFYgF
COw/sWiVQ0AEyboLmCGgrNIsJhgXkRTtdR+WFeou4GQFo350+Q25vkgRl2qYjHjY
Tr+B19qEcXYtkFjH2RRp6CIBAuWNPL27+Mryd5qhXJ+mdv4zXmYI+7fjkgdBExqv
vv4Ksb62fHAMJ3YW7XPSrPhy3YsoAXuabOlTtrLrOU3nBsIEwgL1o7K4jKLSqeX8
4Qb2aqpVrs3sROzTAJv2V+ojDJJcNZN4rdliAc2If8BAT9+pb39MU5iGgAZO84BO
J2cgFuSfNoJ8twPUQdMaWoTLdtaIEfreuL/D7AhAI5rILRbmHlMWraDRIH8Ubuxe
mi4y2qrmnOTDLt5eecrUxAfdhJbW1/YMcvs/RnbR8Ng8w8bNxnc5BXq+Hg/MbHPB
sxeDWcOJtcbqBUxPE0hjI8piYrVxaTrSX4CZMhOvixaoexpDY/gRtZ2bgdfvlImh
LZYYdOU0UfjEGP3PJvorlmQLOhvzE59IW4+PZ55qZzcn7hb2USqoaZgYl0NAZhqZ
bIfN22yq60DB/87WjXijwln5DstwzVC8X3WeOwdMOxrrXLnOLFnVimtRlJt9c+FD
QgYYGcn/4Vn1nnXxNYJ2fmOBqF7ag0LnQN86kwfR78MsFPXEJ0YRX5PFq2zwsZuN
GFTK3D4RuDl9vNBexMNQ1KUSSOicrorU5epqEcxt+XxhZpkqC3KZL1C+hm+8qIJa
ggStvM3CN+BnKFRxR+GNZflqH0M/SWUejs5zF5VbOkR17nZzopt/PN/nQRfiOf7W
69uWkUAxboYhE4MEtHbBwuGavLDlS3W25XaE4AbYKLnPECGJyINZTsNViECBBgGx
P4LlDq2QJa6NDv52nH/8rq8LlXVmHVhAzhtw0X61pAXQLOCOosXN4mZ+QZ8Vo7Yv
E72jJ7jwSb+9xKwBKzFAXlolw695RnDA6B46ssmJgo3OLZ1hj6UdBTtdFc/c6mlc
hfUeNTz9zmXzpqYyIvZpQnrTXq1vmTbRQyFpPZCZ81CQaBjckRXbvPu3iDODdhyK
gUmVyL5Ty3ko9JirBulEkOU1OEOi/p7b6EX6R4YI0YJo5S5qUfpMCmJW2XJuvOZw
dEIEWFT3gg9ZYIy67Y0iA4wTsm4C8UGB0Abj/IDkasLVBgmTLsff33A+mOAJMCGf
sVa43WELJ5UeZ4clZjbgTVoSEel+RM+y/MZZwur/CtRZakmB9eUHMb+9o0pg2tTh
a/j8Dh47v+IGFxKfuB9LG0oP5N/EFdcnUmmpmqtXaxVTIAnySC1Vu+8NM+sAxN6S
UL0c9Hrv8Dj3UJZaszwc0FtY0kLXQEjirFA6iCzAiBwbQHqwXADaoLY0zzCSY0zM
C0OC4q64hTpuVgGL0dC9kxK7LwjGQcxA0882F4FS8x7Wn0dCnksolYkGJI5C8dK+
R2bb6/db7HJe7jiLt6YZCIxI1aonEk6p9ztlD/G1LjMR5MFz0K5X5vU8IWETAqxl
uvIuo7OKNBmlVT3JYhh3yI2LDni8SCTEeTmfgZV9Tdi73TR16lurSzuHh7Un8Wgu
J+Kqc+Wk676/+coQr87J4ND3NKb/bbIsOdFdssyO+yXwsRmQWKFkhmRvmRkg9K48
sV41QQkkssW571FkJjIEdZtOUqakrU54ogqsUZ1aiAyDDxhNuCCMI0Xf9Z12tNjb
W8jj6z1dA0Ezj0iNmcbqUhDIvmuKV34KGW43Tr3I+7KyClW6UWwt9heor2S+yJyG
asIFQSXqJvAvvZ3ObU7sYL7x49gp6AJz9PCXBpg0gRMoDIA/oEiZ6HYOj+TWmB5C
ArZNUSu05jfcsgsP/jkwN72BXCOWbLTkww7+/aAiK1/XmudB1chRtXqU/TcbPpm/
E8UZxEQkY4FSbN97MIX5v5VKzUaqJ0zXgcJgIBAoYsHo8ika/Bv64/1UH+1p21WM
NPQZd61mwiHmvD/Bl+T9bE3f/31YFv0S2HDoFNZkCKjVjXf0tO3W6/ck2ocgj+il
XXopfhe0mEwLuw7yB6ab4/VxKMyZG4n7Z1MLFcAAfybWXIFcZBrbA+V94tQUCZIo
rsluMNAIS0+5JzYnIDSvT5FGW4Vcx9UXdcv51wIbUAZyL1sT4pg8di0PhGROpb79
xZKfI+ze/5R8WWaZxv4Vl3b9GEpMqaI+rmG1jEwAvx1FA8W2969Nv9E4Snwpri5y
+T1ecduzmJ4UtB77J40kS3dwFO67eP7NiTCiGbUtTPSU8L7bQpkxWY78A87jmxn+
TYhhxh4XUP0XDS29+3bh+bYfwjRwMwnvUIMcoUYyoFGOlxPXvUF58Ya/bm4Ojpw9
RK7p3y8pcRQ6qqpA4diX7lZrNcytFxl4RJ4383Sh9LmSspJWi2BFuaNDjn/J8lfv
COswz6gdbd5qcZg+p4kQKrYlWREivKooC3M/S0jc5KuicCLdasSkT1zGlKBEZD2y
QEVJMuxwNFM9hsoGe3T4WSDJYYxYZK0pzQiYHBokTsA2J3U0e3RxPSLglN13CLOM
016PHok5unettGd4vjpawxEQ7j4nB2fUFVLSiLmhp2p3tPYmB9cHwksJ9vGfC5mU
okKD2iyajgsaQY8BIeeWtA572g2JfXEKiOD6uj7GWuaTLzI0jjicyQlZI+AbIbqF
TbHUAsublPYHq1JPv6O0GeEn6ku7R4NRpCDi7XCxoJLj8jjnEM1BML/7uNAMx7aK
l/9ahfO4q2mdiChTnDlGJDr3xcTh/Q5Oo1ac284VfRVwuKYktA1FeKFSCCQ3Z0S8
62tXVYnbNNd3zp9R0/0S82yAuTJM3ZkS28WeBYUIwdJMrqLhe3Jb2CmDROU9nmGK
72LvpHgTuOxxECCpli97SZs025CBXo+ow49wlhU+vB0n0Q2cfwob8RpRl/WZ5TVH
aKCdVQWSSfCgrb8NKBj9tPwEQh1l1sj17UcrGyuiZUERXUHVbBkhTUclKDYPpFgl
P2f87819qKWEhQDY1xUwk/ieRIkXWNp3EoA3MyQay6IIA6O5Q7DBwjzEQMLYKvD8
mFPha/B9h9o1JHsqR2yFuLQFVSqsytSveTmG5sY7eL1uTYHRb6t25mcm3gh5tj4X
rIX0aQhjCuTdM/yjJqa/UbrVG2BE7q10HQNtjnZD590D2bIzEDgUZ1Yg+LOsGEeb
Orx0T6b8UxrLnJL6bhWF/BdP6JtM4BGVkZQOst5FCnQbPqSREbH69TbUAcOtI8Qz
Ql0p8wohOySOKrAmAW2fuIFlqhqew9Ayd+ieWKaoWixkDtTSZGId00kjyt4ElhGL
XNTFlEN5tGyEXF8w3LT7Pah9XgRM/S4G6nVpdNmPA89RzFZMpD3JavQ3EjQzIJAL
pWEwBNmp2lqL1rcnK4DS8h5KRCXClpZew5HEXSKztHO6+WF+4m6oJGEaY4F+W02P
pBkpZjb6XexQDDRhIfI4Eg+d4FmNsPPKt1KzAwDnztTwtwfxhPf9osDZnBNXmmOx
CA6DEnpx203ThV6+/h3oBQ7jvyNuf3irqUb69MoAeGYae2bplTXTpjtGRYzDbgZm
GxM5ZUl6FjJ+QMbrGgFSuPCG6D/3DQlJ7XLxTKJegNeW5uDYugok0EfCyksv+l1P
y9lx4jk5hcD9wgodYWQgpum/49qgSkk2qKHwWVRY+NKfIse8773bZYTxGFdve3QW
phQ6CoEQPwMIFlordnU2Mjsni0i6CYmr6yvnKm1THrHO/t0PCPvJ1kxxVu6HSyVw
YZOqZUqFSbUB0OHQPqP+nnnpqN5xyxxeK2pWicyCJqbjKwqo0EBblVQXfFi0IVCe
zeDM5Gk6T8pC5hDQOevpuY2VC4iCUFnQeWNudwvB9W5+I45mzWVVbRpvKBY7IMCS
jby5oIkqaGKv//g8FQUAy+jg+3yAuUHsky/O8cLugTQH6qeaXwbeey09FTTZCeBl
aFVeqnJPG8Yz7wPD78hksqohaCM78lacrUViGSakB0j23Ri3upXSy7sQuMdgOm/E
twxg8aZ824FcTUUsEBJ4ryFLYaZT4t14212Dq1U7FUGcYS0YVbd9KRB9sk1g00Gn
uK0y2BgX5DfY9WkXK5FIwNcVMei4nBY4rrueEXOUFC7GqvKxWUpUiDhVjo2kmK9x
Ssrav6BRPzwHRLH2V+VNbxkp7oaYNMt0dx+2B/fQQToAumOFIj36JNA2G7kiyY/6
ger0fVDgHlZCfEKKuXWGf8guGUkPjsLW++bw9bp1eHqxVwwL96ByAEbO+yYwH3Al
PmZ5eNJsArCI5f6oLqmiALnWSaEaZIAUlEEw9BZYOsyUNaPvyVTrvV6FRCIgc+bm
rw/0wVhWeWbqpjFhOw59soGjrcBUe+I5mI1uWuzvDDWZ/yDWiua0eEDC/0OEbBFY
1mjPL2KGXZk4YtLw1/lToZSuKcMW5L65h+qcjvgNRMQSoqPOsCGoJfAUGBJ+DmhB
0x8YJmHiA4pSGALMHnLM9q8y9Gv0vv6vxa93UaDAT5MqX9nf5/f9wnh42qieMkst
OIgtEEMztyVv2gZ7vh/LA1tTGg4w+IPxuexksSyOhUZ3/KJ3wwpUA9RkRMDBA6dk
7Gx62KZzrZulKpQt6S3XtoWV3yIonpwQhb92mZH+zf1X5COXh0Vvk2Iccbgak3r/
EXRl11cQKpoRdj1DGBFzZFStT2FyAK5Z8/tpOiwmbJa1XWytTIPbaOExZUL68Rqv
KMwYrUUtVBME6Kc21p4Lzbvt0o8rl6rbNaMB0kimE1TYf1X6gmxxqQFaBXGCn2TN
y3oQbE28noUxwo8zln7ARWIEoy+kfsRFTumfHLuy29S3xDkmszuplH2W+nzPTW67
v5JUcrb+apl9m/ZAa0+nCrGlmUgrZvcasMPWj5Cnllj4GeT9jhkqfRF/ZC1MwZUO
DOxTD9ii7T4Ib7BgHMezEQteOYs4D5LsW/VTHg15UV/HhJCJLt9dq3eoG+TFEzzG
EHRex+wbWIgMd27DbmAh7Y/egISIdEi0gZXBCotIwql6GJOQlQl++8cB6tWVAYxt
kJ2T6sgZAQSOCUP+NmEuttpLqKCrBNufdsliCD3EqSg4RVIIHfhdreIYG0vAzF9T
4I1rSZs9EOFnoGjvIXBmAsmWhd2z9AOtUvcwTVhlsHGMmEciSd9+JSHQv69FAW/o
XBlQGBcHDK9WKID4s6ebJVVp3YAiwhx4YXqUWPRKpttrLiHsU7X15Y3oMoP4uDS+
mO5cSdI1h1eXW38sFsQfv8dC8N7/uCDlzXwr5dZdIW5Jxo+PETeiDsMPno5Qf0pt
cLPF5nVCcAcExPpf2ZW8qE0q5VOy9T0feW8q7D3zmV3PfxB0iqmXqox8L+FDzJDy
p752PTtqQ4WEsqKHIklgCXaq1c2Vk1tXtdkO0hLwUylFAXFkdP99U4Nn82yiItXI
+u0PsWqcWx96FVGpjl6a6SrRBMxM1Nl9kFP/ZOBgq86esHoNCTRi95vEdN0eFLjT
t/HuW0qaXHuRCx/mzHNjdZYPeJ756jpNufPocz9FDeK3FornITXpN9GF3VUP87sX
qQlCSqMD5YhIzmv3HU1kECY2CjmHN7gAesUl29NODJf/KV2rdsop4vW7bQ48ZWyG
7NdxAwUemokpt1IH7qTqQiB3NCpXQBjVDHa7/C8uyHeqI2zgujVx/u7qiSD1B8td
/fUQrZ9UBEnqnaL+jHNi5QeAP/h0XsTfKBcK6TNpUB2OX9ojYabUYyAGBHhg+A4/
p7VujpKDthLY7oWQEErx6CjlZ/8+bYEKd08sJQiURPWfJO2FRfBlp4fRuq/rhb+t
NG4F6YvdBilJ0A3f7Gcgs+iT2+Eklkjjx9ACGeqTgLFsd3BYvWO5O9JyshKsvwkH
ZPpb5xmamJDp78cMqC5R+LGx/lsOnDX69ypZAmmkSPmMroWYnEnH8/qbdj3DJqFi
TP+O5uC5MqEYtzQB/TZIgdX/AwONtC8ak8IWekkUrWpb4gzDM8sFbX9a7mQirGOe
cO6ZNhXwbRemCzD6VHlDpmf1pGINJ6QPMYugWdrRCCSlpNItfR6ZAhnbwIMUrIDS
jI488jFQsFZkLgYF4TKc0g7bUZGJT47Mauvsw37I7bsCMn9J+tepYnmJCTB1nFda
tPf+yYhXoOmkIaYMX0Vn7IHGhz0fMPvlbA+Pigm3NVWbRezk1n8Aozp3SCE/Nxf+
pUnr6WQvXP4N2mVNI8CpgvySxBhlWgfaDQ0vxv8VTzHRNhcLEzwxLodazsY1SJqR
meLKigaq9pB/ULLVaiw12iC4+6B9ryPkmixHlsRJKCF8dheo3KJR3KSs7CY5mwfH
HOCng91oi7N3GWQEwxapazR5/NVzuZNbgAqVerlJOq1tUANUIzSa6uPuEmKgg/uD
sv3rfEIz0DNIw+oE4mlM9RS34Lz6Kh2bPefRADLSv5uapGnIcfnBtwHEQCtdUad4
NFfTJDw6DVsv81gDG/x0mvd2e3gJNxebytY833GYzpXyb5Vl0kVA7/Z8RtI8F1ON
rW+HmGPkbY6hnvBPzglin1HRN8wweJVvHJIBUkjhkl1f/fa+ktQRAW2k6l+c4Xa+
W2iQ7VAFXyVFaxOdw0SIrBafAAMEJHE9dVFQ9n1stB0cOkNw3YIFgrAjL1QyrmDh
eLFfMwT81h7WYrW4FpVcwI1PX2yIaPIUbqyPU0v7RHwy+P5NFWU6CvI/1tIXsWH1
44qULtnS1ePG2hAV2WotuPGrh3u+8wbpwsYLQseUkkLZP3M8KXM4hYWDqFhZ/I1c
5Xb8e6jvC1wk3UTgqBB/p6M9TKMBsgBDGq9rv/U0JRJEEOW4FWp/Ria+nTOCC56B
aaowUTpDp2DFPaXa7IzudnfhFc48qS+SCPXIzr0zuKJAE1WM74oUSTsaZjMUw85o
Dpz48WM3qtEU4ElODImHl/wCc0l995ZdecXcPfTbYroT7TP4kM6e4SMpKWdaMq8y
+219G3HQyWACNNETLut8s60GCO4VrURr9uNfDusqRXTAxpNjctuAH2rtCpwV4ZVS
ccCuh90jOfQARbps90CFKRBhpWTZCuqCcMAFDKljLFm3yUJaoJVLg4kuqvN4FQ/U
uckSyjlWhRKQT/IkUM8oZXi0mMFGXaWOHCSHkjM7NIDM7dSozRWtRysoJS1WzcMR
BBC17QRQfC2uYOFGcjcgHkUXa1D56KXPFxpAaUZQlFN9ex1hkpLkKoIkl9g3GEbH
xVwDj3yX84wc9JHQAkIAwh2wUIor4L9A5OA8fEnLevRuKVSz01rX4Wh0EWbVYPue
7yk2CIkQO1EUxBAe2fZIdoDN6wrZPJAWkCRRBmoGjtf5Xx2PHHm4WpEOg1AM/LUO
lcLaEssouCvL/A/KyfWAvNF96j6FUa7Wd/jgRd14IeA7l5ytL/WW0bJXggb/xXH6
34gY93xbLUoQNNo9JdHw1Fs5KLn4LiUHAIWC2FnSC7dIGv4Dk6HOMiWPJaDtrd5P
Hv2IVAwMOdwoODqEFklZFdGQr9K7Ynlw4sDtkc95q3NKgXdpT1fB+i2OJ8Vv6SiA
8dnyFs29W8+Pja6yuQML6MFTmWA0yUTMHzTFjZd4Uhp47PWO4Y9dTxwj85mlNy5m
vcC3ozE27ejWio8bENXO7+Alski5niJRmJ2xfGwJgr79WmdXRo/R0YYt5NxeAKFi
DXBjmS/uOsXC9keWgB663fKcYh51ADmZspRI8WVy4wlPcKTtgc3v51Yw5/Kq7Sv5
YRTacl+K/EWio8yngRF9/32c4xMeK2PRgcxCAImDa7+NgByi/v6y+ozujGpxKa6/
hBZo/l4uCSuK27cIOfUHJIk4t7s1TBAKM62YhvO+rXsb+m+gpn/Ebfp8BRPTKySH
Vqo2FsbBy7Sa+z4Dqtwc+FeRL9RcQhAR9y4boC+kR25VREVNdL+aSKvFPWaemarv
nOY6/qQ3UIaVhKurkVRetY18AaOnTOpXm0uplaJ12Itir/SwzUwSSvl0JKmDAJGf
OvcEPlzrNguxShYUzV8A/d0r0o1ezfxZHxRA1ZvBHyb5FLe5TEP586LFUBCcpSjS
STivNiyt9nhklPmu/Zto5YOLKnX6e6JqO1RCyoRTS000GFBoSO/oq9KUJOIX9+fp
573wgeElgOHOv8cI1z/P0m0ZNkrK2pGzjSZcEDG21KvhFQ5QGgH7mhEb16RKmF/3
Ss+pFgQumz+qPtWf3NdTTufnkirr6RKSNckZHxEGp+/QGU5JtI6LGcudiuB6tl4Z
Ry+BxGfK27nYk7+UAsqWqVU/COxqY6dnQJe4RZclUWAAOXu/EMcXV6h01PaI8xRA
AWQYYURBkxQZVEKmqxQnwlETnpG1itwUwre0iKCY9By13KCmmTWRLtHPbcWB38tc
9W4HjopPooxX0W1hcw5a1hQF6IO78aB+yJefYH2WI00X4hkF835HPbuqBxtqfXeb
i9PrVFnjc1h8zELNw6RRSIm8jXwOEhe4JFtUTolvqSJFFijDePj4Vs4Fug268obW
njdrlmNkomckaEyHXrPswa9D4mzUyX2sM40zmZxOJSjW6GHbjdHkiuxrzjry3/6q
2cntywasA9j1/gGIarplCsoV2wb2PQhKVr3SIG53qXL8DNmNKuGBVI/YGea9n9s1
1FfMknlEvCAo/P3dgjZDXOYxLFozlwEE50YzYp97wKgQ2u9hd9HcL04VcMfOG8e1
1zSUlDGxoBt7bEpBT8nexbwfNFR9uAuVbMuzYhe5BfduRyr+Z47kmJg+JnzJItPr
HHCSGnyuIUTZ6NYQOt2QVOTU6hOHSVU44+LK+ipNoxOnG79S9Jdb8q7JmII338rV
Ls18B3mDmJ/1C9GX0jRNWCZCTAj1bl+0r9VJ40GB56Lx/U89o0ioQcs3xNwAbRi7
qoSVEJzOf4hhPzomJyTtrs+BmS3vYDprze9KMiTfZQhs7qBbbLLs2youu3OIaVok
m/5DdFDCWqDrTV3lzPsbZpaILIqbWZuSq866pv+33SruhGtinnlLqc2eLS5DGa6m
Hb3qjKmCmKfgLd5wPpqWSH/2b+ZgYqxHE/Hj9UmkWnzBZfqXRy0xAiKPjCFnaXB5
BCKJCCzhfpBxWfyasN+LymByE+PjFg31xvL2LGR20AFNY9JMAb55qzaDePmFaGKc
LcISxPthLSnIl3f/l3ojOL4P5SiP1murJTjf0v5oQU8IgN/l3uK2nr7VxxOwwfYr
++C4rRt5tLQqQke00pz675pfkrSscj/0c5pnkHPadAMJIPmgcNZtni+aYn4RCh3q
6UuJLI1vXobdOeIWU7hx8m7b0EfhKVmKxmeDHKI2EU54F73L3EPRtYJETpzPavX3
7GCbGnDmVA13OQdCted9EekJryDano01u3peZ3yhUrlThuHY3QLKtNT2PoWX16og
LyH5pxQEmU6B+VBB8Ch9A+vImco+6Iylaq8gm61/lyZMBZrre3Smjgxuy+p8Lw6u
gxpPpRFm+RdJ2eT3v1BmgmjKPLYmnmoZlnReo6xGNP742JHn06gVTnEQItPaZH1G
VdrDevlEwfMJ7Bn4Gggu4Sni8wMrEXGpHsj7oym8ql5JCryJmfFXZJJBCGN3Ad3J
/1HKG/8l4CXgst0PXuasOkJvt0/4d9rFW9a1M16D6BZG89m+JUVRhV2UmSKeBXNb
V4at3K5BxpTBkQIalhYo3uy39eCw39H+WX6Njg3M/icFgNZPMu0mIGL22KZbQzEz
KEds/tOhaUjW3Z5ecddQEYU1p7Nw8PDJWJ/fChKK6zj1hIOT+bkXxJNXinvKHXib
JDifAaOELTx8SXBttBW6K9vrHzHWv9ywznQySkvNNHSEfTUv2ZU83Y/ME7ittOJA
OfQr4cMuzZDNKT2l0mFgd8L4PmpxragthU+W4viH2CEwTkMU1nswUyAeOluYt/gC
f/qDrOIgiLlsvGY0mPn9Y6y6PU1RR3bTkKBFCPzAmXbFlMiXAaTdX4rBm7c97Iqv
26tRu1Sf+3zFTBTJ/HwYMMVvgXy29+ks5ZUAw01b8LPB0YlALb7pVLgVjj2PrLbK
geLnYbyGzIcnUytgtBnwDyRb3q9X+5nMYfVbujKxdEAyWFfJMaM3qWmDDvCX74X4
FbjZLZWNd2wFuu/imV3UoS2pdn7mStfWaWNGUo7cuWx7/kEy4e1vBA8FIxsaN4AV
KXx9CY5IbO9dvaWzZiJU+aSKQiM5WfHwreL6nmPxyl8lf8VHYshnDnzm9ncyvcR+
TV+fvCdBty6y2cQVwHmw1kzcYHOKsEaeR2p+YFdIH3RvPI6hfTXteQvDoPXjSugD
cenKtlCMj4HoQ7+WfFnlpH9fSwxxU7VNkr2GCPGUxN/ZUTpErx0DrfLmgM9lDLWu
xnQyFikeTrW9UiJEvufb6uRUOBFRtzq+N7fPfnGnmG8VdQMJHC6EEg9p/W0f/ixP
xj2UtOploFtWPIoL/sC4iyPqBiN/bPVFKMjevERtuZK3PEciR0ejhRqCFBezjBEa
IXard+oxTb04r8X8netDXgqjuoumkAyAGhQPAML0LlG+N67/6qIora9gZ9Xt+YAf
nl69cpLL91NS/HCZy7U4VAWdwi1mYunqtz0uJYIlm8krpRfqUziLh1G7ZTKJARX1
juAbC5gKDIpvNxjcVByo17x996XJIW9EideI36PuWNTb//eSADT0sCZArw1b2NK8
Wq3Qjl/XzANdQvB2t7v67LX8R6xWF1TYLpwZ6OvhrwUzyIoM9FefcWHlKONbaq2a
I8tmoAv6lRjtCTW9Q9Eb+tQRxnTNcxb3LMcddFy6XuPsx1FJby+EpsujcQZvkIJi
W1xXbkSDHdcYPH6f9dQNwrAxD2G8EA1FApM+NpZzrm2tl8ON/btEVMHbIPJX+aT3
0R6z0xptOG5q/8Hjxz0VF5mz/8R7b7y65o/KKCztKziACF+rEkm47gw7mPJ6fQz3
VuM1sDNHlH1MftBnVTtgLHC8dz5GRTbLTEb3KMCIxlDNy5YlQ041Bu0epmooEVdZ
/uHuyI//eNgmmrj3OMX6on0KOKUvUOzLclAxKvYK6ARNktUOAHNC0KyvCxAUxJrF
U2tl5QZRvbzdL3XBTSWC1EQ9qN0hJAYU6ONnAdnuTvJ1tohyuM4iyG9sxK+ZEKZd
2rX7WgqoGqinBXteGEEmqsIrSiUpCsJ0+jUzrfMJuhEaOn+vbTfLIH0JF0/yPnw4
k4InGAtoK/DR9ND1PzCwtoGqMe7TVR/2dz8awBpkD4rb1VDcJAj75r4AWClUMQXr
OZEpqD/b8ZJv/+pV3sz0nVNxQFfVzMe3tOhV97msWiGmWIsYKqEtIhnwiz4d7h3K
Vbd7hn27iFaVaNgmG7q1j0SjKr6e8RXtKR2fdcQDmafPwIM57ac+WuRq7RJsfV+/
Xx3fZbocxG1BKq8IS5Sm6JvDPCNU8LUkCQ3PBy5Q2MAFgOfPZnHGMMsESvWk3FSQ
2S/ktj5AYGOCfwUj3fGttERB/zaAv3uZfdzdqFxLiJccqievFc5ZjWeeJor6r+7X
rfdp5s708Em49iSs24qDJsxp8QyKCaVF67e5OnOM3u+kcuz7oDAZWkTkAIHue4GE
EZc5SD3UUS6vPHE+NJZg8pEQKJEcUO7p5jwBNUKYQ1ltJUkmuLtJ56bumVMrdX1J
TjfiotewyVShz+vZGc4pJ0/MgcQ80kUrbrgJqa0ekHDNFbHVtH30369MB8gnUWmW
PjVIlQrld69XX6215X86feE25s2kZSbiNSeXcMYfRw99kxLlO4PDFM60+icVWHCI
PV9HMEEpJJMmst4IPGUkLt1qprrFYFIHg7Jt0vNb3ZNnEb6c/hMGFBXR5nSKOAeO
2Doef3VjJdrOPZwljjmi3LtmpbvwFY09aBqyGUBdk+zwhnavW5XYyq144GAsm/cT
fadCgGq5kbRCtvbTsXt3iIFcDIaRiM2w+0GDdo6h2OKclgZTGIDdSg5BySjLBa76
pADAAZyaKL3i0mv2W2YNubyPL/4j/V3NCF6Ly+/shBLJsVA2g1lZljKJIZnArgIZ
NuvAaKC1iNOY2+/7+iHOFuaO9u3xYeYE0yPkcGGKgRoblmdlPU5BaxhRUkXxmYyA
lGFsRkN2qwx2GkzfnbQft5pzWFhzQuPtQ+Horwgs1NDKsct6hL/EtasS8g/ZPoSS
wMZ+wWhn4AA7VPVasBP1uUuPc+E42RBsLGCOz8uZCG5qNvRJcm+PMK52HykZe0KR
2KoEm+9cbZP1ezKoh+jgc7GaTX6GtacylvRK+sFeI55/tMli0d7gmhSe1Okcg31e
pSpHqlaR1jt8Lwuz/RARgx8PBdQrGcu9DronbqpxFiplNca4yCxa/txp8bwoPNZO
CcpnfPxqi7OVdq/4yvU/lM8d7rupiWOL2e0a14gRaBE2hQnsOZSVlH3+yxceUQOG
Gpt9GyXhjNproq9rX6JClMVc9os2f5eFS3EdKrzGfwK7uFX86YL+Nzq7EP9XIyP9
tzDqpTcCWydEXaMUFvBBD1tneer7IiMiJ1PDsbbZEBuUPMYyfWEGvzyuU57nAUqg
QBqf44cKGSwcdcK5lyp3UcilZKTBSNk9yf7uYsLLabJjSgHEW0J0WV7cwslICY5h
d3VHH2iiuNJE1Iuv4OxWcF+CNafCy3Q8a6jHh4c06mTaR44azH7cqZ6OXbEHt3BD
Kst2oiJkW1MGFEWbLDkzgMk8SDJyn4xsPbdR0g5zYqfj2RbhgVdHljTYdZcUhY5P
SZqjh1bOkWa5/JvPhKrQnVPCO9hcHHv5Tv3N6vXq19olccU+6iwm7tzTa3j1yUNt
1G8eZK/279TxU6hPhbvvW+8TCEC/ZsXhgrGt5aRfaIDojkg3ghie0bG2xdCbwyoa
kUIm0o7ZIYjEl5ubrxueUfp0qLewBoDMPezNXoIVF/1nKUOizkW8aq74rm6CT3Yw
7JBRT4XXzjaMwFvJz22PUpkvoS9/Mz/8hQyim2M3NLq/lKz/egL6qZzYK9fkfbnE
zgPuD97jn+ykxY/NXReXl0PVwo45JlcjpC3hlSwgwxz0hOBZZdbrqLkjXBKXC+fr
Ws1VCktbZ0V8XDgyUEacppiH5bKe8G0YJUPxeoEuFQm7THZlsZFdnL45MxwMN042
YU8Xd2cBMV5nxD4juhc9HNGDt+JuVeYVBhpGbU9OosUdh0jujSg1Ndo51xnH8/Vn
l3eAlhUqJABlpKvX/mqVOdhzLX6P+/eo1kmX6rVrFpkcQI6uhM+2mFGMlz1+CfXB
9NRz16QZXnFuiTFcqeIKhQBM2GOyE4eLFZIjCNUnwlmz6I/dx3EQMFIxVGdyQsnf
AqYcJ2Ed9aCh+p5rZUAPwPjXZFAFD+8PJWGlBClA1RsrAvylO6f76robqT1eIAFM
26clQeQUURZg41T0Tv9SahZfRZVl6KTGbbTQObvYvLiLzjag3RQrIKRcRd47WJYB
NP1y7EYftQqkVXlCQ27Xn86bb3vmIL68MR2lz8cyNYrvK1LduMSpGJ1ARZHqywvx
iCt+7wOXpzsdpIGszY2fT+tmsxhhf9hT7OPTNEkjiGxC7xUj1KpJTe4hDN3gS+P1
hGJFyCI4Y7Ra/Nc67QTMmCgfjKMHFwYZvnar16JODEGWHC6iRj+FO7HUTVIFfg2D
AFY5RJW3n/NAE/SCqREUj0mgy+ZZ9tAW7CdrivRpfdIVAGcVcJnoj2uALYu+WnZL
TmYuFx/V7VjbMrbryKDZzJixCa8yljy+NrDj0BWxEnM86L+8lIcjLaNMAoW0vlYj
F6IrKHzFB4ncIyHMHfV1iopCCC05lA90HT8c4L6xOMesUT1SsOaOsxgKxds/qr7z
gT9yT7MNyK73h2Xxwjq9oQ07Le45AeTuKX86YdI1q8n7nc4hbyU177dSxrBQpMgv
jG6v8DoiA1xX1rgoMIz+cEdeDyHbCDJb5IQ8WHJ86Mt2T7r7kuFrF+OE6F2Z4+iF
4h78e6Vi8qk5npKrzzQq2zarHLaSWljkNnJiI8QDnjiC75VY5szHdUZ1veHJLczd
GznLigSHbUUgN2SalozBKtZQe+MvNyHlA82c+ztNjtUMM59ROuE6Lu7RID9y+K5p
k1WpxAE6T4DTwkJcpNpdOGlranIwRuoSwc+lOWLSZABfsl+BVolaoise9SbDQ2eL
Wre6xorPoC+IZe8/oD5lG6HYTinXfdc4ybjGzxLp542OPDiWFBebhYRWMkcYfpLG
+1b6bmaE4VdJ4gTgJEPstgXGpLJNexjO5WnZeqdWSMxl2lNgQpwVXeUDkhSou7mr
ptYv00TI8bMqtBdyS07wvHqhCg/IIB8y+PTgYgJPXL/7YqlduFErC21/a3VXmxRc
64uqcCjQWyWrChSGjFhM3xxJMAUPLPBpDSbj3DNjhajg6S6heJ+dZ0ChqukVejFe
/z+RixlKOIAi8XayykU6KrxrJGCeFF0+sasxNZhBm6um0aeN/BW3dCzmnYBQwwb1
bQtXPKI+Gbppe1u64JEdIiOxR4gLqxvWih4FFUXFuhFthnZY3XW50OwHhmEH6dPU
g/afImx4GD0n4LEaCsd/SeLYcSj+vrwnsbZ4MlGo8n9ZmRbmiemSaYG6dS4l4LQL
BmZddjg/nR+7Ku4YwwiuzE7KMZ9aJqLsOdOu1pWGIJdTZps5BLk/zcbs1atNoAKk
gMLK+1uVsU2nh7dtR+Qb+Y9V97floxpxl8UytEwgMe997NoeYM3mpeVEg1tA0P0y
rfRZDQMbPlRUHBD8+l9frvTH1Y0aBUEKwEtjg3kB8vqu2LqEcOC6xFIN+IOZc+Lp
2Zkq7JIzUpuNXcseBrhND2adNe+dDoqBdxAaW2hbDDQdEOkzv/7vwbw1+ONCB6VQ
27CtSVtZRAPiLhn98M3zF6E37MhSFKOjVxKueD0scJyxwX75BSotKiJEpXA1n3Ik
zJvfqNf2wfm3MfLTWEF7z5mBWPLBbA2b2My8jyHxm4SHWOML6hvp8fu706pTMIk9
wGCRxlrxZt+4aduWctnbvJwRxjjbrQKHX8fn454oKnRHhmcMnfZtaoN7UUtoHSBn
AWDb+yPT+yV2WsYSTaoCUuH4zqCPyIkBfpyUOSxWVbgfHSkA8iCjRmnRrW+Fo3t2
KLOTVX1gMpt/5G2SdZXkgukisZb8thZzKdC9FlJu870L5NaYhmj91wv7SCCvToVV
dzEINM2MngqDbOIxgv30nB+B8V9gkHPo0h9ipWJs7TonXQy6yChtpw5npv4/W356
0Meq7ZrE9bwzeDvg3y4sLASHocOFkNz3DJOXopRo+9OmTmQ2U7810Cb2Ch/7YWLw
GaCtYvW1ZxX58XcDkGbYMjuX6usZ7XOhgDuBBUaMUuM+HoNVe9Fru/oDSGb7td68
FhiXz1TU9U6+4k3Ycp6UzGxhBdTrLwNKLpw9FdJgioshFtqai7SO/8Qfq1ZDF5K8
ypgV2hi/AwpcQ2w1ae5gxaxJWdbBOjd6oSqw/Tb5QLjuxHBddplFJDOM6kv+7LM2
WGWFpEel3BKpjq8s2F7wHQNIoEJ98VRrjrxOX243uyGNTpGwDRhR65n/hLP/dsRe
JNMdVr4seXbk7xxVjjqW8S6Mnv6oaJxWogB9/BrWtAuHVvF64nbXen/LaGfyxxGq
P1KuNEI1Kd62Aq4Qkr0RGZfHc2xvTJ0CPSW8z8mPTBkinPkda/yz99/c3WmsUexB
2hOpRhiI73nAcSUkshCwaVSwFqkUvIxCF9HGISbDh+3FzCfxli9aPQXiRAqtWzgY
EqF9PWg8M+iYfNkfkf7WXcGfIpye+p8ASQoMXz7C8KW7vnuRo5T6qDfvGkIJ3qhf
xHq0gyf9AqTsG3iNNi1/o4lHjLtj3hB6fpc8Jio6Z3xPz5Q7/kZUR6ay3hUEAFhK
zAHVveO0ei7acNA2O7EP/oLIh3xgfkCxn6xrFiZj9VCalEt809YVTQBfSnFGx6WX
fhCCAPxkWh9rUAbE5yfBZnYApFo5EVbYAtUAhTHZFBhZKCtllMEowE4m5UWIRR7X
8dltcAWz3rW9XOhL9HPAkHGE5VkJafOkFFWykb+7oSKtE8AqwhAQ5mOLq2VcNBhg
BKnOHlXxhhHIYHwnTw9fGE6pIrjWnpN5d+2tffOH4GXtiE19ZbWAqk8auZLjvdyD
wLdbnPrNKLSBmKMe8KVDFJilL/bmWEs7reAGmfzKzTaRlUsHhcS9Ax4x85gwQmMT
VHKLMd27z2evSrX5SbATubpn1cRH2pMQxgHg0viPXy/Ylh7gfaKoo7okB+ZPlcti
fjsvVHCDtDnE0tlkJ7NfN6g3PWcVNcw9foyQxhY8Y5rhBn3StukoRQoxTB5HAWkW
V/cmSvbFgmRK4ONe9r3xxfiwZvFuyLv7+olvFuUFN9jDgbYipmsipwelIMwNGnJM
LhXBhyo2ydQoVyJa//a/Ledlh7Wg2Cet8eLMpuRnPaB76iPtFnWOF0avZt3iEKO0
yaw76MFS8+4Fh1JZNdFJymADZ2oDvXV9zNEt3y6LvfdTw/WYWlMvgqj7brh38hhD
YMhZ2aCwqDTuc8dmWr+Y9WzPUvKs7GLEQbs7GNFIktCd4Rlmr+5JdydhWkoq8A7y
HdbIkTOUuD3Ar1F85ZFVaLo1TlmOlawPFYBxZFoyIApMf2lt16dFaNodRKoLuh/t
5NS6Ca0uGmeWy9rkH4Eqbtc+nFfnNJHEbMZR6gHSO0+b+x7CTRCaS9n9D/BDF4lX
pfgq2kOJUVmjbsRdcL+JQyBl0pJwVFE0oDmcGdy0d3GC90AgK8GPW41rh4pYnPhb
VSILWAnhsrOA0+1JUMO7zSxjezW3mvOOmMhq1pcAVWR7Xuq0HUzSLkYy92eGONZP
fXWXoQ4cRcKDLfi72v1nJlQems2vlVXhnHpdHz6vrWa+EOgM9N+e7piKS1X6CnoO
DIW0d9Rb9CzD92AJmaadiqFjgjIPtBjBBXjVDT2AMsk6lwd1olG2Jh/VTqO0e8oA
a4bKsCJk819cKE3tDOGShHJqjtUaPbJWw3DNDgfJW85GaaP1B/ghL5AsVl+XqXVN
NmIawRiAl7gjBzO6qcbQy99N38xF/+AgFbM3FZxhby45skNd9GEghDtIc2A503m0
mX0Fja3VcJ/XoydBKsVcrH1eZHJYNxuLDnwv4jCxSKmJDFKh08F2uGbYrBKSyB2h
AHSgmm3YPe4RqRqBRoIMop6/e5bmdt8QdJI9qH8WSCPKsVLt1rkZsnkU9Qtb7RDv
+oYSa9EXl7fh9mTU++cAgPtbGI0mSQAZiqaQihTZqXMDOSbEpm1WYElAlN+eqdpD
c3538xa7JGJ4aTkEBHugkK7ajHZVczuBceJSdyDDzCUzumpBJtYGyDGc9BjzXURl
ed/LbPubbmkqmFvOx+vftFtzlA/UTYx4+3B+BE5LLsOIA7upIKbPwTHEje6OtNBP
sw2cKE0siQSEApAmmUNvK9Qjq0J/k8L9/s75SX2nVJvJLI6mx8lTVwihWlV7ZqLg
r3l8htWaj8i4t5qTiyp2StxcFFbeSgc1qkFJfPgv81lse02bSpdW4Khbl9renoy1
B0fbYqmJSKeOHujOTZSN+UVfOrBbsMTp1ruJUR7MmQOMNeXgkn93pSdmowRUM5wG
SFymRfe2xyyYye667Pom2wgr0A35PX7CUVDIIUzK0B2dyC1OduUjz30ks87cWVly
8NPsPaltUhOHB0W2wLT7o8CxHDHPIN9+Q6ue+NKdGJkhzpjoDdpiom8NWxds+KiL
/QBcanGnwCzUiMgZGp9evu3biYwwnLTU19CV5KdhOemMK9ZuFv8mneKdLcjZJzD6
YWBiB65XPlJPJHfv31xQEvDpxmIQosWdCiRq54QDpDrHn9FfB6LXw/1zzIwRvsAc
JNROcRoPsueAThGNYkf/0iI7DgyOwLvWpztmLDA7Vf1RLnZLxPGN7bLNAtWiDrh+
Uc43z8wvf1/t14AHOBjZdmsDRpZD1mwRvy//bdo4SRonY4hcwDR5Qb91FhR1HQp9
jy3krAPwpV7rtjWHvG5fwtjqK15cC1JIKMnFwJyalnBvY2C7vZtOd8jJiBCywJY3
paIRKQSjn7Cms8Q7EJbtVsYk5hP1EP02srJlyXMw+yczhLPYTqBbB0yhXXPeeuUQ
wRhJTJcrGQcAPty9S++FHgIlyJ/wqs3lZlQHkbJ88Ym68iNWrmzItJ36Qh3O+RAM
0hVy2CtAMX0QItSlR5r5+4SE2UUoqkKym+K5QNhd1XLnlOl0ZgZ1PcHx4JdrNiVI
VBEF5QknLlpsR6Fz+8nkv4PMuUPWhNXSVTeNa7xAvUfjJ9tsYL9NIg3vxVa6cjnK
UD0QZW07XxjDY699iK2ociIj0/pNZGBpEIiBEc/tN0RfvJ66xz83/BdIBLnZfu5A
SJoXlUUFuyZTEnnVu0GmHw3hgL3S2X/58XUMvXNG6erMyCUGvtjaVtOkPr6EljrX
k1RJbtuIMhgG3EGGEvXGv1mI+ErJeySPyZTl2soohzkoYeVbHy1OquBhOH2aLXY3
7sKy+s4cvwao31/5vPwaZhiaz85cdkrSoKFsw8887Lq6NrVkwx8wkyMO0xTqi7Pd
KLZ7xP4MJQKnnNSKugqc21t+xvU1Vf30fUBAz5uHsL3/0HdEcIG4m0c8Bz5AlQ4L
K/ZFEPPy/5O6/TURvbGRQqHnBRL45CsGRfd6cDkApOFHCNZEy6v9Pe6Yal6w1SzX
BX73KO6nSqb9FvUikRibIMY8km+QShWf/h0bX3JuLthV8BzMgtCZVJ4Ut04evli6
Xzcm/XjbIPX9jCCS7xgHmEEAXBLeSiRkhst2f+/xyU3NgNHBaa+QtbXKxYC3Oy1N
9UVnkYpJwB+gH1sHtq1ZJm+Bd9JhsY8g5ClXXIIZh+P523z8lujUrwObxwSmS5Be
VnaflCrQ75MEkb2xOtJj7GEOhJ+haoT5LAr/T+u4sopw7WvbIGeVi/s4yezBDhUe
+NjbJr7LGF3f70PW90wrbIpICkDAPcpC9aVRkXiP+KzDS4yfdazo2/b3UA4j8eZx
DJnqPFP9RboezwlIM7nd68ycszDbPm51yL2bs4zrcv1esmepu7KDZ/0a5zFqPEqH
IV3yYnsIT9P3XhOAsYF+Iu6vAgPcSdpZR/Z8uGqdHbR5b3P2nqediwH214hSlXiE
BKfiVFugiyapMqK6puk7VG+2n9FHTfjtuQrswRUbCUhPXhXi/JACZyu2VYP9GYah
GH7E8ByblrYVfItWcw1IvMDyt0lsmsRkpjjfH4LxZlq9UazsqCi59HrMy59S59/7
zKUXHpsuFGILKkjDpq40H6TzVmqDqgJyAFJIQECE4UhOJkO7Wx0kJLmhp4aOhEeT
fRCeObulHU6LmmIw3oH/BD/oqslxzyTTU+XlhACivdq+0w3i07l2a0sqWdGI8zS6
BQCwzFyiNP7PAO1IoEq8JePSu94pe5EgBvnC9cT773Ik8g9+Ic1xozQcXEyl3FX3
UNUS+2xMzaXjvzyYLcEYbVr1o8gqBExVUICf8TadAwqVFpqCFocngYXK6CltMulQ
33vrCTYz2+IxP75var/mkObqn6eDBQ/Pnr60MiFQycrpDE3Qs9PPsDalcsVljL1S
k6+3D+UX3M2pAPDXHHwyrVjqy6atOXUNP45KfG9sfbU/n+tVliXPexlb8m08xi8F
HD6XwyTrUGvH5C+tDG0/QVDHSiv3l1bXngW7tu4r2NN2SLmLgHBkGqRkPXMP6E90
QPJJBC1io6vfEciGHJ3Yyex3eGtO5pnWZYGdujjTJH7VjvYF01z+QJ65bUgOMsZO
1RY2Lx710jYG35BHd325i6WAfOSn4MU6f+ciIrqyqq+hNxgj8H1lTupkNaFq8qhU
98T5gVpWsnnqkFh0WhiVuQtfrx+JQ7yCYJk51ZNJaE4wNlzhhdRlzB8BfRLATzKV
M7MxISLlI1uUB744pXVwLKnjJGzT1S517tiB+Xi7i58msT+FxQbFkLCRd0PhoQ4U
oaTeEzrCSsRC/KASYopDiI+Ivl1KL/ha9sUnwXhyrez8AG6X97HYcpfpECAcp2Xo
ljfueUUJMxHmZhnWD8a1vGfLPrvAtKKLatLXzrTtAhtMmkhZfP5oURsTLIuyscfc
MzeMwtlC3beM/B55jAQEtF/s3AqVuajzQyAjakpf/6X/CLjmFcskjDmPrb8ypdFj
KGjlW8c9jCWfVAPXEkyb4h3TrVECmuyIKzzL2X4Rl4qUcrn6Zq/S2wjpnSTLsKTE
ZiDUG5qbWjiu22PPoBQt+R7o2Cbhx/BUlDhR/Adutx00vh3sTfJYRfy3qvOeoD5l
7XUCKIUdwMTuvAnMOtwFsktzYc2KLlJcERorKw8qxprowy9ZGVwZg5T6CSpqihWv
AZJ2Y0UF4kapMSyJBndkCK9BkfwAkQXmW3npHzAY0GT+uacQaXgx678G23vRu40z
rweDxELVw2Rk2IK/qTAFcWKIqIyR1JZLWZUY2YGcnMcOabHgBWvk5qcCzvu/JKIu
jVaxFzoKdZRY+LeYL16RuCzx0LyVzwL78Qn6FyyvBfkpDsAbjwAUaiAxnrSJVYJq
w8oiBcblZElWdHgtpZZqvKIGqz2M5YQJby0FFa4KNq6Uvx4UW40OKK748hBIjF6k
lLI8HEsDMXOTimX2hHa9kRmj5nwzEw32ueOSt+mvl+Jv4GVY1vokkk9ljA2Bxyl0
h07IPRwya/dV2NHdKf7aDN3NwxGMsbbZdFWqO3As6V6or9Chw6Vx4Y5uv+7OjPsS
V1zu7ihR87dTtkwPHRW6vR4h4k+wHalrF8X/SLurb6V8c3QYUaiqNi+fIrTX/zfw
j2agJ+5GDajE8mnyfA/CjDS0rLfS4Nx2NmFGi11rR15vO6OXISoM0GYzAUcMsbZy
lSsTY9Qeas3/5ZXGoOxDL4DrpRl3qm82cezUxGNhQqJhH1Xy8g/9e0dJ75xmFQGG
1WZBX4o1MzrxozpX/O0f3in96FWCizBXA0JlQ5Lg8JtR9Gr756gh4ASE+QWpd6n6
zJTNZY9GJqiqzNUhKKb9JgD4gcv2OKslttV9CB8QN2TKuwdqCkMpdTmG4mIsZ8NX
2cm1iiR95KeJdKQ/lF5lHT2FszRgV/dvr9WdyWygFxxrJG+97aRjtMkN8o4I/WIl
iVCi2sJCN41WjRp0WfcKd6s9DGi3Gm43uE1dwrzO2+PiotXwzSm7R1UwSbXkXgIx
DvpetAMQdfcMUFhBU6BxCBDj0l1FOubkwj4VeT5DuNKrZjRbWZFXJabjlF3UUGXw
z+AWKVWgBKG49EbUZ5tMJrjqaZW+VinyS7UqFriPs3UxuEERlA/4MDQtiV6YA+I2
SCJeHdbUSl8jKMEvQYo/VlU9E8o4rfcVeS2t3rrpRvRYN/YKmb3BJ28J0X/sWsXW
QvuxAOy5WcTyGNGEPmtTFyWURWKzfhb8OZUAtReTpG6xHPZX7VVtrf2sPehiZH3s
KtnNE20egKO7Icg7vxR1iMiPPv2f+dxIt5asZ0A1ZVpJDh17MzUYTUOIcH/d4EUp
VB2tUbJv4nrbAe6pUN6RtNZPp4VVUAQpgoxL/Aim/gTtMz+GFg382mkV7JZkpow9
HzKSP7S2wVdjgAHpptsx467V01tWhqPqkhwDQX/mMsYlHophsk8i0Wg8bkTC0iLN
wU4TgwcejcMSKKVGxY9/pBxc/3HBUX7OsVQAx1iyA0X58CbqUoEHJikhpZDIalue
WY36Ssc9RAJXEVZ0eNxk0vXgN3Rd5etKxqTouKaP9wmkt0o2Baw7IRDC8srO0Q3j
ubH1q3M79uLGnzshQ7YakkApCl469+VQXXPEetJySO696/9AnEJGnXZcC3ySQcRv
oatJfNIcnD6RykZIXAgwsqbgaHNyxBcgXCFJfx/x1toQ5pDdht2kgYsq+C098Xza
OH9eZgI5kCqNg5EumLNeMCSCY1pzVpHvTmiwK0L3kdWGruYmT9tnPc1UcHsH5r+b
q/Lbpm/Fc1dLg+t5p2l2veUaDlVsp8j61eTXwGooU1IwYzzCK0VDPGisSmbTdZJj
N4BzbqSjVwtZ4Ks0AXIpSDQD/V9U0NFn4Inqd4+/dQBpoQcrKbtUaAKmqI8atPMY
y4FEdLu42RalMHKBSs2u48PUlbfEwXUfC4DGfoiY23K2uObN4uW/suufNOWHdiMN
PE5OR1QptDeO5ed1mR21GUZFTop0dqA7QTRLxpF+LoVMMFzFsS4h2SXQV20Ix5cB
tEPE5uijq00cxjNCgOGW8ANuojdv47zh3m6AzHb1/9CLQJzQeyqRMTKnIYZ4e+vm
eV8asUeqN3aJYJLnAY+mepcdQBi3f3k+20E83ADPEkxUvX7MEwHLHBXvEK2iV/cS
/wuHGMdIaJVczaVSFbRDjIr5owQfHzr4ssB3C843eUKZWucI1LY7a+cLeP220HYL
sa8fJl1TQupXKGTN/a6dGLbyzS1ic4yi9q2FSQY71XCesjPlQpFxmB2Dem/CXcC4
mgkA3sX0kphpAOZ/j+utlIoXUIwcbOPeTQh2g8CaXjqoSyaad49lBhuCqgDkxM4x
W8OxzVoNKp0wRG8mXNO2FZdb0OjbIg+hKHq2WtPP4j0MMQqDMEBehlntfrg0i1mI
nk/z1tCkJu+BgoAyFzo1ysQtfOWkAoYeQO473yogIUD/y85URIAtWIv0f8vY5/bb
yscZDry+AklZ7M6D6N4iNdswQL+2Q1TaS5kCi4NGYVl6hFXmz9FBQ+UIufswfR99
Aw52+C1e1OnSS+D2ELyJZdGbY/1GqyGg8MPOaM/8VMAVmwx84VhA3gV/NSoMltj4
DQ7P4ur9KSKnHjt+VKikx4pHQIBmmJXslOkSbwTSzQ+dMMaERQKjaJH3KZNWlACH
4eUDvoRpZJpcvTzYqLUFx50/kGvsReT9Txo4gf7hhlvg0KSK+0jS0kQT7Hz5fCaD
2GfWbmEw2+wxyfadRJGQW84buEI5klzKRPzPj3CBNTca48CMDfvsFrv1bpWtgNek
shZPkzcoYs16fzNuZGNVymcNSTRTnp++S+/OOjbZJqSl9Bgq5/JtoYgDg2GHxAxE
iE7In686ZD3/ofrRLJooWenVs1/4jV56Lnclm3V92t14LHS0cPvyeCQdXB3KoBGO
Hay0xsZum/tQFjNC1jy+us+bJhbXfG77ebXsyZeFimTBgK4goYN0GYKZPWcuoi9V
b6iSIBPHEe+oG5H2EckQH6gcoLjSMjldDNmvMBN8vmSDk5jHQobiYKH6PhefMSq6
qNccBcXZRRlkZ6v96TNmj8JYlqedouaYifjNpQejvcq+Gj6NIf2j5kLAwm0UKC4m
nMJwKRIZa95Tbn9HmxOZOrDVfo90s6wMopOouBYKVogNwTNW8hk5wyuyUtG1c+6e
Z3i77zu1nR1gv+veAHzwDprvTVLgX4HFjlYH5Xl4GmuNIacaOuxVsxX9y4h5Vfeu
lQjmOs8cPxUAYw5BfGUimuW+ZVvgNplTO0ACc8JooaHWd34HdDuo2dyfeAVPA9dF
eicXf3LSbZbzAqyBlObDIHnEZYIQDLc95jReNHeQoNelii9GjFtxFmtSxl11jI6Y
EWEIu7OwONOgIOZ+K6As+OmifD9Pu7zlzvJwZ6Oem2Q1wtuRVlNCDNG8HD78KGgN
7N7QAYkMel52AzCuWIR+Yox37TuG9Zoj8pnSmjKlZzqTCDQcWudAuqKRAqmJQ6us
R3S6rm1Ksb8RnIGtfY7h/+U1lsQZ1ZMhklAQkc+/slXpfjhniQb/fPume+yeP8JJ
3E8a4Th/J9YdzNYP8b7NWDolC5kS9Ul6QS8qWS1TzcKOKUIJpOXSPyW0PRwcu5U0
FswCgHgDDknlqj6zKVbfUiIQgMmHELrbucHNAa4qt8msEFoISOidTwC5sxiElzN5
oGk7uo9akK/+O8GTe8psXXp/6+MGPT+ufCuOyCRNDahFNfbbRh/cdFi7HQjlLzXr
xy7V2pJGCnRFJ2g19OVACmDj56hCSKdPDCmYjwiy5WreMCpIh1pWe64WYAWln22x
h92ZsFjbw6qDgWWovB3lDhftRrv0rnEDo0R/toA6bG0Af3RjDR+z78mSVWQVsRL6
6V061rI+WaWQICc4tcDSvcp4h+SpoNm9okUSFXidz8yYLCmr/iy578MGOBWeNF4P
6ljoxpqJjq71oOjMXvYB2yJjleOvNwCRiLt6JTIIYulErj5PVOhH+aeIBMe/FG1n
QS4O1+neHLiUZexiNtqh8MtRdeDkkTDtZI0wbtCJbAdcvqzFwYOQOKCPvDk8UaaZ
2h9oCTGtGCEKouDN0tl1qyTiv120FhO8A6HlUIrsj4gmm4+vVyFDzot7UFBWg0qT
GDN52KMHU1W64yi+oeuomZPSx8LHWIfKF3awwCKe2wrBj6/PrIZcD94wIeANez+1
HcYdy+EQsBAu7aMSb4QlyGNAhUO6hTQqoHYsHIjj5+zMZtO29a5uKlBgdYcpynF9
pCpgu8RsxiNd32bvEVO/y1fLgNapPnv4BnL5k+Qu68p3ZHBO7GbV9AkjIj+vmSca
vIzfVXGEJjjTuy5liaouAtzen4euPpKSV7jKf2/8few0Y1V2CgEbKxKLSiJeNdzo
46RkG5LHtO4q3VWM0ucuXV/Hq/bUXSzE7rv5gIe9SAyJ3xtkiYgHIgCtYRWnGjcw
eId9lU8SwqNP41vI4wZayeW1mtVb3w40H5Lan30Gq315505Phm7jJt1jVkC5wg1Y
e51c55FacIyQS/cTfENsWB8UJXhs6DlOf9Gv3aHXMnlLcwQPqac6pqOCojB/nRyM
6pPSk8NTv0C1kdreRVt+2jnMRekmGShTdVikiFgqQFZurcLyxhEIabvn0j3t9g5H
fFBIJMlFh/ckgcr0iNN/Y0bsIyX1lDY8f5V+32uDpRD5O7qwceYNwPlxp+ufMOvh
nHR4Bk/LJBsxUxMhJeeD8b7LJEIf4r3rceTn68efTyky6VJso7auIAkMFPuWom8H
ofWCFFbq+O+a89xEpyw+iYKdnhh6kkabUXzIcHDT8+QVgcPa5HD1Zq2Yic716kfc
hS0LOR571TdCWE8vfUBUigqsdR6/Ky7lhVF68qCdorLe19lxPYBXOkuUGGdRw/q6
2jeUBBMQU7d8Mi7W8+IVNk8kJHFHaI41fO9KclASreyT+6cIzRpe6svsE7bKCEhs
glGV79AZ0iyi56Pm9dWLyrR0WX1ytkeqgYNOODE7VP7c7Q2Xq1DdV6htPDBprQbS
5gOaoG6NOJ5SMvp6Y5P0DutgMxWW2Os3cPlR7j9q4y598/97jVMdVETWK5nhK9rL
FN4rP5NRHjtvhXUYNAtHG6eLjWTsrz2wftrOWMv01p+LunazLHFUOB9HdbgiD/dp
fqBBUBLdaxOj9ObAvIiZEWveD3MqvU3e9FjXG36WyzkobWFPoX1nmbAkQWVVemtC
KjPD/8yWhB+7F/q6iiooRvatrfmMZH5pSF8it4xFoT/R0pFr4WMfXBEXPutmeo10
Z3TUyEP3ccg40hwbtgE2YO70jmI5VbNiBulH3cS5vc7wvm4yVr84DTZLzs7GQFEJ
IgTYfzxdxEk0u4E2QxOEXSG2uGdjAykYaPkbtETWsQzxaMNbiZIOOKFpa9k6FoZ1
f1qIlgiWmgXrFrTOpN+tr2M9SqkLxiTkb1es/SnhNlbSSwWDPDBJ08PHsThEt2C3
yq8jUyV1qUKlqLQIchOxbs76ITNAttHD64kCHlphxiFaqAIlr8dqq8vXcL/NJvRg
22l8AFYTIfSDnt0Gxv2cBusk/gkONNh87mfJi3I/wbJ2cBHmNQ5wRSICzCWkNj+A
aUfBlCGg6c7hjfLO5tlxkWOf40CFCvM6He0C+n+ozhr6f35RoUTXY0K71DM5kAg9
hQGU5jNs0PJWRQf+CcnAEM7nyEVG35BnI3L+MzMtSYLGp4tOORayKJHQoSAWfQB1
ZA+iIasaAIMy0G29OGm8tMEW8yA8vndMhe066MOSYtv4jEll9LpZVoup09SbFwjJ
NLzy+aC7Cjm2PJ+QEexHP7vs3SljSuzAH+HRLRRBthWcnI6oisoJJp6gwUT1BHvF
huG7a2YwoyWChUzPPlBP/kbsYRxr7eKoLFGGW/kCj/bAwSNRod1wH5w4C4g9xWAw
nR0ybTI8vYxv75hltvjoiHcHSpLtHwTSrd7Vd6l+nuNUvJfRxHUrkcArTJ4pZe5i
pzXIC7G0LxLoVYgECZz1i+9wPD1jIiffl01RpQz+dL6aj1V+2puj+xjb2d0gXmM2
LmVBJO2XDwGtgu1D4RfI47n0j8KetoHcAtC3H2CGZ+RmxOnlIhzHDaTxsqAu80n1
D3ZBUV483YrAgwLlkYY9NeOPgMktqaIeSM2TbzE2Orry37fNuFPX9EgjfgvzIvf5
0DImXLKUPgpVYXZ8FATjDbcaDuhhAtGvGJWFvvwb2pOropH6E0lLlYTHtL8Z0zzq
WqyCeU/zspcy9wr2UzAFu/58PHVORqUZofMbw2xOERKVj4O01dO2UOvFMjvO91wI
RfPih9BWLwbuM+ReVoYtfORRqnJWe8Tjdig5Q+wMbO1il6BpyqtRotJ/gI8o2XUj
3QThANQ/xfa4YKc2wZWXuMgmM+cotuA4s9SM/QpjBvnNka3hM3eXRCu1ChpsiAQd
wNCdpcRS5nII5S0MjHmuAOeyGA53x8p0RINBVsLNMrkoQBdMc3K5ARKDnHxpk/Vp
COITlZAsww3s4Vb3dgb/pv2ZNGEZopRMmqUsgrKJGXaFvA3zVqXf4l4fMKVZ8zCc
a5RidJ2eVC61Xx2uwQQ7ds51Xz4lPi02OL90R/HVjolduOeLMtcA/ft6w36x84R7
EsB+lrVQPvhSFhr9tLRCJPnI6UOuK1IundKiH3v4Rvgyu049caSkZbiVbI3wO3Sm
Vh2wOGe60uCaX80IniRfiOtXyn4468l5sStxLQ1uiKpCRiQVrGzSRReQYZwQiBHl
nSXBtA/4zmDGIu7+8KescATdASjFVWsOKC+vFjLJeKYk5r/UzmB0pi9Mhl5lu7Pm
bWjSVk/oYeLQkorMLCrFExZkKnpwg5TUL0Ty3omexes17kdUNuroeA0DuWGNdGFM
v+/dK3xaLRpGNCKRNshLc6WE4eIiqPSLdpmKUvC5YoSnPt0jzxM7TotEVpkMrJef
/MlWmlKNWxv2LCZAsAvfi17EpT/Ur1FrF7upi/eQRWOeYReJxoem2fTuxty+wgaG
5d5JAZ6heemxn4Va499YLrj8dAhQg1ysPSQmqUuJKZwCfdEGMUdz917oZJJnBXYk
dhXGFb5QLiz0URmUPT3fQplVEdY7oX+ZrCjXr13UoSMXrgnUK4f9uMxPgzg+Vbrg
3j8n3aNWw8ugKc0UWCmjyHttGqdzEf2U0B2HNa1ZcYXV38MfRqKY7jJebdrwpL/4
PwxJ78fQhL3R2UXbcvbVME9iMP3kgkLR1CBoHSDXgoh8xofHX3mgid9JV0PgEoZL
TFgbe9dkr0n8I2UxpdWRMaNkqJIBAXoT+8cCJQ1sAx13mR6aVlLOE2b/VWncQxxt
YZa+8QxCoSXOSqRvM2exn7R2lL2/fg1AcwmZlrugsVt7dkYzEmtsYNUm4+hKV8v6
myrPR+ns7WzkXFQQE6oDGi7Gp/0/rIcbOTnHQdscbTlXSXBJJjRanTTjshucKz+3
mRPPZ8TxIby7qIo3At9ifNMHI5ONLxe5M4Xzcmtp9MPjQSL020r8B9hrOHGToAfv
P+Cb5B7F1Rwkqa6nTUc6uz34sLE6iO/PHjVdgNfwgrQht3X1z4e8aj2EWwPgYBD6
6lYJDEuC1oSzK5c4lDTK/y+XV8ZJr1c5EB/49MvKOUgnljiw3ivSPJMw4/O+/IDP
idrXAOi0nLd7mgRAZoIoSeDtLAg7pLTgzHSBjYRak0YmLWYbg/MPZCj8qVjCCmSx
eOahnyzww2ZKA/6K//4G36KTGorPqTWyRJZcjuU2bR6G/jzrnlKjcFFw7y9nf9ae
JJPb3gmQLB1ISsn0JfZvVAhtixUejeM54clo4B4Uy4EhVz0wzOM6jDYBxXYzJleX
9XQAKWXuaTr6GeGq+R1YfC2xb2nG/LkxfZR063LulU9Pb4Mgt4z/rfLyoEb/rumN
9z+DEeAwdvaZ7dX3DN08YRoPs2GGIQJS+P8zYMGEfyQvPwFXuBnH4q20wpcA1wgn
YzsbfG/fSljz6ptogr7dVUSbQR4430te2safrmHh/hVVAsGpsTT+/YiHdZWRVdFt
x/1jr1Cf4baZHp68ihWa+itSMYHzrrXblHWLSg95tXm3BeAipMrvgQ51rdaURxcP
hWjB4AuahNuSwq01g0iUjQ4Y2dtzDW8ia18061iNKKTnEq7LxWRCCFjIMR52n46O
qWXkPodDPGcawTR1FFJLX735j40VgBmgU6BDQ/met1uf2802ElLzIhnQ9r3ztau6
J6ovT+9o/tvhn8MnX9AElG49A5or50HCNvzahBqpzjtR+P9nlTAhwDbSLipZLDbc
KGAzsyxRtQbgj3HpI34o0uFvgeoEjkYcJHYui6ulNW2FAfw35l37Uh026ve3kNL6
AXs4t005Euid6MJmGAv9cUEneYWfjfLgkOZimkHKqKPhuQlwk7fHZV//J7uTnU4M
OJQebw8oZWGnnxjXJjSESEk9wxWeln/DGQn+aX96h4FM3TEqaUVjW4kCBFMPoPa9
rHp2WC17pzOVaaB3y6zs3rBFyJR/u3voh3F23axXRhUytdtKYRCYxnrBEAlzmOGg
/yU1e4YUp5dM6bPEXhSqUl+WtiYTnd0UV+M0hos9F/+Sq9mb8PvsFSfCFSQPT+3X
cdv8KPmsrbbFUZZ0OI5c7SlTujkq5Tfwu2VNa1T0HrIALmvLOzx9xY1dgwmINd9e
n2ac69+F/4AVC1MzRZqaz9q9f0eoscSZw/v2BnWv9/R7JFwBp9bkHoROVjFTD1xa
LKhPm8zmcdJbCRysGnWO5Nq+iTi5975MueCn4uQxb1sCs7KNB1qkLfn8GizTpsef
Gl3/gUkdIZH/Uqr4W/HnV5bsY5jRCXWXhX0AK27wh9fpRNiJNE8QlZd058c34M9n
R0Eoi9oD5zO5Tib1AI5f6998QwOvYu8vUUNF+1mZmRS51i2+TF5fWVA006f5BtIo
CBT2A6Hame0+TRNwSOCT/CrkwFsyziBDuacQ3cO2JPIR8oNbkmI0Aaje+Drr6Zb/
gvkB8qQq7EsNppTkSYKxxBRB6T+HBzKN/hrKgtwxEionKyR7R7cWVYE++AuOXas5
N8Ij91jaZ9HyySQvab8SZqxmO/P3XB2Lx6SnANdkmh1wHi78kefM9GuaTK/qzSPe
9K4fIQdJ3SsD0342dUdOkluawiOM+U40Un+hnp0y5kBJeLPCf90PAi9GjsavoY1E
H4+MQIbipo6odjFEM2quw8oeVBH/lh+cNLhee+ouBDowoDECQlirolVcGqY7aNd1
RdcitFhSG7DmecxjO+sUgIHNiqAWBJkrFRBk7t5+1s84chQ+uIWIOxf5YrZWso1/
7nlkEXorhLSC6YTp9v30QLLP2zP0B9Jhn8ppHWqInqfgDbEbsQVpsGxdl9bGLBv5
IHJ647CyEDkXOhNqc2fRvrm1DyE/jAwq/lVWuvOlK776je3hYU3amx6a01nshlZV
lvCXpS1ef50kZa87g5x+qPakb9Isu75vgqXRxXVCyVXaJxEEmuFqxAl1+MqEBkfK
oK+eecIEHagMPWqgTL2+idDhgEBlvekikH6/egu3zzdMx8rVE7MYLSyVM0Fiwwzt
1CWl0wvewOyrNid5UdKmpSAcA3obLp1B/JOHlJckcDIzhoerhuyfbBXzi0llzhaW
VfJH6D0FTvM77m1JyhE6Xr1ZulbKG7dSDK8ScUTPCqXEtyUgWEfDk0hAJDXzow3r
DaejBzUOTtxha+0+sBVW6CM09xz9RPWgNRdJ7kT3qDf6ApPJnynX1NOifjOKOuau
5fYBzNcr6daIwA2uCkpRwlYhx4VYZyV2EZujVXI3ch+X5+zYEcnxDoegUarkzrje
anucz6ihN4gu7hlCLu4nUDvfprz92JmWcklFNYUaEF3askBWRWQ3VgGwC0Pdx2jz
qfs9J23gsechEUUJzV9yOi+y09A3H0FzYbcHpasfG9Kd6m9CF2Bs9PVG3nPWD0sS
/YwsewrRhD7I7FuQVY0/xctWrOa6owl+yl40zDWbGQWuLpaXc3g6S874tfLZns/W
FLWlN+IDl+wvtr8+NCSfQ8XdQNET8PRi9x7JhBxGcmhCvrf0VCDScUOQJ0YzVO/0
MkBlR8P375lT8yCYm7vlKjaxYqwbql6V0pApxJVPXZrUmDWffodH86BAEqLGdS5U
EUXgRoFt3zTZO7hMCGzJnrWGeo6AZm2Y/ZeQAVPxhqP2x7lFRqeGUPtka5Y81Nxh
lTHnvkSZYFZG8ljKtdQNz6p/6qtKuYdYsTvnbya+Gd+u2ld6KfU4UDeI9ALlE460
YajuIRZVxHYdyPbvfC7MiUf0ZQyUddisBJ/Ewc0riEWkz2P3PyjQTMGUHXvio/ID
AdxWUBjfVM4SYuy2tNnt7iSI1R6wme2s6IE6U5+NZldMKRtY1hkXwn6D9lOObjUB
psRPisqzPx+OVkI+umRXFzTv11FRsf0IRDQxsg1yQmdmtvzCPueA9lR+jlOaQLVP
+6zjx6rmgXSLWSbzH9BgpVgrk6GQkbUDa5DgqYjI0J7mZC8Z35NCVvqbU6IMOzBS
HOEm86M4bZ+3/kmuLO48UtMq4N5UMGla8NQiMK5e9ggMdXn7PNetOGmQwFzvp2NB
5aigHfy1EaE4FjIWrGIj6N3SqoOVg1qvXHCX3dbzcJTdhllEU1Jzyw6RN9UPnlEe
EB6Bhf16Ii0biKmOW2LjmIdbBGDTbEIvS6bDkW7WUwgV6JJ/0TS+KNc4oGVtMqHE
FAHfbv9H2tCYMMMIVtteTGVsIEtQ9LPnPEH87vhXhf4GY+pHq25iE4Rb+6Q1kLvb
TrkLDeyJpN098opSvwv5LwOwiscnofhz9jEw5SnITcpXfGcC6PtRstYfrIbTviaa
XYDmyEfARgVcH0xlG1gpoPsyyZHfVIyxMxE7j3op44Ehd8GTXl+rUrtrClOvHOlb
/C0dWwIk53ddRjzJhIvR6679RXKFgFlUIrQfrJhhA0N20xXmqq+H2XLKWoVFPvIO
kAUOz/csrNyKTvJD3zLPj8F393nB7lOsUDRtsXLXHGmmujOr3GHH07C8HmHXhohX
Wp1pihwbPGDhAd87jFeDsICzpLB45KxSupHuUxPPmMtIRtKvU7RTJqCBZcHPoxwq
X6qizZ6VcF0y70UdIjjmrQIfs7RTD+drWww1ZKimdWp5hhMJ5jJzV6v3+p3TPG98
lx0cvhpZGy7kGYBjnWv9823B43uS1jVP+9DSiF8V7nv+5fqxbN5MWM43ttaR+dhh
vJwdF9saqN/cTN3E3307DF2+kdgu4xx/aJbKbJP8+kRDjPTwcmJlg6Ippq1CikgH
oRnbLqpiWNBjTSU1as02z6ypeFZbwaLLbBR/hflIcH4izLnKw9ssblH3xf2JXP+w
qsiBuwOEieWnltWYlzNSjU6ghivJ8xOoaaOtEj8y6+AXfhMt6brywlbjQO+xZDlS
nEbGHuOfkY3jDUeCp3yFiXzQL9zRHEED5SfSCVUbq+PUgSfEvAyjASg2tzOLs4/x
OSWBX9pInsWn8hu7Sq7BJ+SpZ5P+LNXHiaDE9t4aZP5VL4dxBJHkh8J0OwRHuykP
JbY7Wguau9SK2xCmAxaekwYeMvTvUqV3JEQfUZdR6VJxllPjLKv4uz2WYxDp1LXV
mctSIM3JfdyP14ci8jF1nvXxNsw/csnpJy7tSkGCT0D84zoV+9AiWG0xEEB/x9rC
y6ZNdnUQDumLsJc560tKGI8hgYMU89AtdCdsQddGAO7O1dyP9ljQzH3IxHqjR6Xm
R7qGTmj2XSdssQnYjSgtoCwN6zPtdpNP7f/KprFx3us69iQxRMKnHPqFzQ4QIlMK
jd3wKHD9ioMK5QQVwRn+O16cbHErEwYY1DhOejShy0BBQpSk4Yp85Q6//Ktq2bA3
7M9nJ2iHiJvRGlLWX2fwEP6UKl/BVdcdh3Z0kfrpWBRmoUzU6RywXpy7diQap5uL
NF4b0V4zIUfQuuD5vJjTSwO1rndzfv+U18VYipONsaSPkD2Unfm9Y9JcB2bZ49pN
7QBCUZ8/pCfNR2AFf3KaHF5iKXTLL094kXdUB6P7bWoBGA3uLT+D/gL7txb9JkWg
hi6JM8me3xvr286j04wGI87hJJG5CFC9lTrxzk36ja7kubttDoSJpYYKiYsq14D9
OeISPHoqLUY+HuczQeu8PdoXXzyAQf3VT667s7dwabrAhVWSm2eTNOY5NmO7sTSJ
6kRFw9k89M6SH8v6Nz9y6qaSXGnVdefwpchgLPt+X6/GWoWXMCdo+KBU2iQ+VjMX
V+LLMS+nT/nXy7ST/mSjvO85/W5KkxTYhnohD8L4pHyl5i+2ssIhN+nVhkJI1PzL
34qQlEC+oLsMPWL9W432BFi4nh88y7y/mvp+lxLW7u9qrFGV60xaI9AOx+WWbWXY
irj8Rx6E8hoSn4su33FxolnguZXKR4NBPG89cIDe19GTqRBi8chlup4dekRHLloe
sxHu1dgl6yuFV20DbIYDlMxTnzm0ZztYxhWF10cSBEZtey6pBGvIIEZrKxM792+q
ZF+33wmD7pMkPlDDU5hn35ZSnKSOEON7klRnIwxY8cQQMfc9F4D3bq7uXGWUz7z8
cCFttWSC7BLMmstqZHWU/O3x/xZkoE0ol1+frXW9L3XccOSCbwWbx2t+m97hUym/
PtSVV/o9B/iUB6QHolCLbZZGrdujnyWAWCKRJdnnbp9ZjK8c+4E5WcKcGRsfU0uU
TbVtolqOgCGdn64nVJUYEMYGYx5fjEeawWR1a1YOPHab18Y2ncdcxvWwtHWg19yN
EyqU10rbVzv1l9eGhUXbAui68TX5PSkslbqKDxeUbFpKoXahHdCSZO2N0eiZRWHM
DlmPhiiezsO0k3ikOEy2DVQRUBveHQfbth5REa1WTDhWZ5stZsfwKmWbPNxB9lkg
rai7yduK4/GX85DJ1qhtwj6l/OXwY0XC5uUZmvwmORNDSvf70BYIk+76tojX6dPw
SM6G6n/GYphqj8Nq/IqwoOmUZqxZB+KEY2uyyGurVTnq5QWhnxl7XuCdrlxm2jLI
3nCdODAg6b0zUfVmmVGg8LKZ0eEW4PKbWF+fkWQCVBs3okAM/cnVSaO16k6Qx0Cy
Z6SgSBKZ4jSChwh/CemL3pmeNZ4FgrwIuqWDSwV90+/z5kBuLFkKq8LU/G26/nGd
hsaUgqeHe0joadTWykypxdZzpBBSHWca2IyKmSPiFLYikhr4W/BT81IVWs4iNP0e
f4Im+rJP30PeEZHPenEvgAn1xUOezr6RZwoLy9nNcnzKownJk91Cdywg/WXnQiGU
IB2cAxP1ZTZ/aBkhxNCqiz4DFFYcnxTdEO0QVTfywzeHIU7Vf4pp36RXsct5DmRO
f1eXib1ni4MkcnLxw4kTRMqMm8qdWsKbX+Rk5A94ehjuhMpoZI0GXYBSWZFtwtv7
X4F1SywRiOAAuBxpiz7K74CGeVWZeyM+fFcPHYa9sWgsYD6hVhKYEtX9U1+B0gMZ
PC1rC5x78UveGFrD8L2w7dacCgceGir4sqOP5x4J1OpxWEvoecu3rtwXzydt7RQF
mkt0vnspKYMS2kIqH8H81vNLVpyackcz7+FMfXHBeUN/+dHKVuuqy1D0E+VLfOD+
2UYKukVq7y284gLxRj8A94wOmimZMBVDbACPbzHyZj0UO7gqvHJu9gTejmvjP6zj
Jff9DFEWlstmiYUHUp1xA4vFE8vcIGDSEW48z9TU01mFhiYYEfqgb7E7rsLiCbjH
31/WVQ3o6bMVM9YISjzi6FjiEogmmf3HkffzE8DRjGoV5LsG0Gmvp4oaS1frqPO/
xtG/Un0tW3GMvW/jcjyZOEeeUtZxmZHSw71R9q2FsR3I/MN0tlU8bWa+jgJik4Ql
JmWGgxIZuqferfSn7AHIYRsFfYZObhLbLw0VeQL3a482sE42rAzZmrOHLkwL/46L
2aYUS0TMO1tDr4XmH6dT/D/4+D7hqaaON0AcokuFw9faycM5CBOoEaJucxSfDjFO
9lTGHVn9sCV/Heonj2ObnAut21Ikq+A7rqPrxjI8d4UpGYIao43DFLWV4UQWsTg6
SNCzgZglstjmSpedrb7jVRneMrd/9EgG7VlH4YWMqxrEWhRmx0Z2hx3RV4H6wUbr
Nhu1DKuTptL3kmSZn2J6ZLqY3SfWNBwCcibwt8vNMykm20YBf0V9609jevqoDfId
5KAU7STrkyvGS7XBDP4El5qRKHl77pcVq37FvaeK2cASjkENnyy2dytgh6e909G0
3aiz9W4SH1RhSiPqZWQyQP2N/BxkQ6jhtWxUGck5NlU5Fi4bitjcIt0KoGhjP0UN
uFjtgZ2TSQPqGNgQ7d/M157eM7WagAwl8ldQQtuq+W/ByAi+Vf3/UZnZzjAWPN5l
+qGMRaEXMRjIKa2xrOCtqNAKwUK2iSeLQO60fyRKFY+/cCMWbUa/abjszjlDc5Lr
WoegfG9IZYV+dz30D3wUDq9y+IElJJmkY+DLZmtsZyGzPfRpya3rR35pBP3lF+u2
bDE3Gv0lts9VXw5k1UPRGBddBQXTP9/7EfKRtRqqMg/1M88JoW8dEAT2BdqN2WRp
zMz1+6rOSodxXxzidRY/TC2bzbzb84hKW+eASqjXEBygxBSaWR68+kQlHpsunSqh
rLkSpGQMqIvrRwLSnm3ZaNoLfaOx/w6erVWpcDZp+rm4rjVMnzewRRpiHKbndkW+
+IQWafCVcQHsvZs80nfUeCQpDvnwjqw594D2vx24J+DYqo57VO7nGn2N5x8BZ+/d
a94rb1kkI/SjxcsB7seEYy+EN2nC3OgJUJTOZOiPUl6HbJUxv0qEAnuUn0ds3cOu
xo0+a8881DZWJXk5TI0MjnUKqnI3FT0u0CzwJF9K5DgYKfbMIpQEvdoeM4NFcjH7
oUS+wbXiH/4LnAqzo/3rNlitJ8t17PbpZL5/4Is/icaf527ULznLRKzImlhmzci6
POdd6Z8e1s+9nTpnGEQXQFsRLix1cw4dz6Qf5AakjMSeJ0DZir0RvX5U5djSSRZ7
qU4IRyGO00jKHwQxGDmR5ZBYDdcFFg3LMhK2rB0NnEShFcLdWAy+G3vKmKtHpVRK
eHmFaoQyBrIjalC6fM9MWnzrIR43f0w+vBtvf6FLmSa+o0FKec/3PFmo3vKc9FDk
0RplKnIZm3r/e+7l6rdM/Nk0mqlzlPMZx5gI3r2IGnOEN0ULxhc0qgpxApVA/dsE
uEHBNXCGg+ZST90d6acb5J4q4R46QtUWfF3ziU7cqOwKN5JsTe+2duko/rwCLlyG
rzjMwEWbVc6FWvMjJssPqkFKuzFnVLp1w0ptg5SHHpREXoSEdLhN6F/od0mLmaK+
EP7YYdTDFV3fdZqjysLSGDBQ34WaIP/ZdqhBJn7DGHXSWVtxvbT8Dp42StGC6aS9
/s5R4gKYTnKMpzCEW3jH8p4iK2Aydd6lg2kdByB/ogZd20+nCGVElg2asg11KvQN
+25QHV6RH72Iu20Hdvr2DLgEGQxjSwLziHsRifpCsNKHFQdAmJ3tCpQivriV/d0e
8uaZ2YQVvsMCcUnBe6o5gQ6ImdoEItD6POiroHW5ENen0co30mnvEk1hyF00yHYO
b+IAV2vqtbCfKQoCTe8EVzFWe+BW3G/ABb1k2oKsNAhyjOdC82XN2Zn0XCXoXXWV
VT4uGf6tT7EuQca+Sx2sgKicQKPBdS5+vWaddM/Gc5aG3bPFUOLxwFhm2tlH/E5D
WIra6Zr6nc2fIFOy9Pqe//fXR6hdnpOcowoUMrLI5TS9LgY01bL1pUsVr/NtMIUm
7/Aewo5kfnfQkgvddCQmlBTfIraeHqgip3/CSViY4GYKXEBkUqxGcgP3ivXWQcRB
mNWz27Tc0tVYybuoTxfRFs32FYAx86rnMOvcThEKFcGUPofR4Y+Mbj/LI24z/RyX
Frq4W73cO5jILhGc/MrRP/U92Wo52Z+mzxOLIqpEVxQcI6V/N4c1MDi8wbRUQJLh
nK9WxUuPq3iioa8X1DAD0AkmSTZCoSkkBMed7vSvCcMtpaeQzMPqed5av+nGkGAi
YaY+B2L1QSklDuX2MoM7ceN8ijlg22f/ysrbiP6Psxxr4AAD+nQzWyVZoM15BwQ5
QrHIEJUBKhj+Hzbv+sTafHeKLV97mLQLZ+hJprR+md9eVR15Ii4MEQ/PsuJO2OJm
5AzOMiTpD257eE65FPWQFk8MpElTR/mJvOJi8qteAACwdCiJIi4iank6DnNhcKJG
yRr3YB77cQcT1wnoxJbSxEv0KKJXS/y66iKbVAjRcKdU0rDgZ3iP73dofKXlkoBw
P3Wc4KNQ+Y7mfY2oCN8uUtihhAnyzsdVTESrbe5iwtnofJlO3Jpg3vGEMi9aaK07
vkjkZSUtwa3yHX8LHAn+YSeSH3tY66PMXkRV81sTrf9Gocv85zhwsdYB8ANVJPDw
k1SYefR+3ATf8poQKu+d8hWrLpqpe3HH0VSP9ABI0lQuVqsKJG/f8bQBi5jWp7vj
ApFV5DMMEal9D+d0kkmW4GVeqC6l+0GViXFt082DNVN3jkRj34AK0LsIMy5kcpXs
u8u+q/dNHxutl94fSnr4IVdixr8WiYxqShXThcLXlQSN/QMrxlqAUgVsuxm9CfYV
PJksljXn3ReCb0YYgdaj0A+FC43s5ZuBw463g++p3QsKoCxYqAewv4gp9z8LLAft
cM2ldT0tnuiqMnwKrI92a9QhSnRY7jzA3Dz1YUG36QMf3VEFaGuXgroaeMOCnzcO
ETdcXhYiKeBdnP8yx13me0qVUUfW2yEUUuDMkPYotYe7ZPIxPBh9AoP5aJumnYDI
2dh1i0JAPOXj6Qa21mP9C5H+bLzRlbhxCzlbS9iCJgr7uWVLDVb/oHmhiibESuAL
x69Jxm9elXUgWt1hiSEV4Y7QoYQKddRI/7tzHarY9K/Q1wjbYXAUXtxcBqgFm3oK
nZILU475kVjhizazejKwEtRFSFb3PtSvNL4g7YHXZj5U662fT07u7oYPmTWjl2oe
dBJUOwU/XtrBJ7fPGKa7RCWpIjchiyGM3n6LPeL5BXZipCFRJ/3Q5HR0jGhnNM/N
CMI3SKU2BXv2rBh5jF3+VOXA6aZvsdMKe7s45rtltHS3m0IW+n2bLCOWL09rexVr
Tu+vaZRE9Xwdk/DJ/3b2sRD9Pw16VMKbJwbxTPzenwc8cMpJT78Y3619qEZYtWWb
PVvG1BsD5DVR8dE+G53I8+FlvSLKgBkyLYpolPqRfeA6BImZD39aJQZKPouIQDuv
bwoRfsIjT+qkG5V67tDnoKYTG/Okyu3MpUwLFl5iyUsoQMI+vw5QLsLFR33LOgz1
YeIV4XYc1zdzXoPPvZ7S+VA/qW6Yu6W9FfLqAbeKcweMfYCl1upEihsFwhCJdOS4
j8bnhOrvaXGkUOMRaIMLKAk2U6Ot8U0ZB8lJk9g9f+KNn9WDryliKYczmi8CKAcz
gtKgwfDUdis+zUpzYkve03OlWbRwg0nA0xPi2unzAiz2eQXw2emZdKwXKYXeH6MB
xYIhcdvtDjIb1+ABF9yMoVgZtTRShAjfnqyyqwkUSxatCQoRPJC51kcXqIt+aKo9
WD9H1MPGE93FPwkeMcik6mVlCqlPEmjIQEqHYfiVmBdsEaa0J1iK0eCVWQ6QtV1j
HUkac59gZNzhsSXbSJTn19Bm3O9ORKwLW9aOUSYfwoModYLPlJwR2I4+NuP5fitf
/Rz5191V8TPO7p6R+/1eiVzlupE/qAgDqu3B66wreVYutWIFviKRG4WT3Lfy7P6h
QR17dftORBi30sbkg0I8uv/cnaHGgqza/WqJH58oSBkk4HC+aM6s0+gqqhGNiFLb
nFmnrD5xlQB1wsFNJQ54hQjS+9I+CSNvYI9/QSp8a8m8J0Yx7MRdpsezwENAS9U5
4C63+Wb6/zD5RXTapcWc9QFivilZ0a4YZ6KnbxblXEsfBx2uoWIsK3YB/6TUxYei
ulMZcqDpvdw5kb1UdJv12pToFfepY9uEtVtZ7b1OxJEKuH9NAUtoqB8N/RLkmvwP
wnu/psWPDqrseecpNI0B/XDWhmbpOya3SW/OWqXIDvpONzj+Tz2sZ+S/x7YXjMSy
KhDiXyWvjDcvC90toldXmNLiUnGzV31n4cw+jl/LYE/FXUhIgz3/izbKaDZM/4Nc
NeMnhJ4k2jLctAVsj7quqSPgzMA/T8MHzyZko2arPcOHoAR68W4qgQZBiC9532Ba
3uH9ETUGrrwlcykLHD3IZixO1nfNMkMfjxgNWhiXMhFoCgxnkGNmKwAFSX/t59uJ
RQbVHSRRjHQaaDI2vNeyB6aNXpl5zl+H7i8Kbf/kdzCc8pkXd2GqVy1+ClWobuRv
t6WWJzwniPOhU1uGEFLTw3lBoIwpw3esTLoIw6mT7iYO14Rt5ncfIFmR/dBhtXf8
JIyRKGpGtptgSPUbq/9/dx9k3Rm0amyyg7ny0i3cSA5nsA9rT+OAkD+8BjJNIJL2
gCaVsPtdKnPr86NXTD6vVH5tP9hPN6qy3fI3c3zMcQ2g/PA+jG/npTHLTdr7IlaI
RGKqs+Zmlpr0z7pbOwk69kd0v1QoB8BXksza2Pnp9tWvWmzZ4VryxkvmzMuO3rWz
MUcQ5SL+HupPPXgMuzDtShLFBNGsihl0gy6hWWgrap3JoxdbB7vePmcm3YUIDmXs
m9+fYWKQasdsi7407elAjde+UNK4dxkcvt3eo41NqyNog/wST8h+ZdRxxOhHRNM8
14n3yIAczFFKAkKpThKZgTN/A4yLpbwWrlr+Ggl/EgwrgxKmxBJ4+1Wkp93N75uw
AiDcj3yJG2F24E19u6NM2guPd4RwXP5pCtb+9GHriLOUveqlThZfcKpDWSYvehJd
gPyb2KWv6v/mfna0pcuZrSxDRLp7lTI13sPcM0fJ1zS0PQuDgFQx2+WNvXBWwiUo
ltmztsSonmXtp8RDC9v5KNgX7fA4mhhJKeZOAN4UEt+55BsDeMHJzDkYoITLUJQe
9CvSYY6gkrqI+CWUsFPqBTHhvg5a+2Wdn3z/+5peAtINB6IA9C52QqDUWfw2/P7M
RnwBdAwi9Ei3esenj9NlVFzH0KRU+aCY2j/a9dHPxOaO+WE80YzNbGzZszNMsvx5
85onTfSBoU0m+R6HrbbgnPXxqfVdwaetQiGGrzO9ZF8LLbIaQm2G2+VuyD6rhtd+
pcLpxi7bAkxie4oNtiLL67oUUt11OAsmFntQbYAVsNV5qR83MaustaMhPgd3WNli
pgk9SNHAZCy26L9BoiGMJt02qxBj0373QiocpxFeAUg+HL6jVD1VNVo6zrmpj8Z5
oDuzl7mP5X1gXLxWdoK2xrVWxyZSGwGrvlyT4Uf7solOuiKENypxvWZ0aw36N4Ck
o8sDtZl2WfouUs68OAEStCj+lnWZfDJVhllfhZoDUm6ZykZwnuBWpKmKYnRQnTDh
68s0qqTKJsw9EJxB59c4KiJiqVWuj7g36itZ+WQp6WJLfY9oxHz2e/ATuswXxQ3z
Vw0D+U1qhgmmWCSLzm6E6CkmUeOLrFYXun2Lxh9W7VTyCUJgQqDFol/nZvaKorty
8H3IPezQf0rzNmM7bt3PLCSicVipcROO5CAE8/NluUCv2hxt3NYayqwacPpTr5Xr
aNp563gYSxdalCKQzEwFGW5onN52DkK6/6nYxY6kF7+vEhOkTkq8IRaP7tHgBkwQ
rP7vcQ842IWp1boq36J/zaGcuSH2+kf6mGrH+pEd8xSlevaERt653naxTiVaUheW
zRA+CZYTnFdtQ6T4+k/C3EknUF+TfSBMAPoHp2pi+0PfJ2AqRugKmVPvp3DNyiJP
FOztravk4hYhrlusVkiMbWb/CfTcZ9YbYBStYfGsyaX4gQRmanVPTPC+tjD3RHd1
MGAbjkrLF+FJ5wbxMgNfJw2jis1Dg5uqBCt6wyUsA9nF+1mCkoCE7wy50Z7E1qd1
bISYgmhCie3tWvQKP+DhBqi5fQgp5gMOUb5/ZSUEanyIqbFbLjeW9a4Wyu4XRVvA
YD+AGtrdAaDq6352anJ3W0pWplF13qx/2oolns7cbeiBWmHpqqngESqWYcNF9QTR
gEVqT+r5ZAgac54m+8DRmbF13ci6+45zPm2KrHGupZSEfdrjfo5ZuT6nPx6QbGB5
RldtXSR7telUFGLKITXunUGIQBWLdc4FBY6W0A1UFdtdbNOtLXaWTSFAGfXVMi7G
6NMj/yYSu8rgJ2HTJm2NXokhWzerIDUyAw9Rf+4dxBZBrH2Z7x9KTWhgrNtgqudx
qMMXTZsSHUe8C7QwogXN2I4It09RPMejMhEH6TH8I8xekElyh7s0uZuw8OXoyLTL
+FlvmYACX7aOg6TC8XblrR2Zf5/CkRDtizRuvwgm9uvnpwLi/hLBJKUqg111Zb/M
K52o/Cm9SAuDkQB0ntF0NO6B7OthbHxYQ0sZgs2899Zp6ltgqe2kmYosAVieCcg0
zF1DKIfsQMmxvNK9lf3FVR6wkotqGavIUWNHzZIAUGw8Ib4rd0cuErhk5KdFIkjt
T50gzqXmsnO/yhxzlfms8NgGjjZbtq5eePumV5+pZd/K17wl2kn+D6HxIDi09tAS
GPwZOxa6tzyYAmHyRGRKzpWwWHZO32R7b3M3m4HV881uDPo3EzyT1QzJWplbiMO0
QmMx21/csoHqg0MhMYYTmcgpnFcyQ1P/TuWI0+IayUxYGlxhzCZP2q769jZ+u7Ml
5wlaKYuoZFN9XBWpypvC3/MA4mRSowERnhsnBhLtnGO7lKoUki+PrZPD3wqvqyiL
MDF7/2j3ZPSrZki9VVLPJky0DebzpUuiIm6zhniA6OG+V/xJ/S1PlMMtXZCZPhMJ
ezIn3QTZrETlQNvwafdYcNpk09G7PJwEA4o8/FRZ0gzStZXY5EdKsg37kvuZzqWW
v1ZdxRcbKPzQrzH0MjRQOCTu6/MzOyqTuDsdYL+pYJLiknfUjphZwpql6oG4Idos
3dqFWE5pQ/VmTW+YjDytWM31FzbCae9wHuCGsnatbsndNAoVl03yz2CkTeiH0fte
i8udXK0znh/i1/Jbehxj30W/sBzLdeIPIufIgWMNM6JwLwi9II4KhhVbCF54hnPl
p+NTGGSfNw5t4FuQqwSZfd+r2RnIIWqcGlvSzTqt2VB3wSccD7NX92bqkiefEGCf
P6fJmq3BhWdZoNo2wlqLbJjbw3j4REK/2SmW/ezxhBiN/t02qYHZDaFyJuvhUu52
mzuaZvqmJRD01kdAEE4tXjodwj0HmAXqarOELasNdUO8w4g6yKAR+Yv9+TCyUeHZ
cupKozrB/sJbknuxJXEqE25+g7KdSOsw+LpO2+dmCxqJi3jzTvr8p/1M9aMltHS3
0jwZc0O1v6u9W6SvFA5/nxDpiLmQ1NHyXWpZZtAE8JN+NyYXCiT8+HuXUxaIsy3X
LAb+IypMBJnJxPp99eJKtaNywv2fYWrNRZsMZqtRty3zR+ckd+J1dti76CJxvYLx
sJLtUb6FC+BZEUNmjJkVT0RU73eTwZArCU06MF2nm+5MQCmfXtj/A6AXktyTYOT/
lz8WpKnCQoT/qYmVM/fwARfM5R7GRMXPaPQAQOnwwET2oC6/jCjQQDMFQCMiQu5s
RNtO4yPBN06a7261twBsG7PD9kLn7TmASU8BaasX+GGJN95yoNiyDjPJX9nuaboa
q2ye500QRHYoU6av9hEGqqnz1Dx6Sk705c33QJ93gwV4Jhfq4MDD/smHz/a+RrBS
IkhiQEsdydpnIHXFne26WuMFUronBsf9phIhPeDp8Xavtie87P9J1zM6BTujUNZl
q0LiS4fr6GOkrgdShb64vptRt+UoHsT28U1SGybehjqwAINYZUnfNKon7c/4HagN
Hsx5g7Lhy34sm3xRyXfGyfiv8oCCMH41XWyCuOyNj6pc1LyJbD3uoOvTab0IWxXc
b1KohBiwAPhXWOhCh1N4r7ChQi0ax9S2Noxf3HaXzeWGluE9hRMCYC/LLFLKTMmk
Qh5zYtxdLznR/MiKzABL+s3yQ+iwawjZliNLtMMtLXfdKYdhWAQ1slyE4nAAXSTl
Ex1LWfYRVn1QGD1S8imHjUF0dP7x0OJXPIEJB+Xzo8X0VXxZU+FSS9bPmx+QIf6H
2GILz5/tOzTGPWRVESb5P1eosyZAl9r4GFTP4QE0S37bopIW3jbIB8zrZigQXy2j
USb0DF2Yt03rJsvaxInnZ72ApamqV0geWSirhYRIOE0OSdley70YIYj+Hg23NCqO
AiEzNIXK1ZY20B3EMrIJhcgXEY6ZX6g4KLUVloYARxaK8sIbL8bByKURAhx+l5ty
OUcmibdat004o2+OVOkZU+rG6jPAvmqNJO0pt3yuC7BbUiJeor7zLWInXdVun9Xr
PmW1wBvl8JLY3SjeG6vbMEWRIf52vj8cCIPJfYzm+YWaDdZcWrm759b1hDGTpkTP
c64hTuQ63toyfMhgPWlL/MeAW+h9rDvyUliMclROtXiwLx6/sUxeaY3F+xrnkqHy
d9k6WjaT0UpjozIJcwSz/bXHPtLLom2g/SwfAkh7xwWDTGiqIdCQE+xi85XnHetD
iOaOUTB/tqcF6yRxCCNf8jLB4QH7INIepD8U+FSewWIE5tACkhBYugNK/BTVZIe6
F73tzvbkGZZtKDoMfNaMLZ1fli2hxIgTYZct8yBcySHsmEWewPX+Z3s+dtTYrwtu
ejJGAbl6sw0Lx6HE9HGzMmfleO2z1XPpiodG+iOXf4vmMcatrg37H5zQZUqxoiW5
kwi0aPZwKqzcA6rQ8dIUMPS0g//k0K8QF7HCTcNUXwRRJXDxBYWaLB8wYivCXBfE
Zj4qEU7EqHJlnA3BkQ0KGuFEJpaO7NCJzD2Q3fwSupYwX6LxDohJ87sJxOc6E6fJ
EzumXUqUfuxLqbK9GdmKgUz9hNexgESwb6ryGTObrrk5NDRhJbeSRUYhnWBqLIT9
lktfB5ZywzteGw/nsu2SLxgqKJ1AVSvhiHHthpxkOlGoN4qIHanlUM4b8Pw4dh+/
+tqcGYtl9YnfcOnHOmLRYx+GNsHjcU00uO1Wkpib85TXc2WweMGw8/XTXwpuw6vX
0jU51cBUtarpnNReYD14EnJ17dEMFI0fCPmhs+bCPqttn6JRa7d1fAmIXvFa7ZFJ
V7jNVZvupybRHOsblnGfGi+bp6sdfDoTMBfKZM6peo5kFNR/3F778FcXXT/SxIDC
S/rxAGDgqnt+pdbm8Asf3KxQhaN5nbG0sfNBO9YKbqb5jMc8CvTlM2Rip0Ygis5D
xL3AYqqfFa93tPFxiwEIEQkiSUG6PNw20Gc+9W7133ChUo+bkluhWCRTitoemQ69
lxGZZfsL0nnqmhTKkqemq8AFM8EFCGvE3AXq/vnigbPcCtPZn4xptqcmK2Ea2m2f
4NOKdicOwmVYoW4t6TqkYCSxGFN5pkex9WcTQGHCS3a7BzfYtPNP0eJGJn77QI6o
GD7DSdzWgUkjzZ77gJmP04t8l4KWTtIpzT8Rd+tcDXacMySh3MoT2o8OBPilokIA
GKG/JBD632PYpAeUC0uTiZtgrb35iKU46PKwB/6oBDzV4BsQ6YzVGWWVRASz9Hva
llULNTr8Nf0HuodrFQwWY1i75TEBmR0ffT5vJVvo8lU7rBDDTwbPIh489meXo5U3
t24u1AbPz1DrbUInIwWgMR5aHUpA8YK28gzH7Js/GFE8Odx/ywDivzm9HfsZWdwC
fapm3VwbVhdv0KbosBTOG0Vg+tn+TqEsrCzA1fYdxCw0a9hemkG4qeaGR3AiH6HY
uq/91Ghcu2k1JrPhDxc4TRPWppTKIB1manmFoHvf6JDRhcO08cd/3tbUZT6RQtyM
8bM0FOnHDEsaBNdSmPRkZHxl5e85BX0Qy8oQevL+8+9r80sbS8Y3DWVAgfa7VN6m
PpqYl0rdB7ixgo6+Uc9w7i2ETh+LxROl96xio4A4UAH1GqGsVytTZnMNU+TtuVrK
liMh054aRMOy3nHs+8IdxEr0j6ndPGbC9+T+X6NBLl55LzpU1nCAHl8nMhN9w0Sc
Aspjt2D6elpb9RlOyN/1neHvISVq+NQEgt1XM2a2o9pBeMb/E+1EewnFtNVgMrqs
+KdY24OguYPbdVfd29MM3GyKeYcu6VC8/ytclUj5sGDueY0+lRwOBFYgIkE4lQJk
7OEpB9D9lnXS9Wx1rdt5LJgUzxtla7ZNCaXT8wEcCQuB8RgcMU5QPDYRDcYMD4O5
lV46+ObdkVCwmt+JdD54OKg/j6w6dn3Lo+eVKgkYuI4x9Dv41Fcj9uPR3+LGXtkn
5Y4FXlIpWd8gpPPcB2owuiml6yLoLjHLEjHsw5Y+owg4ieIsEk/7IpgGmjOlShdd
Ff23dw1PdYepFp8S4kscCskN7Qd3oMGd4SnuYqSc66XYyPv+UvflSZGuUv+1UHr7
dz/VvPUrY/vXVMEb5+Krp+edUFh+5MejxPW3gzWgNRkkcYa4cYlvTOEjXe0LVF1d
xSPRxjddaz/lujJbJ2zod+GdAFFqvSCXrb9mgbjqa13EOWVD07fENVV4MK1uts/k
R4qxAXWiqvkJbPKJWthzUPLZboZy44o4S/8XwvusNOO1bpVHfiXbdHKoYHunxdSP
fTH+KPEwLygWrDAp+zihtFnZuXPSh/ZBozn3gyfGHMD4ynobHeNKFqDrBwL4NLvz
XrlR3Ecz7DU23YysAsXMS+oXYF9YHGhV6GQCi4ZXV17spMI6ZZ/jupuc7xgu9hIr
GlnlrZ+iNVqQ2alEp4r91czGep8b2F2LK0WrfWRNo+ReCUMRKPuzAtI4PhYvSUQK
P6NzW0J9DDeWuSRUQY69mvKqOlHE50YxOYJ7yAqudlkIDaGcZ81Rc/dSeiAgRyfj
knxff6USgNLOJoPmzXwzfhUyj3gxRveh4NvXnBT502iWBuQAiYWkMS/drazLnpHa
iXMnSbfvjm1yVf1w+4i6YQ0UAMQ4D3UZi7YlnTORuz6Oy3O05PjP18x3Izn1gr+b
st0EbRGdKDNl8sWVzMnT47k4G5ocXSCfIkBU9VHmFhwZmBGjma+0IDHdBsC3n+Ho
T2gQ5hBSCLa8StwUCupa9g32vLpZEQiic5xIzg7Zq83z81SQge0u/kA/tY9izyTA
ipBG1GZgZCy1N6gRK4TirxrbZ2laU81HvUALYTRxKRr45V6ti5kBg9YR/GVqYgDk
2PBYE5w2KWrncOR2YPLu/ztM+yNkLTqu5keyB266P30via3V+4Ln1t6T38Lai1ea
NnyIPHhQLdOf2j03mg1foEN4Z/xB32SnMdotXiwVhrg4HGEhxWEE5+nxz8yw5JKV
2Ne/fYd7hs/NLize8nkjJG95JGzSd7ISXLIX2UOlaGwT8hdHYZO0kGTHtixHdsmJ
efT9ygf8MLALstFbNYFUwpSF8/S8tk797CtQhoBRCNkB44243KyUcyDmvmrsqGXg
IKpyKcutOhxLfaBndAb0gdw3W5umhnFVQILN18D8I6eyBEI2ZS5cjooByiTrSuhP
sEKb66Lu/i50cBOIlOh3SdApMheJrc3Lg/ObhRJueupqR4wINj8tOgBSB3CHH9sw
3XFf3jprVPpRY1/XSw9ZBad1fMRKmR9PUfN6alI6NmijpJRUz8wqbQv+yLh0vHQs
1rB5UUSXMeKSC0/ZI54v2SSxwn8kpvI2jST1pczsv3UYL8OhNvwQHjomp50cwS51
euNJI6I5H5WaN/FRTD0LZsl6Ta2rtz/sknug5a+pHEY5NNthBJ4eAtRzbzdROKn1
Y0KWvSkwsS3gMzuZc/kR4yRVHMTUIl5+Djk4xKxqOizBxscbObCwmyGPGT9KxxIs
tbDzl/iOqSc6rOoHGnV8uCMjFClrsLIFk4fUUua0eia5z2M9RgicxMuFMcJQtQMV
LDWhUHfskW9yx40PH3w2SBuUllxYWuYmCQcGAXgFkbOp13IKDVm8KzxQ7BHAPguj
Q3NPLPqfjOBPx1RWATM34wh4hhHVFJGnc3QyiuRXQpl3kUw9owLXNTWU8Ak4GmP5
BB2qzS4JPF2Gwz0LDUNBFsutLQe55ZJmj+ImoHzkNzEFn8YMm9A2vWcSbdUvmjQ8
PXKc0wwnB24+/BNtcT9KYhGtT/4jXPCNa8unLyRtW4IXopF1PKujXfc6MXpD8xW5
ojnwlEU6gaffDTi4jdU9PvX+/h3Xvgp4Bzym3CEltz+uZ1QifkJI0dYGVmah3PTg
DdXepMwWUT6yxa0aL+QI/l/zVjLwHchVHjdo22dsGe8JPeN+5wHVSU6RN5bpVdBd
xP4mz1z4dMNMsxuYPeqCdUpznqOpvpDYjkxAEZhYSJHx8lzjZz4bRBVfnVGxLmJo
X+EazEymD3Kib8Ol0gtYpI1nZo7A+YaPr4RR7ITPr4qD6rQU+2A6FZek7pc4wyMh
0tuQrUqXMTYZygLokglf1YtZCSELHlZBoa9s9onbyAaIX+uo8v92eRXThvlNd/XB
r2AgBFoneZ2uUEKcMHavyCyKqfqcBTvEXmeNrbKCct6NnVFd6I/xt9nO3WbIeIt/
3LS8enOu+zMg6z6Dnk/WBcqeorB9bZR+sTIu3jDJ99rCaocIVXkxMmnICE291J+F
kFYgObK5slAqqLkBJj+LnEduICDz4OOAJbRp0XT6mMJOMU94Cwwock1KeGs1Jf4g
wC0pnl4htFK51JxHj9ZHBK21IfNP4fscQMRURYrbfF/DGzg4TFUm4wrSgqurwfdh
gUOXHIz2NW8eE8zVsZKd5B7TzIUhSwPN0vjXzMQfYPUxub4UtDEjn1aATorwMH5l
Ebi5Zn9QNSCAFgnrCKQMs19IZ9gmY2FTasi9pPlaGMqWeUwZJaJfCfKHfQWtLm7I
C4N9mpuGFc+rLyWy3OXXUkuUdLyoSf2XJD32j49CE7KzfWH4SAjN2u05zv3V6xDE
+w9d41p+NrMeuzlxvnRo8ISbmOTb0HzFaV0ZVjhTN+d52IL+lNAXr/AIY5uAVEKk
WvmNrjTvHFRafgfgAMnCXxjy4E1XAk1lxAeIkpc1v7TeBVf6VUgHOo/L9+JYsmPQ
Hmeq7Rf2TIsgqkWYNnDlXGlWt5dU6Ya/FT9IOaCTuQQxGJGn4DldGyfj7aoeD46f
0pCDYYO8iHckKmaKbHYsBzsspel7HZcGfRfd2f9SNxT/9kZZDf9ll3jx3+29opqn
GAKwJaLil964e2IrlOQjBBjN66qu0pklUMPBpIGdSquFPPdtIrzeJjjDH32mfsC2
MQP6QFO9K3WZvPLVyO1AS1PvtpaFbU/Jaxu1ch+WDp1PYBa+mTlw/6c8gtI28Dqn
DAA1P4PDUWGYFqwy8r6KkWIwFSk4FjylGfP9muDzfjRV9bwvdLi2FDG892criXuC
ZX0kCb0bNKHDCwqDQ6CBQfZBmv9lNPno2Sxxtxly534Ak+MZ9f2a35pJxxMgUeQG
W0GOnLrooJv3mLa9Z3Y4fcpWoHRH05FD3gHpwUbgM7foGH/prrzG7cRtrM2wobsu
oKKag+zJmmEUld/OEzCJfupekFZt6z8g5uutQqEtNijbcUGzlCV/ZJ1d1+Nuueke
/jy+qIyZfgfi/uR4YYitvuJhs7e8k7QOV+YIUztLeye8PrbSlliYk7XIEJQtAgJa
Oeq177oUWaXdCbGrHqTiPa3bWMIanZpDWWEd8gOQ6IIVL/siKur+POdzzztOZgkL
XNfwNssPyruOr4qOjIvTLctNt9Bx9849sjce6wUOJQaoYr1h7vl3ML3BWRsxpg7Q
ilUfSc/Qzno7NWxViETPOQqa0fLxovArKM+gSKDJTRxLldX/5jiigeiwVBK1lpgg
LqimbZRee31YVPR2S641v7Lu3j9adLMsAAY86o2ky1jAwPI8CkanQ0xDWq97JJD1
hH2Mk3k9UQHlxN++EzR1hlxOfilTDXLwjtVnCsyvxFbIqZ17WQc5gg/gC5Bo860i
3DHQbf9/CLN6nwwt1u6iSMGHgYpoOPFRBoZqTaKiopmt5FpUKWZfs392x86inVgH
NyrYfqdUBR0MVUu78QKdkr99hxp5WSHNMtF8M4uzmKg4CY+3RFTd+xRkVwiuDDJ7
9P+OXiIZ937O4HGC+J0dk4UbqiMuvgEZY3Evi/K9HsFrMxzp8i67MDGy6maWih3Y
kOkwCL5zzk1TkyNDsPcOODYH9GDy/Q6WWZftzDIU8pWKaCGNUvXitYWvsEWeI2er
hZLR93POX22Y0Vu1Tree7c01WSVfSYYdWiTwTMavA8pkZZk2VgJrgeWjE2TCLrW8
/XEA2xhzGZuEF3YyZDjqUieh0JTE21ibNTSzZVbaj/UorCmdIZ++DTkREe3UpHGe
myJG9uN+3jz2y1rOTlLHNBSeOoNE6XJJJijRJdZRzrUo5bUr4fAE+8wXZqdFTXbC
pugtVhziXKSKeiz7YuDdn9HNzs8MoRnumLrVf3LqUfh88ryN7IUvSx3xtv7W4hUW
zIVtd+sRjKIUQXZgs0DHNA5YXH3m6LkhvPLLmG3/RaxGIpXGuAjKdwwblus4wRfV
z8NK2zz/a7rMQLKLi9R5ayYJxaTHnVpAk7BeKvmvM+VVXUMr6ltLRBEHzbAtIJHD
Y5f2o+ewHY/WWQDC5ph2X5/y7AHxtybwp5k6UEQGWzDzWsFKflVxI3DDU6J62X6A
5yQWqM+xFKrsDJrtIGCSqW7z9iyEO4srwqzgN/IKztFGip29FydwXzr3HcXcmnMH
HwW78x6Sm3qjOKVD9UQ5z0EkW14qxumB+YmF1zgEhhiuTBkNavTWoWvf4tR5FOt7
Y4n96xZGngh5GkrfRJaH/frq/tFn2/zXvVvoKT4YkEFCtOoxEUyoRgdSX15nGrJ1
RWhww6MMcJZSEosg6gDUdVt92lM5B5o+Lch/cWIsch3r1WMrEyIxyXgH1gZtnySY
qn+fwxOWf9vhDIGuRobcOeqItR9MHvycFFjYl2opeoU2wjJ8d4tQ6AW6GAYpCRuy
Y/+Pc9ozbk51fqk9APH7jLlMkc+KV4kEiOcrOoOXYJUq8qil7eZ6Kl2h3TT9Dpz3
pklQJEaw8P7K2GAKhORqW7aQBuQDwvTBvqsJYsJOa4U9OiscIS1MGaS5xgQRj7Qh
GgMvm1pJC34Gyl9rmVnI6NXlhyS0FMSJPeC2mFCK4y9RTpVVwyiy8/Jmxwb3Zsnr
6sLnkKX4kDNGOyNBvaIVWujfIx2r9vwiiwbyBCv1IIKY3CvOY7SL01eqaEsug1gZ
TdHn8auvYmdj4P4L5nCTZF36MeukmSbSJEOQe0YT/djO+s7/+mX3fl2WeCyzF+Ks
l0yqzhHCnlr05b8vBGQ8xGhIbn+/JqtYfQOT/tpn+//+7D+A1u1Su8lxaUCpEgpg
4ZJPW6Tw6YqwBQBGQ4cKIMtDdssVwkfnqMwMhiodpPSvVIpR+4PVc6kIJYB1q67a
yigVHczQpDF+Vxbz5vdgdxbPSz3uHbfsPzxcGs7ibgfkbgiXfxiPHIa738LbNBDQ
gnqEdF7NSKzirZhYsG0e2cNv+H8eQquxrb8nSuCb6TzmHf26cOI7idmVZl2YpoQk
H3+wa7fZym7bCfxCVbazhId6vWF8IBN+kPekpV1rYARw50dyDmD7lgUnvRGZzjx5
jKqyxDQH39HkZ8U95KMpx+rVpsLLsVAqpf7UPjHvin++OerxAJlp7lH8ixROtbJK
vHkpjp5FwJvFDVOuSxipraYL3D95E7ZvawJWaOd0gXpGi0u4yPM3Xw1qatZ/Ga3c
HxLEgou38gqI7tEcfAYpGvZialq2ynno7Ygwhbitx2mQ38cLc78KJiuwVGNTeyk1
irJWUfuV8pe2pjp+fD/jGwkzGSQEqs+g816u4Vv1nFbrIcMzkJwAzysnV7/cVjhF
6bt50iBQvVEH1niOD5HNIIL7r+CLuFn50AFgPvWvBjFCIw4Z+TYadhz5MY/wKYTt
HBun9OEg+IFFpCr8pgYbuZxIx1URNlH7NRxSzg63TiWe3HNK3s0c6NCSmxsWepgr
IglbMU/QerVfPxTK8X8objzId+S9BK4EESJ8NN6wBHUm0juTpIFNehoRf5O5qmuh
Mcws4Qvyl37pjaG6c1OVzqzpIVGVUr9KFQMOVoD+ynCHG3/XofgEJlg3wyQkfch/
OrxEGe0t9NteGV84QdphU2sPcOXb5H9+tG+YROv6XHPF4TTn2hk3kuDTAOq5WMqv
PFYE+re4ARhntgDeRHtVa+yVTnzXYbqz8ehhDHV/KsaxDdTtG5PHAUXauAYpJoUZ
kjPD2xLdj0EQHDbWCmBei7juKEs7r4yp7WHa4jUfgxjU9AfsiUG7UG+oWUS8RaIE
+ff34XgZ5fT5cEJZY7VYeFOG61HcGo1hIULUi6tUTJSOjYIioi+K97H4pQXtl2ch
cdyIAlKrpnyBF1OEyZcZ23K7R1W3QkDODoeWr0ln4Ct1+PkLW0fyyUz8RB8G0Xq8
Q4EG2u4F3bmxqdNpSCeGuij83C0Ive/9da60WBoUnm6aneEf5sR3JS1b7iTf2RPU
b+Rvn/2dtVSG3mu+pD1GbLhWu7rxH13Go9864prpZRPN7uemeqx5zXbKyOiyESZG
qgkdn0B5709LPpgY9BySwpLg0N1uDTYi7JHvmxZ9GFM+Rh1Q8j6wSgAHw5btJ5QJ
OJDzfKI4sAIyfIiXO3mvYlMhpnoOwu5mhMuEYXao/nqi01XA/JaNjfq+1ePjAxXL
09UEY/FJhhi9QSIyHkyWtlXYliS1ddwahSqBWIrPRc4VCLXdjI9d8QOTjfcUmMvr
eaqXSUm4NsYX+pzoJcZQeelu2u7kDguncOJ09SjTYbg11TIWOZjI6i9iyfLC0p0+
w1cBAOU19rAKpWqxPN4ihxa8sc783M6Twa7dXsLlJsAFxU8CLYvflSFdcaUuYJ3A
BJgaWPVtgKT5RVIyh0zVfKK9J5D9MioMEj9UM6BBD+zymIDdCT58YPuY6qIKfpkT
OWxOvSpPPLibgu8Gqp9okeguvWGFt0e+RLgSX+ODueYHV77ZigNR0B19Eh4adDTS
t2gIm/qjxqUdM1JtFPgmK0smqqaI5VqrfI6NjkHt6QiQC1oTXmSpwadXrwFaPd9r
6u4Sc9PYu2IAfTkFflyStVzd/wn19k/6OR5qFz5cG0ygMMB4+PYo02HmIfsSoeJZ
KGe3Ldaiul9/n+qrHDSvLBcq6XklK1acT1kWb0DlhP56FED5/R0bQFKUj8G+s2Ce
nqnHld0+0PhNfFp8ooJzv6mUDRUy1O4rdPvyn7HO92w/XDV38bBwlTMK0hyNzI69
xEVc8CjlQ7MxCgdi72u67038aAO2S5LnULEM5onz03J0vAHL3aCdmlZTiwAkwQ1/
oYePDq1aTDoMHiMowDNGyVEnMXpqEu50lDu2tknd3u1OWo7s05AQEZVF5AfFqt9x
q1m0PmuSyAxsCmilRoRmqlo6va4ncU2N63rUEZfO97hLcGitfXeDOHx/wQWWCxDG
gA+tNza0bseXKxvOvXz2PLxjEsfRPfMCIJNOmvBel89XPhPltJgoKKalVHnNbEhB
sz5gizZfunTj5mnzPSlTnUSLZ4LQFSVGj97V4+4ckCSs54tjWnBk2N45QMEFpcdI
BWF6vtt0rsxXDfrvnhxF4aJyjvxptGLpmwpM31zrAI/N2z8SnUaOliZmb1y4R4wm
8LsPQJH5tDy0kh3lp6WMofcY6W33EJkAvrVtrEDcshpK+w188eDAhnIDYeaEvRnS
EWWErTkoixehY+7hRPDa4jCFdUZYlBY2RNRWf3fp8gpBomuHp91vim0yopxQs7dn
RZW5iFYOw2TXkgB0HRcVm/pNHbih/g6wMy4aV8T66+cpsSvYjEJaGKl6aLPzLXGz
DLr3elUZjQvR+m0TYOwZ4tVv9DE1phNeKTla5+Qf5wUmodaAsDh4O1E2oO2E8nfD
LxETr/Jftuh81OJCqC4ZKWkp3O8fNjdi57xDipnigpfQ9gHeCgvSA47rZVnYl216
nb/ahzCwWx18PSgCvD8n6N3DIz337QN6pXeqfzc3HKlXpvUI40iVbiygPnrBWHKp
v9muPlHOuhhHCV4giuFnx9s9IP8WD5snzWPsYE3E3S0LNALdJZ4ASXoWc20f+kGh
k4LiflV/4LamgQaKEqjBTUg9LLBTdtCLIO2s0oMTChs2xouEdJNPbs/eCaSci76G
RmIQ2E1b4eKQ/bFcJqsyiaf89S3nbHoIlWurHN5koCdfk+PAQ/tSdupA8q1oow4s
dw6cbnyMh5nPUMJCVC9uyb0QarpRIA+eC9TPjQFJz8hdV17QO3XYDhDYEH2urmFZ
E4Whjf3yDA7iq72bXlkxwHcFUuE5GGqW42zOxViMNVsn6xYgvtdMR9rKekema9lA
cx25qJ/bwjxvCUvo0SDFPD1zKgp1ptBHoO8lc0RK61ZUSy4WyVvJTIP9iflyrCwE
qTzjf0cxVROB8b6eVgWWNus4cDy4ZXR2PIQmcsJFRad30iezOTRrvzg6zqajNfTh
UoUHGeGqvkjIWYXDhh840+8MScj9MPAusDpdsbJtlsCtZOIJjTsaHRZtEANNEfqn
5kJrDxmnfuTphOVz5EolCVZXQDt4vpU8NxHo6VC1b829r37E7vUOAiVGOpzZ1/Kl
w8VAOkPQi9RFVWi1WOAMdw3JWy5s5JLrVehOvLXIRFojVXLRSR3/bY6rEq/tf2Nw
83puBAujKWoEszk8E4CSqlj5+WdmwGDjsoAWvPdkrjvlJtGSHpgEPeTQEiCmD/FD
s7Q1fsQ6i2JqvllVT3QmX/SjSMb/Qk7lEX0GE058ktBk4FBzijihpYlMmSvVCwJa
8UB50p8kuoOMHkHxf9VDr3o/gPLBN9sFATsIfBZfoCWqqvsrh2Rf6hNOmWCwS0B7
xed7mdct5bF/sGi4qY9DCnvEy10iL6Ndok8/NfxCwXvNacwgccw4OrT6nyT2p3DT
8/wQFYzbEJqHSNdnIKRQ/fcYQeNRgD/6plgEQ/Ozrr2ApoHd2G4vGxohWOYJMhJe
vEHiidruidrwU6Kaf6bmJ/1GECqoSTK726aJPFR58CDnuJKBqEVadI/wduj+A8nS
1WrabupT1wEYhahZg8iHk9rDwQvAMXzFAVe5hUYErp6IGUKolkmTf1uyeMhzt6+P
DeTNZA1MNVxOHJsD0ym/8wSAy4X3mxCGv7TFOIMN/7Hcl8gyGAax99HzwxtRU4ig
cJTttbz2h2HbnNV8beaZ7QnNaOy/UwsszuNkGTKBDM8sRPUfP5cxqKmsFJ4IGnTU
FDTrsFU4vxjsxsk9XQLEsdnLB3gPnPyBcj/WONRIMcr9P7CgiIHu+QvZQxe716My
kogVKJ4F6A/s5HeSkxknntERchytsjF49JP2Y0pHrVFocoiagwbU6fBuAcs/FUgI
iVRng3aRyC4GHEEP3Fm/JVMGsEtVqKpe1Cwhso1EWIMc9TuHz+acARlfvTxPKlRT
B19wAxmzHp+La2neVPS7JnHWBdLemOqFrF0slQu5vP/JcmKWxGaAcahmn8I+bZCk
TczjuRChmBu9YpnmYkakRD1aFS6/En71wYMch9w44RD2HGH5HAv6j0nV1Ujt0F5F
4FWuv0pvB5nXV9D7m5TzHWtNjCLufDCPvbOxdOlVKgLYlxDLs3OaIvm/NYdi9kHN
B8mRLc85LAdpO/ijxhh+twdItMaGLerPf0/QBbuoSzQxy5duV6a87xGTTo46IrIu
fbxtrQHZflGJI9NLT41K4GHL0NlFznGYp1DABZMCBtbpmYgGipPmxtqtxjgmUEPq
cJjnMaUwyta+md6D3650KK78wKtaT+3x35FeJrCKD84J8WiypesX40CheHlLgkPp
w1OdN+IVPQ19PSEDqz8BFUSiwowAfdQJ0wCMVL1PPU/EVwueuO1cjJovmKlWHLNY
WPNoQcAi/XWyNBzIhQtuRHjg4oUoBlvxbil5K0Xz4Xv+L5My/1KDpKTnHXdruj18
EhVF6qG+XRilK+M57GVfUf+89LvUEYdgWFUL36NSusyXgq/BBSblotxwsruyzskS
eEAby9ziia+nsiYT3xDiUl7XsFdFscennbGBgq9SETXXYeehYXeQ+LteR7FyTTJk
yqSuMNYUjky8D2PAGYFGdJsioF9ZSfDKKwYCPzYhPPr8ys0BHM1frozH9oPVIk3q
qqCrfyrnmGBh3auIRvZWkUZywnGbwMiF9ECtbfzNNva7noldbJgwlkWUIW8FX2o3
WgNg5iYc03cSELxYwHrENWlcVueGQ8YJbpHkJnGKxeeSE4yVM8nERHh0QfifUgTF
DGw1W8ka83GolhqMOI3HMgN+11LizaeLwCGOmXTX49VXgL7/OrF0RH6FLMuBbFlW
IiG/zpjtx5zZoGEd6etn7GMfLeQn/mA+eKKw1HNtpx2+OwtC2HXJd63d/2Daf5cr
/VUqwg9/16lT3x65+1TzV4PaqIzGRfHq0srvA2YgkZRhvxtvc4lY2RyQJ+Du617V
s1KFBB230pGQRLBrWHxk1/UN1J36WRQ/OB1NCvkrn95aU4QQ5ORr8+9ymqWesrne
Jkx48RlQ+jtJoGs06xY3jUYwvO8lrtyr0NzAp6YamwcERPWdSxwv2l8hZdgrkIO7
BHlm5MRS2hNWGYEuEH6qz9kO0oWesCpY0nArF7v/BjNGcVQMjDrMGSN5oOQ3n5/O
S5DKv4DECcaRoM5FSflyU2T0Fnn4qrc4VAJ3hWfZPLJdcnAq3lov6LXctDbrthMY
iQW8TpsdJB8J/z7v8dGfKom77g3529KI/xs5OanweiHuLsv3Pjtnep1rE4Gxnceo
5EdIrgsgOP8BjPVutr9b6gmeWk+61JHCrBaxHcJGJ8jUrJT5UjtKFL3yPcGEsUBs
AEgnFCpeZYIBqQFz32WlobR491Ji+gSYUsDbUk470NP7lsjWF1ETc77QSVF981Mq
UQl0IRg/ECkUICd24mG2QRCfx7FaTsN0np//Y/H5cGODKedhq1IbsofKIC5VWZaM
2KQHb02BrvqdmUqoYZXP987JlkIqRx378qrfCtuTtQ4Tt1dL+UJtq3pnJ4pZjK+y
tIKa9QtTxjQt7Snn4Z+aB4avD/0o6dJdkmjNWLKZhHMVm5a7KbJhcOrfIGnzEKCV
tb6zJWfJ3rcPH/6Usd9f4DAE/6a9CBQK1YooVRuwjo8cfeYSb8rq4SkUblzoFLNn
XZiMzlUkziX3y4kZdQJcIcFF8mqQJmiH1JiNfGZcZ7MfcZfU+MPa0qsci4/h4IQx
lRiCsBR2C6oZK1AIa9bpAg1LtXKp38vRRSMCNv1MmjwvDBC0kKQYfsw+K/fvJCZC
b2AFdA2WeupoWS4RjnphfgXnM6WADKSEPgu/LdGZOSXC6g/Tjfa2GUD6z/h0GaPR
VdQtrB5b0dJM9i4miNE388OQM+cr+JaoKdG1V5rYwXBz4bFf0jv2AOiN/BGydUtH
04Fay7We0msQQm+ELnPFKWFoLYMlRqVSb0YPsAFb9g6dO5odpiv2lA4pv+amS3hX
DMZC1kw01vjMTSAJuUx+6f++JM6mNpWfN90m1SbSFJMLun8Az8yqjHpvqaKnEt/d
yk75t0iVc1bbY557UwqCcIrSTDTIqz3VoBFkYn5NBWWXtURpS6XCgs7uo7LIkGA+
2pAo0cdaF2OtZN/FCQFC3w2oQAFVsXUPVZVnRfdoPbLQoaVOTDqGtsFe2Ve86DGw
t6kY/zCeNLSRzJWySGrcwZUJljw+VdxsF8SmjUiW5GSzZ9QVQ20PzIIkYVK8ahYa
rk0ojeRoIEG2XJRiQXt8yQCP0YjPNsH0+ObON22pQs+KrbLZ+7So45W53iYiqbjh
iqc8GwBqsljXG1G1EI8Pl2VjlSDAbjGAIyAxYHHxCF/DJClNsGyioAxHvqjsT7lY
5nGVy6ZuXXcEEiFOXaGpPdkpQaA0F8qYs4Xmuai7dSzDdum+DYVrCAT5GpU3j4YD
I12EuHmbQxYt+JS4WGtquuvkpTHCEphZydj2X2BVHj3mweuVuoyR5GLyGxa/IHvb
kIC9K57byrsNvOJJSClyDSdQwUUWRqFTx3WVcldrwCVv3/UDH9esZaI5toTn8Rd/
Gj5dVVoVu01oVe6jJJ0dtOAKmV+I1fPpp9IEcew+iTZj9zcc4ACuRuxPwfrWO67F
BvHUq6xs5GiFvSTSkbKkxTxTkM2DljfaRcu5tAxHfsjQzRSmC4Iz3/qAaPku+sSO
Sw46V6u9O/mccR5Utc8xKT3BrhXn9qgCuRZx3X/asDk4HTCSnQMf46nkpRWKJ0bK
fopaYNrApp3CAMmYwxcA5rryC+5CbiMvaH5NZV2SMnZGXtdI8wAT2IwhM3SIl4wT
/Xf1/ElmOrR6siogjiFaSv46Tuf/ardP04dGkfiJQMvsn/y8TzgOxqpG8Z7aDpGE
NEWQStFriXSlphSgsSUPNYfXJGBUjRSTd930+8rqAaXv4F60u5mR8MJ1FNh5z5qn
ReGl8N0Zjm+iSrJOY6Dhpgh77U88C2fKlECrcz67eMRsneIFj/w4wO4skLSnQ6ZU
gKIX/Ctg2boygcy3X/7aZQ96fjsLtWZ0gQPA2CQI37b2HoZz/nVw2rsyA7haewN8
SJr80aVtnFmwtU6FUeKNetoFZCIWy5SKD+x6OC/2RrG5O12kWdZ6JyFXwT1viSAj
AaFyJrn4U541YHmSjW1JJ8IAXTezVWWMHo/d/d1nkVjIQceWiV9ENTBd43ZVJMXD
OtKhSSYFFerHipUpgCXaX6OqBSKsBKzNhO/5C8dpvMa5tZzCPJSPtTuVVeoq+ahQ
q5gkNnV7i85p5iERro7OWrOCJvHH2Os6N8STGWkeAcz7/ja65yvyyg6zHnvG4zoY
BgdZIlBDfn0VE7pWBYmYi3XUx4y+16UOUrsgx6Kr39N303/I3vIXHhdBOww1Q3st
IiafkMdQdCFjhNjfhvnH/+pd/ifEBmmPmp/IIs3GJpg4qV5L5PJAiqh6w5t0HjTl
nSLjGJ2td/ALT/VOybT+OHiwBsqKPdWVZ+MItKhZAkSSRp5VVxF7VsXuQXUMyBGZ
7m2ckuRv73KNdaK68WCpYe7DEJgGaPNHuwCcx0ib/hTpXcGAE2sff7H5M9YIqMa2
N77QTotkmcjtEcTFr7hPUIrKMat+Heg1BZ/7Swr6is62b0aYftR9GALmJ0fYkYpY
nudpiQP3ASgc3VIjwG5rKEn2sLHRCzHPSMCn2IWGZAD0gwBQRQr70dxMFGbKWffj
ZKrPMSDoI86hXDHEpb8ZW5n6N/jtkFOGL0EVmRQkQCDuMaLGCIJNygaI8JKP8bRH
Mo0w2X1aMhwniKdfIptI3D5XQ6y2YiPzvxmtwnithgPv5nJra/jID3aYrQpqzqKf
bsQSzAhgAzQpycYpdNqLvq59mRFvUWvZN/Sd3z6FX0Q6O4jjVCDIZ8zAIJFGP4re
77bM53ebPKYteQp5w+xQWrFKYHOtDeM3ZOO5sa11Wmoahj3EtBp8aw8cSXXshqUv
9Yt1zllqs938BWk4I4JJDF7HljWMb4318Sk9Pkt+F9BbggRJGiuiwxN+3MyQ/F9q
2ZCfpx8mi4fBrD0TeAxleUH008wBWnIn+SVAXy5B45UdfL3i9Qz/GMvBVnxzgO0V
lXt0ui/fFZ2KDkCDXnPccce/jlwMhDSE+JE3237h558nUM4uO/oqtGrLbWPO66q5
IKSHD2QzmmVTXUoiCeJQ1XVd7q+yVERRuVqcMXEAcyY1wMxoD6yhLqq+AhSorLrO
lpjMvYakeCtQKU82XFOAvvxDPNKpPyt4riMyJd8EJ6J/il1anyf34WEtb0ZYF08B
dcFbCK8skupZZ86LPikNWHvv8+2f9OOp57v+nwvpXUteV4Ycwp2JfeFCP9YlPcO8
mUjoZc4LAv1P2ZWd1ZR3yFaGz2u7GNmDM11xlqUAEfEMvg6CnrB4JINPtdnviRZs
bIjgi78dzy8hgUKGzmg2w2H5f2EkTfJrDhGrPeMSuaNQODsOnnVFVhHNXie0MdgD
No/KlCNcjYCIQlaW6BmXuD1HHQgD5tVKrlx3erwRodkccEiciTeAksEC+qvS+VV6
3VFiLR+JqbKR3G/7hbB2kUEGFzhXAf6m4LUHPH1WCtyFIXJj6ukLQ/PeAaaAyTxH
kWYPin1RlwU7y6bdWSXr9xmeV7ab/eDr9n6vDJBm+4JTMXwuACp9fDols+k+kQ/V
1ew0Ije+20Pq9VdhQgn1rZ6BtXGLw/1sGpxMRMw6Gg0sSc2/OO4RfbQksKR+lDN3
HF2zqznPiHChYcZgAxRKSvfgAKG9QJa9kl/vs0UHWfIVubP2Mr1u1v8y0JaM4IvU
rlQIMezp1es7q98CuZ8QH/zH8/03tRVlGmcLtR5cK0MXDz7LdzWi/HjShra265KF
7zQpo/blttGUTr3ug7FbIkXgxp6EXv4d4hMA/CujuECxd6vI7zuaiTkjBELEmPsa
8bWrvOFfqidFrMl37YfgdrhOT36VB4IQ+mmTVVZGPnvdI+4t6Ek41YYxyOVf04Fk
T6+PkWV1I8mWcH2ySIvAqz5fcuIcA5dQLzZBUdjTw3/izOIs0UxXZ74uWAzTi4vm
tcbPTOqxFCvfFZ62sC590Kxn/JKfFn+zmBlirUcde1iRZzF0kvmpo6rdKYm4RvFU
KNaSgs0pfYsAtoO60aAz7RJ7JBD0aR47EQJ3cP21M68WyBuiFa4sQSQjDnEJJtOP
QaltQnRUrmnQInKOh8OahiRf9C/ygNL07gff9CEmTVuKpVEmXkEcKDfhzw4RTv4/
rqKQiSFca0JY90oy7FDnLCr0Uh91YtW9/fgPx8lUha2ghXPkxTHibEFpK5gm4g53
qw4jwF4KgeHX/kDk6JDdkDrDQBZFAlBZd2T3IpVQhnAPRcg703yF6kWVvCK4Ja1R
m5st45BbQJgqDRGyrdSbDTp/gcb3QAZOBt9RwSK4lcyRABSrFN23JIC/Ki2AnHfM
wk05Uj9Q+IIbULCJVHoa6YGHVqXDqxBtSGw4iOqT7N6PNkOWcyABUDJAouyNjM9Q
spLbwE5Po5Mwy5QvQ4iJXlQJGXjWE/5i1aPlTqOau0T1eTnuvQLEBeNyFuypv82C
O6zrzJDSq39U/VrIXQDSesASaT6eUlqocMcA9hNTs8ej29sWLHQ2zjTBoLWUIjnt
+D/TrfJhIr8sGXPEOeHrupvBof+j/h0GbUQuMJNe4DoGXV9n3Bx8I3NWgcbnLWmZ
iA/SyqCTwKomR2U/HvuVk2uIA/0dpuLmGp153+BnNBBzP3qPE0Rz3j70dZeCvIJ1
FEFWjvQrWXxKi8GB/E+bt8pZmob/nCOtupikRZnG9HJaQ4xRby0Vb4D7hrz6hfGQ
uyXhIPd9RglPMSc2xXf/POYGS7Zf/O/d/b9pJ1d9pp8+f2u7pD/C8jAWaYP2CiVu
t9/xX7pqFl4PKM9D+SGm2YeFCSiAvJw19hK7Qy1L/oeTZik1PaQ2pvSFutqLZ4aw
z/eY9vV+okr3EvG7cfe6QRBnSygJFCLvwmWi4/5g6IOLSgySgYDjiJGhm5vIUifM
K4EWcTd+x02Nsl3w/ZL2gFjsO5z+OQG9rcOtBC+6G9yL+ADfnUNnoEbPUWtABH4N
XZP4k7HNkd31+BbJG1FhWi92ffzOqbDE2PBHO+h54leLSYEnUYNqyeGoIiiZjbcW
uy/yBT3MX9R6AV40FLsCW6e419xkpj9MiMjk/HsANWygeyjIYhQ5mfnYbTF1nfBv
xk4jagP9KRUHCalrjWLpdjT/vyXtJ9MJZLxIMp9nHjA86qpmfq4lMSfwOwvOfbiz
gEvNJv+lgpXjlaN3hXXIZOUawCpSlDNM5hyVjIwf64y/lNEWPurzmXQZ7RDcBWS3
iez33OEiOtY1Wc0+b/si5H8HbsmGy/j3doZ8uwAVjZhMafOis8Ndex3/WuQEFR/p
rRzjI/iiF+sAAL6BoYP8PLSg4+HSj3j2IshDUMM0CmBGjTC1NmbOo7OilJHFh6c4
3q+wZEpWVqxBYk97kfkmlH/a/qrG4Q7PJdJZOqr/mVbj60fghIdIDebjJplAiMVK
/dkjaZE2usVvs6OteVozxwFW+G1ZBzsb7tqBJTOWP9vSxXCpwNktMttilCMrWmre
PrN6HMDVW/6+RQCCt+GqGEXAScyT1GVHXUxKCeXhxWS9HlHMViAuNLYIJSwD2wqL
bQPMcwh45XXFuzPRifiTCwnchoZFLe+zcKmbYdPo0bi52KDZaedee1ED2Q6Q9TTH
i8b9OlRNu6AJ+2hP0hSN+lOL7oXVPXnHDjWLOdf3Yi08bFy7aWbcp4YPV+vobIZR
dN32lA12kTNr69GNtZzTBkz3NEckMNGKGMNzSkxfsVmoTBT7MZjvDa7734rkmjMp
IfYGWLpZUQF0wF0be7k5PATfof4O57uYj0Y3r2fBTB+mOVSifg30KFfBmU53Wki6
znT7+SJ4Jt/1qHhJMv4Y+qJytiy9pyT1vpUaPjq71z47olN7lq0mQjb5t8yQ6949
hLQ4OYlHkkDskvpu+LTOcgV8nHn3EgqzHKCFF7NkNqVacIufKhY9LbcDC+YdiuoF
obMp8ff1I+bGrf35xB4eql2Xf/m5gBBU2meuJfd3IfvnX7qWukqbm/Xgo4IqSg27
eLyRZ+0ySdv5TQbDZ7gNOwnihzSKRtpbWS1/IBzj6e/mugHnzux6Qlc0qaEq+zSJ
hmwj4RniIHnWCcl+ImE3cJrF82FDTI/azUx8+aERsNfjJoBn2EJ9ZOzW4Mal6A4J
8fjRoodRn6MAS7dCACUBP2KmxUR+EsOne3O0XFQJsgw70ha/hEE6OpTet7sePrMK
JM3IsrXyefZntZNX5mIWXuDjuDq/ZoNpcYjYBIkOJ2pG0TmDoj0o/ccKGGtOdZ//
pG5Rru/Y9OWAcHb52BjRLHXntaFWBB22gEgMCQta/N6BiT9yg/VrEClQLkSvkeX8
o8CjZsZyM/fdYUaEiA9zOf4VKKPnVtu3HcILmIOCJz6LXypaAg4o7XNKj20OORNi
bOk9egyDbJDy5bOJHNsWhercZ6EkO76r0v2WA9lB93Haon/h5w0wAu7ub1xSSO61
EP+kWHwp8yQNbOma6krKp5Z7KZhM4m8pL1nh5gf8KpQh/8vrXNjOxZ9rncOEbcGU
xalC59m1UBJURguqYk8zTHVj752XriRllVTOBIlMlCxV/hlBKsRDT+fosC4ptIMF
FizzkAX4Ij4fB56TJqVzjMNnpy6lZQauuKLypXp/ppZiBq+HdL0IytpdfSJD2Ozb
u0N8sPnOfr+LgyM8jaCodx/ppmmO46U+TCLS0CwDOti+raDd+2MSVjIc0DPbC7Ry
ioBwXxw66ymSzn8LBuDX1/X+mvbzUA5itxjU+b47urSUnLReyoYk7TWe76WP5qmN
u32mlHRTe4cXr15u1wc3LASaY/p9qFyHLH4lItk2u4pcjGyeRIsPu+0EK0A/+Dzp
zubpI1YCSR3x9JCXsZci2QZTu6U/REr+5f8S9Df85RgeyP8DMmxDCnwc6JcVJ/d0
NVZo5wFhr2GVRqy5bjcilu4dHcBi4MM5fcfHIbne4xEjzNU7ARG7dEQAlaKL6iDu
7mzpyURZZiYRVIy5YfVCOFldYu28OcnLTAPMlzwAFjxwQYwrUdonmEYoVt4bmbab
2aH4Ob+XXiZqrOxCz473vcPNlz4ZwhbPk8Dfwq/cSjCR4SPyIEtxXoBjo1hUryNg
mtINhPkCPS2tbKHuhzHPn/m+UGFtaRRN+LyWAEQsigNg74ly54vrTvO/82494aXA
HC/FkUFgXDIm9XfOgLz6R0Wft3khUMH1MCYscY81yjOwT5sEMHODKrciK61jvRpr
/lyWPlzLu5ndISEvjbYXoKjzLV6ffyJp+X/BdQgQG2oOd51pjw/8/UVP4fsXhuSl
s4xs8y82irCYTT2G7+zsb15DgAvDAnzdc9pw11mBnxlMngIYYtZZJylwJAmGWAc1
3TflSkW5DxrsHcGXMNEkq3xOG2DX9UnGHAp9jeQ6y9ll9gKWfNrZapLnQQgchgHa
AunADZedoYws1TatovZW4r+6D+V3Qs093raDRYVOLoTZhrkM3NI2neTAwOTFr2MD
uPM7RdcAHmLfF7Kg9vJEZlkqna/2+Rit7IvTtUyRNdY2IEif4cKHriq84L1ASr72
3o50sawXOkBKio5nRDS3cAy87/A3Gm45wrE2Ullj1E+1sLWb07nw4z5YaAwb6lpo
fUVOZQ6WMsNuovflPU8Vp0eNWrKvoM2Qt4iWGnmWp4yH5M+9v28rmP+08t9ncORt
4QbKGZqsG02BCmwQdW25uTRXZmW2bmqOjX4Rc4tSaKFFyfdC38yE10cDTokttYEO
Ill3Tt/N0l7sZCJaz44AbIMMk5r11lzjeKElZiN6dl0AUiRytN6pa4zrXPWnJUL1
Whs3dLDM9sGj56mNSTwCC3KFFy+qiqmKjI/JPLs/CA831lMeuUV6w+ZpG77pUYwp
xTU/pGwWuqJFH39tPuKeMsvz70Fg5Blq4VjuEhIpexCB+FT8K+TnbLPL/vr4uk/S
kykAEh4MLGOWHyIXgAx7ukcDE3RSYOaG6hzZw4YYMoxkPNXwTPKbGrp2hzNEIwLc
/BUxF0pNxnzrFejiJy1XHafXnpY2slooBzLV7zXwzACh68ib4ylxVP7muKIRKMV3
/4xPzQgPoA/4denRT8LxN8RS2vC94p2g+lCna1dgog1/6h7Cb2+RE/8N4zIsTNgD
LsG80IeGJyof6HPmi04cx0sImfJlzfKIUEhtDxzwc9mQVZJNqN/kaY6HWkD4T+lx
a3mvG/L/iW+y1zvpwD0sI4bqKbsSzXwNONF4yianKldfsXfUcZ7GQ9/B+AF7DTy+
39TaBMuTbap8cONVZR58uy5WA/nBC3QNtZazrS3PExr1ChLnsuIE7VxKg+QI/j24
ugpFaCgW78/KgVZAqFjgWSBhOVTUJnshon0cdLKCC3PDPZrmBnHUGBrHodfcnNKR
Rp4vyerz4fobsG7+FEGMJrz2I1so5kL6S7j9eZtJwdBZv2H/q40PmdZll3JIPEOs
CKSkX02ZZFTD7nsgmk/OJILI648MxSHKVLUsiFfe2U3T5kmmPevU08B2NzSN3EYa
I1C/nrs2jbW4xv6Ze50QDVh1W1mnaE/cFId+wheM7Gz8SjiPqi+zmNeablAkrbfz
25nyDAfa642C6YKcZrgFVe6sYKW506zVuEFCEAlCkyATWFVPhJkFQsTyl0ycf9t7
fpvdNezBA/zIKP1SZ0SAvEDyR0Y0mv0VzF970RdlW86BZv2D7B7nkRynME/oE/hR
0/TbrgYBxD0N8TTV5xoRFX32qs/I/XIf5DtOro71AKxAjHmrM9a3Nu/zlXwIUO0J
SUjGcAPhtp0gvPMtTDVgZqE3QWqmt4hcqSrV7RcQmcXXu6TFKO3FCa7eQ6moEYJz
UQo29BTRoy5x3ydUCWttrrliq2hv1EgpHWclie0w1+Jaue0dXFMiAHHOdKoVSZ0r
NpBsdlIO0XtZL3KwNU6Q/KAU3/qmkgw7i4ly9K8EnGtUrzxVYHmeiuTXJSj9R3he
zClP/6h6SnpwWcyClt2x8qZQSomQRJV4gzYBXl4dYiGFtgUrHf6TaXU8F6fLyF4D
zlwh1lg0ez1RW5yL85DtxsQGI4XsLAsJvhgWIsBJl+Fuhx8tC5OC9UC6vBtxkNF8
gQe23fOiyNuKLzxvk0HwzVt7Gz8wZiJNsqYznJEl4lMHjk9c3cBgW28hS1ILFurp
4tzNeuez7jNqKlpscOYnQEDwxL30FoVHRpwJEB6uLh4vTgdOe3H3JP7p+99uTX75
9nu+mTkWAGi+5T6j7D3L9B5pasOHBdehcesi6JTV1mBq590mF6HlpQ5oU20Y1Zn0
LsiADRjNyAFjxFu4r0vwHLdMU7wzxSZtWuBcLfV13HM0A5DR/tEuiXWAmdcjNfHa
xQfchUAtaJY/n7RdGsOwcV7PhHdM6XYplPNghRUuVBlxMewovP0UjNTG8ciwt+vm
aVs4Ga4R0e9ilOZ3yF/RtMnYuAlmEl/cxsv7mhA8B06xoV5XJsXY8G+X8IIitDo3
x1ojVj8WldpR2cIgUzEuCvd0HDBtcU13Kk07BUoHg3D7xlb/CyQ5ycJctnU6gt44
81QJey7W5tDq1sYLvPwCKJUjFROgzQcGoX5EZs1iPHC84fwwyrGkKm3kv0tGaYWv
5Ctii50eRKO+WLLhozZCV3+JrGb8RXfjQOnFUDTjgXEuP2ZsoYSnwWnR3BrF95wm
tiEthx767POT9PaP7yM6ATR0XjPT9QWM/4pi/gaDijKHga0KHotLH5NvNXHxK4vC
4FKmk0tF0t30KXa1tA+E7QZqkeVeH6By9vvkDlohSkWEdECOzVsEqAYdmg9aOs2Y
mqhy1yQ6Muu7mvZa7BAtmrdVnql/GvqEe+5FI7I9kBsDgsrDg5XUfti3VdeEGCAC
rGRlddHOSgM+zR7nEdMR/4jBZAaS95HDgXWL8u3CZwnifOBDPfnctnFk2jRiE07h
ImUXxja28XOPe+doykkMlPuYCuW3+gUnzhxATl+cTXgwvsYN4Sa8suUjw6K6NL5H
d1I3SdnXCxCAg6Wb1JaYVpR7pJzSYw0ZB7FXmJSjzePIenkTbLJC6bYsnrjL8nWA
bus5GZjFGWrq7Lf7OLc3ZzE+9PNmL51zcFy7tz6dXrS+wHb6946FqaWW1f10xSLq
YKQ0wGtkewB9HPdEduNm8Mez/jXTp7ZSl5kfLj4/+u6OYdfh6yivMxb1HInhGSTP
dORBFllqwA0IYBWGEo5G88ENgyQ2DaWNUX827jJdWh/i69MGr32RBLJwSHvnGbv2
M5RHdyUXB/MWtq41uZcT4qvab75UvqfHuklcu8fiDmFk99733gROI107TvWwQShi
XIPJJaunCnttqqtFdT0fM7R67vBgoqZoVXogjI0lfT1utzNwyaTDeW53o8q47UvJ
98RwMqD3uwmbVlvsxewsnPDkAO6aUB/MLOmWR5ool5hYp1mikRai02o04980LU7F
N1+zz1EzX5qyKdWm5RPlQIx/93DPH9esz7UCOU7TuQJ2dmiUK2zK8p1HIv8qAlg7
/WO1yyIIjdc+Qq0nGGwoPCr38OQCi+G47e2WFGoAfagEdJMhVqGyNRong7ripfj9
xBbB1twHWO+DvA0RkHnrXfCWJXooY/pjVMAxM6VhXZ2erp8EjTUZ3BMbhrl4gxVM
b0xFwPI77sLFnOVTYIysck7nHMuOTBXXOHm/NW6qIsiVAaV4zyHzH2Pbpn7gODgV
AD4LD5DaScwTulihhu555pHo8+z7U1GPv6ifm5MWWmy/s1+FszTm6FjP4QIGAWiB
Cyvr3K11yOUlJKyQ+PRy77ECGYeWvYeVW55TSfLFaquGJA6rYWHzPbp6RN0qla5X
+t1WnAFeKX6saICFrLVbxGf8tTI3KnhvAJ4aprQtwxRQSPeFIJxtXHUpOh5dsBQw
wHEPOpRTEHg6K/Sw9aFRbUdz7XCD3V3duTa6IX4E4+ZxcCugmQTqsEZ+5xVre51Q
5l8wVbi64H45QgA+n7ZDH2lgnBbtFBsXTfkzGFPZCERXWC5P+OM7Keu8UpNZDADq
Q+Ygsjxejfj5Rsa2FV2L2Y5lP+UWghHMLRv5siZc1fU4ZludFK26sHcDuONPBwuo
j5chbvVxlSYSVvKWs1esmyI8IC0eaWfyNJyVEwqQJL9S955DhS8EJ66v6BoyYb3p
O+iKjdeAXQjNCiocoBBmvhyrNReAmWOKl+Ol6gCwDaiL3IlYm2SCEF/6DnAeJYa9
3E6IatYcKZOlFs6vulJA6p9VYtpV6uhKyqUZvTn50FseJnMjZGo4Rl81rCDvGc/I
jkrrFp6J1y59FTto5/1aQ0DVn7CxfeWAE8tjVgklUnzOpH+RW9m4q5+sdJNIG26W
C8u8mRmclvG9h7FwGTzb/p9fEXNh1nCWk2g9k+fd9hiNihMJVki7Ow6mc9NLcO8D
hSNhDf1Ss2zu/nSZ4GHAp6RMwd92n70YoKn5sjI+EJm9B6xUJNJdiPxArjG3jOtA
7IVD/pfHWBBpwzuA0HB8bDMOhyH3VFPCQSSHR/JIWfCWqvS8oGMXjAwzL3X6KREl
efIR/MwZMqsQwWYG9P32HhXm9XzciL+aqknr8T3RUZ40mBIxIIR9uKkoTjeqwQgr
DyuMOJM+2pQxZekdROULVs3eWcz2WCLmZoddKdkScSiDnBg2CafygcRB1rvZh/TE
uxSVp9p6FVi0NuoWGFK4SMp+PUUx9KfkceoJaTilHUerIXdm9ywbGRkgVJwzVym9
HHii7al2c9YyGiLTsC0FLUWIs/7SBtwQvFybI05t+yy/Ffah/uJSMHECO5brn7cx
EmEEh3mkzHmkaxupmURCbYxKbEjNABeTEclBf/v7E4yW8YULzq3ns4QGiuQu4V8Y
oJkrn9ckKCM4Ml5vCyEy1N+Cmd4QYXNgcVnqMHHjlRqJXsqEkgan1AnSvYHgQDPe
d6WVAj04WtEJkAFmyp17/b78TOMcltXJ6lHcHNtkh/YMnthx/YC4a67Eq1XDhTrP
eypZ/MxYiiNQjWWuGGmMBvsoezs8cRpJK50BQVPyDZ0ETRceEbDec8i3w1BOCk2z
swDtg7yK5D71t+sJSfm4qmC6MVdrEqpzVfkdW54gMmC7vb77P6C/xYaH1qJzj0Rm
PRsSPAdyxLQC9xeBdsGEfXyrRT6vWLJs0mATHV522BNX4oghZOCtam1ZD4ZJDj8y
qZldEH8khZlmsJnMZogdLGOLnpDf0cniHZn0xNMCFhwErCeNotN3WocMixiLG9pv
zOCldelMqS/J/vqdgMwFaQml1bmnTAn76+lxbR43+AfwlIaWfyJM3cSUwKw1dvZp
jll/g/PSJRFajdW8jA3RL0h7zvVuRZdN74C4ae6pp/GZio0uUHIB2wTqJg1jdqrj
oWOP1li/Y5mXjck/etBSOMoGTKuC6cyIX1yJ4Vv+kI7DlcQV/gYGNmG6y37eNBBf
O81BxqWUNuhVuet2X8iunJH5lVySf2c/oQEGD0fPa8CVIFM9AN7IESXOg9Jb5rj1
MOruvn/GBqQWE+pYpSbaUxoZaPg+TxXKHjCZ5DiQoyYDrBeq2/PSVmd/cEF+hgoP
lN49u9prkuXCtwKPN6bRhvkMLR1OZza+WfPWiDpO6W8qo97nSA6Y1nUHpzxPRfI4
pdhcwiZtl45sEO1+6nl8iJKh6oyY0ekYvievI4ntw5HZPE0PulGXvRu/QLXeDTAf
8Uh7RsxCKpQYaGcbm8XRdTPk810X4KjUgnXsLGrPEkhoUk31iwI71LBRwhcBjNDy
imFnh1EbsNOv+B7wFJi1pzixai6qRO9KF8rXVTNubrx3yWshPmkyLv4w8HVZFd8J
4SDbdCNvP+Yvm7HMBW4ccsuT0mVCwZEPM923RtPNAFgI9RaFDMMcs9/yFDKBkhok
FlIye7zJw1jGLg+XDsjvKV0YGBQEydrCJ50CEHKnOmqFuZ5pjpHLScJ8tbIwFOW9
AENbJpNmlDmsJ7HkAv6Ylezhs1EhDuwgpeCiXsKZvjt1SPdj+4k9P/14VVqAuIwW
6vQLt/kVg/cQ540PsgwBnk5rZnxfXr6XRf0BPEvKMSDdizUD8PW6jR3gkHMxFlRp
p+7rMTvhhgacnN5IHyvISqMh+4yGTVN4QL7QCgA2sBwLIKnry1qP7DbIKc0iXTpt
uh0Y/N2zGzMA7cqYVJFBYNXurR6qh+0c7eZOevV35G/h7otBK3jTBkCn7EAAlpX4
LH4duc2vTWM5q7gxsQzkGLBY/y7JChtgXqu6dPCgVegajR+AmoM2EZBE2Fb60o3O
Ej2huY3CTmit0DsNGs89KBB6toqfGntdASDqNHo1339bHkmR82PZJsjK0nwUdLKE
d3fP31vFiaRsvuDRjsOEufWpc7MTrKiJA65z45AbryqwsMIPHp/8XoE+tyVYLzqh
BYn/JGglETkYvCZEu69lQRbyXZQ021gu09biXwUmg7AAJ4Ss+S6POSyICzBW3+nY
pLe7uCejzd0sRnZGJ3u+GULVrzlawF4oH0hU8hTcFaa7wbbclFl2TmRWFytFZusv
Y5NFxfedVnuqHedT04QWCeCI15jJVErjljtJMZqwmGmuy/GYJcDILHEFHulbPzfT
7PB2Q654i6wW1jRl97A+jzJOtOClwtQQKb54FHta8eYO0Cdrz/BiiD+RBqixACZA
yQThaKD3385mMh13cIFOh1Vn9J3KqO8MryUbaUEW1mP8Y/yqTmNwd3q4KBjhOeHK
Vz3FAwqrs5bOLgzCT6grwhBhxVnJjbw0JM53bCSRz5JBVxNd+OW89DeGxVQBIVQG
1m4Lb8J00Mfen7A/f7aq0RkVgPAYOYEm2JARMGmNQqIEOGjsMS+eU3yMxbgroA3m
k3vQ8Y1ICROARUc1m/UDry5evDt+bXShozh3GFmFDv3qi6MuE7u1+ivd2p9w3aLq
uQKe7yeoVrCqYB3GHuUgKhZQ2VQ+vmKo81hQLV9Z7EpfS0l9iRjDqsJ4hnRYRdx6
WxOY2y+Yth16x1uTI/Hj2c78ET7UEd13CUPC9mxObSPNlfuHxZiD8az0GblSL/Cc
9Y4eQFvmJDaOF52Uv8h5CsFzQyTVScXK7DwEwmskf4fxY2gCFQAyz3NSjvthlZkc
bf8mLq0QPRS7Nb7tXfeQgb0MMOz+6RLzc+w/Gcu3lAXwugbNdVOxCxNy3sEqoapU
7FoVq69G6B+ubvA6f8kQJG+7VN64VxpsPn73vAY0rv7jbBynj2rdD60/uErSRXV1
NPhxJBnY0E0YChr3rkWJv3o941hsm21av6pWHRXUVrMwkiAfy3HZVqRdNIK6RnX0
5rwb7xW52bNcmD5wY6AQviVoHFmCxXzXzyBqkWWws0VoSW7TYQMqrsK7V9fv6X8o
z7dkppmFgQXRvfRLfP8JDNRu0Zm1OqWAdi9ioubSoTXllU7KRiGpoMSyCLo5gBgc
Q9ljDt7G9Zjxdm3B4FDTPt8UWalURMK0EnNHMjRtE+RCzTJ84HfTs5QqIAGiA6Qa
RpE9fmAbyD+gkrlkTCK+/AyJ03HyHQ50MVngitAgw+GNVFnLcyvMq9SMyugq71Nj
SSntih8OzpgXhmGyKKlY7q5kSTCQUvU6jDYMri4jDy8UZC12zffMNPDMQAxN+BGq
GGiOquE4s49wiFikJeHVycdvzH8R7YY3lP1wA+IK5PvRJmacCYZKvT7bXY+C0Zmw
/WlXppdGFDQgl+F5lO7Vg09Hj5v8/Tkj3Wlfuk8mg0aDkuLOzZTIbCbNudyuI1Ej
1w1xV6tcPjq8En7iOp/1Fhy+Px84DLVWLCSnghstiDw0lnYS5KHtc3EEoDLwR/be
2nZuYjrn60laGKXMNDJ2cyYhZOChjU893MN86diB1BZW7sh4KXIz+Ia/1lDNH5Oh
f1zYs43PEqVYDUBvzlJgjqsRdl5wTHC+XVKPovwku/SzAHlelfC4+8YJOaO1/e69
5hZzoDaCjJ1OOOkeLgqsfC+S27PIuxF/xYnbCumeA9vBGiTKts0HCtXSsQUcMq6N
SblqFO6xNYgGTGRQ3WPnEaU6cHah2t+9wHdTCpF4W4Y56cidtEDoskw9aF9jtkUi
LTIw2r7mOxMLs7AdFXo0Ld32KqlgOBeFGzmpxI0sLgyB1dX1oqTITgOyDLnn4PHq
zm67e0BhdASm2p50KyNbBeZUc2divzSeFEynalS8pcaaGKKYTwVDi4K8OuLAGL6/
G+XksYQepeg7Rx2QjD77WITk8C3hmHa35maJJ2TYA/DaIfVcR9BTnihM55eA9WaV
RD4elXYl4Crr72y4Oy55WArpGyAkeIyVou2fIgL3qAEQvGpQFsKSowB76RSLW9zk
c6/Y+cr5ZhqZKvYw9kzmt+0kP6Irze6PLXjDin+ZAOFmPND8c8oXnMAb1IGAYkAH
dyYHwMRYxCjgXcUfw33G1plXcOpvssQL1oK6bTXZT0hXA5uFaPEU1Q2eoT+p+SBS
BLxHkItFcWafGPzLXyZfy1IIyKsdGTQzJcZb9NvJVt3YTR/KKp+TzV8hQNiGwovo
ovmgxvIUloKWq2rrASLovohIb8iG3Jm04DmiG8gmlRwhD3SfDWX+opdeWy72QIhY
PZ89BTVFnzjq22eVIE5G283ajVLvlIJDjgZCdedXQXI+tFR0JNHb8r+HvSJk4dSM
VZVy14PHyzuDeg6VCgvntV35ruG3yMJbEA+HD3kHDwK8bVvcSEqV4p29a3DU7KM8
UaE0E+7w6JUfW/39BeQSCcqGwfXfYpsCa0wyTxZ8r4qDdvfPua6GA/UlUJudeDgU
hfHDJoTAHb61Yh+ZmY8xKKGkJ31dUzDpPPYaMdcD2dwnnLEy10QCI+f3vmX328/a
HL1GsSSSx5yg90Db2W1glkdEtRhDEQERBhsKsp4BGu6n8Ij0qDWepflFyQxFnfIT
62t9jnqYkjFTcVmRxn+HQtgsaWJLf5jza0odos7WMGNPT34RdgdsHzZAPQw0qib5
JctCNPU1u1pll8wDnjmrrfFeVe8cEjCsK6A8tC82RB0UyK4cOrPnVI7nmVQOsRZo
+xGKFaqozGgZ6cL0GWmfau4QfkgpMhUzjKPyJF/T1b/Tww+X3weTS+8joPtBAlER
dV4QXnKRmCOs3Zeq1UBKkIcmvBFVk1ufXKW9LtqHk6heGO6JGhdjh4qIbuzI6e1b
PzJRsNAODHuxxY8SuSwpFxKo2RCkTUpmlA3rVbzmSWYA2+pcYbTNdvN9a7vOnGWt
pFGOeqRML7c19pqZcbXlDLRo3kaXQt8Doz2sSWtvGzHaLML5r5yg8UwYN6/iMtg+
Neki0yaQ2vmObLj0b2o1N+b5OFXZjn5nq9OxWdZSCp1Rao5v9uAi3HG96R3OOYRM
fhBSMmJHY5ihi0ZbKyOl/QQs3EbZdCH3eBovkYrGAzydj5MjkMT1y8IKOxK1x/B0
4KERWXck9UbHxL+Ji3u9sFN2oMX8tz4n+VmcZMDFbRYnQyZsqfQXFobBhmohY3Zk
3S0vtHat4/fJeiFWNIAhDWr6GeG2U5YNhZP/Px0qUoe3UMETTaU3ll6P0+olGyau
r7fi0UucvrQS0kIdzSkLbXMmCoeIgDYnXMLP5NhdLQukz/oix8TTHnHD7yfBehfe
Ck/QtRvC2bglMKsg/LeVAK0NTutNqmPhp6U76vME9AIk/2iAWXA2T0zQTwzJI+ef
hitahTSQQ84dNwVpibW/M73YWPtMhZnoCiF9srN+NuaAmQervPYwuIU9Uk3BEyDc
Q+sfZsNv+Jlkc6w1wrrithRL/bJzzZGNB0cIDd4W/gkHkEL7NxJNNi3iQck95f+8
w8g1SLasLUFrpaB3QzkaoQUZbvxKog0eqxQjHeIBd9Y+U9Pij19TdA98CxR8r6d+
QcoanhTi/B3qpMhKHSQvOO30ML0rLD5/T6zRhjeAQ85otGDAjhZidmfOUONij59r
3A9E2eRDfOqKzXRUF8PEcOdBfTzxvHLAQh1MKAfKwZlbP49uNaxhrXvODbo8Bs9C
Q1yfvg+uEiYS2Oj/F6R1fKB8Ab07F8vv4gRqDVa0nSwly5dagKIa/wXbMTvDUWpU
qbUPit/8T4rAxqeanz90bZmBsAlZ4pl3uSICgfZwtSnRyVUpk87A8GchxiTadDeG
6jlBip4U/KKA7jAh9qa8tTn2oJYcv+mlAEC+q9jIBg4/CZoA/KYNo27BctvFjr08
nEMBLXN55m1eUExxuBVVayuLUOoBYCl/HNmGjfEjA+0QKMAdWNFwGN8Az8FpnxyQ
VURFlOgUoUAhKQJxpxEyDxmM6PUFgAHL2qABs/WPd/6jNiJKb8MY/og48TajshkH
qhCNz13iosvr6rM63iwUOz1Qc+q4uN/7ylqt2vhKNs1p3xq+KbOJ4MHIUkXfiQhq
k7XUHwGJG/tygMdnY/3b+yTQyFc/QjDCWjOS1UYKKFrIydOKxF5GYhQU1TpFsLM4
giUXs8xOvRvaJq58oGsBHzhZQqNt666BrRLBLYadKcG/K9NcJ0JJTk6OKqOGif0X
RSyvt8f/wUq/EJRFtKBYq/kCLGw8o1zrmO+m0Tj5cAQe3PCFtHGIal6xHvYo1ml2
LuF4I3hmmhviRucRUIg1JZrzo7Gdblof3BaPfquURxy9P8De2Bk8u8kRnZJnN2MM
K7T1ETthGSs2e2dstT/Wv3lTHKLFecHJuW0O2C8lcLw9J+KM7EdFfePG6QKnVbM4
N7icG+5G82BpkEsx5kS/9VrgVDiba9DqkFAYnOayxrN+Z6c8ZR3jOdkLSydK0m4J
WJu00hVpK0V4zBZ+4gMVwCXZ3eUBXSL0JIdtdlmRmHYVHYfBFZ+MlWa5H0EUuCo2
0fTPsn1Xq3mEVP8GkeghSoyd5uYZ3Z1HkaYhvLwe0OkYk6yowh2GcE2M0OusqToR
/L5vRv8hqjFshq9QwM496TvyDoBb+gAqzZKTHAvNWc5o8tLEP/VpG9sR5WQ8/3r7
e73LEzKDbIPRrZ953W9SQt8BPVARsuYswFhStTkF4zp7Ur3ESkAONQhmSzyReCA6
vj85NrlXWO+jSyabMf8QpcMbK/G3l9GbU/sW56Nt3KW1Z9k92+J1zi4fPVUd5dG6
+3SRsCQADWyaEJZd2OlbPNKWPoi4CFg0Q94kbBdRYaoe6HRoO+jhKd6TaMpgAPMA
5vYK2srgNwlAKTgIAP6v0U/jUH+rOHs0D03cgvNCIsEL4yJERMxLWpl+nQ3Y/7e5
434ip5PBFeweXwhKYdEDPUBEcj4JzWkR2KtRX5ptKKf/seIySiKz3v3NDo7uuOm/
+2/XI3eB24bMIwaYg6FAcwDSYT/SozW2Q5lgezOOaymhRoClBwkp+uqcFFF+Gdu8
PF0WpBoKDHU/D7QHA0XogJ9o/2B6tOH422uqS3k5Av8g/k6EOf+UHFjZTzPQXaqj
NiivNN+fUfTddK69WDdRpZoRArZTUoMRJ8P+eeY6fcAEPjk7fsqMW0ikgvmwfbZ+
M/91HZPWKJocU6XqFvOOjOSauH/YK42I9Wf1m9IEwjNWAzUJHN5azZYD4EaLDm1a
96d91h5cD/0O7IobltJB8i9BonQMe07fe9wYzVcDMo7jtNO/yrTjmTR8j1OmQGAg
mKi7kyDKea5V11kz4o9ckA2M+Mz9wsWlyWbNJJ+vgyYCBFcOMuq71c6YI+RaHeYY
osp85bUlBZzuN74BdedeHgyvBkoMgx2K6Qu6RjdZim6l3KzMDgGX5/yxwS/ElVTn
9dOvyvHZHNbZA/uVVguXTg6FkeD/NlbR+0Kx6Poo+kFeduZU5C6Neb9Ax5mGmvU7
DAONj14btFk9nJuDrgL8yc81aunfHyF/D/QVi/qMe0VyaEsoANkUPDAu9kGICnRW
EuSHS0Qd0s5oJJpYaHuzlDzs7+QtVwf/unhqD+Kz2tIDEtVHurBoFF0Ge6WDsAVL
+gFKgU4d5ik7v1hdoXC3LQvw5srePonQNcGav4iJAJi5SQ5rhAHCN0qEp1CtDrno
Q9/0eTuBnsUEhBpXTeH296A5TeObb4rBsJWT62sUnDhWtceSvdLWCWim0JkvjxoS
hNQ32EnCGHfNO4j/uC/DQmrahCCmkAIqF5zfU1FMSUIEjmOeYBH3eNrqY35bydeA
qtJgu6O9dUgvh78mUkMM7TKjeK/Q0bEuqQkz9QKadt5uhYca7elW/YqdYEPXm9+X
PXWtyIw43sPvSBtXSn5XfWQa+TlH8SZBrKbTXWI3U4msjUST454+FuoKkjtqxZ8c
pMKi8mmk6v/vHp7nzHrIhr1TEiC7nMcrMafbBSK1d3/vZ0exCLbZl1Cj0y01z5n2
LY4Yb8hyku3Tc7t2YZcTe4vllI9cioCrd4hj0n2frXqABFRp9D275JgvnBYazQaW
RLws0z/8+TjORPolPxa7NvGC1poEh7HXPuTmxc/VukR4telxZU7Qk9kWmDixZJ1Z
/2KXEMm4GX567wn7Gop1zFC51yb14n+uWzvy6AefWjU4I1ULIuIRCJKYIROpiZdx
3t8vHEyLf0/awiSxOS/BO3ixcxb0Q6nSWznE1MnZ2Lx8DF3U6CbvTKzCf43iozrw
Ez+XGIuvEpR2HkMSBzkZV/7yHxlwteRLTTlmOKgjlLsnQ7mJmLbKa59hAljTGZ2Z
cTynGpGxVf/00fg0I234TV/IbQxePWrZSItetLWAI1RZ1kB9tciKE562/xuRLUtX
M9HdAh10gWSAeJtf+DJTkHK0WUp7SLfDGeJKpTqZYuBp+Dyr/h7B+0+D5vL/FS35
lnabcx++EAFD2t/95fU+awulsMTRnIjohPQs3d8gbLnGPVXv7R6IeiWTP8EQrSD5
J0lJ5kdyLSg016L+TfAwC+eaP3IVEQWJ1ev5V9m3UqC6WaWKIQdqn21EqHT0N4jp
inmH+bnS5iLfHBtGy0ysSGGe1ZQ35yOq3ahLqhd00scY9NXyDSSBPJ5EFq7FsT6x
fGLY9VS/4pSpWQCYqFbSZrGc/tVIdxybTaXwEgjWQztA9+ixZFlHSE02oeYxpNEe
ADjB9X/NKPmBF+dCxXO+93baUHWoCRBmsiqtim3scOznx0gspT9oU8eKgozRFWzT
f2vXw7h0yVlo+PmizKKoY3F+9hLd0RTV9PeNueXU59UXINC1yqWGkF4YkPP1iQKs
PtMKqyoAwtJawNrGvl82VQUOfDc489dHXzn3qnlaX/lvWeX8taZ6+hegs3ODHpR+
IXOnlHqmcfGJ5sj87lvcCzdBe3rDLQETp3Dg+UQFlOHMmXIAsUCsTNWcofyqW6V5
bv1MVa3goH3pwl90imshBv1FagirqCqRyTLxiVwY99lLtTT4pX3r+Re82LltR3Av
IvdN+EBlyjRuPHKDGtirP5XgCyN3Mplmqcaneo8gP+L3v0ZL+JnfyxslaF072tce
ZaQ25W4cUsQ3y8PvDggOdg5ytUK2aSJJDEVCBPJizgkmq2rAY2DoD38Io6Tv6vo4
IXU1KcNCvaB2gN1nedkLyXuRBzLdC3bVgb0Kp+UPDo7Y+77/jVdXBnLQyQPiDnKQ
TbDnnLYDz1sjZf/XsITC6wipaLP1sgOtYyVHgUt5MGnAQ7yOGM0KSq1Aby+9QMZk
nQzZuAjCLCjByh3iJr7ccg2Pvy+BtF1o3vTw0Hf9uKkJt6lOEd8X8VP1PEqMmSI3
76lgfguneHv/V6hE6M1jH278MZaKOYiEkTaQaXcBFyO/aiuRk6XSPYZkB/hAbRZ2
vaqJyWymSwt8QxkAKl1D73ZA8JtCpMo6PGLrt0uxxuNJ6QfS9IY0HjKvzQNEM39j
lT01xAtg2PlUTczu3owVJoNDK+vv4ZOi+SD3DhUYLBm131llTGe8FO4cb1AeawsN
VjD4F57JtwpBSdCJZ7s90J1KYKm3Z+QZcw05u5YnwOyxDU3cYvRL0+dqEw4tztG3
AjVZVpbiimNOGxWFW4ZpxYO4WQGwG9t7ULNshATRsbiRF21Q4gGbwOiZN5yDWnPK
xOJ0wNTbvfiWbJgWFe1nbX//J4jAiOlQgYJem+KgkQXjDxKZHvB4xBzbNj7XnMkm
JMxI9w6Y4I+meTC/0GF8jMSxUAoR1vAwjcgN8k5bJoNK+/x5JovQC9uM9hBKJF4E
G4FpVH1ZTE8ejby/DqSZJirefBe1923KgX93lVqIuzkCxRbr5c1Vzo0ct/R7+S+p
f1XetsGZ94p/+bEfK0dThouX/vp7KOmnB+ZJRsknrmF7ZZdMvf2i54GENclsaTPt
tvLBZJzAmNk6ucorX6kCmI3oDX2Tr4Rkl+3vT6Ao4H2jAXf4Qj+2LadTFZQWQdK2
A2ODoCw/1Xz+h/bbGIA5BdH19vfEY+kivTp7Bj1FIECEy50JA7o90mQMj8npoi1V
KneIZMhlSR7B2P9MFB24fpG5SE8uaEgRgebgOA2vSm5UkQckgyrMnqDVSbtyBAse
xO7G5IluJ/KfLI3ZT1ar6wahWdOWY1jAEsRuuyLW9HzNfZsptb4WPgjOOnxKZVz4
zXSecJ9lD3gagMme0SUwugbVHH+MFMAt+r8YkQ5IJGzC3OcfOEwJWqHpl+UZscY+
j7gVhARRy8oOYv5b32oOnuxyL/hLOdZtaTf9CFrixEseQ2ltZtywjUAptuJ/SD7t
JgJEXWBxfmufNUQpE7UODYXCKMM41+p13ZRuL9VG+i+vqaP/VhaiQ1KCY/rDv4AI
dkX2UOb46tvrQVkJBgHgMT82zdsAXXDr4ZyWZJwjWPWsUZ1kRa1tUaZ/k4I81FnH
dP7srjoDKeba3ELUeECzwPoW773YTwXSyQ0Kal6oWKbUD7FLb1L4ZLPw3Y36/3bP
3yWCpFHBIW2cW4m5praE6WwH72GHt1b0YXejOOnLln79cQFyl3V057t4oP8SLsYw
wqE9nFdFycjZl5z8K7ZG21Lov4t+mAw7B7Bb0R5qAlAYHhtvA2cy8FzapD519gK0
4pZjBsUqy/bqOBqPQTMWqaM+/YEJUWDcA9NIdrD6WWqovhLvGsTxs9G+8T5IG8za
JMgARtjE1ooX6BFdIa2Ew6vR6Fc1mS6nsJMgRX5Ugkl8f/78sXXZ5vuUE4XIF9R0
h5BkxMz9EjbfaMHvm3qyROoDYmivndl4aJHPi9Yhmz/M6jYgb1pUD2BtUT4cjadA
thUIHqOn04vtlGeNW5k8wzd+xMJeSbwZ8+UiMvDwuSfMvgVSd14vzq38qxJ6YLsH
NRZqY+MdQBzEWnu7jpUUPhSme7tnspRzcY3/B84desCKhBsHaF5hAuoQSldF/jYR
E7pJC4PhCk2WQ9K0b7gPQNTv1vFHuB6KNmMFrwEptlZLnLPK2rNZRR3+CImOmqDg
BJ6khKGu4ZOJVckPNR/QfbNTy5ZCSKQv5kStfWCUffGiz5pbYbKh9/7RodQ1iIha
9XpLIA7S1JcH9KxgMz30pQc1y+vY50yAPMTryTXNTyQF2TUMt52YkIMvxqev5nn2
Zye/vUTqcXwRvjPl6NjktINgukcfG7s1/hHAsmSPfzMMzqY0asDlIsqksTPIcWt/
h7GeopfUM8NQHVUSOBDfoLNgiEM3yTXZwfzH1GliFjSqCLoKbEbIUErgoCelhUy1
sSFCOkEIepWm39w/xUFj0BRH4Lsn4TqxhOfnALCQ9ukWk6j4frmjmYQK7WrgphOq
x5cutK5PHpGct8JTZ2hG+0c1OfgSxpjoOgh7iH/1YHFKE2T14PAJl6PK97f+/hMe
H+StUfugZ8Z6kWCWq01ZxZDQTrYS0g2JzS1CGK0rThBMhQ5+lgyhSodA8vl3LoNz
xRbXAumw3ZVtqfIp2Yd7B/7hQua3jwiZdglJ4Sb3NPKW7v1xoKx0Rn3y9/QxRekb
2deY9++X5QwT7FWDCHQE0mBYwJmaNgyAHDJ8vgzaYxOgouEzaNSlv6ojarPx4E3z
9jIqfHkx8IqLsGA9Wk4saNWQYL80BRwnOm+7CX/y64uY16JO6cB7YeI9ecDU5dXE
0zfHSJocT2Nd/aB7EK/3pa6oo87E7j+MVZIkHcSU2vKk2sreky4CMB/PT3+UgZtm
qu28ggAa4QSFouYApsB/dhYN+8hu6JzCsK9TjJ9rPR4PzDdmt1Ouz2MaeDe9IV5N
usXF9/6ug5j1nlGq7v6ju/GXqLMe3VepB7h76F4Z/XnkkOFpd4Wl5sitkcQDRItf
ixqgZZQfztUoZmaoLFfL5oye5anedSWTLIprNTGuqXDUVd2XwNaH0AikI0pochLJ
WFr//EmDvUOWcd6exYlmIHUs+O56rFIIffyYZs4YRSOV7R54fEuiVOh4x0uvSodr
g3JM45mppzdlVTFQ6YvzWcI1xeXdqYhNYsJx7YJq4T5BxGYJSPQQ9jwOGXMLyiLW
ztBWGEzfRxTzQvY+HxQ7T5O4fo/KWAOHGyC3rI7w/0o9mUNISuvUPOF0y21vihLe
AnK3/3Z+W4Iq2eiQJo3M1mwyMf+qZwcvz/Q3GGWS62xltw8WrZicrGG536tbzxdQ
C2do5ZNYqhhRxZDs8RJwHozpMyeWjxZQjE1dFaBG7pCqq2TBHcedligefiFfHYd9
KxlXh8JJArHBwy+8E82ZqSL9/OfbrTMKmdibfYK5eE7bYMRCTeJo5jN7b+kukJQA
dX3MkQ1Cw/ipxULbyHX5xbQ/KfP8pe7D4uvRnfXwtnWtDe9bpMRP/MUj08INUORl
NPlJx8D4pJXWJFE9DhjcuRMbg3riQi1el04frJ9fnX8gcVOhrd0BYDl7/fl07c0n
QX9QhxtNCa11A/2c3yMmw09aEMTRKrYwAfMDVOBPRNQY6sey3Vz7ioCh3BgxAo89
rnZhtdQp25f6EAkHhQrU+lPhV09xQPpHGXdJoL0647emuWxI6DbDtazg0/32IDIs
vcUhAsTeJ7Zc+Nnsl3hUk9MkeIIWCjasjxpHznJ89XrPRgcINxP5wGDYI49p+v7/
al2pCJIL8wZqvqzzvYFCAQtzLLTTb8jmyHpuGUQ+R0iCqj3wdQ5lTz/JXn0QBXDR
seYGxVL3yocD5RPNygqt4uxYhiE8Eb7j59cnEWuQys5PbSthR2y5orcPpw8cJ6bb
JLzQzKyH26jD26B6be4NEXAtUUqDyY30WuUGRmTwNjbR95J8nnvHEw/Zvi1kHK67
MGewuO4neHLoJb0qBnpXZPB4BS5VhdyVVBWn0vbe9p+p5luOPPlYim5Tmi2kCHYL
aazHbaoZIOpsuGGEVaRXDzDtrvyrM7sF5vS8TwG354q0uK3O5B4nkLP4vNJ+UcHN
Xy+plWMS8OpkfCmaM3/4Gvb/Y/HReXu2ImOYGbtwyDP8VqAOnUcYo4bCerruEYTJ
iPOzTKPPBlMypZSytHfk6pwbYap6f4eCrg2nRlLFWPbsSLreqt0ydDN0p06tlwz/
Fgdor+Je2GD9lpNfGOJOXJs2AUghcF22XLSxheByw1eW+kWB8U++l0wDrQKYabx8
XRcRji2ESvTLHDwmcamSAHfv2G9tHGyJ3Pli5tAAsn+AHzk/8/XeiAijUC2eA/XV
1y9T1q0o/eGSxiPPbmyZXFZPhYGVij2fgNYkcajxjBeALa9c2RVgQjJkuEgas918
Ehi49+Kun6+kQu1sSpBCzSVOaapqtpgHpz/2CWYTgVNKwsrq7dKU3Wx68QL3kQpj
SPh+pL+TNbtru7XZM+YnViHjRhazxj1VKYGIAO+GTtb7W7mNkTYTZB1WW0jYuQ4/
C2T9HDPo9xd/FajZQyExTefYdpWdKT2DnBCn7XxBbiC6mCNCBIR4rWBA1ntWB3yx
+TmItSe4f5bpEUXl/ol7T3HVwr3cjPsdW5Y6V2OCrHMPq73ZRdlKpjcIBSQ7UOvz
e44fuTAh3Fh2mh2XKh58BE8uaCNzYFNhONHwh98il7sqbBid8PTddM8H8yxiwNdT
jPW1PKkCmQZL2VRYi8JRf1lVxw8827liYgRxmTX/EFvBrGjsOU3r8TvY7t1oBMzc
FjWcYVOWZmDxTDQSxMcbLbWL/ZuyqcKSs802NZjPZa8wZ45+CXX7P2jjNhz62mTE
76Av4MfPT1zoV8gcrtjCWlL0xZSGE8fLGFpyn3gZf6HdXvJSn81be7Hiap0KmIZV
I+iU++4wkiVP/Rq4oXSc++hJ73Y+YK6r4tnBlmlPmIrtP59ehMF+BjlJFuCgyzTf
FyiKONtU1bDEw1OggXFaw1n8e4Vzn0uAgCNjZ3waYAbpKuJF4hxqYqoOqL8Mic9w
K4+omTbXzFWV/wK8flr7GROlPD9oT7GNB5PsenKUvKfGlFF5rnMIrz3LcB3pI5cc
kB0HSvN9BTpXt2W7caGxze28D2RH8a484GVEJHO5W//6EsifPJvJpkmVh7AafJHn
AsMeCA7hFIkWbpv1Oh5jgltHV2QvrevvnmM72Z1o+pDA/d7zqqvQpfmFRL1mjgBU
RdFnknaev5VTxlXK9p2V/9GslxHonccQhj+gsDdkHaCQzOgQVLzXukbtBL2blCw7
HZaf3oD2WhTAJqf0gNY7oqagPHeIhFm7ZUXRt/eKHb6AqO26sV/0T7JBwWfVFM1h
3nI5QD76LstG/cWFzDoRw7c+CRspbjRST8YC6+kQg7cSEOrm9QV+ziUgZ+8Fn4BS
p9YAGy27NLhI/W1Ib6VEEbkFRmIkTHqXZzWsaiOHp2VSeCkvhVvRjx5Kph+KGJtG
yESLN/93tC6NxpUCGXQeF+T5GM1SfDh+s+VdFtljVmAkvqvypJUoH5z/ceiJN6NL
1wSLKDq6xAfIEqtDjJlUysDTHBRCUzXy0qOq1qrjhSmc3qfaOzRqRERc3snRkInD
mXFOy/YjBetbli+OvXDm/2exA0woEk/JALPa0+I8mqoqexHJUti+6efvBnbDj++S
CSAc5KwrrJ/K8365BsRWeQciyx1BdgwbIaiQlEDjfsWbrFSn9ot/wpfpsQJ8hOhl
3HMt9jvUua1IWGEwBG3O+NqCD1Qvc45rIwAQ1bYnpEuNtFRx6yFXzkkAS6U6jcnD
PcLuDweu8xHni21gxVH+fOVFYxzku+5FAGTyAwpEUKoVhmrFvur8i76NfDkM2cul
2y5QXRCZWEsWfNsl2+ywj8RZj0emH4GVfjHgAK3fLnCexiR5PYhFJtpXdA2lZO9G
Y9JBCAO+KNOLzaub623vikMswNeu5x1K/EgwkxbA37GBg3B6mY9TO338S13NTnGa
N90VmwSDXEx7SCHXncoyJCs8pblbhL4Mucumvn1y1OnqjHWZHQqL/lSyrZXv3Noo
GNCtINkIGSoF1aTWK8LQbfSXYpGuc+cZLoWAbNmpNQltl3GVCj+yPqVNrnKSEVkH
F+612oGMWxIKfyD1fty5buS4Jhe0jalUCa0tvPuwK6bCbsKQl95Oi+g2exUZTpp9
OwsXnsokMqC8EbjKczq1LCeBnVMZVDpEcL30S2Q5jE3gFfBPmSub0bsb8twxP/8n
i0E2vKbr+b7c//rR3nwuJQft4KBFq7Uat+5g1MsPL28Z7aq8y6GQeKZQfnS6GUVw
E8tkkqVOLnjGwcgxGoOgusHnA3LC1sTQ7e/82qm9wQeb1NUfRoLlCue4GEM/rDuI
D54ONexAFYhqxgu9BHd4e8MUjv7K20oaoJGLH64W2aDkrIxZKY62lJ1fb9xAa3l5
2ezRbn3sGESTX8vch51TPyJ3sj8bfrYgioCfrT4LRa5JXH/FKyRPfKwc1Eyd/zIw
23eukb1yWLaWogSedz9p9hoWBbtsFQ3tx2WQbKarjKHGy1lRqaYbFRLW8VmymUr0
9h34nAE+vQmpP914xvxv/jZc2LoGNB9QyrZEn6/U+jK8tg79NMaXuPtj5YHmue3X
xVPFWYpOVDo/IWEFJBbRwk+XKgre0kr26wIUGbAdUXyy47c5BqPLej24m0QA4jcn
KDn+LVvy6kEox9FOBVuy776zP3Fnt5KyoXciyzbT7g2DttPKzzqq0KaIDOzRdCpZ
8bGHe6YqX7gJJVIdhdxgFifC6J/PjZD6OLUS59dV06QrnPXka+hprUzODqT+TRlU
+NjaOecoUVdoDWGUX4+jBO6Q/0eO0JWZaMkwer6zANjq+wL1FOcNLYmd2JR/1vM7
5KTX6x1KsE0sOqokImwwb4JCDCQ9Dcv1x+80MUlpJ90wQkVm6w4qC9w3t9W6glbW
bLc1adDC4J6U1UJ6dxYwM7lxWjzE3XzLpkfUpl5cDnhyj5Hkj/THga4YO8YjbkmS
+7CHWeIfK5wxvwBUf+YywBIik3JC9agfNl+tTA1g/b3RBOp2pX28XnMsCzRshlIK
STVrUtuHR8KUneqWBBoNpRQWTKI8CXG/8y2CThvWQ2GIVztslW8yGhC+9epHom6w
wq1ed2zcdrO6UOEUj2TCr3CfuEcR+uS/b4PdAqKEhxxrXLyNkk+6WSw9Z4xKfeDM
C3FF8z5jqbgn08Q/im6cCtjdBGMjOz8X/wUhqtkVGDUEVlHD89vd4BPYDOHbTm1w
uYW/tOXhhmMtDyqNXQ1O9jpQ60/ME8lN3Zm8RWV6LZSlelQoRxoPvhGBkDply+QO
EE3yTrQ5YhKWyRBY28PGGPd5/4O0RFyCyFT/fHYYfcVW4gOLtYouCBjEAiT/r+aP
O9g+VeDLF7mlru7Qtthl3utrtBfbQzUFaRGeP/vYj39EjHpt5UOf5K5s/ujpWa1v
Ang7T40QwqOeH2IsxFhbk6hF6v//rgVPWImZ9saqYYCtkO6menCfvDrHfVZSD8B+
5VD41yIJD0SYC3Ra/4KlnsUtc6eUYeyGI7APCnUYjvAXLI7h/RFByjZPT6QfuKpR
lMEp8H3U1GYLIPIAIRrdqba5QEQQJ/mIippxTYDpJ9LQ9a6nXHDDge0cvsBUvz26
73ia14jfKPigNSu1FzKyd+ZEyKp4JDV9Wq8UJfrzZideyeOtX+FhzMo3pdyfYb6J
RegWPLDewW+LODiDf55dXFY2Kn3zl3yCoAfEO3xOoke8q4BgJ901B3hZLznk1Ftg
1k8ehBJqVyyYxnVQk4hAdI6KHjccmjUmozGemvvEotsCjrXL1TJEihwdIrrm8gbf
cpy8LW7OR+E+ssf/f4s9pQGdaqgmxaHQt9AEPUefoaTf2AxNR16oxdkbuD8CsA/Z
S+1t9yvCLgVdUaGz1n+JwTie+Y0uE/qCJpUtCBDIhm9peGlGuF9LE5fvJS8FB44r
rZhxuYq7qtd6s0SQLcvw2+HnTvZRrTorwvEVF7/tVbAW5XJv+IQmbA7eTDN9+AqW
8jXVOrqk18P/KiizXaepJZIPSIwaPIRVRH6fYTNJ/So5G+9YRuCRJStDjf/AYOT9
i0rd8yftD004qen8uNLNmPSXimc3lRNzjzU5tFMoAoQX9qQ+XQUPgmF1Bw64xiUS
uWeVAkI3n3ra2oKGLQGThIUZ1ERtOEpP73e8o/7CXkuVCDyEzxwTrjlMKAkc0tAJ
79WT33FcgWuG/p1kZN8ygSKxJ8MurtAvuBQ8sug9EHiJBLAG6SKbmuXpVAn20qEy
QeUKTcz1w4QCjUtk6Ok47roo3f4veI0C22xb0lzzr1Ot/pPR1Kf5ry62ZYSESC4A
BAzLuClVGQu9024+W123Q4dFoiALpuEHl6+4ohWmjaEfZ10olRVC3VYjjmRn+j1t
qt1VwJAscQLjQqO+gp4ZR8tf1JQLCA5BU78pZPqXRAxxZnt4f1LUAhxnQxOCz+tQ
Tw+NAGpSeiVLhRWZ75RV0jOnOb5lDgy9eMjQJOHS1BYAeZpQ0jagdhb0dn4zChfS
/C1maXxXzDq8bIYRYAhQVWaoRFG8A8oHzCqM9VYP94f+6r417a9PNRLY3jc5p4K8
AFbmprCpn8+W35Rs01nzkKdb7CUoxjyL67P+eDUVt0OvN7XCAB7WqRkY04nvO1xi
JLnwrBLVyyJcsI2RrPsaCIT5hjKXgHx2BkHG8vYPx/+F0bxn5GD16dgcBkvNK1FH
S7KHW6q+TS7jw5Fiy7GLUZbP0pCo1tzVyHYkmkmfA3dzIWpowsR/fKBooOY3ZLvO
6vLCg5NKRk2DthRAWSr4L1Gij2Cd9fFcaKtz3bFv1gsK/rgIgK8nSOOF5xDbYg46
llbavTwQLczmnr3AQ4mY4GfJUwKPk7GIPEUYu5D2tgHUfSHWUShbmflSbD93qs/N
taJais8azEb0lagxLoTy0Dz66xb+AbU/paofxDwqTRZm65DvbJUfXaTiW6mLR9si
uVl9bUyaAIpSoxM2e7i5fG3kCUwcz3oYgqfR+mSz4xODMShCSz4neutYK1PAgJ2s
nSkMFLuIeA+2wKJo18gZke9vd2E4UK9L1+5MMPDM4TGNT+hGKNgYyl+4HEx8jFCr
fPNgZLnPLJItG2M7SBnlai1na//KZp0xBd0giVHckE5enRhK4jr3Du/EMvoVOHB0
23KX0vyoBwtAlqQKaEwWTvbx4l/pnHjITQrENv8NV2K5wOF+1re+1O7tGMylk1CG
dEEL4CC3pGLUZGk5DDFTGofElHLhJnxoB0EtwjN2SKfDN9jNLYGac9UiUPTicAN7
IZr4vXwoNdeh08C6V6aK0CRl5Bx4p26HoUDuW7kHDkJXCp2T0eIDeHOLHvKVNLHk
wGUS+sSEujgkt/aYqfI89oDkbDLBf4Wzi/DS30YLs88wn8bUYPvw/dlnTH1AW5Y5
QkRYxF7xu8EdpvhdDH6auaLd8w0K1qmckB62N34qalejjifMkz6U+3olUguo0MZI
h1m1pQ2BZnn4tjPJmSTgwxcB6aHr21OB4gXQJLFxh1xPwhMSNHlvP2Frl2tDHQKl
0qQI1yF78UyP4dYUyHYGr/kp919PpBN43r3ORFLytag5zrQNs7LPuP6agYhIK3xD
pDhXHqM8P15Np2Si49iTMizv9a62yB2yG7QDdFmdQWm6YeDaUKXoa7DwMHwZXbFx
GhJZOLKp0w3NbL9Xm0RxJIzHcNkUAecs6vAHOS3/zPTfxRggNSfslDq9I+S0IpBb
EOU6RjSIUThnlPG++thLMVyjSDrVm8UTg1vzkBD2thU9rzLy6eLioRpdkl2J2Fki
RT7tC7IeAQEsoFmyNuhWbC5LRgqKnxHrsf/0kH4Sw2P+2dxXbB9qXqmi9fiBwVLN
juftglGtytUQ2l1O5RQYiW0bjtj0OAchbTDO14MrKIJI2StfWKJOyh0yVZ8+RkPO
ZdNEVYgTp5QBIVUGWTQXRKA3aXQftm9mBM5i8O5y+mAHPGex1BQ5Kw+ZlU8618JH
KbHCSfB9wJdsniipiLeCrQRK4jnMGKg/EAbXSjKmgZVjQ8VJJ44mpNMRLhKBD692
dvVr15ZaNALavvqL8ytduRQM7+Xojk2ymqcvKA3a4CRifbDVJhX+fxKMyHYGONmE
X9td45u3tb7ZFyzxQt+Q8CuvRlh5Gsbm/T7ME4lFfh2ZxORFpXBZSicBTyyzs6kX
lEuD2VE9T4frfZWabA5BWTamLNs/TEUtPnPyE9gM5sVdyWPlDsSieCf5jXGL9fk2
UYqKXueE3bpa8k6uVsUTpxi6he6M0svnzfDGM3lvW16kc8ls6sLgLoGy05UFlxLd
m1dd3S3QGGoE+j9tptwhfD1YSooDLQNOGr6LAv/vuCaAM3BLw6b0VbTMswXEzOOD
vyrYPpaZz2AqZzJbYjFSsak1Dj/qtYDsl7dsLaQzUji0HNMx/2Wc6F2UcH9CcBQJ
JhwDdfWXNYtaoJ/1+mbpwmc9TSiEsKwQweNWH7QfpbIwRmcLxLvQHC8UMD3c/OAc
nEtjO9rc9vNEUGNjHJ9sEanqNA9fx1CT0+BMyVcxQSuqCOKEZcifCzP0+qdG71Oi
fYB39CCrIKj67CeT7RvQz10WORNETfy2ZpYcWARsixwSaNEI/QVQmwendMtwbiCO
9HNqVKQgnsP51VlXpeOQTqIqnMEGpowhM+rpR8ilA9ydRuO+lZiUaVb8EKiCqKzR
7VbnUgOfc/iewPZcWQhCsdf/XMne3W18XnR5s8cIU0jQQ82UObI/zZuGN2P2Ve4l
tucSTiMjJA60TJiN+8xgkV9bYPxqJ8ivYw2ifth/kDuvhBpXGEXwLLvX/ag1jO5r
IbRQn9+TKSTZVgdSd1jcmxDzr6yHAx88cYkc7NkaFVsCKihzXr88EGMsW6Zsu9+K
Uszr8h/c47ddIn6ypGnhDlyqvA63K7aC4QPpc+OWBECPvcOYkHrVSGUYvH2aahat
KncuIcFiKijnPyOzJ12MLkbzip1pN9RQ/BQbiRmj5Uhgegp1gaN5aA92afCwvA4h
014IQmxd9TbPiApflm7sZnphL0s6Osx7MaoYVMXObBdZkT1yRzL9q4NujcGjamLG
lGmLfITNFHfAmW9aawaQGDAqeb96tjHcNoH4tE0TIV44JMBktZOqaQ1kc1omM1Kd
XwEV/Y2/4MZ5/uAryPi/xkME3pFMgyJdw1sbMkgCDZdsKfE4a/nOu9kcjGPrBCfN
o83qRi/XGzM0WcTaErZybQi2w25iLSyBOYyWwjFe9GwHkS9e8LP5z7ytNXZoZxXa
XwdzcpnHeTYmdhZLDeDgj0rrRaVTbytbkSfOVs3psCRH+HIeFtRKvpGgPW+uYxlc
S34aZ5/DcHgAIkF8/0+VK9Y0WJ67l/0YJlJWxeecB/p5up0tzkXKj5cwTXdkDXuy
URRtxpZC85xxd6EHmOhPEg8Cts4acGULhsqQJCFlFRsNAjs6iDIjR3o8VW+bEAYa
pidlvc6YsRPVRUx7yJIAQ6eyMzT/cmuG7DJS9hzk0aFbYL+YwELHRmCiNG79OWDs
mfYMIv5dt5k2HVtJ925c52KHBcoFaQU5BoT4nr/V/7TuixSr5ZL0Wr2+qrfmySSH
bqM0qyGWOSEWb67NUxqIq/2f9LNM/7anrLQDMDeU1rpQUSCHGTBmQrWg/QVUPnrt
ac6Vsw53542v1YE/5SLfOuz80cPpAPR3KOsao6qTZ8RPDRDfmwT4LV+o8kbyurcI
vxnANCQfXbCZuwf3iJTJpNxbvZ9jWrO63z6h0P5r9UlDBNIWdKznWSy5H5qNR8vs
MH/gwTIYQv3f6cu4qUzmL2awO3iN9ZpYgo4tpUh2VC2giUiOWSla92LOCnFlIsA/
S8DG5ObGuGe3vMJTk6/vJKMOZ+nwIWSk4S7dcNqGd6zXd+uhmfawZDm7FhECCa3j
k7a82B9UBq5jgwpBeWtoukvYBUfiCymC+5nyEqjRU70ZB0o7fadeS+oN2ubZwuR7
3QMDlHehWSfFiuWY+hU7VmMb6pJcwc8FFuUpxLawAZAS1Fm8OMyxWG30SriUZC5W
VarGHnZuBfkvWrJnIDqftKivIKrKs8kSH3+BL/3C/JSmQ+nDC5j9XAVjOhmcshyw
gZ7FGq4JOk1oloqv8knKrDohe7J3f9yzOSW30vl75OvFs3UPQ4u5y0fkEHvqmyQm
DVgjbJ8B1heIlmij9gyH/mLRwQJOO/NiDj8fTSoRdNaE6QExd85SDyvHG2W1kex6
h+yoJGYl3KVRhTwf+MHt1fHvOzTZ3ViyDxoQURhv1z778Ha3zZAE50EvytJz62RE
2s4Agw+7LX3TXhIAHGcQkxsjBBU7GfBDwoJ0LN8V5qIgs788W5pLdTGeUmXMogE+
oO2oityodz4R8Z4npSpJrQZdxrFQZrDCPRipHQDNny/+OhBRCVgoqkKVm4zLlQ+e
wzS7p3bZKCEHo6sNY+Es3uzUDan7s7q8ooEXmHJZRMcYIsHdoWKiJKP+3OWlnWjq
ajgtwxzuyraeKyC9E7tMyuKMQ7KABub7qQnbZDDlSdFoWjD8s2Y/lPAX4nS8B0Ad
Bna4XRwpH3yEwAkCoU7N2RwtEo+ITFKfDR8OLel1mR2LTX8A2jDPG7KBONuJgZKi
xX/kI9Z+6psSbOPNZTt/FRTAlbRjtD6jSey2n3eCQn9SmC8g4vIqMKJzHNj2j/C2
bvF+2oJiYo2CsUKdjTaAmqC4/cIqFL4+iPfcG6MHfAQkTOctuszgreKkbJIVKifv
shBaR9PoBJKv0iY++wet9uGbT3Rl5F+VwfbEiuAZzIFGRIy6r+IyKwaux/515dpA
V2OQMOdDNWmy+1JHvIHKJUAQmeWZrkXd37ZebgeBjBYd69IilE4RGViwZG+XGHSb
vKkonjoPZiOP5yeP2FqODSVsoThBmb1CbuzTTYTbTHrYg9NCk+MZA7EYTMUXwLnn
NS6Ep1XKVhdxf91jkxyzoMtewvFciC78INMAUDL3S3xgotuBiIIuBv9XvQ+tPguE
ShgbtZnQwyUhuz1kF4R0vmwtnFHKiiKtfDsPVQmHXByYSgD9rnqT0qDQoY1xVwoM
fC77PPCKKD1+W8z/WzUemytWZW7WLUwQPwECGUPF5OD7LQvSM+ME3vxwh70MJovb
XyBe4l08sDiJMTZMsMKS0zW73L1lxFLEzRnlfrR7saWRGvgbBuRUzKB9I1iidn4s
QIZIUZYk+JgLzXcmThr8x4Aaswsz5XqC9GeXS/BUxKeyBOyHc7LItl5v0Yr+DgWn
KhIxteIWw+gCZ4D9aPvetusS0eUiK3Yn2ZVyZTev6uxTd4yMfUtm0PwDquQNZhd4
hwZ30X/TtIOhygqXYyFOg/qkh1Tq6VXVZMiLOcQxvNzgmn2gg+16qUYS8D/aBESX
vmTIKdRROcLEtQD9LCxAdQyI4uBTlMPHKewnOUeewn0lLd5Omz7BLWPlFKqXL+jb
Eu5Wqt5YemR7Y/282JC5ORCOTrVMqT5yiuJ6BsZKJOYDfTHhd9lHGm4gBsVaCN18
8bH8beMF3hVKMAg09571i2BKKO+eM0iGjScsWRELhcDqqtopD9Ot16XC6dyrJaAJ
gxZLLyg9DcNVzerak4p4ciaeuomZVtNk8wS/gQqqaHmCAOFFKtBz8ijT4cGw6B3E
wWzrpVXsCwJ9outEE3SKy4PZjia/K4B5duJI5c7gqvK6knY72CK69umx2B4RbQvV
QShnXBroLHhizgm1Ah08Sz4qsWaLUeq32dkIBQkB5718HFJVt+hsRVySQFTV36DR
wivkBkndK1uf7M2PPGnb+JKvOatRxB2CIWCsHY+H4jN+kjqcRS0k58RiMUzXtfQ0
maJF1YXAWQIaQQeOJdR26zPd9d/OHAYOeLCCrM3fz4w7ATz7CdpEP4Ag9oZ+jdeH
Ai1Zl/ARPjt6S600qTNTZRAkLHhm0Ov3qa6oJSRyo6O9il+30mmDvJYT/KxuCPnD
AXAMMfAoayxa4B7QBDMoqWWgkMT62qA+85lBBb1uGO078uVwt0Sk6LtdDaIAryUP
xmd8AsUTtCie0daoIV9MsTE0Po6UR0feeWzeU3Mfv9ay9Uh9ExVGyV5Kz6ufVMHw
gmAJV3ASIyIs4g524LlAi2X6yYtLK3isjy2oQKK+U4HItji5Q9SX1CSDQHkBKdfz
jY4UO9VEpYEDlFsET1MLOrJVj/6pfCJpyAhkZx5FwZNa1kNnFVjoCX+Mt5csWKvw
nsx16tRVByKMNVgziMN2hvQ1YBk+4m7fXmi/j5MfZab2HY86uwrJzSd1oW3JdnPO
v9095/KM9BgFma+xUCLQl/N4Z1Npm+NsWZMHIqri2p2NalXLm9IpsgM2J3Zn95T6
MXHNPzz6Qo+Qyfr+Kal8KvVQF/Tpxlu2V7+vPI+QdV6ffw8tg/BakZySUxI0TL3/
XJ/NcGLGMxGTUIOa9oYAOeri3bkCGLpKEZ7BpDd5aipe/JExzdAqbYMsI0gtyoAP
5DahdHF55H6qXxlZVODix5f6xrAB0c5plh2AX0Xn1AGazybtFtPtjneqYjUnxzNZ
2chcg4KZfQp9x0zOEO4Rhqzvh7CCNZUiPi/fJ8BH6ggjpH7R6oP0YTxCKBOxpicM
eGagaCqrlPyeCQId4927AtV9h+WLykSkNR5cD5jUV3MA567mCP/5aO/lLgFYcSXz
uDK+6rCoBiDY46uyXb5eyqmZEv5KD3gVxdjCXlgaOE3XydhcMl6Q7ZsM3aCDcSFo
YNlC6YdvwAZY7VxRQYlbO9fGBjg3zfplp9gSO/w13E8mSZdHYW6d9b9V9z8H/K8D
uE7oiU5fCbJFk5HJO3zzgGVamKQb23dofUK70+U/GJjqFWDpEq9L6+2LNWJAS6vu
ZXx4ELq2708XS4UBOfccXrjKShAM3cW6fy1/+lAP6xQGIRm8aG7B/0P8986jNvMQ
44wThvLYNfuCPMjh58apBXQCjsMDUJbqVQAJUyxYraKe6gGBuYjHyOUGW5LTf2d9
fA8NAz9cNHY3Ls+Jga+r52ZMcjDVahOlJVsDKJtnBuDTAlU+jh47zRV2cZoy03+6
y+OgsmTVe+Cm7JndMAwxr2O7vZPnH0kxM1J4x5FJGmznZdnIWuLyQHyUjw+sm7KR
AhzuVyr6ttE3xF4pp0bNH2Onaf5i7W/qi1yILjGzspiV4yiFhpImLMSavtDyiFZB
Hms9CwfFIgTDlogp0aVLYPsfUWp328tIzzBhLoYldZzY1LGEL1GyMkrHTMywC5L1
dEPqRXjUk7hZRP+ielHIF1olyBaDb07z8Uk42QUvO4zX9qjogIomY724Mk8VwmwH
mYVUEybd9uTGZzI5Wz0Q5GRQnHMa2FAEyNfHAeEi0mJ1JL8m3mVFT46h2qKCmgD+
HrqixUjChcyXjhW5ISxi5dmZZ/8zY/dp4OoTvYgQqjzCiWbjaoL/x4UvndignmNM
Nj1cJ0/eNOiUnEhqQGdHLjLTKULIKL7yMxXtvjVFcOthrcW4TBg1rgRGIisOxAr9
WTq2blrzm3bLn2pj02yK5FjZEeQ3iQ8mWr2XDi1S7y01fBLbBC+pKOmmIMnd/GBc
vZWB7jDTFIdTpNTDSeijiT+p9ihg6rXhxqLRbIKKHC6nVtrIamxDBKH1ckj9cDQG
9XWNWPUsiTM1dZ6FK4T2wwjMwdk8xT8lIbHCDneor55TbJzBrNAdD50z6KZDG8CX
yNwE17P8Atm0SAHl+uqhcDFnYfNlQ3MLp47e0i/I6BxvhlCYvmE04QemmFGdHvBg
QbHlNislErUJYp8lm72Q521jTgUtcVN9PEl6fzDX9/jfQlkxiP28LaSVQjN8G5fB
MskuC7SbycjQMpWVf9elTyTnvKXEkDnj8+1sgL98BFIY8d/9vCLG/XFvHR0580S6
jtDzOChCmgmedoLKknqezE1h+OVs4y4KGjTUo80w7cQ5qbR+6pzYBnMFH4epS+JT
w3wSTQOrFlk38raV1GPrIgcIp+j4s8FSjqKNuqBJDnIy+Nb9rW0L6UgznXFS95RS
jn/Hc7bb6TXRxXKgndzMbVrLbHhS8Iok2/GfQ5OQIRwSUjIOQRTPkXoHqAYBb0BQ
cIY0pnOSEb5mUAmSjForxjx2YxVqBgOwx0N4VFwcoWTKnQzphflMTJCsNZf2Fk1y
tkpEFBOst/4M+viowXSBGVc1kQDZbmN4Rf7zYb1omoFSmwxJo66bOB/AT8tTHXqx
tkPPWqJNJzEhU0ex2Inu8vHIgNPR+hgorPIy4FyVkxSBDIqPWexYClM/VOvCRrGI
84sLNJMkSHDv51p7TRKFk571wo03LWdezGIMqaHZUM8HALqehflMolsWFN2/dcjr
qkp2cx2eXP53QtNiGnTWcmv4vod1Jfr8Xm7dCjMnp6+9oC6bIiLJM+MIrmtA52HJ
U9KOiJ3jB8UQYeljEb+RBJiAc/EKwlsRCeYBCOFAdUuh5FLPM2Mr7CEQ5JTH6rm3
tQH6Sc4UOyg1ntlpmo8StpkWJqb7/aLmHY8W21Tmj6VcSaEVMkUHp4xWz5kzVDi0
CpQ6dJTZPg6j/pTH5wJENpyzAsovh8sidR5fAdg+AAS3v/oaUKnuqsyKKSsGHzuT
Bm733KjrFoT8IqJRGNVHNY81khtiOihroz60ELVU53iQMI7c65UbrzwKBnSqWw92
8vZdcYR2lr6R4LFGCNG2jv7kkszoVd6NFOVIQAXJJjDBJ+lPeX8YLRS8a+cSVmGp
06vdAa0YVza7M/f6PhIPXkTZhRMhuWA5wwh+26TfLjGGWISI5OuZjWYot0xsLMCi
0wB0H7ZJk4KxUhoQ0UH+8dkQQZMA0h7GjrOUsT3qCczAIcPLAKLzDf1ieXxoH9n5
/VwfSXgzRAx9x3b0I4cYz/KZCtmHXyDy7KlAD9cMOBtoz66ffA3uvjgpSiJtsGhc
R3+UHvd37qM/PtHyHlzkwhdGT6n3SwCtnPKK6Sh6BQDWqgxaL4JFgtJGjFMTa967
WvuxWsGmDpr1ZwSngHMIWCv/TYWPl3Qs0nu9eY5/xc+7M3GYs1Pt4ApZTzONYvoN
/6S70kI8PYsYTUYUBP0X8025KeNFa0HARFR5RZocbUiIWnHAJhImTb++A26C0pa+
9b5kIXiXJJi/qckpOUGnvzA42kyG6We7wSvp6+e+Ij+UKNkMJCv0WZLn2HpX05gT
NBuFuPLgfo9Wungcg323HHI5oT7TztIdMMqJxXY7g5xH62YSKkDMvv4EbBFLojwY
eCdLYxtNL8yilMBYPjBi9paOm0dsyeKfi66nesYMvIk1e4HgCZM4LdUzVd/sFHBk
xIT5axAhVBa9nnKjqmlJ613anfj6NvPreHDcAnrqv2Lg9MskcWbV39viBWwY0cLz
BIQdpfXmegyN8WhcjLlFBwJgj+68go0szwoC2VvhzFqkTC6yIgLYXncB7FPMfQss
AQKKYcgkzymJAx6XCokvSwvsjd2SEmrI2fPb/qSwFZjf37aXTtjuTwRwdXdZSral
eKh1CTfsZhthk/+ggjGh5ynoOnSPt+/bkJkU9rsefzDIUqxoaGnSXtrnE19yjTQL
mYsPMsIet3JtEVRGeNXkp22JvAoGGHcCIBF+Y9T1XithkC1bLCtTZszrAwm+CsYq
7mtNXVbJqVIjb0Lx80FxwCiQTWOmzW8yxlm39z3RPzOjQJ+cXZZMQXueQT7cqv6m
a7SMg3fKXy7wrUDU3369IR5CZ1s2i6Xpm/2UkokG/b2QfPK+T2uPTN18/6R7YxOO
jQepV6KaVcON8eI+84LyahXczFD/0oJgqp8GUl6nKUozXGBL4d8y87WEDUaxr9km
kyEbX6Qu2B5Vc8XSZ4A8/nRtBZxR8fAhUE1X3Bs7a1Gf8DLCarEWr6Ar+UhmCWik
sbUgr/3bMlTMj2x4DEZeqN+sUWTt5xyLgH0+Ppz6XugLMDlc+5CvsyLA4NZZb4aU
8fvoU0Z/uwA9QTaD9o/EaFvkqQJx+ey/FzDb5BpPOaQHhWgY0zqBB1h/1oHva0z3
w/VUPjPx+6DVVg02yAop9z6m62CxGexVyvRi9c19M3fmgAdV818dfVnITCjC7Lig
LEAjBwEAifYVU3yZ3b/t8X/TraxXI/eOTUcWrljn8shXIhwvzwHxpHyA+rnCEuVq
Y0IoJHhCmnT0onI2DTw+UG6I7czg+YXmLWPG92/tJdmRHWxN60Ysla0XANcqem/R
k5oErUWZ5ASQkhGhtS+iCv71Rn+XgpzqszLMQps6iL/yPRqrZ6ZplOUB4t6qxSS6
3QnpwYobWbuLrR2MrZLXC9PKzaAbCDZCBpRtkpFtVxBNMZHVZ/vwu+9iqNeEWbJ9
Anur7G814YmzWMjwTmrVstUJ71tFb3yDbZhZxY7cy65SR4fzVIqcEBi0RCfjF0ZD
l+NGZXfDvkRZSv2lnpg3+BB3h5kwpg2lOgjXe6usV43ksPYXP8Sc8jgp1772O9bL
/Czw7GboKh+wtDP1COjt+tQZp0ZAsTkeerYaRz/r3mPQqrOot4YSx2m3VvtJcNTj
w5PdlUEndfjTA/ArMAmNCDPHGv24mzm4ZGcWRVsrTYJ9IrNr7gMiUQNOps1g7sKV
/2VqWzeZcstq/CNRe1mooA7HcTxuKJwDypEdF9b7mojpJEaKLHibo5xCyb5VSXPL
B8LtOWC75k6qO8fcy34w/ImaPg/kaPoodnmzbeD1EBDKdAgRAeftYn5T5/XJEBY8
Hfj5bnPPEcIGkvY38js1A3nzHr6yZqkf5VrYWUjGixfpS+yMbdxA4yWJdxHsYAAt
iaw0IQiGtHZF9hv5WfusJkEv2hD3kkmmZFO78N0S9I3UngHarnBvGaIPWfJaFZqA
ZMkFf4QJgOUYDp/Y/I2+aJRiMWRogwWLjlUxeol0iqlYzoeaEdbPiN2cOFyYnjKz
Ltqpt3ciVhGZ3x8tYTeZYN97224PlGXQ8SoYWOFnriOEkpjz2QQNIsizAhd9z91o
iGgMRsk74xhJp768N5mpTxkeddC6MKwcHJrxmpKlqU57oghRV9+b36cWShUCRdWQ
3ANutQavzFoHbybrrekIyEggf0FW5FQQENul+4aI13TUKHb+k0S69gnLJFOBnEoA
ZCKlw3qO7HSsSNeL/knYE1QMxouNiiGyw/CjBSdD4T6fKY+65QJxgprWpx2xEm5K
IahgTADoL1aM2qFnh6Dfc4Dt1Ic5pMA2EBN3az99B5+MSUcgnD/bhM86Emvch8ID
C5XI+OsPI9CvL8qyt6BwjZeDC/FqdL/3nh14WrFnkzHwSDED4ONEP8CxKFfno8OY
r5a1PW5q9eZOpxDWY78Hjd1h6kKD1/8gpte8k6kaBhbad4NZ+9QZZcJimJRKJMaA
5HyrGLjeJCSlrZt7TDUMQyZd04RnBFgUFEFAhWy/gTRpXbqj5o4Ybfgz/5qVzIb7
bm/Fnouzd9O7xEEVe5ccCBPgig7sdObxEdgbyQDlFZBcVhCE8294mBwvNNNTVNe1
gPDcgbnnM4AKm+PwkfpOyReR4o8ktxJuWwVaJ0mwIQUHAKJQrXmVmJbWreJL5uQe
CUXLdbh2mGQAtBlX5PNLz1QRxCfcgGbCYH2iT1F8hymo5L/AfYEFKz3Bk9V5OKxh
532505/pQPCHgjmsc3NiqLrgI6+BXo7HeH9EFYt1G0W291lwOu7Pmczzp0VJRVdb
cQZt+KvWmzF/FVJ9Nhf+8264F+g4VAKU4cs3WuepDVoGsJZyYnnuTeilRZGNTcq8
9n5xxyk9m8gtDXxxC5aoScrL5VHCkC2ITlAOyWQctSWNtSQjw5dyB4fRMDZ5lUEo
+bos/OuVNOv+xrMCFCT7kbSzrN9hu/dksixqsS67zxxWdpAeigGNBA783j+AK3FA
fMb1zXWVg6WSHR54OKfe5JZ+jxRO/zfjJkU8sVp0jHFuWD1BiMG7KfG2cTYtxdOi
E4go5S3kgpootKTz/sDjIyyO2Xsno0HqEQmULlc7p+y0Y2gXTD+hnKCoFlxHE+HJ
yF/tm2xUoXIejOJqUgkjHkDyYgW2U9q1hY1EjyW1i1BgDtEQpIylTTrxqiE8ELp+
DH9NOQeUjHWkWFOAOYqhBsA6Yw+hAuJAaawGQ1DPxonmRah7iGHA7SJyKtZx/tqf
4nNh7Xd1BwmrKFZ8f2thPNW3lGHU0Dlo8/MCx/xnk0+63mNLUxtwLMKoGyrwYLRz
Fm/LQPsy0H/J8UZj9d1PpmBQ2UeKRFiJhBFfUDK955SJfgGVO8aok0/3WlfwXFr5
Q/ACq3M+tcp84TtbD6g7XQQN1iFS9bAeIdzDeOrl7XS7Q8gCA2WzlovH7XPVCxGm
acavJ9GbIUoga6vhRcAOZ+iPF9Go9ZHB8T8qr/gcfYHlw6MaEiO6Re4AF47w3rXB
vWvgunD5SjvNAWZWQWq0dgKjzAh+hsjF4PaWKktUtDlLFCqpWr+R9PjR4+UvKFvP
xVN1I6rBOS+v3o+n57Q8GKzc+mHYlZwto7sJZ5MbgKSzxwKvaw+iAkaGhMv1lJYc
LBE9HZCXCKQfABBYNiBPHjhyTan4/s1ZKvncwtdVtXbC7ToHc03ZzkZAWc6b4RXz
fBu4f39pHCDjvHlU1daHO0NWBKzYZRtIKgKlqOfd1X0857/g8/e10iV10kKRMW6Z
qRcq8iW2BUKWlw+7XpFSTwvbCY0fKyME/tqtKFFsv/574qYxWf3jpzbaJiyDoMvW
qsICQ52E44MQ/B5ZMUB9YbHZpEwEUlOGXfZHYuiLjMXkskIOSDMQvl+7wMJYOQsQ
+6SBlFiKo08PUHzvGO13eFEDBWZxW8eT//qM19DJY254ARId+yWiPL7/Imopc9ZG
uDY02YfV2MSyYKA1iBd7dS0TddJRpSy73OUMQRdMgAiZMULhBVRS/z75EjX/BTO0
76is9rOvPsvWIIe5newHqBhNK8c5OSuq3c3UzhUpEFMrvgDFMtCxiEPHYHqikAHg
+SwR/FS581nbqgbnX84JABd1nAH5q6LkmGa6PZhGGKTxG6+xzA65mjvnElbjs8OT
mw+TM1XAoaPKWWMQ1+bzCWQqSqHYIb46PLkDBPhzJqBuBMEiE1aEO6lU9oet14SB
iN1CJTzXRBeUplJU3kGrk4bgwNjAa2AKqRulDHmLwh3FiFgh/nE6Vz/3T0ViCc/1
sYSLRUTGv72fdq9TZq8hHhirIowHx0CdZ4a2rP1zm25kB1u9tGOAX6EQex9axU5q
q2XPUoAAh5DZOWl0QC/hgmV5RBMwmqFnyHgubRSITMUMXIpc4hg0UqQuQ5oW20Rw
QaE/cVUcAaMpu/B0egpyd0VGpUGcLHM3tZIy4HrIlttGMocAAqw+uHBzykgStMn5
Prgjh0gE+/sJoI7+XHsppULUEm9TkJMMkm8uhppR6aPt69stZQ5ICbEflo9suRVm
+Q998yXcyNJXdNCGcVXvQDPN/vsIGaiTK2xYdbxWMPr1qxe6n2t+mjQX84sDAIII
mcXIn9sTCgDPIwE/Lsv6PJQdhAQ/B+RnzwovBgT0F9hixOaPhQWUkiT26jXG9qBu
rjGGufa3VIJISJHMjlqzx4eFmI4mIjfiuzzGztVExAxjQYBlYbaFvExR6jgs/E5q
/J3VDOM1A61b5/zuzw9kKxdScVtRYUlcdedNsAK9BV1YNyWmNlw4+aVlda/2P2fY
CCN145DE6mFVUGo7cl5qnSW+fCGtrMhko670F4G8h+Aci8kZC2rrXwny3Eo0r7hI
C77QGNWePV5q3a2FC6e0x0PZK0vfztDLiuLxzW5h56GBaWKGoieWLHz1JqN8DfEy
zD8N791aZaZz3mzruSj+hqDTO24It3KxvdeaGgWC2+4+zsNbJHDdocxX+0qDO3Bo
kBnT/uOmck1McxcJoY7CUDJQyzVoCBS/Swly3pN0/eRFJOLZpAzkLXN7ohWCdZ5n
dbLsJuSHRsi/Px5yY77379GwVz9cbJzCTX+aCDVBncnwx2Abfthggx4mzgeJPiUg
Y+iv8JuDMYjaKF3VZBHGeXvWCVE35OHsJTcgspDPVxW52rUgK8hvfSRQAxpZ9SFd
vwgVhcWie9NGk/hVJOjf5knnrpRP1p7boPKMUx9zxPaBRnsj3djEcNVtw2Z+O+Vr
gME6/1ixMPjCv+utD+Vgccgyfw22AEX3+ofQdRlTDEPSxs5tPAYByHFBpoYAkitb
1g4iBh+xWJH5kDZP0/fEepl/rm1SHTw2EmhYK9MzrjLx11N53oMDmorO4c4Oyd8Y
w7bZOsVmXmi9xzPI0Sl7dKD6MjhRUzjKKclouq6sqfERjtOhD1o5147EyRZic8Rs
uDOnSV/SnGOi0WVKQN/RCrXoWfkdVKn20NUaBqdhViA9E6YUkidjO1AsyrymrsSV
tZPSG2IiP/aXSPmkkp3Be2C6qrJxbTfG66yV8SWGBCOTpStfUNFRlQnh/E7T0R2Z
fcGizICo12D3vMrUTGBaLOff3b73gMloFxuqIz/56+rwIfVUdOFDDe144ip7oic9
poFxA3GGgGHxFo+lkrkqRAMFanSt/vXAOGWkWr5wHgnDA9OaFlKSBNMlzmnZm9P0
oB5foVhCWJubkhZ/To9SPht4MDx0vHW8tuHYyja12EbZGWTO3z7ATbn9VFa9ClAO
5JGXgmyUrrb03O+LvII+21iHx+pfPHkMvWN/rtKBshNZIDUy+IDSgst9+Ck+593y
O9YABrDmJeID7DdFbo/sFzSEq4lO+eae5/yMptK+s+2SADnIE49PFRECGJVAFh8T
FVFrbHucH65RX7SVi0L1q8yF03i4PfkgkYjQ2M+2ZVgPq2Psr5P7GXNxmmAvtVhs
ok8Xwz5i7ZxwmmIFAMkj3ZUKdb1v0/01FM39MGzRzXDsCFor6hs54lQGYiIScVUU
FDPnRUZOwauZb1lvztRM10p7ikId3cLjrUTYOTKTgXFp/ewUfRWKqBRasTh8LCv5
EaQSYJX2jGH7jjowSK03nVEem3Umo+PreGezXAH0El8jmU2jxhAZUwRfeCc/0YXm
3jMB/JCjzhLdHsiL0CmutD/Cskh/cB3uMOIVj7RFgUVpMMakk00GHDD9W8iu5jSC
i0bSRAOHgleggUhenydU3wur259hAWm71p2pxqCa/Ghgnoz59Ya+GXIKQq6513tZ
1G9b+IZov5X/OkkUvn2k2f9PSs7AnzIxqAx91dlKncTx4BgWiSrTvWpn8HFbe+X3
gwQAzUYZZtlXIJI3uBRj3EsG4sZ9IQePPBtA2bMIuaf3M9u4ruKpMHWk6CjGwlvw
fTyKdqa1Pbqb0zC8sDKPIcKSMOzZoIr5QgwN941boxISzdQi0h97Xn+C3vTZA7Rd
+fVcRaZcuS9JMQ3TdrHYf2m6VO8VFJQezUMfYIig0/+uoxVWCI13nMiy/HjMEDC+
5YjWh0Kw7iNm9RkXlUwqBKHf94OUrkMwR+8cGZ3hQItKvLm0yqsQDLbO5mZi8oCo
qDiC+6wh+aBpqWptLvzgh3IgUJEIYGqRz4PiDFtGYH4osG8WH5AIolSbVTmE+nMk
Hj3AaGaPBCOCgB3UhozZq6Tmh2yQp4Ej9jzcnbAgg+nmoiHJXaPe1xr1PEXmDJRA
RtexN8F9N7hK3bEXahDusqItpNd0tBGP+qgwpX4TFwNSTN/1GHZzmWjGBsr1Ntm6
CFHBd4UyggytdHdRcPnXRiMwIKAvIsMMugTe2GikYMtONAHqj70vUPT3UND+qQAL
4clCgS85Lx1K/qEfBwkEzo7yac0Rpr4+8AKE3G9PVwFoFweT7JRKZeYlAjE0wG0h
Gtb0uqU0i2oppSrBP4lCz2OzwdboOLpF5Ggf/iRbGHHWT7mz8TsIQ9X4ZKm9x7xL
l9vaTwMaa6POK2+XQBngfzWMEEQ66eJIOF7EnpHa08TolPvR//UuXsJDMdBz37Pc
49LS+jbWIBxAir2Iv8wnMnYZFbYvC75UNi/eI3Ig8Y+I+o+rwezFeTU80jQ8COKP
Ksy3xJT3f53xvsh8qtTcpaFV7W5VrLk91yu39eJqlBeD4GZc+sB6kUTET3eFhfTV
xYeA4sdimlzlxuI++Byw94qnBnHOx/jJMLmRQ8VtJnYIrZrTmu5chiPMhIFxcVCr
POpZ+CVgw+pH06q/ATdKLji6Pzf2eaCnjlBOw2zoZOLx3Ql/Dnvoe5rTK3xShBHp
5eI/ks/TBac3XBnvu3zDv+RC9UpbGmblUbRzqyLKbxrKNsUBRfFlBf4P6TcUwz3m
57x+sO1/1L3/HcmvmG1pVuQBDnGgr/PcQegPvKhwELRUl2SnOtOihoyIgDFJi8Y/
j6d3aV4Z2ihmqTk4BBzlT7qK/VGd8BoOH5rwRc0U2/iqVWNlnxGZQhk/yYocQ1Fk
rct5S0swDBlSTVlNuEOOr3vAR8Qe0t7gQbUtZhVKkRzC+G3UnfVZxKoVoe8deU11
T8rJscotO0miZIqRYpRh761KzE9XGl8HhYoMysWUTRMjT0FxZjbJaLzK4gcGAh5z
BJxA1AldGHRyrdmfOjR//3wYnfJeoDTmNXaYL12eW/oZkE4qTM1XNmIE7G6HNlM8
jFKjtutU5txhfeIrpbDXPUN2o10qhOPwW+/VMUH6Y/cpG7Q3TP3DOmfm4H2XsxR2
sjXkYcPI5QZ67z/rsBJpAkaJOEgi7kZfJyxV/lhhRDL4KQCowky4TGqVpFUFjvpV
+SxJOaJnbOwSAwM1waMB+Lo7UcUblyBfhEnQ2owdAN+XgxMmwBMnIEeCo4QR56ye
jJG92FhA5fHGFXcJJed/qDxZbnN4ovRf2z+tXsWERnLqy6rUxnJ1wv1A1szQWL0w
0cJt/bI38GtD7u8dm00jdSRhl15kwOaU9RK1qxpyRChA9BY6kmp1qd5RaemOI7LS
kqCQc4oXGvofHOQZMUbBL0A6iZjQ7qrAt7pk/gd4fl1kClLIIwMHJqEMr4yBsJvE
6NaykXZYnRgQXOPy/Nj7KmO5fLkmB13roMFXcU/OMhSxKkWZd4GsWv/xRoV1+7Nc
kLE77ebl94f18sodiPvLFDtLLo5GcJxCnVsZnbWVgZ3Cx5FNL+55HM2k4UuhEIEM
D1qWF4USGOFUecb2PZZ4JF8J9v7cYwLFDIo3p9cTNV7+3wjTCQ5/R2nWpxCXqUD/
fhi9tD6m16dNX7I8dHaDP7hhG6NRoHE9VCqf+yeYxFknUCP18fMjwpJhmn3apoEj
YbG8VyqWk4IZoJ1D8CHbue3ktRsNuXAxWoDkKoYYjIwbKmzbn8gQdo/p21CUyCTy
LIWDqRnk3dhbeds/Jn6qgQUh1Rw5uea9XVbkuOw1LkdSyxiDU7cDu5CZO6rWML9S
BHnToew0drWcO8F6TozRfr4SqnW6tewf0IewSch9OdJTc6aG7mXwqIwxlE4jmr1O
2MqGH/RLaDBZ9oIdRnQcsIvrfgVGmFv4spgRpcxrLkkvaWSymRNMHxH7SixUKiR3
yJKjlKDpKqBgE0GBlrrjqeSt79cHAg142ThrirexSDCDdj7FjxBQLSi3008347qh
0gbftTo3A5tFG+OhRmrO7aE3bfot4eJeqYlzS8pp9bZ+shyqLz4+j78uxiQM9xGZ
kP54+uAVne3XwyAuA/0jMs8YnbZZdTsEi0Y0CDC0zxBuu8asaTf64+WijhL1Sy2O
BtmeougcSgxShMx+PqDEGubxZ7EOchboUpMtaQ1Sl4N89AzsEEAmb4REPen0CE+O
5pakTbTsQKEUzEMAhqX1oBgo6s+MrZRcNcQsdNmiOfPLKYyWlnKMwiU+6UAE6Stl
kBXwTiH6kenMOpKTML/ICW42iiuincPR2dSPE0k/l21yvoZb/0FB1cT0keolrQCD
Ru29fUEexosx7HEO8ynQt4J1P+DXp7A2xw/YztYpRWjpQ55MVf5iQEva5VmSpUI4
dqq4/z4C+AUXBm/9bxQE4JN8dnqhE8AXHgAlZtasSIRJ36k9cM8WuQWjFwHN5Fp0
8tD6Tnyhv/pHTLvrg4WrggRHKKsLasxI0u9KUuYqR8BOiFxuxTZt1yO4Mj7125bO
/vnd2bRte2fW8QBeoubqxquiOjdqkcpa5Oq9KJKYHWTF3hGFiQWHqPajCgWslkWy
UVfVpTsCRa7YmTwuAJTvqvebaXjRLc69qdTCipmWaSD1Kgc204J+6ovXMoKoa/sT
NyIFgEeqHeFJB3X5mjQilV0oGbVh8lTSLmmjQfwTDyDlf7N7pCQyufE+hOgufb6M
5TUK3Vg9i0e6tbn40ahyryuVcwF35L9aTiLUEhh3AotvqTWNfZFIjhZZBvglsL/9
J3kMJjOky+WLI7xrwh/SgXP/ddV9/QZX5pISYicw4ORwahbP+PX+O0wKoZafflwb
NUafiAVL1NdihF8HVQQjR1lp++NCAclJ5yjwLFO32R8tn+nmFIysS+uujSlsDNNo
E+sCcBV6zEt8iHtO8g3o6FAi/YBARFnkZ+64v0WbQvQfNEMIP28Xai89BLXc/7IV
bw5z1t4N0n71IxrEnjRC513RZF25Zy1pbOWPd9pHzBVcvA+ljG2oqKgPWHcrG/Z9
55xAsWSG5fwU9HB2VTcpd6V5kl0DbjuZMh53NnpZs1fu24Px1LHiJyCE40qD6SP/
jjJyeKtdaG2vAdORvvTD1jQUr2TOYAMyaaKb04ynuFqx6ON+y7tTATMAXL7/pTDY
2Hd+BVb292N6o6ryuMsW2QIREnF1SCPnXXDHLSkDmUvJuT8q+po4QvD8sUyBdbBW
tJgEdSHxqf14zHiok2u1jiizt6uiKqBjkZsBBNYF8qlIeNUvJ0M93j4usvudKCAc
EsRMQuds5ZKCW+PSWFdvNH0eo/O/KGBuUKmYtiDBRlCf9NvQA6dOD0sG7MZnZvdP
nnp6GyYKJvmSgiTbsKMl0RdLupfSIeT5EwNQffrm0pt9h0ZO/KV+NdCAF4AuNn30
LFNE7gPGV3pMtDwJG6B2viLlPQvSUrDgsLlaLwFGBUp14DYt2SSwUreYbkAfkyN4
E05QFexAUFsst1BKx8HMJv3dITBu5in4fDLyP5o+qvuCBktfHxqnyIgl6Y/NJ+a2
R36xk2Zoa6SYcrC531I5buouuOzfX8U35h0UxRAagMJji+qt8olBLwK5iVSoat4z
rP2hSgN/Byvw4JAaMMi43UCh3C8ogQuSxFHa9NM/eQUC0M65VWD9bR2yFfMOqeIt
c4HrRdmNcTX1pM5dEXgymeYvlMrOM19WayBsiC43eF2IDLZdiEaw4beeuwwSVQ90
o0kE4aZkS1ZwaT8WDr254np93qeGWDFJFsWMs/dXbP1l1dvgg6jmvqE6EuejSG0a
VOF494jMPIeUSGLUnn/M+z1ht9M5xrcdZrjrs+JeEUfafyGhN8pj4TbQsSiw14OK
bpprK59SKTVuCt6EDB08Cdv3O5ppTVamAloiEbV03PKO7ObTelJx8/dWDN2simEA
vkl8EPnOWY905QYeXCjeeF5/RtXtm3yDVizHwz7u/r+I2ynN4SCVFz4HAZERMtSy
QQ9e/iy7+gt3rT0CeHrJ609t+JztgwqrUGc9dPMPblefiy1tCculI6ZDiJutxGvf
CiELigeVDNwmqskgeTEv68qtWe3BdZCC4cAOxiK3NRsIPYcQIwEEbxeuadpetx/N
WCpXCvsAysBbxrnaE8GP4HLPww8FK0TYuJbIhF1DmCoeMgb86qEwGsxdbHlwgDgI
ERO1dhHIPTySCTEIIXFx0xafkrT54v3VHWXlRD8xO63DhJqB4EairQBHup2LxL7d
3TIcNslAg1o79r1N+0SADQDU0v5JgFSR6TZVAAdflv9B9TnCE+8RRSltjv+ElHH2
09YurNmLTSPW58F6sj8aTy4DPdg53jeLWJ4NnkElAvcaq6la19eFml8o2pT0v7Gf
ktimDwuJzybFqXsHa7T8JpQQ3JlLdTyck/ovQF5jncmabSU8fpYOc9wiRAZ5Igz4
NWj9z2U82ITo1jKI8lTIAW9aiYlu/UZdcMk2vwOTvbFsMi+5Iq4A5J2ek9ohbowE
ns6CU5h3BjXApvApLtrImXEbsti7Kj+dDRWAGNkxceWdeh7xqUinUBj+vQ5L3c58
tQY7MxOtlXHLnmPCaTHlMn+unzUwBqUhPkWyxmWFP/5Hzr6nk7Jod2bNAxVUU5mJ
TWcnmsd154RDRtpZA+LVqNdGp/tVFb57VX3BWmz+3LDDz9GYjgzdZT7eUaaIoOYf
foVuFvVAswpz5+H2VpzUBJWomRuxvAUgRvb6yvmtay3J/QqKiKF55G16GmSY7I+D
Q9QBMzUsNN2CWdF5WNMtpb+FHzH8nmegtwBXD6eKaBlXPCic4T7foIf5OKu3E7hF
g5Cy2cqTbqTYZkS84zpXpnwG3O5VmagKT5OfQmLvhuHBdDPI412TWEZWzoUjrBC1
46iWUZ6daS9EOW/7A6qL6GDrkb1y3ahdKq/mtVyag6h559mm/qWpQ1qnhi5koKaw
VCO51eBJMBj8Jt/E9AZ7atplSxa4JJwY/NKdJyLUdawRAc0rqeqB+zttXxSI/ujJ
oXo5b02bcXsQ2MpXZFfMJOk4+McRW83WPmgZftRwym81I6JPWWBGNNiCo2f8dyQA
W4r21ZQdyErBCSo7BuJ+HD1pNNStLfY/qSUD0YT4cWEqRV+S7QBVwptceCVdCq6t
c9pzebCJbW797z7zP5N9hYwBRwGwkjZBPpt2Wp0GiyM6pWcbkOe0oFEbarO55mP1
kKUeBQHkubvoXdZpEYUwDy8yBAwCEsxrwlY/gC+fvKWwLDKrv26a/MEIBOs8+p42
zvnuXQmxRZ8ZGhbMPoRPQAwo0A4J31Nw3Wt81ZGOvz2mluKGk/hgjIIMtgZodrK0
/wn5qDJ6h5GK3NjPU+ASPDxnrU/62ocxe2FXehxuz3x0OrzDBP2vR56bgxmdAaCG
FRGR60oK/QZ+UwUOapZSCVMMsjuu3Yi3HdgUM+pPXP8/nSUrTP17FSoNPCTAiGYL
szkW+hu4QwtyhYbmwVLySUwbn1bysgWhnlrxcGCgJhcufz54/0vo7T8mARQ9gg7a
4ezq9J0qCz9/Jnh405sPV72ns71EVJ1EzKlh1w04ZEDV7HTLMSpRBQMuoKwv38KR
B8rXSFKRx/612FOCrE3iBezkcqrFttkbI/ctjFopjiVP9hvV26UhsP/arIu5KDRL
GkYIh1ORj4dpX+VFM1tVB1HBaEQo2dv1m3QnMU+tn6OS/3u64ljHsi9aUBELNu8L
sWoI30IxyD61nSoK259/H/C2cx/j5yWUGKOdBHj7v4HmB/CeBNJ469ekF4vhIKvf
OjtBMeUEOv5Tkb1in4iz3kVK0zB+VhCnCLnqMeZpqNA5cVk4Fv6ORRuE3n+LAl0g
NEoBjliOl1mJtbLgK0uw3J9ozkdJu6wpqZTlgw9bl4G4vMFDRN6tem2ybgtlfDRt
Wz6OETzcoZIXJWF9WU+164TaHI/utl4RrLiDL8uEEQjGRbZOIIpb1jkAgIXGI+RW
fHb6249BaWbUpCrAgpDfdkUGEeNwChMAjvq7INzN6fNUUTP0CTIaiX4fflCrblql
nnmN/xE/TUlJ8Fsbe58oNlXLLRE2IeyriukP08OXd4jMMn5Q9Qce2snrQWyZTPDp
+M94Og5u6Ng3Sq8wRDGCw1PHJeNhH0RQdZnLQ+cxS7fxybU1NdImfOCpLUwajsVY
MwG+XcwJJOtwK0XZafQvLzvbzcM3ujknT21DJ3YUk3OmyS8Vhi2lse5K16g4xyxf
EzTWsxiB/TXy42d6ld/hdTX8HwaoZn+WLYpywhXprXIgK6A7UBuNgiJ82c2EBOjt
ZaZxojM9VOax2BOc3D8mk0QpZkAF6xkykEmlt0+6XWLPrUqcrDvHhqHjkrok5rMz
Dd+hJ9CmdCOLhV+jlj8E8KoCOgAAxpXKAezFIpfmDBRKWkLkrqnltQ+sIWakCqA5
d96Ppafww3N3kL5tTvxCzcF8W13RphYFpdCYTrXHkKhtwUgQAh4/Pqd8EjbUYXPQ
6F9dxKv2QVBAp90bbrG8fyfvnvzcdLUbu+paMAei2Zn9vgQvWLH6Ds4oXAFZ8H87
lS+uh9QB4zBo1o4AUUd6eQ8cxSWxji3VOIRM8hih6lswqafCyBUfcapyo6onOlF5
nzRDTOufFBb4asKnEwgHrU327WAGJlx7OOiNWzvkEcPYiCRwAf6JTFCyL8GLPQ8D
HsD9kF8Lx4HqgOUqrg8DIjCxygC6ZomKm8bkhHq19IcLnz/ERa1cgefH0Gln4ki4
mYuIzWf28B605DS0aMr+8TCHBtofE4Z6jbNHM8LOaK4M0Llritic7rP6LjKICrU1
QY4BV5D80J2fXUDjhEzoWRhmb16bphuHn3APBt0OasRLISfOgBpQczXMaC1I68Kb
lSDMz14oadaiprutkiCNPaJ3qqQFy7cvaTrvSIRXKu/SjOjwcMIT27gqlBtjJFOK
EMwqQzGiN7hPkSkaAm6XTDQHX+rKuAUb6uL9Z3tpsDKnmU/pXdj/1Sy0C4EQf1Mk
PpITbNyhFPMHWaj2w2iG/zGasf1hayLxHmCEWqb9v4z2prMmmXrvqUlsMaWhJTG0
kJNWT6oFb2fKzz11Cxd76VAjKR+C2ADIAZzAF6Ifekb3VcsGApSc7SQLo7PG5Drg
HP4hC8pvsR0oG453x5F4FXOKh74ceAeMPDmINTe23hWC+5959gOfl10iQlEIeL83
xxhU7xZgnOWV1kr60CYOII+B3TO8ZLuS2HPqGUD+U2tGpn1tR1gobsa9WBs3VVeb
e8ZPql8NeE2VdRWcN0fU2acfCDh6hfF/w+LOmqKC+bT/tVHC7Xwsms9o4fe3scxY
6cd0oUkYjfl7oeS1ubN6avsIPdA6GwWcGAHNnm6mD0oOamcHedjF4xx2jWfwbagg
UVNh4333IQeZ0Bb5C5y3fKb3p0p+guavn7/ychuQeM/NsnOPnkSpj5Lf+xh7kuOr
Ta7kNt9Re2eJwg1I2iIaQs5lcARj/cOw8W2uKM/4AOzjdRbb+hJoAnlQ4rUIUOgU
569kpyAh0IEvy30GMOqA8LNnRpgkPawEsTAh3fsS6vYFsqN8LTtcosXnYGP3+2Rl
ybuUKQOHVD7m9agHDth3ddZi4pIYHJ8sNa/ryWYU3GV7/riOUAfzSoxyA8wbnu14
JsQQoLHCOASt/cXnwsdnm8OWiHRh9ccfHRqxcwRSsIzQuCHBVeYLMXrae6/tEAJk
KgZIxe5E10hRjJyDUM7GGmBdxJ826TSpV7QbdsL2KF7+q5mG+FNGv/LfZXmxUfDS
GEyyRAKECu66H0fWdSSDDWJ4Yb5w9OzKqcmdI6+5i8FlWmdVo0tAtSnwUA+o/CB+
p/gnbt5P7rTv45pO7HMiVL6JeI6aEu/cJBjQ3WJCchvewcA/4Nbg/+rzwJm0sdsU
eiiKWQUe8Q8RFksMNzmA2mW7AKHbP6DtI2LYxOxm7igyxXErFgMlWFmu5xqP5dG4
XahNoQLcvby6Uj0IW5IKdK0jPKh8tMx96s7OX/srXWeOfcJuSpkftH+0bXGgNELQ
UiDtQCLGfeR8toTYPuWn2HWQMbW3hWVzuvGlFjLttTiA5V1V6pSPb0aCFDT37q/l
mAPO9hbq+s+uTCxiKLqh+Gts7gKIfWlZBSIttU2Bz2niyu6mPkv2c8a4wlRg0WQZ
6q1R5B5Tmi6SP1W5aHw04Zz9UV1GwcwtDns0mIm5NO7Tzxh5nVZbk7bukrsD5fX3
ReMYh9ZeX4RZWVGuJft021rKLWd5zg4VWB9BZLzLsZxr8cXQiG/F5U1fzYTtehmp
tWNyC/dzOY6r9nXS3W13S7pWSHAyLFsWl1N2rhdKO1hXPCW5azVNcl8IYeR0EiMZ
kfqfYTuQgxC+VBNMDCYSkIeXdsUhOSTz0jXP5hfLQ0DYHnKKTWEZcUmnoAqXN73g
62OXLfloxAB31yI7ujtAnPnKXiojSUrE5PGH4w/Cfu/JfDpoVfBF+515gq7o5FxW
Cz7cF5ZtvpZLbl47xNh8CVltIb20aMJi3ZxhioOFE0JifCj2bUm9NVtWcP9bMOpQ
KIq5Wx7w0rYkAFfhkC0CQPM53JHPSI1/PpAUCdOWrpWWqDMvaxEAMKfCC0NcpXNn
08Iw8QoPPHWTOSwjW3Byqt9STMVJTj7MT1pczyz+f7Q0PdMwDAcZOjgVX6o5Hi7J
aF7IBwd3mxlgKzVIfcvHukpT1/oBr3BryXdq76OGM4tooaRFPL4SJNl04L4Y36IT
E4ruUOFgkF46zqaYjUEiFzn8cZRQ3Hx3IxTAIkHiQC/4MIB3AzrhUmqyCAuNyIyd
AThNLKv6m7ix8Z1qumAmoLtuROPoCI477Ekk52M/f1vOHqcL+n6Ug9wpPvBfTg6/
9zbndivAdGCy9rg0RitqUWrsXySFrFEbAb40NFAxhfe+eSZMNcjTO+hyJNLzf4NC
qHENaQ1IL+gud8Qb5ddb2J8Y7xzt6uab6xzsQBJLRGLaTJmJ4e+D/KlAnRdOm0/T
6CX+pQSMtVzX8YhqiXW7kHHv2xwsM/NKLid+QY2xTx7t3dqDpIBQnMGK69wC5lZ3
VH7IcZyt3ZpkM/TjfBojBdi7zltX99oRo+4Xkh7DvsnetWEIAlRA1X4LwKF4zCuT
HkN18uo1eftS3p91exvDkLbA1Z0q9L+qnufBiJDcBJC8fWVzTt8+pEu8lDyZxJ5p
LD41Ri3P2djrzNUorrDsoMKH06gE1d1BlyC7kSSQYARY+0uJRzMKmUy17qEBCHBC
W62VWvA0cNUprxEcUS+n5ebG/LV/7JN5v4DXyxGjlyRWvmUhN6Ad0znmvutASkpl
WBuvrkQPH6D67X3id1tPfFdtEAE2BQ3KcHdOUmLb6d+pA/FwM7JvFci346QS21nN
wCNXfeCJEkz6toU451O90v+Zzj5mFzqfyGDxbBofRgFo9q+AmFZYgYGsRh3SQWQU
cpCPRNHAx++gtqRZeVZYmcrtdoJKJ0SLN3W0oX92uzg85/vWBdtd3+JqLYHxCrRS
reJBzZQskODiCNCwEIJOdbjRuyO3P8O5lC4TftH7u5pwGR2Kwp/N1B0vfiA1PKHl
RZ0iYPYPwl27xsHbf4/KfOU6GMu46YrMo5OiT4L8XImk8KhK+7fKH0GD5vnUUtfC
m2017ZknwF1a1ZF2JIEzFk/bvoZ0jCbiLFYGMMfzgHI3Q+pptvqp1sFXcXSGqVRB
FFdkwYLeJlAH62PUUJ9VJMlSIp0b5i2dzmtTu9vLBcBjPW3Pe+ZJv52hZyoyelmX
LhRKim/47hxVNCK6iFezQ8Ifbrsn4ASJAL55U7DMr+CXhZuFXi8a0fI6Y9VTrDW6
sMJfv/tWTFy7TzqZ5NImXx0EXKltTVLD7w3pEL4hCLNt1MT3H9dvkXD2lepSxiUJ
wGkzBvaVKFqLGa7L2No4dr1tvwIlMtW9VfGC6TqeNGwDqFxkX1J3Qe37mH0ff1YJ
osPT3Gg0ZGBXKKKL1DBP3O1Ms37e113/MN6BkZDYSCzgCl0ucFPIh1ntjbTwt8KY
qg/NwqwLYabbvs3deJQEOSRMyeCRydCOtwZT62X80MItA3S/uvH9/wWcTZcTT7oy
IdNguly9chdxvut9GZGFiAPR5BjUrQYSO4apviZJwYo8eCLJ8uQOnztvdqhN3zsT
2dcdwCr4V1iK1ia32pbR2Sse8xThZU9ITsZ13OHEeIPe1pqoRpDvZDmaZw0WJmlU
h8Wwm+2AzjCdltJA0PviOPDi1/UsjeTpJWdn+ah37G/j96KJ2Qup+I0wmL6iQBq4
arZMeIMq0bewlO8NW+DdRQeBAEnjLG4g+JQLNBy4HJmFpzKHaJeTnbxqVUB21Zbj
diaYUjbmZ7sQOKvJ7aAVW87a01LNBikN0dYMyeRC89qdDag9B73Ul7Xza1ZFgDno
sgW6/j/xHSNT7tUXQU3B99cacqUQ5xrKjLyzFymdC4iVgQc3Cfe3rbJpa7jeB0DQ
e+NsOUzkQT+86kKDQ9jJRRjyPixCjS2/reOUUdUUKC42kqalZ/t65WEcYmeqjlAW
Xhxh2cuYswiK/Jx2Mzk9XB9DBUk2Ndv5nMmBM8ZyjoVRbCR7P3dFAAcXNKVB1yc9
WjZsZ2tVGXISWQo6USoHkY2QoZtYOA7lBrx+fBOzWJAcdFaGJJ/XeYSv++3h3a6V
9lQ4J3UGIbW4Lti+itz2x/XO9s7HHulKZbCZNLkeOOAFVzANzYdrx2shDtP7tzAR
/fVKV+pcXcvehVpvRti3xBQyWnZTngGS1vCXeAf23VWZpiFdt059W0yybkAdeq84
uIZ5rtrC7ssR2hD0qPPKmDHj5DxfxuCTf04oDhjMja2oE+WxngvbEMusFRLnRFYf
MjzQDTqaZqyKfjThMD+eMF8DngMv+I0ktQ5z87pL9TL+uTjpIeiVKDOjCY7tjup1
+mkYPIShcZwNcMKqtGmCPMsm5FtR6hpOasPf6dUapOMJtK2D9ZO26IWJPobbNvjm
HX6lstnT2ok7yFLwEziyDe/fP2TLjoVuYyRt2SDVtLR7MvFdFy6sUxeHHFYDACNo
rpXiWzEI0HIpPzGc/LogoC3iLQlmbjv3xgud4H2Irh+/gWkiYf9KROHi/tHKU6R0
onfCTAU3OBhRMN9efDdCBLOt74Kdid/IOK41kLmbUYxDq8vnLZW6ibYUQfGrXDzc
xfWWt/HcXbR4J0DHiAEBrR/xW/B2LZaFqCv+FlN1c4sIJ8H44WEuApjo19nU7UPE
3IDwrJjaDPHw5pKmdvIbwy20U+mhtUdWodvXcz8bKs8cwUHMlTxmnU/XCkpDSi+S
PcKC6tpFQVEWkcfw6DYJjtGl67QD44xmfioj/7ciYLq+lqyiYiwT3jODGbwtlzHV
ukFomKAEARYhMAPAWi+FT3gaKie1lOSdl+1Hi4pfyAplXhmJ87hkxkyBS5aC+mte
uhuna30YHqclx40n1F0rnHDxHT32eRONX9RVOhCydw42x3nBzY0sGZyW2ADaOlGQ
+uDJEtQDpU1yASPKXuG9u+a9rR5YpMesQSRbr5OlsxT2T0yXhES/jdzi4J5GJjR6
ngf2Yu+Ym78vGOFRmiYGYUTSYV7qRqOieYEWh6rQ9MAUo/rIOuo7Ot0YLz3BgFwe
AjZAFeWLaYTmzpluHThaAlw5UTjVFtSkmuoA5LpGb5jniLaSqcGiIMokmKfIfTrg
FTDtGRmMdbpRyUDNBCZN6reBXA7CT8CbAfRZffDm3FOIhMuwUjPFg+Lhb9QuL1Q9
WuKl7luFLXFboTOhM0tHIHJQZZwmwLSBoJWDxV/Fe2WcSBfVlCZrCzCYxEM4EBlN
OkwahTup3ailg4hxHoaA+BbAFnx3gqXlfrqYZWWT3MZdJKevzCd0p8KWAvS7MVoC
OJZl06Adehp0H/tpG8YCJDZt8GqWlfJIMzG6UU/F3WukM9zwGV3ZzLFhFMaHhSWy
jOOeyEVN0Pl3q/amC8RKaS+k500znJpe2jzXQeLnZX75R0BeNeDHGeTvKwmoyqyB
o2l6PVUuJ0jXymKkGN+37CTxmm0XIDRqV9BSzJNG3lsw9hU0alOBozN9LbIGlS3/
TmFFhB9jQbQuf06Ym/GprLWyHXvJSf69OIoDd3lNmBPDfhIgYBA0+8k/iy+6YxFl
zjfP1IIO0m09Y4hGHfm465mF2FKT0EWSdMo2r/Tv6CInhZBRfrSMW/lNXswbDYvw
wI/LWVwUbqpYD0nATUcK79cEfKZWbbC+a+G7Q84N6Vz/tz+khp5/KfxASG3ryNMB
0xwL4O0XMFh/PLaSPhXSEP3wnnDOBwCsoCxifH+jcj5Bw1pxHnhzyOgZ66FWRp1h
aeeJYhHSd+Y0O+6eryU+o6vmL5n4zyieI+4YlOJpKCguO8/rGuvT+6ZTWzKp6tje
iB2hsHVKTsYZmNkNF5WPfT20CMSxnKu2yPEkCacJu4dd0lCWuyG0fOzPWal+kEYS
2SRu4EV0rbnFDPBwr61EJTOCTdNI9LxyNwosvbXGAoNdq7YwUNda1VF8ooMa9Mue
BcEUrC/eCS17ESTdWol+1UxNr7BU9MbcS40585vV5MBL3RNxyNdCpk0VeSkn4EM4
O7gITsZMvOQ2RW+pEVqYyhvyaIek++WpUmqFihumIiBg9SjAamC7+4SK95aC0T6y
mKRKE+FMwKLGqDIORVeXPfXJFw8oUOvf2NYfc8uxe2FdnhbLBqs26Zu9slPecG6W
jVuuUYpRaIGai9aDp02dFAGDIy0emIbTsC4M4kHVFkDIpstxtS5EffQZLJRL9+dx
0rKAJxuNTrHzHLSDjbmm37RXpZ2NZ/lOhCZIhRPgnXabOvfIPWFhKTLCR5ooD8KB
kKjzNlkv2z2yocjm6YXodlQuGzRx1VJTo/NUrM17xt1V/leliv6AAR+VJbM/Bh3P
E0yzLNdZUWHLYTtUy6Jd2Z8DuPu8SRy0JTnGJWjGqbnGmur31crI2NJHchDyGhiZ
emA9V1GhcC6X66pWiB37x0CNXYEx9U1TqV4WDb31v5kYFTyRNF1anIiknDOjeRZD
5lxrLmTVkyqim5pf/v6nC38CtTztysn2CtktAAulNXRW89o/EW782d1IT5e+d17I
zNRYNu9vYAOk4c3mRJlGJAbsG90pHrBiVyJCbqGdhfBVrT75pDAn2djwvCuLTdnO
nC6j16lOiWEKH/PF3wKhhpI93Oaja0CdSUcQCwLrV29if3cTe95Y9Mi+zdtOSAFC
/7lGsT31D3QHqWaWusG++9qlulY35Vap2ZSKweUxtW+sIV6uyFhkY0m146ho4zHb
Whu7/W9qii3+QfEtr/yKvtK71TESMz71hZIFfSUf+9F5ofx0Qwui3/NX/1gQiycF
De5lbpdsL1FRsFUtJXp+9UZOVvwVqG3mhwj5vBZomNxdg0ztpwkIVGvB2ll9v+AA
mumM2zNZ0PRR1jjbwq3frHalV/iHvKLpVmKZHzPrRhErpsUJqOHs0fjbGcw304Av
c+M4F/1kyr4nsdLwtlJDow9mm4vUvB0gAf6EL5loVej07Z7134y/wQBU0l2flGJa
4nogEc974yZV4b6FomU95Kna/4Fd3OpFLdCjSX4InC88X0qjHf9gZO84fpcFjeBd
a2XfX9rPv4L+uTR8poZF3cRQ2b2jFgSGfQM51DlEJwme5UjSXvFQqiihDAPSxxIj
5LwvYTN8U0rJzHrZLGI2s+mLdnJXnFMtouGY6LA+T6BDlZoRxehxKlNplwClyZxQ
5FwwQ4+kZ21Yr6rl5IBgrAheY1pdaxD695NyGcKLTGGt9CcEnk1Y1pBCgcnK45hs
J4h6EAovjdozIrXm+1viPnCdUHSF6+mrTKwfQ/ozm7YuKSyjL44qkd/Prn+Dk7GR
EwFKVctZFHMcEjzEA3Hk4rd+mCtcMJkdic5Cs+wFy/PUJc0PCTn3Alq4XhPbrETt
bZNxtlndPtGC//nLSIRnye4Xovdz7TuzprMQCMiWoPs8KkbmtNQPKf0GfjrvnSFr
I9wa4PXKREVEapOqAvkQwghWvH51UUfgwW3o1wKXa6U0YYxVAQWyOdHocOC+nsLY
kfYU6JSzIGYNgvecQtqWSaZW3Mmk5ThWvn7dXRV6hL12gtCmtk5Hyhr4/zoUEAHK
6Dj+lPRkNOfwUdyS6BSzElVmWa/3iHvzxeLHmen+VsxdTQHilkzX4I9tM4rWq5kH
Z1yZ7DduuI+eU7KsgL8gglwro56su9vlCEcWZWjdlWLZS5IHOUXvqsu+gjLkVLjP
clOUIGgr/6G/1hKgYiJXU7XL6c7b17WM+RDEsveLKh0viOtQ8GH0XFLi17/KZZDA
wW0namIZc9L7xnl4qhqkWSn7sRBvP8Bbb3v79l1no5GGJDfLDv7/TN+Y4m++6cyC
DRILwmmL/d6a3Sd+J1BaUpO2Kw9vj5h2+UAUGCjk3kxyAKhPULW+ZnvSocXbfHRd
+eD5298xSTr+GEIIWVeeRBiMn/ju7ABKASdvOH/dlJJncoWJEnNN5G0emCPyxcvE
+TBPr5sFqzUHX+53KaGcVb4v4CtByiv+Ow1Ifq4Yk/s7VM60wwmV74QYaMByZIBS
TCHshLe4ozDDQJc8swmz+KVJ+pKcSdxYYbMZP4BdJVd//zibgTyM4hJjt/zTTVBJ
eaQVy76HfyfuYuFdvcVIiB950Znt5kcRq8FYWq7fp1Y5s/UKcdVMzUca0h41LjNZ
/cpvYE6ujX2VRc1pxFvRr2YPkUKdi1u02X9zI3rRupAET9qeN5tLPEQ1vge4GfK+
kNryrCBMqCHoM1DsIftJjSlGmcB5lUasej8/jb4bWdXZLVIYZE/LUlB56AsVgGyA
YkXBWYptDEFWgOzBXeYWNiDSFD0UdSgMJ7RKyputKIU423fGitjO1qS1MZe+OcW8
S95+9DNA3jnyy9iHt2+gWfZBUa56uWx66T24Um1t8FGraDAx4pVEy1wqj/nYi71h
oHB9TW/JY9yyEl7GDSXAZxfLI4FQl73FKja/SJhjinAXNYtaauq88o5w646bM4zC
E9vEAo73CLRqQ3qoxb4RhkAgWZ+KF/DVZUbPXd1LqKr2E/fyT1WAQiAgHR67FHGR
hlWeRw1YalUxDgWvFcswM9U6Ps4XoALvN38PsPjt1432cBhdk/l/KXEuCvDFQ5jB
JTzWD3X3XuVE3mZ4JevihqbCqP6Q/lRlCCkV6cVPQUl+6jye2736iASav6X8Y1bS
gczoShygEU33xhx9V0fMj/GZtS/rqmHNOIsS83M+q90JdL4AILg9aO8VPglor7uF
FANNVkodCGkx84vc7oK/2zJnnWJpHZFVM+P8GfN0Opwpudl29MFxs7SDDCFKWblK
4U46+jtZYKelKag9VZobemENBV9mRfm05erR4RTlI9SavCLX6mdMZeOPYJVlCnz6
0Q5HAU2bYysPIVZCmrkvRX112QiI6fg3aY974jVrZCcq2Nj+5SDs/o++BBkbdUJq
aN+MHhbK55pL5nKWh+55+2Aj3eFsu8prpagLEhBLYAWMxJlQkEg0LZq/G+NRsqsC
DAsllVv13NYhlRDHustduSjgCJ8SdYq/hS8mc/MBR01VWy9UQf9AyC+ZCTEqCDA1
miS2I/EqByDTcBnNxKWkXRk0xXtCS6l0aCGZULZ3SZnBJZnZPaBX3EUTRfMD3cv8
GjPWJ2AWiSBV7Czzjz67/uXvX9prVkLoKLIdPHiI7scSJooZsQnMsL9iAdsM9Vef
/WCW1sEYTD1QVbtJTtJMGNdBbKGPUh8M50tLDL5FDtJ5A14Nu712m6sjNdJYn57t
OVVfJm9zLrYTrpZ9bDdk30oFyp3NEuy0LuJV9/iRa0KbB7lHuM1AcPZr34qDmNGJ
Iwq8DQ2QIhPVCSKFKvT/uvIWpBmQZk8cZ0JDH/ho08no6eNc5PQ7RzA6goNUcXPM
qZRBu4nVNIM1g3C6yBAiZUhlD1Q9i5cEm5yHiTuZzlyHWQsCXDCvhZ76I2hsUtiD
gY7F6cXz9/Wo06nlytffxtVW1bWvZcqUuAxQbcBkWCUdW5uVHCpCevgIwIXZbzA2
7DxpHqhECkhY71CDAEsEjgUEkMH3qOroxHyTT6cjwUKYaiUpOBkocQEXcwEKqS0f
dtKBnhpmeTligBGSIYOnSvphN/p5YYD7BCTapoewsPxOTZwlTNeDl7pF2BPLRH3R
O9ZFIoNK4sTg75aN+zgJVOUwbZN2hGUfd9Eltaf66nVZJ1bG1kGsMJmX8dSY2Nno
oqhUqzLZVeRe+DqdpYg/lJ/EqvYE/Swr7wm17CrdVdwgc04lsVFKZ57xkjSB6YzV
rh2EIiuBXTcjEKWN9MlGfb1D7i6rFKsjjCJavqebVY//p3x9LquiFgiLY90bvTYD
xKcqHk4Dj9ZQWiOhe8pt2so9/o7jdVH9OookkeNhT0i0u3mdKl8wSD9LVWvAEHlE
HOqx7fbYDtcWohDVvgYbmH2Hw89/PPMijhs546kfeiOWqqzlbY0r11iYVArSK5YO
Gq71wvN5dH9mV2J6Yvoxibgzg/HwGa9s5PItMCqdIRR7xklYnS8wKlzndsZNTr1K
7dK1rV1/if7/k2ou921wz+R2tbPkrjdoK43673y7GH8kdKAlMPl4TP5MwjDiDWcu
jXTcMYQDsto6kP+ibghruhOAheTKDTaYZLAawBYw6Qta/0rKSVODVy5smqHuckdQ
lGV8KIPZ7M20RghL4+bwY7vXLcMQZ7npz2c8TdJCi3xxvF2dgkJSV4IZesQaDqmN
Xb6yTWEy5hx6NMTaBgx7cZt9T8wyRAK5sixnBNz5t0g8lSVU0fx9lqdYyAg2AO8Y
zjJpKuqdLvetIifmvVZAMq7dVuW6VUgFp7kk8WGFcXzwKzwlv919O6k2123NA5yu
STK7fk6KDeU1jmjul16ew71wcQZqCGVTOAxbqi5kWkc6JUd0e+FpXtyfoJpr4H4D
kC1KLoTV2GeZ8AyRwqA3oL9CxSFad131YdAhevcDVVqi+tVqMSqKVwWwOcsR6qvF
FaAFv+XSJk++3TPOzT/2+F+KejYlh9seLfVxjt1/IeFa2D567pP8JtH8ZaQpfGFu
Xi3EVFyF6zQowuYPjw2VhxciXD6hqDUCBdiONzBtBH/wch2PfHOvGJr/9wuWZ+Wc
6IF6UAgni8xkaCfqPaxv8+dN7Y29/zmNKqqCSVven7oloUElXRsk0qXzKUHSqUBm
M12pBMrkGx9XVajFpeSb9Jq92pf2J79wTNvFjES8ce3ZYPnSDaPWncKKpVu48Bgw
8EJcxA38OyvB3zQzEgKqk7MzNPJ9kwYBsA8kj5aJnDGjypUroXVVfhxQ//JLhzdJ
qnc+M67McwjUDzvPlTpx7CTDEULxg3GgWtqW7fKb+Fv5ZBEwv+ntsqyXFKrebT5I
oVm59bUHwrMyPnOchWXJMLNw6IQ6XWWNjgvCW9ccl/C1+GnMQwB0N6m446Z3y3Zm
ftRJnSkbo0fdY9mQHPN0KixrgyaryBIkRbClgXyNYScOdgMQxaBVgdMdeKhHuyx4
8K2P3I8A+MYqXUDQZlfA/U6+5KOBF4KNEbhyZ4PKwMGYVB79c5gcQvcW1EXlpEHW
7G3HjKIwH+qlU5VtA2dYKK/pvf9RP3T2zYxoePh5Tu/JLl9zQT4F7IjRZYCNd+jK
fFQMZbcSGI9rHGkxtqiSH7GtAr4S9eXMpOTIhvyq0cETimG/G57lzTxkxLKiSbIJ
OGRxYKkxLKP07+58kaEpFvqeghJsQCVT5i8GH98z4tZIIsHG8rhMUR3DlmFX9ueY
vPModEa+1wbMeO3Z5vFvFwz3Nj37qJiWx+N2dPXZFHBflV53fyK9eYEuH0VULYlS
oXrK2gnrNBNflmbl9JZgLugIPAc08AMB74WlvpMdpoVrTA0exAhNq1sqsiOvNkZG
7T0700LE4jvKjG3G17b3ECp3OA5pMU6+WqqTL8qKQTXiyQ+yfPCBK0eiCV1fdQRC
2oXq1elLHKQ2TRCp3dCktMh8jkojgEAQHLFh4obxhFia4jxdG5fGVA6Cqh0Rxvpn
HhQtmP3fkJ51rhsgoHIeP7XEJtHGnNvnEwG+64IsLpuuncCDJ7Q7QK+dDqenJxfw
0/nNlZgnQYZMUbl/iWoWYdKicVkXRE6q9eDsKcmELJNNaoT6N8aXmAV0a0/OYi81
Kh1XJE2HG+doqKyo60omE4nfwSfiKM1CJktbmjdtcUZ00+TMkrsA5HKzsAarZeEd
rShiZXK0J36Q7u1UsDlzHqIrBVjV2lmFd/owO0xcFj670AogvenSh4sGivs4Fzd8
ez4QP1HGtlFJcz5jK+kgXDsSCtXr2zY/C4f1Ft1w4C/qIKsoA3wC6+KY6OAIk3pJ
RpWIiRyog65NBK5WZB+Eyq1/0JaSHZjm0eauW2iYm2/fbnuN7czp7m5jQes9chJX
+J3MCqE3TT2w0yQspDJiXpshHdvZB1QCjLcGu95EL59Dju1DPz13Lfwp4KXLtVpK
9/JXWhoLSeBz/UcpmIBwa2jPq2vu4qHn0v2wXPi1F9LZwQK1+nqKSGYvwjzcbedS
8h/Dk413LvhJFDCPASns7mr2k0HFMxwnTdZcu3HEp1BrgK8RzBdS/hDLXcgT/EEd
mppNW930QIVc3XqsChBOdgR7yOap6X/cOVyNfBaG5isZh0hb+63sINCAUwgodqBQ
ECYCZl/bH08AamMvRqwEf4YKbjYrCGXHbxO/voWBYOarE+sA/2nsCcK4B7RxBRkO
hbl3Y1Al92fSwm39FntLwEXcdFIQh4OAP4Z73ZFyaCCbSYufZ2bAzkJlkeW4Ib7T
kPvXyM+1iQn8CHYQng4t7K7kgn7+Znn25F8ieABFjpQlceTrkQ/3+TLU78nZnkWk
K6oXNxIl6RYBavnk67QhgGsXmPwu+QMNQREI5hykoYQKZ1s6aAgH8NesChOVbcV5
V19HMTSLlcsQ5Kpv9cIWPxvkjhOcomGjgPIK5EI75CtNbR8VIMyYkspeD3EkmWMu
6Nce1dq4LEo4CA4WMN2cCBiZGcvYvEvqBg4qmiuFRI8ioqFnh+gyzPNtOaKGKFJx
1xjiCw3xDwhmp9SiK1sWtoJiemu7/fj27YUY07sF71Q1g8vfyzgO3/DKj36IWGx/
kpJOdnx+yoZlrqyJD/YHyfhkAeyQ+wdvIrjxoIUzm0ltr0+t6c5wJdQ3qyR0cUyx
vV6LKPaZTeBWUKh/FAN9NZYyui8x3Y2D1dKVE2GWMIPrvfBuUAO6lFWuce0Vy7TC
WwAXYXAHwlFLbxabPvD88h+oRVdNTcH/IBbklpe07bWvf0UM7YfFqrmIPF552QR9
QFqVQCRsBdSW47EnSTdTzreUWt6U4Lb2i7W0QEhcpXfAEjCMQ3EB1gkmA6ee80tq
C+gR0YxHMuiYcOUuuEIA4/DLtBuo7JKYXPxON7FrkDoO50zuaw17bV76JZfL3IIt
W0F3XithTwFidl60FHROC443Ql+EB48OaBc1Hc7JyGry06Jy9xxDBRxlD9dyYNi3
kEue/mvkuZafopU7PsYhlMQdWC4e/2I1WygSj7aVAGRsD6QF4N4+j6AKGoBGWFVx
yMUGhVxOsdM1W3JLGu+6Lj6nyd/BmdD/DYKT62+cJGo/upKmj/yYkAI6h/dZh1eT
fAaJybWjFo+T5S12VRIGCuR5RGMcmFShTPmu2kZjcTt/b22Ps9Bb5Uw79IgixtXx
wPUA0gdG9hTNLY0L2QT5+8zuz9JEGV9BCI5yAXThnhzyaSG0IpzV2O+HJAS4YiNZ
B5DFqe7T8X/xf72021ZdCY9tPRaA9EXeJpnsB9/20qqCdgyf6BkaQG9wtYz15TPU
wSNwTDFwqyfZjBZE3Zsi2YdVy8pgeCkk0bK/lxipR4wxhnW95lVXXiCvJAlJsEO2
RzWRRMZVF7bYcJNpmo7E+VjjA386GYJKVHdOr5yiK+9j/fJphYw7/4AnBAatwRQE
CaX6cUxgFUCoWhKWRJSZ6nR3Zf4Mg+MQs8EsBSl7OrjneOPUF/0FY5j7ax3RY2tz
RmZ3ph4Z6TeflFxTAMCCEisstcaWN9cluyochnapqp+NWH/CB/XMs/xHawJ12WAC
fK4ty4ggGUXCvLRaBk2TaSIyJ19XHfmirO+ItrAalgh9sTEYLWqFd6iAnn2kxzAT
hMFw0wZt93WoRy6y1udMsq/Mc1HCwkAQAhhQj0xEGn8w+T1xZwH0F+I6mJoDU3ZT
UA36fB6vDea6vo829iKqxtiYuzXPx1dYaXLTy/LJccEYjrpvtPWc/LrkHNCfYflb
U+4HescYT52IQwZqjj2ivXddKjQ0gzbqJLG9oidLxS8S6DqBZpF16UG7jftM424b
2bl8P8ls7oD0mug10HKd7hWsVPmWyTR8qoGhPE0RAB0GobuEC+GxPerwYP1reNL+
sDx0esfEBj/sIcDjNuabFRdDepJSmIefAJYxdodjAXf9kwDrpI2gso6RWCzgjo0P
McVvKdM5KWkLPsjtR5MVGTkrjwSquFSYhQwmVKWvmNDXbAj2Dm2xLFV5r0RAheyy
9RIO+t6fo2fLUi/Pt4eMzkNPh0lI/yVcdfmlNNyzmG/guO9dal8ISpRXLaZmV5xI
QTqhqj7lFp5c7T3bWqbyz/OAEUm9FQVvFMpuDIFmB9aNR25U3XgK29eArkUHhgj7
Jk4NLldzsvL0dDJuZSHEnFZ3X9pHpUa4ysjsVZ46rMucQhutpphCkx9isZq1lfe+
Kssi5RGWHNqR3U5B3ZGmzGEsI0FxarXnrEqEIbKGcpLaID7vAOLnJT6+ojauFzYM
OR+VHJFGHAFzfT7vHbCvt7GMDv5eM8JgnlQyV8C4l9SaXbuWU3gPdE2PJPWGbCgT
jfkYeYlTZJ+jT9+Ilf/hEfpp1pU7G6T+HmFu5uN2+Qcz4vXvNeDkZcsP5h0Y04au
vSXfaAs5IFy1JRP84/77mBVcsACpqP0TY9fGYI8pGz0wJVCCCY+d+r/tBcum2GRt
IqDq2efK1ze2y0Lm7bJGJwGHP7V+rsbQYTSVxMNbeuKqmRqDbeX3XGpiMGoKD+3Z
xMLVC6z+T5iCCRYUutWQKbrI+2khC26ECsbJMdwlIH8PRP+08AhWrodKBVyPFvkS
8lthhKCep1ny9pL8mYpnNRiE6tzsd7ioRkglljh+vvvkow7GA14IQ6BGGZ5ez+5O
Aq2mUPw5u4tIroDWkigFQ9TSwDb96c8BqnJ4Z7RqMDbeEPz+UbrJYwUgDqmFip87
lwYce3ALVOGNlsFPRT8goAHAmBjqXZw+rCFdSItyR5/N+NTM0ehrHdD7vkWfD8sO
Qd6seQDCUeL4aDRVxuQblihRUscx/7WpG1mWWwJWQpq45wrghYWtsb20M3EQBs3x
mvRoWqnAyDLBc3EKMUQYCqfqvdt6TGgCPm/fUfcqddJVZnxIzlXVyHtG3krxbLjG
0czfC4b9I5BUqBvrL8/r8HcNf6l2NMF8IWlu0cpfxWylcU7KCFLaC9Xjs6X69lz2
hT2BgeB0+z4GZnPS4ffVG1JUEnMGSu+f71eQEaB14CFV8gJ9PAWcBVrIhvWq3f53
lTrAaWA5oVoynkkaMeK+g8r9ME3HbIoWEuNQB35B45y431jGL8TBsF4H/aCqWZnC
XCSAynAwqBA9toVZ6kZ07SViFmiAmyf+OumTIotnxQV4PexqVhX71QC8GGm+P4Dv
Pp6uEVZ/Q8Crk6zUSAhUHZEM8kIifebe1W0Bjll1hx1os7du2cSp/XUTBNtsIcez
RJ1vU6OToKv+fQAlcjoIrnLA2ZhQy7Y9LjLDZwBBhcgXFkIvXDmf0Nid8BjiefW1
p940ccyZuQ8qZFEvbrf20V35H+8oIBhx8+Ik4hnrh3YX081n1dhlWnH10evujh+q
Hx3xNjHdqWxBu5TUY9W3w7Kxf+yhFmBqBOFM0QGoqOFoY6wBfYhODNmjBXbMyVg1
8ClJ2EzmTKdH8LYqVZQDbQe2MU0zYukeME3GjWJ5q8W4pUnVzoWgRnmVfZUZO325
3zCsvsryM0YNkrpyCzmFU0LwPV12xBrXj9JzYtlfaLy8QZQngs3JjJgeMwgjT/8u
MZl1ojnKwbk+ItHPyl9diPx2etuNC5ogatr7iCgBWrkbal1TaZoeL03gzjAAgb2n
bnXLpgCJ8puOI2bHD8Op8dZa03+d3oK6CdtnNuPJ/GR0mN4O1ZXzhG7oZ/64yJmR
PTIrw7OCANcGy/arrjjseMJhchzRtX4lNMPZsxhF3AOTAtk4d+04qM+FK5yYsk4T
Q2gbIknE+yugDh4wxbnwVlFdjxKoWgoQvRoRYUox2ZgeCfLsQZ2RYDou3HBV6MXS
r1mhv3Kt8pdBGv/Z7tAaI3bMujZsdrWl2uHGqQwaciNdtHIyXdlgemztDj7D4U5K
ySMTdLh/NJH4gzwJ3U4qPeHzihNoWTvKO6V1+k7/Dh4cHQZwILtjGqAHQaOtuwpf
bCvOXFdVLy8vU/8oomyA9AzmYAOndpebNZyl7xfA3tYOW0j8mS9vIyPGtcBoKlcW
rE7l4LUmkcAXry3Mb2v8nTKY8R9vPpanmzGdsolLMwatYkuZrY/o+zKoDRg0z/2V
7sp+5FO7eFMVriUk2b4MAn4/VVahbljdPg2eKnUUaMpFjW0tCz7FU+uV9QbhHgqp
8Q0DY7nO2kaXVSCZ2WFkXQmghOMLjHTwluzCVWIVc9xn5YymFGG08tIk0KUaETv+
RslXb/fZDfg+AOz+eA/h02V7rNM09LlR/4RHrkdY/HN/fZJSyiqmc4yZHhr+e1w2
81mPVKaxdCBeiJQZxRlQkp5y6P1GS7Qu2NEC7R1l979Oo/Qip4fVyNLbNQCrWlmz
fZB2otz/4Lgz6DcrEiqX4ihHCi4JNwOo3KZtctSPYyb/Omu5t1lCVc2f5bdIsrDQ
+HFjrH/j8N5oZkQpBVz27EcUa8Q2TgqK/Fm62kaGZOT4pDrbEHE2WxOGRhC6bdz/
FDiBVlk9/lIBaG+/pzgbPgXXAKz8oGQE9HsKBf499ItgWXLezu/Ndi+RirIsmM5T
yDBFj8irNKp+WvouEo5KnOIiny31xCaunxCepsmneykOJ93jvq81VgW/5EgSALky
p9P4F6NozRwQg9WyxgsucleXHY2ly9TX5C+6TqUdYhdFhNFG0eva2HD7tGAFYknL
ODzRMvBPKOE0XzErWIkp+TwPh116Pp0KwMv3WwmGm9YKYJzwDR4bZ1/0gtfKfMxx
7i60nxShjfWoJXn28HlA5llLnPDW28xes8DAtfiSdrE0xLm6SY5ZWWXyEfNuznM4
ZTkE/ClMNZO8VWVOR65HWdrQyc2xeYhfjkiYIhMLbGsJVuAttHGV2zorC+/zI/au
WxnRAkux0mZAV9cVhHALC2TTXB0GKRw1+AD0EgC6YhxuGeLLZ+3Yrj5QTVoXdMBn
HbiADlzB+V8HdAS9hkzXd7bpxmOtXiXYHFuRypBOlr9nq40tFCy0dShRF1hP//OR
mO9/I/bk0f4AeI1YFs0mQ08U0O1+ODDBzW6Jc0067j+vHK/EUYHQwctEVUAVP8tB
29df3r7jG73YXgkDPi6yJq00/+Mi2XBadGlxcGzyLRm+pF2TExeOFKLn6ceIjiUI
RphFF6unXv1ZOsTU8IkcYs3rKdElYzMNUtnM2YyapABJcQmvoU1lJX/r8tnNIoM/
Tn6xsb7D8q9FUUudST426J3kjWSAzbodTg5mXvEIDP1ewHSOWZ8G5uGHRditGQUi
UcABD3komIK4t2UZJ9buODhh5GddtNVfWZOav0H3+aoKBrMmubibo/suURGENxi+
EEgCF3VT+grEuQ4GauVKiB/Rn5KdMdOCGf10RQ0l1INVVBQ9saq+8Y25MdzBjJFO
B7G5P5ycTXQxzqzRzsPv44TOfmnTq9CjQYRSLcUGgK2rdh0MCJ8o8zhwrePbyL94
BfCr/gVJUy1WQQR6Z2ZzkyEOca7+0RIIllenwsE1WooIJzbbqsvHbRqGmz+weZt5
NpNipLWqgDya7OPYpQPVU076gIq4VksjrM0HptII0oIPhVOql09ZTWojzb6X852m
P2dZVHBad55cUjNGlE+JlAwIYq7ROmRBZqbN8gQdf+edC4K7XcDTGMGFpXJKoGKb
mIFHu3pJ6v8O27bJTR0DW3o5+2GrXYHnxnF+Hbw+K2eaqtPjXxyx7vv0WnAkhtR2
gftZZKNe8S23BOIqtw/KCs53t/hm2aTjS9KBQvVSpwQmrnRujY0Udtvob1H+7HK4
ucgrfin3t9i1g5yFkLpK+hPtk1x2Nf5enXbBgQrByMIklfkGhoCbeMXfAPkjRZAD
si6GHbMlci6nTlMKvJfBmf74HpuL0oYZpavA73n3pWWRFJDPPI/neV754ub0XNFu
8oZSaeNlO8hieH4vTy5reEJiklqpgm8AUuj/EaZt3DTFOmBWnF6fGJymo3NHYVFa
hukZl3kc3y50oo1yr79SG1hrE4ztcY5Te0C0/YwWTk0TJBGn1gKeKF3dbLpmsERt
hJWSxd6hZsn0KIMk4xwC6HnHOa5w8hGKeRnbGlPsHb/aISbN8nsKOmEcs15RREvs
NvR5H/G1D47kqcNfo5SacMHzOC8n1WpwCl5UIeonqnK2cVcnpgpIYYCBv1riIW7u
thowEXfsBj/bg1EzXhMmFLsU6I3fUugUpn7k66JKsWl1rkfMBPZc7zbB7TlBeMrz
U2NvJaTFxgoamGNcRl0IvJQSPh8EvqAsk6z8WXLcg0USAh2bHlt46fM40bHAQeGx
AAEBPqQd1ILL80msXtmLIJcRxvZ+kRSEKseHt5Km1e9oshTY0sWJI9+8c5GNjm5q
2h94kHJKYKkDTZShwhyghZ+A/9x60Pi4HJxPvZOu6GIGHsvOAv7lBPzRqIdNaosj
F/Cn8UscwJlMreNtlocxkkYqc5tFjwqcqAz64BgAbAca5a7JlG1/S2ewcMul09ig
IHvS8qCnKudSmliOBg02pxY0gE8pvwgqHlQpXdh6HdvXJ0qwzhi9FlTFvbzppa3F
UPVDCQpTs9zRRyGkPhuFzLIgSQZID6uhUvN05w+RRbSa44juSFIKzunI7pexv52f
0AMcbzRdwGLCc6IIrlksK9dbPMCJY7Zxq7Bf52sFgPuJ/lgx+BM/LEpVNccpDNBV
V7Z1oaVokiRB3l7LG99ty7tZklMnGekor/ktkjzUHjwTWC0/jQbOPJXNMQaVGyCE
lGAHQI/rCWpw/SJL+7+zG7ECo4vlhfJ2B+he24HuyQcIxwaJSudaGXyw99GhPqjl
2WT8gi9hwplfY9j8eiVhycsQy9gPCPWmPg5Nh1nNWjVNQvN+GaBs863xuQw4vxeO
MM1jIuN+Ou1n1YJV5mRvh+freXjX4xxdT6KAqLJtsE7jfwoQXGXd+MDE7H7yRuoX
fmtBTd2sCGg+sNJZb2iaL7xV1cQ247+GuW+bD75EaW7gDBduLKKFczx7/QWWMF6R
hgRHM+EWl9XF2/C76b0B+8Kq5KJwAPob7yMJjK4Ob2gMIrCg2Fdrs7ObmDsR1Hfw
nTDank4v9qD6RJ1F2p/XW4NVmIkMb0gQ5S0x/FH5S97qNsOX430fpVxb17YphT2Q
yYWz/L56YaJN+deYk0ZtYRW+bJYYr+E4ylJt8QGDfE5NLxRp9H3LW31s13BC5xSg
ekVAIS9+98zoaHQ07EzntwOaO7oO8Wwgs3AUXopjWmG5z+e1f4+Fn7tkMjOS6QwV
DzP9z522K25u6hEeRvwV8MFOpPzVK4JujTg80cTcmVMo/1IIT1KP5tqZS1vmPP7p
FA1HTFBV8L0/Hq1Ppqm2LVicW4h1bUT7dNQFzUYovR/epQ8j6yvP+VxD+9l9cIQR
PIsjSZgpguNZs3GMpc3A7ZG1Tl7SP5R2Sy41xQuZYcBLVOAsrNkxr3u4M6KU//vK
8raNCVdjtk+T960GfxBAa1LBy/7Hb77uxhbfIqKYwNe6Z0ZSVPeQ2pBUXilCtq7p
uDNoS3IYLn3EvogG4qyDKBig9k/gUHq3dqQCzVltEoPaY71Yo7XGul85FSJfMfZr
T0K7qafZPXStB9pCSCdnZad8cXhLoA7k7F3EpkIW/yIsZuEs45EL9WcKjh5RfJsD
zoY/GZFMClhHjgCZ8BDP9JLw37QAqeyLVbxIlvKMOhHl58aA4unIKaDP4IIDYbBE
vPJzqm2G6UBe0otxkXSCAFpzgAaPvVTSaalLDCfrjVQyPCr5bEVTzkFsx8eeQ7no
wD14U/ZRH1as9iwhaLq7An9nAT0NGBGPDMxhMl+/Bfocem5km4CZeokTI2Du1b7x
V78ui1Efz1TSw0mzAM6avnOSmw18eMcaU0RVG48L2t6cFOfQAU07WaS9Y/oAG4uO
TI9slRt48RF/cdQSUjPesjH2KH2Y4IYMac1EAUgPPY7R0rXmhYdwX4SvF6pcS83N
g6eXRi7zgcZVXwc5ksbCQiKYhcj4kP7q9y3RXffLhl8Q1RUjY2Wi3jcl8NxJFVrT
leC29tidxc3VFjOTkff6n7q+ds74Kyx+7X5bWgez7nZTa9zurxtHGyeI6ceE0YJm
bzKtHXjQP8Q8/Oiu8hcGuEF9ICzDSjPTu37YhVZVmHYWOYhzGAnwbS8x/09iv5ez
nmtFdC1bFdLQTDbMl/OEv8wrqH7ELexEXDYAq3xfdzinu0KIzwlHscfPdFlxBtla
nuWTxVPDSWCFETvxtWLeCQ+Sk2NzsW/jBW2NFyBezvQw1/ptLS/+U/kjzLdNQ10T
Fr+io0VwXILnh9QEZ/1AHnLUSlAyOg+pQaTTGKiLJeuaCrR9JUjqcHdgtirxanM+
wbu2FNBjoZC/HEzovrhmE0YRb7JFNMGQTJXemKvEEFaKALXykya2yug66/6jprj2
z0Fo3qH/1hr+I+dJLwqcUp0QAa7BnVP0beONXgUhZmvHr6iaeEHSqQWAIONXTpuj
mf++2lFhSSpuuAlzGUeUON1hOueqk5TSn1lpPbH1Xq+NkeekA8ghcAciP/yFdiRH
H9PypxBgXjMqbHWLU4Jm/mqteY0NM40NQJRSA+/Vm9vONfo/4dJMCrZZ2tYhKsvQ
x3UxfcmXadJJ/RksnOJ/AP++34oAKvcdB6xHm1BK7suLTqT8oOpMyLxfYIrSwnVd
1N3hmw+q18x2h0PpJJzYABSwI9tgR+e/Oq19GWaAsrIxNrVX03Dn/GAFQ3el0N8C
xlGD3nW9d8UfcMh437TRlhfyr/pbSGEjOxbtENpSTdv/Bs1JhrbbnUg/BT/DF0ER
cWnFTyyDP7lo8mUvHmTaBKnI8ust073agiUJvKZxKq1sS0I1gjo+7t4d4Ro/vMNo
DwkSh0yPXnn7BYo9duKgccEDQZ0pJn50zQtoRdCVU50jzcrh2YbLG01AKMOr2H0k
3SEl19BneQf5Yqpzi6VmhlgHklDxCWcJL75n8hAx5aEV+d3bXYlXe6WgvWNUT+BK
UFQS82FW3LH4bOCNiQLDNqkF6RF8fH3nnpRQD8IPZtE6D+4Fuqvlj9okXNHYhrPx
PWbLpFEv6t54JRox1k8qXIn5xqeUdaRk+ntx169RDFr7C1B0QyANe9dK3WRYwM4I
NWVwE7K6CJHwzAKVjyz7+ZGyYtasG/IzdcAmBtknWyI6vHpU6G+hSHz36qcSLPlE
7XH/g3r9qi1ZA8fx5PdWW4X5GkPYjxR0s2CJAjNDvra5yuiN+m3WPG+/Fvi7SMFF
KvMaxoE/IxIqoAQ85/ZVeWO4DzvB0Sg+8+k1tdVn8hzrv+vHxA1Vfchb/s2Ez1G+
4Wrp9gGdJfIVzqTMLGetO/HnuTr0An3CmPXaolnhBLg/tyqjjB+2Idv7JEVvtRnK
4XkGhAI6KG/wBseN8xHZYoSBinKoDbBwflWCBedUaSjl+Rng6DjCFDCE8CISgGo1
Gu17XbzPAZdyUtRPMK8gOntSZBeZrvMXfaPBEJYO4H8gBUqFqfvJc9YiLgXpViXc
PBBffeODCO59UbzTdXDtzlY7wSExIDzQftwrlSrs+mcgcMNg9JOpnptDktuS32lt
LERwGotyz16Nx2Eim4LAALiAaCBaEw2YsvmDavJ91rEgmk4y9Np48yHzAhbzP4n2
e2XzSWHtcbpGN7RH+8p2HzhVonTYk4k0eUd40y+d2HCgR5xxZ23UnEvad3JEWJ8v
8OQS9/fUuwwu7B1+XDHwgWQ/h6m2jGFJKMpm2QydMymlPGYgJrTrd6tzgw/+D2gI
lltXR2be8enGTZHzjrcAJDbN95nadUxNY07Q1rOcqPyK7ejjeSf4f2pn9Jx91WMn
kOPflGjoygz35FZeU81xmXfpdiFmiuN3lBhp8ti+QjQlIqXvTwK1iL+2CXo6nq7o
yt6O7rUVs5YOnN6ZoZsz8x/H2Jx+wrl01n7hsLMJyPi9azRz8DMuKWJh0Y2nfHvp
UVW20pLvohNfDT+bYllH+cUAOHcgT/tBr5WgSmGtP6e08o0an5+lWgh+8VTwIaGV
aXi+hOiVaqGk6Rh99A6xIYmSLHCsL1HyCgWNAM6222JK/dNawUc81c7QilANbWGi
kvHx4cZ/i+dT4epWetZTbn9d70K6nhhSkb2xLdUokWTKHp9j/0tGxF9PP6JReGnR
tCv3Cl3FzAr4YUdN918eB4k6pabElcW43B3L5aBLmXHHO1byyTSVnytigpoko6fF
3AREyM9bzIF0I7sH6u4ApzBf3yvJKV3WuZBCDE6Y2tRcuLxaxtWJY5d8QkltBt66
E0zt6Fd6kRQujWtppW7GTth1YBh1KZO6b8dH5TO9jG9T8+0iRgIKJyTftR+4MGhB
5erp9IvSeN1OvQwwH3J3U7LuFg+JKZzpgrF4pYrZSWpR8zMdCWtYzdizr9a9+XhR
i8ffm4x2uVNahL/IUO4QFPVzmtNTDKt2FtxKU4fqITebn9Wc71S9TSkpH/eWzV+h
ffoxnGksyuiAHxZgtKT7Zsw/EI1AiVdpq4f8m85KjvMfIs0aaL8FVP+trno+rcMo
F5WbAlg2CVDO2dUiAIkRD5A9pocNtQMb6yIZUVCjI83397XNq6MeAyWUSedgi+er
9TQGritQMayD2kNpXAKVwNThUc0YJrd5P4pfYsEIj01e6MYaJLNC9LQhSHCtoj/+
ONvU97RzRBiQ3eGBTTOny+yotG5R2AHH77ecjnllFwQ94N5dHNFi2+wTQJxA2jiO
fyKplrk8ndhVngqQskXGvjztBYk87m2MpZAO+rNbMgGo8QpKN2P1PtXXtg+VqV83
rUlPF8HWKkrUIBcTPIcQUhsTg94SbXa5yrA/X+VZFdQllxWbQQsXnldv5gQ9JLU1
oaonYKXSv07CBVFm4vSMdvAuK64KG/ZBNa0zH4gQu6B8HtXP5yeZU7Eq4W6yOcl8
FXQKgSwAaMFUtqPwrfVTPbTYqYqcclZOX+zKUgFzQ5AKZvNKhdLTE0GuSdmhjjV2
cFVRatwrPxkPoUD7dHkk8ytrAbAqDfujqvvKj0VKn5jZmHKeJeJYf/bptNtMGvGk
PgCqwpZdUGniOkcMDUiG+t8Cse0GwMTPf6e7mjKCVu/RPIBfN9LywDz/B4rXurQi
bJFH41hKnFSMU48ALvqaOwHCB7ZY5DmHcBu6tvaPFGtCy17MmvwiqIAfVAxPS+Wk
iUq5Zcst9mBCg9q1sYAGFzurPHXodlg2Ilt+nM+s3ws9FgjbCZE+VYII+nrjlXKD
FBi0kkFD8D5ea9mEifb8ViA9yYo26DFARJ/4fcFQ2mtDdX9agfPsAvN1w3ybYBQR
VYF4sdQtoxWO2jkT3vSLV/5JvQrmlFhN8Z8IKf6+m77WitTs9eWNYx1b3RQQFSVw
ESyx4NXojh8XBQ0NhDkz0r9rQjicRrQjMCvHkjCc/rHxdTGIt7vkJyvYluFatvEv
XebcQ24T74JgmLeSTDUF3GvrJrcfii5m1iMPTpJLiogq4FqsSnrPPI+qI/GDe8Cz
nlWcIKFoMe8+MPAgHP6Z6i7MmncZfj+qt9K1NdoleKIPKzmE1Xzg+BtrXz034CeK
vDe8OI/qjHO768vza2OWC3Ilp+tAwO6R9fbUi5gyN7yZ5uuYQ2yC8HVmzlKnsbbY
XrfWRTCd99TuAFwVWJkE5YapcNYpOKwoTd5PR+fK5UPoSNEnou1Yr6ODflcDgBsz
EfLE/bIzme3kimyZAU3OIW+mAPBpu1erKJGs/uIUgtlLQ2160yaluu1sBWsJl8em
VBREpuLAAxFvfMQLTBEbawFiTgNiPT2AATaN4/nMo4bavn2SwXyRknHAgNc8WZwW
qgRcatw833CCqHj8fb9BPSXvznb1WXLDwsB7bQjBVJdx8EOmeggIuNjONN6xjb5M
hrpvBKzrOFTSXHWHu5HuenO1A81mm0CTuOic8yme8sm6hDqfNpUVKG1Df3uYp94Z
e37xr9triafawl7ucYwyq62vyNGbwk1uDBeZIfRLka0yvV/R3OYl+UHi8dZ9Bz5i
QZEb6YZPwCZLpz0RavqXTIbNBPy7iTNZQok+mRdpP9StrF7WOsU9yp4c5a/wNPLR
IhzdCuYIFh48CsIsbL4M2ePhqbpi5CrL5PnYwtZd9G0ncggnJfVFZJuduCMSMZiD
1BwTH6ocqxfFJYJIQpggqnR/yW9D2rSqjLR5JjTOMGeZa7cmv/jgnR01uksr85Eb
YVRRm3jDHNgmw7NEqk002cr4XYqjgv/iVbt1Bac3/K2tXwD8fZRaM/rvt9qQP+u8
Kq6yX41YRqwspi5butjmHdhYCxSijhE0L9vg3pgd9MQZRfsC9zW108OUY9BS26qb
/Gbb0GbhYDn3MmCuY5QPEM1z3L5Kl6FWEVVuSSg5Gs1X1lSUChFuFh34aoYpKpbj
36WfLq/r3+/jANIq7a5BtwwYe7fzyUqWt3VOsVDa34VC9KC9FF+7JBkHS6xi/YKP
O3QBDzPi8sKvY6QEty5pY3LIv/oByfgFrfo7aCtoowkOL+ZVj3N3JFeri54UYgEn
DQy67qv/ZefOzUuwgEBOLizaySomaQrv4oltehbtZi+bf4zhtnOigh5b0pzWOry3
zPQUX3n4i8UwZTtCjYXtKIQYRvaGfOURicjsIWdyOFNkFwUod7mt19l4cOaCJfJJ
lEJlQX8uBKTddl2Lbh5RZKyYW3V1LHopyCBwSkPcX0OXgOk/MndGtjm5n1fBxX41
4rK0oKfi2bdo0jAw415TS/LOO/ll9O+mM14JjcDGEiY8mz5zkMf/OeeNL4P8EcCj
Yh9ppUZgxxvHyDH2dfdVv8AAWtQ10w/rTqrfn0oGhZ6TbYc9E6okoMjFAoxVWXCu
nl0oh3nogHOfMelgK8EBuZPiI7qaCw7wetyzsNQTMX2nx83s7JJj12HidP700LJ1
n378UXtgX8TFgFZzkGn/x8pRf5MQi5cRuo9J1G0NLznfitBEOaOUMSdbn5iCY5xX
eE7k3KrcC1WK9zWz67bdkG6J8xR8VwB6pz0zktuBv4+TB//PnVHushGN3ZyxL8XN
6NeMtQBsDhd4CjhJN1duwbdpYVQpOZLfW8ppOaX1Vgws+33ER1oXrrMDBSUWlyLM
c4RoFBz97pKZMhJDWKrVQirN3GZI1m1lDlK98z/8NCrf+rsO3gM5LuFxFQkBeaZ8
V+J/aZ4A7Fdz2cnOe2WNM7kZabtzcajzVFlwexjKlvT9LjhIUs+atKkm21i+NacO
9Zzg/7h7yNbyfGAZeaWjuZAZpZ1ZT/MfaHw5CVm7tB8YBnUpWoh/DnFg4hvwgjkt
sRNO9+DhyXe+1OfdQcJ+AJNwpVCX6eHSr5mYIyt1T03Qdk1DzkuwXkZkP8W0xigh
L0gGcURQ0IjQM5nqLh7IrscmfmaRY+m2+VnZee5MKlFVJOFKAH9plx6RcU+F0K18
mmPxsjGXu1W037NYsxJGXV6XTIWBX5tZx50GB3Fx67oQAJgLnZgs2VdtugCTVrI1
lxJeBgFrMEzxyTuSpm8bTFnTXriPmG7n2TIbI9q4+zvlXLPGUsEbAuqdf+V/zmUn
IyaKFgVlqQIUUcUjv3hxa3QWPGvM6zaNL0s8e+dEOedBDRfvpY9FEC4IFgOykz2i
DIzza7RqQJX76HN6rdHelfI/P6bJH9wmFaRf5g8APSCgTJxphpVxqGHi9JBbfPzG
kkXfqWvywmrqlHZh3LcX1VVcCab5YOCGpUn8PveGXBZ/n/BQRZuIzn7PX7ECiTMg
JKD9uO90ShWSW9Or60h8f9xZtR9IzV+ZkzZA3hXfq+ZptqR8VI8wghJiJsYUP+78
2zaBxee9K/e1c7zU64PjGSTjqVmOrxzs2kf6U5p5yk6fTb9IuZcW7DygPEO5MUtd
YePZLG+9vxsezTe/Dss9DGam9rKtr2EEXiQKrABXM+XHLCp+MPTz3gVBcfIlrd8u
7D7yEmigXgensSuTdaUqitpuX33KZgXDAmBm63CeQC/8101Uj15F+5MspOky234D
oP5QTLeG4sFbiftD34ZlokInsw/DxuDjlSdwezm6il1XLeoMkBgGjnKMTlUZud5Z
edVFZI+Szvn1eBfDqBBpSJnQ3V+Yt63N9sbJE7fhmpp6xHScfQtRVxsRCuG+7kXa
+Nisp4En3mCNQETEt1EKOKUnjPKXxxKV4bXV4Z2vXHtgvC43NWD7bgW2/coLSM3s
cRFZNTrg2Wih63coSNvrfkX/6UMgVygliV736CKzcJZKSQQ/hQxTKPvzqqS10w7D
VVqDnpsQX6vZrRgSRoko26IQlep9Tujrx64urewLS2kPvlntpIDBo4Qz4UTVMFyb
KcX2uU/XbInPenMHbvxAFB0M2v708L5vEEOz1RipPoyyog2xD1SG7i07g10sn1Op
pgfmoYNqKlG00rw66TQVzOnEsyaivQxlkPtaNe33M9VUsj4n36ng8oQMYcscwXLe
coYoZmGm/+8QgYN9Mi3QpQqwA7e6pr2o4QLMlyvrVUgDQpSBLhw3tRzLYWj8Mg2K
nTZ+xUec+9ndqHeDNOh72y9Wp17c4bcQx7/7isO7CdUQH2N70qwR++yvIolFl909
QP0ZjbB0DMJ1DlAoSAlZXdmpfkbgRI1viTZN5PAeCGruO/5IrckHYw12iELeLCMG
8Yrp2xcaAVbaQiTpOP9nt5oaWigNYD3To3WDUa+Ifmhzzr0nZkBbCzNmSDMHdx+R
PMStlZtmZs4GKrSUtAIbciloYGcXQ31auekv2wfVMLRaJcR0e0w0KqNOIwC9aB4W
muNGTzjP9sBy9wSPhiVSWaOMBNi9uQq53DLc86LtwnRrxjxKfJTDqARsGlI0KImR
qouTKqniCNo3H44NcAM6inEgZEdCpZ2ekZm3BDEY8NJ5B+FjPq0lCUdQkp0+xiWN
e2IAltRJYJqdGXfPmcD9MS57GFG3gpTeHo2CUbGNIuVQ29CyoDdY6CDiJhrDU5/B
tv8LNkekC95PTfNUTCp2fY1/met/XrpeVkI/DUnnbMTtLYRzqcRlsNK3keiRPY67
/O7xUtJkzO4VE6QMbNnJbUemKIXQjoXnsUhoHkgqoPKyBb7ZlqhLDrEbLipqQSVN
MWlavURDJ8wqSRJkuxIwyiu58Jj3BRnwPdMH7gLI/D1Yj48rNai8ULAWeBB4Gf8d
IlEoa+ES6Qs0G2SMj8TJ5tuN4Mog/MfQAkxI/ZYMTY6jRU3XNew5ZsRx1+QVV+DL
awz+tMeODwK7zJ5XleLlMg3zhL/1zp9eWmgeShjLO4zy3wbWjCW9NOdf9o1SIqQA
tiKC+Y6WI1owQ2HBowUfYcuUHxBzktIMPFo5BNYrqQA1R9+f3gANSk8Zfk98quUP
S5RzzdtEvBh6eLL6rT33MG5RU9ADTOKlNTa3QmvPA1zU4067C5OrtzT+nrTyhZWn
8RwAGwzFOhh9gno23kizj7vYUsy/svgKUA9GmPg2EE2z40ybID0ZIZdrRdB7yS9H
k2+CpsPafwnUsjavhk93ZXISSIyOoTY++9ui+/g0ucbBpGYMdJ2eFYN114teZQvA
x41biSzv8FYUj0AdDDRrLDmeZXVEE2vzAP08dvcLyePp/Y9aDtffl2wq0y9p/M87
Hc6/1ckpkWU33oK+UD1rb4zZbfQ/OHLK24hb3mSDWZojQ3eL38wogo//dOH78oKm
CnnDwdURK6u1nojS5ZT8lyRl0wOfrslr6+I89G5zKidVTncfZHxGyDrFewCrGkcJ
SlblzoIIIAQS8J0mP/jVTaHbRUreIEQRKodVg8siTH+URaZg9BFvmap94UlVIJ1W
+i9QNU3ql42CG4lIwPwNPlt3rvfEfCdrsE6il5ZRJ89Fb0TL7bpaJ6buf2vuBdy6
lRdbVI7mEbcA1f3zWs4LMLxP++umvWeZ2i+iOuU5PrjyR0H2fMDRw50WoTG423oB
BDJu9eJ8AoHg/GwLjKTXNt26t4rKCvupaXF66Siud2uYKj9PAowbj6YgL6NjMB0v
nDRuzfjtlQg0BhtBSM454yOQDe62sn7BBifJ/ISEbLzgPWROMom9DZ1+Zt7bRR/e
V+JRm0wKNo38Ymw67ZqIqPZlZsrgJLJpMW4MZLZdkplqfzlSFMQhNFhoENavRCTe
uOWeDHYtwlYZSONNbET+CGV53b4tAjlwBsxaL7wh/HM2uai/dLnSBo81NEO68wAi
+ov/oPBkv7oIKHfOUjxxbxuqlN3ZzfZnD9rjexdXYbuMl2NSSKxsdcmK8X45yX2p
iRU7FzJMXt/O0Z5BQbo4Q6Eosnc1OLgOBTOigVZnulB2dlACtNxMC0uCzROcJTwr
c07N6bnZYZtl6xhn1R241RGK2xn0PKsak3lBDrRYrs8KGPKd6ENsBqDk8uzHLjHm
d30O3Mi/F8RE6ZUJV8bYhB1KJKzE4xB1CBe4lg+UNO2HC5x426atoh5COb7xJd3f
SPaNjji/JF5OcGevZg3Pb3+uDVBvTe3hxhm0PwOaYK6OTEN0K9EZQ5/KV8WPbq4E
dtZr8OBH7tprCBVY1YQdV86gLxIoRxhLDAVuoEqipiDXrcAvsYsw24StTCvScbQq
4ovq19kD4yEzjlQLZCD2xYrHvA1bVYCTY3iHa0KAseI1B/Kyxw03bhKylyRwxitN
F6PaDLaneY77EHom+Pw6uV0/kMM+QWN7uQArScqXdDnne8IFSD1AK7sxSjLIRlfy
GLygj5B2zxna7luIkB/IkU6ttbZ13C3qTBIETYSlJCCpK47X0mSO0UN7ojSL8vJv
wNNq0cES+KiKUa9XR7zzwN9QbtGZQVZDLHnb1OkWrAYlEPVKbXxOhMYMSVKCsptC
Gdz2Eg1OqgiBpZgmMAgC1e3OcK17K3+E2iACqiAJL6sArlKmRhK9oTFTdrjWqo41
qvdeBiGtGPi5dZQyj15DuMxDEbndk1mSrWctxpKjY4fNGECNjjh5Gs0hSt0UigF3
np4fmymEvFgleN9UE+ZM3IxNzH/9r0s5CldadPf3cqE/gJRXcq9Uyre4ES+ZGlHF
Zh3BkvdC6xGD/+THvPKjeZ8r0Ox1N3Hi/1H2qB24Hn+VMm12fQlkcXjOLCNwwkTG
PyqqFlD5t1PSu7Vlg32waqbXpfh0diAUR7Hl6oiel6lVD87KFEcSGzZbesAEHhn6
9pLbLNt3T8rmO80cpCCAYqupWNDFFZMzMB7htPvIWVF0258hfk0LQR7NgQljfUy5
e9+61R+izzpHeiM60iN4DJ1W9vGvifjOOhLVpypb3ViCpChlX6g/2aQsKVODlj9q
ctLpvO9YoRUs1F5fTGUyce8y1O1RdiiD74GT9QqL+F0xII9KMc4zU3q1MuVblMWb
DC6KGiPCWtth4tObRZ1AZ1CJ+/dngxZb6OakCA3iaPtrOshKKV7rdCy+2lYepzcA
n9VRMR/2VsZA3UNpa+b2MT8W4Y4ejZ+/V1VUHVIV8CXtDzh4wiN6RwAvtLll5eT2
cCvARX7Sqbf8WQIDmtWWYvx4H8PbiAfcnJ4R3YbxtkjL+Mu4x6Ch+UpuBVq4Hu5Y
CVLP8x4xIEm7zXxxvkH7rIeibfQxj5umqWgsWosWQZ849g8aKMoCwCVMhzYV3am9
tgV1cZ4NRyc5E6QYAvKXbSFZgl01yxr/NL0QMsxP4PmhdaBTnuUjWkNbdrfI+1CU
UC59MSy4cdhRmpmOeRFiwhW63MyOaUxwFY2iK0sdJU1RCrrPpEtLXHeyW4nuVn0H
cBmRIH/vbYnjYzKjqTcWA9gl7/UH3E8Eqo7+3GqTb5HhUeH3KqKlivcwNu5XYGzX
apYYSbtmLQT3EdJaeCi8185ALncV3EYWUcGMWqSkmSWm68L1xbuSvw6XOKllXWfk
IQwPjlCx2InqkSYybx/fm+YmmT2N2IzYKQ1tL7xL6gpE0lvrXpriTs/QlHmEOj58
DI9zcReHkfWQRoZ8iyDfnGC3Bm4gmChRFZthClevJEqW9ETOAfbQ1FTg8WrewoBM
rY0NCNjTU3gx4RLZwOYTI5hLnq2RSKBezx//wII5R8X6EUHJnWQnjdWqu0Cu/VeL
xpcgLbDIcw/0zTHHAsy7MqVHOreDOgFxoErun+3BtlI2GvgSG/4ozprGLhwJNCgj
3m1JUzcCe/o4Ue5FIwLC+drKbOQlb7SqgvM3qGxUlfc9mmmyuGGdT++6OxPDG0+a
F4AdeGq/d8CI7caxHw7uTDENGNUJaD/pw7k40vTuzY+H+Q+/xWsTcAq9+CPJ65Eg
JLP1ynCYBykqhjPyaHpQ/4K9He3C2EA/sO8b3P634pEvCm4nMRZ2u+PtrVYmCSja
Opa0f7zL82jMQpsJfeO1lYDwlH0mdr3gLbLEeN2JWFWPNfnNh5QFKW2+D2f4+96n
sGZy5Rsty0RSiKIZRFF6rmNgN5LWoMYxbPNhKtwxBE6GgJ1Zv+QAHCufpi6zpXNq
xcNNYWTrUh+6f6oFk0Cm0YniJnEqxYMkxhDdqC/s8Df5RdITOFYv/Kg0tDRX24XC
4ZACrTZebvkNKkm3hAttvs0BZexzrli/Z9CgjB/DcpXZxuHofo3wBxBH1bWyCs5Y
4haBaa3gDSe7nJ4DWYoM9xiuXl4sqng/WXqHGhLyo3knw6WgEfdXKQsIeeTKGHhK
rD1xqUxjZ6L3nDPeWTsCtaQ9q+j01c3rlmZG9gLQssobh7mE3nsdR+Qi440/Mf3u
WMGXt6vH6wPoDa36KWUiyenLYBd1a6r37gD2V6bqZDslvoz6hbRJWobQvvbkVmJV
BMEhO/BU6D1gDYp02Rtu8EwAfj7iB3EX4O5eJh6GutdDWhIY81gtJwdj5JATihCj
CXAnu9xDMqUKCs04Cyopr30F5YXUL1a93AHand4tDbP66QM5mgFNJ/lb9TCcAplS
jRVmqUcHk7yX/juGpKs4Tant4pBb3QOE5F94HPvauuVmc2olSkWuynrGVThoSraA
If48TR01kFapgAZsDXZPuOQKdC6EXot0Z/XtwKSdSBiZVsfwhTi+wPcR+0que7uS
JbJh00DuvB/uZB4EhsMh+cNZmluDCYU1NtSjiZ4XEM+O1jD27hvyizVjTgX4VGUw
XEhFPnT0XtbBTJFjtZH3cfCdT7HA55Xi6FpWefNFuVuwreedftLBTuMgAczM38Qb
pWeF2rSCPVE6jvsJhlNRkAEJVZ7dttQFwCpzC7D1suJr0q1o29Ysktb4KGfrPxiX
SZWjoQALxwn7XUH4VVE3sj9dDsyhVAIdYKQDxxqrqAcFjrgJymkNSqXFHgnyPba2
koX80eaTAXz1zSJSeyCHy2FOTDGfQ9DXumhB7eScMwu7HY6wC7GrZF3bpkP41Du+
BI4UIAhFFHqUDpkvMjQBHzOnmG4NJd3SEemrkwirsOvEQ2fEB8r3TY8nCGYzi9nf
X6/51Pr9GLOgDAsMahWK5nxCsequfuvhBkF6aANmwfviuOMIUudF1JVCbER2/9vC
ajPt3t+eK48zbpuVSkpQqh/jMLxlV0UmeW2CPmFSckKIGwd1k1Mf0RPkTbc5LFZL
20Ti4mMU+PYq6mSQmkOHBE+JOOWz/iUvzigwtSQf+FeON4Vh950tBYpylnArCGhR
9JQH6ydBvJM97vldeNqupv6KSxykKr86+UVtzg7RhM4fKSuCXqQFF6dxNwfmi4BP
bRtfO93Hoa23SJKt7Mjn5iqkER7XZJmMDFMNt4NA0QSohSWpygPsgJwwaxhzW5zN
3CfrtJcErohz0c73ZxxA0oGjCz01i7bw2WmjV0CkeJU1Gx5VYWVUhygH96fqGKeS
Ic77KQuQepzUSKOC5Brac2dBdmvgOnZrpipgLMD03RulzadNLoPRZDoEdoYRGHdi
MyUp9C2M2BWmY9GjfVLbj+x6xj9MCVm15E0LUGCiHfNZX+zbNwREM7eCC8cJO1T3
1woGLBNy7+IUfl2ycbyWTqg/tipqTwLHR2xGST2fy9DhHENBzOoVG8Vg3j2/Qgcv
symaXzSbrzvXYa/LVMXeMOGtjIGxzIJui3nDHz/I9I2JW002b4CQLayC6Xv1Fn+i
BmZ3GfXu5G8hIHxuaeZikyYS+myq3UxNaLqh7Gn79pv/Jn8N7Sk71dvVWgKiN02Z
5W9sVtdo0irOPXqs4qAM9itUGjUXCemTyFg2nPRPYb9EKK1Oy+C1DXQhjIu9stHL
fG7qUtu6thrwwAFU/Chz4sx375JvE5jYFJWP1w+razB4NhxPQdz0aiQ8RUbjI/7f
/W9AAzfcbsQU9ypKy/6r4I0SBzGWjQLgdtNCXu1gduUaCq3qNDgwUbhkPL3XAMGe
M3w+q8rjM+XKhFrcM6Yz9L5c/lFxsFej2kPVufWYURkF+oh2sSchs9RQH/Xy9UlG
p7QbgROLd4Xcg3oD97mvTfdhvf0WI6m/rvX5scuIbF94AkS0jyOzILQxX5VNZ8zT
MkJTIz2E/29Dwj5WR1sohe8BtCgNQZpR0OLWVBokYSAnHRsUpZpvUAmqCwFUu89t
Q9MK4fBFM6LyAkLsEN0uiGTxsX0fEjOaU6i55yrSiaSkEwrFeG82R3dd8+minK+H
3jgg5aGIwbLOA6TZ425cYZEGuPIys1+T/x+6OGUqBHclt2q25C8kLliDuukZGQ0k
uB8WxCX1oXglKttrAN6srgBL7ulC2lPrH4d1yDzI5kSATCvMpNzJT8CKuMfyK+H+
QjH5cpRp/C0Jgku4/LugWknABRxmtVa8o6iYGpW2S9Svn/14BfRv4PNOd5NdO1YB
Hqyec3qROchaA259yXxnsT0liBJOBFRkdwTWmG+b+LFxYd5JK8h6LisBc4UGJI3w
KMLzi+vHLwjozDJkppNOnSsrZ+sqFBAefHI98ZEQxKgQFvGuo+60WmO1uZyXW3rq
MHDzL9rEhYYHYzpQEStcQ0GZzwHkkyiHGbFxO5sjpwiI2LBpjTYP6ncgBmjRqlls
H02+E0C7zYZ4IrLhQdqCMbo+BLVyOOotpEbX8yidx9Q8uPURe/tBV5AMO3Vpt2RN
TX/eDsVDCySsQRSqD9uQ2heWe8/xEb4vv0kDpO7d+Hycw3yJLx0GutWyMws5POwG
MWZghY97zWnOLdbddONuJsZmZclADdy47jdBQpZGcWeQc6LlKdFKDu4kNCFXMkMq
5JfaQ47dAyWjFsrujW1xkeEYV/pOlBLAZPt2hOrFBgShybliYJ9cocinAeij0GsB
mPErcPIVHPr+7NWFaUzXgS40Nq3RTlWQhgJDsVMhUi4sCT4IQqF76QIWGWx6Z4Ps
inXhvUfmi0kdVK/u8SrASyqeUHYBLHfWrrJbErIxdltNYvGr3sVavT32DR1//X34
HnI7BEYVpG/KKUBgzCn3Xaq7m48Mi6dT4HhWyiOPtEQhBta+AN8rWWJ78T8EET7o
rD9JvYFXEmKF4ZhrOoqcOmZ6AvUqZlfCSTBrLG2mk+rgWymEhSvxogSs5mOugRCA
5HnFYzcuthjHoFZZfummLC8GkaBXVvq7wvLSg81cg+s+SSP466tb566Oej/p56qJ
oF/H2hCngxWsmfXbW/8+EpTeETfy5+PMZYQZQdpLRFI5aYCfZ75Kn+AEK3ZrRSUz
86j3wZZYwmZqQ3dIXLgf4dEDGum0+1WWWnhemvHnd38iNtAOuHul7ORNOHQJCK6P
gQR3AK12UceV5aJLbWIxgTSRefvIoXXve0sBbzIDYrFdTzeEsCZSKb32rok46cUc
fbmpA+5kKbtCrRKdUUiYi62rjf1cHlX40tqih3GhBVjPAxG8Fyy0prOA2i6q2Iia
enUaleLYUGym2wu6YsQ6DnMfxA6m3k/Nt1Q59jtYhLwEMu7ONYNI6i6p2OJmN/n6
dEmDQS6F91QcQfB6AbXEEtlZ8a/Sp7I4hN5pO3l9fJSwXw1LstKG2HIwJTYbCiRk
jgiNTDSGkWd1AP435qEPQHZe/TcujldAHW0TGaYqo71vJIItLfrli+GCedg8ifr9
YGU1e0xIbKplhEyHKdCcXC9uu0in9kaR7ySq4zLbM5lXpV+WC9J0vIQjVsFygeUT
WM69FhGrvFnHt1B4W/o3mC662Hgn5kJMh/FIo//flCXBjCY8yXg/IbuufYMvaAor
qXkUMXDcH9OkjrlXAhqo5dXKYFsihfEXTh9Y1FlRKTXzH83keqRvjV31Lz6SFsB9
8r4zqBsbTJOy3Vaa/+vYAVogIv+QfFb09InOk0ob7sQpWTQmwDUCk2PrF+hjvZUw
z3jtx66pkqfrxGcsHROZJVaDKOVZzsiyJ55lh25Ifo57G2I6ZnzIAxo/LBfxRcC3
ChOvQaNjoMG5KzIergtx2k9BttAvTW7uKtOo9rHgqydUEu99FAXWtfuoIpFEx4oa
b8vnIQagc2yqXDudXqZu7ukqEeIz2Hsu3cVT6EGeYLh0Tl8m3MAsZMnxlEhfovLh
ZutRsT/kxbfo+OK8mvJ5boGAPA0mEvVNf6W0W+RON0F450JN+vw1whFS7ZRiplj2
d2EMSROkX6JJG6HT4bgFspXGdLYsJGo0DEGtO3ypT6iR8mKKVWKciUaJA1jB0+j+
VC/EBpYACbUggtk4ks/1R2Vzn5oIjVvv5KohhVXw/mh5NsExh+34Thlo4IOwU7Sw
aSkJBVLwIwgJ5YYPq38e6Vbi+ljpBYxM0I1y9tXAK4HnQdOSpZ9FXD8gYV+L5M7D
jBy7YX9xasOHkG5te5lvB6RISPefxtyv/j4rYK+R/05SM0X+hFXkSanPwjWeQ45a
KoodmhaTO8TolYETNvwF/OdU6RzoCtblo+gquaWy373XGpUP2uOPHLJa5vLaE+4q
LuKcnELwPcpNogg+QbowopEKiMLy2HZLQDHKRhKvSHpCwEB0aLCvNHtmkt1l+a6N
V34XNvAJQ89vrxfV5cbpmI9EL7kgQN6+ckoWhSE12NDk7Keh/7XbZ2gpXLKPtCRD
iqqp+QPU9GmBTU3EPAAUiPJkcU5qUO2xLV6jnXZ8DXwEiPlqyCjpOG1tBEm+Pg+U
K3EGgQm8yvmaDk05k6DeZQWqGC2Ps6qMgz4EvO4lwPCQBzgrvpjiWu/tCmU8+HKB
IjZgCUphSjeaynG1iSC9yzVHA/k+CzSqGgftrcXSn929usT7wmaGYcrJK8DcYBJ1
pfpAjYdFAiNkdzIXqbuehnOvwustrnVg2KjcdZQJTFSbvIzIUndn403P6ukFIHZi
Ibl8LfOEVsSNq3Yu+hg+UnN/O8ESDHw9ewH9GiRAQkdKcw7xe+fNe+5xGAI78gUu
BBj/c6GL1CsM9lMBsEgL3r6u54mJ1YqdxH3AkobDxizwZnWT/gUrk7vVwgrFFLlS
7lq31gjsn84onHFNhThJPpGXKUyk1e5SpgFWJYJkI8XYke0+ff8RP1mibEKDXYER
DMpCzpMrtvOPp1JoHzQcr/wDfqMpdM+CU1TeSYIbHQucvygY+jhC6wopMVv8WR0+
d2MXelSJ1RKJjJ+IP7NJq51npaKumJ3xqzZjJ6dTqeiHX4T2MJW/reYktNuhGrco
KMLbcCGzn7yCZj2aO4lZ0+1WFxn0Bccm+hJSPhpcvh9WU8A1d2B5mHqfTPvQR5A2
Y7bn/yZ6oXkai/5wOMTQRxV8Ocr+pa1U2blTPOtZdBdufgiMhrD3jWdHuG9Y1Ymh
X2VTyvyGcFI7jjW5hWsb2wDbuIQ1CUAeDuQWRMa3WKFcDei9J2kI/MEJV/Rq+4Zy
6pPTO3PPvdQJZ6Gf7eQY7pC2+TA4I0yNQ7mM0tIHQwQ+5bGHnQCtBRReW6WfKu+G
DAueoZuudV31Iu1IvH5bGcy0ZvQFfCErHfeAtA8/9+Zx2TlfCW9SKA/RMYnn7tWm
rC9fZ0uQbw5Vv4uCQy1pkshUghZB246oNzXxKJnWz1LFRe/bkdKO01uc6KVWrCwB
gDMa5llxVZBqimiieF7XJa94SWClbq6d9CtAnQs61vRcpVEFcWgyqFHM1LaB/roU
xh94SuW7quEkBb4LMA7R1EKs6E+HgaJffvk/rSOnfsM0W9GW+GG1Zz7TQTEJF7PE
4/7ur43dxlf85MoVYhexrKpaF1MVqtVhR8q2WnBXiIiAQfk7M0VtkvijiET+9W1I
ARfF2nYjqWpInBi2mt+uIXA1+6aLxdpcYgRChSbFrXtkj1hT0LhKDFed+M6HECre
6AidnoZPwWzegJ2trGW0qDeinmJsqzUc6nbbRkNZmVBg47PEmVdKkOnTkedm5uhU
eg0qdt0Hwh6ToNig2nw7SyrwcEhsBVzUvvwv08RfiDU0z2msGpdq00N6kN+HkQIg
mhL1PihLe1pfiIbYJmxEvtCxwjCQNsBOm2nRyJ7n5BXfeHcg0o+s3Km2VKMSQQjP
I9TERJ62qOndKfmKSIMg0RDm/AvIOyX1tp61ckMoXVTYG6+mdwB9L/g6vCrIZgF4
vlf3LvqH/lQWKscCXrAnaSTlgZTFKGohw4huGyOR8Hso83v/wazwjt2O9flGutHb
/Qs8ZilwohMrEUmKSbKgOoeDiGvOFsni51E46jQF1HkTBJ/5cnvPbO/oBkC1Pa9h
pnyZv8QMXAU+/8I4pflPj7pizo2rjmqjw6kYnB6JLh23HlVjv1m6deuvgxGmLcj6
GAnjwkRXxxfMA/qatd545jAjEDHQ/2qfRzTVU4HCZSlRvJH1/W2wth30IbTevrn4
LCG1sOCV1AFdqdHkPEk4+Ln4NG4GwWx2GLvFRVLbOmMPWBJFX6Vy2hvnRfEtH2x4
1giceU2Khr0CQ4ZKidbw6Z4HVQ77IoBVL8eF6/GwKYmFsDHGEvZwgwSiOpzpbkoq
L1LbO7slBUkfrNjdMY2H/Zei6up1MpNQeDOHD+I6Q7xmNQvdB4oT4YONO6L4q2jj
NtKqSy7oqf09aoZreA1kuIF4SxXab37HQXgdjq+gGCENRdeTR3p2/dyDH9oCa3Ul
Tz0+WtUoj0nDKHGiz7r1WOucmdeB+eNFTERRk+ollgyZc5p5UfvOkG0C+y9ZH4Tv
QMQsbJfhBxonIJBpYQD2NRlctMPeP6fc3yTMOM3l6iByzdoafbDRDDjszvG31IBA
X8wo+pA0Y5PVwYKD4m/LkLWdC+HhXhzBwjK3Qk+RTfOCAdYEkaybhBHmqJAR5vtq
DaNY0aNyTKHWWDsPtlrquE8COGKmXAgrVBx03dPO+yk1ssQo2Ay7X0xu8Dskqd3X
nwZIyRTG3i9/rvqimrqhfNz9oRx+ot9leqRE0pRLk9QCyWG3EfI5pf9DXS2v8kCH
XXCOAY1AkBZxKFcWs4WI6Mn1V1ND+yh10Wt+lO2Xh+y3O3N+5J8Cwy6Y3886gNk5
e6QRkIBbkqtqqQ99p3y6wLRHjNDRgSsvH+7xUHOtyHUQN/NX22/9yE7ABnTG9fHA
zXZL4rVvwWfGt0LU3oW+qOsB/+lh+4eBavlnXj0l8NKcashXWz1vEPXZSWypTF/R
/5xglAUkaZZbDv1bwd+we+pEDV05QpbJ4feYLg4YiGhGp/9tPrMBBm18ZqvR1GVa
Y1EPE679NphLU4XrSjDRud9unsf35qQKhi0jveFN8a+TqKln2f2w+NOy+WGm+DBR
4HT3K2bLQ7BV/Uv2c9+o99bvN+ncnYkZnYlTH0tmcrAZRxV3VxlSSjnBw4EY/KHF
T0rXT0435GBTWq8IBrM3Rz160ThcwItt9U3LEVqsXXGk+lmEtDfNagM6ZPiZnboR
rbWVS6E0QNjHQOSyxMua6oP5bBD2HIE/tCpWEDNHP1KTVuswIOxSjIz+eqj3uPFs
DpKZbMieVXix3DB+Ql7tXpwoFx0mCKt6LhmGa7c5VqOV25GToafXaaS/AmeT1Pls
c6HgppsFJAOsCwwTMV2Mj9XHqMRk4uuOLPVLI8KGH3/GfrTBAtQ1II0WqJpvDfBp
vyCI9yI1KrKU454lCpvq8tCBWQ3P7RpDEuIL+9CDZ5FQuy1mm3I61H+DMQp/trhK
k011+pONns7BSvErEm3Ak8ickJfMp/Sj4MAZi3diaKxf2qpuchNdCrFypdzP9/4H
QNby2C9dgPAQDpg7qodZsv/QVvrRbgI5r6XCxkx94BIRgkP1QWkaRt0P85Htzz4/
wk9arZ9+KLIz12eJD0LAxPJBll3/WYaYYDCTQy6v/5mtsyl6701NWL7e77JZDxmf
vKz1v1negHHbBH6UbGLnGumSvYZLT+iPSrAn8ugnEke/9nmmTmWW+QBErASFetCa
DnFPK6XIS0m7wajeCRuGjhKEVi8x8UAi6YwFolVNTmWWm8Vquugr61x0Hr6gfcB5
QBsosFnVYtrN/9Sp+0uvN2x0PlJlfWMhlIsFZFDEqGEsKla3j/1mQDKjmH6HEteg
Ell7mTfVTlszF/LMSCGlPClWCeBT8yepOuY9IVVvZp+gZghaIkrlWlkvtRhjGrqL
BIRo/rKcnfaFEONhqon/61lRAIqKL7IH+i/Q0IneU+r/exDQSAxYBcYmndKtfYT/
y2/vecH4aDUWP9SgSdL5xBBwfeI6MmOd4NlENctJ+b+hKwCyN676reYV2jkCOCUJ
1IlsRz+2AMjAtOoq08k1wVAWzffxyGPJUQsCCaAvq2QCoC6ZhY9yHi/7udC/AKqV
ZZoq813nr0t/Z2tauszgfBaCHgCsMfQxSYcZ5uV3rZpQ/hoIGzQcrOGiWWrjqLBf
rW9d8y/NYAhqVKebkNE3KiWLoWx2quY0FswJ22+z7F86CFyTDe6ZUhvJnePlvYm/
vk8oIPulf+mIlk3eLMYSFbjkX1bESFOv6nMeMmTGY/gqvM6CTf/R0P+wC7GQ4013
8LNJV0u6wERFNmCaQpZ4McdIEMRmvn9bioSbuq5AoU/FAP08g88CobVmEUU5qPry
ZGFa0hYJJdYN/ASNLL+uZgo9P6gOwl1w4c8WOTOf4bLYmWJTHl3SplbsFFr31l3r
2YTlmRnGxZvgoLvm8w2FxIe2s2Xt0BMekBKQ/8BVB2loSIyYzt9KOMJky8zikACJ
xxaiSPQa1AtT6SqPkmRmsMjQwPUqLDFsFLJrMNRzrLuVehHxbEaWqdDUZcv/qyNG
U8iM9hwr3XfpGAjwhVmTmkeeiUd3It7ECMdvnqpTaQWXODrKSEfX71aDx3UkiQKi
MLCDyvE8vMZCfGyBaa6y1/nKkPSBnaM5UNr7kY3T9/On5lNmz5vmiik5zn7RNB7x
gRPM43o8+DFLBPUzULbLsazt51TplvCyV3PzmewRNCVvZ3VWFZhOhYecy2s7tBSM
au3VZ77v8g2/3gokY8N0nzlf9wO1puEjmxF2/AvZsRQUp9X8uxWWUSzVflX9V0ta
eUmusEkGWdCVJ/K66nCYXVrgtaWpMGmZV1DelO9Z1z1lcAaTRk2OMWckZYlGrawi
1kLjB81S4wkkrD6e76DhLe42XAjA7IhZpico3+S59HwvnmJ078ipOKkuOVccsYPF
seaYaKo7mhabYS1fLTELP7ObP8zfhwDFT5WTdcE4kEgFedmTlHKObEJPMyhw2frt
XgXTdLzHawrLlsX63NFHSkNrqtblCtvYWwrQz8unc64JXyAeVXEZVhhGBGfOg8Uj
mgV/3uLN0VkTCKeP6oMeRzx2Yu7KLg931Y77/UWiTnlE+thKCWKcYwOiJmgc/9kq
E1EN1aDp5WuafGnkp2/8CsZZSx9tcEpGnkm4Kv1u5HDfMYfMtgRWq5rgIVeMl+0X
RZFz9MkzdSkvtzdfjZq8uiDTdV+77wXy8hn5rBQdQvK4XM3lDZORDQOpmA9JZBui
xrBHuUAhR/l/LragSDSFIOXTfzSunMAhF8S7ykPW0GofHrY3GO17fxGJNf0XJ1gy
2jCfdJvJvtLP1F4br8h2qvjGN7zNkMh7GUcDbocKjcL/q0lFEbwirtgQX5RXyoFq
v6ho0+Kitar9ZFe3ZNLktKnQJdqtpATR0iE5z53TZUBZxUXF+njt9cpwcve3j/SE
lv0xwQDyumqD5EIW903PWyg8UZpeVTWlbVGNxmS7ator+QVbM0kU9zEaMEel5en0
Kh3MjgyHTE+qImd8OMGGwioUYg53k2XJ2NmzxOClWuAdpS9dNGPgp1dyJ7JxZRNE
ZgIAhgOZhxhf8W3jx5ceKbCQ1B+0xL4xYuKFeLfsr7ih3Ni+1T6mistyl6XISKbd
hAhd8APkaS85Go+DsrQMVCVehJkwDNOai0MkScDVtuUzT0McNaL8/X1zBVZB1n7m
qky3+jIf1V7QaqH7LdozEwygAglaLjkuF7d4TzjmH9/YX0Jq3eJ5mHpYnfpH2QBd
T9kVTr2IWP/JncQJg6H6YLMRB4S/zRBXWXEs3zibxhyTeK5TZJDqFMHM/qNdAR0P
2vn651eeM3wNEiA6q4XIXPVmefAcu/pn4AuBJvW/9Rrm7Bxs9y+UWqz/aXE4kugu
PLR6GSif7rpEkTBEi6XRqK63vPBVZxqepzvQd1nZKsFOaMhbpEBrqa2OJPSN3PRE
F6hDMdvPG7vEiaC31hhj5OXpm6Rg7+NfrrVmOY0mrOATmlR+d1wpUSNu7K6GcaYJ
dgxdL07vKaDe2Q4Bq+CtDehDlxCLMT8E39EztMjqHvGBZRNq+GSRWZQJxiBmvFE7
xJnVMX0+K00aeSOUW9RGzoiqDZ1ZepsNxL2Zp2NfzPa+d8gvte1bMxAbRqlp8qtx
qivgUjTjfoLk8IwWtWwICqU4bGNn+hx6v45osWwH+itWYNn7bTpkZv/NTTxZPUFd
8C9qb8PSuc786Roo64TSQt5tBA5ju8YrD3TTbngB+CxCJh3zJhRYDwigErf1S7A+
TpIU0K0mSlxrnJH3NEQXfIqRMjBzj1UX8X3G58tDI+zknxBHwNJZcjfiOJCYfP3F
ZdSPF8dHSRfx2+NxtbCmQL3O48jfmvpVh9h2k47iGO9BPQpD+67Z6thmjogYLGyQ
xBBqBX5OT2mEkGVrvfiUkrL7n4DCAbmV+ob2QYFqKzTIJx0uwcRGtYbo2Cr/OFuv
OnsN+G7d/sq61uR2x16xUZlCHEWkk+hAfrGD1Et6RFiHc/3MoecmY2LNGB3qfzwq
h2J02NhlRmNW9fAla/u/vZxmNzniV7gSsmpuWOccLfToJzBqAUw3JXAeq/rI5Run
gJgykPhzPGawslunVgNb6nPpEgSAPTFGZwecL4MoOgLsAVJGoW1AfW/mO8TZLs5f
PX2CoLU6MeLchHYnr075D8q4GrXOF0B2/3TCOXCn3glSDCvYY383vbVlc+HY7auj
hQV1ACJ6Tp9PLG7/LA81GSmSI1GKAA2+pXW7XdDt99k0g5e8D2Qx1+uqUhSqsQBk
rihSyNZnEh1B/Fv7YvIV4lpN6aLUMK2CiUQ3BgvFxRAhtrWQq3jzczU7B3yr3Hl7
TrnHX79211m1b0Lf6Ek9qr8FS49G3bQ5yiOVeWRArQOrrcU0rKr+r3WLocH+zoMR
G07Ww1Ep8BikyQ42EAuYrCkV6FfEN0ZR7Nq9p+VfLJf9T83gqBMYpD5G5/WC/W5S
v5SKdHlndC3S11J9W1vLWfYvliAcMinj5Hm/z9tYJcwFHR05owBnyWdOvG+T3ElJ
fyofDKnNwW3uugWkg6ZMIMrdJzeuFVaEZc83+wCaM8HjvMWz0F3vXVOoEUswklC0
k/LOw1tTwfp21sQrwXVSlvH+scw3vPxp6i5dGOfE6hwwwYsLw8T+GOYVCM+jHOVE
0Kr6d+1j1TqZiKeOjLWOzyOzROyD2GgqPkyjCcaYTHURZ2v853us3C5yxqk+aso6
BN8ZdDZBZFNDyXAWB7q1l9Ydp48bCzPdaxUWB4k2RLRYNlxvklDWylugf1B6wHtK
NZBfJ4R4TVlrf9XncDkuoqlraCxK/fC0U8kEQ2J3GevfuipU95DJBTNsx9fILtJJ
V2D80pFb3NjH0sn/blJQCkOhd5JOwBAIqZGNzt7ya/bmUYHejZFIJD6rjAC9K4R4
3k+NURZTm3LD2hHT7wTIRg+Q9vT8RdKny/vidVTG/Fp2v3vnc+0WzC8QA/IV5a1b
/1g68/AtR8w2i0/cALHvqhPrrlGDkjRnR0WRmsD+Q2fWbRGD5YBKZ7b+ZaxXQAVl
GOp5JbcXbQxqcfTqIII1BiJK8X6azugDmaTlRq+nhnJ5Of4T5h9qG9GoNfUdy1LM
Oo+oP01ijx30dJto30rENscPLifhltCq6XQ1Zg5ZIHvWlG9QfNqE1y3PUnPOer00
MGb0YPXksOhD/Gy6tnAwtjbkHPSarCHab826WUDLJx+sN9XOJxmPZ9oNutV54Bdj
ci6OIudRaxK4HadhFiyURxVTDEUpJUx2GfQjhrvtYYcupWW750J7oCABLQFpZZwg
TU20LNKtfUgQRXBUTutrY5cuaz3LL+QyP92NJb8vvUlS6VUC07H/z5ure9DsXdyb
wDDrU19f9pzTz1flm356nm/GzZoySHcyffh8tdg91wgWbhhfhc3+y96/FRZ2Q2vD
1+fP/d9KsDvytmj5zR+XfYbWQiSsa2C1iPIav7FXrt/k0BTkSipTFkukcC9r4uS3
9HKtKkj7LMkdUaUl0MRANHpAbV2sakt2K1giJsAmeGuB7fVznLLmqDw8uPSfEsiV
0vNudn95JUsOCIkB+ZQfj6HZ5zu8jtMBPqZTFJmLYkd4gnUGr/Fiq9IDaMvDPyo0
PmTHhPjIyobEIidE0TKUmjVxgY7m4JJguWxJytDGOf25wktB2XGTU+a9D0E51el6
O1raGFOIGWDaPgIkkTBuIQVdyRlqrQTQ+qYgEJ/R68No/W+1sUEPJNyJCwT2Fa29
bu/zLmnWvVCPN3jmzeP2CCa36wesndMuTqehtiPknJ+R9Wen0Ta3ij2lDhamXz5N
zZrgd6msMKOKC/DlfzRl8iLrn8ylGJckR3kye1j2iCwF9tHJ/99vi4iDWMhEZWgr
H0LhpmVz49fJ/fJ4v6ewr5pyX7x28lG0NZ6mm0Th4WWuZooS7lx6uF3wxa+dapyL
tvuBQx7wLmBOlp/DN/gl+LlPtc9NAj9OeM5AcKMJCUjuJ2sXGh+bbs6XmvwLJ9cU
bLel/qAWuHp6odi9uK13AIVEK3QdK+D922B5wGxlpRvA/f+0FgCmTCxNLiAz9bB8
yDnVFX1x+43icfSqx36LLzjoY3OkMUvXUSxb8vOyWzh22Bc/HRF7hfbpq945ZLxm
ytP1gPZeJB1TB5sSm4yJMYzm6u6yit+/R988w+eCuuuyphKEjffazfwjAm4c3cwH
fdqGZhHqSLUmRhFvng3bA9Tx1L2pohWj5lsI/nqVw4/xEQmX1LZ62Nh8i2ih/JCw
gIBPZ7ynAVvSI0ziskMQGtyMgMApbIRFAyYXJAzTh5cuK7sVA9Z/7MTJf43Bus2o
ao/pgT1mFk0k7sY4eK40w2qyBwYjlL/KXdzeZ9eyjuJtt8isAmFo+tgQIfHFE7Xl
RotzasxmliTqj6C0zVABC3iBJjk3tEao2cvllfN0PCJVPXKMq220hrSdfsKdofrK
E7dsAxK3YIk4HLojFtSNWzPgZAPI3Zuu10hJycRfSiDAuagdncF2SvmF7fCJ4xvn
AGuYSg5yXBc8FGS/qdh1MsBnL6rmOs9UZNnGxON1TgTJ8lQ8PJmRvtiOAXXIZ0Mk
2oVlZ/1AxxAGSQNhJU+ITeXlUvQMFIvhqt6F0vhiALlDvrrdvmw2oczNx9kwvzSF
7gWLXl8yC2giNtxAhbLRJ7AhQ4ajOeBIfXv5bYfNV842tBPtsm25OnC/EjIYe2FN
dT4+fAOKoXyOyV+TwD4LjiAf/4YEViM1rP8fZ9kY2sCEfduVscxvvqk5KNfVDbUn
nLb2Xs2tI0SiULeZikbCeyDXDRUeHyvBZHJUuiQvL4iojAIk/c7SGjH2KcbSqddb
y0Lx1TECJGw+uRqeddDn84z7Q+nPnzHQuWcXFL3ntcI5M5/YmEvvWH4FEAQ3m6jv
fu2zuoIcJMIXIGNQZFJDA2my4eYmNPxkA4i708U0+K1RjAr3tkbN41tFSu97ss8R
ohGj7j+GluMWZqBZACVtEt/AwGiTFezaYMOCROPXLXNC4VfveYEIK6F2D2Mhm/h8
ZJ5jcPAcuzn3aKV2uJ411vYyDNKixDASJ7eZPsnqigxq3CBCYzmoyOzzubjeIG3i
4Sa+BktsIqQNXR0Aw2kNLqDEvLLWZZUqlbfDXsn7rkS4UwCyk8/jj3cP7DXdYN4y
LKHajNr9byzPis9wlj2uce9Z61NXygCZ99fqUgA07JTb3ksOFJRhVprcAKHoaVa0
9O/zp0ry3I6pNrdRSOKMs0hkTfvDmugzpmH6B4ibAjMlmpmYvclRRXeEaJFGFxN8
v2htQ7B0bLVqco4prBD/yDo2kPgCIZjxnFad9W3OWyvt+jenJBWyu+SDxjsL6bfB
eGNoFIeBZlbMFVvAAAW4NGlyqmkjtsUlV7aYGKlakY3E/5QQxv0YRWrGQ3nNgbm0
muPwXFkVwECdQ7ApHpzXSBGtD4+bi2drWssdHfUmOGoet0Ah+dNMBm7VUZvTDtHk
pvESwEEValzdVkwFC0DRGpIr98dfac67mBJdTwodOrPg/3yCHJJCt2WZ/efb78ZK
ufaEO6y3SDrhT5OaonjL/x4uuibMoW5j6ChqVxBSMcgqUkOkJCxC/3LgJ3PejX31
9nXXeVW9ZVqXMaSC/G6oK1lJ1rPjOt45VbYMJCYSG5J4k0vy8+t6vADLXK7xXVL8
5Usfr+J1rc0MIbRa+uA8KBbpFJmYmA55qILw+hWtp2XoxddT9i/guBRlfpYqrJ7p
QLPXcotHyqtzLhekYHOiE2qKXPD+zTFZipzs1ZvlVkGo5fgk4mD87hDmH24lPMpG
iUZccqMP9FrWb3vZIWPhC+lZ+qXJTbZnlqkOBB5yfEmwqFkbGNCYiwmZSBo3US9b
D9Eo1e9Bky8n7nId3W9CoznETheH3HhxwJUsAVODvc/F9KvrK6BgQT81klJmwvGT
NQmd+1NfyxNdXf/8ub6tfzHeA41ciVUOPyKwoT9y81SvSsufZE4cKxx9tOrWgFqt
79SYHCKPzlSa2l9MfpT+nBqmg744f9jVrn8xK1+sHmq/ND0b/ZCXk3Sycj//rqwM
m5pcC+Wf1KhOpPsKP4xCz1VQdHHPek4Bsly0cqx8MOtvRqBCM9Le3R0jDBAz+7m4
7tzOvr92Y+Ldonuf6PEmhJ38GHiw7nYWcCsgML07H09NlfvDFUcYmYF0jhnE2Jxd
RmC0T1Ty7st46Yhe9WZFcOcU766twa6DDqxIaDPwHF6QrhmHpc33paJxuhbsa9QE
rXyA2qX8VtrgMhSgXHuvDTHkLGRE2vBZgd7jKSgg4tAOBMiZjec19lB0cu5KuPEn
QpTgnPT3FgKrAaHzBg8f78mDdbGWh4Cx2koyMjO3lcrjPuxAcENwKyLyp5DVArzQ
M1W1M3NgqAqO6KDcpYyquJJY2R9Rm77hYCa93iZpYhJP+RCLbn5uEVBuLRw09wlg
T18aC02RhvpKXZml5KBF+26wbyOXUb39bOYwLhfbcugbQPOSHF1FHs2jQgrPxPWY
e9lxs3IZzql6q6jZzzF5viBYcL+wrNVCg0VtOr6gwySuDVsDYGddbSLjwV3tIruJ
3YvSkIirvsD9djCNN8X9UIV2oACMMZToBjr4/yVoiKOtqtnoB4CzkHh94b9ZUWI1
jK8Z6JnkxU7AMAXa5dWaOw2oDaHpICkwj77PNiOz0LUzLXuSfd5UWZbpTTGj1rhF
+devX8ni6CK25BhWN3PJM9MWlBFy4BVpr9Ll8KI06crmKAh02S85Npg4R3lbM7XZ
jagdJvZpeCE9Fc1a8ieSfoLAdZfCTo/KpIemVtHg/OQ8FgAUKRQPuCPbv0tVYAec
QTvcEOH/z09fDDHb+xIaoMHayP2nclVf9zNqmTcf4vq78t65wkUWSgMMh1nCJJfW
jkrk82JAmBrTQfBzqnsirCJtXnrnBp0sgjPcNDvALgmHCk46J1ESCEatJifB54KT
HkL2eibHDXenPGsTy6SXih+42M8+OPGcD35l3kJJbSxZq9opW5P3gqDRxYvZ7lYE
M1Fz5BUEiwY0ccq8Cjx/Y8tJJpFcVqYqW8m+o6PTg6VgQ1AbJihQTwVwz9jSNy8x
VlStZ/h1u4DesOxI9oRl0UXTu4xs2s39pOIQYeNiwb9YfGmp7nxlaEAbsBB9Gap9
lB6flaDB2njMDSLDnPuyfqNahJq0vcTZJCU06uG6S2k6oowLnYKasi18UM83xpP3
zAFDMum5SKcvBwEcmVmUo2fYMpeOsjZZky7+GO7J9DCzekpzu0PboZphlW+iMpqy
JD2+/WeXH3vGMjeS04aYh9DvGn8QJK5DYP1s7R0bxMJmi8lQE/ip7rE2oBQRhPiI
mUUYUu1SBnZCHtvL9asqG76eNsVfn+xV40GJXMTJoht/Eh0qEb5znqnuA2JaYrEM
U2Ku0Vejwbd6xZKP/BYte1kz+Kwhgix7mvWUKy3pnGZ0FH3d3goPECxqpB3fdnTJ
2TQGb0Y9tZ/ZCOffeZdKyBFpvm3iFCQPUCSYONI2sBmKZzNEApB6TNm+TQD0mx6F
wECy9aFnfFRXF4c2XUgX66ndcNryOJunNaGDSha8XFVmQ34SezWQanrL+EHNYdVt
r8T9WGIleNLFP4iS08D+fSqbhnWeLTtUBQ2RsqcRMJZixjfLwO46VaBomVuDJRUV
xWVHjHc/Lb72cQAckI2232WkyV4zKPQGkZuH6heF4QPT4PSDPU2wKY3RApjDBJJ3
3JTdnoz4g4XaeYwEb4mmdLjtwYMuAVW1f+PGhiKceXRVKTHBZ500AT96BxaEE1uX
dPwWstpyeZnltz/RrAH+TcSDUQGHmJ04zbsPVmrl8DoCsO5CPK1KYhLKyCwUH9Xk
hDqFQJeRtmpoR3WQQUuiFzmBRsWSjTV7U/vT4wH82SUqbCqTKdG9DXPtzLvHrKJP
f5VZPJY9mGvGfbwPQwVYobd1bf/tpGBe0Ggdqp0qvi5xxPnUw21ZYqkfCBoBT8mh
mqZixsDtLrwxgwawAOsYqnk235vcof8KiAgpjtVVQ+OsAsefI5NQr2+JHP3c5aYr
G4EoktzuXuqmuHDPw8Z/q/KENDfHvs2cU3ARtHo4wsl+m0d6ggbPuHTCDt6oeBs4
UMGSBJzHjOWRpPgG4i96/MFFkMGfJJo0f3af3Mv1/J9j+BCn7AYr7cY2QqTQtFCx
G6NNFuUHxgvFKhFfdKx3CyEcL9UfGVCKQis9u9MBYfDxVntDBrcxxtcKtnuh1ea7
ZGuHXaqw3upAh+li1ek6Vu2jNfetFocdOuVl0O0D0n+LThJ3xD37zaSmUyvEH9O3
zz5fgVpWvlTnlZhRoNWu6Nr3U6suoOwfHd5Yw1qe9rzGeHIvSRGspDJKth4EL7JS
SmMMpbM5WBEHXZQ3jvg7Z98HGrEEIWd1PvnHqOYyMBEhFp6cNz/m6pQe3xf69IZP
t9NYJPLioGQX4yjBhJZPr45ES7vKGA2Xz4Y1bOvYaykWWUsaFX6jU2iHxCjaRtU4
KJtHGzpCKX7HdqT/ITbVLkOu6Nd4N6rH9xkFQKTyD49cQSIP5zcwQ59Q/dhT3zi3
iead9/nn+Frs4MHp66oH2JdN26j3iik5xi6U/YZkZPoaKLSsitvGwxfWxHOT27t2
9SYNuHIQGaYnWD69HkwCfNav983LsCsw5PXRHnvjdwnOTMhDeo7LY0eZbJBuSfeu
/bcecKEbwrZ/FihqijuZDh5a/LZPCkIFsIX9Iz7GGeOQk9dd/pd7Guo9cBXQRFpM
/zMQWLZl9x+Z4e7Nrc6L3XFOWPCpNpKEfdg98OCPYHrykBuzyXPSBixnnWlP3qck
Wfd3/aut7oL3DGnQquDDsLg00YNVq1r3k3XLOSzgUFfhvhv+VdnbDW8xDQxyuL+K
sqgIrnhFhOb0xi3+rC6j52nDzk3j2j9qmC+6p3o6i6GY6um/oXfOcijY47kRt9hh
HjF/jPnPFXda3s5BbEhatBvRqI+0mRpvypnMCfrp12sEAXY4rxZitdo05X24Mk6Y
zV3PrIDG8ppJ64mJqNtEFdcQB+bECkEDvhfiKLKe7DkkJOb7Pyj96hj8j6uatp04
CdZzrKZozzB60oWqAIGZhLdOQ19fh/95IIqCcKSVjEdtO4/mnbm1j4BM/XxYA+Vr
/KcX04zaEtRhGpOx+qWLmHlGCjdA5ApSST4d/ZKhadQo2XxtpO7i7JEtjSMUJJ0B
eF0Z8/Umk5P9m3qyPeRO1KXs/ooIJqVRuUtZvTs7hGRkYgQGU0MgNc/d+ZvtYP2j
lRruyAVtLG9i8ohDbMNqRrYHRP8Ta+hY+lbuphcdUZBDBRtx11iX/c/NOCVXaTvX
YCNKGJR3RdfGAEdIsE0vYmtv3BZfWraja79fWjdvwZ0pIbhBoQs++M5TDMlHaPHq
/mn1IxV1nJxoWMBdl9J+TCfauRvtmXj1Ev7ChTHKc7alTCTue0JJfB12ZQAdkfbu
CfYPT5mhGn8toGzt/kw8n9uI8ikxZgy8YyE+RryIdacFsPZIcNZ5gsm1abegB/zT
2jb7IdlOqb1sQhlr0ELiponsG0iKUR438Ubg9tY6K+9AnXkcNRfceOn/Vuq+rLCT
pSU36Y+OgaGceRgx1q2lW26QGylpztrJfUyq9cvbpu0sVVhWWFdf+kyuh4MpuD3N
Igeuu3MidWjZSfLTjZ+bPtcWzVuf3AVHag8I7b/UsOIpw8cEx8vj2eQLsfdRK32E
NosQ1qMlWaC8ZwxQvK9q3GpJp4hmS4qVs0zRzY0mXmNvq72vDyJUoZBGVC1qBk1P
UioIqOX9VQxbfRnafDDyv19Y3qSIh609TTo9NerrnPgzaFbW/lsF9iNmftrIhkoy
puZg2g6SAw3HFoRnsB+ZXIGY+YkQbwWe4ic/S0Ddi4ezfGUsp3A9N3R+Qy+gWD8o
q59yrANZa3xOrfWzHTkatHyU1OQHXyfgQNVp1vvvKeIt4iaKior01UCGW5p3ckd4
6usT1P5Ojyp+aHrVgNPZpo5eqsCkPxHgn2WCmyLPQzC9vVIMiGS07ae3FrIXhNzr
O+QUbDEx44qZix5usFV1wT5xdzfQTPVNFtsgEuxIm70LmhbqBwaX+K0xbVZp4mN7
MKNAzBd9IKJJs+252oX0jYwSoEy2XMbKLT/gcqJn0R905RMAnJVWl7aw/qirsm4B
ZlpzAOj2zai+VfWvd3bsvPVEQOK0yntmT7zQjZuabKJuHfaCoaihYDrvjvR0GyiF
lgEToZ9dZnIYouf5Nsrs60TyRabFZX7pfe5RnmH6hfm9LLOvXXzU0ejPJIOj8Drj
IxbJYP9M1BZ4z3vlloGcWpzbRqABjzm6tKibTruo8Ns4nVDbZEf75ABqHZTzocwc
rIgpkqyf6MJHNo+gnDRf8PqSOtLI0W2ya/4RPrLQ57BJRp7Ej6uW2ykYXsRg1OY9
j+b/XimiP58BQf1NJEosdj2ydibmWPDEbLF8o7sM0S3s2YCbyuIlxjb93qden9K4
sTa5LVbgiRc2vZA/6TlEFBd85StrvHXGtP8oph7jhkdXK/HIGfiz3KeZgfVe+oJz
8dM9DLRB4TlUt/Y13bZen8zWpzF5d/N5G3xJrsEuaLQTyRcHhrpdOYYF54XB64vm
hpsp8Tx1ftcNwFLQ+cI6nUT5GGtnGSROJ5A77K5PssbeNyc8u54ubJlaCytXEcS3
5C29QsNl1GSHaCh8EfQ67dHAgQ9WqdAW7AwFFVyO7B5jLaQu1Q9oIkpmxWktxh1P
So55mkSB9xNZuiX8dvr3ms115aSZBmbC0u6iIvp1X3GgPiuVE1OGXvGDwu2iIALH
aOOo/p2h53myICVQgwkR/hsoPUcvN6NqrECyfC9+FYu8MOgSOzZtPc+uN9+DAq5f
Qsd0QCjpGsHKk2Fx4HWC7R94yK3KSMPYG0vVQCE56IJva4gnaEGGAPPNRVUYIV6X
VDFz+LpA1da7Tg+/31cmr+I0yJYZY+6TLb7ZSY7bepre71+y35if6Z9WnEnN5mvv
4R4xVUCmDYsEEcTpwiTE3Olf60fm7QD8+Oq2zgbtAbyTTgoSimVZgrMw7cte4Z2w
FLmNVtAhmOWsrDFrwS3C8LwgIONHc6kipgIatSvPA/TmEe3jFjGJrx3emieYc7TG
Sy14gJEuRbU5BNuGO/VZ0MKfEtV8rtTWhtPZ0g1Sn3t1neh0dkTJqhRfb2QQRgWX
OcUA+/JiWcOvpxQKPOo0LVsgWjHwgXniZJYPhf1JAX1bVJIOgVqiRcTjTzDV1QNR
gfDCBOzQZ1HhmWr51DP5cD66bwKar+ajolUfGB4p6GL4YBtd8fejQxWjYMWEPew6
kmrfBHrkO53XnHnK8DelUvepYQumqyDdu/VMzFeQLc6AZvCeGA/w8hw8x+Lu9mF4
dVlvt0Q51J6Dj5lJ2Q7vAdwUYB9/to+G8JjtYk9uCm/XWemp+Ig7qxbzrm3ZQHYB
3lxL8g8V3wdX52tu9dpVBGPU/Fy9QqMluMQMVim3KlEsHvtpoR61fU1WvZF3U3m2
J2t1oYVgJlXnhyHgDwfUneyCo7/HyznCKZ7kesGaG58JvqEMVBiAAFBPPAv3mm3N
emU8oAkhLcPC22GUhdBVbD6uVXSAeS9MRSx3YdzEZUhdB+u3CbBpMctVgdbwAHsZ
I1ZzcLDfDKDx4WaaBg7Daat30QQy8KD3/GDhf9zG4jLeR+JWIhC01bhvkLUJPkfz
DX7XcME9LHVCN7ssrmCPRnJQyIaxgqOs/VrhDw8vlK7bbjUytT5rfWJ8svYcxNeE
lNHuD3Ia1C60gRJu1fluaFlIZBlBYnwdyvwyweR7YcVZkeXVXfg/D8/+3J/qua9X
f+4bfG1XkG/cb+2mSw4b2bkSYNCYKLNraLdVQEv2+87Fh3znaHVfI+e9Ens5V2C/
ylnaWp2eismQNprQHKtxuG9qYA5R1H1ZiAMw3ipCy+w+j0kAqZ5h4Zm3HHT+ZiFb
ZAcJ7l2oIxBq2hKpcE8jbPNBFKJWxF5NDWurHjLTOlsOeLMiUnslfY1pgytD9C12
cjZ6Bw1AGNGExc28N1Q6irOPJxEcgY4OVjG/1YrkAEFKnnUFX+pDEee8z6praCLF
FAUMTinfESOx5eFBq/UtdNZQDz2Ql2ijoBKEeTdf5dAZxZ1chIoeY9Q69IyG0TDk
3Hj/XK3rbJGPWXUuwqXORAod7mbck8EeOJ4Rd/hEOoXTtRlY2TuadNnDFjl2P9en
2uA31PG+n+RfQ5E/b9r70xa5UUgKHrNNkEvlXxS6Cm+tfbYnwOh2rgXPc4H9XxxU
23egrxdFeXKRyfIGd2NNgEUkQaVxK2j4ks3aUXg0IwnEJFIovm+uXMtUMVUMRrJJ
2yhIW6gFdUgL8ZiiBfw0kgGu+RqE5j0MS2Y8gpaUbNRGU0a0N4zHKnBcytVo2qdz
nOyEwSqu0wCUuXplCftlFF3np9xSQAawhTtgKt90EWkd41zHZgy0Jd2ig6x/ReoI
Qpwf681lkV2ifYYX+pNjsC5Iwp9XivIyM9pEuCNI1tF3nou+sm6rlQf9kdWlEvLU
A/l5oWDQOLG+KF3XTSVEwRDpqtujl64S9nABX7dekJuir9J1/xb9ZNR3/E7LhD9b
kUUzMT5VGHfGYX39BylJucW79rmXCr02OW2VSay58EPJJyAZC0T/y5sgZG/hB1QR
NDMJyKIPsWye03DO7IDc5Fp2OjrfghweBin6dLaLb8TwzC7sbLnlT/uuWw5mT10E
s2xHR9Jrvj3t56cL/4LF8y9n0HOj89inP3LumSikuEcDNEowd+5EM1d6mKuFugt+
O+H+9KFLHP+MWkt0mSvpsgLcLPQUTqd2WcQTIDUamLhrBCrQpT9/isaAqai503Wb
aElbXoODso8rhdv2TX6Tf10oHo6KcnAzp8hEZMWa34+ACTl591r3LpDVe7y9PYYc
QS5Byn75QFlZxgSNlxeKpuGFFB5cgtjMUAy+250tF/N60u3EiNR812oMlR2VslKa
1Fj+XLgTkXS8cuFiItXtHR81C99ojH1+bjvE0GW50uzYekC1/Gjmdj+QDsfV2xxc
um1IQPs+CJndPdeUXopvNW5HYJBkeK//k+4Tn4rj22WAGZfOkJ4HO8q2Z+PITUfx
cQvOFQ0xyP2KkxGUa5LRGF41kc//8RTcKLsyMFLKmtFlwL66uSsYeYYx9MuCgFII
cVCrMadwSD9NOivDtTsGQMqb6ZjtkVrBxRV2iU5Mc8J/vuZIJeV/YphkWhR+Y5cu
oojX/C257tDyD6o0ePreG8j1AR1V4C60lA6XaQV0nkmbtMF/859iXlk4yBOersvz
hsm2xl3I2atgBdk6xPbRGWwTQQYvGVyql4fKLQR9io9yImKZZ0WCfy23NkMVK/ox
audItVJTdjx6T9l5UgmZct5Go7zjkbX4gFpgM1LPasovA4l+jGXwgw2ivPZ9Cyo8
W7z9ZMvYHrOwmT1T6p3gn40VRtee1caDeAuijeNXiu0Ffe/uogJ3bRpPQDg1dRES
R6IfsoAfNyAB9G8CSHIX/doGS5c8oCrUDg9XgPltCgOuzb/7wnjlkWCPWCWBWrUe
fJjSKOrAYuoXAK8zhvU52rNa42oC+rdJep0r7OVgexP7HiIXkkiNy37O8B2zMWDH
kYEP5XmaV31Oe1SnJVl4qwOAgeqYwLDa/9DhXLdzwxPcfKpKp6CaYhlsoO3OU0LM
IkICFXA8HVrJ0xATuS1IQucRpQlUCkAcfGiVB6aK3cSFsAbkhIC/IgeF+9JlSyRC
38yaO67aiSlJQdwns9WqFma9XpFVAJfBn1mdpFYiCjW+PraHYKbTqWhfjpbpS1lP
WUbgw0ngL3CGyefE7yMGAqGZcwVQfgTye+6BFg9+sxKY4wokXANLqdFKChm1zing
ErRoDegT05pM2rCtpcGI1WZaALNUl/alHKhs9Fy8DkTDqMIPbXM5fl61CLA2LP87
KQ/xQSdgmlZtpzaLr8CIOvMfzq1LnGq5QGkOwCanmKuZ3PiY4Et8CJKCj0kIKMJH
XTd2jFg6anxbR5maf7IteIyVtd+n6gzx2sCwl5e734R+qmBpOPlJ/vmyoMFAyvfg
eeWXbzZLFohMfHZ3ZXVTlahmF4Av3uCumN9YCvZLr0xjSdjr3wSiEQUMTWk9dOrj
PsssBsgb6IgQH03fbz/jANz6e1Mo4yYgGaU3RApgdY8+o6CuRP6a4Mq2NPCjIza5
JceuhxYPVh2PJiX5g3e2A2zl4RhLxocemSFGBwcIApkmEbEXCOuxA7bEhvOcotUu
is77Eim5kVtuelNgbhc/BjfpH5gLoOkf/j66EWKQkC18kSI4iw2fixv2MgYnqEnO
V9qtuQEDv/mpY1OMWzzy5IrUtDs7wEWDzDm0YtCThk9aCespceEpnar3u314nWsW
wKuDc7YdHEI9kVe+ucgqqHSI+gvHT+Hua8ucNAv5x0P7D9WHthxZAJCRjimTYIFS
o7FXKtPjvF+buEBrn/a0QJ+zXR43NrTReYQC02paoOM/sGamwYtouibeDRBLYj30
T4NYkZHLZ0ySug2I9y3qzKo3hYna+4xG4bRQSiGrxDHHVSCrOKEgBBLYS+s+p8Sc
RHEdZS53rnzdrwETKreLaF+oK4GzrTi4BNyOQLSs7KNYefGgmlAfMKLg6feCoH64
RBSIv8IPxhrfEBSjDpDEQVii/5bG3qJ/az29GWpjQWKwZCQRBKiTv9eiyymcal7P
rf1SaUtFiqDX77krbw6HC9yv8UvcFY0I3BmnZeGfpzV1JhQG8MKzTUGZMJSKdVei
wLun6BrkMtG6ih7qsls3obJQLhK2J6bzAb03hUFf+XTsVSvaQqQpD36iGACz8th7
7q8QezU+cFPB3qzgToMKJoMP7VdHjN0Gd/9Xnw16qjhU83kH5fUwoqVmlD8MB3eO
IqgbJY+gp4lRtqUnfGQqENa7JKV50vDG3kyzUHJNtXqnji2nSjbpM7gymul3yMkn
lvfldn9dVecjQxm9NBsegYr7/U3GTMJ0QTGeTEP4NGn8JSGdTMnat72SuPbzeI76
WIk8AjOzdKXpPjPyI9Yjz/gUddZpPOYy8y77fihjCHqBpeLMTYgHqeEirL+MwDRy
3w0Xk+Oofhb4K3OTb7ml09NMVpuMG/piNxrWwnycMHOjfpFT7Iqn1n7L3mXxgLkq
eKomZ/BPHt9ra1gV++F5K12hItuh/u+Hf8ypAro2y5Rx9UeaMJe09VAszADZufwA
HkliAS/0QzCiVwD87AMES1tZb1yIBVAFKMamzIRlKwGqLqSXsF6BbTmfDK5Gmy+b
Al932qH38zbgZMN3FKWBwQRaUUPbrl1e1HaDDrM21+OTi9XLaShmWiYvhHaH9bbD
HCq/MFwXO1fweOgutWfjtC3LGTzAeSp0JrkJQ4rJa4Or8K+1dxKht8OL4rx2xbYn
BAzRvDSm+CHA5y71Zp6JCGh92TOApJWSUo1Zj6+FqGPjwwSGSIp2HgQBCLSN+1Cj
GlPUp+6SQInCKytX5WbvA+2Mtb4MqiTSzTkC6m78CMunFeH1glHjnVjNyu19AvmI
2CqX+qf5w4bacg71hw81ojpqhNMONcm69WFq9EdAoux5sXGW/XelBkXMxDaS9VG0
AOw/6mxDqwqggWr9GSrgFDOtC9VFiem5Jx85zs5yghJ3mSB8vq4l6b0cLF22nP/X
/NEsnUESIScgF+sjnVUJj0NbQULnc42vaIx9q5xvRi5fh28pyn+Xv1+Cv4nl3VUG
zxuvreYOvXt3ORrjZQkq5FYNMu8mtmh9i5iZnXYgqL5HOpsghqwICWxecMhRQc9t
JmTTWBxa4VhKwnf5T+SFGoO9EdIRoO1HNVVc0tTnZsWp0J6X/lPQNpYHRYPykCKJ
6U47vQtyjG8TsRCVmeP8bIM3mG+FYGqZSjeCUmndQvBoK9PP+5VnxG01D+4l6EnD
G9DGWhIzYHsLkKL3lzvb+SzYlP8UN96ETh0n/f7F68tTLHZ5zPyBUHGHs+DVX0dd
ATSyWqmGE9j4keU+6o9Crft6HBWjqOOzf/EyrQJgjcmq98j0M7lpF5/at0jbdg3o
E+3riHuGdDfL/k1iTbM6EVoPJ9IwMhxdnam6jMM3wTpVOFcXFnaIusVjwMZtfEon
V0KwhDFAywtADrfq+baUI0yZKIe0i5sXGi4X8bd62ue46kbdhxDW1ZG86tYpYHus
IxItLFRi6DrR8yMEfEDgAgsQAKd2V1YR2KvUvSGx4zBH9mm7OBSkTlvAErnSmHbT
36Rj8FbIf3xG9yUmdkH+YiASOl4lEMZow34gKe/e9bLe8S3Upa50fprnf/WIz6BZ
M8LQeXA0R6p+AcT2IJ0lMjldUOfv3uyt+N0Jw8ug2069CYOBF6DoR6DQtkXNfUai
69QVsuS+EFWwvyNN7JzgZ7S+BYoikNfleO3YYahXP8Xv1G9ge7H5cWxLqP6dY6I0
G6ICnuiaR+nzGcQKokAw6oc9yZZAOJYFeEZ4jCVDistWcd4xzawbCVJHG2ovBFSR
mV29k7/QTJ+LWwK7xF5Ex9UmPP6ETZdSmoLhclvRFkhkKJ1pXvNE9je/T3mF2pyh
0A1KOgtN2GPtxuWf6Ofa7oHoWS00jiovhQMZIY9AEaYKVFm04Y1xG/bQiPi+LHa/
aoA4i0KXuVsvvZTss/MA1HTwyqTrUXT4XUOE8y5a7+ctbsw/SAj2quq06gGY+IUM
TgPdKfOGGf10pP/KMgLxdgaNUy0qW5JLUks7KK/6+OIZGMXzpDneKvbFGzhEUNBM
EA6v78RyJ2qBFW4nLsHrxiyBvHv5pvPF8oz3lJnCcHbFPgBhDdh6Z7xgDXXV2zTP
omSpC+7HbWhkevS8H6gf8qqxkJqd9W/6uOOVxcLhZvyYHcRzaiucTFd2UwGxl9qy
ho9jvzQFl7rFJTPz9ksAA83r89rp/WhJpeUzIt7eNkZKdy3ovkViDUYHBDSmDls9
KWzfL8Ak5BfqQg7khlGM0w0me9TQwy1ErrTL9rkGfOMwTnsieK1tBsPvyk+aS8AV
+QeWIJKUyogFTrbIHtpOG3R5e1z9sbaMjNoWG1GG4w0ScNWhhweJgLaH8vrQPTny
TD7mehlD2Qdcd+jHrPXNomfaSZf8PD7bRfFH5XHqhPbPtxzy3iClAkmyDqQp2xEi
ry002te7P4+JuTJ7u4r1dNHg4lN73jNp02gCVDLWVrYEJtNmQ+3pd1Avl/Wimyqv
6cFkMViZlNj+WzzujudSRX7VSjWzh4qcOMp9L8Ew3rdVNf1ZKkDLM3aW3Dc7pq+Y
eKPqeiT5yIZ3doYXGRDgJIjoXYBkdMMA8GV/TfhrO+yhEt2XNaaE6/wiUXnKu1yx
kODEoWqGvSSu35MI2fwzZoIQua0k0FROuEAoxUPDKvPhkDfWdJra0CHH1SWj/mwS
4CrdFuBvti4MvyQFSrBxD5T9UZQHJ7guZFDhBl2Tr4rdhSI7hjRpD3g1OGATaov7
kK1gOFcsDNFbmNER32iOnKqklmXowUIeIVwwOnWzzXjciZbJuOgQHeJX3pLry+VL
3mBh/QLRaZ9Bgu2tMO5JpoTodN14Sh3vSU9BaUayjDj3eYPU5bII/fiSRTMDlsjD
BX+in1U9Gf/y0k+QLC4ygZ7atvq9hLUXs/FZcPQRcRkgdqxpeSb40J1lZHpjG+Jf
6Lo/6+yOwCVBpzbILzdrJ8XcMdKfrDuaY27KiKLkOhlXUqFAJ1btlv2h0Rn/4Elp
mmaWGK3f6eMSlslrvPLzhgvRlvGKtpcy+fuDJZ0/xnfFHqOsktoDYDrvwrtXXAhH
AMKlnsuR2eaYJDzfSqbmndWo0LU+/58QRWlsR+m34iUBgL1Ehb85xB67e8acl9d1
Xa7501c75NW3qq1kOuDhFZAHa3J4m/zQSeZmyfKQVN9uaHv3ST2jHu4oFacL2738
zEG6xbe1fw07N0kk5eIhwumSbTuXkVsFLSt+5hkL0E/FAN7noy0R6fUM9tWfaVh/
+90rx9NGzgsivhHMYAF6BDJYsZWPaM5ebPr419PJUFJz18Ys6d8kcTooXlt1jCR3
x5zWc3lC4ZATv+2FIdH4tW83CJYp3vGy6Na3axSetUw5J16Bf6vzcSR39RcKhH+c
vrtybo1jILV1e5c1vYuALC7OUiB++kWArXe1EDP3bumeR1uhPMxzIaxbdXSQbx2z
bVDZIWjE7TKf5e2QZDJXwHY8rLn3CRynAha1MZbIbxWAqhqotz1smuvn5ue9k60H
LTP81idMpMb1LBXadQz7Wz+hROq8zTqBcdmIo2mLMEsKA6KGFJYGzxH0hXZLTYd6
AhU6ExMD+kfJX5YfXIWccr7JXMZSZHZXTM2pbmkkYWt2rVuQ7VMIpawaIHSs6czG
d6GP0e+GdT1qAU630ajBq5cO33Zn0v6Og2EVDt6C2MF5kmp2iqrvkbxXNNZu3zmW
mV+SrsE8MCD2+1x/zJYs/+5KG0Y4llRzVGhWd5aFSlHSYQml2BPQOfhJZblBr6R1
f9a3CmZB7vM6Ni3mvh06WwKDWlw+s2GckzU/87I/lWgwNvubppqyNjE3CH5UcPq4
85rkqyYzf/f8pflYUcW2JNLRy3TijJrPjBYD/VhzRGXhHEdGinBupaFqClQWxA1l
PADkzPazUFVI/VwodMmqqPYvh7upaUuiIlXH/wL1wpKz8c23+OaHxLs5Jmz3/ILi
uRTpFkgyO1ifehxpXpRYjbTW9+tTDp6UWbEKKV+8YocDcK1YnffTPoiaLozDMI7/
vQwMcZyiYJyFnLX8u1w8ZCYdTjsi8ka130UwWLhAKMYfP2fsq3+7WS9zFwwxbTOc
9SJhuoneVPMREqqS8wMH7t/oDuCZkCSNMQhdzSScZkhojQzf0N/JPbBw+nw9joV7
pbYjjwpoOlTDOYxwx+QKKvmaD/b2ZhE+awrrRu2dqupePq3DC/xNxcHhrizisS/k
grgQHHhPDEvXgfYkOEV/dIZR36jW4N32jvF1BmsTC11Sff/+PkJNbROad2tqtIOF
/CmMpi+G5dxDoHNZjXz5min3gCNUXvijn0z6TdPh3XicKTNMxIourQ3FnDCQmCzH
bKR4q15K8ZWl3phHYdLApZdl8a0Zg42A3JrbM0CRi0jCjbhE7mWSY5/FN8XNrpKR
7lEe68WwND5C7t38iX5X+yQ+6SzslprCPRKKRrOj3waFEUXWT7SGYoYuCxbtYyDR
ENSPqlnHw8volBI98cbDdK3N4wM9JC7UJo67RY4cZUH6rrw5KxodD49CCWrLV28T
KLrTXmdTovty8WlHW9uwUZeOMS8CWbf3MP7HrdFQew8NyQd4b22P5jievec34G4Q
6HfZm7kxBcmyx5CWLbUqCiVJexIsEZ9SXnyZ6SoolD2b8zWApXpO2OBR8NksWD/g
tTvkzlitVteeT1qCxpFS8GisH0t+UHvJ6EY5//Pm7yfN39RxkGAL/Iug7eEFlndw
pcxQmaMUvguMYxM4AkAwuiVYnH+rQ+8xqOqPfPnaqte8anb3oMwFE30gMdAXTMDo
B8c4LOt/XfdXKTmUFGtLEGdy8+J6KSntqe0Fe0I2HvMKBB53+qdyMbBQWEktGBgA
0/imEitDJsgG1XpSNvzBLAAADjfoKk41wunuPEaebKKrHeKIt9Z70sGBZNWHxmEX
cuycxfdNRgro4mpPicHS3M/wG2sOTWVqEjopvpY1L28fKPRPNX0ILyic19FTAu98
CZBgXiP97e+z3eu0JQEndIqdsdQ9o4DTiqqtrmMWvQE0diN2JBv5drkxzmBVyw7Y
ORnql+aRsopwT5vOtpAY2gVIYDPDhwadc9tXNhrWUbVBVPLoHQUCG+Iz3yGJy8cL
skrIw9zqmaa90LhKNyzN9jq6MiUGlYmeok6Z1pP6zwlzByaK7JSd7u9JQ/DYiXTB
I0IbqZIClyzKKBsKmAk0e2qmmL0eXSsrxFbPFs/LQocliEyjysqLqy3NtdAeIhbJ
sPJlN+Kcc44K+NkuRqChsdxHjSY+82atbFod2xWlX9AJsVCyi4EhQIc54r1f6hvM
yYUAOvs2xf3yDQp5xHvxbpYh2Vbhh0rOb0EZBIXroBHpgR8941llTENW66h4ThK7
Si3DiK2CgiGUnqUo1WXVahPmM8NHpLf5tSJ7e6cXFNgTPMPMZWIZDNtTXioLaiQq
rWfNDqX68wY2BCp1hHvDd5cDqcqF91T74zM/Qvt+42UfY2r0ynIMK4bd9l1TywkJ
LugDsuKWwO8jAOr50l8V1gnIlq/5ss3NEqMccElP05adeUScDC/I9BZIUWm9XBaQ
keoOdoracSzG/KRs3AVVibMvfDlflZV3eh4jJ/OP2DlNTQqm9FPFLZVNLWOokEHS
NYtmUPTDiRVHOB7coLlpk9Q7qGBsmXYl99m8MVPas+xevAsN0QdNuAXF3UerFifB
XBMC0XrkI5s3m8mj1YiUHBggSG/2mTdHIqXyEd3bSaxmYKFNO3TZmu99TRfphp0r
WgJCIQW8ShxbDeQU/5//VL9Hi1vaw9f5T4W9V8u94TDEnAiEZbk3H6G8M9HAMY4Z
2cofjZHHaDA+QUt257DTlxJNbx6QztaNkV+U29ak+YM0UKdOxS9xSrDnekIpc2Y2
Zv1iilV/WiDsVuZZRPQcusTK1c++TDyywAaGcRLazrwmqd1JydZ3qOild4Rcf2Mp
xRuigtNojXuEtsXEw8kkcdnJ7NOadkvXIT58lNBoceiQkkjdpJFODQaoDW+InyGF
wXD6MKFsCfdfD3w+ANXxdKaBSROjh04gyPpY8efN2wbfH1UvxYf3fqGIgNcfu7e/
KKJ5OPLT+4kmJFCNDPHmEoRbGmV8z6ipMwvUuV2GobYG6ul+kvLNvTO6Qaf7YtJf
V4TqPIkVHI5mgsre1jtN+/CzH1V7a0N5BECyEfooMCQv22PnT1hIajfuvgWZC2q6
Yem15X2d0jHF8SjXSXb/HTDVJpRN61FL4PfkKvfOumXLWl9+i2KaP4MQW0mh1nC7
CGy3Cdlb6js205Lh6F9VGgFuPqDeEXePN69BhdR8O+N24f5qC6ql5mwEovU8rqcn
D/CIb7fWn98/TZTURbSk/ruL4TXWeUbThvctwis6AHWNq4wdQKWUQaKKLX/k9JSQ
0TQUEBKHMwVBcMGj3FMACgXYr7ILuXRVqQXkXDV1oMK3Z0qrCEXZvGTWGIv/BJyi
xyybxz6k0mCE9Gd15BbD6xlgODT+Fv7PkwtuFTG8Klc6wFdTEdK/17WasugqtrY4
FOVfs1IL+7JGEqhy0D6UZ1qWg3UQuY81zxYntcjXjetWn5QzTzwD0ZebrYkATZZX
Uy3/U2qL4ZOAXorhxkWPLZd3D61pM43iBiz5tzyT5eNPZUh/9LblhaNroakgZFf8
X7icZpAq3LNrHC8LRfEvYiPdJvlqmpgOJZDtGHjLyVuaUwIo/LsEDtpor+zrVzZT
/yHbbS2iXEzPZrb3q56fkq+y9FDWB6k/ltlvfqeIUg/ZRSRQcNyB37iCjIcaCJQl
7Wtz5BxcfQHjiOMZA5SfSkjy/8QtSCEpVOefQRvwBr0Hlga1bB5PlPO+WLIgeoIj
7JidHqsW0d3mEspwXAA+5p69IEC4w9HgUJFsWPUgdTVEkmp+u2R8GRJ1OCdeotkX
XJEW099mRd5gm0P4k+WKnbIQz+g8sTMWe3ZmFe7IkDxE5BzYnti7aEtS/aFf8m7q
ENAGfeMP44Fv1TcVqvyI7ST/r22g4lnTdngYdTZ7JMeOGcX/5x9gCwKO4xB+NGuG
ip0S7GByVKE7gSPxCEUy4VMwuFxy95awd0sGc+tHlu5uV3xP0kg19PrSoIBAE2nK
cUku+MUujehQb6exkgJGRF2CH752RsWByVa4bOqxhD+zkEpUwlSer4ye8obk3tAj
pz3fUQO4uPRsSSdRfgMiH3b7X0xsz79yMnVuWsDczBXohs5Kh+dl88yE+tzAoE4F
ZxQhc7YZJzcyTHNvkhnaOiSKW8i0/dQ30pfLwVkVwzA1eUlXqSsEd1Z7Z6f2dI8F
1SSoc8fW0kYnotk7+YpE4ysqCMfuQBohXOm1v+hOkppM9zTn9q9jqjoZW+ypBFZj
YumS34BDpwmJFk/nIK/cz/vSqyXM13flDjeE20hh21uSxt0PKpdxVekrma5ZiY7a
otPzn+Nufc6IiBgWaNg9ezE2uKPTYllyNQmY+SZgTZkd6UCyAYj8KNXQAB1o2vLg
SJB+2zDY5o6WK73BvqOlDTUzwQacbCdjR71QtdRctd9WWgPWMsZEFM9PXt9Tup0c
hxyzsJuXV1pVtdavn4EyG149JoV3il/PjIgg4DZ7uVaAqFGAgEe0g7nejwdA3RSL
E1xwC08iB+IS6xFWyaLw22bidTqOUk3/1J2/ZoTkXfFmePzPiRZ/knfvVDvC/kQP
WnkOL3nHSbZSXVMYzRF6JKjhHPcjKafNCTDwpE/pk9M4PPuTyVovn6g4NE4nC5Mc
kMXu4Yasun2tW6yKB0eZWjZzLwkjwxpZNc5ah/SZaBND7eCkhdONHP+7YZoIRuwk
Fv5NYR6IdP9AHvhJ5/JmdlngbR6sWhJ6zlpYCH8jaC1Ai+NRv1cLyydFj6h93zHh
jtc8WudMMYNspzyVUzIJDq2QoZnSDYmXuB0YiyDo1aziCrhLcHNSoumJLXo/6Uqg
OAZuh9d3Ed+0TbtHBJ2A0bN7eX9+YjvgZnR7VHWp6p1MGudV5hCVoEanWkARqMyc
RRneVJ4VLAyYVHY6ojo+38NdmN5AYzJPENUAHTKlJVRo5AGOR+fGUg34FIUfwpCA
b3PS9II/cxqqEfn3HE/Cx9z7fWO8AZH7hCq7yJ9fZ20/7lciqU53Kkf6rWqyq7lC
R7O+7uzUHHWaSTNhVvYRv4ZjFb/D6AqfT4cxtzMXZA0d6MxCtTYslmxA1MT4+1RU
Wd8soEuPzQyAuZ8QsqFA0+1wFKrGT+Q+KZMK/YAGPMCf6uSMOoEf3bxAlJubQV/J
3Nek8iaf8f13JDtnHZ7z+acGagjThuLhpHIgEIfL+TsTPafnE0jYmT3yDKWeYMCc
q8K2jP6GyRVT2VrNysGOOe8aYiOJTGc8H7HTNkJ/hdJrc3lrLoE2hL+NGqVQF5x+
0v/bk88GyvOVaweUND+UepwAqOTI1Hyt1kXd2My8oVRMhy2RbjBlFubTZoqUGuiz
R7WsslEDSfgB+n9NBQKpBb0KxkgBydkwbhKFEBxBMj1jQ6PBNvCwjfXb1gO9S7nA
oWpPcN0N8K/yXLdIMEwDsHg3FkzSK220RtsWKVY8KSuQy6XSuMgc7P2peoAom81s
tDq+SbG8g/fcbwxltciYfxOFeKqynKuStLDAwuiFUs29k97xIiSxW9EU4zVN1XXC
nSyGalawceiRPuvRZee6CpPHJIu2Eb7ZCXgO5oRJEGrV7FsmKDcSkStKgVNddIgR
lKF47+/oo9roSMMb0cJ0MptedpqClbpmqn++/t9/89WM+XmZZt8YzsItj32h+Zbq
Sm/cG9jrp8lJDf3jd1vggLAoiqtSYdYy9kOg+04Vg9pb8X3njHAI1L6UUUN5KmK0
FRjauqhf91w/vS3rn4uJHb3u3sbEcJddUFds+7Vvvyn4qwfAhvBbks1bL8PeOP+N
1oH+CASEGH52E5J2LseVAHmlyyUxJ/6XRQ5XVa8NFiG233y3mUDHrtsOGuwJgTh8
sn8Er1SJdBnp5OLPQmIY5GFn/SfIM/pFzZR4IdcqxmpGp5eBOaTZuOl/DG8wFwQ3
o/JaGqGhIkjshD4r2vYJxQSn9WK1FHYVBOoi3hjly9Gd3zghwYQQ3kuUKRX7OL6z
J/++m1JZaU+VaKuqo3esTzM4J7f2ioVtF8k8X6ynBXYK0ihBVQO6ulYXM4jWscNX
xE16zejpQKpQgzOBC66rVXHszuHdxPH4IStKjgubjhqi9YUNEtjN9hPWnMKhDZRA
KaZ1FrXa5OU9bpem4jb4ldot1v+lT1+W75r/6mCYwqb2SK8kEEoqaV0oQAA3Px5P
cezkEqNQmALHBiQal5tf3V/8xWz7Tic967jTWQAC2A+BykFWHmfxsa4V9RetKsW9
Qo83Hki334+GE5Emke+52PT4HyT6kKI0RZrOtSdp8isUl3mn+/eiRtkyhD5thKRg
QwwuBzSrmc6iZZTwlWVu7Y6Gi4mYxGj4tuTdUAVjtYOl3hmCCvWtqipsISjYVb7D
PRbtKXxRFCEHZ5D94AZznxtOFhypZPWCRfFVnmENGc3JHOLuwr7rhTtfkKaYA0HM
EORHcubv+tnSvvTKDXD9pit1Ll66mCTshmi+OMyrdmrFuQpSHbxPSbSR6S6YN5dw
fmx+N65pSZhckG8LGnBEZLXol1X5L5QR7tLKVoIoAwH6huBRnS6nMrRd2QNi/Uxr
dSiZPLMKniWgtQLJ85embZ09HPOLCD7MOM3wk9u/A/SC7Y+ewHlmWqOw41hsJOr0
h0r3Wp3UMAcMyqyPQ0QyoCFhkkpYoEqgPep8BSvA1cvIc3S05ZKxZ8+ytVWT3kpX
Zi0gIeSC2rJI1yoWcMzNVsg3XPlynF+IhLq27mdrJ7hA1tsuI+tu41OrEqrpfgZM
grhpPLVHi3tc4vNDiCWl0OQELz521p3yAwG2c4QNwNum3WMVeROHV8lIeDbgV0VK
UhOqb3RS/h538ZbJcHr1Ds1OiCrzPv2dcESsGgelLu+APSidbakWh0Zb++z4Dh6t
ryX+9eh55VN9vdHYwr2FUL8fxyqlrov5o6KySsEf45kjSJ5TlOc3QULWEZfn5qlj
JqbtGxO1r+Gkdjx0ROrXXJrHKXNVmdB2yYQzQZCU6VfhD6HyaRKUK+txIikx6a0j
jkIvkpUNWFDsNNnaFfnXDadD/GZMg3w8MUYaLnnUvi0xgEvZpogQ9o+ukbRwA85J
Gv91m4oNADdlvYDQ7s84ljm0XfkvLCS4csS2bCIHi1I2UWEjd0mw7DhOWW80UDL3
FaDIzPP09bBg7FzzPhjg2r5zEqcTAlnZn7bzKXsx8FfUM2Njgpz0TrJKA36YTwrq
tzC6FcdAyJMg3klGRfzUx1g+sqZbKvUlEFN0KCWfip6WG0P4sw6Fj6/rn79VwudI
Wqz6Ip1cHGfTZAE5AJvfRKqIfI+5G5PEozUHsLz98moHyD0tV9M+XwfqN4s9zkD+
xyW1WDVgfMEsadMfnzIt53gFEliuCUadj62Z6CRwBmIf4H7ZRNG9JiqDU4Mvb7XI
D7S17RMSO4EmDzPOKpro/m/cD+PNVPL8kgwzxwE0dhBbBbIiHBtUi2Cbv7pdizrP
Fm7RRzuIji9hmg3mIRpgmr64WL6nXYaNfatj+iSEGlG3QHkMBkzUJhx4DXuipM1o
gkE4Sxopcg4iLIn0xXLWCFKRPLE/DP9D2kxEGydEnOJ7WZUij3lKzrIdyFXjrZf+
WgIf8LddUNojr8S0GJcggCb4Kn7gL5RVcqOBSz/TDwfY6+9LiYEoIN3Ke2W76EeK
koGnZz/kTiWNiV3dhXI3xm6AjJkAlOOLyWGoRV2EIRO7Hew8ciwugPb6g5NdGf7h
STqF+gdElnQs0EMKRkU/Ae9AS5uF/ZqRrSAQSp2giNBDn283l8+WTDsrciNwEPgn
gYA7y69Y3JSyqAy5wLjxgtj9zxp4sgWmMNIHS2Mps5AHnHzDT9Vt/HiWsZBWJvTO
nEgMLmSvk5fKNs5J5Gm2ElAfx7xSfBmMWfoui4pEF10khzFLJfohjJwDR9v5blHw
yRREX7lODN535NOZPINYkESLGyb7Ukl0yh+7OnypcQWaRMbJ7faHhEZjvDu66PMr
WHlJBRCGZoeGh0sis8qRkVdOdHrF+sj2TpwsjaBNgIK3fJtDsgt10wDKLZmM06Fk
Y6R+HOwsEJoRqLgs9Ny6Tfs/LbSba3P+FMCCCC53/vdBwit8cBUu6FhDUExzjz6J
WpzK21v5CksuzKbRakJlLorn43Otw2ZkvYePPdbfxR+KaMJeUizOmmFb91vECmWH
sub3wkOC0fqVK3nukAT2Q/kxYgQ+zDaZ5nimOoWlusGpJXpbEqt+NP2UcCpR8Txv
IBcTGLvYGU4a4FtbQbLOTBLIzDkp5u1T0AzXqulRaSuFLyxGz3aYWIl/0oWpHQsP
002XEhtGnSVk+gikKtBXH1u2KNcKOwRgVncJkLT30WAKLxzSsq0mcnn1W9VtUp1l
3apsohzcJED9K3Eqvr3M8TfaJm5Izzn/fD0U2QeMjE8P5LZNXT1ggTgiqDxi26qR
oNBcDnRqXoySmmrhAbx5EdAXKCiXEDRjN/wrtN81MeeC34EKOkqydenq7iZc+Gg+
BHLGbpSePoVe0PEJUy/KwBchuVt4xjz4oEC9GQb+fc79Q5mNlU3VsKA/YO9FtVTr
9lWPqocYwJQltvU6djd52MQ9JoBxJnT1pTbPJ85xjMMI16gOKOGsZSzBbcY27vJu
kSLqDFyYCqCXDLTTfy2avaPjC3uc0LLCDyUV4tpShCyu4WULZAm/bRYV/RibNHrV
EqJzQ6HL4oHAwWFYiRA5lS6FU/qxQ4uhuwYjIgFr8VR048W/j7p/G/EhW7QSxv/k
A0YHeFqXZP1CEc2hcUqvFCHHPY8lj2fntGXIkTm0iqIDnlifcupD0P+DUgu+pgA9
ZNfTfkEs7ICCFTwz8HJPiP8gYIc1O/g/ORLclIZSIZ++D5DDgZg16xbFfnMOyCYd
mFWhc66UG+tpIrBA0ylXp0S6ISH8ajlEGRo2lQlMRsOu/caLsEUDoh8PLPwBGB8j
LEQdp7fJhGIzsLfdugRNepP4tCibvTzNHPYTz1d6Ott3dBOZjeMbhCe8oO73abyj
2taQtVGqX4Zfx2AJ/nVGR1C//rzmh2Iv5kttp4Wr7bmvSjYI+nbyn5ARAmkn0S4B
yMQriiOSX+WR3eWAu85PRhGSiVhlf1EC4F9tHFpkWjMC9KHAzQ6jOfkCemOTdaOq
pMEU/DQYEbyT5pmz5SOSR7e4PXf2ks9W+ZgLCtFNGYQrxYEKNxML3U9iIi7KPhZI
tc27On4qY18EDNeW41jpeaW1tR988/AK6Jkodv95eSI/MIuz9Ig9jub1AskpL+F5
+JowdvkYv85+u8YDMy6b4sYcAXdEILIO/3rI/CAkL7e0wujHHQIuR/4SIWC9qHBV
oqV0VVJ4kmv9KbzVEUdTUcL3f/olxqwdEjJdksMvfpVEWlOP3Ucw5xeaqi/fHHBF
g2RUoyHD61ELb575stO69hl/DV3bsJXMKxcyqUdy5OD6azc0ybi4h6sNw3DNQ8n5
BYO6QnE60E15v461DPDP3LaIG+p6qSO0z4h2nv6/SGU39jSfRiRLj/HaDHsFjNKv
GJmiD8jlLatQX9J+I/X2iMExozLQTXr4HHrkZAeHXVuYrQvdbpOxB1QxrBszE/6u
c/FaCiZCn1zL0L5HR7e797fnxB1syL+ZPWl6pom9rVQDHUHba+3stWyv7QyP9Boc
UeGxQCj/pq+45+EcHOyMyxBgM7+P38yA5TUZPXV0Ket7Rx+ssAQVwuF4UjEay0UO
Qmy/gmyLnD2AWx2XNyh8UKE1c6bzAk5L3wFu4uDJVrw86iFwSQoKSXnSg8iSWzey
XOVJ1pdtjf4t0N6PefzabCD0zvdMeuaFZDc74/M+jY0a6y+UQYVmsQvtj+iJs3i3
LtTVqKQ37jpAbu+7+UsE7Hu8WGdPgU5xmrtqGHK+MjW/RfwSO4k+HOpiNV1FfeOX
qcSS7z9MtBjpf3KCvMq1/Tqu/6RmtrO2TIEYFchNmVGZtNY4JQj5tWaYFp2+fzaq
T7DMXDjmfpck6VG60TZj51cZt5yymsgBx+JK14fYcUPhpEv7pP3pNAwHzmyLQfQe
r+Iqa8/Y3j1uZxZ9d0alRI9WwkvunmKIw8nnF+xRsCtwNlC0Crig9SDKDcwFqv0d
64J6xXRiyKbdopnOdfHea+4P1c9Mhltb6ZAD1GGXgmhJucA7gL3fZ/04HqFVyyHk
lhfB0vqxcmnQR6FOdLEFdPNAmyTWcj+dssvREQ8/FpmB14jivhIvViNos+x1NxxR
ErAvEUgXE52P2I+d3lWCscZxPSCjh4j/fILBq7J521rERweumT+MBfFvWaCO2g9O
/74V10BHpJ94GzN1lbp+w4pdoDdYfuxBDqHc1WvTItEhKPMIXYfKYo1i+W1Qutm3
/fWTE4nDVgjHTbY6aOl31n1Q8j78tnr6AcRZogD6HddLzQunoAumqNIs7RjVQ70n
LwOnNzQ9afKeJhS3VwjUsaNZ/ciAR17xf1kw9CTXCPiJ/fLg70ojtIasSQt/r7/z
rFHelELfZx3oyuOP22Xmh7LOW38NypaNbN3DMAhUf9yjbIM97ItxS7JZmatW6OHY
LcMHI7wMszE+nUZje5BWKYxtt7/cOGTGJWc40GiEl0gfr+63OZYnkjZxC3PXfVxk
Go2+I5qhTyWkaViUpsVUuLdyW28C+ovuap/Xh+NGXgbj4eoj/rWtd28RFFi14Z7O
KJVG5qbS4xuv91YeHCN8FZe9DXrbEa1sZEKOJX5K6+RBYnI6hK2VDYwkiqiLEuG3
VRqK1u8g96ROaNqUWEUu4SQ/v0w1McZs4zK6OkCUCZmBaAm+NyftJaol6GHDZAhZ
QcCLdojn+FHUSYZ/B5BNqw/GoYFWe+35BfdOUzQXNqB+UrvK2ApHH4hpyXJb5VDC
ws7Tm2crqS8Qr+Wpf8aUUXdYlNwID0B+aSIN9dekDAwPdqMgNg1Zt5neOyNgVho2
R+wL/kUa51zjejTWUfqXptq06WDytHjMN+nfdpiJqSHSUzxNUVk19BGIAG0+vzHe
8i9RmtkhWGTeWDZvzu0VYVmDmYvM0LuzyR8ccGAKiw9R2WZbMgs8ZjzGCzWItHyl
5ACHYfko5zbwtVuGul4DX3QI260Aq/xcSUssCJc8l/sTwrOAmh06F+sZ5bNy7q3x
vp5kr3tMJfN1w4/BCR/raBr21l5OTW8hBv4sStIIAZ+kIM5wkTrKahRTg1LaTAjX
Hiw5fwDFn4HBU32yAhjSFsaobGI9AEDB+1m12e4hOKojNfncXi2pA1aLwMmjhn+p
xj7HG3MA6uB0DRwj7kUBk+y5LPTJaSoMD9Gdqry6omk9yccGzZE8DyJU3lWW9mM4
ETzxwp91KAyRk2uZk3J8NGfvxEEgk8xBshBctJOfG5KThQevHFqCpDL8AxTjjnWK
6r4ilLvaQ9566MdgiuSL/r0Nb0gRdQ0raEAheb/HfXws3/WNp3ZzXMQ0+MMOftsd
DGRYnGiV1FWG27jTtGVn7U769lzKLu5wha5fWkc023vHrAUQdKvHcbslE+LVG/Ux
jkFXZaz/+UVKKBvIsmv49B+WM8S1m+CmFjsJKiO6r37DeNUXpLgr+Eo8rKgbYa2s
riP+vSQRMW33ANuZv7l3BPTsrMuEfUbFMR6zhGzXeHGkfRzwKgpS9Y+GB+cbMdd+
rSEIFXYnf3uOvfNSI8EuXuQBf57kNZ78NG47vUpNF5WTghiCjbuyrOco6oLBZQoa
yjycaQSGXALaOdpbQax6ttmOUu5YiE04BaQoq1ri16hfHvO/CoPZP8e6BAJojY9I
sT46ZdLSkEFVbqBQ6+jiMOZopjGFkB6NWXsVrQswV9NcPPUDiEUbwZgK64dulFmf
tYDEq3PtcHJuc6xOJQSYwka9ioe3l2pHHqQzI+1NLJFJbr/QxDv9Sqh8rdXz2t5x
6wISAcyv1kkz8TxkmKu0Z8G146hzK0AnW5HmkZ+MyC5wlVEvnbB5x23FT75N2v0A
wiapXg/QaF8M0v076b/eL3BEOkRqqsHOsPxSRJx0bhE6llv/bTSJ+ExEyMiuOqAf
DEkRvJyJ6xHMXjeQD2l4yr+l65+Clvz8ok2MjN9Nou4yakSl1B8xujTRIf3mZ0Mj
59JRjLKvXieuHhm25v7r/RRXQZcUngUnzH/uw946T2hv6Qi+GLArw3TNEXKrPQXR
CfpQRg9EpCYgrgDLc6yDpPcu13vUcRqx90riiNkIRWib7X2eywRYdkQidJ1erEpD
9MmE6WmFFTMs7QctnHpa1WtqU4e7kezzIaS3SxLvFIdvqWxZ6QqI/a6ysw8G0Qcf
Kc3jS7JGt5jcYY0+9BVH+aQ1e8GWo/sHIS8iPnaAH8qzfdbNYxI+GIfFNhlXKtOj
4735V7l+olsvfZSVA/dJazRFAINoSLGX2IYDTcCsdFIKdY3yYzrDmp8aEC3BH3cn
6taVyVA9TxOl17Mp5aH2HIpYu7TKaWjvLsai1jtUd17gSmMfvdlu2YktKeciL7PO
9KlvnHIBUACmR0wTYhZ8bJp0NrT3iFpKzLPxi7cP9e3AAf6hO7TxylsAkBEORlEl
BiXi/COdIzisemCMd57hTDBxDSnc72WVfZrFkgfMjr8vCCQilZVj8gXdgsVeOgOm
U57k1BbNW4M0iEWS8XqbviCUNaqD5mCfEUiEyD/HYJqbGDotb+87/ZZApECrC1A9
3WKKlVbYCbD1KIrntDM/mWyyRSscurTtgDdlZ2Rb6swNqNF9ylk/ZzsyL7ADVJut
lUHUL5BqLMRu1AogEgTAxHj6nqdJnT4eYn2GAzAIqtD1wm6BFX1UtZDJ30qd9YAI
WyOO1vYkFUHGnfpTU6+ra6wfz4h7F0Hs2cDfD1W7AITq2bAi5EkMIZQprY47UT3B
hG1hb0nOS1rx16n2gUmGxixFuLKtr9ltOkXOhd7PW7M4JzJdnt6+Wum9F75YojpB
faWzC04sBpJN/YzfXZY7B5/U8zXMwRqnJfcmm1ViRssDHRVRXTbTI2IUF8d7wyBL
HlD5BWUUtOkwJ7gtpHWVDxBcozXQ0H4/uYQ76ZLyvr543oo9m5ZeEAKtx8POTKdI
lU65pdxXAnSBArOcLewecatYxPEkwSERXv+kqLmZOyN53TLJ37V7RkI28LvN8vU7
rfnd/1nQxv06hz1x7asuklW+06ahL6Yoh+Yfp3JZi4xcQY5naWvKO2Hi/vPqx/hI
yC+HbT8rExU6bOdP83mIm/y5G/x6FlD3ydLKOHNJ299LRQ5BGKqzLPHB1P5j0+CM
ao9IZS3VkMOIx6vE0m4cCtHWEKTGL4m/yRpW3U0oFvbDHf1D5SUW+1Zj7Jl2jdov
9QeftY9x73LTIQD4KjNLF2q38ZZFkAYTBiPQv11Lj9dwwlsXoyR2Sxf21ucCM130
PUA51+VRZeKDCgeTZmVyQFxlWQuV69KaW5MlG/FAlx0uOAd+OJB+RnlVRePFHPn6
66ab3hLDJ4rigFQU7d8G2TKSfPept6X0x9Yh9hDyZlDXvy+aJOcbJbTqtlIIEoce
nLihoN/rtNR7nJ2oyxGjyO0gJu1nGwX2fb4hCud7l8v8h1LT/5N65auYEZkCQjLK
EEprc5EBmEC4zVAxjBSizO7nM344nOxNylAeF4Yi673yGbm3sVmjG3J850Q/IEuq
xa1Qw47xQADBt2iOztVe5k8HQ1E45AoGdws1DxiHSpAkkI3tTopkoWmqWtwEHFs4
o6hcynhvL03IAbbGNgK+5EaOLGDg0YaKw67FAdLkLyjprvS2JVjARhlnaQvxsiYv
VaVy0dJvIVHyhLlUtRjpxyA1eTT1w9wIMb1G5J3ghDboaMbNlDdWbovYEAglFlou
NmOPiBDJZbgl8HQ8FfTuc8Fl7sqUW3OiPVthpMVKGr7QHfqTkpeTNEKLksekOH7T
MlZPzQtH5EeNzW5m7IIG/EdolgNHctbJTgazhR+Tej3gXf9rATjk2Cb9DzMv6WMf
a8MWg+GLKD3CQcW1jvzhhU702ZasinPPhaYi2DVXtMnFRklUll/AvNTIBYh8dqcj
zK36liyrnzc5LcIAjGXTDQZk8+ci5PqFfRNbcyIK/nBONFlpJq79UFk73UI4OHjg
brU7Vrq4csc25C7bdJj9oHxY6R7i3xC7wb8y9gG9eIXXnz5J+3XSOF8HsXlCHq4a
zsDYRFBB+PViMFI0h3yK/9xXse3Z6/xkjghu/IjgZ2BNFnWwcITmVR37n8QsAq57
sb/0s8gIHS0E2FP4aLEkKCDI4FRX5ARVp15QPFbw6rNAEiZh8b4DdJ3/Cc4OG8px
OQKt6LNtWajTnwloCcLVoViMTP+DJ3QLo0mBZEkt7RxkB85OKTYTyODcNoYFuGx2
62713NU9JNmxn+njRsSrPOLEhGMWEt/2HQonKQ628em/4Wgwj6qdrcjxZmfzBXJj
HQsH/Nacr/p+c0cRtEqUbgWBLgQ/UfbJoHQCMiHpbLRVNXMHviAKgqGCf7If8c81
zX3fkJG1IMZDTryhy+crnI3HjZBsVgzVIfBmP1J/PLHofwKMpsPuWalu4ey3CbpI
E4426vjnlJOJnr6ddVRly3XMuKuSBFBOvH+jTaLaOevt8EgIn0Y4AsOc7I0AoR3G
me/3giGe63WVHldL5+n8+Vibh8zwUsIILXJ1EF4ePq2pbzQ63tFU0MCcQG+XldfL
9GfwWlO3cRKHx3XxuGphQ7Z4KQYarW/xfyaJ+7JTO+uHm2Eb+KDPhCgSiyicfjsj
U1SJkhDjKMphh+Df5MG/yiycknmFiOTAeLmVNjC8xWunezyhdeKUQlx5RxNEhSkD
Jv/ngDqqt2naWhDDaTdWEREDr0Lp5mxt+rYUbcbWMDiljVdkIpYP2onMN+Glto95
n4XPG1QBFgHa1O64jxv7lVEfgyP7q4QKU2rqn2mB/XDTKZWhxaBdbdvOzywFK441
OGfR8XHITbhY9lxXmrARptTKDMe4C5X03qVHI9vsA3YVZbUqRODc4HkliPy0fTcP
hDjoVtrARq9GIDVjUzFgP0A5srrfv8Rzj2Y3T4OhgILs09NvkWBNUGg9THieD8BU
OOsI91U6DQ0EPadg288zEjM58vXxi1sKCLn1EzBo7VAmBcDsv8vq24n5e+ht2/6F
kHM6aLHFV7ASMN71WOYaHAK+aWu7ZgvZ6mqJ/Tb4UDru7w+XhnWfORkbWNzT6/1e
/2VKn4egoLB/LlHPL9aTEvMsKl/9VuS58+V2n1G0V38kI0HyELl79vlucITL+NJS
7zIBiTbYJg/E9j4oXN7TFM7yy+IJwUHCz5/4wMH0p6Ma+qFn1GVSlz565lEcDexz
fk/E7BNBz4xnW01t9YCow4is18GD/58EUdH9UXnJlAJIpUy2OIg66Cef9WXddY3P
9yQdqKgi1Q1bpKUIzmtdyIpTmG3gQ8YurEdWF72A/YZjSm7BkkYd0OjnKD6zbmCI
mIMRS6Kpu8xhU8kueEmVQFQrbEIcBz41oytDmhnEJ1GFrGCZdHLHrTtXiivAilfr
BQ4xkIKYXkdWoO2BziMhcQfiBq1FY4gc1bmroATirfAFJJ5R/oJoIn+Pt0txaTUA
qO/10eFwdZBxcZlttpOqdbgwN1KudrUS4yzHQGdboRHQQqJZdA/eXO/84yUFc7YX
Bv6Ax5XlAB9fvxzzgs8XEDgEJsS8CODlQ8nlLQpnkhFuyT0Ld4EtGsL0nts7tETt
9v81wgDPrRdVbbM5HqdlOoIbAXcD3Eqf3hKUXVVHNL4P13jJePEVTX8KcwJ9z+6N
yD6l+EXFuW/27ynd/PFeVWYLXuYQfr1x1tcUWEChdxKhFU7l6wH1WN0a9bFiFQVt
CBeb7D+lIxmWDkh77idhW8uZCS2tBl3VobByc/Foyq1pvS/nJ4HKFizDqdx7vzCw
/KztyAXDGcd0lKEydh42LWcAADFl0T2k78DxFxvbHfJNtoxJIwAZ6s29P6k5deKK
PjTijYC6xNw9FJgM3s6qb1BhHqJzkJGfVi9PDhc0WhsxT8x58gIngHYxjmdSTYhC
8RFVJN4P+gahYkB+zPnnMZNsZqdev+PMS1nKZnmECVGPHk+j9059DZdM4tJ8ZuYh
g9IzMnACXdXZ4RinX4ZqZBgGNYeJuBBcy14I215U6m07l20IYDiJiMayRlHHU/s2
nJDcD1AyA8HBDrZbOm0E+TZa984R0VXnDeHByWncKKeHdAv/YhykimOK5M/zK53I
EXcmNvJ0waHm77dqQ5lGEycz1DYncF8Tqai/vqoavlseQ7qqq/rb7wC3IsPyTXCF
U4faArAAe2iqy1Tzfbadqn+X8Z1xH5ME5oQ9aIILDkmoyFCxdRbslLCAdq0GOJvH
0BXhnZiKYPuA45hQ3gAjJkK+1JLwNaEq6l4JBBAnSi1Vok19ynEK5CmE/nSweENl
bOqwL9vDWbJM9rH/Mt7onsnmXOatwQR0FuJtYz9gV7Sssnp1gCRDb5T3ZWSCT6TV
g5UdhPq5yFWluM/b14lWdNFp04K+Q1ucZTW3E5Lq0ElJY+GIpTbHYJrDHgKqnQE/
YqqZE9LX3IuN4RPmNXgiMFbDmMXomrsTOLxmctgjTYFbVQLxGA0Ot/omOnesRkth
FK1vHgcfKvOmC3hSiS4uM3jDtMHbmtOl8HaQjfCeFnAzZPiPS/Ltgt8VfG02Bcx6
ShXV5CgBhfEuhXPLRh3Nw5l4Z3Kt3xQG1jbUK72RPFaqFjIoJL0a+AP8UvaJGmrP
5VCssygJPFuinbucb1HN7duUNyeWfUjz3baKhYzPGUch9mZVdwSqVVzq53Yd7vEy
cun16h2uJnwg3fD7HUMWRW+qT2DU3yV5rSua3VvAfUCBaatdDgGjVA7N7P1zJaKY
6LnCL/6/OxlJhdnUxHVPpFzQUJHr7Jb2nJ7DEX+1bn+ChzFL3nD6OjacYjc0q18P
qfIgA0cFXHoY2NKUEWFSVlxJRGZmqJbO8177pH0vOsyRAWQzepOCy0D6dY2GW4YF
kAr4fLo3z9xXzY2doWTcKUoZr6o5RoQpGC6yGoEtQfs1N7xWAiTDDJGkmR/hmQPc
GPV7Nbj8ldHcWNeJj1Pmz6snBCFt5CGYwvB5PeW2IGCkVbxpTSpgFh89cICAuOx/
AD5ouPDBRJq2STsiXFqF6Ex5TSZTJCzXgc4Jekm91hxnlBRIgxZEMYvQJbC2dGeo
xULECRInVddZYM9ci5rNW8bcw24ZyQejQQBFX10RyREymkl8fPPZe8qVgBE4nsok
PTMdDTKQy7MPe1vs5R4xqRJ/fzQrPFB5YC69XPYTyIgKLssEufriZKCbItqQkRZu
fd5wAph2JW7dboAWbo4rIo5lY4rQ1sr6dQQSMsvWiLotDIPYfIJlBkFtbTQD43G+
M1VE9jiLDALV7fxMdzGVWrIkKkwjdPXP2SbM1sViCeKNEIB8u0BetbLuqQ0gMAAv
BhH4L4SL7jemJ6MliQvwZRGvBwikxT8flGC8Upy2oWMrKZlhchNfYuHAB3B4SdOt
9sU1N9dXl7SF9vQ0Rs4qIA7ZRytRYAunuqf0reAmKTPmCNICtQ2VV1kAU/UTNs8j
ybxA3mepkohJ77TEk+knuRRtnblH1UI7XoAiDJyJLXxJ2xthbwugSVwrzhYikRYg
VdGTTOsQzSCpQDuii6tG8Y5JADH5tpVluw0YRY+aMPHTIJj/mwDuNa21m0W9U3tl
9YPcwn28iUBhwbydF4eO+DACv+tKno7WzZtsYMGnFu/e3Kwy6DtuzxpffTgINI/R
korTgFZhTRIUmIVg67k122yzA6HTvOZFl9Jt6tLBQl6aYBhK3VX8pLRzE/aGBeU7
7kWAb83ChB8N9kK5oalJooAbI0D1OmMPWpkklRXtxUdj+SyKKfkj01oNoNNzy21o
YYsUfjZDHxBT81wwIX02uQIkCv0j7POt7x1KrrPm5iu1LUt2qZBEd49AuWCOuqNr
2dcQvcCy5AY0VGO5/mUUEkuRpbRTlm62k+tQp9sNNrffuxvgsD+NOZnBB9bu4Bh2
UsoYXbFqN4ngddO9F+idjydwJqto8gqx1qnfR5nAT3O9aFVEigpAebQk3SX7cnBv
pAdxmodDjrZD2krKmRtS4Ea3NG3Elygnto04e8Ru8j2jqnijfch5L6W7FK04W4Ap
MVYEx68ZIePLww/LXQqJrW5oQigrJGMOiUFrtrWAvK4VGJQ5sdY9Ggl/SPw4qa0i
ZjBJSMzpQBXhNaytFwUaHdyUDTS7zbd5MMaNEptSouziXbunRORPt7hM3TINWHZJ
YUhuhQfHt6FGLN+CQnlOvvFEGJUS1GoQOBJVsg1yNP9Ha7tjm8NhtstdVtFRTYf2
88XaIR6/Ge+IK3R/6lhxeHOosh2Rqd/mvBPTm4PHaqw9Zeig8or+w0TnXIXI464B
gsuSSW1C4wZJY6+FCPenOKWdU/0kZLlVH/HapD79vk7a8sHY6+5F0Iy84TVe21Tp
2MeQtgBqOAmvoeLtKdnXEyVD43OIOXr3DVyy7/e9sUDqcl3sTGuHp/yylm+pVj2u
o3GuIP/Wrvc1q349MfXXUWWwo20Rgn4QBtaN41YGaYs+LW56sf8lzLexEFIByVVf
qPkYDDKATDg+yAdV9LzrSOPsYm1/EGyP8fJwJ0i5u8DZRjUStvmc8NqAKaoUTSNv
YP3s7fg8ZSTg5cJP3kAqyeGWqnnCiKEuOlaLGboN2jF9TQA1M6ljBcY3NziVW5hJ
wQlH8iNpwz+I8FQq6rQPDQ7wJXVfuqMrLPuAqEI2zborE4CioqLOA3fH4hH997Or
2pRSFWsaobahZwQ7rQ4QhrXldkPsWkEyOnxioC4H7QwP8NhqT3FwuOZK2nUjSkgj
o+wgQYn3gtl9O4tSmTLOU1ig2rj819lOJfHWYZwOduZSUUBtgiQo8XY7YBNXXyH+
36nZhqpvEmoRrfLYUq2Zy9PTP4R8MdNcEQUFBN6W0mYp4n1t2yeYgExiqgDDrNw1
LNR5RzosZ7bmzFwkj8SkfEfSIWzjN2lrfPh6jrbk+fxoNc+JHTczlag6fEmF/d3H
7YL8XxgN2WnvY9hqEkSaG596si/Kw0cs7Aau5dxH8hK5w+Bx0QzxWBmqKhBt8BWn
3WBnAVuYy2e6PZoRYm1HcRbrt/R6FJ94MGrwBNX6o51YDjjkly5nlhoc6Ucgfw4k
MdXn4FFxPLqqBFLZ3DCSQykKWCFfQ7vH2YrgCvmykCto1oHrpbqJeAr2dubzvkVU
5jKEahBxi9jEx6THGE6VmSyivXBzfuBJDHOCymsPbel/djKsP4E7DLg5ro6YarYd
6lJzFbQgVf7fbxV4y3BeFq6bu6KItrRx2lOEgH3Jdsafp53wTSK1abgO4mWkdIQC
HOSv41aeXjnhFHpVmoBm0MWu7/i7D6gPCzv5pvrI+b1rzeu2VBV2EQ6lAlE/LJ1n
z//uxSg/iuzHlLAGsmrASPo3iTQ3PfgI9021vLY622KW33S7DzRRK1+hKlQFxMZi
ovQEyR51WzdbX/w9gXTsfHpXN/qROUCs/bRSjdp7rSTjDGeR/0I+uDrsoQlbw294
/p8yUHI+kABOBUUSyxN1UCmmVI30AioROHrn9qG+6P6KGJBFwoKzXFIEeCyLyaCW
afNizBjT2SLns575KVr39r5j+IZVfWcLMWrPamzZWxf4RaTuTgyGOZewouB4jVS8
OyyMTQdCXgvJsj9kQhNekf2aZUzeGsdicu/KLM+3Ia/5d7vHhCWKwX73JMe3YE0c
S46hZvIbgx5mHMi2l0kQ3du5UfOgrqo7x8ptwbHMsCh1kdW3yOJN0KEzkiPnksI4
sZG1/4ck/D34BOxVDU1yDF7Hp+19yd45difhCYGPtjLtZTo7TYZBndRNFZtFiCEL
QeScoKRVhrLk0BQp+9tPfQ8NNKMGs7qCdgTyg4poD6G8SFxuYFC+gI7io0JSDMjr
lX4gRLY4io6Q2/B+AkzePvdU3PeUr/aYeJ48jKTfIMU3GDzEi4f2ETvdMp7nhd9A
7KWd09/i/wNFStsZNyLIXCQ3NZbh3mnuIAVxMQaM5lK/tJgmBD2TDxNMAK738EQr
7roAQDukEpsFsClL5cQaBLsRubtzILIVKGwCFCSfw9/fBC5XixtwiMuv9TAVZFfs
G1ZBx1nKz0Mtu5ASgrHt0KtGhhVdPEFLIu+5Hkhx5Tey672b+DCYzKIn7Cab1BMp
Z3DoBecj3JjQTBsB0E2+Wtqq1fHe7fBGZ1EoayyRE5nfk7jlPU5aqaPg42yfkGS6
Cq9dAbPp1umsTOmW2vXGVEuMjXG2X1lD6rgaRez9C9l0cHiHPPmKe3ML9Afb4dvp
iDku0snpA4ElZoygm0CwqefQuC1tICKFXzvQ54v1KwU+CyLllRsmBgqwCcjbh9na
LRxRp5Zk8Awx0ZBGnRstPlP6VjZjdUm2mHvyAMSQOkS76awCjfTbws+710VpjUgz
bzgOxzJbU33p2THYqUzUgrJAKeBD7RGbUDywNSacPJAMSBIlRBynNWaao8PaUNI6
UI/AOrfh8SIF3l4CELKOTsFE1CZoD+6EAs7FNlg/siyn/qMl9Jt5WVKsRmcpgZb4
3m3t2aDauPntMhIxBvx5PxV1Tlp24QDczGQkl3IbIGv8UW4/kOYZEsvjmM0DYQRP
EA9znPul+m+ldw5Sg6wRy8nUPMDPm1w8ZhUV6frQAbnqZRI2mCoVl2unGvZPFoPw
qUC4gu0SZt8rLepDttCIBEtcpXsr7OMUzsc7gGVCxHCV1T6YPSpc16O+0wPOZWUg
WVmhSPhoAYHPX/oabTMWSvIwsgYtzS7h0LzMdwHB9EkbSWHSSGbL+Ix9KpOI2FaW
SPTEzmLVDxGZUQ81G2cP+E5ulVgG+dAczOydzHV/xK+KVil4bZEZEUOMYv2X40XX
9xkCHKC389WpBKQKbjylwA/b/nPB9u4+V36QP8fePHruNS7wGj2ENu5LAGoKANaE
AkseGtkaXKeudQzyJIIDUtdOSmIL3hfzs40O7d+eGjDvjQ5qNCkbN4AaKLJdg0sY
DBtTbNeEKiG40P/YmC0cRv9SEvKZ38VR2dLeC9QgFTE/DtuqN6JythKa0HzOEw+B
gATdrYp0Kip6RVY1LJbanqTifyTX5bIZ+UFqrjqF13lQfVNCV6y+29umqvSSoo8w
BcYLWYJwpWi81M8IL6mh4KlCOxmVs5QcNw01sWIvDxMTING/7MZkoR4iFWCeltjL
Luw5jv68oucMVxT7kSIg3JEt0uEIVm3QyG/gCHTGmv8G56Bf+hP3UHAFYJtzRHWh
1R6LqZZaJRmBFL/pvLS+LmBqqZAB70ubFxhnQIaVIJOG40uFhHSAkWQlsxrqgv7Q
C6xIvQN30cCzMeyVKvGJdPNBrF5/FiQQXdPaI5GHcchIX3gnQ2LXBEh5UHVcSqtr
NQ92AYmDKC/s1GBaHOwY84IcJM0EmEUOBVgN6LuDgLd07peeP8fX8XPzI+2SCugf
qC7X8F+Kpi8Wt8MdTeiHOE1bdNtdWwgu0IqzzkY/0J35tCqQUJCrEIOevvkI3UxX
MsnfmMMZP/USVW96+EX2HhAO4v6AF8Qk+hNNY8AAaQ/U9bFkD7MYc7H96APL1IdL
U8yWjaOVqQ6degaokysAd3uK4uRQnmsFhFSJ3qZ5K1UcM4YJln0qJV6mxRi8LKMv
zHdYOOb82XqIVcD6nCoNDaCsyixLJXHLwOAwM7zEnhT2SOusu8Pef9xpSSPh+B5O
uk6TE3ePu/lk+kWEjJXAnm0zPdc4rDcPfQKIYkK8/JP/WLq3BdTIOcFhL2h01Tvw
hiabF6FqoMmDxZcElbPXOWv6HFTE5ke5m187+pANyVE73ZthwnDrESEfT+kuclll
tX/7qRlxcpaFVmnYhc/s5SehYO/N3Bf3lKF8e1P8Vsu1EzYRR3vINBzxcZ9GEiNQ
semdMhHd2hWcBDbNY6moQCECWD6KqzbvKvIJzqARXxusUnRf3h2pNfy4E26NuXot
ElWrpu2cDHg7hH83jRLpDjba9lz5LP5SiceD+nQNHpq5GdhOZGgf76IeLWPp0u3r
Z4gV0JF2gZ54/NhsLPqaUqmFG8Rqh0UR272M4tu9xxoFMCJglEcuDX/N1p9+s6OH
TYMOySargneh8ji0T6FA05ct6rTtuuGo+mYVWafMOVnAJbNX7X839Pk4BsA92W9Y
hCKtI0xegyAbVKUUq3MdRML/lya3zPLGnUG1iQdktWMuQ3lSDBCSKFO1WuG6Pg2R
pavKy6Bo74dicWWSB+xJcSg06EUjuEfb6Q58gGooe/1Yh9oFMzLqtUKOaPrWDV75
LJrB75nUNzWFmpWY6SiHKJfEWKdQQk2VwfihFIsL6ByLYIkpeZtldm6p6r7hS6Jz
Aadnz3KHkvftnil2pCKqqN2KHan3gRVb9QL/ugJxZBl/MXNlAVA4+hQQvTX1dyD+
k8o/lcMnSRqpe6w2WOgIr6iusq7/7YIAI2q27B0upntrJmXX7OG4mAGrEUhJSqTM
i9zZCh7FJ1kx0x/AuxWkBBij12IFfnBXnthnAsDK/+Aei2xbnsOx6Q5l0AFScdVs
Za9r6SWHFzqCnJWuzD1HobfjH8NkQk5A7wK1EArQkt7kCc80EK/MlAs8/l3M3Oiq
h773HODAfj6pShVHJUes8wEvcw15ptdpc+wORY3NO6NQMSrYrdaFFmSRAw2PLxDr
PjD5jNQsyTUN07VWoaycHp/x0zq0DDiO30HDJsa1fyH2dFE5DWQsLH0E3cKxAgZv
EOZTMITIw6L4LH3ERDt/8O6G9BcPS6WRX4VRg4289eYBHbrSsrOSmVVGIEVy/GOh
mRKh3UcwAOcmYAIkislIhlJMxotr73KeosDmRxSHvI28TFFMW4q4PiNbgvD0bWwk
0GFj3FDexk3cwv8HAGEMCXlpHLp5zK+m4mra28KMFI1bbjA1m9eH0k+9CYVfOIy/
KmPPL/oPt6bDF4kkjYfYmNC5DSIQigKTMUHryFzlK58AD7FQ5GSSoyJbFoSoiYOa
Nf1/PjkaSVsgzrls73KtJpxXp8Yp8Gs5nXMlZRyvBNUIp9hqzMGu3guMJgRPmUcu
K1ZXYEzukagZC01NpByfj7/H89+R/npKIqUl6LxUTE5JuW09KD1jJPQvqy3Rgjrg
HgJbvdRLI6neEeARLHnGuXELl8jI6XnhMaPUpm18fLYBvjR7iPatvbsX0HHiUuxz
FvhH2vdFke5YZMWNpX4bLi8m8xFHlKeVT6WTrsL84Df39b4FSTWX8oisq8Kys9vw
rr6ONJKrnekCe9kag/8dUJWDfnt77PHIiuwMtjovjn+KNhldpvoq5Ww71Xr5meNf
3KbrI3rqglikuI+behUZkI8iN6s7qkGxW0YiqupIXajujLJPcIE7RpqDJq8PiAwX
Jj+lqP3KaFL6RBgLN8mKee22nWS5GMPYXyiUjUsyML9lA6tI+pvIrDSKwTkNrnU1
gfmDa3ynTy/EMBj58lyZ0Nn3OUQs641Mlsjrj+4GmOFtTErThpKglU34023qIvas
Gldim83y1scSHDZ9GIVPwpnlqaigh+wRiYuksB4oKFSoaWR9eejgyeNh01NA5kSU
DhQ4ZGlFPqk1hpCCCPZ3EjJ54L/HFRJm+7ZaxdR2c0bARet8k5//nR6/R/L8TCXA
ZNwJouJb8QV4aDQkGw3xOTEC9FXiIoV3uYjnOn9drA1owG2Z6Pkc41o/5YIFzaGS
k53Wt9NGF6D4GenQ3ER2kquW3MWMVU/t3tdv8eQ+Hl4SvE2tKse8w40dhzw/ST61
aQrFzi/wRSlryxd53K3fM1fdSkgT6NfyAaOKGxmX8iyxHceurf12LWa1fbxQd3BA
UoqTx9hV313a+/8hIzZvFo8CD95YPmiRSp7Dw6dlXKP+HLHEHHcPscImgdy8v7FS
ovBSMpFhoqttHwDfGl1zk+AI2NLkkejY1KeejFQ9dKVqNdvHA1PY68CuTYAttYzQ
tvlvDh0F8cj97cVlVyDPejv/GYufXAL8oQJ7WhrCFdGJZzWIK8VQ4iXaJb5lCE+V
VJ3zQew0Mglv0xvTPdNd3AQSVFEXJ14AUvAqRQv8y6Vsra68Imn0cvqLMobrkuP8
BSv+phg8HXp5RAmicIIsTJ6r9/QMfi2uDXpcNFykA7bpZW9oaESodFlcf3UhSf2G
Aow0u0KXHzxl30yIn9G5eAzY4mRPNd1UPLjfagX3nleBmAldxxGpQ+9uLzvATVn4
qoUXypaKTqqEGl6uhjZJC2IIhyv+Fj9qUhn9K0Fw274rv4p3NPLCpvl8Tjm6b1m2
p1z93UJPicpnrv1sDy1E1Fx7aS48wbl+ycd+W5n1I4Me/lOAv2yuVtz/rmzqb1g0
yaWC0fPjHOhreVPqz8zec0ccX7KDQYzFWuoaSkZTUwAxo1rdt8COOt+AX2XDDlLm
XbG6wLnuVNNEPgETaM/Pa/MWSJDTB1zU+bnKHmW34MBprecrqkzBHxMNBxN6710U
04TN6EbU05nJ8AcZbOT9k4pgcVZ+i0K/6sLwibfZ4CUqIfdSm11GKX0nchSUUdnU
V0ScA+rgdtxiCx3oWtZngZg5ZD4e113nRl69wXfzUO3XYwubVHN8S9oBx0FPNKic
skjuBiJ8/oMy3iF94c6obtA1P4J2bKCaBbPGdo5NtKYF2GG9pVzlKU+RSNVdSASU
gx2/hU3a0CAZuiZQXXs2VZWdA9jJ9pODOJMfZVyc5Sy9m0i/qIeSHguLfGPe7OGW
24iZBkjo9Kkqqq6pd/4iCtPbmd1k2w8TdeQt/zg7cYZZKhwCAA7V7sliOpViVpcm
pdpRVF2lu2HpeQhADODiLPc5NonvZBVU1H7/ycxv4E23jbs1uM9KFUlI4yq7xBoe
Axde7rorvVyi73p86PBMbOrqePN7ssTAOEJOF11x46rSGUc/+vcGogj0A8zmqy2O
VrJeT9sMJ2WlI2FzxWD/AgjUivfe2+c4W7L25q+/krp9II37K02S1xjcZ6kP276k
1o3rxBxSCG75zRaKKIcdVpFUjNHzllBlf06IxgIhd3V87tMgwLheL6DDiYsJA6gk
hTu15RKtfUpCxr8SmGP1UhL9vJKdkpN3qHwdINP3LJfxaOTwRB55z+ImdGFI9IzC
wcGXcvIDA8IvtBWNpOt8fmNEk8CtRMQbC7NmO+lAzy7es4uaP2aGtiPxe15sZPzl
TXrOmZqbPH5/QHDJpDyCLNAoeMpMtQlNfAJX2CqHiM7wwZtwihujolsV/TnhTonF
MCFmjn9q/gyuOcH2T68RSavn5KAJEk55dTvt/y2nSGezrQ1I2XJZb53mf+YLU/vz
UwUM++JDjpQTWHjLaUzDg5UdmYzO9RClG9Y7ZBj7BSOYC9ChQxsQyJ74SC8aESBp
aUZrvKr/UayGr48/TxEGWkewEuybWpV/8+alOxiG2xj0trKwAbgghfAdAmwliEzb
TyCJgXJ+NQxbDg5WPfDV9qvWBwEd8qGrJNurzvjNoI59qfQKEKyWNCqSZ5Qnlasm
i9JE54QQYgMcBHn4K25jpKGkoXrzTrK5mcpSGplZE4sB+ZZFxkV2+gkYwgJiLC7w
KvPBYUxrkUW7LE3aHIQzSjR7BVdveIoQiHVbHsVKbtu0dmGPX85oBkHk7iPRqMfb
f+VuKyvo+i0YBRDz1jZ9ptfEbynfnXXAT+ET1fqzxq7lfGpTiwToFPp73MMTEYxX
vTJTnRGELwCVpWdm95RLNikwmkxFBt0pyVBZC5QBeMF2RTYWYbqjqwi6KlqM34kF
RYQWzAyFk0GGsIzIspycjeb8mWXISRzUSG9xLxytgI6qJcv7ohzzfHx/7u3g7lwv
jsU2mlFl5DZQHHeGEZm6y6Ypo5r7lPVthlvwFzipm8lFOapNbVmXwD+LrKelqIAu
397h2ZiCLdjS5X1zoSqzMa6BAEYhnmzI77lHG4RBgbClFbCQK+f8pD/14seJVqqX
zRq/ohZG65VoYO1TYUpfDrzGZkibTFdQ18sMwoqMvVhyOk51vVsG2y2v94/bDr6+
8Tm7uPhs94Ntfe7dgTr35d+/RdMHoQK7vT+OnVcJ8sWCECIphVvyGeVcBVsieYeo
/P7p+zHSmYCBKVyyOwjUQwJ4cnbUtYJ6jv0vniM1GHYFRr+ZliXW8HD6686JeT2I
DLtLAhm5e0D+fsau8T/Jq/iBhpAOmkajJeb+o6/2PhqyZy5XNxRGjHm8VwTRZ3xZ
cWec9eVBeyJ3iGq/zZaN7i+FJletR0FBWSF7gIqKrFU+FK7jIVorGBPq63cx7IUZ
Oghm1aV/qonfUa6QsY/eTCECFreo+L5JakSy4UBJiLEEz/360bAtRpXvzipu0wmI
gtpdmP2At+oIHPAAoMj4JIBJuiHQftNrneUv3UmGgcC99CVLFLe1qY821PvYflxV
4SPXrr9/bS/2PRmqlWbnJBDWqAPBPicBnxaTWYfdvWTZJIgtIN0l1r2RJapxkFPw
ab+ERx7nb7BjOhZy212p24nk1dvOXWUMA5rtKXqtlS7KvdrpLb6uCkyhPKWgV/JV
b4UV3T6vTjtZV69B/XI2bIsFAOT+k4fUe2Ds09f+mki7WcsGREbl33TW6MTrH2RI
8th/6T4rsBf/oV1wzS8r7v7tt2UFLSh6b6sb7YtCgavugcgn+t7ULWkTmuo90bxZ
37qZzwUj518GzwLszfkk07hhETXVinXq//slyw+c3gaJIcmLUsnLsoQu0hWAYtoZ
KoqN2YCWBNaFrTDVma5ayb+gNBJ2PthHenfnSWZLvCLP4dZgHQ9YU2ZHVNM91tRQ
x7oLYFiTkOqDnCDL5p2kWz0RafmkGUr81PUhN9oyqMuRYZs57q4LuRJu3bA70pTc
uvStaQyjL0VqTknZEbAA3S400mR0OFwgc8ndJXce6rkiJSJLCgOU4OXfZ/rLMKTz
pWp6JEr+0Gu5rIxM06AdwzSlQrEtaqQEQsCCABlRSEb0ap832uG/Z9ov5CqoBrSq
406M8G8Im6H31sECT6FZRxO/DHlwcKg4ej7zRz3WFItII2xY/fT/qPq32Lc2/78t
29lc8mXoDKEUhQO5yYerdgxGmbnMf1+h6lr1aFE1oxKf7prWRIcRWX2JjPJ+WZSC
Ye4jKRBElGqjBOBFCu1M7ZHuMv3q5m9SLD0QaxMcYv6giJbh9fCdfVFm3VNheN8Z
wYQNGPgNx+GlHarzxD0jkwwhsRdcib1SOjsHrhF0XsTSgoDzabfovcvWwGsBSMvO
4hr3o7b8TwtEL8km/+kGvTonqrGX/G2dAkSClIvZa88LsQsN3CNVBBZz9WWQrrU3
FeW/KSCDx4kP3tNw3Y9A1fqhF2cvPsMyW+eY6cvkKpk5XgxbEMgFMpB25xwVKcS5
71fqoDQkIjkzrOZOLixN3OaL7caIJW+A0s1NS9cFHGFOIOARM9uLzfSC9E9AjZUL
nYUdTye90bTh5QyY7el7SYdic8LzvIMQqqFvKoHuudufD0YA3Fcg3kHZ9RWbu9CJ
UChLYdwMG+pk5gdLY0JnLA3c6acijDdCvSCfnReQOg6OXFOXXkDTGcCC5h+Yo+49
qanXQpVvRylXt6+bJcUQRL3JIHA5nn7d8zibsqVzfKMGQHvjsrHgTOezu6WdQDnj
TsGHP13EfjPVX5+mQVX4ZpjMOT4ZrBcdbiny1Cwn3pmJLUgQkdddPm5NjLUAkl9P
LA828nh3TwJNYQwkFFW8hYo9YKYGtYFTSd3hj+Z1VU6cax/anUIZCtzbU/w4L32W
rzBTo0L8KvaQhShx66alTvONe1/UOeVRY+q10YXPqSfUYMPM7AhWzZcbMrwtVi/g
rLauvMtmy3tzb+Zc8Jbq/wG6YABEW7zmOgddxIHhay3AtLoQkH/khyskOHHknEyG
dEPFaAYNh/bVR3nt4F0K8FdezfeYbxWIIpff2uBOZPQhePxsFpPv/e0SnDAxoLDk
dyXk9ts/7WEzfNMheu7ODMn4Wd0jn93kXAgqesCJM+dDyxEU/iRCQpU/2YhlKvFt
K/w6vvntiGcbIcL0EEBw+LWPWhtGd4N/8VBWD6fAcmxjOY/8hEe11hys1n75N92J
wsQnQK8Wl5dx/xl9TuldPZ9iNIxAoCXZS+uZUYe9UHHf5xj7LyqG+VdnS+qIKDnO
0GJEP3HWrnQoEvKuIOx/kDmUMHyIIWlSIgC02iiMUAfP0wHmK5UmbZSY813xi09i
kLl0QY7lkIOpu/818XhYXO9fwy5ESRIfsb+iWfybfZ6oeHfg+/Ct5o8nmdMZ+XFV
/RyCW0VJgJ/P8uId+r4tSrOx8arNoq0dwMqb0KOK/YcGzSXkGszYX9jFN4ls2wWR
P6Wg3Z0hRZptOQu6mPbeLVehtVIFfxCMgtJ84lAOTYylJtb+Eq+wZIAbyUR+koyv
y+4uGcH7SFpv2mU4+Gk7Qf1ng4GbkLU+F9oc/4Dht9k11qs7Q4R4F2QL0ug/BHUQ
KXrx3rLI14McGITLIwbnH09bZLDjyrxoWV6PnfUdGrez9MqETBoODom/mdDejb4B
HQF+SUhjmggSX1d7d+QYZ+EnYuTRZ4D5km9w1Mko23ILnQnhuBR1QYobFfVby/El
MxpnyvxiDh+WDm6w6Ldfz5+nrw/YLkhxv23xftqZJ0RmQy6dc+8w8D/Q2dsKeXL6
1+yN1BbA2yy2uDTfGUPsERy60/XXZJ6QdZMrPx1Y7fVjESIIC6h6wUUJNjdp8rrG
fN9Ru+nx/UfjbW9EFlo73POWfcrntpZL7HOHYyDhGcf5Z8NPBrlNLMSgoI08/fEL
UVULXgKdIG91PLpZy4NFDvszPo5o4urq7BPxdBJbKfj5xc247Hy3tJYt2VljCLFy
6CJv+KBMrvM8CxQjIsfTBXlfBk4jYJWYcSTool0JgBc6HSTa+7jWtyoIDzOBqb16
SHiioK5ZNsaQJkW9twf1HmvG7OA8CE/z5qyODI+2BKacyvdZ7Y6x/Omhpma3OeNO
vTDTBVTDpSP6ZCjEd/spW8UHdQT/yeW/COHZuFMBjKZwJwjv/K7ULo21XwG7N2ir
8j5kPT5l77O895RbCJSkXPTzL7OLKdI3SDxlh7Mlmn8Y4nzTN+ZqUW8poxJS1Vsf
ebu3ATmmJs8EHo1AdIo7YDCiVfaacy+WqJe9bGjFGxfp7Ah/wR0TBrAWzb1BoAs5
vKrScP1d0JfhXaKbokRyv6+Cz3z0XcOnnfMYhmdQGQTa5B1ggapdZsHzsGTc/5/7
NztvHGioD3q0MUA/d07m3MTmkw9gBBs80PUy8VsiK7umzVrdNKKDsCLfsO9ULDTo
zHs0c61nlhK8JHYuu0v+JvSu5aNlejgCsZ05Y1QaRtjRMd2rsJFxyUniRH2zKIRJ
Puq0yOpQQiGV2VziszEtweh/HrPGIdJSGo5u+5rA6lg9AjKBNeu9jKg2rs24I9Tz
woiUI3qUwZ0Og0vRF8xbTiqWQ6mS98CIcv0gCKBv7OvqdwAopVWo9S9n36Q1do0A
tOe3oBktGJUbMqtMGQd82v4S7u4L8vbURWUeMfIu7O4NeVlDE1jM5F0JkOHrFhW4
grWW4aJi4R8bG1T4nXKw++J+nbt0uTWL3jpuUTTz/raSy0d7IsZFP2dD8n5DO+Tf
qotBrR5w+Erar+1FQoYbkkZHSdWsPrYTkmA1zI8fX2cSY9PWj62/y4pVpoOcH7ox
l/n0ZlU+EPPKiPPFvUmx3dnu2jodN+iFk3kQgdcijRiJnDA8lXadDYtnG0pd2FAF
X6T988PRvNxg6BXjcKU1USNt2cAQmfseUTXb2lY/CGQLd6wikcEZLFWBjhypvIJf
JgsRqpnto8lVU0LzroKjDK08t5765mZhnBKsNJv98PvsFMsvSsPi/EHlOLqlQpDi
RiAYqP5h/HLMtfY28GwTtC7GlLrE+q25NWqSxKo23ZCsZRRCMnciK1zWVWQkLAop
nbeUqGwNbHmvaG4H7oxRE7A1K05+dUeElCrW+9pKy+iTrhMGjWFeUdzUYAL4HW0A
xMbvZC+8OtqHQvBcGKKgtf3WKKvhfTksyRVJNIvAgkoF6Q58qGk8vmT5816Y8J4u
C87jR2+nfkChMYKNa6cHT3OqUPYvct6E33wup8f9tU8GFIUpiHFEKYXBAZte07gC
hw2JV+4b/9rtD67p5lP25XjShmzkP33oQevvDrR6pnT+rnmCemcAzVreqd52RRIE
mQnatEtB/xsycKXZwv6zdVCi7rY8w2pYqkGuF14IF5bitzX/1k6dBP+zNRsV9Wsi
HR+zqit4vLRDakarRCUwHiNItMVpkhYXojZyjY+4dYtWfKI0N5bk1bixSJDxJJ1C
Tf/+gHx/52g2n5yyS/jfbZaMZleZJY6DMaI42gfXLwzOidqrXENmSyBYuxsPCkf6
99HM1ACUC5mkaOx9GLOpNKjgM8gZ0r+kANhYhIJ32/GkjTmhsQ+yb4ZpKU+SpMsg
rUrjh6nmgAca2xWrfk0KaNfICBbLhTn9layeESCfAVeTNsiIN5mQlV/BXLqwLLRC
W+fay4uZO05520RZHGvN5qhypQYbvAevh82CnN57TcDQk+4caC//TOzTdGFfPGN8
Ff1UYLplRSJkFUDaFKphoVVjMmkvCYYqsniMIeRK+WhsHaki2sppp3tq9vr/3qxc
oXtuBgMaWhjpnmSeTFC4jsc38xRv0yeQ4hwjJzBkzo6GJjwEZFRoDABvkyRBTLIi
G5yYNc7oGlBszkvnRHDU/wyOjoo6z+ODsmRryOxA46zmWFP2rER2PEtQmLRCYEZV
aN1fP5W0c0ZiXkYqtlw5xxorWWrIdvWrsn29oV7tL1AQKqbQKNrN9uIMb4Is3h2h
2u01juU/bEUwaTU0Br4SRpwvATnu9QhKv+aBdpbH5SiDGSsaCfPi1GOr3LBejCBK
iBgRMHzUtlABmGjgVqxRYnUsvRJht5hjVHITB4zJJNhiimeoodqxF4NLO6Go7rNF
+Rtu3mDL/XdMHExI1/WOjvBgrIUTooduF+S4f/vAlNyHSxRs0hVMlK6GUkHWbbNn
HqUQmghybdgesfBZ0J1JTDylx/yGsf/41O+JvotltGZfOsjoQ4C3HsFC7XhCM50o
ihTXookWf9SJ0IHGMCUCUKk2qWTvzYt8CpsVhTPbmofGjPn7BoQOGUfgNh8dEYVV
fBbG/XxGsaKsw3zlUTtQYC5TqeihERSvwR327rbhqAgINLTpeZb/l71iYvz/sguC
//rqiICiFdXbP0/k90RH/OHxgVMYnK8NmalLPodVVcOva2sGsjDu9PNsjq+OhLBp
NnX5hyw2L+u+XgiYOL585/l6DGpjgY2fQd/kjHdeAalnz6GHY3U5ukZ9LCSJARFw
3H+kOS0Qi4oowhXUIejpjoWS3ZdrIgYPVWVryfVGa9jOBPQmWKlcpgzrDtwU/sNj
c/b/uFUYD/7JxPO3qW9c2bFLiQIyEZD0l4F+bv38Tekx1oRdZJKEwn6oRkO2nNZQ
ms1eE87WMHyujlGNOW7pX8oDRDDN9iK0qCMIh7mHbzzkD0kwY6ssCQW527lp3+wC
FxTzhMSUWaJhjYK9QDiwpX4wZUODSAgTxUeUAaxUdqbYweQ+qpIXFTyoqfFX910W
m2r/lcvvVhRNwIhG5LXi0Zx8b/l2cQ22CxzzjdCixbEq+zGnmZL2ySazUaP+yENl
ey1UDWQXVvDRf6qWuA8mqrghqOcuaV2hytYWuWznKjfxLBGlCgvQ6p+/WSH5dbV3
SYRlz3nlPoSBZzGly4OeQ1o9X1kgLBrVETH1gykwV/IV+VQh9d7b5hltjjSwHQ4/
1S2sTDEZn8JCbqD9aKkeiMixILV/TJjSIRoKPadT93XXKhEFmNM0HoG6nczy9tHj
/Yr8aojgocwPWq9Lb3EFkatsIXSTvKiUl0RN45x3RA3PhXlSqvJYH5DQ/KQgy0th
NKfK/VO3N4adntQCSMXrF72Wo75iymZAGkc0IM8zf4jsqE5bCuQjR2PxxCBhhagZ
7FFHfweehcqc+0V3M7a+0iUza1l5tFJE4f24PrXt4FVr5MMruqu4CyrgqQzfAIWg
hg9xDOppBD3iEKw8jgGjSCJ0CupgR1XaFHPUB/3Gvk05ls5Owv8MmY+8OWci8hw5
z6aWkUOOil1I4xajO0naH9vdi/EA9FcwYLWQUYTqoyrOEoR4YeE5Z2kNfOIvH2mO
2k25nWLt42CDmPAX8oN0juu4E9zHdDi5JNG6AJkQ+prwM8xdxG+rmYz11+RAYbzX
pTrQY1t0xrRPsGMk2qR2zpI+USN6Hw+5XV4TJ/+fjJy9dekjJCYBNhnpQCy0zxFd
m/Mq/I5IgYDH4z0Ib3IuDJLpFyeZMsdOLPov6JVd+dE4+RMGopMHAlXeujSy8Jxp
ap6farP+L9N/ivw10aQ0Ifw/7MQjZskJvZ1Hee+RMacEQQNN7Ngp5PJsX6sK7jO/
x9EebvCqB7dndBEZ1VXjY41k7eIVqxdceDmVeKy+peiZ+Z1d6/jk5qlhhFksJZxL
Zx+grO16uSBeQIP5bL7wmCQHcqPuCXbSC93lw8amDZPkMTGRmxK2pMiNf1CEktUc
IAtwjqZg4lsRahRqaFn/iGFNOGW8f9nSU2LbiNaEXxURr5QRHZboSOxcMV8fPpVe
RCxSQpY2NvDZCJk/68iykdOU8RtwrOeLW5RO63Mv6PBqvGibw5xnJY3u5B9uJjFK
FTpO/RoerZIIs8Nr+ecFR7yXZCU2xee2X9Ik+4gOulvI1bn+9yY7Ri12p063rLfa
0WzbyZTWrObEJBRCznkZUhQThdiqV/hgp5bRKxfFinQdGcJj+9aShDX64L4u46wo
d1Gr0Awd7PQZFk/3XZ8c10Lhpx3xeUhYMt/uG+VyX5zjfHBdhvaKL886gSudSG4V
zDl/2j3Mp/nKbAw61FRK50N8UNdggLFPlI1s4SJejOb59andc7PzAffS9QgfcT+0
kDSsLOh2GAC/NpuqA2Hnw0ldSp3hj8oegyW0WDS35Dyzp9ySFwaPXVSAtq3WsbPb
9a9Z4aVt7u96X2xQRdeGn81fuXPQfKAid0PJmEv2GrCkHOG4tgc1fV9LCRDoiZu6
AhnEQ41j/k/OSfz4BPgsTpMnCvmKjWfj4h44EpjcjjhgY2nQkrkxJilTqmRfrgmK
YDRd/QMq6otWNI0Atv11fF5CSd8FTlGGhQ3GYFdI/diDQ3Nx39UexBuJcIkM2fvu
UNov57aWc8roTpLQdqGFBDMdBHRhm/Hn24baRcSoGewKPj4cgtRLSUWj7OYRAQAL
ob49dXkucSn75nE7R5fiOLCXqJx/w5MkGmXDvM4e7dUb2I6w0guu6BBTGfxIUMo5
UKVxbxovCux/MhUmwJDHNDoKKl37Kmy6z7AXSB/UxNH30nL/qHWGDaN739pcXnrb
5zhGSmvsKhA/B5fh1QQVkaJDLqKyAulsy3WSultAnVWV4tJ0teDUMUJCTt8R6pqn
3cBv8gMGUJTKAix4JiAiGCBbMxiecXw4JtJQHNs1o3RDUCeeRbgDTIuJL5SXY7OU
6dphtKvZ/bNjmvGTx4un2vOPyatt62JxM4AbsVratf6ky3JSJbUX++uWjpxE2nU7
gZZUi1/5EmDmEsno0CdaqytrFm7+zYnwC40GLOwaj3ugcwM5qbBQMCzKLCu/39Li
eSgCpW7hyZRDTXXChpVtnrRtBjqT8+4ctRAkBWSt5fHS7b8vXiSh2ln5sY7etxv1
hBoa1RHIik+yO2016OaY/vgvXUFJJ1i5PJSZdjo/VeYRnPCnh7jwtJbZeJv7vpFK
/Gw2y4bBd0gB7QwZk5X5zymyKxtlJct1K6jTd8diJKGf6nJ3ar8gDF8pW/9Hnpyz
SgChjdn2Mhv1rmAs/77RjL/HFSuqDeiEjZs/0bYiKzHjAGgkhZNcqkGFOa1PCCAu
U36rblgDw+KznHIfFcBHsA4n2Om+CxiWoBXGZxlg8SooTQsDhGHqDe3GcQVdM5MH
iBcAtCkcg9b0InYJzvlYl/Hj5x2E9ZNV4zcC8e7LQvErM/hkemHOKjC06pKeC36R
wxfxv5fgSpcsD4oW1DxD0rnw4MpDsbSsds8AI7tCAy20OFpIwHJZH39GlIGuyRjl
Ui3fSd4GKZP0eA/0GRB9S82dZkTNK2/P8bktmlAtWHaQrlCv1tFajq5VRNwbsjWr
Aqb4L+b2aw/092C2hn5OJHIk53EjHesc67DSMO6tyXfY1yB95YwureZegYdQ6vyn
MHiMtnlSpAx9ujN90xu1myJFnaCTZn7EyXMGQmMqYNkX1h2IJWrHE2br1ty2Zv+l
n8UTjzS5ilU5nzCk8IMfrkKxhzD2Za7Z1Bol6EJCOkY9j5VVJMonYyuTMVg/46x0
WPCJaq8ygnebhKUwb2D0rJJGAntCECDof35np1CTGrRC5gN+VOu8Q94SZjvEn+c5
d5vcxWr6In64edJqriP69/Qv2UrSCtPuSPd2Yoh8ki2Jrop34uTdG7sPnH6+PmBR
aPkS9PWmgIBlhfLMAP4jYRuEnh1ItKYV5ic79lQwYnlVVls1faC6TQM5un3wbiYa
VpxQu7oQbaBQO3+TGIdYMhij8RD0gXGOfyQrDtzWan56zgXgVwjdeI4+c4WVOqPC
SaKLMpZY6xqyNK3bpamda9aQ2l7/sXn9UKJmgy5avqLwdyxBTWCW37AlYP1vn2w/
9/onYG95wLkrON/itZ0h6nDKcLJfsu89iYrcdHsvegV4QToogIzHhRY2GAuifPMT
gQ5G+A6MD0gJ4Zk26Ywxw0QxOrDDt7v7T48SMYRJGhece2hb+BbFE8ljlmU49rjY
DAg5A/Pg3uFXJrGcMEpAh/JKkgKE7iLqatxu6VzyYs6dyfNbqcIFZ5Vb9W2nSIsH
B4Tb4u9Owwc8GWd+C/1QUB1m3SbBK1XwdRMJTC0M2pXe/RZPYOXncgg6z3AQgWuT
oyqLVvqvZDSul5SWU7cIQjYOO8Lyk04vO0KqB3VlFOosDuM4WHRjOFa2J8r00CYm
XqH5V1c/DPNB6svU1K3qcNVFTxEQSDlToYNVwlAbF1KkiyjiAERe0i21tDaX4FsP
/PfojKLj4pO8dhvT0AEbstIpE7ufXoGJw1ACmKpvFqA6yiPzRwodPUkrgLXlAezk
M7Nw4cmwJZj1n0II/vIpWmD8cTh2OCt3QZUW+OnWQ8t4b1UQBFYhP8cwJstACWsG
CZO7CZOJ/y7rNWQYrgVWCWMTtUdVBZoSBRrzk/Oalote7Lig2IQfKbBIgvbt4jNU
zEg31GzHfDdzqomKP6Y+jJXApS8WJtN62ccGzgGFpGaLenkEE7ttfnMHmVUH/b2D
9YycoxhwopfECZ4Jf5hDOEnD5ByxwJbjKhLtGxgwNdzof82fN+/aXulP4MNix6n8
a7T0zZXlfLfFVwe7Hgm9RWJRrBNCtjIDv/JPHruYe3I2fhW89QkvpJ91ixAk0PPx
UYc97Qt949mRd0tlsHnq8tAevx+sEnJ9/Y0MzMDplbDIw2BhKOC9ilPVtO7PZaVq
xuac5cg/ELTUdv5RinCCcCv5lPLJnYTRjO2f66dif1du0cQKOuPlie31reaFBfnc
zzlwUrOL0vf7FA96zaFnYyZFB6iwnmd7qlFSpW35CcgCLTuTEcbhaZhBFfnU3VLS
tgztR32UGFYuGN4Atp+1Cv1kKRfZqe6Ss2j/Gb+F1UItUwgDRxgTACWqRHCW8RX6
f13kcigYWKhlvRTM424KhB6FEGuvi0yVyFq1UsTU87nCOBNIwzxFpT36diEHjGKk
k8xsHm0uOjG1KAqY3MlpPyARf0cKvK3CcXv32U21veLJt+FMLmo9rP6NDBzu3jRd
bfgYOfkX2obnj5AjEne9da8EW0Qj5rg/2yR3Ey/i8HbR1YJuvuFXgsa2gn+9uYzr
qSjhRjtnNByfPpPj2jGCiguW3wFMu9H6PNUm6XLwIwt+eUa50v1bCD4QlGOSA5F3
eTXiiIg2pilZVSgVP1EKdzc+g8AJsVEM0QqCXxnJhbAbgTLXc314kIs0Mfd9fnAd
v2zwiKFv3XfCGSo4kNu7bstANb96rBTYyCMcjGd9K8RBR7zWG8Xj7z3cSWhv8cxM
BJSGVHOTkdl9oXvdQ9evbo4eCi7Q2he0iGiGaEHcAI1lOD1VX2qRkOlZpDlkoBDp
gU7oLYRoEkaOhnWXoKLf1la7FwhCuHSYkUzIHCabNycEUBSK7xiUQExpol72+R3t
JxL/bMZiPJU5rrSn73eYCzWuMbFMaIGSMou+YlWtnWYTt7GH0aNPCtKb/Eu1e0Qa
fGvxk1qV3a/GI74xJzls/4T7dMlbYjL8/rjUwWetjTSaomL4SPNGmAKiK/2WOsKS
hD6W2eDJyPNYCXBAggWyxcs8U6Xfoq+F4YRcBvemjU3w7xYjgkhnqyndjNc8QQzK
Z4LBhgRF7kcfgM+zJJLDIsihs2u/oW7Y+m8r0Ui1PgdpGEn09dmeekXMeUBo4S4h
P7xdCtHmKRi4kATGCRlNdEAflzqGR/4i12k3HPDPq7Ff4S/+cZ6hV5FEro1kNhEj
A0ct4SIXLubPBVk5DveekIpxJErewftBsjXymVDvO6JbKrVSoj4GrmPzs6Zefyn4
qDfNSC4pXa9it6Ak41CfsnLx9bCsoxhs8sS3Z53g1uifxlZk7DIEsx6hxozzYCcD
FrSfYnspo41Xyr1UQE/N5as/M8TxcWp4TOUL/54O41zGeFI8pCZtx31oYa6Ytg8D
wAlx8ZEtiDm0pGhrWcjImfo0wNEs204W00zpzEQHxbb5KaYBdsW8suPFvV9iAmVh
WlEE1x5/pR+9ya6kPAeCE+S67g4nFkg19+bx/epJ8XgsBPapzkB4N1knXxFZhFfV
HlEcoVe/MGlO46OOz9Vvx0Gk2Loe0gyxcKXgOyHL42AQP6vkAIaesYgTlkMMn1Ic
WBsy3SQVOB97b47H5r+omiK0d+VIZAv0dQnS4lho+5L+Ywwh7DR6oEfj+R5+lZ/o
vp9XSK0InAx6eF1VIXXR5I7ZyfIIFHOxk+mSMitmZxIKVp4LaN0tp9sGSMAd7NgB
ds+ySAiXKJcJmhoRVBjdOJXiEwaVm8NcBqvqkRNhv1As/pSGHlZkOA+W5ZR6aES5
mK3K/5YWg+it1JoSzoie+k8JnmOsZI/xQeIqjtC/GcXDgyC0H7jeKN0bgsNyh1ZS
5zSLAi0aqX+cSy4r5PMGJhCXR72d51G7KKAkM5yAHHnzv6a+2OiAbuL23tnvosNP
eXSe1v2Osv+coRqzZCoLSCDuO9put2RmK/BVo3+RhNf+uHGCfAxp8kZ1fX9CmxVg
FA6ugbKd/nS1DtkhxvmFKQG3kZigFDaIY8lit5AdeIB283hy+Yu8q/WROBqceEK4
nZLFyDOe1xp+AJU60sqw2bNz6Ou5tQw8yY6R6NpaJdGb4L6EQyUu1QfhgrbcuPlB
Ui1v7HrbmCs5/pDafENvJ4GKSpYnJ/wlbWxPgJCUZrlGpyQlUQztDWtbtaQlkyDa
H8eFNXwZwcq9i85eJPuXU8w+q17tgxAm79eHQv7jy7TjlQrea4mCoq0aCnBOmVLa
T/10ywNufuYd/pGORkZfXk34dP2mUyX6AGkjqvRXHS+AlcSPtQmXoi3No1cIFlpK
QbguqYbu1RqVgXkw1nc+AdVhT2fBMVI2DI3yGvlgWrRptntPzgJ2BGxRIgGx7XD3
57h9668qxr9+9AztKVmtWjZoHFU9Llmq4lsZFCFKqR4gQm1JQJ2Np4+lhQesX7Kr
KnvWwR0tr82a3t97kM98bFW8skoM52c9jZSevg7FSeNgGuai8wKqw8DzQxG3XO82
jjibA16MyppAuzlLtpaPuts3/sIXRJHpMO046dRjFzW2+5qJRGNNuDGU+ReTjvq8
eWkKVWtvZESx+36lw3Hqh8S3KUEuk6KRdqRw7Ez8dCMYZy7Rt9zXz4ceH2uXnLM6
FkJpQ4j7Ie8e0YWF9sUSV0cxOP/KUSBrirnM3v+9+BbLIaszNx8gWKomciyl+4K/
5n0ugqSNAu6mlkyWtg7vjg6yIpmHzFxra3pOoyai+XMeeuJBmV4DaBCjk0lSpGQA
xX0lyNCuBx+CYOtf6VH+sF61FiGcZtrL7oEWlCsQTaJni2lJ5WeRSJ0ALBtEaotG
ei5KVi9rElRDAWSBHbx/aLAqDTyPfY1Dswjll1vhT7vZgnCyt2MkrJsFqfFvZwUf
fgXJKNtL3YwSt+lprmZRZQUel5c6PPn0GmPgxd79bGzkcVWZa1ro/q7cT6IXBffr
kZRn4aOQzcbxhfeysM3130NYmicQ1HDm7hoyTxYHbj51NpMae88ymrP8RZqlfY2f
Ojqj7aCBOXueGzu7LyuVr1YKZMRXL7Cm5geQ2mmWsx6xuXLYgUF7Ffa/ir9KYeSO
Zn7dZEAr1bZtHLeguFzmJjEp4nr64tf5rrPgMqP0ae0nfe8ngXYsIwIabqbBvwk2
7+an1+mQqLLPnPJGQgVUEeU9iib3de2cqvmbIbQs46+mGGLMEAofKEaZSjaO7+uF
kN9dy04S77feircI9DgjUQhTjZtCvH9v8eaqdEDSE1RSpwLbeD0ajlpRanXgfwd9
W7Q14CWRIksA1aKkcyuntJcy8EgZbGo2aS2Pwy2eERrqxux157w2lzogHMyDFLcD
c81iTAVaq6bCqRiKTaoPThJ3Xen+hY3IYpx8WtoBQpzREhvulcnvTX9xUDu9rCFX
2aTOYj0bF3o3s0Rl/hKLzdzp3zkkMxhNrjypHgxiSZSoaLmdXg8EC7KM5nzT3okz
Uu/ZjSAEAzAAYtgQVJjmU8QGACgLpreluhLjaygku9i2NkpH3R7uRlpd7ojoLpPj
P3FjrfYWTfZcyQPFf/AS42YEyBA0USNBEflXIwiR5DrwA1C7Nw+tfhbWHJSDh1j2
3jubFxnAI0boavN7W34OUpjoQhOOn3f0TQoUaziqSnM7zZDKlX0HJZ27cafOtNI9
YhlZI/Svid+tLK1BTSzVQ0OMPpoVyS1PmCtQsCOvRyoUQn24S8TFAZyDCuC67kep
l1pY5MAfEvi8D9uL0hOCva0AaQYwNfUozGJ64fL+zRrO0PIrKGScENskMudU/bOk
7HA6gG19U4r6DpVvKqH42Fq7stTAmhf0JCHnBF5ykXnjh+ypUp2ovxO8miet5mJp
WUMHpHKXAXrR2mYpAZ3nISeylSXhIATRCco0WWgNYBJmo4L+yxDxuK6CE+LIVCTK
Rjbz2t5+nQGIHQyZupZB5fncEONasQ7HBr6mXVAPpzOwLC6qxjB/rGupj+wgweqg
DycYDyfNnWjA3HCCrgZpVqW5qiMZ4IK6A8zmFNEvmSuTsWIRAZ7uyRhNnssIMNGD
vDk+I9jaolGsOgxXEt8vnWTqnn7I9wxn8JhA/Twfvicn1hWjA1euXBoqu36qKPVJ
2KKHQMSjCthyMSNbVcf/4mvsFIozI3UIy1Z4b+oCvvCR7kK0XpEl0tVUqSQdaIeI
QYaA1cjJfkLhoL9hsnDesT8gYl9/fRbmXv6+6BLRw33bxrpkgEsGRFzs+Fp0WhEf
gaCtNFwbK5Ayy/GGK8dNKzBMepfDZk/Po/dDcdbmgCHcfOoB1S0gyXHbjurlBoVk
oGC35T0wMuV/+0wme5Kc0PmtlPaRmE7QWhHdFwdr8rzIPZwWw7MoLuoBgVi6TQui
tyCAyG/wKNpVRe/D0Yfj7DrrocKtgtByaHEkzkcV8n9tfQsUzXZzhSZBHXTlD8zy
O1NxeAqhXLSb0EzF0O0IWYmND8wozUluV/VNC4ipckLC22N1dOtAxzOLw55UKVjw
EPRm/qvaxHdGQImY4nhU1LgQm7NZpt7whYdnkvZR1X7x6IB1KyDFuvcJA2uvkgO3
L3M9DHffPbU8cn709rmu37p48GsQ+WZq01whEiedvj/FOfPxmDjyyMs8rvc/WLSr
lRIDtG/ha0/9Vc6SzY7DtlWpVZaMdyEdsHMUBcBwKJBk/9uN6q9upcXs+jBbso9C
n6glDN/jnPA+LNIqmvpIl7MU+lGAro3BLIoHv9zMTQAknHmgz7wJONmP9xFVKjWo
tbiisVsisl1qoF3N2ZtJMdQ2/xAIxi5KLScuapuoi9CGY4+gyU7K3y4IgbDP11D4
ieRmEnrItq+/6CVnmubrFnp50uX9d7Y44IbnnUrSE0q5RwCRF8CFL4t2KcBgWrav
GKASf8ojJbwwIm7vf8DSuAHrcXYyhsBRl3vKQjk6vw7zv07+hpU6XQbyPNzogKSf
/ZJexWt1Oi5reomar+cl19HaJRAHR4L9BfdC6GLshALW6qsFxA30VpHAZs681oQC
GTbnmY4z2sWVSn9dcu/8B1RVxhmsrHYMVNX+5n1E2jSuhHuUJLfzlP6pmMMgNF7t
Q2oxMf31k6UA2FqLV9dj72FOOC63YHDQPkBLRQOlZLRpmtDjvOb4QIdfBOj2Mpg+
YjezFP74nJUf6QiciNebyVvgugCk8lzoH9/2ZDIeo5yyT1lYEOWii1PXt8Vpw6Dk
pG6bp1mB7y1ZciR3B9nCXoUiSmSkTzkWh/Q0y7dOrF4qzU8Lr8K1bV09vJWl6mwO
L/XGyvW1ZjAb2gHh9g0PKLN02hM38/f3mk754ws70Bp57I+f1XIpFOAWntZ5MT6o
zJ4C2xrQeQt1T59MRN/oJUKH4IsaKhFukdRPitCyzuJ4MV/Ei09ezWPZDlx9A/oK
vZNZJRP+CyTO5Pynpid1+1OJx+RQy7q5bT7ALpViAxxPSMwNi720UQM+GEJ4xk63
dEhkFqAOp2qgp9VkNJMP06UJ1yO3CTV9YprdKWMMMJjKomnLJJDpS61KLKzX3O2y
d3Uqw6LpoxlWhxpP3Ql2edIEPCNt1KH0YA0D9b1ObDw67fTIYYMTWVYw7GuUE2J8
7noqSYZs5tusoDuc/ZOc58PR/9lB85+i3q7MskwT8mkgw/6h81dIZO53uvCawe0I
s1N4WO6D+hExZYyOLtTWxjk7Zqu7D0oG1N5NOzF/iJ/A5haBeovAKc0ws2WbyQ/K
LmwJSt3hE+ndlKbQTvhjA0WnypVFkBTMhiXUTziGZ8bPLY6hqfzkLBa9pEASMK0D
YVQOP7MOp9b3VPinUfOt3SfwgrZR2Kr15Vcs5LfnTnyADCso8fGPB5oUDXUO4GF+
dcINU+jlVAOBfW+xcQUFJF5uxJdEGO66kmhoT3Oh/W8KNXGoWDZt36dVugP8fGJr
o3+RaalaLUBKoaHS6bx8ot8kVLB3KRAFJD1op4N40HApi/vue/Dc46YwTlo8OczG
2FkAoBSIsIJR6QJF7E567+Pi9zF4mWK35Rq0ka8bp87fddp0Nzjaq4KOJ/iZDp98
fQaXJo9YHdgW4+1wEd/o71wlVYI99VAKAIsov3KZGrHbaJgMBMIOPfmuMevSlPqn
4LCsL16ArjdrLaIoYIyexnoeT88vSumIMroon8LLJHuJyz5igNnnMsdpfbOkCs7H
lC9tGSWfkQoLrMLbJE4gsG6rIsND3rmHWfJ4ONvD8IspH2MWqU9wdYN2OGpOSRlG
zRW9d08eqlg7yXg6Od0ZJG7veAsHu43FNW/by2kyzNthh8dMQ6Xaba0qgXWHk1GF
LLfYDZpSOLi6xBsdZcaYGIY4fsMeG89vcBEhIzYgtrwcXw1Eivs0iL4fKY4QlPPF
zHrN730w3hMZ8ZTQtf6/wDAQ0Hh2wxWHlihbkYo8xTV7KYEupmueGVGtzp+AQfKU
RqE7oWpnmBnxm4SOQHwuOaqwrjrvfUWKyCg3ejX/+QckCn8wTJMI2DwGTYUKPkiu
lLgBn/86p1hq95x0t0TLzTDhGcQfDRqDKk8onl0SlM2RW+sO0BCPp/RqsFEKPxTp
Y2lv5l2zFn4u/I42Y7J8JrAuS/nPYkZkq+CjYXHhCWil6tXJiHEM06pBS+eHoLjE
Ul8176z043kBbX4pfyK5mtjGw+4/NGQqNsGAmGCPmEam/gSvXVFlbnBjIDN7sVeA
pR5xb8+oMZACmSHdM/zbgg6b6pQGdzsylQtrrb1aMgO2a1BBeePOGLz+/UjQk651
zQmmvj9rZGUXbJaHY+OX1O4EHUmvwKv5i7YK+XrBZlBr4uKjlVQxM9JgLxe13hoh
WRL97DMuSenoPHj31e6af5gixOvgiWbrHD84EFlGyLTYB1pPTlwrdDoRjbypmBbO
0/FV1l3snLRVFaxyTx9dLe73NWiB/Idt3twq3bPcAAKvU5RKN33qy7kYwMt0Sr4B
PaXByrfAwH9E7/ZIEifHv1eGNWj0q3O0U7V1AVyy7DHydMKrERDzEIa02bDFlrCn
uFU2JI57HzHMGSHdCnrFAbLtiwfMqU19WiUyKU8fGQXvrCW2PEk4cEBsuRdO3mwg
RTrwYcar2Md1rZi577Sm+ULV2KTbmAj1B8+5eyMhNQ6g/JeCvSjCvw5EslqWznGP
pRj2lwfcszzvsgJGgJqCwt2NQq4yfczTAzIsHgtqY8UDUaCQjnW+HAWz5HhM4Unf
hTfCyO8isT1f9B1sxHxOX7rBv0eBLsqWDhST/+12tioFzQu+UYSQ1bZi2CSuk3q4
r4mrVzyaD0oKGBowiQBHR6D4xJqKP83gbRgeN7ZZeX2AzC72nWY+K5iGz0Ojcz+w
jOF0yRiYTNbvTrpn0WUlMcllT36+5qT4iX1FtYqvSgcTb4fp3jFe+Hr0agsfYhVf
LDw2AQcBPzPHMrK/Zq6bu+eDYiCvpybBNWe8CTv59oDSnKg1c0uZcvSKi2UKrewQ
yInFejPOWryR2snPhnuJe5htakfW4yUTP3V4y3pjj3z7crUb330WxeJ5dDymQ8Sl
ChN69FUT+r7T/hgdvsOkkb0bi9jKrGVp+HkgGfyMoDtD4lGuHffVNzUPevKPlYM/
3CjH3l7xcOKKONcKZfSJfyvLCAg0+3gE0DEnxYnAw5HppImNdgjF3OBy4wOGr24a
ONIKPJUhCB9CJiWp6BcDezDwBqQBn1hzIT3O9PAkKRj8bNb5npPJ1f6WU5eLx0bl
wAewkC7GyI13JewLs/rkeG6V/bOGOrylaFRGG7HN1Od5/XbOetVpOH9TLjncwUF8
/Zmckqm34ineNkNdCCib+iO68FoiaGCBy6Sa01l+PIr9r5XUv6I/P0YmSOUmWLTy
ZbxFBXALmSyOpoJ2IXP4UaKhbUJTcFpvUqA6YIjQ8V/5Q7AFFBIvGasdRvVCxTnu
lhkj0qaWz8GZIU3m0MRLzmmSRY+STjF52mFEFuR96yCsFKfjkFD25iXHwbzbqAJH
Kgn7+eE5f9M7faEoKw7vmun0fpx5FwSQfqpsrcfxMYTm0oXItTtx38dIH19g9MB0
g3ZhChX/9ErMXmcqrZd2OP5PCrJifown9i1AFL0G3kZlmcD6xL1Wrwf9bF5iZsvI
WoE/6FnLYXXTpEGiKuqcBmQF1AgRNUWccDQdn20TtesrJOpaDJrCOnA9YEuD3VMJ
M+mVAuJj3Ehpa7wPKOaHObnnIXUHan60fSoNMinbKnhA+GID/Cu+vRZqA/K0thHP
08YMmJtl5PxlwIbWDXp0kfCl2gI/uCRLhDxeNVW3WXIT68A761wfS2LxR1LHNZyA
ezf2f34V9UwexdL4NCQVn1QnB/xAPja6X0is7WBeZvoy9rwPa7pjFvC/sLvreKzq
1V4u4HkXSYTl6yb3TBKAMmHlLJ2jPo1ivEvbWI5mUqGvv5pW1m6smHdtH2jVtXly
Z/jCCQ6LcQgk/TNKowPFUOE5IhZFihjhpr9h8BgSPHIA22CQDtSqum+wRbvJu+nx
HU/qurdBNGXhnRnJZB03zSlB5xOI512+iKC0rvBZvu6I8Hbqo/O8aa41iZyUxx9L
NuLSWl6x+815+XVFbUj0RmBCb4WV6IeC+OIOCSEXOd50br641ULvHZQD46oGTBW6
G4t/q95Rp4iQUqN1K166QsMDCCxVaOVx1WsXLhozqIfEFiTfcnGhxbVu0lEyFf4P
4e0Dd3BIVnwN6psDECRAob/WnbI+CiL2swmBUbxISx9fpNtTnwTPPR/wVXsvv+m5
KXwe8jKxm/2iFfgVl75WQbLf3QmSZO9WlcERr2tiR83s4zlo6vMdBmku+rso63Fp
lqsyUDZWF3qGYwl4BMFM0DqpEv/fNTebherIIMmxcZHb+L1ZKmhN7IJwCO2ojl16
ousOqKn4fagwS7nwwBsvhJDMbs3OeaeR0gAfrqXTYCD/yQ3Oq4lkdGXY7LHFLK3w
Lgzy5nNoIMDLqP58qki5B6+eIoeICwKWVNl/fFO/HY7EUj2HONmDjkaeu0CnS8yC
l7uorEZGCxzFRh8TPJqbM9YKvnBSk4fQwJlmWVcGNHMGX1ONXEytllThhcA3ahib
Ib8nrc9OujDX/hcTWgHiwkWBiKsLQbngV17f3nEZKZ+ZvpCkOOlMaNKMSMMEJyWF
xr3cwQdAfLcbfPzCevzENDeepP6Z2+N+CK+nkVMgv0FuS+Yi0ae/zdFWF+tH1aqA
DMNyz0mrwbFKctSB3n4RY3CHLx/fp+X6AdmMtOQfQdW7rpuNbpNplf1IT088C+mU
Qa5Hp/weelfWaW68dm7g7sBVLeMH31qBSV6txCQOQEfd5ckV/4zg5Cu7S3T3sRIe
dKAG0vUoPZd6K5FjCji3zSCZTM16ldmlB3Qu1RiV6vlIaEhoXYb5SfPlwa7eeMLp
I0m5KYxeB+MupMiyCSMAmghE/mao/FDLSzr653IwcY7+wx9IMXe+JG+kC03heBIA
iBuDu25qEiRlHRPO+CQBDz5F7JvpTMoJO3eXVYAafcUEZn4407YNQ+RTy6wv9YUa
ST3QpZm/WIC6GoLgGmncfgr+9ln9u0VmX5mKkZfgSXiMhn33/a5I48KISZv42rPH
RadhPnCvvR5etosvQPhgbw+LSLAGMuhvbZ5mTaSAnqWqek5CI6r5bWM7QtUfdwnM
YKNuL8ubbHa9Y5hKhrAq6d4KUCr4p5dlwSZzhsTCr4onaH2Lvd6WOm+awhsdW3sZ
q191hGxKzNZReBvvGW6IGNAObw6okfZVpxiftXy/bfpO4RrSFqdN/v47i76o9tJh
AvQJzt6XWox9KRCjIneb/Er31lNDxBlh6WGiBgT1MZloearexQ1XbpbSbpEVHDgy
hJSzxQRY7V1PLLcLEGO7nyOtr8QkXQ50GZwj2uLDin7OTw5yHM8iMwgs/RxJuwV0
F8cGJ8rA6/hH3U1yWc0cJqdeQDdkEBYgXGiMobA0jNdVAMn3J0M8PeeTB3DBuvMV
2YCTXMIe4K99IBP/NPxN+3PibZ7dvwb7ncqQo0zGo4F0YeTrkoTqDdXpQ0+/uan9
PyRuI6EhS5V6iMEwLDeW2ozE6KcSpc25BwGoQ7HWJwfYVk3nxjtSiIiD3XpFSE17
nQRvqW8/4ad9zw4OCdUTpzFl2QT7Wnr2wrf5xy4CLeH8yFOcrN2PJ1UjdykBH/Zq
+803TyxpfaJbrCnm9H8H/qTeJ7/HuST8S7MbZ+9mShs0VWGSuawpMbTJvfuPpGP8
0eocvF4JDX4yv7MsWvqWkdJp3kPyHgFSTjMuwk7HGwm0n0EWrxN4XiQ8MqiPkTrT
3snX5wB6AXpsZ2m6yN5xSAD/HFAuK9El5i3lbBndVqQ1jOtOqxmAOeB4g28zamme
weRVJucYkamvFyy8beeR2L7PlwOtefg+m0nwBhSPOUBXpeGuTrKI49Bfj1cE4zeQ
AJUfKyTU0GGInrOK8jlND3MdLJnEYw3/2f4PZiSsAk1sxOJBTiUQjFf/BZ8JbXP6
Kz0/ilaHgcKvBbRHOaScYDq73C0j1d5kJbd0SEaeW/wc0ciCFUsp3kbnqh/vbp4O
rzvCrlaN6MN9JQlYVQGKJ1oKn/8KSUx490ElnS7dmMluTferjopa3yGNZ+y7wIzy
EPApsuAkL45lxJ/tsBhSWuIpZf8cgMI6GztpgUN8J61hCv2vAPrUH+7j73rE/VKD
81xAVYU+W0DdW9c4pyH3F8rW+gYPvYfY4EJQ6dYaHXf8vC9APkKcIF52U7Zh+JY1
ZrDLy4ntrvegqXYir8dKAFRyYCbqryRDOCmVa4FZL8qjHaBocZNXxzeKn5tQQUBC
ywi7EceEBvzYEl4ZuKNXRfDxsqOBZTeH4mJh1x+hvafBW20wOHIBD5jdN/CkFibj
vzxC+UNnCEGHs5agL2tEsqIsSyRJlTHUD5nX2T0ssWC5QqV55re1sQhCCMka9NPT
s3UlB0Rtj0aB6NaqYsZiI2ZEa5KhiJJEoCUNfNo1rb/FoKexToLTu/GnJNubrA5b
aVk46Aat7gEVxF9ffRuYJp2lwgAT+GnVFHC8fdCPPHmobnNAmsh5KIoPTMMktbgD
kmgSSoWMA5lu17JMA5iPY/7asORMFdqFGbSvxymIyTn7xIiNAC8rDl/c4k3vTPG1
S732gbfu6KO/0p94XI05Ct6Q+a9geMQgVPOFY5RKKe3BuRD0j2savmzq2bjIxuEE
fQxE4f2UEVraQqwofZn0siKgiYEc/d4zszSIDWVGx7ORSeYlvNa64tkgW6/FINp4
bxyiHJ8qcocGTABxx88CfCBvbhAyPbTdvq/kJOs7WI/4+uHjuRgzNprUsrT25W8A
hfath4l/BEIOx15UdcBBoPim2HvAZqqbKOw/1F8nvnzB3DBmlVLAL4Og99IGdQii
ZWxoNs0A5rN+cLleJHtyQh9DRa7wO2kOj1OLHL4JXpiz9sf3vKVZWPyhfYZDWhfC
NespIq5sVoohE7EbkF1F2UHKw9SEyNJuRtHH1EsAdgWvMNF+DYyQS1dMAMdEkuDB
Lspn4oyqKbgBy44em+t/0SXoNxjU/m1EXjHzvdtwh4iFpK47KVEmSTte/37oek2p
YGj4m7JaHMAwpA82NKvVRqovIQZUi7ZNTpcVN1tVBU8eEtv53Tl1k+osG/TIdU7q
jeMb5LEH+iz6g7Tk1nC830oM2bu4DEk/hBW69OoMV+4cx0l+RNIzFOdWfhg+02kh
Xb4mkVUM5zdYOMnhgfj2wScofXnT34JiHuhGwU/0nF2IbqgINX1QrDP3KTU9z8LZ
fIDLXT8LunaERDy8HJoT6ul4sH7bTzEOEhgq6Uhh/bJaszSuek7ntP1Dcj97RfGM
yZxiGKa99R1484uHtsFg40eCa4OsTmTNeqpGrpt6DCbxm0EYkjzXlnxLkhQbPhXH
iUDRK23iBkgNtnt2FfKz0Ki7glggii3ZNlVI6kM5p+lhmh6uQSAx0gku1h88k+Js
wzqw6WMENKoKaZAywFZ9JHCgyI/1oZfw7kgRXwXZgMza0BsxrP+FFLApkgWiDRM2
rHn7s5VBUyxsVhSMmyqB/IMQx+/sHoZM26G9H2790Jc71/UF3NMaISCIdAInUHlE
1wwhjbGZqACEWKWpxOHvArVa7c2tQCBWeCh0rvIXJd2cUVmPhSJTM0maj0nS17yQ
A2CvlZ3xA0K125KeqMYfqVVpbkCQZBJG0TWvYrOAeuynZYHJ66Ynnp1J2O5eWm6n
26PemvpIMzSwOuKBsk7uIEyxosB97lvAql6Y1JF92M0FUn44pX1jiHR91/2qZTPM
S7C1zRnqHVX4IVjBbFi6FJbDgWYqxTpisASpdQarMm+4WjUOr4V/e4cqzIT6pqCg
7YMmUYWrlGQVcSB8GLbk+LC1YNOvPrbz6u83f7OwbJDkbk22IUWSXW4hKAr+q67Z
o2ieu4T+jQwwD+5bZ3riaAEkSWEYhAtMj4ecuwGMDAuprhQQjiKOmGOirWaLocaU
fV/hvalDUePX94WKvodU9JQmkhnIDtJ3mNUTpgwsZ47S7x+yQUkvyeFL3JmXMc39
53R99ocCLODj//fQkyFwtZZSBuH+gD6hTVGf1z0g8wLjTJnoHzOKrOfTiW4F2QmS
9ehgNf+9SRfdagQXGluMxcuFAFOr2DI6py78CgEDLmJRAKjUGuj1puHRssb6a9sI
WP9IDvZCXmaNRX5UVAf21+l8TpldEEqJlNPUNC9dtP+BGUR57DXbCaR8oxJsOfTm
hjuUFrRNM4VIe12BvmVDEUEC+r3w1YJBpFyBeGNvlJ+aETC53j7mqb+dmjzfuiAo
JqSn3qxEP1OrDxTqicgz59o7gbl9qJwpkjcWm0CLQUbv2r3be9cb65bD5Sd4tbMV
9z+EulirCMDkv1P8t5zlbItHF/bMlCF6S4Od9v9bI1/OoEb2JcwjfpCcPHuLV89/
Ly8Rb29m2t07Vu75GoAvjDAPS/u79g33oUy41U9lTSxw5suUAyIcA3KSIXbJHrnN
0fhfPaJCuJCaZ32dFuvxv6T6WPt7ZYx5qa+4VR6dcccDnxqDOI052AZlbjYK4jYW
v3GQqFpT9TSlr5iGuMt6aZIeiEPexPL/QWsEi2IZa9lSU37q4RZE9hkTlBttHoKL
IRpO7IlylzF15z52C49yYvwblRuHKr0U2RKaD95o5IckB1360MHpk62niEa8pgFU
8n6fe5oQeGPlnnIyXTRdUnOJH158Kc56tcBYSUJguGOPdu244hdhp9Wj/I9mUiJ0
aYvnR2wMIhTvp6c7jsl0TqZ5+g25lFvCp1Etnh+DqdbVhpJjCsWpBETXpUFu+PJ3
/icS0n/CmhAMj2rAoDkzeE2ZPZ0wpoz2+CnygziVyuoF3REa86qhI0bdREO66Qtr
58yO0u6DXqlDsveUiuC29oU6DqP1oho3wZ2X3kd4lo3jexFvf7ZbCXQ1M0eLSDoy
FcRvSPgKCx4P4D76eUrsBfRKezcDe9rwc5xHPEmOpR4XPybj/+3AO0Cn5PfQ9pYp
KXHBIuxAobBR6xndWNg4pXQxLT1CV6mEb5o/PwA1uGUOKXm16jhJDOPNpQrK82Rj
EU2DXTh9GKZYWn6lDWcA2OLtHnuwUBwj0g5dH7UF/bvFYdiGQkyT70raY3R5m+iT
lUeuM6n+he0GRtS8jPUTs+Eq7INcgvsAxs5VRPtJfOfJk/oPMHQGoFn73OL6RIDO
JdVI9Hj3C4PUXeY8md7ehfoziLqcrAoJZqYoDGbR5lSqxOPWRqvb8FVpTXTw97K6
3FyeaLponmywEzd4Mo+2cXA2T6Yo7xHvdbZTeFHFr7aGwXtzj6MNzSetdTA6XCmS
ChDZtP3azsHXNrAU1ktxr+D6YDNMJFLgJg15Pz78+j7bMi6iPkAddtVULCAhXA2o
RAjLh9aXnBB82DzZxXWHN5H34piYh642UZK8qMTveu95nfLPVMlx57Ex0zHTOR8O
ZDc8LrV1XavitCO+ATdl+a24lFzInYyS6nuSioPZmGEBcN/7EtESgA8hMxdFzdkt
sN8bJdDKIdEZs9wYsEdHwNanuytPZEEkjAOvlhJZ8ihMjjDP6COWriVbbcO231E4
DXs/En5KVwHbnBJBXipbcEjrLOClR4HcxBM9EyTigh22CqhX5gaJ246NbPWGeJUX
HQGz/QmypXiyQXC+xv6K2VltyqsMVkiR+eM5CgSB7vx7CCMVBMP6fRahUAqp2n+1
D4yyGcsdk5pRaEHemiE1iwCHT79oVrn4DhBuxQ77QeVVhgFf6u/dIOz0dZuUioPC
aPhLfuCOME+NzII9Eo1/Vd8HinkCGzVeoYVVyu+1D0P7PMvzG1eEVKuRMQTxFjbE
MGjx51lKl7lPXTWyfRqQkKY51ozWwaj+Rz4O3iKfK7+us81JTT1w9SzSpZrx9K80
Cgstq4ePsMGX+ZaKx8gfH9pQOSNcGcYqHAXEa57Xzne7LPuufOIQ0W2ER5Vp9VRI
fB2cHesvMH0zibcnn/HekZ5CM9fB2pSclS/GnndO5CiP9N+OnzuYoTc6VmS4npju
62Y9nqAjXsY2tNDS/AOlOR5PYLCD/jS66Y+vBjqHiCyQmgX4NaY2Z0wO2ck7k8DM
Io0wiR+swYn6BsmhJvVDr9b0nOLmh1Zj5WX6DwmkMUDoMlCVaNRXbRxZt8TX9DB4
UW9AflVRlPiljcvGAZX+HhBszW/S3NPCL64pgi+h2sVAgoGyXO7Wz7fEtZV6UZgI
hhHYq5FJH8CywYco+le6cT13q9bAR2C4B68OkVelG6N3uAb+c2iPoyVrdTxJ89Bt
fsjpVO2O5LFXbJmapSsaS9RmJ0qnFlTCkrhyr7E7d016yBts+Hfq6ckzN1x47Qj1
Amqj5KL/YiCyvjBfkiCoIwp4Qt0ZfBSZN81zgJDbJS1HUA33eRo+NOsQgBmmCJUO
yN6Y6UrWzSh42ZkPuas5vlnGam8oWwwurW4vgZ2BQJvVrtx+sj+udUumcmMj253X
mtouqYRosREYZ9OZ51vhkZwU8GnplL1/sNMqiyiyfn/fkr2ivhMOFTEepI8T2/U0
Z97GfpRapt0sM4xJ33V2cWOGcZwvza4fi+OhKeeCUvkxdMHsNRQUJNu8LmrLmduV
LfHMDglgUblFLI9QVpxhMA+AGP0ISsjF+yvEIuNPoOJFa2LwyqlqpZu7Cxv46Eiv
HvwDc0EdOebbkuzgv1O5nDq4Jft+jmmrKjuO08R8IJfICabMQa0EDtJ3zu5xKCpd
qcOdMX/9HeNw/G0aejsJAUDvzDT+ml4D+vx2ZirpMj24Odg7W2CPskcmoi0Y4V0w
fby2g6WVvs1l2xC6XJtH0CVwHsEaYR7kDqVpGYkZi44BtheNbHXDvDyAdOyfICDg
794DTgruxz9gxYolwg1RPxSF+T6MLddeat5a7FvSHq8+aMqgzbpmqfIjgSzH4FOa
cnWjWahKcqN+xEPDp/86Dheyautsqr2Uu0DRFcI66hEba+Bpq+GFBY4zIvpfiCBq
B5xRQ5J4sWuhmlLoH3vtO9gf2i//8v9XQIY7jvYLRno0xfmlYy8SaKJUfW6eW1SQ
Lth6okSZBMkUBERAyDCVwuUr8palHE0HxEdcxtFBcPERC5SWVAlutcB/WjlJ7c4t
eKxr9qIrDsGFNSwLpGx7sOvgGaqpasYk9e8BkQ+OgKp5xoAT/6wH9KOZeuA9LUfT
gPRaV56Xcu8ebLc73H5SH84aRqP0LAcdzzDL0LYHlSwBepsldBb6MJ9xgGsJWFr3
gzKWQYswX+u77/gK62+XpvuXh/q/5524XOvosZ0G2yooKZ09ESa1culjRUCxO+m7
UXT1V2C3NrvI/21W5FYQYdV4NmNEwttTf/HLXUbTuJ3P+0L5CYAQ8oE5K8OUsZe7
+xgzTXxxYjrtdRSAH9/0Lxt5PvbkcO6HMsv9JnVYeNhxA8yemo4zxoK+RzdL41nX
i3GCkYJr/sGiy8RqPb4tyIC9aelrmViDIHCjBDdObN7c2PdrnnR+aI6XBoE73Wf+
LS7Zhc9YLKOk6iPOTMj64PfmmKhcxnLR0iE94PWgzRg6zN2pc6bexXwN4YCwhbCL
nyqdZGaClJI7IU052TOGGXgm+TmTsXNiCdwpO0wl5wRyEd3dqNcZ39eMcKAxpkXz
HE67T9ARJvYXVg2QLjYrnqc13UWkg0CO1S4UQGxJx0iSDdzikF6pvXqJdvxvrh5D
NUr9rqxDYUn0FLOnsnKVxYjr2XU0UjiccdYIHwP4OLu/z1HGDns40VB+ixm3fJMm
ay2Nkv3oMvxtFQx+FwhNLy8jhvqV7TSr3NPgKciFHuzvuttAU53aPH/zyxBXpiZV
igaOm+VpmelZ4yiMWrAcxFmQsAHSC+7V8jImBCBNyrjWwEhd7eyP4NPH4X8lsAew
3LqzIM6HCCiDnrWVDswkXuE7zx+QXfneCkA7y9bkW2pfmp0T0xGbmG86oL5HLR6p
sfWCynig0BAI68+t9pvgap5a/u7Nhovyj+ydYOhOye68vj42AsoFM7RDztZg9m2S
yLS/Lf2yKEDV9fNapcruFHMF2rpFw0Zruj55+8wfsAP68+UJBoUpL2KjopUG902Q
ZNhAZGDLkde9kLaKrojKbvDrqU8sUwqgbTQ6LOR/r45fDAptsdYTFaq+ZhWdLR/9
x0Fb3JA4SxlRKzREa4QMUKoJOAFpht+QfD+HH0Y4GPAgPAwtCSaLqCY8ZvsLJ1oc
vtkmmPTnZ1pllsxEGVAl3GhqeDGcjzKT9H4hrGl1+gq/3cCXCGH8t9HidUhncwxB
/jUqumDVRLkNKYp5onM9YWpQW01wqe9r0FeaC5yKyl25Qjd2Tb4Zn8/s5BRzspjO
aB3heNW8g913ihlQb4jnbd4y+tDpgJxpuSDomqob2y9RZ/OTadujOb0ub+rJuIG8
8ZioH6b39S+D5AjBAjjE2JeSmXNxRGqs1CqCF32rqtZ38rhK4m4mmxjX6td7wgKi
W70HWF/Mvvt7VXFVNlsqGZCGvBtYq6NKz/3YhUKxv5P9gLgDIz1PLdfMw3E1FuQg
cI3pJPZcSnYlngqqBc83dFGVOaJLo7qBZ6xPGwBif7pyqQZMBhPL8j+cIn9bsWlw
HGi2kcL0O2DPnLGmos3jxflQgBzqxL/johrzEeLyO1gBD/u22gvFP2En64v4kGpy
db6yS3BuelmEH7mPzU5Rtk8XRgx+UDE0igsns4i0I9C118jhaGfBdvEdKuOxgKIt
Qex6LZdq985z7y1S6IyMzY4LR+MFZqItpJiXuqlwWdY1bozZBYF/iMIE7PWZ9qLd
oSjQMumY2ODimtqf8F0jRvuJFhO7dXOn3wzYWKTLAp3EZi080dVeaJzIZN6qwuu1
EjB5McmKHPIzWYPu53X++q38nE77Wnm5giJ8SaN0xYXpErdKKNs8uouFOPUZ9Mra
AzPgXSJJAarMdUzSfv5EEDa46FzsFILxeh4bGxQaE7PiuP4hQUPHo4xlrU1roEy1
dV3iPN4bJbHkG0kE/veEmKxWm5P7nQn46o9FY242w7eyx3DTkoyO8daSay6nrWN1
32wjQK9Z3mdAh/3am1+do4UhSDGgYuzRqc053u5u8EtNqnhlZ/ONK+O5pVkZTncv
CDb39+IddnSdwPHX296T3L1+GsA5uHlgb3KsEGDlexRoqpiFEENC2C2WEFN/1jOA
qD2ZNdOOCLckHHnkUQck8ANv8FUzB1aqw6M5GjC/ztyVftEpPTR73uBtC2aJajQy
VfhI/1YgzenwWfYzKbHUdDBfUmUHbz8O9FKj11iY4pAWdRDVQDYNeD7TjU0FVQM5
CfwFrY3rgwrBnZOowduuE8p2Wtd2fkVPBRn3gW+Rsfo8+YtdauNovKNgEbNcgBZ3
sLUxjXhaSfL95eQuYYx7gOI7zd21mk4I8IhWZL88jTQOBF7pMmY6zBjzifTKmZvi
ol1e0fXCdji7NIztQ8r8AQ/+FAPN2TPIFvA2x7fwIe0DolbpGLov1rjtBYCEBM8L
A698LIvpwSq8GnANCib3bltIIjT0h3QHTsWS02rPRSIaol+HzNukClRwWLmi+dhQ
53RDIDHwarmzIH/14gNyX+ifKUov71rA3ifyecFYH3JCFZMGP86M3bKzzuxW+8+t
2xwsKQeHAoqDiChzwV5Q0oGtRIWJDPWl4ZCFuOVfHrMiAe//49kKcOqA63CMIMNH
ZtkQ1/qtFCduS4/5k7N2EJZDSOCeho25ka7FQ7uusJCYC2A/nnfeGMaRUUFWGP9f
nmKlRfeuFkdZ8Iu15XchzdpSTmmTdYgSxd6gsV2mxONTQG0ySecKw1qFUI058Rns
T9ziqbI7hQNBVYTcJqA10K4ZLV7Oys4SpWRCRB5ivYa71GUNK3Z5uoVNo6XCopGJ
AfVMSHwfj/CDw2YxZPdVZ6q0U80PwU8YAXQc1nlW912BbbR7ZG/7q65DFc2qYAbS
RySBMRBN0jJka5MxX4GZtEIcDbcrhPCBxrLeiqbHfZYDqQJ0Jt/vVQn3bpcNEtEl
d5i9JuLObtejfCHphLJMKmUIutBK84+26Dk1mjpmYQWcJesvXsXd1G5beUQUWH43
nZClYLLnOWwhvClxhirdoz6oQ0LdFVh8nFKNSwmtpYvW4MUDJFuMP8UDEzk6/WTH
GEgZyd0tlweAx7kPY+lye4hbnQw9igx7FH2HaoPIhAmQoMuqyuiUzvNsdgkjB7ew
LOuj97+ANGFm88oalFGGupAvle17SrRjn6TmRNmkdiRbRcuSQPq5LBOyXXqOVhHF
VcIIeqKcsR1f5LHyLRtppoZrYJLRtunO32ck2aZNlWN+AjnBDeKCEOuZNf3598GE
h4P7ROKmqPuBrsFrQnqxK13IMB8NmAKs2I6krBYQu33FZhmNfnbloyxUmaP6NRTw
nEeRz8cI8TvtW03SIqxJ+Dv6LVi8o7aWqWV46EfOk23sE97wIO9Q30DO4l0g21Jj
n7ZoxC3MqDivCe+ebV2BHR2SMeJ9Fyt2/bORR3ntxqA5evQO0iJMC7PQTJ7NskIf
lOOcDbuKTBPPeAvfPtdh6xKSfu2L5Rqm6zI3wRChWa/uDYeBbRsy7l0u8E5iDXPx
sIqHfN5pVZMTBw7yJqsREPmu1eIMOVBFkadPO2UdQYoLQjZEMn/JCbYdySlELLXI
KtPTRMK+QFiXrAwh86EvR6F122LDUOMx+R19K7r/lRz2yfXrrMS4MG2XVbe9rs95
UfoRwj9K/bcfPXhICjMNiJdq/RpstsLcy7PaG/eSY/xqrrQMHxMG+hJBETyr5Ekf
O2lym25BcaK5Qvet3kksAgGXPNYHtGOt/ZAWywGderp9ZjGjFMegEUcJEcQ/gRO0
YHXEpqh+qJyOz9HynrZNJfjd2/x5GdZ+0tLDohXmxHXKn85lzXer+kPmAjlH644I
5TIOxoKWF5AdAdcq+ttSb5Kq5JUllFYXvvZ2pnAaEkMwtAtsIah7/geiz9LoWZLn
aIP4m73WAR3vs0HAGFvFqcHmONctoK37ED2IE2Fk3R57omWzB+Bw7+0Y3J44XISe
pfKGhYe81kkb3/4um1JVkt6FaUtf74XjfnQ5Uy5gi18Lx/+O7h9mQh8c5wCxcP6G
XipATpBKiotBz4BB0Iu2ow502oyxODisRMrBq8G5B49+VCT5vB4rzaFpf866a+gO
iAnl0+fSRmw0ORXaAk0I/qUJivkGj2CRP2DXVC+6j8lodEIBlHrbCMt9uwUmjanP
3gaBOMBU4Ur4GpTXTAKQUBOLyWg1NzyVmBmxjeyAFJOmXhFacLnwyrnZMZWYC/19
B7VFQTzbvDqIFCHcQht838rVFJ7MNG5hOGI8jdQEKuRNMS05oVLzGz99rAppVPU2
3Kkhd70TM7XWvBsoOm7xxGkWI9/hmpojp0LF9cIcQgBJw5SupOXDdMc9/Thk6F8O
ZUjouePxh4qfYBtTc3foMZ7eGat4miVC1xD6J4jjvK8oAV4LNfo62puECYlyzd7d
v2TxBkyNwMgOtO6aLLOolWiraZ+BUvxlJQsOylP5/JubT0J+GPZuq0zDQUbSGYsA
GSh5k62sy+T8LQzsISkkLQzFmCTjx2eqDW5RH1bpylAUBTS/NdNtvAdScL4UhxOM
UxDH++fDEumjAZRKWPzfrlg7IflVcAh5ijUczRlcUeFQk+9RIw0HFQutDSt0EJhD
bX/JmbQbJTT5yfYPjUAesZFyyu2HWo5nKH9y3E7sxWOmPnFaGOWBmNlO12xlrFdA
4l7HWCQ0ZGavttBwMzE6LdImXKfDQbxEiZ/HVQqDUUly/m8lrwU/OBejGnbFh3Qb
wFSF4HZgCeuwpnJ03EcgKyMAHY2VXUq5uUqMfor5qPsmNIUUAgAlXPRuxW3P/OYE
1XuQxiIqttLA/22bRc5l7dauZwNXeujQwv2HgLzRwm60fmNy4NlBK38/xZCdiU4I
wzfNvcco4zvwKJziTg1YvHBrQPfalZz+psoCyFdwMGittIlA0cKPXJTOYoMWOfvI
VdfSvWkE8E8uN/Zkl6eC7GSGLB+33Fw894Ygyg5HTivVOpKXApD9yJ8vIeWmj3cj
whZfJe+TEFXLOQBtj/JSPkcn6QyKPCW4TK3N8eB7XEZT0OyB8QMQ/OAHk5tWbLb0
t1kC1QtMeCOY164BDvNTk9KTBB2uZwIsVX+PniuU1nGokB3Xk7Tx1qk5meWtMzBj
juwgCLwoZL2ajGSv/8BWDXk8kHo6vP1yNyG45AtxIQAolSFbbt24QmQeEIQ0WYbY
P2m2uUndQQ2hojXOnEnxmmYX13DsgQTWJyfKdwiiLOL1bJRO4sbKZXA5rj6p9QqQ
q9U4V/Ug4jUEDyhmud0whD9A9s+qmT6V6ZwzBmcxg156eAD6uxo83gI37dZFRDQ3
JmrKUjXLpy5nvdWVoj7c5ggHcs5XK1vD26Y1tpO/U4zjjSrczbWWBNTWPakZ0zUH
6/8K4qcwOm/TEls5gQhM/pRtrUkFcsruRDWO0TWsR5w/MTOt8tSB3pWV0e++hU1x
8FwR9aZBbPIREAK06/GH6EnQDCQikvwN7CCSWs9BTIZYJBWAQ+b5G9tmiJKi+wqu
H3aq2jeFqnEG3wVtPsxBWcjV9NCn5z+TcaaXBWjqcGgGOkiavIJtoTLhz5nSnCD1
GyGvHgrumVVF8VREN9SitHv6EuhlZQePj3emAzCc+UZEPFqTot8SqKHQVMtolcWI
71a/H1mhCvCsnfuPnoKanyqO2NN1r0mhmmu830QgP6L7dROrvVmqCCtPe3QInatk
zkS98zu88Cb94YS/Yq3wPhfEQ8gdVD53FaEYpfz8PxnT8oJsYTw7X0Lobaf+nMCq
prMpZmLr/n9dt143I5gbKavq3xjcUPUFV8wsK6dkLkt2GDusDx4RMSONhInL6P0R
DdNLX94ddSvljbWlQ6XS/pcZdI6S3G232ZVELsWvJsMCtFB7Yi2dErX6mHxSHASy
W/cm6kU0wIx27L/mjUZ9SASkxJDpQ72RUUNtK4movlHc9LH6lRGms9EX9GtGrJX/
OqF675qx+vQKbNXvLlsK2nZC2YQeAZLVOHRVBCHnpXAGUZVCRvOPzQ50SuiPuGLe
Vq6KsZtTL/Ld2RVHfDeqtJ9h7xYDoBBSdGnHbD6i0Yf1F0bnac/SBe+qZES0gewS
0jK8aVAHedePzlRYbJF/LCEdKVusAetVaPRaQlwjNeX++b0SxWiN8lTf8TJEynn3
1MbZiWAcAuF/B18EvJ3r/GcXB47wmVR7CuBUBAZWgbVOMCHkeFk7bdcYVxKWT3Hl
H+1Hl3uagLyqXoUqrMxDHZcL0tJXAd38d/2u8ymthh//9KV7HFvUdFwvp9NWTEfx
QO7wTVdXkMYushm7IHTvIfTNHDi5oUwG+aJOzLghbP+0Q+y9XjR2h35k23ohqWXk
Y/A7tuABP7XE9CKx3FHFQC/Tf/gwQyRLFrSdgbufBaDWXzjOQU0FHP3dJ2xLTMTq
uCDXv58RUd2kn602m7l4Ivpc/ASUM9PsT5CwZF1B5R+KsPvwAW0+qpC+EVtZ3eIT
1iq1a+mWuhtyBK9Kd9vHsG+6p+xW0zFQrOBWM2HDaBCiqUr9khsn8RhcJ2FXWGmL
Tp5Ow7lzb5QhNPYEgq+O+HL7S5mh4kY+21EpJLZ4OuFUEJcu6Ckczo1ORacsEqPl
5JO/DtSYy8ANaUHv/myIVR2+GC6jjQD4i9khk9hRYYWIqAlkfCOE3HQ8R51bp0aU
Ewvb4HhfM1hqhLijhcC1Zh5AhHSIlYwn9LNnJ3g8kEoxNhEpcsfy4CRVNQ9CJZqe
4A4B09GKQ0DoyDEoWTWExlF7x7u8ll7iJV1P8JgifafCFl2/s26l/rhQQRaaHWmr
s5/l0vW7zlWSl/eQTccskWhSk0Jjd5FN72QhuplInoiUCZ+0E+14aSR2Vg9KNEcu
4ShzEk2WCU/EeqdfUJ23j4QlsbA/PGrrpr8fd2Po6rwDBGppMx1ZJuM+sTo90owD
RWnlvKkuGvy9XKyF1Y+EdXyJan5UGxkui0AcLquq7P5iX5nikmCSZUjJ8xYca/yY
INvtSuAPf22U+Jn7NFYB8Yg7X5bbq52JC8aUTOEXLx3hihqopeFuaJ/OfQOGe6Sr
esMioHtqcmgHh8tG0r+2wfn5BjHLTSISuyxYsNfOW/ImICFFYXajE3iiQMx3HFeH
TlKpNFgO7rhTVvLEkbTImBJubbmgn9r54jB+cXZ5h+2oSC1f233suowUYKhSbSr6
ePysh6jyk6Mgwl51A8SL5et+/+CrjVAj6eKSbzQ6Blpj2uwgIfpcp25DkY2Qo5rt
RTCrI5N38jAdn7Pt90Fu76AavPFHxu2/463kQ+Nf6wqoP2lrkKUhQ1KjLaR8k0gq
wDhOcvof4SlBkqfoW8F9709yXrIUQ8CoRBWRZP82oSmTe71991jkZDp6hPHoS4rn
W6xjxp7dCSgnS/T41MYLeORSYSYoMIXBR9FAKLpgkA9biLZdnC1rIANTFfUU/7KV
Q/WeGaXoU47T0ypkO/WDr+WtZ+rlqf6Ub8VRBRbqQKi2/pV659DnBRX+UF32ytKr
1vV/TRYdKVLjXFEn4Oq1NMVEzYog9YrDT5XYXbbz7HBvvYPCKOZaF3BJXH4VmDot
z3qxyWiHThLnStjDQVtTReCebztRJE+DkXOZXNIzNzCG7ENhkmjLsxFT4/zdZl9o
y6Zvh9M7T6sIFfbv1+v28NlraKdzSCebeLvWIyD+lV5L7G6hBwy9VCCANjTWPSf5
A0DdqcadgCik7vmdtP0YoovC5CWlzXko3MCUgeVX3zCcuPVqet8Rx342a3dCrNcz
6eFgZkOUqaDbFxI0sit9m1pU0SJtfOsV9SJvKcaJ538u1EsBbHF2sVCxxDwa2BfN
V38ooipEErcsd3M1XWIH5AapnkmOvDS16UYtlVRh5bbt2AVNKoH2umU2tIp9RuSe
8/XgX76+qJ1SdLi9W5XL8ualJ0e3rYs5OFTjYy0/q8NajoeiJEplpWnls9Zj3FWQ
VY5knK2TEYo22mNTvUeP7IE+a31GkhyIOenlPl1+VZOBNR3f9rZ4FBCrbMyTLmIq
FynJourjjtemwffc+N2vt5oTQL6bm67NwzstErROznpztKYWvBJHEMYRFEIhdQIi
a0AyAw4NgqGoehUYSlHjXE2u2Lkyx0E0Ho9T5Hx7P33ToFg5mBz1UIaqVpm0xKr7
CxG03n5qhsBsc/DMiVrVjB9w8kHPqa6OAugcj2/QgzNMudTk3E0c8vZ1EiOIEQ9D
qB08JeN04SWi96OSjyL48yWyyHf0DI/8bqZPp3YwlxLmsO1O9MBLz4X+k6z1CGxp
mHDCmKlWt4P45o0sxlhVSZC3zFysOjErXrv1rvWn+vg52F4cf+0MvaT4snJo/9qi
w1PRZR23D7uYgKdFIIbSKqmcdNEUgShTAAWdfq0OiqHJDniwxu/bH35fr13YEdVc
qeHMMR4OFL5mpaYy39zTfmr7zTIMgxMSusP0H0dHN5JPXJHCB8y4NjqNXp9a2f0O
+hUAtlGrVwLAajs8MrFzQXd9UC0Qqt1GXP7OtY5cWNMIa9uuKiO4k6VrvGdCklFa
01YlcSNQQkqZ3PE0M7ApukjcQf3GTi0esdJVZP7ex973k8k6o8BG0mK4SuJpBqGA
hd9mI94nXn4SrImEQAHbFX/eMNQrwRIf9pjav8zPgsAwx2ZHEZhWK5/FWLuI/k6F
xruY/XYWE90RH/FX5U1YRzb8a5woYiXhMmQAYU7DP5Dp/2Q3HCND865Poa+0vuTu
CeG06fjFYWdcDytEYcUTaHN1iZz2brQKuO+E9jJ3Np0TUppf2vU3BDjZ0bmG+PMT
4pGM2BnWREiqsZFOmTeqTmyL2nf2kb/3aRS0R2jj2oCU3WMq02mNEELtgVtqBFZC
jm2tnkf6iDIYTMUmD8KvOUkOeFGMku8QKOJR1RJyIZsskD64LbOlq2C+Bz+2nixG
PhVp35+LuGuKzD0iIrtWiNihy970OJiQqx8a1IkgheDyXy8M+dxEWg9kuhjDcK3c
TQqw8gHDMtJBJJ7LIJuu0usmNwrlVcCykHWpuIlT2o4JQbTZ7Q7ICxTcjU6BZqSx
KK3EEcIp2VucF+EwLcNhh5LZcrGmKvgdn5wQyK8sA/jEtMmlSkWoFjePTF4aLE4y
UrE8KWfI0m+b7XFEVMoINwlcNghdZdAhq5Wyh+AsY9YqhUXuLSUh3R9f2nWkihG5
c3B5deWLPs2GowLk4FEEwKQpiuEGMQVg4kezfqCJxZIT40/YOzPInDjfB+FpUX1p
cJSQlsoFN1Lvq7hOwnJjM3u7aFsU3tv88TpSnc0nhrdNeOqEglh6khX/vBHGZk3w
Y47Ucb2qar7q6i77L1iVEzz5HydCfBWs7mDZi2Z1Jr4YDAN+exJaheRS1vCPCQqU
EQQ9Tsd1wu0u4his2ntzk6hamzE0BX2rMJIGJ2cDOADh4xE4EOa8XOWcIFJ8rofy
IhuVpUmf+TAgelXqJh5VU7DtJMZ2RA/4weJyb0sRD7UP3M3gE2DpnpCoTNz9GMGc
Rw1VTSGx2cVXeExnhXL7qyHOdg7LJbOwy77zaEMJLOw7SWGctbo75eu8Gzav0ztK
1JxwN9DiNEc5+jfQ37wqetK3Ji/qO8oPPI8wsfZ3PsKE4LS2xrAAzHjsnJSNv5SO
PV0/Qm2VL8/F28CY08jVAE3Z0lUB1+TJKOYnC/AnVbfHDYypo9OW2nN8J0RQtwOK
JwRYhQ5QiV+/ndHpyi4pvi/LORu+dRDNKpLadCNISh10BFUgq5rZOSqqjmvTJE11
gKKcMNFpIm75ud4UP6NwPyDaYsr+QpxDy0dhQ6wRZT9uMXA4R6xvJ7EqwpOfYknj
7mgkCE5eVr6q4ZASd0otwFHdqo9qFFx092VPpLu4gj/I/JIaYeX8TA/twR+2tvAo
7sR09ISm8+Xc4RCBOF1olkCqNqsaVyQVZYviy2CVr38nevig460IKS+dcaaeCLKi
mm0JxTk1jC2zKlm9dTf8TsAv0zdMl4SAJYaJcpODoRus+cA570FKjwavy8T6+gIy
HaZx0i9TbHRgSdJAEuA9Axogc/2PvqKsAfBjbn/ADwdjZPn7X24vJGY9eKMm750Y
ZfeHOynYqDeg4k685fNUh5xjCLLATXpEoyPw0kv/j+vntqAFepCVwAv4hz4DtiQh
ku8bzzoufKpBWKt6wn8oJlrs47+exiogr54YF3OuYF99gJyvwTX3bL4EduzMR0yO
tR1cbYnOnnlgZWAJ9xhxPkWv3Oa2P3oYVPLCLrpLhYcyKiHFTvTxGVqc3OIp6uXp
G57yecK8w8M53Fq+rnWSL2ZPKxl1RFVXKONPAsnMWPYZRPePG1eH5ervmcE2ocdO
gsKYvCnk0PFqETWtfO7u7McAW+T6BuzgWsIVvHmg6a3QBhAlRBthj3xWyFBc+UZC
eXBKxyGL7DR0wgq8vRpuL06W1vscviTm4He+miwikEpf1hNXaUXnQG1fBEMX8/wf
WHtkDk3RZgwgrt+ofnqQOTGLlyHRsZYfsbeqoBNqroqUAxf0Logxz1u0KxNX0bH2
vRQUmy8S1PM2hSh9oKxnFl1d2ol1ke1M2nFSkPLIjV8eGo0+toPE/HfoDLvHhe4y
K9e23A9DpoN4twzFlITY1NG2XF5nMynY5CMU22Pkt7MtJkZzUzwPO+j7aIgPixdz
x4qhx2nm0vWobId3TZ9V3YUMEH+b0rNEZqkQOJv8ipE4QLINIo8EPhzckrmWtYLP
wuGpZVNwCoWH/4gVFuqpWvuppNV4xCNLx4xGbNYsA1z2UKYJgfql7GPoN72cVJRG
utPDX3kdu0BveU6vJLjUgM9GIu95L/mT+0obN67Dj4gLRgiEh5xbNoA0mZaRdof9
KbG4E24160J9a3oOaEwStcsZ3TFdReTZT4v34R9FRHwsQmJRjjnM8OYDJyNiKUNa
oXhRFZSq+mfe4eOd7NAwAL9jdXzcSMHBlhY5v8ZSQqWR7vldthJp1snL9JLzFAi5
Z2yykcNWNV1IjY2hV7me79mWxAwiOJcRz3M/vLDKb5dE/8djQPuoM2IgtFvEJptg
lGeBzpH21DbTA8Hf3mUvN4V/IU/pH4aX6P1QuGvK/UkMpSQgQtP+MEZdfi4qPrgK
+JKwrX6LMDKXSYVL7RiYcKauue1mFuOaGQe/onakzmGzaaCsaJd5Jeh4FBIrB+Z5
vLDRqi/sRT304Ehr1KRYuw2jqcuILfYPWopyQGtWG1GMEpRrm0FzIwa1H2KIojEA
ADre/rMtmKxN+ZNUQSsxWdmZKeyqzI2hIWl+86RFPwjJOnOhvWbtWZr6iO4VJlhH
OpbDn/mWKjfQpl6rUB7+/PXoSO/SntyHn4PjdN5ZQytRZ3qZUhtJLG5Br5SEcCwk
uKGzjL1W4bedZEyE1qBFFtptuSgZlVD7gmwp7JRH4QC1ORnwQg9Bvll3KwTu8Q2f
6fgF74sMNpMsEiNLpjsfuj3797R9QJGy0RqkMDG9qNa0VakanCKbqfowDbpz9VX0
ca5OocRHtXtdchmN2g46NKkT9K82djn1SmTjMDOfCJTkUPVJGY5ZJOmbmYptYy0S
M5LPpKqZ4sUz5q5xumLi6YPpUDPbOfdMjACHlqyUbHF9Ki5ytt0Ne2R4h7TgHqRG
u+pk3tv+wN/RRgNMjzsaXtb/goe0uo+nK+AvP2v40ggaISz2s+/+jPqr9S9MfQz9
rXRxQgyfGF2TOczLC8kHR/vC8l/yG8P8+2rNkktxZx1s5F4Zep/thq14PAYSZA6s
17gPTGYbz8EbTKz9ULP0tz7F5cMYWaRfsmIlIHjTEGAPViztX2k1SKaxJ3qhY7cx
duEC638h6+alwlPrmWWx34n8JFEsIeDVDcDqXk7mvdAVtuLUMkn1XSZAcL2LOB+E
txJgjBfzkddgQkYumKIDM5z5xPd+HKtScrniSRF/VBHB+sTSNTmfx2ELzB08b58E
RZkPQH7O8lxLNQ+7kl2wNzA5yLiex+21C7hFDopAMzUgRbLoxvrAqf4DJSBrSUzA
kmPop0HimLJAq51PENsedTQYWUSG6RjIIzKQ32ViBdVUWB2RXocSY4vu9vlrzDCf
XarocR4f4aW+DfYXWZpZwyrKrP2NtH37Gbs02pBhQ1P4zE//p19iOEmT9bn4mVRA
flPa0q4v16UdfPqoQUD/9ZUSl8FWQKVtYCjv0YKF+GKjvoGnU3/zLnx4frxUMm0g
TQCxU2ytJtoRqTb14PnxexWArNVObuvEvlh3v9vJ7aXrbyS++NRHUvUSvdF5MmBF
z6X3o5zY1w3OmVErimWvmBY9xDH54BS9UiSHEDPdz9bOAGIr8S9jrtaWVW3a6TQd
doZ3cW7R55OZnF2tUigxxYxEB2TQw314ARthZdjbkcLw5+iVAksTTsBrUlsqQjMc
vc8b1b/sl1eYlYgLokk//z3tzOmGczvty8h+5Nv0Kiig35daGbRyU6wtsJYwbtnm
Km0x6Njula5GBkqKzXYIb2IL4++GcWpId0CXculLIMZOYcFlQNnhOH8u2PBRVc7u
iqcGrVdEFVl1Peyywnx0tilptbDPHtVZefOFbj1T1dHODXGSYrIv6MR8vnjCIaP5
/q7Yq9yRiTvYG1yunPpiDycqnEEJ9oYtkF7SLsUS3Hiwt3fa9QSExtFKh33aFyGI
rssSPjWncWeRZYI2LZLtIeJVn/stnrDzWOU9TBWpU7bIKfwcLl2yd8OMWI5QyGs7
nUgSfFv5YRkKjUQDKhIWq9TFciA2bOr9FeC/wWGzJjPVtt37VjlrfvR8b591b0qM
bPuL+Kf+ir13QmruAT6dVtUCxzS00j6s+vFe/ypA9M5Xwhgoeqzi4kT8lMj6RnjT
JKA51yo/DlzYH7ckP6JE9XoJSSnr6yeIn/RmZ9LY3R4KEc0fzFRyr/r/GoLWz4W4
EI76UBnP8Xio6shkzDOcFYgmz5QKO1KRivUkLP8KdYV/02Nn7nnaayUKedHQRDm7
+S9xWFQFEhKOlkaoWTb5HOGa1t0Ss9awirGeFfZhQIOoquG1eIscDEKMsu+mvIvw
u5MBo8c1PIDTl6r0bprFK3X105WlgCe0J8enRkUs9Oi32UO6T7G4W9ZvI84HKPcl
hQduuQPpgxfJJYYlMpOiRyX/UZOKYhDa1q9bLJuZNhItv5UNUxBv2sq2khE0z8mV
6aN5t0XUodf8U8Gs7f54Zq072CnXlnBCe977GsWlre/UgCZWTpcazhM6WhRPDXlZ
BMTkw2iW7i/EQoC7FSfkOUn5oNTq2t+LhqjM9Ziu4QJqlv1r3hXOtFBhma6GL1BY
99mtPzDBr4+aw5omUQb8thpvN+bUdLdG+jpo25tMiKmLCnAdkIHm8uo9sbsfghue
X41o7KLCj0yPk6C71i3c95nSnqjuCFv+A9e/vYSAfQLfW+7Fg9GTy2DNv7u3VXX6
DofTuAJIyyo3VlrO1r8namI9Gdm2zNI85UhtHU/+W7VIkEwLdkjLun5Qm2J4LH7S
wl4LlC0C6fQNATynr2b7YAytz28+Glz/1Zxm+wkwY9RKKUDUn1UWbQFpAShauHf9
Fo7VyNYT7dxBqj8eCjI9bP1tVeJ9eIvy9XBc1de1XKTL38XcU7w7biujN3b4rl3A
i4k4ggcE3X8c/F7l1UU3Vh1bL23+nCzlcLZt+OtGJ0cje57T1AKDTUVwkyjrmCAF
0/voM/q6/mKfyalhNMgrvFm2hszr7U64HNC9hUeDKsNliSTPNt755+P1nWMgGyJY
GoqU9Vrowtm/xTHSFAesm9gziojv4Qnb6mJM9WShSdIccXziK+pwckWuoHt5YZ/Q
G+wPkMSCurZssJ4Qhy9pESFbRGfn0gjeq+Snptiy9TcDdE+zbDfp0ILWeDUCUUi2
xUFxq1s0OkOTIiO7pdmiKTSM3HZQjrV+bVSKA3DgCGU4NBmZhR1g5xD1OIT/xjRS
EaER8lx5tdWUo6zukdZEYplUlEG6R/3v8OBrYL6v3eZnwlTIJuXaNqnGph+DjVn2
PtKENhT2pmNbPHlpGRn4v9GgCXF04w4vgYU1ayUCJ2tDzTrpobpJNtFP9wHFBT15
nuv0WSpFsgE4ssT7mn64F1zAnXYv0FQdKtr3QyAFuhRInhGGL/HXpxzQtp/FPsrW
hP+8d6jnZnYEyIFdHgIi2tz2zSoAeUJ6IltYgM9OyrxtlEl1nHjMngkLmjw1qyQL
WI9E13A7GbjfwQSnH9QplezKZBogoYmw4csPBJGlwsPAb40C0fma8BtP0MBEoPpt
dAvRzvsra1P4fzO/EpaItqmCdp6k/s7W2/D6s/7uIfUfMK359ZCYKgA5PBzZvPIG
PAf7H/qiLhdmnIJF8Sm3U38KAqNsI85PLCy7k2YC4fgQv5HhTZmoW6KQ52gxUTwr
8OcfWMxmQSTYg42/8tkulOL43uYfIQ3KcuZjCuO//aly/Hu+vSzZJ+jw6gMmdBiO
ntY9bfyrVt6svv5gKLCx+4sDokKQPXFJeZd4Rr0HU20XKBUImMYuYkghFUXzHDpP
gRYULAN2+xcA/bJKmzKQ8JMhyaEqMIJb6OgFA3qxAgTjWzFEBJNP2q7ACBqWtZNC
QVcNxKDtHhF4uDph14P+w/KQJPWFhTyMPo3T4Gib2HHGD7tazkzYZCt664WgzUUA
ii2bkXZdDrDHXFaLWGRcpjsBPc3xKBgD1LTAwXTgIWv0rc//fEq1i+IiZSKHsJOD
PdNACE2MZvBWIlkP8XqhDNNy6R0maivpA4vjXwPheTpmRYz+pUnS2rPPotBz+9Fs
oso1D960t93X76UMZH8vVQYMbwVcj9yG1VX2ZuEdKTo8zpDZgSBc9luf5m4jRxy1
tV+FOtc2E1G6yLv7nnH/kvsocaDRgEoDlHjtKYOtKxZgwid7J+TImMFC5EZlB4Q4
jhJRcHPHxuEAx1NzZwpGokMKTIrh32kRAD1EG/TL0kxlrt+iVC7rDrAoWzWDDa2M
jL5ju1hxC/XUOXvNwqTyKVdrAjbuCnIrz5/+MANavw3eqhxw66HX+EoO2h053RT0
cb8tnPpUhYKpXs1JMtu+B/U2VvD8HZCOjeZLXtu6UqS2fJDH6GuPqtqYOq0ygQdF
SwLKIGnw/P7GE1XqU6JsnUWX6IKKohVif1dn4DQ/1bKWGc2NAjgH/1L/QfzzUi9l
/j7yEsBqQWuflEz3Zh3uxfYC9cMcnCA54ElJWVRroqrCS2x7u7SPwVJMAFxiIdiz
ZfSWZZrqk6wJgvzKzq6UJtu/L/RndZvIxrdU4Crdv1HV4dhhTg+NJKug6DQsJtmI
LDcsJYIu3CPX75Q2uQhyT1FGuKwnY6U8L4MviPLfREzTPlC7m64SPTsHTo6cSs6E
43PSQpLTxLgAzN0kahK9enbaoM4LbEpK+TUvgcsLdrsNWCogK4t5D0Gp1gixLmmT
Zvkx1oO/svRAJay5RWC+sTN9rZyXmbIsyk9gaE+Gqfd0AIASVcu6cqWtCoGQ//li
tJ0gj3vNLWIzkCakTR3xdSHFdklK9UkXaMj18i9IiuD9poAsh1otNfL10N7AbvTG
MBaQVvDmzOe5xt9lcqfZsI10JYIbu4AbfRlYPi+C2i4Su/3j3SYhjgYO8peVBhnF
73Vh7oi9A4Qp1lVxFM/uKks03IuQazyNnr/Jyqzav+pBf3ZS9ScVseAhDKUpu1Tg
+nr5z5R+Fkx1sbU6FvNPhwxlUZglqcFawOeW+qoHTzfd44NL5OVp53nHv2xLvYOP
caMY2i/JYhJvNQrtjhFufAkNN/rQKEmaEJjlZ1uKIJ69wApLTq/XdIPNBo1twmex
m+oH1qkK1soQ58thAVkj+6wrjQUXC0k+PHtTgm0ssrPZQPlHNnsS5bXJRTnAMFs4
8icNau6eXR9OT+Jk5EQR3Xcf/kqB690FaHL3lEi9PD59MDJJVMeaek56MaP1WSp5
tvjE6q2g3m6PrfE4liZjuKUl4EBIoEe8GUPRryjDTjTlFjLUYRn1AMtyq8Ljw4zb
9G1A/0kdgZ26EZ0IEAaDiTOFK0lBPsOxA5oHW2dvFDg2jIMgwcpAFAie5lE6U9Qh
BScpy9C/ms4ZtOXRWbOhppQboOx2smA1aI/P0+OYLm814B7yjrVdbseJ419equ12
yjmzY/2LQW3URyCE1YR/3vT5L/7ThsDDxV67wb1uDqlXI+z5oUOi8g0xZiqIKIP6
zfweqvqOz32GdhxSV09VsyPjEsJfZeScWa1ZZ1Jh+FcS2u0EVGaLuBFoERAXsNF5
sm1kFmpS3QSot8szZ+VLyi3qBzBoANPeNxc1CXgK1Q02jGaOmHkHNUm+PUb5xNlb
Y/7t6qG2dLz9FdDczrbjdhetw/nQuoGiklk3bXc8xkOOTQ/4JHcSt0usWZ0TJ7Mp
bjOm2PZa2bcMvOyN7wR8oc4TvQF1iqYMzyPZ2RRHRe0fQHqTi9z8GByAoZN0jnV1
7e6tA7B64wh5Iamc9zDPdJx6F1YBC27MlGVw2wepVdf0f2owwdpVD4G/MlD3rNJk
/goBdGk2haI2gBN3SSzIzsYEm9TVfhBBRAcyiy3PfB4Gr7tEiyJbqS39ePjvYhdw
daxVPhiYvP0HuxkO4isS3uGJFIL7cR0FF1vtBP67745hsK1xB7odATZIk/3vKAnW
o9Az43uFaJmx2+HHBL4UfP4Q9j/HVqjvhHsHq8Y7xlR9vjsnlOph+KX1AOCkpAtU
XuUMI9Kyq3kKIcL1fggIFZAUTu65YupsINdXGVMDq9Py8+Tenf6PUEL3Aq69xxXE
5C1aIIMA9LLlB6/4ZggUC2SrGMkzCTa/Bbh9mY8M5A2adZtI83cfrNF9mymNsrx0
wpZGDR/LPRvgBUpCzTL621j0Hkou9AEhRslM0mdHgYSZDtiQPgbquede2b6VGtjy
vB/KpLbrfa4woA4YozzuEMa6+fy+odiU8s0a0fSoOkGiF8p8AlseyqfC/FSRlo/W
AMoGJ+as5creujpf/PCApzMdd52a/gaMVIii7yRKP4CCTBeEuhemkOYNakV7f9XE
F5zYPjElpn7Q99fgkem5O7WaCTCssKYhXBify42t2HjvfDTCj3rmmM3K2cYtUe9J
TkYGkyQibdvzzAQGkfCzPtPLKKFQubSIXshN8dWOG+EQStjhz9Rn4ixGJ4SSlYVs
ZdXgxg6aLcvwI81xSYq2sakcS2STFXzF9hKE8EZxPt1tGsna0QYKlSFF49oveCkQ
l5E1uF/7xTbzH3xUOn57td/V6hxhCjQo2h2QtP3/dzeEGucRQPn1fmTLOUQXhM0x
h6vJbGJC2HJSDnBD7cFpig993+Qdoa2lH7vkQnRzQB+UAZQBfRJ23N7YNOKa7ehM
79ZCRf9yyjgfUW9+qYM4b7xJL9hZFCflXrKrnvR4Xr/r2/C4v3zlxBbvTEdpWfg6
UWj0hTZRVeg4Yr0idnEbMOsOkcwQkfGH6X0VEdZpQh0sp44Ia0ISA0KHngsPpS6n
zl2OmAxDYi1b4TC1Xzrn/NW22Q3gJRyA/iXcsOP91TklOJVK97ZHgWoDt/23fx0F
SLovArdSZ0hnyuhVoq1r9Mp9HNP/96AJRkLjpurL/t2Tbh37BSsPOz9TRZpkL4x3
rtELVPhzjsePvcVNISBQCCEgd1yKZKHCmC9wrEzCokSaVNc5P3jntdT/ZSKfcodh
riieTN4GNUFqRB0ln2+wKFNIU5ahBweXPQzef0rZmZVCa0XTSWkiPmZdkSx7tO6T
Q3vF/8BWc/E9MLBsPUVd3/LbTueydS1OVKOmYVB3uiVF+HiVZVzl4lKw+q9RM/nU
0VxtMQZFC2pdavVr6BiVbyEKNuLaAaZfymHcEWgK+N0rMx36UUi5xsPvfzYcARtE
fgzaAloR4KXZx3B7YgxvRI8uAkj40ULWKYgn3Uk26DFwqgze6hcsDXJnnU2vi0Ki
YrS5qX8KrIbPdHWD9CEbvPkl6AhaZaUdy3WhO42qvzkzN531vZnfn0Oqn1QlXs6v
GO9gZmWp2GjCx3sCdUKv8pwCxO69x3qqsX6kWkjosjK1wBkf0569ZsN0xmqYfdeV
rF6s9GQAhhEPSHjQXfM3jMqv2BL0iZlXtcec3QMCYa9EmCYrLMTZi3tNeE1pubwx
hbQe2fUssex17IB2f9VcozEFOWp0Vbb0qpa8TpdNEQxkcI56hNwBILaq2UBkT8ZE
t6BX5qjGRK06908RhxoxJzIKKE69ZjRzK1A/xgveQzj8e3dv7vLqAsa6jQPVsPiI
yIu1KA3QF0zydRaEaYfvHo3+bLo2ErjJuy7detFEFDGbC/YdPCxLZ4KuJEsjtZlc
CpazUjicrYgi5YIRs1x9LctGr3LT26AeCuMk542UroDCxZkYsPxzObXOauE34OHY
Y9Be3Vb2KbGuKa/N2ZIo3dAN6OW/RWgCJLyYL6KXfQk/tcoROT0TcvuKR6FYO8wn
0dRWeZz+XPLPq0SdOGWwgYGCzlF25VxOcS1TNIX7Jg4mEwugAZsKyMr84By3fLHK
WQaUzrD4Npk2Gy5hPW2g9pEzuoZZex+lPejiXIZPqqULpn2/9NiV5CIGxjRYogVp
Ylc1fklq4V9ox18SqUVajLQFsvE7j3KFfCWD2G+j2op/syjmHYAKn/uZRd3Dv4Rr
QK1enkp3AO8K8DYpLMvNIV6je6pdN7aGa2aNfizOjstrucUNqHZZ3QpUkMB37bBU
j1AdQ826GzQL93GT6+F2NdlbgVFAQov2QgG31bdHyKKHk1IbXHxO5KqkBjvJ8Wds
OJZ5H3w0bF+GGe7Nbuh/8JJF9IVJrG8eU2v52YhZsRrn+XBDkSBVYi4kDKiNpnSg
cbMJ38d8RuBlIEnoeKgtd0TKegurG+S14p/94v4zAzp/YM8zfC/R0Qtibq4lH+uu
51Mw5zgtsWJmSw//0P4+8IuPJ7aF0duARbs0zGBYdl5AJNGC1hKqIIFOLaDJMEZK
bs7AiqZqZnocg8MBFWOTVsRO2RQxwMWNFfk1i5i1jRyH8v8g1NRBBnS62VVV/Ab4
KH5jWc1uFCb1Q/9Z1m49Cv8biaoIoZ2j9TeA/DSAREk1c4lTSpoNZAZBQTyWkh7F
kLpcXPYQ8+wKllKnULlS5aKiguIt4Z4s9IUn/rvxgNehJtdt5TVuaLh9yyXMfNZJ
V+Q4+3amSBhFXY3crA2E7fwcs1ts4FI+HnGA7CVMljHmYSBey9Kzs6Zj3Zdrsls8
QWbcPT5jF1Vo/b16Ur2PFV3WU5Ry5eQq9vE7u1CXcfTl6RecTgnwwkkm8SWu1qjd
+wEUslN4+gUZ7bi3xnMA0DClQYLuldtYOIMIC13jL+BcSqNt9C/q6/tXY0jPmWs1
O+gIC8Tx2wFJdO8ExqtRT+8SlXGLsHLloPCeRq9mAQOMzZB1uRe44Q7m72GLrnLq
C0B2qZz0vgStVFIfl1/K1agCxxEnXLITugcP6t4QDZwPcHjqllwlBa5h+WIDpWPa
Ki37zbqIMXzI4lX2ZPR6s9eOS9dZ1qeuy131cxLlesOllynMUCe5DLfqYnqUqP2D
q47BT+Wnv/JruzzfH62hkZ2YhM3D0reBG1j+A+ZTLD4getRpXnMnva1NdYwPSlVx
AMCKglxHlTIJH9iSLbfDVzQE6whKRG3bVf7OorB2XPfNTsCJiMFS9ASTV0Zc7abK
QmkuwG/2mH3qd31Y02wqVH7IRNfu7zkzgdPG5Rv/dYGEUvEq1VWhM6vWWVkIgOha
4xhpi0RMfv8ZsQGM8qPvc/SA4WtHf2533meLhk//bFgI7/2Wg5qcRjpBauR5vupl
EzAe2bfIYk+1qv220VsG33IPCWjQc22mE2yVbsfomCSg/wF2NGCnNRU+lRHsIxne
MUNONC/5bX2GUMOfon/e5WtTkQTgaLP3pJB0S0cNRWng/T67HD3jye3ZXJzanPhc
ocHLZJl4j9qfpNnOLY5F/ZjjvL+o4JvjgrUlQVXwoPzX4sDPVL4S8ztlxzfPwuCO
kfG9iNklT3yvxmVErUC5j5l+Lwl/hDZCCyfnPGuvpQE1E3Esx75fK5Cic+jBix4a
EqYCBXDGC/PjuetGRZZkIzHf27+nYvm0tRAQ3BAI2vLYzUaf4fBXwyY2FPDkSx6n
VVnviqK/nKupiqa3R7P32CFBgxjfiK/o8AUCOG+cwErIZbWbHmeQCCwqoXxpi1I2
388cKT6MtCZepWnClDykaKPUoxEY8zOFZSPPNOD/KAsdrRx4lfrmgVNqXWFnFAAv
cwUAAjTpBdvA1jOz0/Rt/GvgcrExslChz0av2AhMuG1wrJvTG7sPLQ6hn6iun6Bc
yyQuvUnY1Py6BAzWac0DolryGwHlPekjgEVm7JQNliVakw9AjgXcWKf827aY+zH/
oLF2c1oSHlim4qqnJAVMLtacziGEIQVu2XpB+fnE8dfRkh0jMCewbDUnzzv1/oDt
ybZ5t86xADeP1DIYX7sgWmYHTBlH8zhDrcBHOLWDNU1XvOccetSRZwID+4sP2TB0
0102ZWZxlubd+rTTVX9JIU3pPysMOOHFS+JMCivwmWIAQjYC7LHCtZUItikaWDWl
emKzuoSnuhIwOIFxJEOw4pRbdB022cBAf0Tv6KzyR3xOXlWkVODo/tlhSgO9lk3a
R6FqOYp1t1S8Ylxednuzvf4B97pmNTQTCln/vzXo2BGtlA8N69tw64kVBg2ThSmR
lBPJEDa9/VgCuU50okIvgGIgitf4jnHun7B/RAbiac+4ooyjltCvKnIMQ5cdOF0F
Vh92V+oQox6bFZoU2xhVt+28SaeKhd5c09HZxxAr5u06iPGpDOuNNxgmB0kK41Qp
i7D2Rc/7sz+hKSAueNduQkkRoBhomvWQcR9+KpIrTm0EI8cFdFR8KlYvhpGJQeSZ
i5hsUIU1QodspDNzpePZ4XrKrs8FuSzLfhvhcFWPS+q/pAqRCkZqPUmY3z7HUCci
y+71IIae0W8mVTbCE2k60DIT/QvuwYUbA37ogwr7XMzykUmhf/s2u9Gah0qDFEcU
zsUBerucp3IoUB4a+ZgM0G9db7c9AvFgz3qYZrSSrxzUUOAz21Jv6CaiXBHwM163
51nm35kusS1C8kXolGzjVr0jkW1h2bZp+gHvPVaZg8tV9qdZT3Eq/MpWt9DgP98Y
rueznpegE3aPGKRfhVtrm5scxn7moF1YSCHzUZjHWgTrJ9NDJ5DUzqbSIIaH+TlF
Vfxh0FK5/Ev8Ew6LRftI0bY4TuFPFb5A8YhskkP3ZBDqMKxEa+LgeMJfTGmSjfuZ
1d+eNC5LlxgAyuzX+slDjLQ9+XK0LUeu8/wLlRlmnr95iaqETuU/xdPGrHJW07xa
fGPNqILtiiorIdV/NxYYlm00/iB/B9IaOB6jANWtBPTGXCYfn0js7ehFged6BRJZ
hUMbmKistIE4ssYNNcfxhC8iSnUyhR3H5LzFxIBzxNK6PoVROrQya054d0+fYokB
n6I9/ew4pXu9cYyoBJ41kc7CBp9cL2XaZAJ5OlkDeqYzEBnM1g2HIy9DOCtuyWsC
38Qn4MKQU9N4PPpFgMsE6u8Grr8kX1NxhmkA90lVU6hivQyUqoNjblAEJpTtr6II
mYfDUW/KH+TmgkXFh2/6rAdC5SEdTULt9auMkwDwL8ZF46Z/MtInc8F9b1p0tu4W
D20XgUQUbb0+PsOKeE81VFn3qja2IaZpuKdR6ZIv9yLP+6CSA/A9Jcq+DA8vAZ/H
iFGntbRMfhtMq5xhjIMwGl5ircxcEZc4zW+L9ZdF3ShPv8URd5iDbpRYed6VZt5Y
3ZVf1SR6Y1ZFAdCfIWT1ZWuhYGj5snIsryAhaIGLtTqqBiW0VC162LUii44xjpI+
6HeT3/yfDxoimApCj9mtENILn7JH/I4q/UQXAJCZu3uhOjCGJGiX0q1ipdxhDQ5D
Pad8rI1Lv2mUniupNgrUK6yj/KO8v3o47kChfn8ePrqhi8ghzki0AABq1mHYfV/4
vgp5Z0lotzkt+v2S/Ee6UpwIkUb5e0dKu5d+T0eEjCGUop2tZ2N9cLJKX0sAADFu
gqOBcsH+w9bmPUai9oRnBQMH+CZ4OqfI75J4fPjeo6p/vmdMNcr0BnDRHcTq8nXU
FUl6iTw0dIgucSNwDOZpAJUpZbr9CaThT+AcTPyEFLcj3k406tvb9KpamAAHRhzq
YSfZ/6rSW/hHyB+V0zU8M27u67EWNTj0KlJMIMDLkZgNLsPNBXLTlh4JeZkudQSZ
A+1QkaIvTBUosIuq0ph2jbV0sLzZ6zhEkb1Yebk2zA3R2zyOWlfy7PAoGqOvkvw0
fkDLHSnicOwrPCA9ZnP5argj5NeQKyJH382KgFY7LGW4W6LfYGHdj+Kl9TSJI6DE
EK58xJtLTOjGXXE2LoF7xnN0FMxu7u7H49dPk/ZIYLDeHk5Ez17ilrdHmZhPINbd
19Clu9sK1Dc3dMBA8uZ3AyxufkyQpw+Pf1EBYeX+Nr4tLC36JmJbxcYK8twgql+0
HUH+ZxNYgogMyQN9q9/7aEcJ6arjOmStfDEyYrodbNy0ZmLmd3ftIg5M6cgiexx+
1477IOHFMgwH4a/r006K9Ojw5Q5JPqRi4zXi3A2RMp9o8pdUvCCFiNmEfaNYfCE3
QJ/UNp9N91i+cZqU6HxzKX0q2wDhjJ92z8jNPvCsyiOgWARhaIQrYSRfBRkPXaCu
2ATRKvbMNOgxKBZvjNPGVlbDPB//0o7nYFubHOyFd5YwiE/t1vRmJr38J+c3OdMY
7B8v86bn8khthIPwqIjkgIUvOexIWRNo2L9Pgh5oqFOgq2PA8NItLSoNV16FR4MW
0a75RDIgVpvttfNFyvOTWT+L7r/LqJUoDB9fh0erVfp9abUwS6hv8+KTttGQ9Z2L
XP9lCsFlOjXuohTGTRnVZRpHWn5BG8rAjdJn3CBnodDBY3SKi00Tsl2byGcsXXcc
Ij8ySfOi3D5Iy1CZ6H6+mqJ0ExYh+eZcQOwii3jBDK0CVMRHMFAnx3pQ1wj9+1Gj
POIGT5nxjA4HsOGdP1jjxnuELQKcub9b6inJy0Juv9K3rrEiGH9IEqfeaXO2qmBE
+5EM4IXq6FbKyhG6KWb9y3ebAO33RVyKaEuTfYgMAa7jyZVfSULl0ZaGib4ecdXu
Tl/+FaFnnVpjOPXNv1i4BEiDfr36HLHpuetzjUnXtaPSHQr0X/VB410D3td72E8d
dtjEhb0D0fRqQOyyvWlesOyqp5pEqAqBeCZ7yvtysjdV8/W87Sw/ErPqLurmCjvx
0q3uQi+ZPX4DvEc+jQPP3Eng91yYkp0UUgQD7ujdD0ThY9X/yPKjWq1fM5/IItPT
B6sdXl09L6Wb6l3tIeAn6cEzBolXH2ESyUjuyalp8HAPjLysBDKQFukfBRj0ucC4
/KhiO9sEOUbM6it0c25lGr7cp13l40UHl2mXmv3OJQJ7SAkNLo1VCV97PIsx2znu
8fuSS06f4ltIzCLv114R21ngpYSWq0f1z2zBoKwq0Cu8kTmF480eefFwJad/vjaI
8gyKxjM68TqK9junjhynQ4OazJpX4LiKdqL3420kFXTkuatRxDLIFml7CG0mJGR3
IzGtyR2xHAsdjKRnvQcgEFENgx0mFnGcAmvSYri0a3x0HAZW3Yk30jlAQ7lszSVx
qzCrA4IRsyYnOwrT2CWseF3HA7jKyKb2/t9LrhjwijEjRBumZ6XVTb1Xubu7Nqo2
SlbC6d25BuGfI1cOyuI+V5wtIf8AdGLIJ6wadpZ8YpaFm9IcgxqEBBOjcLRFof3p
M/K42on4YhbYvRUy7/PlElrSr4tpTBoRCa6DrJV3mk8kAGo6jWLBOOG26xmZF68x
Cf7EzJyC/kBPZzAeVUAUjK2Yq60DBfRi38rHzm5KyD6z0TWWfelNfwsO2EE2baSR
lx7tP53LAi6zCCL1/hkH7sxqP46wDDfMBdZz0D53KO+3TkJnvq10TUjXFdeuOccR
PXP9/pRYA/iRt8xGXNmpppPfqsrMzKJzyetWZMjGR2m0yGzMqoj/pJzdTcJubvea
P5jZuSDKTP9HQWtj/CU55O6rKmHUJ1c4OVTl+vUkUZZWBB8/lZ9x4KsjX9jHYGUs
eWitqdPqfFbsz+aQB+LNVswsGrg0eLZvS1iGJBcKaegJXwUXzn8RTZ0ysvgeGh0D
HHa14vjTQyBX1E6/GQaZE3n4bKrCud1Oyga5TV74zqS2g51tKt3+queSTjTqjEDH
B9bAxH5r9qOkDxgDtz3q99SVPBmfIG5Mk97i//RsoF5JhBAF79RerAEAgYZ/E9oa
CWkQTGZfj/rz5DJQN2ARR1M+7yP+3OkTKmZ0kNUeB0u3obR0+Vfl7kEEKVGbQMgs
Q2XyBojRNMBBs7qi29KCX6QZh48KsUIuZ81NFDL2cGx51jBKkDL67NRfe4+EPYJw
C+GjjnEXnieZJxPQYxZ8FhUVU7ma1cnzV7fnB1lYj56XEznlQ+FjY8D2h086m8br
6iYr/fg937d0Vmbmhdy/8/gknfob7+xbMxUTCf44oeK3kyD88smQvgN0oCnhIQR9
xSVN/ybmZZuuER1JgTJfWb7Ug7O3cS6I4kyB8Hovb/rRFb1MyfBpM59FYsH28yDT
7n4pLfJWXdt8aj6l1JCLreSSjwKAFv5quHaTopDugXGPZke/6izxx1uUkLM+qPXH
9YKi9V9t0NERCtExiVZp30dPpl/7BWlJf4R5AjVHaA0YMwTrncbk4GU1Tjugra/f
3JiEmXSXqalNJVd1Qew7XpaYLGytDvms67J4CdVqHv+MW3V3LI+mJA8wM+Ocmx8m
Xd+fF2DmetnbNbiCqyb4CqZbWjQRIqI9dT6ia3alFzLxcxmqgnWCWnCBz7G442Gz
a+pUf9sP72I9NzTCi76VDfRNv0ipAVQj2BLgFICFkkj3oiRt6iO3qxm0Bf1yy21g
LC2TEmG/FyF/fJtUgVncxRUFNxAKZI34NtWnudAr99BCU9T56NMBbFNGNpO5Zly/
dfydK9cc0Y200ckFgO+VsjZ+mpIBI+oCW9xQbux7nj+x72Rdi+zOX1sbsX7WG3Im
QbRBTGeTgtv3dBEmIRX5Lo7dYW9nul0441CtHLh0X1HYdfVXA1+9OYoGpJQtLITL
bhu90q+C+R9leNcE5ngDPSnRd1UMB9X3A2oc589N6Gl7ywWzObHHm4v+7pD7MPMD
glWpYhji6NW6DXl5uzk7pwBH4FUCSVOyx4+CcqLOEGRfFegWybzsciGlFFSpXJo8
Koe/Jz00vo8XoSa+PHagHRx0uNveQgf8Jxve0iYc1cIsVtW4rLRvuMj2JkDICprW
U1L00lTqXijbIuvNhcx8YCYWgfv3DgEMRPOKdkfFa+fKjt3NlYoQZL5woVa3P8a2
zCG7gdN2CQtudGIDvUc5Rs+vucn0mlPgXNQ6HB3AeTpT2i7pwi6fwX5bkblphCUX
azxhtL7uAQKRq7LSgWQrJzktfXh/hFrJc78eD0NTuXFMudU5AbdC95Ba2CW31hvz
GhcCge3l7NSkKouMLcKOiOXuTmvOGZcjOvh42adKCH6vHZeK/DkYJjcRE6vIRyiQ
xwCchiKJZVnvgFSpiMrNPHg2l8UotZ6gnAPp8CsrGcen/W3Tnn0xA9LH/cYWsepV
4lGlE5V6Cn5Um8DweTd8DcGflDKGH/dPJWK9EDEkKcRBwc7XFegrmOxWixpW1R6g
+nTrHLLnMfpheDBa5+LGSI66i+LXnZ18wNloTi9j4zt+MIHJs36m2Sp7NddUbysT
lxY5WdtD1giDDNPMJvnTws2gmu2QpV2OeB4TQoXEkHLeEL/dNtsr3qT+p+Mca+t9
z6JoqZbYAVErb5Ka+k0pDU29RmfcWscxrBDaI9bx3m+6u340vLtkJIjrtcKFXQQT
JKxswGpxgQ64pXBG5BPiNSZlQJgWXGYByfSC7KkalYMG37qmFFGxhLkC/t0saAie
HqXs7elsxvYgBEXBk6It6Rz3R/SLyZwvZjWRI1aqdp2SlzZKTpAYjK8Q0JoZoQ9L
EcmBYXMS5aQJ3IsA/f2zkoYSw01TKY0QsaenAt9ygr3yfWwZOzI7piKmDARJFy2F
sUzI/O8pc9DHP+ac3sjO6vhaUn+VW3w7E4ljAKFNm9h2sWLui8I2xa3tV10uJNjs
Uep4qrnGnQmakzn17mw+r8/mAALFx2Un2CEHr5BMJ8lagQz322HwOVHFmb64GXpt
YXdRQs6aQ1mzJndQvcFH9oBzkigOse5U3BSmW/kO8rz2BE33X/4fP/xkw09MRAT2
nrJD4jGlgOT1JcDXtTWAq2kwlbKayNpXk3pLH0U1CxAN2MohlakJsjdmm3GhJpN/
UmuenAiNOSaUWWBWbcn02J/Eykuw6H1oVO6nclu+LVCm7+dEvTK+0L1xiBw0JFBk
vESprSarUOv15U2oNc8lMeXE1iYextuLrEV0bV5CicTIHLbkLyB3TdvIN9UDUdiO
Q0BqutEebNI/Q8Tfbi1H/aBThra+XcDZIOrFXHLMKMBuISmyw67xyX0ov48AB42d
T6d4QQ8Ga1bPnQZgQ4IYB8oibioN1MCth1R40toviQS9oJdtKtEEdwN1mP7k3ngI
Scbd7mFYD6B7iJzoJGvQkeCRvlwBZ1QZ7Lf65MgrPamTQqF53m59U9kZFgdXJCRF
98+7UPBdnidFUZt1fujfbHXafL1WmrD7RYYz9erDdTqyXVQHYIRK4o11E+8LtlTU
J/3n7RNuMkqJDTtRcdPDQW6Pr/RaMRgNPhTSVyWIwvFaRiGcFRRb+KgpyXpC7cjH
kygsnzWLf1CAQ5smxi5ljp1gbU1RRTutD7VDuXmnK0vj3lJQWeVCgmD83aqtWz6p
TCaMJU3UXH2SdoiZsVu6x05Kthh8mYNpDqcwLNqYui7E7LOVeAAkqGKhb7vTWTPr
368WOpLze2oAtoUSG78CrQqgkIcrgWekYi8VJVaaVO3icp6yVkFXdZnl1u4/8CIY
jVC399An6jjzcWRfaqoMCtVzQ0D/Xc6Zn8C5wcuPPADXplGKCJOouaI4NQIS5P16
0TMmQJ6JFvCRrStc/+xxKREyIO4yE76wCLtu4F4aZFBuc0QXj3dZbov6TX9qt2cf
N/Kec1V8lwF70jnykA43bJKOkmHF1oN+RfObVXP6UoRhYPhhAebVgMecLeODlQeA
dMbfQg4RdA84PzGdkjQj182EPP1D4if+SfWFdi7pgFDD3UtMez6HZKIbYnNbQbQ+
6MG3u++nIqnj/2SDzIt5RGmmsTGCKRHBa2twK2KEvU3vBsAf1CUbQc2hJZAOj3wQ
lyX7YLqKRjTicTXIHK2ptrvpl1JBgom7Q4VsQ5GQVUs/eXxbwQyW9KuP1s3VXRdV
KTJcunqYVGMsjVIDGXBMaSag3pDWMPisrX+eNX6Z2sHIS9RCdvft7Kg3cNMTSK4U
6tOKzW5ZU3IJbdWiPuLyhR4StuBS0gmhnHHv4N3lkZ/8rGKHqoT0LHGc1OWbLU3y
S2PWroUaemTLIYZZ/VurzvVP7blGIoYxVIY9MR2m9XQPToLP2BOd0fTiDknJohEe
AFPR2mCx2CqcBAOO8jVdIyXR0Bg7H8daCHum5PE/Mcs4z13HnWTk9NfXYGkksrNQ
ewY7OEx8ZTLJohCVLPWKlJrFpg8sS15/l+T6LQKpbxB0piDBQcMIOw50YThrAZAX
tijmpmCHEaT1snDAUwLrDyAgMNIr3Bq6SaCtWSWTXpPbQcqk6eDl3LJbmqOj7kHv
epw+9pXT/IaZs95ci9xVCK13VjikmgtxfYVKqhanyPTZrQKJhBiTmxu0BESc8hyT
2a9FQYwGUmlQ/T9PrzZjm4SRFeMVHUx9wOTpVTSwdR5cF3meQr05aCDRFsykVB8O
Ky9A7sHdbuQcaUVySukrxIkomVLaOU1c7yHWzztwXmGchHAkq13Ku7K+bq9o3d3x
KW3Ipufw+m1XYDWvIyDn3ZrKOh93PPHsqGCO01d8bfjT+Y3XkkESuAoaiDlxxQWv
qGlJ2feDmm/AQphbw3zmVc1N5gYipDIyFcQdbeELyJmkNO6EEYbbCw+E3PeIMznk
H1Qx86Nia2i3Y+kcho3rJP1TzNh+m44PwHmCHnTHJCu6CIiq6DMSi4qX+EWAvOjv
WcJlOLMj0y2pllspXl7/eYs1XMX8D9zpfOftk5GN048RRg28gbRRXRWn/M1Ok8KQ
CDVM1hjG1PLskcmONdlgh3Aa1rEbP3E3Ga758uB01sGFRvTVbZA7XHlMcUh6ZdPU
puBbw0QqtViYNgQMukupZhBlBXhT6qwkkG2eIkPmRzT8ayn/2whdkphyc489Z13Q
CE5oyaVSLoINgYcsVX+8e2luxL9MnPT1dzTH647h0qfuI7RpwQ8ChhUMZN54qFWg
rOdTCPoC6znBN4mpF4VtPeMruyX+aohnr8B+xLuSMUh5c8XGeZ2eZ/mpAJN1t80n
oLBF6kqebPy7CvHYXeEAnKoIEWkRNUc9pP1BAgXfo5L7lW1YMF0tpl3xRKqwmULj
klWRFO8FqzUFY6zTSCbkLZ2x95PbxEF7Pf5ETF6pcDl9kkKY3ykKNx1HFUQcnEFy
GXALHUYGr/j3qPEVmbXjY3tLmzVdSpibM8NqyoYRPirWKlCUG6GUFC46CKHl1FLl
fXf2I8zcljcekiMaPP/RXWDVs79Iqk0mkLmsqyQW6UsjLPOMQBtjhsXmRamRxv+w
4PjrrHfdYzPoxRQhNoT0z3hmr4iX0lUqsU4ay8f/m6g3CvL2pHocVb62JOIv2GOj
vzU2PRtB67bRT2peRZeZtgnvgJSBIfzZtWQKAB1Ni0TVb6plByXI5OOxW9f5tlCI
A7T1M+YJvtTR+d3rz7pFCq07r4J+zTGZ+bUL8ePozwTqc1f4cIvhPMmxgYWAm2Z8
g0aL4unt9Njk/It+A1i8oI50LzghRFPuZeu25wtUq2SvJ5Zkw8mnyi4pOy98IGcu
Qq8JWmCRGiMKkagd4x4jCoYWXss5UaccHVxXs19JDNufFJPz8YrLEUTj3w5g6lpq
ur1E6v4e/LVHraGA+IVi8R2Jr6Jx17/F1pPr882lPXK18OtzMCFB0fhzUOAfMaMd
bPemZhcIq90oyXdKnngLJxzckgoqY7LlchcHj6V/4LYf0k6fUSBX1+/90ZNqXHtf
DtCryXJaRrQYkfpEXFb2A8EcNiCjzGGvWth6J9xPEliTm5QFhAb0OckOOcw3KYEp
ZGjovTl7HR3UiVsnPChGhPnSVf+ABsB9dyqf7Newd50xBaiHnEQ2d8xVq/Wnd6ao
nUGTLbYR/Jij8F/wfoFFiIf/gWldOXGjPdKP00JZSSV/fWyAnjEqpBaMZszUYNuQ
l34sRkyjeEQ9+IiaZ1R0nfdNSEmddMl2lwV81QBqd96o87itMf+kjSDCbAand442
owksdTbkj+rOwq+T+BsExNnUERHXkWJIpKVa1RGuBQyHWQUxBW77bcVSTPIcAxPl
dQzjPC9uWAdU3PXj+huJ/QutUG61kkPxJtv4H4S9uypoNSfKpUTikK5cCk/RWQa5
eeNY5baRP5A9B4PCdhQHFtQ7KF3ux7nePt9gMxHk77FVoHl49kAvLj3gGWXtrqXl
I0Eo/uaVuAJp/Fy16saaYuUU+YRY1zKwIOf6eEKBjTzLOrUDYHsC9OmzYmSqTyHl
7DQ2KgpijCkhC8sh7sdvTB/0OPY8d+0N+Ng7GZeWc98E2Bq3frFg5s9IQe49gHMf
AXiYK6TIBa8yujewY028EO1sAXtb9WlBiNsz6PmOKs7v1xmvMHeiEvjM70bJZVqk
rbbPul09o2hUlsKAUbhV/NB0outKVSqIli7snyfnJ3PNmhT/wpIiiIA8gXTR5IkT
1xUoD0QAOTV86B1nF3asQ89hdLB0V/47vvQJS+J9mZoJuQClPim09j5Ct3zQTjAp
QYRbPd6bp5lVxFMnoLS9LLl+SEiqu1W1EHOh4m6MmRey5tEv9ZCsbFk+cmp5s64l
12VOuYQYZblRzfCXGk4uxM1AAmw/hRJpw8rY9vZ2p6iedmtSXDYAk3owfgVqVtBW
KMTuVSUpqLKhy/L2Whti19IpDxN1kA2Hmt7nCoJJikz6tdyhgA4oFJ6fjzrkSgBe
HI1ig7lEEhMNed+HMckoAcGeD+1qJCTMPmLf8Omx25baJb0K3IMCdeV5aAfgoSLb
UygJAVO1EkDl1d7wrEbFUon7Ehlmac5Y8IvtELZYGKDIFv7inHPCe+/9YK4wWFaU
9btzsQWsSUu0W4aOa9v2hPtsNim30dZQMAJrAIgBEQdFKt8RDmsbKT7Hzw/+URSl
L8CDvEKPeHAVXaBg0gYpX6c/T/vk7bTPcKKD7UzsKZfMXGYtmBj6LvVr5BbtmRJY
Y3iKYbemJ3v1/rZmFmzjfWXcpqlaDC0M7hm94aRGAzHo89a58nI9+FF07hrUAya4
Nkzt0W7soc0nyXT32TZgFzLchYWzGqemsq9TC4FTiWQP6ftudG1Fby+WmRrcy8Mu
rIciFZPu4tsxSA4AR3bUTXqqT42yaFLh3PG8naZhc6bzEfjd2ud7vhC7hLn6NSHi
BsJq/tvs796oPUOLsXEdyTZrXLgSnIHyAEgJokAz5RaQAQLeetFRTo+ZJ79tJntb
uSqypb6Jrq3vyRb1TcmJlU2XEUJk+SL9cAQaZ0PQ5h7HAN+/keUxFDxA/wCLy0Na
419E8D7qAT8+Mp/U49h4RbDYNmHlRJZpi0Aju8T6EUt1csgNJMMtxWIU9oTe195g
hxgKQpEHfj8aIlDuRdEKDZiefpPm6SHjxKxCl99ntRLZ1x4QwGslQ4nXhYNFzYxc
TUvJr6nfu4d+FK+U+mmti9t4JyybQgNgB7IO71iDnDeNdnGKTNpWZEmfYTJHVY6y
mFstJAdiSBoBMr8xhG5E0tx6IQ55j5pMgegqmrQYE/ufFLcpf6TAwWqaMxS86Txw
nn5JGB2cu2wE9YRlDtThBRbTpv0h+98t67nH8rnxaVQ11dD30IwaoOq49r9djVQV
s72Oo5e+TwR691RLyflq4tssCZ0GFmxVulj1coUjMSCRa0fv2gjdn07GQZujlo0Y
5VWaDYde53TvTYO4DmScWrHcztfAqo89P8DKrL2ehO7F63YK/l4nmMeaKQuNmi9T
Scpd3Y2hgR2FOKZDeKigHnvC73dMt/w+2u8GfluFMP+ttmQYf7iSv1gvtjlObMs3
aIQCRtGPsHi94d76g6WflreDYQPxek1JMpnG64N/QwDRTIwgBhJyLJt/8sa7UCCj
j7EPUduByVKF1vwEcq2zMOyLP3a4TTzWGGT5OWKYO6rlfYPd42oPAwtcTces5RT3
VS/lq46mjzORITQgu8wUtPUT40J0BozAIFaOjGlbmjMbpcvrDE4aNQYH8PolY70v
ggatM9d7RUi/fJrgsdLSUGlmyNYr85V0WRsc+Pu7npRlGHt96pD3/4hXTt2rJ9ig
BTAtPOQ3P2cgJ0eEAgeyP7WSu7qsSCYwWacfP7O1ZFfdMY1vf3UsURiQU0sVG7Ju
XJN+R4clXaWvhjve2iMCbhEIfOZle00tqXs4+zvAkQk9f8jUjpUlrlL0C67xKtES
DBEll3Aa9lSAEIiTo8/Zax5vGM/Mbn0meDK9ynTaz938HMdHCuXSh8XKKZ3DsgcT
dCUcCCYC6CrLNFBC2id/yz0oN6Pgjyfv7qyUCwE9oAFGyRQDyHCS4axW+iw0RlUg
8GRNuHfa+v7VMLxNjTFMf5Z/I4yOD3bUtmooDaAoVYmc3hlh5OyLVCO5DTB9Td1I
sISXgtFyxKSklQNN7gc8z/EyEgra0cYb5w+QNKNW4jGiWxzliIs84IzUB/EXqiOw
zImDCSkwSsBWwA+oURXnRDtSvr3Jk77TbrGbnmmYU/qvJLz9lKnwXQnS9x6TzBo1
T/Bihy/dQ0pqGRajh4HCXrkCTXgGA7hmO2S1XHGPRkSDzy+w2Wm3lchYvfywGAZc
22DgWv6fmwgqKyBWJe0AFVVQAxi4B2sobKmn8PcfEUKhLVci2VZiLJzwSdYdA5eL
xNFW9TXN9SiJJPN7QmwDyEd3y85SZrS8UFTBHRq12ZWbu8fj0MoORBiaixlV3eXZ
MemUS5eAmBIpzCqtXlpuKZ57ijBIl8qsb4kgGEJL03BakWw9tpFqDcyyGAypj6vD
Tfw7QM4rj642UCPvFHZ2HO+tkJoUEEO+cbfR6eO0RrhuDmjlJ1aDU4INqRSmW5EX
0mAYDemLY13hW88ScTljMtRNj9fcYri0+oJJejhZO583VuL5XxtUxVDxWktXi/Zz
+IPKChHqT6SZ3err/iY678Z5U83smitdAMR7pXF5vS409OEt+GvCmi9I2FQrAEbw
yb3fMy9BucwXVKHpdT8e+woQk0BDK5TzhIAtMCkrsQ1fwxRHhbm49XGoNenbcoiw
ekPKQ4kV85Yd+mQhn8el/BM1OgTiIJ4BdYiYiVt7gDYYCLlA/dQHRqYu6mGlTH/x
1DooN7t5FUOch+rejX9bMZcH5vVWqXpJ8YJKqJizq3e9t3UShVn8czAMk63Bo/f5
fR4DmtY7Avx20JLlhFf3as8vQvC09HgNmSVdokxBY7chX3H03HgamcBhLpT9LiDJ
kFuHqxtMPcUuBecyt+ekYJEJnQJSqaHI+6OylfYi/uQJsvQ6Sh/x46TwBr0QC2ut
4MKDt98+b6gECp4niGwgwlCf6AKwBvOCvSw2E71755tGLPhCVMKdLyARTCw2uXtp
zlDZRDTHTKeNkuf0s6di7iEuQN3P3V1gKG5kbKag7JUk5YMWwRgBqbzvHIs4lzZc
Ih0/t9g8TVdF//JV10S0qFuUnc/Qa9iQ2TzZAG5E+MkcrUaA9NJ4bNlyp007v9BQ
Rd8EOB/aIF41xmY+9auGHcqMOVidOnw7slZuVc4dOhc+qRVX1U0jcAKFbi8XRd4s
y7jb5EdALQDQ6NqcR2y6C82U8g3aJinyGTNEglRssDMKWoOUmFaiaEuFHJeH7XEN
JPaqw4YbYRKJZeeZ6anqWLpLA3kRwsJFPpDf0v4EBCi88fE6COXRSLYnw6wSW/fA
iMJHOupN3xbC0425DqLSXHp5B2Vv2NHmAaTxon/toTYZfUmEMDWxk5G8XMUdQoGa
8dmopbekW5fUCIPIMYRik6uJk7HybyIP52z3gG+noPp7qaB5EGVv7Ou/1+QvGg0j
A6eXt33U1rrluX8uKic3DAc3Xur3T7V46oIKLkuSg2Y4MwxorxEH97TX2T1I1HFr
Dr15adQtyXB67zQzd3MX3lF/TMcxgwbXdZwcK5o3ak6ZpQ0wZqaK3zL7f9V3g1yU
zG0hk82f4rhw8tiEPuRt4K69yZqxBwN0SYnSyLn9rdiR4bGMaoXKKjkD4uxSx02/
6PjB1ujiYzIk6zIR92TGL4vTAdALJgt95pAoq35h6VZ0V0+hbTvWD1QlEsj2wmqw
/+ucJCFzoPVi6ZBTgbcmtYch4yXGwvo1MrINHJbhsGZbGcMFjJ1gJPtZ9YZWPpnT
GW05Mjf18WNsFewZyowf0kTId9Hdsn0M9Sfn3IID7yRzci94VoWB2pQDlO+LBrA/
lM3gPk7uhU7dMCVdq2UzyJ9gTiRjsIcov1FJXhUJqFSUnhVdKJlK3L62mifbxXc9
3qLbt5+Ncv3o/BLEIlV6SXiVKDmTimu6+C7FFpioUax7LQjoA5A2tPOqZs13IsSX
gaJtMmT5hC8nXO1Z6eabhcdvOqHdtVzlyJtfNC5PruCTNYGCdvqWc5KpP9JWK/IC
YZZoE7sgGu9Xu4V9NJZztyOC8fLqwpdstn5+R75RcwrEsdU3x26ExwMtEiQQ3cTM
MbG5QwQyZGLQ9fRwQoc1zOfeTemMiI15JUWmGTF+2mS2s9UBLtUTZzZSblO7hU1g
eK+avO/yKJDAjutuBsxcOlo2GYkmY7OUkz4+82HSCPfZ2BzrYq0M889fhHYKUsCR
yrKzZ7/EeEM8cavQJxqFtIUw1v7cU2J9bLolzkN8bTe9a0ADyBa8ndrex/omNDvR
gy2hzsRIdveX16so0fv8TqFXkLOrSf6CIho4bbVbToXSxHKLgzyH7LZdkWFJr3Yv
IDm0NXv/8+tahvc7EXjTQxc4IvoNhAQan0a1oWKe3JNU78g+bCqewh/XY2uf0ust
weps1HpoSJsusqh1oygU+4WJOldzRWz8h30NHhpHfvMkaUJHSzaQnA28igXvZV4g
Rsq9mEwmN6tuvlvk3/uYRPctMXTsGqZQA/l9/vuz9NB0wVUPUEgzAAskGuynZ6ts
+8bCdnKAmISexwuFXg4i9EQLo9++oaNfpE6jhQJiB64n9r7yS984l56tUAkGcPvw
39+vlfWpltn6UnLnLzJUdUvgImpYhO8qQOThjaI3sKDnhKznM/Q0O0KiTOb8bajb
UXPy13ztj8S8NwfnbQVyKbjUjCHeXLFr4PcLkvKG+YNBsoIPCElo3Ts7wdj0QUrb
wAEJvhUhc2+cGvVgaXREFHsJGopM8X2XpfApEnVu8BzT/sffwNQJnX4ipj+HZ+Q8
MgIJeLEYV/mRAA70O2OYFHrO4qSsGQoMEuetRqA+/GsanULcHRiF/q+rVw+wvnwQ
Q7ehlJjxxzRcz50KwJzQ1pETJVb7LA6E25l1+lZ4E+iBtQVfYWAlGWk0vIb64cVm
dbVCwSNEIUu4JNUn3XemtgKOCaJFOK04XD2lGhty+hD3sCjITPqoY9VPtR0lNlf6
O9Wn+cfG86nxUcHmcd92s8l4nShyTp4b9endSQdKpbOs09s/mEVj+Ssg9ggC+Wgp
YEGrR3bc/x2Da25HXciMo0GDwhS6QyTfaYsYgbUcDTkjl+P/wAbtzEnkAr6vTZqf
z5eV9ce+EWKYR8VbEeKb7ArH33Ut9h2OlffRHSZkGVLNU5grienTEJomfmUr5E2o
iZGaDF7oaVwRYvtZj8C2dGmuMJWslmhX/+1Qg6JEBIisJsgclrs/7U4jIQ16p1Az
MYrTNGab2Bj+dBy+2lGkiksmYwKL9egP2EN7MoNqCM6MrC7WgDdAyAb6wHa+oBrV
p80ntKSIExn1kbI8cp9UZVvK/S0lQE/ctbmQPCzmud/LUF1Vi8tsysm8JH12ACJ/
B46KdrXIKejs6v+4iSBaQuxUb9L/9hQoh/tUWdI5H1qwZbBsbVEIDRys1N2KsfvW
41PPvNVkYATo3CgXefoScFItzGdKKR6Jai7Nx0hdTnlzi2is9+fwejLaMN4PMr3D
t2SAik0ZhQlzGS+bcDXhwxrtIaCC7PfE0UdnUF+N+rr/NaIIcnmYaLxq/l1cqiKx
NtLuvBG0PoPGqWG+wEufj0ZWD5REaoYVdsBLCFZ5pPT0gL6TChgEJcq5nOn0VYg3
WHCtVA5Ub5fG3mpQc10tMzC9BpMs3sPEmy6C2vHee2VSGuF1PNq333rhESD4GCK4
d7Hi6nJCPBFDBrnpjZaSvEKWHMNgEVKOwQSpbbjR4HIEfgr2Je2lQ1JXwlYXjiQ8
iwkitzfAjmTXO+Dgt5bsI7kHQNRKV+GmXC2ckoZC6Ix9aUn0Shu78rAVFfuQWnR9
IipRnuzamZcJbAOuSX1j253z3xLgcqyeOg3qUVY3b3q7lMrWK3W9ap/udLw46BUq
rZbtvWYDviUPSppJMTcletEFThwj+FbycGO1KwedZAh/wjHr8IT5lnEVCEhvbdyB
OARm0k2w9e+DXJMTWiIePpSV6NSWVzSYzPI3MiQeyYI/4b5sUYBAU74kVpp8U17Y
FTCCBu6/MyVAwdlJW92hHvNQBQEs1NQ0LiX8ugh2e+Pjz9tjo3HoCCyz2TKOZ2er
d4IKLuybLbuhuUVy0IvcFeJWV3e9awK56O8QGu1Mh1NpresO/o+n5HRL8+voQ9c6
IzLB1nPyR7uIWnZtzzKk5V6RL1TFEDAZdc4iJHt5HEjLPk3tebY35agclplFnXFu
yeO/FGSv/x3Rldr3cLDHpx9y8y4TS3Kar8o9kwIkj8r0qTz7bCDvYyxejVZQ5uUs
zzn579HKioXTGRvC6SCcti9qv8GjXcxd9Qc8WeicinaMTuL/+4EfyQQTQ5bbdd1/
gMpOlKVyQvEwxFWFdzr7+3PXOFdEyq+pjmHAyCmoGOUi9uwAT2QPYdUcuTpGr5Gd
/kjfIqsNyNz7tMDN9VgkCN56XEGdakq94NNA8YM0R/GCXXYSSflIVre9m6PmFqON
OZGDX+hP1BxKZM7p+a6eyvkgGF5AXL372IcvRG9e6kIDlaDpKKLeivtPO6TQCJQn
wQzG/zTAh/gZ9g23z2yjTduFgVunqAzPg6uxrTzh7fZQns9h9707/Hx5vegJ45Y3
cIcHThMoKjbDD/oT1ux4enUftSvomd5QcAuePO2qtDRzynIa8EL9JbM757LAy7v6
e998nRBc5xZbmJhS2h3xfw0R0LULFInR5iG4ZflB3CXLdoShJZQ2Xgc1+9O0XF3M
1wTv15mQ6UJtSXby1Z5jfrFlPH4AfP/0IERTYncoOKJdNLH/pbjdwZVCe6K9EWW7
fINTA+PtDIjtvHvY6/SNXMU1YT1pdCGrrtInsOq9ZXNFhMmV0Tgyf9vbDzk/rL5/
IK/EcL0dxOqiIp+UmDbHXMzQL4VXTLO2Sy29ITvzUiqMm7f22BcYCCp+XGATnkcq
t3wNyOLUISdUtMsCmDNcCLz3eP5edDPJpIIYqs6KpU85X1TJcEse8NxaJXqbsVID
ys25/0keGaAyXXvxhu3Z8Yi7v71bjLQjQK0zUaZcK3lwrZ2WD1kgSqV9jH8USh+n
JIFOU4x0Zl8gISQth3f0LVQOK3CgNHR7lGDejj/PGmdK+xNpos+EHLrscz0XqPTk
9o1UgyQ9cQDWqy1+z18UnLDTVObiTmflmVhk+1SS05kYWBgFnJHfQ/HuWo8Sp5uL
YI0LEzaZ1+DMx/lTrnJsKHYML+BcCCglgllDMSOpXivCNGnOqalKE/7hJQdnSKXu
yx1pOTg1oLEjWwy1ti3iSBi9Ee56ULQAaUOT4i65EaX3yL8l7UANUxoTLJlQJBPO
NJXCHrc3t//rJTO8Jl8IA9lVY29xDRl/PDRceQ3kNVWcpE8Rs5IT70Xv6AGnTJ0w
uqTbl+QDjHxt2RDq9iuE6Su9QvOA8w54bjV1DE0iHYHKvct7ih6rGQ3q/YdDhWeC
o2GnwWG8L93OIRAalAdbNjvbi8c2xEjtHo+SKPm1JZQC6cs74TD2TB7DK1ikVkyo
MNhik/i/ly+0e1DATG0R/jbNV2eErnauwklrahzr6/ZtEkkj1iKgBbkxJ4U+wWjI
1rtkMq+NgqxAPyybRWfy3AQJBzN8oF6ZgHvWq0LK+Aw61g1nGRcZ3R5O/hu9i06h
seb0CzK1exSBAeYvF5aVSN+k1E0eK/qJ3etLVtLNqwFLRkdn+/pUBLKQoyCEdSyv
BZNvRRVZ9gbwC5l6tC6vD8sqCmRGaVJcUUv6ut1XgZ+5n5zUwwj7xr6qAdfN3thd
GBISO1QNFhSZrk4Qz3cGHoIqi7gTQDilM8o8OIrk753Fxt8LacG+1YsvdyoLoWtZ
hStR+nClHJd4Lvpu7yzcwj2zibQHpIB9DeC8LGjGfJBMeLYDbYrsyl1ciUgsrIdB
L3vsJXDA5MVLdDRhNbkhKH3X82f2XIs6uOXDvZKc/sDULKd5VM9Q3SER5ttwxpAS
AfEbdXiiZEUS3q3MrLCR4+pFy6Yt7VBi1Y+CtTIWEaENet51kl/WxHHGNkWgRhaS
ym54kDjcmxd8XvTmA6CPJBC+EH9LPkrttnR4U9E+vJ/+kAhx6e9zvaj/3wt/EVdt
qmsWnp++i7chIYzTOS/attBhX5CRDSSigVpF/gb2rxbNDRBAax5xnT8Tw9uFQylS
FO0Y+owFlem8F47ZlgI/kmSJRpu7Gxi3uznWykJs6JArOFL/NV2x2Hb2g9JNwBRw
Abp2QivyDUSegrhoo+nHs9rTYhwfxZy9ufgqiO5xIuWam5M7sYepGtxnKeZF9EzZ
fwD5PdYaP65Ai61wVKIGCSS1I/nG3oOAE+mFDq9ELxfNs+IHm6zID1mieJ/JLyos
DDUF4nuugbamRrSSy44A9fa4PvfHos0Yfh+uWyg3EzYtZ8yby/pWVN9BZZi3bKfp
+9UwRGVKkysleMctWV3qWe0wUYa4IHY7TXwql6nTFLuWoa8yPrM+keMAPJSz4l7d
132csVp7gpJHrWHW5KQD+Skte5Zhxueehyauyep8zNhmloHNeV04eVXcTBxCzEC+
vWHPfrC4ReZ139OgXeCrOIuYW0avW3S6vAo1YPilUz0SlrvZeo5rzKi5UUo2X1J8
ZnEZAz8Fh7N4a1M76hpxe+GoaHkWfmG+Zojb3amie5RaGD2c1o1T66IDzhf/ydfA
8pbeeRKRKgJiPAPnYiyWrEEG0HcW6rWy7MO3ddrdU79W2s+J9sQPn5ILbCJptyPM
64kKS1Z41yVu7dhcuPM00sESqGLfkSyATTP21R4C5G/I1HbHV1t8+NAGzoKjDZLp
b8CnA6FnizmKiOrz/Mz6eLSlLefKhmC7PkN+miIS7eZMM4Ygr40V8hCbvQx48YjN
oAbmtBJY7jby6mRwF7Ros0Tt01D2dJvoo0PPbMAryYI2rp1XR0g+10RHAk0Fg75z
W5lSH2vnuZge2fvIM/GLdZOGB91Whxr4UtJiAP18SQNLTjZml3f52wEc8D67SVN8
wBJ1J2x2l7Cgw5nb7A+aBrlEQL/Cc7NntwfbrgQaD3Yiy5sJudGFkNHEDB4KgToI
ZNa8uXwntqO0HGOiuxwjWz83uHjWYJ/UPyzWaFsxKEJMZtqAyJ2KQRlz0H6i32kI
63Zt1Mt7J1meMhXODnWVdcQmUuqeIXr4WUE2SGBPXZrd4nqGM5yIi9QrQTypY47S
4Uwsuvtx1lHeSjgXNxaOjxEziVuOW1MigH/89Jgvew0F77cHnqvWE2YK8cWAdp+n
TFbDVxOrR4RdeF6bLQ2nhnYvXvCi5yUk1sxwFLFQPs/gEWu0Zpb2tYbGJDwOkk1v
EZS+2yjl09fOZfHEJM6BVEmnT7+6tKjkpT4Uf4N+Y87AG8bEf62FvvmHi4n39reE
Oo0Fmu3K0pIMnxzqmfehMbJEIrehGv7Jshq5tZRRzlXxl1+P4LajfEgAGy+vhrMk
7IOBfwQq4aSTKRwmkIpY00JMAz7WYiCqJyvJgfOpjBBX01mQIzWfAq0vSb0OwChP
JHZKPGCZon7e/abGCuKneYHfwgET4Od73VWs5zyIK5LjAy9eOXtSVbEXGuoPksNY
pjCBI9Cde+bqtK/YDm9NBQNJKsNBkIx4HuW+2dyE+Nr/QQhZaNxgVE0v5fPwie+C
WQsmIQD27/oW4V+TVvuCPg9VAcmSZNBxtyF3sgowmpo1z6GfnLDFre4b+I9OsL57
6vYQ3A4mJMym88+CSoSXnu5jBFyCCkaoDfsQwlTWIgImRNWpe2FexSl8PCKiasby
ukq1Z046a2pKc0sL3LPlCMO1dG/gK8M+1xemQbYSlmMHSwAgFwl/uIjJKKGVgG+i
s13YXIOOk9JM4B89mgjcblpRCvw1YHjwF++meRQp2NBe/S7r0jukXlNMCL3TXrCr
5+HtqYJ1iG81EBu7FLdE7xnEFvKgPtya4FAxeseTLdDF0Wv0X2HGpSep29HQdIi2
UX4fhTt/l+MjPTjYor9Bet6Bfk5O285QbgiyAiV9HMmOP1siFJ/X2X8zUUL/rvai
a7xsTzk8ZsEz1a1xVtfG8KJLln+4w0kQCmv4PkQu1TMcyGAPM/89wW3VQBxRlwCa
ZkQ1hiBVyd2pbjyGxiNPAaeTczWzyEle5MFWjdSg18O4ClxhAZwkuTsvekvL+Dq2
Wwj2UpPc/lgE7E6H/hiBBAi95MieaThT9pQp/8JdVAiB11+Ea3fDhM0oOHQ6r3+b
rHvV9Nd1yKlBcoHTGLG/xEmgDI0fUwfB5lFUN//gDKIWyYic/mnmdsX6rTnBavJa
UcihSQ2SuvmpPIJcHiY02HRhaVP7bXRBEt94aE5zAkaRB4ew1dpnnTu1X+rQF3v2
/ciWz9SEyk6qEIdoCvI1jLf/vynTAoAXOftKOzw1ItGyhK8+KMGOglmB2FnQ/QwJ
BnCDY47I1GqFkItdZ0Nvmlikr6SnDmGYxCkZfjCSjVW2usugE9bMioidmfVoaghO
Tyr1gT2ro7Gi/cEqehPSeVnwjWdtFCr4SU8WoaAtJiPjxPmsJ953o7sZ1vZQFBnQ
IYeHCv6vmcsCJJENFaNjHnZ9Q9qSH4aqDP58YYjWczuuZ/JlBGEulSIoZi6Dvh5k
/7+P0csG+IV0rFYAh5sbIayV3GjP17d4JwEpZ/k/k26o7PWnW5rb/zN/LcXhclla
yxxxb0i5E7N6KGRWZi+vAAhBZ6PW4Ym2HLoAM4OemuThXe25aeGgka0MAn04Qt4D
XzDqQxn6KH0cyrTVPxzigbgbtrqvleUTtvGbMHa3Noxv/uvtm1xiFSGFuCx2/Ws2
ROvS1JjylVRVZmJOLfID4ew0/1yz+9HD3/1hMJiT3qYEBcr/UU8iK2BN/kY71iaB
B52mQ7qgcoscVn+UHGZmXedN9HQeQHDuLA7SBOJnfdLjWjIM1XhK9D5PQsjcLJ0i
0iiu6tBb+11+yYCANCLVfQ1xZ5xuY4Pyq1fRSXUoVhuLy5+C1LO237ZSCcTjLunH
Mrjvs5hoOn1X+e3H/be5sjDF2aTpsSDwFbWsse2erV3A0uXljOS/aEkIy1Jj9w3S
NuaUijOxH/OFZQpymo+s4r2Lat9TXa276mBf8Vy5iVpGnQbc2ctAA5l0dSlu0L9e
3/HZT+7BFBXvllDb4NJgtNqrSt6ANr5ynVcNBMuFWJ+YxnpZwlP8m8guLkYPA8xD
N+fTWGHHKSLh87r+ySDJfrW+x2vMZXHyQch0d7QABNna4FkC11s4IuiFdCR8od/J
uf4svRgiD4o6LnyzE53RTcCHKP326hKAM237WPBWlbLLX4P25kVUk98faU5AXAah
obpizIC4W68tpfiaCI1bugM6bKZmovyUkxd1gICnjuzIVAvC/NDslqcbuif6xpLU
Dqvan3MlD7I91y2KeMplOQgeyXxI172icpcq8uqd4werl0NBETwxelOE7kf4Mr/r
TgouHTRmHJV/FgRZpMRw8lfTfWv7i6cVXYFShcqc6VWD95Unp+riUgi6hW7EGJWz
W3HPyU5b0ttvPSjkM6pYZoMSq0EDA2Bhn4zq93rOta7+5pjv4z6/h5BnFqamTzHB
B2pkUDejDR6zrigTadq5Mufe20g7FK14/hC5fi8l9WrRU8KiZUbTw8O2QilFB/fc
wmBga0T+62/28hgn4t2nskCXIccFpXm+N+rDoj3HiH1qYyoepY05F6Mhpt2FZqdD
UgYXEaZn5YcyyEhaI0V2h5KZ9JqaD/O7xzOhCW9Uu7e14KPg+MISmcQpEQii6YdT
IuiCzeN9kRBR6OQ+1/xCiRDTzeuvfamB07/UN0bQr/Pn89brFPKrr3NGOgfW0WcW
iTxxMqJFqxX0NkZvYEjtL5lofTO5/xgSm41GfpXo6VuF6/XBSpkrKsYkVTQQ8kZZ
MZl0re75Cd6HI4eS1H4iThFqTNVM1a9LuvuK8eo1WHOcAaYR+t/JDBZXi4Aqaxnk
5S2s8kguKhlkAvTSlqSrCQTvDqPNjzEL9uqr4Z1aDwKIAGdF53U2kyb7muMBjk0L
LLCjqVt3Ayse/5VQtAC1J157RyZBR7c0YrD5kgTk1fO5/V2lonFV6BdZTzO20YpN
Q3+VELaARhSPmmoR7PRsvOIqLBpCP9idNyMnJVoxCe4+2y1zJkRdTA6RcPRxAjxj
2rbyFw3B+0460HgWBpacNEyW85YQMM5XEwzU/pLeexbGI5dIrbkmyHqyCf/hwapF
pqlvCRDivyrTBJm7Z+xCzJhM5akmysqrUTuzWOi05QrIifQf/SelpMkd+8J8qY1m
VI9/PNLPtlk3OBqQM4r9xo777NgYDpmJmA08c58VJpLvCU7Zpnm8cwWuqYrZMdBz
pv/SgPlnex91HnMtEzJUzJnjxqSEG0VQUle7N6+kTJOnZsuvBrGj5Mg/hFoE6eEU
M4DumJJJke+pu+yMJyxuoM2caYx0kdaorFbMwLakvyn5ilxxwm/nEdq25R8oUsa2
Ec9p6hM9fKLbGUZR0VjX0EAJbk5vlNweTcPbPpYii+KRrLpVQBOm5kZcQeG3RZkR
i39cPJDHpuwqp19J9VqqHKK/Nej5cx1EFfNNbK21fNCMSViWFqgbecR7SJ4fO4zV
bQVl8Fcndh9GMOsqCoryJf30P2Wz1kkz6xU43s7+Zv4fWVs1E8RMl0YDAxl99aw1
hHUtF+t3LrXJ/ICyJgKYuCKIZTbwn1nLSpO0n+pThGx8IguRzkcfoncKnlfT3+KU
MNKcuJo8U2XSyxUaAd2KupWWiMOf/bMA/Kkbo1QrrkLHnnuiql3Gipb4f9zTus8r
fjD7jx2hRDjjIvSBvqyydmHuXhwIeFVvrHA8JRLjj1t8mnW7plECdhfh9gij7m4V
vkLHZ0Qbx27EsA0Je4pKWgkYdikSwT/5xXFvh6TCBYupROjEDYXc8cNsEvbk37yK
SK9I45cpAT0m7UPPk4Eb0jSUFM+hVoEWBBd3qk/7F2HPjq7GLB6kezMJU0k3dJZo
fC+Bmf47+6uyWCcf1uIp1kl0UdWxamyUU4C5HsoaglBGns04V6rkf1Ro8StlYhbn
7Lz/ypFiZeaqFLlzj31HiH4bI6O+hX0DQEXK8GhZ0q/la7bO/B/ZmAyUV3JtYU/V
cJE8/VvWd9Bbhegd3Lu/kuWswjwIJEwVnQC3lob7bKUFlHNkoVq/kUmMTrdzwojr
tG7lbc/pygv1w/Zcqchpy1/B4muntGJWaowZXpe7EEDIXg51a2zRo5MOkVHC5rv/
2j336MCYKMq2NIUiUIcQ/3EX5J6Y5kgudIjj1e2vKGptAM1QQtnysCoYIznMAkhX
gjEvzSMNLHC4GJ3Vv+1lJAIzAid3O4k2dvIJgoaFhPIXcZuKH43YozHzY19dmWm7
NvaN/0W7TYijQIDpibBB8UadXAq4SPNNt//LbAZgUtPJqiBiKb2L6o5wIAFPB/Il
uITBVePMGryIrcBg5EKuUj+/aKIcCjvCuFzNGl3bkhzDTYzPBboaAqqQKiEMFgpg
0HvxPIXOA6vanYNyZIrfrfOe7IcpH2BCSfh0wZX11L1WljPpcr1SYgO45Y7n55OE
2lYUbthVdsn6CTSrpuO5zMf/JRKPlbIVM/F39BBDhJJAbpYXEs2YUL4xiF3eXvhu
XyhQe9j+qJJt5EJu9ih0Q7SWq0enY/zT3fvyFSIReDVRA9L+xpCdNYhvq2hYtOBa
V9lpiJTpJ11dnv7GNuu2MdcR1a5N/tHuzvtj9XeP4gdNWS5EvBL1XrZCRyAzzsih
V6dfFQfX1KJpd25baouJ/034HML8nBKKh0Set4zFi74KOnNAaJDrR13wztj+rAy1
byjgTIiMMvGtjGqvx1EUoYDeDPAJWA76g9aQ3ql0aHzevhDyV0wQQHcZnuP4yrY2
pwm+J+TlTHUY1oUwS/iFXtj3wVC7DKTMdy/CWYv1+9D/GHFdlMldtJ/4far77esY
Jjwwb4jyjAsLr0OLF1HEQ7dSqgvVT0BJICub5EFT+dxYfImlcSUkcdRjBZpLYncS
WY/Kjqy04Ms7tJoN0sMyZz1mb4LmnU7jZUmmTnP2ovC7FBvQTL7LBTTmiee4B+zy
9opggWcf+3ScKn47V6+3+X/hb2RVt4PRO5g5ZkiYkbm4tEyvJkRRo0sYiRa5JxCq
eb3mVl6lFIfSwtInX3SSq0dAbCXFdhSaWrAlta7p6pirvwhRirRG2M+KKe6H98NO
JoqSGu8UqTsZ6whO3kcTj3Z+Qo5EwWfcYYc+kIUHofEaJZsh0BGkKEMmz+a6911J
cE/ueYRvnbfKn10RDorjQExT+eUd2pHK/+To5CKNyOY2Bs/F2mVbiKg7x82RMXnz
/jiz0HrNKxp2qG8jjGTGNcJtWyRU2JHkYfp9xtQWIrx4X5zZP1iZu2EBQy9IxCtx
suHmKKpY4YFybLOFlZUB5PhxrnWAPg0s4veslbBFnYgrT+Yav8dHnBK+okIqUWoK
Dm82TyicgV1QYHgcwlnn0ix8oPQkDxgcGNpoijqGip17r8kTHIKXXrP0NNGoNqX6
owV6LdSLkouB77VrSDjyI540BFDYHBubWNUJGKui4tg490KDSLaxlsdDgTL+SHWn
Gsik6f+oXHuuI9yCmfiAqnWUf1Atk8cfykKXJKEXOwjghzMQCFq9nhG43/4ashzF
nN3Hx1G6p+HJEBVzuKW4SRssvQHCFXRqsX+BLZuu3iht9Mgzr0rxUaCUW+/df9f1
/ZIX7yzmVOOGHdKto19vDns6i51XxcI9tgDBbitSXP5HO2O+F6g5eVSzqkMO93h2
oNdHKjqp8u0vsS4x5Ha/tuU5oNF0taZ85TPYdHYA067i/I3Dl+XtUMQjbxK8eNlQ
ugZ13iSxyO8mpgGXhM3pOv+fNk7asmxGghJgRjGiuxhWZTA1Mrjibxy1O7tRMjKq
ODXlg4rGeqG1rX/yW2CA/78yvKWbGR1nWq+MLwBxktyStmy56JwAvQqD1t5nGBnE
Ri8yjwJBex+488kVldJqMwb7wF+6NHDQkIYyTpEIRcP3+fxa696HtYcmE38vmE6i
DoxvaAtF4ocklu2lP19VhPciDLLnUu7j0sg4asNuRsRD5UnhNkwA7gtanvrnt+63
2SKg7ERU/oYt7Cs970Koonz1ontnwVbIRWESbf6I7X9wCHFw9OVNokDuo4s636Cg
cVl5jEES5puyRaAq0mrfjExCZ423NanULt7sxEGPQCQv/6nWl29Fh/dfUTAfMt9O
YfPJ3HUaM/76Yi6UUfOteTTYNuR8W9W63U5Ta+9Fz9wSSlxJX9ZjCivJ9ZcRnVtB
ugS/llWJSq8fKJpa53SHiQxFjyXEiu2MjtNtkfk9NH+3SGcla27fHPyCwkyh41QH
fhUg/d0oCqSvz1X2GyqTYt+7+rthVqjF7I8XxloNiifgM0PjcNNYHpmVuRNWFoHl
C0Bo3NoKKBtFYZnDuHOnHgZLfky0mD36ZtOLr3PjWl5U2giw6IgPD325CVRpb2lu
g9EpNSA+8r92J8+n6+gJj1axskU7jFKnU5T/DAYhP+YenZGddCFIniLc0YOfDClZ
Qv/DKsS+SOin/PJ719B4h0r83MJtShG6yzJHHIkp/mKbdtI9LAode9WKhpuIckBl
FJwu93QLpHc3aQYVxKmoYkwYgEU+aE+gssTMv5+KcLyl2xdy+4TgRjbsjWF1RjS0
qoiNoHCK2h0WbUh0dP9QHaQ0S5m8aa+r8soGiLh5LgH2JhdxYN7ZIcyB56KGNA8z
6NKMiZ9p0VXFuUfX6RouO4Fq6xxsLKpQqWhiusJvSlDe0Y2xVNipflAwqQxmqJ3X
fyDhy36l+PohvAjkneYPVRcQqDCFh4Gq9gEx1Og5mX0EXRy/RW46onBh9ah907IT
Xr7sE1Q0nWSvb2a02+j3Wxp19hqIES0xUEfPhHqFsq1QYxLmvev3FN/dddAghanu
0AkFoEZo5jnfhjXKB7MQLNhYRmq3CoIJ1Ol83k2wyNR5ZHfef6R0Hh8WlSuJkEh7
bsBtPZl+qUS6CpWkxK0j42ckQRtbAh231T+MTVEYViDuU0gf+yPq+KNswywFGx6A
OeaNVa1xOgXxr7feSU0vgJtENnxbnzx5MbRfMb/rsP+vF5LEmYFJpJzDeqtBhKq5
HFTPoYuIToVx6K20TYWth5jM4TMzNnFeugNN50BonxRkeq6FoCXeH/kF/I4nLo5d
xTSf+lON68nr/miCbJcaXKjBmEADVAbqLbdRUAoLZzGQPBd8E0xwzkIJF7KAhkSc
8u/zedvcrOKeQ7BJWDikTrnKjzwT0maRSbBivNBs+ydrtAuCuDZJl7Kdg0Ujvkbl
Ko2XmGu2v6VyXfUXvHRfH9f/2O0E5kvU6aPuhbGCjmICty4wXRdSkmxrBde/AYIF
1drUw5su6UHISD5CGfYMw2tK9U3XdiQpBDnA2vJSG0f78vIRvZ2CJg61iCJAcDD9
Raa5EJRunxQNyqkOuUGqpUI26ZHwMLAHIx9c5xSB6Y1U7T/mHQHKgUZ8FBGdcAWk
Hv6mbUrESZvqAw60Tfc/0bUYdNZ5/VNxAHiozL/rimAkVOjbuxKhAybwrdphTY0s
sr930Q6k0xYDxUN9vC8yMkpFjhD1ZDWYnxUBDmOBJ32xOhnPYEISDpOUagnIP/nH
wBkljJeIRodbv6Pwe9r8ZXiPKbett03chj4al10lgEiC8ff1by1o65ZArxA00roa
JV09gSnMlhCwa5rxJ1xw5FzSozMOvOjSmiu+7piLyZ+ZTVJQgFoQf7fMxQG/SP46
1RphEcqVGlRGSN5YAITH7cvRAM0CbXxbx9W+MH8g3pergo2L98fqFCZ419Di4C1z
ZZcfCq5hUvU2z3L+qt0ROh+rR+xvj0cZ5ocVLixZOl+It9LyJ0DrscsQwrXoZ8Gj
zIR/SnpPUFpwxdUaUyhoZ5R8xUIktYrPbUbOe0xpJ9NewwvcoqjJg11yLmRUV0wb
SNtKDH9K36IIxn++/cig1DbYeoYptDakh+PcD2Ec6pj+v658jRARm4k0asSgB6Kt
V+Vh4cqkyAEDFXiNkwdatWuzR1y8KonvwadX57GgD9+xn1o1DwD6gU4zpgtVb+Ei
WOD4B9MQxQ1tzAdYmLBx4LCWVV2Bk7ruXQPwaHclDCkXoflfqzn9bRONi3IeFN/K
nUrZd6dEWFCO8eofjr0jy3Nn8rBMaLtF/atFMFcYckxhPY96Nkivozfw5NZrQZZs
nW8LPHO3oKCw/gmwjvTkfA93r8fBKpsyfxfWE7e3fudexLFwB/EDR4wQTeNoMk1h
tJh5GGY00tTvNMVbR0EhHJsSAAhzR7s52Wk0/ggQHJ+6pY4vfn2n/6gK5cJnA2dB
hfmxX+7oKGrg6yCCCbD7/fcxEr6Rp3NaYJJOlwzruGdVxITkNugOGbgzKD8Hu2pu
oqjHJPLciuYIbs3kFoJ6NVjVi/AoPI4T4OOyj4aq78Y8JbNp9IZAoa8+YeF7GJ+1
eJVq3/WbH6qupJ9nvGrF1OYEqEwde6TdHWAnjRIS8ULzd0sFFFHy7H5SWtbjF1e5
lZHlb4R0SR4XT9w4Y0muGO78dwyh9MMdZrUu7V1/s5mCTnczEru4d823uH4n3HzC
cpMxRfSRNFx1SCt2H6VmZg51J+OBy2+wt0itP+hyxsMblUtqZ5+jJZnMFBmWAUqw
XZM00wrq/Y7iZat9mX+V8v1FXgJ7jdmSlPjaSWibUg1HqhPKP6Hch+D7cLGtDKDX
N6b/JO8BbfGpk0DpGnk1DiqtFvI53MUhcREsApUtOqg3ejZ5nwORwQ8091EGv4N5
xWLbzNxtATMwldunQu59Me8aaV+arZgzmVDMTE/sd3zQoym+GD7DO1O4zBEztqXQ
AwGcmQKA5Bn536Giveoc6DLFMfMiS5y//8tyTF34TRPX3v/pBYGmm+blG4FR+y9r
1+1R6DE3ckR5ztpFvMgY9G7fU7PORZadXaA0zr7qxqr2R1NVedvB3bIPFz7igu6F
6aNkLkwVFhpscP2IO7RIlNJwkvUmsAHh5u0o4/Tcr4YVV0vNJx9kOvRcLd3OyEab
KAjwu4pQpjzCgKb5oQskjEaxH+vIHTp6+NvovbSrJX9+nPJkUxfwyA/3fXQ1/vpu
J/DTaa0JT9KQLideeiNEX56vAc96gJgWEBMyDA/WGIc5ODd/bIjPo7T1IWlvKEKd
J5dxwhwEaplXm9kcpy2FUs8oFgJb8BVD6yLE85NNc9Bly0CF8R1pDjKBdX5h6D/k
6ut0/an1IyxrbVxHtkP8C22W+VpBF0hQ4f13yFF8rmCnLDNe28JR8mxnhK63get9
f2gAz6YqmPR9X0Wt2Y8cPMhTsJJeiopHvcaf0bPGaI8t5gX8HAOmLDy+117MmaM6
Z4RZRFLFahBeiQkhh/Ewv70VkEBAjIrbwPejTw+pkUo4REvD+8CBngPg3KDYuAR4
C1kOx7h4fgIGSUK5Hmg5oIDHIRTQZkV+wfLk9siApjiJ14q5CpLmgW6NLCt+1Uw9
zCzZ9NuZyMv7VF0EL8IWxrnjndCfpgMkUVXEdbVrdCVFE28fVDXRxtvZd4qFGDQa
XpBfgDF9mb+8qVC3m0LgnceAHnEhO75NUOvpu5tYqTlncy5uAwABr/UaWYmyp9SJ
7zugS2lMqV2kj1RMQ0PovEusMpWnkgzDRdU+nYstrozmEp4FqknhVViWNPZjq+Vg
hQGxMMJCSIQRGP3u41tjS4yEde/PHkJxnNtO+431ggTnuSAAxKAwnwRAygdVNFRG
aQuW1zQmGWAtTiG/mGMU75TslTGWjP3HHtLQn231OhiRHNMLmUVKETZL7mvUKJ7V
Ir160QLXSXHDDaeO03wVKOqxaSnfo0kzA2oD8AVa3vpZZxrX5jCAhCcWzyiWfl00
P7Qsn1+FF5SMEeR/SRtIavYYeUvJ6icgA9Sn7DfMK1RtuWH8Ia3CIMvIeqElVSDa
N13b1ViBkrpcbHnkAXPls+IDbOLdZquJtoOMDswm06M0v9fwDueqkNrqzJMk3xal
Ng+K1WMWmSZS+bHYHOplzZh+qdRp8Wb5QTQTV4LSXiO2RMNSfqXquEOSwNWCmj6U
KtBBLhxhcaWv10lf1zKipKyy6EZTZV7VGuMx/ILFJaV0Up1YmI1qV0AuP3HGEP1x
XNBhQd9qfpR1av32oNv0m2mQxi/udn7ap1wvQ0X4jQuxZnaj9cCNZ68lmaVG3PIC
IaEmumktxIw5ggp3jgpKmZozQ7qKc0/jRGr/SHJv23UGCj4nbc5xxqiA67W52Yic
i+QvLeefmvPWVidebCWlohnMoQScWjSlSlhTPBrTRDgP0linw0ZbXLYmqVlHhtuA
Du0oaT/2kvJLn+HACg9xB/JihwBiHcADFHVhCFSJUwCL88A9Q7d4EnIzmad//GDj
PqTu3itkvezamN7JL7w9L4pTLybfEG0aZH0HzT6KNhf2j2yihJ3ZGsXNhgr4YVWv
lJ2HHnejC8gEPKJ79HJ+uYuDJBm0gv6fz5SN5CvgP0jdDjpQhjO8QSUjBhr+oMOi
fqkzDVhCbha7EBVrByoDhyhDbikrC5ZjTRSWnM/aYJjuX1nw1BJSra41a4U4kgNu
8E1YpUOHFGmDcIXiIh9TaPE9Adz4r6Qi1kpSZC54pwmHZa7+NqAAe/PXCnfkKJE6
Au1JJensLhGwb0EnSLjn4CwGRnbnHyN7LZQB8625RGAAsAkySsGfAjvONiFKiQpv
P1otDQlWLxfcOvAXXzjzLX0S27VA6YJWMNdFLzZCdF80b5Hgr/WpkK+m/3zfsO2A
bKGhCYaQb2Fi+2GCyZN4AOYt971Z11vq1mpgBnqOjb1QYxpJeCZnpBst6HUTaA0z
+WA0Me/VbcmM2pPh+fREhMboqkDLEZo/kXl9ZCBjmS+IQ2byyy5LBK/mMxX3TDfY
jdnkblsGgzY+Lz9OCTnMyn6WQVwp3yJLv4xyLoBLAN8I9964SiLNDHOAsVO2D+60
3L4NCiVb1Ud3eewrEanlqbmZmdFxl4quRjGxR6UjhcDFsFAPj74mhx9ohOAaI6iI
UJEiO6eMc5VbVwdkkK+ETDGumF8xP9r8pDGrieEakFhJxyVuCAY31NoTRXMNnUnT
D2OqozgDpfhhmSwZEGdLm88YDh46CVL/K93Al9lTW9/27W8iAcTAZtDJGq5/pUfT
PguWPDQTgcG9yLy4tH+tjPWzv7LXzIK7e+gPy+YJLUuoC7sH2CJHOrjB8J0ZywMN
jRIenR/qrNtNuT4mWy/Ldb+q98MFTFoKnaCY/L/qWZeMKsxCiGtH+usuwFnLhcNv
i1bZx7jp3So7qtzFLBV95A/8z4rjp4WBg22QGg8ZGGFWZiq4nK6MZcwlHgGH1MiB
en8k84RGP5Fd6/rSSmNwH5chgoY6M+T4VeFr3i06C1whLbBr/lel+AJQoxpw0PnU
4FlYGopjQe5GkPwMhGLiNHQm5W17PKZuZoTk5+ISuzhfCJX2XPf4d4H8CCL/QbE0
lKXgJmdCWe0Vbfe2+wHankt2tV6tq/cETe+AJ6q04CpMoIWvl88XCXlLucjuy/ig
AcLiNUZTCxPHt7r9JZOZ7HqAh6tE3RlOmK09EFWQ9hW5cneKs0hPNaiIJvppwlv2
xtvHq7PuPSFqwmurCSI4D53pW8/6lXEyjWz/ErBx2eqwrsLSt2qnj0IVBhYst1Jc
6D2Uf+c+JKYpfwtyq4wUr1Ra5XQsxjLt/TwyYkupuf5pIyaQwx4MDTy2t5Btyt+0
/OG0pmvx8Mo7lUSA9wt+hEyMJGm31HXSWVo5kopVSP3XdxVxDcTXWflsFfcCR00Q
mcui3clwa1m0UgyVYqBWf/zeJdOHcwtIbuWasMg0WHd8vyywD13JLkV0wt7SsOCk
xFAt4Xg12YGiuiZMN3GscT4HbqfI1KlpElSv8lcOR4U8ZLgC08iBNkRJTpSgNqcb
gKHG43AoOzW6og4iKOiO8+K/R2LlMUvyW13uVoxbootWaGb0mvO1hNte+8o7ovJ+
7u/Pz4yleP2Fk2jojf17+q/NnncppedHxZ9jIQg7+A/VoklSsPOvT+8T65twrJde
KRNebZ4a8EvPe+E9FcNDUq3OrAyN5Z9CUCpPI9B9EMITf1q3CyQKee39FObqla0H
FGIsXSDeV8LvaYqrx6ea+6+gYk+XNv6dQNBSZacPS47J+ox9Jq44izyqdUm8M0Xq
zQT2kwCWyQYaRaUNFJU5Jt1Yfc/jc8Pi94usziI/Mb1KOhQtvMwsp/ijG5n6emBs
oKRqS41wPfazPZf8JijorZPGFqtXGd6Bcdz+JuviT4W6GpHWA3aBrzXqhSgOISn/
reEeivszq2Pz5DhrNZaGOlYfvx2/n7Hf7bocQrxnIqS3FVPA7BFuwUmWtpVt794M
4u+iJ5/FDIHzVdagly2T9xT7BGb2zw09vWfN4LKw8l+Qkf6xKLwy3xHX1mEEaPyF
shwbPv+11R9yAXk5ptyEDRdVsIyJfzVWSRJkavcIWwv9WuN2U7/k5ZKqLfUT012A
muvxBXSbR9MAKzK8rwA71Wxvm+6+94DIBH6PEocy0tIVDCbcsxNNr8WWYF7DeyMC
/R0m4BxVRg6UAt6xaOHQeUjge0BkN7ybwmkMENkj/gYqb+HJlCQAUda6iL+4PIVy
ES4kg5eXoK1Tx+3xe67DPgXqBJwPRgs3LK8+kNrF5r6xWGbGS0GQOMutZjjD30uz
H4/KGaXt1n5wUiC/PkmdgrOosVrsBw9uidGDQgIIra23JVhjMQUfSMpTRe0AHcvV
xk/u6n0KwvzekxeDSQBNRtuFVb1bX8TUsTYoQL5/hDr8EqvL4HcEaw2XUC6XTUd2
ke/xtLkQ6FzqchXMs5ldUDGO8a/pZs+jUY9pPtJOyYgnO1yxZwbZtqYjrpPRBCXY
9PCH6EYKNaxC40tT5XJ5Dr0hAqLFniica2LfGOutsZdzKrtn0TKi/I8WdVjd9JZi
PU71xcPkGBA+rLnyi6k7SbSyTnGpQt8a7nvEjmpvCMV1vrLmC1cClSHGYSJELKBn
y7xgi+BkiLiy/o+mTpftqzhpoHKQXIo8FdpAKJMbtLgiJgH2st0Pj+FHxmjCToaS
KtDUIdOs65PTIl662ekyhTy8+ATuImS2SACAwFffKQZ3Gju7dNpy/qqoWIP/tLxv
Gyde2EYHeT+v6VavWQDsSeuDbByVA5oyfFxguDQirIBVogpyV9m6D4uVE9cjmEt2
H6Hh57GdAWIGWVnCFwQaDoWisKhwzaHMN0ehqe0vzWFtHtjnpKNoDfDkBrFsBtR3
Z2I1IYVK0x1QIJPu70xXcUSXu3Izfb3LhCNohPl+M/GlRv5+VszbunQdFAss6zuv
FEKPXKttG8Ew+H0gVAUg4UsFLNdp5ExaEIb18P+y8LlyvjLILELwO5B6gEP0FREa
OQEZbznVVvMK4G3V1xhSiZEV/y77MoccNlavOS/bs1/v9Q2drYGKsSXXFvq3BxQA
s15NYiCZDK+BU2Ub5C2JEYJe/5yHXzfs3HVdmhztz76yBZuB5hfaiyfo9al9Kquz
0O4XM7A0UZhjFjvy33ZjiLiw9MdtIZbqMxNEWWxKdmT25QpvwSYljVc+R2nn2bF4
Brt5fCEM/dWzyVvvalh/tVOH364b26lz1Om5KCrULlSa9NtQFz/jjv4Z5pqrBXzj
d+OzU+cYS8gG3BHwkLIsdEJ3dp+fnyu1wys/GXgnPIojqEEQAbrZk7FKJdMhC8S6
EOev03NzpiKWxrxsqgVK6sM5wwQdrwptCWeCpAuo2QCCse7ZHoHxXhX9PujhNEWP
JVdGOP+zdbV2ZOg0vJshtopvge8tk5FLfLH21GeMlPIzlMNtQGIKeRC0sk+S6E/H
WytZUwujrcckyGOMm4PIWES8+MwQmqKL/yd+ND0H5Vd1q9Ah3EE3+0r9u2z+0y5U
y0b142xlB7EBzXy8UVJAtdij2jXrGk3EqtAn4bZ7KrwJ36bCCGu+K9PMptB0M01y
mu1gT8kCRXdzxjQrSVgfhlu88ndTQOT+dDQXJvcnIvpi37LDlnwEtuCIraFYwYqf
D9V6G01xJH5IL22MW9+YuiMeemEIBk8tdyNNdtpkYn/q/3t182ptvixUyFD1+0XP
4SSvOcvMyBNHO3qIQIXTorbN3hxggVYWAD54XpbYvkoARXqf+OjTkpYcXEWrGyp4
eSdS/2vZ7Z+n7RhR3k/0jyE3/9Q3X07m6gyVlA5jKvEpYYMTF3RSpA6ASx/UWg8J
5FbshpYbDjY8g51/bDr9miIxuL2fI+d1ivnkMwPqCB6vnQ+0choKyhA5DLSp0Dqh
jEQrR2WsWf3ENuMn7sWnjD+nv8+jBLuGCWh83Ubjmrf171wRzev3S34uXu+dm8RU
Ay8I4N4pry3DWb7m5vzmb6/iq5zTdJM2Oy4LuMGAtW9Yo1N2LiGVA1l/ujiSRD+a
SUTGAiV4gBP6kv3zcae/9qRQbjpUuu1ce5EmhHsuiX2Eh0cqzEWI0wJ9CnUcBrwX
6atZGcWPgeyqgk/fK8Y2H8EmHElh2vPGFHEhTgREZIXDmxkGFqwFNGayEeWURTeC
pmVbPKFe1y+NS+a1bmf1OpJNJ0RW6E14cyNhVHrtPCdUe/yZNJ5g0ttsXpCh3qzj
ncH473DeDsb9ajG4c7Qf+7fQh7SiZR48YCSR1MqgPCtwTpaKDDNb57N6v1drH05H
K44mxyim4ixqWDiVCND9YkcTW6qCsoUmcrmKPqenJlijLBTyiJnP396/b++bZrfN
sltdeXCV2aTrIPBg/c6Bo7xzTRExs9YlKzx47XOZMTj4QcINcOWgy/dyMd/je9z1
upBBo34c/O1mwmntp65NTCwGBbJQZUHLAnO5w/RdqZ7H4MEgOYBYXbgYSP/bPFLG
PWnocvp3Z6dFTTFX5nXDZFt+WdlJw8dUNpqakKxsixLY19L4RK/4vANdnqQxxi9w
PC0TN1GJZ8QU1gX1/GWbXYd/rGIx9wC3OGL6BJuiaKMom4ciZF45RlmXTxBFa41p
f0115OOB8J/QqvT+DbNnVIPs4Fc+lB/MEYlKCCqHgpTJVDG4DuNAvrm1YxR9+XMD
AEy8Fh8hMmz8QtoF5P5Hp9AgvsRArcJZNyDGcbcN+yO1HXWs9ffum1GUMvROZuot
omJ8NsrJ3utL/Ma3YvgaD1gqaf/qvBz3CNDy8lceGXkI8huRKfd3PBJt7nUpmZ2R
3tP1yXgP+1OfvSUwEqcu5pVZx7nPKBs00KzjqSF0wx2NhUF8JaHi8vJAhmANZsgS
B90AybV8XBwM0gWAjWV50Br4S2kvUJWdFlONFp9/s3ybTvvPpCrMXKXMpIIoeezH
DRMVmJXzWeQpQOb1Lpb/FLw7P2jGs8WJX5FU1MA5hbzI3+hnq4Jf3V1CFKiq23cp
uKUYS4mAtkp7Z+bzHdOcoT+Dv/hlmEqslVS7wkTbWK4dt1fH2VP5JW5OHibJ7J/9
dLnYRu075f0s1F69LtjguEnlFAIJyc3DyJbjxkafTjqV5ZqZtOYcguEKdVzmR3HX
cLU2H2IsU8G01AaB5qQXLNT54ZKgULbKf4XdglL/5xU4KVwuuXplm6+Al/Lxh7Aj
9j6XjWH+37UF/QC2wMzQGhvsno7nZ+negQc3Nusr+RG1ormqcNW8KvsPPeqaWTTh
xUQOlw85J2YRBs41ENeol1xMvZn33O8P3wPAXiNhLZ4hH7nQCtqrdGkdJa5lmVIj
F2fP+c+P0XHKgqloOrL0I62rjMUh0QceaHaEPX/y0Ur94TY6qFvcckeE71omKNwc
A6ib5hrtGwJbfO90KRVsdOFPzp4V2jZLu4/dqWj7kKn0jiO3EfCv53Pt0ukF5Z9O
/pdgU2+fCC5ywSLpMR+u6OGDMZ+KYbZ5QKbuAusYrt0qDAGEA6c4ctxfGY21Vext
sBhGDy6L628i0vFw9LhrHBm4KjNeMFui+idrSvp9sm1lr0Cn6oPTZulLGTYRsejG
ygueRRiWYm4GVxWzwMxEVxtUXVd/XpT36j7eaMQkReGfsYaSbwtGNd3yiKCBzMFI
VEHyS4udCtuN/WTYBx8pfrmWCqh6S2eBhUlT9eNGvnyXH5ef8lkDK+ge47wtxPF2
TYvnv75T99Qf54j90mHm4JwtbPd3nq2ZJxpjksIZxuwXldUGsbeDFluNjOdFMO/b
FEUEg56s6uI8rGxK2Kpua0T+KJJLVtvntNyj1PpYVh1Ryp5DhVXh3OPY375yVrZm
7mQ4pB/DFWBNf+1orMTXcBQCRe2r6pSnqyCfhbnLaurXsKmDiBsGo5rvoCffq+C8
DyRK6C0Gpv0btSiBTe4Nm/RvyhutcP2k1Pw41SsOXn9W6eBSpe8RtOYmwDvzBnPq
Ha5qti8IuNyDzMG+cdmZTMHaC7BBHZyECLuMASm5nL5BMM7rJUPSl1W5OFsDSqem
7BxX1eSoRsVZnZPmTkMXGnuVOkBZBkjDmaRadykCzTGpRXeLu1fOQ+Cka9HZVROL
b7QUwlrrXhvRlq43c+frTlAC//lJO2s34hjSrjhpGowHgHtyrsyIU1H2eBA9oRPF
BuYV6bGk67alguH4EgJuPB7f08NiTi6kADnt/dQFb7ctMrr3FLE0bBJbrXhUGF5S
Vq5UuhKaRKHerJPofb4D5EpWLKQrvHKfif/7eUtPS2kII+fSR8H+KOrJaf3HbSqq
CtM+idBbFnWrbT9QJKW3uWDNKQUwHh8W8NiTm/z2aIy/K9+PXUi0x0qFFDGDjLNU
BNgpaHH83YjWKctCxxkEDJTAQNu7lZksMuppjyq1e4krV4XWUGI7YvIPPmV25B9p
k4GfxxbBOExZbLLXGRvlBI+QJetiS8G7Zz1iGbvN1sOYFq5yHKvU7tNUWDpuTTH1
UUiqZffG3+WqSV+0Vf/qGwu6cFyju4KuCYsVVt9+qTzZ7Hc1cymhD4bd76v5VtWe
HvW4uaKIyFV9nghyil4yNXTd75QmYVTw6Sl43QLHnAOqeb1vHS+kCqHiM70mS5+r
hmPX5NKaAD9xw8hRz3K95e+V8yqWRvEEju17kmPzLzPCdOERhWIaZcEBH3meEp3p
xjE2m2mJsMuKx1l5DWEw/na2X9x0DgoIxgWuhFC124ZyxUFrYbyINn8HpUbqSxzs
puNLIx6uXenDcSwS/vPOUmPuy7f4UorAuVLSFPm3K4uWx0/vUqtWSpxPeL3BTN1L
hkIOHKYlZv/CuOvT77jKAcMkbasCe0u9RMcZ9Cpy9oYnrvxJpftgLvkgadvF+fsj
Ly/CRyK6Kxi3xhVkSDsehD/xwdVLE+FncRLuRsYAF4j/aWgBSbnNbDJMZ4NRN0Ds
V7+iC3Arxq+ylkfjyHJHOF0u81LV82h0ABolIDJEb1f4ECQTcnS1eOrYDiAvaGEo
Zy9rPLbYoxkr6LRzg8oIBC1KMlduXi0SHqwt/YjON5l87/WS5W6bSgc3neB4FWEQ
Asqtr+iLjuSdNNwBQIILiw6PeAlMA6TDYtcXFUjLF9ZPTQJntUTABHMXYwNdEaqa
wpp9fE4+n4MasZTayXvTJoMHmJ8aVQbAgVBVgeC8jtzkeSnU9nr7HPHxJbCc+X+u
B/M1t/sCvOz3WEwNViURnORbNH4Rt3cxgioAEDIZUGnjDUARPhoVsPhjR5Uq8RiR
gNk7PGitUql4Ckk3FSIhhlBZ3FWWJhLLnwA7avlshjxI2uJs97omL7Tt8KKJUcoN
PiZxZRHp+pwb6G1wrcOX6eny7R7mAyhYxszDIlVxfbAMD+Do8K4QxH7yBAJkoEvh
W8Oto03MaI9Gak6jbvcTaidgAs1tCNDHVZ7MRTxxQoPpDrF46EUueVjekKI9lE2V
0i43VLi/MI7b3fPlgzaPhriDGxL0q36z8sJNkUAFQLz1UWZPQLr8x4zuHVQpvIsX
H0pAI5azFDS4XYdvxn7e2TyVhHtf7y1NEiQo202/jj8eyaJyEgX7sbEGl6DHsfYV
IFtFI7NGUZs9NoVZEj3MM0OnE3dFL3ckGJFNI67gqfy/lSvwTzA+1aHR6xtERZWV
rZjAldsHK8O9n8DxOoJ+8hLVKXS2adHk0MY6XOirj0FNaf52NOuWYWAF2l236S32
dqmtAgsd4GmmVwAokuCYn+7v346xH1/N6FVWQTWZD5qLtjm5nHwxR7+Flt1FVxsZ
4DTBxyODw/4q9emc5ZOqE7asvitAK6sku6ui5UrRlr0ZbtriD+YjYw1aoiQd5x6b
T02Mv7xrzCGNCtR+bLsfoaEVt8POv4uzQJzbqY44IoBgnTbvbZF33hjhMR1zd09d
1/KC6TQaAo6KTmYePD66N1Pa9Hkjqoqr9zmzgQO8IT5iQnOaQnEFU7lc8P7xQdSz
5hFvb+Pkq3COPR0EewDZBoMZLPCyzjJ+pac1c2IapEnuRCZH8AEbf0a62DeCPDYw
JrkoCgBEPZ/ALfvEanCKAM/UOEwBcTrcAm+/h+xv2DhP4oeOL7rshqW5adpiWZyP
liW0Oj9PEUAsvRI1iqaXOCefLiE3aSqWvCq4Tl+1NuUiO11iD+vlX/V17cYoVf+Y
r1eEVrq+9cuhDfwHy4O6R5GDjsmklS24ZjlwBXS58i+dAFHqGzsYWrfOaA0YFY1A
KYP34z8NqfsgMEjPCeXoyZPVaoNcHLNxCEJyeOHeLtOftKsDtMInrWULQq/bP3L5
cshA1ifGTIAnsP73rjfFuGD4KVm32F3UtJHFDfUzESJDPQUGc6Y3e0a1P+hZHc6q
403L3F9XfHDUFAczBAYyxjshX8NQHal+Pi+wySVukMVHN7m0rAc6eV//nG7quz75
b0yOEmIbLLQEWAuT0CawHX0EN7wuzmwLsdYiBKJBgb6qxkHWnkFDmlEZMWTTeVFb
XEJLjEs9ETcYWSQwpZvtMS5njEI4CAS5YHacwCe3shmhltWaaGLX5IvR1A8Q4LBy
YiM9jat9houjDxJYFBEF9rgaKbLXo5OQvKjV8Lwz+kPPeFmWasBb5xCOG84dwiJK
NCR/Rk5F2wYwFkzx/suHec3ZLCCLpCyHzJuvAqsnZO6e071iXjlZX2j2Hi++jW89
qkAJ/HGJ5P4obbuaHLXPsXM3bresC5tXC2ETsCz2G1L8DJBToVcut8LKRVuKevKi
uzyMPftMg9RvZVIDRhsb67kdRAHzIyUkUrLci//8xGxeAsqq1PHBN+YMSl83I2vo
DI8NkATODuCVGGuoXjuqSeUHsuEN52Jf19bEi7YYojSfouSXPL9atLlmRTTyMUI3
r0KAVetpbjUzp692LNP3Qn5/K4f1ebRSWQODHD/7GVtM4pX+xt1wranKgxIa4apP
QSHMJSk4NWKI51Br2RjdEeeL1fIPvOSfqfO+3t7wBKaUKv3hatEmZ5b3tAVfDr00
+z0a0AnBo4MSmQwjXJXrXxEXSS4X3d5avKm5+9iHfLEU17yRH8dPQCsG7taxh1mk
SVX1kwOV/IxzE6gYeg5KjS5w2STnggXp3x9/15W4NEnM3BWnQVVExbvt0MdJ222F
b+NLYyx/sF2mK5fzG76d7ijEpzy5qWU24PlgCWvWIqBYYHBu5LEq2mMim1g4yq0L
3S6756HIM9qqgeIQeh5oIBc1graVu7lkCqQhd/CYaIFd2BMVwEdv27OTJFMo1ugZ
JbShju85ixFaV5JZgH3f+OXss79wdTfGKBNvItSzTFyQhrbUQFm4xaJ0KLcMFlBC
1cF8wqm4K+3eNeAJRkP4wZC4wod4tge/8As84/8fVCLKgMXK/wc/sjQPvdegnth1
/l9CmGffulQpBNkWMvEiZ+IP4CcJS6UC+gq/Dt200w8ySMJQ5lppbycSKL3Gb/m0
4S+o+MTWznaLgJnkiMEHdvoiNyRftP5nXf4pO0Pur9UryzMlPM0kjLbPuB6MRjf6
b3GkU62wg1/YKWUTtanIoPHxP4U3Kcn7ZQUkp0uHZVgDBWRmoOslEQQpPkeqo/9X
9CL0opbCleT9DgnAaplm7ZKTaOOlglM0jd1Y3CTfnaI7KlvkftgZvInUhGSbPkMh
2C+gW0ZD0Cs5YeTAeqOA4JmxnuUroqhzohunhEEZLags1UJRZIOozM3cl75lq+Hz
pkO0gMtnfOCqNfhUwKq2ovarIryS8NGNQ9MCg0cQtPG46f+gsbQVBFUQSd83ZlBa
YUvJh9Q+yRY3ILvVCJ/lR9YBQFTnspramOW6j9gmtHwSo4dNZhCngmYv/pumFEtt
XPV4w6YHSLQsaap5+DqnQYhsuzORo8NFgSoX2RrMzwwwzh3p4gYYX9LHaHnyzIhR
h4Nlgf52dTH99PXfJ+sCPK+S7aUKgx7+e62RYfC3iNLJbVeE9Jntpt62TyIc3Sod
3LaFZl+/wXdlogEzzQ/5/jWdZXsFMcLk8coIGJkRp0mjs2iAhRhBKFIWJIogQ+D4
RLx1N3xIETbIuUEH1baNu+sOI+tRAGRcBpY2iqvBwnln0qIDZV7a0WGu9gMupUom
JXb18JCCUl6snw3Ge4M1N6M20F27SnCD0Ekc1/0W9b/Bez1ovhZBsX01aaMjHNcW
C1Ngk+T0e0pQFqlpG1IAZtxytuaxNKFP+Ut/MEbQaQGF99qzualBmsFDzNLDzc54
nq6xTWShslVo+z1YxC3NjrajPc/TmXbVne/iJvGlEevV7KP232ueeYunN0RpRrCJ
bQ9+crAD5uuyoBUZHD/PUmuE5Lu3rdwQ0q3U78i3s9XL8XsIe1IFXukNbeIdCZxn
E+7h9rJ+IqIGv+vmlSvgy94puSdjmeerCv/zkiyuus7dCt8QiL+n/a6ys0MbX2rT
EQEW4f1oU0ipXM8h+DOblgP6GYF1HaMj4qVP20D+4OPy4GjXDYCkrxv4KAyPqMtm
XSKoW2jT0N4XVALh8Uh8/ALZRWqDnZOBhjminmCNEdQn8mMSqdrTDuH165fyXCL1
P90tmBeMm2npxiZmY1JGXOP8+GRcSpV10R4ubRkDarU5ANSgoOkEd0zGQrM4nEbW
w93uashif+duFr9bI6JlX7N+Uy06rEqGg82i40bkvCZ+9Kzi7G2fJDj7Lv22v6VK
7RNZ505c5I8HNzmdCMEzCwtTum1EsYSZs9zvO6iyFr84AP2IVicMq/7nncFqjeq0
pIQamSYvlXgQY2ggPOVTd+RaNaS/0fH760xTy7hfeye/CteDuqWJFDs1B+JVRl1m
MeaIahCmEeDy+nalDxpwCbOnXu2B5J5wfSAiuOY3wfyuSmVFEC41c6ZNHUpGBqO5
sntQz/WpcBG4oZxtYnCGh62hJDdjd+jN11ZT5pse9+8KSxMduKHs2N8GiKhifU8P
ud3FdAeB3r+wGfrH6cusgvTJ2duqiOqGAzmBhk/wBrM/GpETOTdE6NwJ3LwhJxw1
OSeWtvqbCA1tRzqLfeW7cVAFHqyFHmFbw2+BJC+Ta7IoLO5YRf9mj2Efvz8fK6hk
PBTOcjDfj/pz8zdJmy9JyPo9pRPAOAxCYqwuYzbxasyxcCWk/l1Hazabld7b0fB7
DBamZEbzz85z1UTqL+gy59FEshW7z3ERDg3livyuRaCh1z51Ds+f+OCzi1gH6en3
GdL/6A1FUQt+4uffiMWOWvjCv/TQ7omKPQY4cwhv3YGoDL4x7MSLmXoLNtZZYN01
f7QhV/U+sd1s88ca3v7shyzRO5hWOsO72qRDLPMF+MYxQ8Tb/ZqERrpou6ELy9iP
TbFhqHYSiI0vIARy6mCU4CIIlDy6ooa3rBEJpKBJYOjSC0toi3QstmQoT1xXUFnA
XxnE2avgDF5o0AIP0p+hvtF2ZtOmO9NYx8DfGCNLC4eTj1H/uS0iKkMpMzA/wS66
SHZ07WEdXlFYd+KLf4ONpuV8x47YYSAs+hrV+dqvAZZp6Gt1N1YS4lFsxdw7OJ9r
2vV1dlPcq4hjiNVbFKBzA6zc8b3ZGZH4nuBCCee78bK6IZx+WAz7piUzp9MRvh1t
qhgw0Xvqbq1BBP+xbp//yTBQefHmTCir0zbBsOdcf6hKTEVJ09u8Swvrc3AuHir0
ZGCfdTtRc5bkpH45P7cVJkHej3lCoYlfwlpf8mSdGKL3T9jWWkq7Ca+/5y3n8cTg
CT4OoFHN65iEQGsVQOqaK05TRkIayTiUJlE9cl9PVOmclOXqwUko2m+WVE/PCp5Q
chiVTDvOKyioVFbViDf8Rr7xhSey/whRM9Hiyr+hjDC8K5ANC7enO19aiFTcoDTd
0W7P34YXAIWvBeki3CzsyZzlqOZ1sSgSM3gZFn42PSo44RcPI6x5AP2m+kzeb7I6
+VXJDWJzKhtKddQ5cm4M2CXdCFVVtVjk0xuLiK3N2R3TGq3iTX53D7/esUCEXKcx
9BHoBy39jNe4NPBQyt0g0zX+FdUA1TEAHzNcJyzqNfN+FBSJiDrtiAGy4LkfI8+S
5AmdgsslA6FNScMupVGNu8rFC2urst8J0Ckyn4ZnnPkDo1CbPVFMbXd123WcPnuY
qMUOXGBrZapIcd58zyR25i9rdeMQLExPnlEzYgnijwQVqvxXDG0YfPNMQCzCuCPu
43IUk5s4qwn0PFD7IHzxO5alugnOhNA76tE49sXLxqgfy1Zq4Ojy5CCQh/Jif+xB
kKL0e/pVyyhceygV0dbDKYp15+RIHv0M4+SJTZkCmX1AyjaGTLZ4V8Yb5M3ANKI0
7TvSDXkXLrGqFiY7odqxqajesVqbVNOROlc+v2zTKLIgEqiFgI/yeY5tCO6DIAJ+
hIBzaZPyjXt5T54dg2GzUd+kbF+V1C+6NfmTjsIWJP/N6t+BsFQfvTeMMiumKxSP
b2eI3MsA29zj3p5i30HecRKhVPUmvijschVlngc4ldVdReJlacm1LRP/F8ZSAXbT
8isBOxMqfNRn2OHZ3bgxTgFfO3Wmlx1c32P625A1y8NsbV0/EL5H6bfBsXJHAN51
tkE+xLb6sEZtdMydgGhCCI7hdNshIzEJy8vs5/QA4JRou4jxj8t1epWhDGT9u3b/
CcoUTQGdbmdKpgO6oqs6Ggf2GLe0HGoxSVfChr+F5e5CgodyrLbDCq6HCyltpPP/
qhZVjgcM72ETc4XZK4USD6Ltlcr7+3U9uiYqRuURzoHv2uv0q8PzKHALgvQAQ2Ma
xPmSRNtiZ0FSBo2Ut5fsZwJGT/DNAvuoVNPnsBVc1i1UnY61wi13SNw9sluUy7IB
X4mOpu2xTRDvLF13bu0kMFxQ9oT3ue3+nzxtmL+/kSlw+OymtkG9Eeb6JSQ2+Zdk
jaFFfuH0kHHXYwNs2yr34cjifkvHJBikK6hF9hJ/MCb3b++PQt9+qZQt4cUPjcWR
AMvsk/UlVHSeV7E5oYEIjMlZpPxWYDO39CPoAMMP0UzIRrXKiZCTKgkcE7SkyYOj
AbsaXAFCdyNX0IB+SVtBNtKM1D/UvxFHyKapPizj1rcKDvoT6v/PI6Ec9keA+tlX
iZ9OR0Ts7sJnGcSgbTKkSm8mpyUb5jM2+S//2zuzflHmalTGA8b3RBHEX8/UQmNT
qvgkdm7DFnDC7rwXCFPSl3n4GS5jYzz1tIm0BX4FdFL0TBi9MalsfZdP7AsvEa6R
0FE/pZZ8Y/yOzkJV9I+aTkY4/eXLiHhghG/Cfrk6fh5VsyVp+6kvTrwmbcuUb8Yd
OhgWpwFaVDEUhH12sToST37Fr6enPixFVxugTCh9nJavNyAEA/qfBYm0XXszb6YR
KGaYzuQJOgmCbOZzkKbNUwZrI3FyXPmGhy4FTX/743Lw/F5rceDWXnJnJurSKpOP
zSyMc/kuh6l+AilswdzKO/pniRYzx6pfEoufvUTRb4fQ7nzhqnJD7GqJEnQ5YR4q
7PiEF5oWlXUlnrOrdPwSunStfhKf1lnk/hDsyrkqQLXYSNfQ9jw1lfyrZsXqQugp
DKpHOAcQ1XigAraEIEm5hMQMK7Phpp/mva/iYJmH7lUUbmZvAcGWRXMVcnLgeICO
jBL1x7hS7WvJP9QZGbQVH6AMHjdH2ryzwvVzuncBG7mt8pQwgYIe8PFVfZ7dvvED
5RsIdayr28+3/6Pjxdwi7wDnZkY455+7u3kXZzcWjkQP/4zchhmUtZxLP+on/2AI
1x8hooNOo2iLdj4RmQUYwqyetWDjJgIe6nO6loTlxGjVw+LNM0EPk43LUj9s+eBI
JUQwprUPXozzUuwByV7yQG53NmmkKjraCLhA3Y/m05ADq7eZA9AFqHh8D6l3CwQO
Ms4vEcr1eYC3N3PautErJTDHi+lSFph0Bc2TEG55Zl4K6rTWw2xWHUkaZPCKP8yE
2Uh3fcWpXNIY1qtRoe2wRu2U7OmH+9FnpQ8dbZ4DgKSyhQSDISVxApXvJzkyGMPl
aDXC4pu30WP5Td3dt0IOAGFt4NUcj2rjxbQujWVJegBWc+3z1gl8iDA0/TZPYzRu
fjoi+n3WUFKQPBhNGRN+Z1hJNdRfqeWB7/khOYExi5KXmv/3n6mTGS9njbmAV531
V98vQnjGyZEeskPCRKcUNF+W4yih053tiGzH02mRSNSE2brAGMt80OPjNVpgrc/Q
ogtgOFPYWRd8t70nIc2Is68u1eDC+vZlNJL8M72qnESF1PezIHE8JIXAccTZT+n2
FEK4nZKx6faOUofISLaLjEkRGCpugV4TxGTMQguKtYWSJTS6ycuTSiWg1KIQazHw
Krk6DZThpl/1zpQ5saJ36xYsA5pUId+6urz+hBYjmSgFVK2yav6QOCRu3OCj2gGk
aOTSgEE4lfT20sNSSdReJT02mnn61lxpFOcJX6xGtDneamPWBo7/GEjXJEIQ2Fmx
+fkEJ3NuHXV4vcH2ojIdkjVFHRo9xItkK8/I8CRhzDrPCMWD+mil+k81DejgmE2b
tsK6VbQwJ7Fl/Hd86kevMbIliyhWyFVxEN+MKi6y97Sc4ql09wtJFe+hMcGPpOit
OzcUvrDnXPxBwSOFhP3cH9PUYMwt1QjZEW1QpR/X9btXfANTfSEAAgJMoaUEUsSn
5dRndQ1n794+RDWdjpOOmQ6O7bW6RXKc8bGA9Uto4fcMf9RtzD2huN+OuozZD/B/
zmydSPxMhh5X3gSi+udtjMPDKBQpjIAG6LgQh7bGuCiO1xJCyM3URCrHyncDw/YL
qVTYri6tCw5ye8avNUk23KWPUfTnDAkIKyylCP0JrSnoe1LDBwRRgPUyBSUCe2/A
Dll8++S+zsbUiIvI3uv8VTEmBoPgrk7dNnuTFFNxq5fVPXYN77WfxYBgf2ONGo/6
B1OTtrUMuQjWpjq17XJd62p7+tbuaCAIeH9rpAgsLV+E4iWtkcVLwS8jOvRlOCJS
l6HzK/8w/O3EiExaXwV58sLigPUTLiK7L5TB7utCloqVJYZLsmWx9y7ukj9595kv
rK3+y0UgfgycxlKizTYKfsTeI99k0jjuqtQMu0lMVx9h1aCTLFsIRBvmEP7o/9L9
w0tW46LUwS6E/ibf7pjUV4dmFpTibrPMqpt9SGfSZ4l75AxtRB4F1tE+O+8ZU+Ei
3uV04mLbRW/wFjivw7CJn0Is4KSHAzmipGsMcD8fdEtv0K+v/Ln4D/slaI8gTa/w
zprlrSvr1EjlqsQRQiM3bEumC4bjQT7uehqeB4ZbGK0LHWQpj2sfl0mnVL5bP9/B
QHJTaLGYGG+L/xhHCxiS914tXfpDFVUc24fQL0O4Rowo2XLL27EEI3ArX3Gpjbkc
tmGkZedgMAn4M0xo9gPzgWjWrVTJY15N1MSauUuhjX+T+rZCbK0TzVgWhH85/JwZ
7MVhiD4IJH7mJFtprIQ1jokVY4bHG++947oOtgwRiQCzbv5AzDGGLv4UHwNUv6i8
q2qAe1Bze3hw0d2O4b0p0m/M9pkQXyBT0uRJozvqEOGfGGNcDbmrzMFgBu4WMGtd
sK/TcnU/EFaq1I1RhtcthFUYC5/SJIihSJGPrrvhVwf7aBJJgWVq5bub4JxQYxRS
nc88dCKnJd5lldbVS4rep1nZAPzpUTAwDz43YDGsaW9i37pBwkkw0gJwywbSkrF8
irpM/oVJ/tt7YTJ/XVjAKQqan6YjV5mEA0icDWygKw2c8lrMdrOsAg14ZBx2rc4V
ky4WxjO7r/OQznSd1yTRf6CEgD8/97JSQ497FU6G4NOgaT88EKliZF1FNBdn3aKy
wpDybE/UxlQPpe6x/5LpgjN8UOemdigXFqjCWpqMZDrZZeJKq+IUer1rQFbn87Di
OAWbYL9TW/LrC2XWkdxsp89cXewwLZeJyXUmaQ+moOOoj95QMBtB7zWmKZMtmQSX
oZwxfjNk4K3lgceWwi+eCa2Ha5gjdH3DZmKvJK1KusrX/8oZ/BrjsFSkKWNjAPDe
MnKiOyGhjkH84hUiKwu9UM9I25kVZY6GEJ7VocVXADJ1G9vK9XZjRiYJWkpNulc9
ckxiqHuPLPKzn1RUL1bI6jaVbltauOjehq5SqMVnSwlvu/70/B4p/Zfa7RsZ32nV
FBF7vOWn/o0md5a1n5krSl1+oHdiVzw4sKosTDfZLm9laB0wOp5japUreCsIcxB0
/ImD3MV+IIdR/Piw24lBBec8OM5BLlpfxCc1H/fUrgDY26RJU+Hv7CpcemyVHyTc
y8COiJyM7n1aQz02elCnyz+4RsDMdKv9exofqv4Ru5t9n7vfc0OkoYbTZq3H1GMu
mght1lh3f3jbE2fna7yXU3hxwmFwomMV/DvxcC2UC1LLEyq19n0e4Y4DmClMs5cD
O55Czf4n0rEUd8S7RQxu9XcB6HH0RRqCOwZnr3zQ0TdYE7AAKTo87gFnEDD8m1oG
ma8HpebEmlCFPmK2Q73ODKbxT1nDAu0FlPoAcTjY6+NpyBM9gtsuMhwRlpWbntv8
4aWUM49vDrxQf02p7c7FzHdoiRhq9qoJjmYznDFvJ5VWg3+0R9V2/akua0p2s1K1
LUQ2PwyOCUwAiU/9zJvAJU/sEZO4YCjKfL19zxpX0ROyw7jmfwZR8MSIw2fBlmRN
1L/8X7YfdZ7JSVkCDRqg+EPtcaHOxXRAdWirTeb2eYl+9L+F5PC1ZK9SFobRg9CZ
CCcjLQUAs+HGSwNpntCSUgvYEDKJKNtCiHfbjJMkTXEWCFdzbnylviGXPS+lSDg5
ahtYsNiyCQ+Qf1/CqnzZo31eEh7g4VySAcmoYuaEVXnoDsdE6rn31/W5vdf7Opst
/gbOMUp0CcIHEptvABwMtymGEpFiNqj7bpNG7dSMFHzDseYHJVyimFNHiQXRcIy2
zsTncEODzUzO0NJi/eXSt2fW2AhulUNadCgdwcgIrsGj2MippY7kH8TQ5VC7eA+B
GxelXwQaBC2fnNb8irtCLmkDqPM1ZRS+lFOIAYB7qVMwNYNb+ScJD43D1E1N71Iy
TmTzHPN1h7pcZbx+uEEbxhjt2b1k0ZXnTvt1gScV9egDnVo+ApDwjSg5iexLXxcL
tUOctuXb379qnNvBLNqEb4NlDH10IX6uFZeDPTWqUZx3d5lsIggxAnLQqOl/9ToB
AIUDE0CA0waR2h9RTon0oNs2ingdkueLhQEoKKMVvS0VHrdj367W1HnovqmeAE8n
gjmo8DA+3CJ1PiDvenHBtEsamb4hU8ItlJ4Vn01vuRJ/cKw6qx9tGGimJFvxbSv0
M/RUWPvIZeZykUjO+f4WGY335nw2xa3bMlIMu0jA2ZP/5e/Fuy8hVS3BNEDPcuaE
JKpVluL2XLHEc9BQ7tGX5frgiCIYUnugo9IT5ncSqJMMcgF54eueIHeQFI9HQQDf
KW+oJYSu8OdXrAUNqmmtyec42g0E94HiynxQq3/Ko/pteMVc1T8wTXZi/7dTHEyY
n1KDIJysnszJdzfTUNg4ASJyYbESOFmqoBtGC2g66Bv2qn+jXEUVXTmj5vODJxoi
VHG4/HyAxm+2plA+Ib0c5c7oqXKceb1iYrZ3uw61D4Xpjgb9Q6UYLo2ZoI3vA35P
ayDYm/a0Pbe6yo010M9g3ku+RZxgp9EkShqnEO/BDtDTFzSY5L+EJmSTsraP7nfM
ptLe8Jo+vWCvgkmDMcacwW/v70ysoyrbzGOWAl2Xwpc0lEs2MJpd6CCTXckq7kXh
4gdbIdf3sV/P1GJ7hw6SjWGMi+oOpBYGl0vbdawDNAPzn/wXnJOj920OO9h2r/FK
R5TfGnTBfArhoPSx+UmDLj5/Ud2fjSWIkN/WJTUx9IRhyEfhkG1JEQYYTXXLNrg5
n5ioIR4/WUxZDAEHMX1WvcnQgBJYiUIsfRaYYx+EZmIAdBEUsKlPcER7uGJWsu/N
6Ndu636vp4mMFltzLk1B44pGVlGAUeUkSn9gsIy0MdIiB6FJIMi5SvqAHOcjRsDq
pe/3xV6ZqPpTxsUJl0mO01iowcOI35uizqbqKBDKN2/VlIhVyfXZKUj6VGBkE3wD
sAbNRd1exNMIVkv6/dvcCLonkIG+ep5fqCFGyhEX3WCz11E5LgR65lPjiFpVbUuE
pSQ57km5raXpzmob/jboWhiFJn1RVq0HSl9taSoESF3mjbRwkHbYh1L/AbGLj1qC
NG/rUUPo9B/LBXtOlGsmyr6j9HEoP/DU/VhusS0TU+IMpafwTmMAJvOGNYzp1cOW
g8Auo9YYyWb/qQmibAAOXNZAys40mddDIT6Rlslp6MAa4vyWVzlJHwCdl7xIRD+S
lRbduUQ9jhzG2euU10W4al5hPITC0J09sEBxoMFjSnxGamYF3UKUSa1tgJDSB5IP
0F4l5UxvzusNE/CDgk/gIcBMJo7nrCBx4koM6NDolCjlqGc/2QLe+rC+6LDuNHE2
TXo/+mRiqqLy756UocQF4VlyEkvLJm/nIlwRVWEY4TlFCQCfYxURC8rASDsYVP1V
+O4T01GJeVbO4zu/2UJyKnNAopQppCGo97zIgSSZisurkZmVFI1cG3APpVODjAGy
WnkXZlbc7Uw3GrmiD+jFCvyALFD95I4mz6YtlUTXaQdMA9SSwtpnzuUI3Tp1g6+J
P2Zio2aIPkdyUIRj+GR+/7ZPljlDGtBZrzCdvgM1BEKiAHv2QGfYqB6JVlfBVKsa
YBYovuZwJ4LCJXy/ctedfvND5QdO13jrcaFCvmp9v4XTWA8d5aKtZClUqX1gBJth
RLItqAIc+Nj3YDpmH5RHpZK8mu3hxb+Ob2gUyl2I0lp/AezDe4HRUjwK3sMXxIsm
w/+lrruThis7+/UW+qhZVywuqjlc+QCFW6BFVZieBNDDxFIHnihsTFDa8uaG3qsB
t0r+N3euLU34XfgpKuQpGz249ApvU0vqeKsY8KnPFJ90P1vXcpaGv12s7bI9uZsi
srEoc8sGJolA7SFBYfvs59h0Hh+nFOpPuV2UeFrwP0da90MilV9Z8alWo62jSvgK
tw4NalxJrkL0SFopQGf+kQDpRLM/Vh7SLsXolGa0uDLm9I6uCRD0VPzXiqB5BSV9
i+uej7bZ+f18EE+Eq0E6mzG+0XWYVlSgOp8dhcvoSFa+rL1H764R+lQEnCpSzJO+
ehLlsou5EX7iH9mn5tXXz0VbAJKxtcVVSN/2sqXYaIMP7Ms8nKM94B1bPOyTzuiX
kbnUwR3B5HZZBvDMaKynjj0xccXydMu/HTDDN1GlRlaPqsMJaxBbETK0p+rSGn5B
ccGtPqMEdCe3bP7razVAn5qgJb2jPsKb29QvqC2L8x64PCHreUeKsdcZkDqYczOZ
l3zSQvg/OVcHKR05ycA1OS+yITdCPBn71G0Wib7rl7xgwZX9G5i6E/I4mBCZThE1
DAyNLKzp5dO0UkTvL282AVL2TGRJnj1AGGVvztkoYLhKFahm3B9v3u4++TGSEwvn
8RldqNISTc8jPJ6vmswhEPWZpky+/UNM+tn5IbB9Qu0grKZPfXr4MhL1lND70G0L
OFMi/JrA49gdZCcDGrZU0ogm/Ijqr/CKMW2wDZgZHvX2K3fmqlkE9X8+9/8ymTu0
G8RDJwYj515+x8foktXRnK9H5DhGEkW0fVn67wpn7/xSlcD9ZlDGnBeYat0GXBOk
Ua99djyCvwBFhM6UjDoxejXfvEp1pyEFUqGa92WBiwnZlQe8Cmz1ysshmMczqloy
zHtNPIpPDi8DfC+SxI7pg1EfsilX9iJePqDdA64GHj5op0+LLhVxVhuYURnZGrmn
fD0lUAn+Lj49II9JRTPSvUXJK0Q+Z0chU7JVgDDp8QpIYBU9ndWV9Ub7R1wnnT6/
YbinD6APwPBuB1Nh8OhoFWBhlwfnujsCDJkE55G8OXvEcqfB7Nju7mPifFPxZNS2
Lt/NGxqnDHzAs1YDN67fsZ5prgxLglgS6OTUwU0p836Co8wJgolBhWNkHTfmfKzM
fItbQCU2c/xics5U0azGUY60jb9+/0JE4McSOffX2NQo+IstUWsRBPpqw9HyDQYO
+Q1Im7O2puiB+GgvVKC5WZgaW7ATRNbFzIEminn4j8ZJ2/2PpGDYfQc3K+yfIzc7
xgBFV8DVfP0RkdtIIE64fudJuz2b240MzTWZvkX0mFT1wfCUUuSXUFr8TbJrU7Zt
fUYFAr7VLIXrmnHWFwLqLXvPkWK98frv8ABFI1Mfr8CGu13OaVsqapynz6nKjcWA
VO/PGPkPm/ZkQwHDB6ew9DVRVFXWKCa9dai/2fLvzpu1et1wSV/Pz/3/nQZN+Y2G
dZp4JnV+Qk6mycYZk3jIiq1S0WD0jCeNpu7/LUEsmOE1CTUu3Rig5/FVknX920mr
1d/Vli6Sd/Yf8l14Phy/2yj1ew0BaaUfGIXtVhvw0FxhbxDG0OCFjHl+i+gEsHgi
U5T7g/8c4YqZfifb60pmyyaRO+k8sfn0FCo2RwjHFnnrCoZjJC5oukpT98CaY+E+
4jdqK0wEGCSpObY7OArDLFH1KhDaiSyrlE41LPrHmTad6TgJ1hc2V+l5fGjfD403
o3zlcGRyHf4iMV0C7XLhCeRr/B3McLAQ+hOs3axFbvcDkI4IJ+yOTrr6HiYBBQH9
mVgdLID/Tslib/L2jw69g5ggpgq51kOGYX1jQQfY4OklxNDmekZ+ZuvhWXVio1Tq
b9jstiAur+xn7vPYYZqF7ycI9UQrzxwtvfzSiGZIRvRQRB6T76lb53EcJ3pPbLXy
+/hn6a53JPjR/aMUu1fJJNzLoSmEHbVCa0pqNC2oJTBwK7NwAppSNEAEp7Dqm1lk
oI9USyKMFEsYWqKEvgcHTXFiEHHaB3f6RakuM7PDdcOfb9Usg8VeIHr1/SA74InD
UwFtrPuFr7Bq4W7Z0aFDi5RP+BhXlEoyHz1Q44nZjm/VyyTitc/qZMzghbhgAgJo
qR+opcaZIrgd9Xg37zYePdODfo+VCsgRiZMB9Kb4JVwENWUiZ4bDibOmUYMNoG9h
C2L87IWJBwFR7eB/RDJDqi2fgpy6cwknonF6ahKwur+Fz4W4QIy+WD4RX3LEq3nw
mObA1ND90Hk1rmqKZKVijQhb+Nx23e23VVxge9kBhu5cbb0pJoJXKuYI4JAwNnNQ
5TnWhXV955uShj2nx6eMFLAlh38WxRFBMKBracrsHHtnk5duK3vUHqwL6JaBrh6K
pA6cGJPmUc5q0fonkcisMro9vb0wJjZAA+2qEGp6KNHCJAGq5LodWLcY2k7LT7Yv
PLwgjX1UYij78Fkx7CEzO+oizBhx9DkcqB6JdooxCG8GxIMJc65OFQxsWaQ3VzQW
JEbjMZQ7BpiUHM6f7TBvn9dbiJjGz5C1rGDC/hX9ec22TWN4YsxBtrjeER6gAmyn
R1AS484mkq9qMkNTo9JZu3S6+E4Eyg70pspGJKRFCK32TdGHa1/CJda1mqre6Iex
j9Z+01jhHaKryfkOEluuGpetn5zLBNZj7PsndDaevKBYHKA6JzYdPwr986nNCeLA
tmtg4damVvjWM3Ww55gWl76ZaGiBEjC2KJ7lrTrzt7Zg0ob1WvjK70dVOn8LTGt8
7ikEmnmu3aEm9MADfDBR+D8lEszyZFbhuh/s4By3PKtKggkI9ZY2iB2Fs1jIb70X
xo4DvSXhCeLDlU1cLbuT7e+Agey2l08XUWzWTH7NCJOs7bjo2Db13DdrT6rCtKyw
Uby8dcxo11MPAirN6o5ZIjRhGCW9SopCPKEqmbfmXIFHuOgTxczobM8MiP+pQKra
FnxoOoAipa6hdKjy1OMWZI0/pkq36TXhkUwLXJ05yTtDZI35KFrE3HE9yXAbmqEA
dE6nQsgMcPKEYzCceV/YA4PwEOWQqVBVhT323my8HjV4uvy/GTcWRzjr0tVMwceL
FmgRrSleMGJ1iWOBSTSEHYEVcJ6ApExX3kP7Hz1BmIP3aNb7oPI02bEz99dsE90E
GmP0Ji6Q1rwX5cN/InK6hhM+wOFrrgUeqnudJgTu1NeBUUJlzG7oqB10/eDjdiEZ
OhxIN8auIhd2AH9RkLP5lqw9NVfhGqA6Ec0u+RdX4gyBavLc31vl0SBd6RJujwFY
WJF0C8yRNiPLxNfcoTIq1xOzezXVV72QpAtSk2cttR4osHhNk0yk8t4+Syjb+O2h
9aeoR0V7Dx4hdtkGJjiKdG4CrVu1CmTr6ALFohgdSWOxXiKgNJO2kAR1tOmGwV//
PPBE3+5yGYQTyEfcQRln0wAc33G7ovnjXwVjBubS36emNkPzAkyhL1dct/gRa20j
QBr55GLPaPJ/ZigqQGCL1nPBgVmLlydg+APAyd6X01Osl4AH/N1DudR2JjuurQa0
tVgOZXkxXokD9TOC7oK+R+1S+Sn3ERmOXl0YJxlmKgutDlyw0fSBanL95OWAdz+g
8QPZRtjjB0FVB/N3jrEIzu09qwjxtDrkDdLEkv4D2zjcthd7X3QmJdWY7XS3KzNk
ERLPqvWM5BuFiBTG9usw+nS4uRzPfqvHmKXEsZ0a73cOBJ+d5kHR0dawn5itnRhD
a/Rv6LqpLNbMJD0SOcpqa89zgAkyBadJ7HeMGn7RMEKiQubEOmTFkpJTwUSCLnyL
SHceaj63/dNN4fazBRP/BT1Y+xHVa3/5ildgQDp/2oeuRAHNVYmB5jpN360m0sp9
jd5umXDeS1KpeU1fs9d9lAE2GpGZCOaMprj71r59xPYA6GTX5m48pDcUVbpPSC6z
p2sWkDCwz4mdKPdjKsdfHdr52ZQ+/YK2D/x1BogbwGyMvlBcj2Bkl3Bu+wwGHnc3
rE49yst3SMtphgIroqudyiX8SAvVsu+XLPvGH8240wHcp6ZFzfZGcL25DO8SqYSt
5m68n7YVCGMr+xvnrgYD1g0Vz7TUiRfotVjFqEVVmSIDdSprbqFf8lPB264dlkrX
JQoyYGpxsjFXBv98mqVRp89GwuqRZz84d8rQRKbEx0LohysNqSpv5PNOQ1eV6c4B
B4Irc7kTM9zEPmkkgr00owpkjqTVTdxoKLR7TFTvzXY5p+B3zwSD35lpp/Fh76JC
xI8fbm4NaLe6gBpBykIyXcfi3JuOS4piAsu+8B5O+yWGeWeyzFP72LhExVXs/m+4
ZoCWZNdjQdDwlj2q0NCc6GaKZKwmdcYmaV/nppNATeZkKlTTn0e2clLLgQM+6/M5
INOT1hWLM1OwazsMLKoNOAImpD51jhgJjUp0jSY0JBlPhODDYkXPOR50KjIUCoz/
s6MdqSxofr21v5vHsfRpn0nTBwp86YtBWnyr8OY2nMdgEChhlgSoaLaRqg9YsCXB
WhguRyKhV0FQGLGCYjYzlDTysJkxQbxKTQ3LpSnDxhjuSuRX5fY4BhATgKL6Ib8I
Za/o6no4d7dHXDCr7QB2LoKoR4FkUC25zkuGeu95EgIftuY5K7yy26MvN77IiH8n
tmEVV9AzMqvzj+8rFYbZx6EZm6IHtmZYz4gs7tc6X/oecFHJVKqyiIP25g3XhyyW
kAPHjRJ5UKgyoMaWFo+SwF0EpYPXvDsHjwKIVV+NLpHh5q4iEb5/BJnLcTKr5/sJ
3E+bzv4QPn8iy7t5X+FCpqpXNb1p/krDDuFZ7ieQ07sWvh2xZjzX31l7sv5fZxQI
Nyj5JgR1Eb+WX1gY6XAES4UYgsXlOyvmIScIK3D8BR/8U6QunxxejT9VCWRd/4pr
nHe+xp2zdbOdv9uWjCRH9RJW6QcVavNw1Z3kQDLeU45xWE5tg68NRYEiziVd0jXz
0pPNgBlcDD2qhmkVQIMybqDMmGkKbydBbkq5UcjuHp8g+A8RuxSsO+tKxKfE3F5Z
vSF4C93zLhL87mEpDTkkklUHP3KBszQDsOqKrsVjqDEp/OdXPPHty50FNYT00vVS
bL4u65QP1jsttbdHOI+SxBiEaQdJgtYaL5ak5OX6oZehT9FNX3vELvsyOpP4bsFl
NQzS7rQh/5tf71BRqcEnEpLVCN7cD8zA0OX+z5fthBiOc4rNkPs+wJpRYchpBMDR
tsw/uJp8SsiJ+LiGDB6eQyf7Ghgir4PZ9xMdCUamVYNjXSXEK97Eo5H3mhPsa4Wp
uF4Z/8JgFsjoaSR3Mso1rcGAUWPQjbfYBRJj6JOEkHgiGUiRltXBFPVobng8RL/B
uC85eAOa53KqGfZxUE2vSHurE1ydg2MEITux43Btqww3hXzmvysJAc94qbFTyJ+G
X7xWnvrsc/+jDEDM/EwEB0DhfgsbV2hSrMuV6RL4GuH6biCKu19BCXv/STuFphC1
jeH6V/937oGsUKNOkU8M663jgMHySyja2WdV6j+3RjHF8dGcyRNoCobZ5AAC+tQi
JV/yxj6O/uszjDQAuKGQJNUJmV0roVV3gxhdrlWzxbi2lGGMHaUONSbk5RvUrrzB
tUE1mrM9cNMN9CYwgkoSiQXphNFdPk/ZHaIH6fbfuWdATEclmN6yPUh78gaQbQth
aWYA9k5kC4KLTWSvs0eAdHNyvy99z21nIQCz4UnwQH9yC9T7dYZ1KM3myq51fsSO
+gePDdwq/1xj4ulhlGriogNOt5jbl5SD3h39kT1c0Tk2IGs4PUkqr0jPXzxVoYpk
W2xjBtDd8OTRSHj36zg0aojhE4Z0aZhQQuULV1j2UsEnym9assSTlyXzXSWAMqEc
bhCusif01Vyo+IRNViuAijGBcRXYkpTKVMPUlmijRiFmDS2Xsdo9Hjzb6zh08MRJ
YMeyF8owjIJ2NFFiAK2Slcoq1FR1KhLj5w305Eyo2McgXZppK0dGk6CjO/p8+kYq
wOuyfJcT6sPJwVmniOKn1Ll3n6YGX0XUSJAxHdPZvn5Jpgv/QuJnJDOW1y/0L85R
tDf8Jet7MI2erOThYWbe+eU84bJo6GOTMMuE9WxMlmoErAqQkxJ+Od7rvg6zKbRF
5Jru/XlVcjvr++9cV5WMzDwwpVunCAFJJk+8uwka97Y/DG/Zm4mk+AEg9szRjaTE
3LvOkaWjIuWKYxx5CrZ4Am62zT8w1CB+QlL9nfS2zHc8Y9KEhMP44nyRUOjXeukn
vDj3SfORMwYBlmYJnz6XthJf6OVxBDFcFmRF6eojOV7Oy++mUf3WTAiKAK8h1//w
F/Cj7z1RqdZOs+cm9wmhQoTrY1aIq58pKje012CpJqq+QuAB3ynhv9w0113Sdzd0
RA43SH6BuMM7MtnLjL8Y4wf+y30ac3qveIh2b9TGJUXgE9gt++FoIJEwQIfhHIF8
EQ/ef6kw1IB19kN3GebfaCaK9NCFm8OfpZpdtkzEDXJrDLvsNh0FV0Q7kPtcuwyi
1YUfuLkdJDXGQDF8QQg4gOdjs7N8DltElT6U0flosNhRAcCqD9/9VOxg1KAjHGFD
D9cDevNaEJrW//7kO2iPOzZtAzKqiCeakPcXuBB7kgdAelAlNv9oVs8SCFiTz7//
WnWI04pyQ6i4gE3tBT4ZDff2VM0C61njAyY+WRwOGULomNadYHUiuxTIlYI9ZeNE
r1xrw0I2CMBjih7KoW7lpb8D7eTsLHVKrH2JjuELXheExY9Rrt0l3JNGM7abLguL
nuJFhkj9Glg+M5qjJzzvHludB4jUAvDf8nXe1CLwYJLtp58qHWBK208f1eH2xI+f
CDrcf4zXovKPeCj1KJSOoRHVLg6vc1tDwtNTsRNJoQYEMp93p+RFyR3lYxofri3N
4i9jdKx+1Jc65MgTbc1ASHpdrC7LspScRpHWcPRHhthAiWoWoGhXLlucziH29Fhh
r0g2Vy1ZYPCy/7qazbQJI+cV6H2gz5InHkZzwi+M11f+doiYVIgKyUWh4xlKu3no
zcIxmsBvMl7eQovZdDWxTxd0mU5wHkAAajYwmYvvh60WvY0ElFGoPwlYsFWXsPP2
e22+Lx/bBxjc0OyKoO87Bj7TIz0z4/vgg1U5tqYOE1aEISIcCdhz3QmeNKtutuzY
RVqtvZIdlNvJjE7+PjOxYke/Fhvtm3z+/SGGqpHElA4IBRUgxpJp2CdaoBWEpWXF
qJOXyRZa2nQ2B7g9s9lYupPzBk8gzUz71/o0b3/zmRj7PKZI7GqdTqTBJ5tC62qd
UyjKA1JhRkNEcp+2/rYlLLJ82WBpG2xF+9J76ofikuJuC09shlJf7rBl7pMv7s86
KfOjuzJe3MXICn+HmNgrxxkkecf2YdUYWEmUHtDL5AogoZqrEi4SkvSuJCmB2dPp
8uRgdQ3pH8Tjcl14vaVArFeupl34ZhXn2OXw+pATAd3q4YVORKNJa0XaBa1OH36a
EMxowb04XAKM9Yj75MExYGYXgEfGrJLxqrgywPhyM16B/tUONvrKqXcaNAw1bbAU
OJYm6lStFQYEm738Fnm0SQg/B4G6xhLXev1kHtf1puYD92M60gGUafs6vHbLiRZ7
Eb/75ha/vPMYMS3lQwUEJIIPOow2jhHUUcnZ8F1Vd6Dlv/dHuPDoBjzivR22iSj5
EHOhNwLYR/attggFvf0LqATNEKF6GDpGj9qGiqLbP5V9qAEs98mLjG64KdGvhEXi
hw04UUKHkMoMBOLsfkKaI/XGGa4iRGo7KpborqQPwt5p+ia9XXaq7sTLtQ4dhKin
w7CaoRacDEi/5IVwPTUeG4vAAcpxc/LJK8SODiuk2A0phiSwpuw4SZnI4lxHpIqQ
Z4xm21exZ5bETrNdlRWWutecW4PQ6qiTRuOlStoOiM8i270puq3dSHIEPe89iddn
zXqtISro8atTq2gBMYH1mO0XIT+bgc6+JXN+K7aayAaEJtU5ZSJ48Bwz1hnDx+qF
6mLwJIRucUQ53i3d/uXkms9FExutHmsn/7P4S52ZUsErJ2rvsFSfrnkNvVqYb4iw
O9lajmGr8BnxiWiS84mZ2alypFYagG9F0icDa/Pn5j9RDT7vWl7/cevxDcsTwxA7
ffbOePvJckntDeJnBiKlTvQQ9fjeKNZ3mzI+joTa1wtkeSnqHm76+XXwS10tluRZ
wY0dWmmdNE5YM7gyv7FXMDRKB2svAmXgCDw8luslauS/eQAxfsEQI1OM1ksY598c
WyBwLTo2AaDz9KD7pnimYJv9FloQUQHP+ard4TjvIRtvSLxm4I5GOGAMYr5syYyQ
o1BawKPUCPa+zuOvxXurP2xiIgJ9D1ne/d+C+ZjTo4FkAjlbTrJ9XSqLgYck59Eq
bpIu0thNDsYHa5/THQdzC4umArtmYsS8RhZcmb+CmhuTTC73As871FHICtwWjLQJ
+xLaJGp8i3PKHP0SNlnbJYwLtAGZJsoupYC8UPACSyr9gUkhSUHn5bnVmdj6oEDs
84emwCn3aYGdW7o2T1qp05DZm3xJqMt+9JrxPkkhhlMOMGwD3tx+xNrsA4xQGxwK
2xbcYX/ukfK0LF7bsQl4y+0w2bxLRl3nE5QDf9he5h2xD1tjL+S1ptr0ZKYbAtnB
P2FaM2b/fMAGQooV57PZGPDYbp8Pla+ZTMp2BNsMrKq2DOhj49yn8+6tv9rCippo
HkdsG20abmPfpP1cq3p/CBM/rWKZu441BXhEzCLqBu5PrIDSC1VEHSDhPONX4osg
7OAOARyd8Cjw5KK7cgB3wB7zEGmG+vq2Dh2ZpnO+euM/Eto4DEO0DH3PU0WkpKP4
jx3Dxvx43+E46KLKAlMUjnymclQxOLrm15d1CtL+iWuproKoE/00glwpLQ0rP/fi
5j/d1V19YbiGe8GN+oUhtslgYUOPfHyPOpZaixdNDOZIPsf2fMyhtIFqfgLZbt/F
mofJApqDjUT8ZSuxDM3aHWlqoeP20nK+1g3LVm+s0tMjcc60jLDZgiBBZsEMB3jR
6Thm6FuwVm8mZh5jpM7ScNlo1WmjzPqDchJHFEpBx4/VEJcPiOETacu4ZdbFIA1z
ZLjZoGTi8TwVdUPmxHWqnjORZR0l6hnP89X6MSWgo5DLJo3arde7dLJ/Y2eccVqG
OecgdEbyetNKBPyFjLd8QpE9EyfYybfe2HaxnBGw010u6hCE3Ky0Aa3zbS3/xFRV
hjtktxet7Nl1cqzYh4iY32uDY+EuCx4jtwzTcbd7NJhAZ3XZOwjL2dmFiN/gZXWh
PDcmKTVFRBPgR7urQD9Wdga7KtdO2jVwNFOyXsHUBIuAQrJU4RhXYOBipubPqWND
7GdtCQSiEpSUzQaiaTV5wiLUUNugmYw974bLww6Bwn244SwMwSZaZsGz8cRB+04D
4FHcvtuZzQX3i4TqyAlS1izir6YEYn9XXOhyFSpXmtyxPI/xPu/ht0+8RFlqPRhz
7WW/SlHnJ69XCzoJgcKmFKRW4lwwS2WBKr4B8pHqXWNtgEfKq82FJQ3+u4mSf+aM
JqoOzfx7kUXAtw6mZMKuKIPvGPzzqoAo8LtQhREewF3GUIqSmqC6eCB65mg/FMFi
3jB8gh6X/N0hOjJ0/nrhtp+zhzxCiynXTOpth8AxF36BbJVz2HClyf1U7H1O2ZrF
vgMxrHAYjkS/xmRFF08DzEZJEYdWt7bAYs5TdiijXLcLz2i1XKCtHvN2ZpxBdqp0
mgVKb+UV8HjJwH+vcYFSQ8X5rJu/INK/Ofz0r7A6djRL9dDx1DfktwhYl1tCElmZ
I5sGdmnqtM7c6dg71aViXJI6FlbhMZqclfdo0coSKRxTIx2LnIn12T8Mlx6MawNU
HvWBPyKFu5a0rPHT8Bna5kjDGm2v2qWOdvCVfoP5T8TfBAeaOF7/NFuac2Zx297S
mP419VItu2NljYGHr3IpLUwrrmLHNGy4iq0C1ESVlfVS8VIaEFjS7JmV8Dvq56xH
W66fEPXwGsK+SaJd+0vwV50bqerpxJgbKywagF1SwvlIUkGP7wGb/yPpttYdvb2q
pZd+TrwXPV9BVKaUBZiwNijXG9RZQX/t2NUAoBKeInUU3D9PdOL0r3hZQtf6z1C1
wLQ4Pn7sqTLdhwXWPTgW74NzV+lgvG32crcvOQrgA60OjaRYW1KHdC93cAxCw+6y
GZVkw5WOM8hoJ0WBzjDIMgSJ1xFiACLYx5rLQx/Zsu4Zi4H8Ec5+iInGQYOUvmuq
+XfcTIyjbmFA9ExGtz+2bRg7lWiYLa8GzKXEDda2zOmJW5EVz7UIlfvvgVSf3hGG
3/Rg5/dxL8zHWhra82XBExzJGcnm+dYtLcaufOS3GGkpXnha5Y1+ggEsO8jASOe6
TB4WyM9zCHL38/Yl21lPxQMNqjitc7A3ybqSNZ8N79ViEYHt1gcD8XOqzVs7xsur
iGSI+MVZ4NlHKLdegutOzX4RbuMBzMT0BpOcOjttshlSOb1CFvywKrZCxUBY8Wc5
VDhIPYSGuNugcnWu656iFKc9n7pOjAx+ysGlsvBI/db7PWoH5sG4Ui4MZhg+0d1F
il8gYBIha1GsttXD9cSabUgeB3XoZZeHJaw1qb+Xfv8GM/ER8XuPTv4nvZlGGrh/
iazICSXZhWYFm6XXEwemkvKiNIGoDW9nE09aOu4k8YjscqLSq01lJHYvCSzE4HJi
JqGH/Yjb1xH+rT9PUWsMVs/mcY26v5USVLtkksYxRhvu/r0a8EJPTAqnujaPmF+I
g8AYzvr5gZ0AIjQxF+smG4RXJuKVj9fNWdEpSYPYV6OueLQrgwRaAjzBbfFIbyIw
BcFxz1HYktCmlCqCnESkihoy6nd5IlhKxLfNlHIrEfYgGdCvEtQwslLeKuAVEv6l
q9Pb2Q2PkcHiyyESe7oLWFBJ5rMQa1fKg7TkA7xVfvRG2wb2Vt+xyH5DkKhWaUeo
8gSzQar9VHfjo5tXwbAaTBdhLfifc2mSpGlk3QkSDN+2ti30BK5TOER1AovM8UDP
tj3XcHLFNTE3ni0AdQ/FS/gIg5P/wyWk+0q8t6/B1FSaYYkaoUDn95/o1pDtCAJV
y1kB5YhgTXnTKwlqJIMZKO2HRR2U4MQjV/dqmqSYFiVQTqX/5J2eLcyrYe0FBhyk
S+6/Xbh+Cx/AYjrc8fYFq1OZvjBRBet478dPyVmGpdsZrh0h77WZm8HMDWUxSq1O
pYMepOT6L9KdTPuAkKIEU+aru9UPMPv1AEHevd3BFxbUOlkObQfTgNFRAsZ96PCN
DTdRLNelZzKzgYyCAuTDXcobKe9qoklvYS4yoGvykaYyi+HS7c9fQtx/jYiGOOyo
MC5Da0o6i6fm3dWNBhOtWt6px+bKE0XmI2clG8Uj8swAzQ0OXkxtcFWURMwReYgW
V8vEyhh12Q6vouR8RvRj8z7b6759zlLtlMvut2bur9RfPO4/9o/aIW3IU62vBR78
aGac8fJYV+BZathSHXOmKm9zISyYxulwJ/xFdUeqXvFuvMYoqahmdXQVyeEuWe3i
evJGTZ7Ag70/TVMnkF6VbHAID4DS3FXQsjjnzMYvFpjacR56/0BdVuBZIkULWdaq
At+Ip1sNM+aHmZsTatHx8nycnsJ6uJwgFWbsTjNWxisqZ2Tqp8acR1i+kE2MBv+T
4vLHZP4FUiAPcDRFDQ5h0e0cCje39bZxOxTWB4CqCIlCxZaMgsOCVPtklNez84GQ
+YbL5GKk7cjaGnGHNHhU9zYR0fBNgoHgTl7TDZv92rZQK0dUM2STMgb38cvPEA6L
4AL5mD189pMVFFbGBhh11uAfgW8bTFvAzx6/C9IQcVaQIu7MRQRJQ+9gkdKEV67K
MQpv8mEMOm6K46CXpkKnYyBRlrfFsOk9Swnj85c87eazbBFT8mlI+F9ygC/TYu/x
NnVYLGfp9q64WYJv6MU52E2mtVP8YdTKZEdKTHY6sygPn+B6zdAThO5z7Vqdc7x6
lmLFyBoj9IAjYSePkpFGj9J6TxMtYLxlYr7y9+7HYMkldw0qufAkoSVYK+guqL84
753I75BEH4gl3Yh8RloFbp1a/OJcYfbVkcUuYkLBGzJ0H6C8mYvt6D3QFJ3sJP4B
nKXHaJNuCMveFdFtLkjNZrHvk1BMLoRXlpO34fyDhctFUlzH/zheyDgBEhN1O+tU
pf61lrWsRlTgSf3emAGGq8A7nkCBfvrmDHJ3r/j/Bi+F9J6/mTI1ccRUpwgh1+Qr
BYME+A//MjFbusn6UuMI/z6kYaGzwlROg5ErNKgV+6mrh3NeFSXRLIaoKjZqvzTo
9Q3kkhzruTQQwj2ocxXdVlfvkcKPixeLDioVfvOeH5jF0chsx3Sf9p+bR9AHqJO3
PJ6fNMxHSC1WTKKSkl30dHovm7Onol9mMj4ybjEtOPOY5kRufnvSjVr7ENJfsxYJ
2Z1do0clXrNMIXVy6Yw8y397PeHQFqPV1h4lwQ/f4ReN2T335bKla20BHvmRK8Rt
hTZwbyCueLIOdrhlVP6adUbpkKv+HG7h9iCC4zx9Q8aRo2r5NImO07kKdWnVIsrq
kaxWGTbqCAgDJfcPt9Qrn+q0iegrC+H4eEi4WWYuc8kWx+D4nof1R30Yg5ziWOpp
8m4d1EluREHad9ND/yACdTUsWb0uUeIBXt+lBcNJbpgs7cJSJofEkX+VN3jsfGtW
OR64pLkevY8hcDMjVMm25R6gUwZ2pXvUzMN8VXrLNJFBxZl3QnPujlHLpXZH4hvc
j56wygSOd0bWkFiMMVdzSbRuBCv6F2QEy3VWLg5gBbsBtN4q0NV0IOHdmQkr0i22
eVub7xov9S7C0Kw6VFTY6shF7b1rk5E6hg8gFlnUInI2hbeKEe663I9OrMWyquAC
D92zKerO+/ZMCqcJgba1JGamgWDUI5Wk1bel8me4IyRTrW02DW4Mq7ThfPmSzZXq
0vEvRktBjkmUK57BcYnB6x/8xmlReKrr7OZ1AY61le/CKR+uklmoeFWPLq1QjsUV
J5Udp8210N5FDI+auhX3bV8dqKCXj0IBzk+IWuHYY5vF28J46EA0dR02TlDEC8x0
nNM4J5+uHk3wyhrZVHQlRgXA7EVedwIuFu/SK2KzGaRt+Ha7UO6M9eKpa972KarK
/Z6jJiqo6gbjQTzFtqa3Xn1LgVrQsh157fTuvjGuV5uWS3YRqtZeVYKZJC08wk+r
jyd0n43OjiEMzJzHG/6tXA/fmf6A1Bq9OIZVp+T7wVirwDJFiUYX+Bs0mA9jj41N
C3nyS2tQergjvSdxlvwu5K1mm7Rym8Or82bzPtxa9oFGCRqo8cg3TFyRtqKhao0E
rSP84vwYBJmqrqb1fh/DcZPzWC/Cep6Um0rmrAqPPJ5dyG6e7qflVa+B9W8vjgbA
UW7E8FvcNssyhBbxWmALMqGIV7gU3UqoRvDl0JquFtorq/EW0Ru86lTt51/aExF9
LWZNqDhO5J6eA8/lcy2S7vZph+rhX8UDVOeTF5mmOwTxunx3IEMu+z8aC3rob6PR
FtbgWm+gjteihiyOW8kMvFZlinwdO2KE/zGsgbkZ/gRo+wpA19iyrjnYhOBo/wlf
vcuWqII2XlhLkVjQvjBb8frUXuJ7BzrYQLkqsi1v4ESMmF2II5mL3w/3PRwWp97p
6FPQY6OXEOynwKfNEE4cBe+JFoom1NeLsxVedwXOxkmmAlWqSpGVzUGBtJU0ci8q
0MwgbljezWFGDPN30f6Ea35cTA7XYatu6sQtaPxE+riLqBVuq/9/3XO4E+jOyniA
Lnt4GSx3C6iSwXdNrb6ycl7EqaR6PkQyiWefGNjZaOJ9mkpdE5L+jXgkOGDglgCj
3A1T6F5rqcxy2zMsc77MtcCnXQnXah10XaatooiG+O0ROjb5dGSowgn3xtBd3sIm
p56kpFLAWsg3aCrUoggVfcYpjcYHiy6Mco9PpEwptWKXIMAHwbk7+zkgK+ck5VF9
cthL+Vsj6x0GPXGsgScosFj9rmHN/14SgkxdvZXHd6LMgnurRRZOehimjL4fRCDW
74QSqeFKkQ7lDUpB6rucJUnhPvl4fMzSkYktFilw1WROEdZSRkm251Qk24cs+HBG
ZsZAL/2Ipn8qy+MGIfY/+X2HOvV4aniL/49riQfZi22dzmP2iGUN61IRacy0fZ2e
HD+gD3YlUK+wSzvp1LFUAIUMoD2mAOpa2yxhSWOWem58dbIx0NwZuFfEdXS9BmG9
h1c53tDABkos7TDeIR8ufTmvhrXIoEhDukX3hGt/DQPANPdLlDIafbjS3YbXI690
a3MGHjk/ZvO347zdyfNG+i8szW7Dr8SEjo5XVflEi3u8laMMXLZhc5ETF0RkJkl6
G1wJA3UcsIH0K7tuHAN0GQNqXqdUNKrbyl7yEXMU9vinuYh8pz5hCE5woMSbvTuZ
VXIOxTs0cjlizXB59/FwDKitXM/eHESmgeP8GTG9bNy3m9skL7+YfIViZ01PaT/7
f/x0Jq+LRwgNHXuEqOtI1w6YH73U8hM+6rqN0gI9ozc8c6qPSRL19866KO4Y6ggF
FrqgKYfSF0lMdUYiXjAGdLM0IQoOWek5K4fhiL9/8x/5KCCcVDpjiJdKgYxJ8IKN
9O0iI/Ubg8iI+NYgXjaIaNWbGqj6mZHsCQBAtICWVdcDvqZiv+MFPzG8WFfAHzFW
AFtp6iWNId2fkwusuj052AdMCXAAkw+9ZoNVGMHozacAGmtHDDiZNvW519ZgWAN8
+WIybYIhgqP8PG9N5f9jwYmyHitTGnovbFvVFA9SlRezfQfOEyqWtSYN9WQI8xQP
GXmVk7Zg+pUFZRHPHrOrLlemFbbQhqqo7XTuj1S2sz6vdO+2nBazkH3kmmkgLI99
//hwfiBRanBc6oEHinJeymwmiqb+KP4NAaOrBZwoSdcCLxymkqVzLWpI+WqCPW2+
umcMvrZ5doQzzqaseVLpcygNb+vNs4GtWO3h3zuI+FAcX0Pj6IRAAM3wvFATC4dQ
6gMADJduQL3eo7FfsC7kEY8CwAErX41mKCduGw7Qrx+gNBaOxqasvslTjv3SNs8Q
I0uUyB6nJ2U4xcd7zL+DLV8OZ7feDKdj3RXePIsfCvpNB3Vq+Z5Dq0znIHJhbcMI
Nl4pcnfTsuF7ZhpjwLl3efhGuEHValljZGBlF8Jj7JJyQn/WR4oGCkKCpUJBd7rc
Hw2GpdYTJS1KA/AnjL0ce90QkZTUkL94TTXBGxwI0E9zCa3BmEK+l/nmCizfbDOH
ZnxXlqyibnNvYIzUGLdDADwFc5OoGpIRj32KNyneFHTf0M6RnXx4Oo4+BLHLRIXm
RVib9Dz79SKXWti1/Jwok8MnlcF/CwuxWOO/Ald7sSZI1XC+zB9jJmGXa0uK7owP
3NMkKK7UkAD9K++VdBz2PT4UBEQ9+M5M5FFqqExSvNVmNAzsZQlpFhQdjwwXn6FZ
jMr9rbpmVAFPUCvWgEA1OYmnNx0iHERBBqj2KahWSH3nAkE4EqSs6jYl+ESFHJ5P
mYs4qdJ0A3MBXyxBfa3DS8la9X9EjY5+vO95T39FQT3HJmb6yJiI+HXip4C/U2xA
jVR2mjJbTJRuw2BVXJUErswrkaj77sz4QdYckMV4tiv2N/ROUG730eFB8ohyK+VX
3AyJn+rmpLFEXSbgJNVKrY1aPOZSdLNk2vW6XTKMF0tVL7q7E+fVNYAT/sSXYO+U
2y/e50+OtL0GqtEUPFzuoIy7o6F7MdJp+v0vQiZ74hgqbbDsNPukc/K3SJq5RKG3
38HwKS93t3fb6J9ASLaqxUKsEWROeviX0gZK9ZCGSC6+l3PAXuuecHt/oCGhlKS+
4cCXAlTE/1Uz2ay1hELmVfLiD01Yz53lsLpoLl+EkxTohR+b9V3E9vXSgDl5nMa7
Yy6fJTwDNDQ1HGmNVCHMqw+U9gWVnz26mMJYfsN7QHK805hdQa1pGU941XmzSJWg
RGJhoMpd8E6kv038rhH3gVsEm1X4rchbAybhL2cNJUV2iWFnYj8OronqxGCWw9eX
uZEcw3xxzCx9kPauK1VfehuZzC7YnNZTR4FxpuG5JpDWBtXNeFjvUlI/g7AU/aoK
ab8ySPH8+1XGQgde2uHYeqrG1TS6bUombPi2TOeY+7LPIjrc7TpHJR7o4Eerr53Y
hnaGwFmzz5KTjYhkK3nIE2vqnJiK02vN8PPnCjDwUk0oV6Wd+4rnICgOH3ttjvpE
Bp1THlc5S3ZDcknVBrgHSLU1RvWOuP+odcllLm7OkX1xklq+q88p+GK9YtAaHmoq
RqBtJcnidO/A8vc7es2BqFDh803vTUpoPxcxscItI5WyUmYor7LCBH4GJNg59RTu
xtNyEOlK58bVG+D4XQ77fYlRw7OGtozjYrbV6IGlyj2h2BIJNn+9jUtrHuIyxxva
wZR+Dy37K+2dv+7bM8EsequFOI4QqehYdWxgE+eqvklCxL9tMOY9qMQXKVdBeiHe
3d5zFIE2d7LTUn9lWFLCf3RW9AHfrAwKZa7RLqmrLiSFzv2nyDOeOLZB1c5OLG99
zVK1U6QNb1LKvvKOKUYj30Mf/nftzNWKinO3YveHnfSus2jbCiu9tfi/cztvsfnu
TdWd4nTIbe/pmm56X7TqyrmdycVYX8CQJUMZ2guLm+Ek2JmwiroDviQ9OTvknOjy
okj8J5X0M/352XsCkVLsUkfNQybzcHEN+tM6s1mDaatk4cDSizcut/CPyoXZV3qT
/7xL/CQYY9D0vuz9Lpim0kgKEH0uA6dh7Z2Gplwe2EWyfFEyxU7WbZksHbHTJVG/
9nvICIsaGHDiD5ZwZgDaA8/5QC6OYGYZ8dcoaG1W6LOvQokASmwVWt5+cGICFeOO
lcJFyF7NEPBMPH8d6zOiV9gMpZcXveRj5wKDeDJ91VHFx766IxkkiHOP6GNd14vV
GcZ+Pn99vy2VahBFz8quttvDO96WxZNdUNb7A45h211bZVCgDMqyh5qusPhB6Ag6
ajyEec0O4dsIjAxEdluZ6uULfn9WRGlE+b58E7C540sZxKIVPAzookI0aINqY6Ih
gSLhwWVOoPKF/3jW6rywWGs+uUE+lFw/qAJ2keMTSKsvgVaso8IfZORaz+qm8hVb
fe4aUSVmHOgcOeH7b87HlhhKWF9XkY31btOeX9Ds+9/vfxbn0zJsloZieymFJJBN
lhVUQ7FExfgNmAwfXp7KSQwL1U3DnRaPpW/1MQvBYtUe2OYE2EqwARup4WD3RS8S
xDdsZY3E49HgZzdkCfw7VUeHj2dUia6zyUbnF0FKMjkDEDxAD0o+0NzgWpZSHorL
hQNnbQZ8gaAf+msgxXn93Yxkl3+NP64RSFZC+j6KHBqBJy3EjsKWfmhzlPc8sVuP
pZ/9TbQ4FCdmvZU3j7wWiB1/VtTm1yi7rnOxNMlfBtxTbDpnTDst/x2depZxNWFV
tYpCboyyPdFNGR84PA0pwq7JnKYr6WZsEbhJ9LFbsHk+6h/IWbOa6BRwiNyUv+F6
hOfj1rg90M14b15lDf6M9mF3PSudADr8VBFRhGM2x5R7gg/BoLtKAue5+Ws7djnS
f5H9j1YKlirwXdNP0ecG7O4AMcnQxG6PUOhS1gOIzqbv+gGHwVBJfHan6tJi/iCD
BPnut3PkVdhUTc4ConWxKQlLaAXwo6AKKy7XQdU0FNaJuo0c7mQIC/w3a82KZhzz
5qK9liTVfPJvyG5bxaFR1CFfvrEuxxO6SYolH73Gs9+3vF990esfqW3yswk4WPUc
CgyPzYdPru9NBoeVW4u6sN3U7Q37ftOEbvKjWXjnMu4r3ipAyqi2HohK9nsJzHEy
Xd0ILGFrhjo8FC/8hoqvSvdNq4/VGWox8N4wl3X70jD8++3MY+ZqJfaJ1eLv0FCD
UmM8I/lHCziwquocOWGy6wPrQVS6UZ63vZd0gjB6Yz5ZQd8Ydgm+o+SjzI8ht1Y9
uww59nukYABznmtcpzlx+lXKHE7CrbJXUi8RIdIVg8+K54MIe/P/7xQHI26PaSH8
ubidvbGNT+/sRtoDDK9kDYoJc7JyXxTZhxQ4vDAOxnH7r7DvyyQRDXaHNDK3ouT3
j4hfED4SNgH93posdGXb8MeNB2gMka8c6XqGOGzIXg1vFSBjU+Ptx2gvAfh6qjJZ
QnlWMhNd1w4q1ZS2TUA5/kMkUE+EX46PcU4YtoKY7P5HCCJGzPNEWLBZRxxG+mdn
XQ/MbTr7npZC2r6Lza9T0CJpJb6oaHmfY/dC2Nlw2Lt1j/oWT7jG/PhfzHGOSyvb
FzFwyxpJu9xk99NzR6Zv9NUUGnYwz6qHjtzsbbdXChzLqx3hitI4n6iSo1jvPaGr
PuILKZ4jVe/fJQtcy/ztJNtCgDcClOTvYFGqNfXu3VTqcbqRAZ8AiGVT+HF4OB/Z
LCp6AdV5RypZj4F6WaMkGJzkf/6x9t4zurK1tx9SKb1dlW7PVzw7AmEFFOdBSISq
7jmjw5ZOeOrw8gql7Ta6iwy4U/Eq1MaiIAr7qdUgZcvaUbVDiXCED/Fj97pBEpEW
GKiqNm+BFmwW46QspCyc/Jc6fgaYJGF04MCqkdyGZ3+fspEEAM7Ff4kWh/eqJZsI
hPK2kYqd/QHn79/FsxhPFg3aF2Pr9xry0oQrE6+6G9tCU2TUR7BhCGvxBr+wUVd0
0vxrmKoSsWFmsCIiXUxC9tuGklGWG0HUnRvrJKhyThOwk72AVl8rPGRQmiknQQBW
r6/NlDegHnr+hlHVT3HEIZEQPzp4lm6JHVhyLeV9GOijhwTco6gHMPwIrk6tZahR
ESk8Tsk9heug2XhN1wJBTUa605axYXEX6ZG+sJ9x8sV1okWU7sPWJKWlRtr66WsZ
MwYzngItZbNtIJtNUFmzXlyJmR05zdWgJ6pWgTK5ZSopC05WVKkKA3VSfP+vbUtw
1XOmdBqWYuZ+xKpLk6MrL1zAIjG5xkky2LkPSe/gHVjeQMhoScz9tDvO8HCJyG91
5cKfleMUvR0mjX28lrq5NPibWCTxN3b/MH3GhZ5YQF/o1akoGI5Jkre8RocRn1rf
MEJmR3YKNEgLGwKsKFNAMexifvZNC9YGeS8ah4UyfqrZJwaRRdbAzJHwrGFpd9oI
Q1RMFPXneytheLxGownpOg+GmStJpcpGyxEGSx25S1K4EbPVq+NdmphineyfAI4D
8br9PDvQ820TZTvKx+A7332Wj9pzILh5MndaP1tW0Rbu6ZbBFA18YxsKVBmV0W+4
nOIZAuXGv7k/sNnT9szYIwzW2BFLbaCnASzOU4KVZ46oYTcrfu/agbVlPnnQmXuO
YYAhzFm8yyiGUGQiOZFd2VPFbZfYwAO1+htorOTc5hbtikXfHFkbHQiSr+AOs/y9
JarzOmh04f69TVWbyMzea5uHNiBVfL3kW8PQh+I66SxqrR+NgP/QGSW10i+8w4Ne
KXMhuDhZxz+45INxgwjiPjlFLbD5E4kTVR20KfiZRudf9l5cF3P/MNtfXpv5jtrD
oekp83vG1ndifiuSAyLH5HUNDvtPyPoAwkSJnNGoIRdH/PEZwNy24MBtwz2EpduF
qKadOFjH2tJ4A/PdJD2dcVBWBzNQy5N8N59CdTJhv9gMAp7KxBj+EpROe3o5bH+N
VZG4qXkrATKdD9QVEQbrurkSJ4JfO2RruEINNyiOZdX9h04ZRAm/aidlIHGdBQJ5
CNG6AYc7tOd5tZi6abjRuWQFWPZGVCA/XUNgN/M33ub6NOlu0YYP2lJLlg1eYkaf
UVWR0r5ut57LkFVlTgOvUs0gm8IVMHO6c9UMo9jrjMajMK/CRgETtORt3jbhyJu2
0ko6Ftji+WML0jTcc2O7QLXvyjgtY9ga8tZCr4LA4wvbVwJYo/zzJe+tzqfBoWiw
adB7GvxSpiE1mnZ/eZyvFLd5PCbaKDmp2BjxpVgpbi3u2VnsqoGsEV3xRd5IDG2V
sezk4Xh8fwCrsM6pJgQ2p2+uJRczE6zZELj7uVwy7afCfpeUqAlA93BkdYn6Rz7O
WJl2pGR/lW5t2YvLOXtCCOIjS8rvxMP4NbzvnwbsOjQwnlUukx57h7Xen9pYck+j
ouv0XONq+1F+hfqZKZQplMNMto51+ujtwm908WOPnAcGkVvQ15WPbrL76pbkhTJ9
fPqonct9KfsnLVvXZkAFh8tKV0W9h7RmCoqipX/tuImXqQ5FeSz3M6A2RaF7lSTD
6pUDK/BQlbap0XQDz8KdX+YfPRYrS1jPyjfJsYhDR9sCq6uoUuiRGv0+88/q3kgE
KWuXIyQqKonFnQMikluVIw3ATEl7FBSx48jZmxCvSZ8Uky0uHDMgIB8O8Q8+iMIS
xdi2n/GRJUKIxww6siynvxFzIBfbYYTxsFrLU+faGQfPUt7Nb0ihWr/4zDkaJ0VQ
NjZEL95BYhj+4hnJW92/sOGToGEaL4KFefLW+qzvDXJejQd/DVS1qOy1dHizjrwC
UOjG/YIokc+uSr2bfocwd8C0xuEIEUhK8qN+eId6z6+I6KB0jRnWx0OBAz5V6+Ax
RXsFH9Ayf++kMW4fQYKM2/mpTT2b7M7BMNirDwbqQzi5wa6DeNzOFJ90fJi8W1rM
Gl6E4GwN9YbA/ufd80CilW3cHluCNVWgUjHJgoK3zFmADcbQtj997bECa6UgXEsr
8XfLQms0Rh59yU1sR5v0XmPQXufERGgS4sR5BNSGzTopc6F+TwegkXRyB+EXTbh7
mfkXbIWzgBjdNx7ihCkMmkfENn2arh2VfelK7ve4nSJAm5j5ECWNlWyXE4Hvz8dN
4XQChzIqpPut2F5Y9SmVr102S6k6rLbtMYstvVmdcl/iQ9vdEkrbNMPSQBbD2zbq
y95mJOf4LVaKeeUJ7PqD2PT0shv3rCS31fattP2ltISoaCmMUp1O/cIutW6aW8c5
7ZPYFUOFHn2wHuulppKGRVNbD9qT8r881bbaLgX37OEcwDGxgVdAIoN1CXdFbqoZ
/8uYG0215giMrNKUji9EQD7iYX2CO+xjZBi6B+ism87qQObmJojmtG8Qv3yCgo3J
qGFof6KyJpMxO8ibBznfHlKiRBk2VTcJcojgOwazte6w3A/U8aUN+I1ZV/NuMrca
aXNUA88aYMIBUvra3OED+y95iEvatnq1d1SpVvZaJnOFDBqKR7EQKEqlYVTAnYf9
XTt0Z0DTIPw2+gPSWb6qO4H9f5SHpnGIl4+XXA2Yu/WhRmII5bXMsBAVpqTfbyAo
Ri1zyZ4X7y55d5IZ6MZXjjHMLbH6NBBd7o+qefSVBYFCJ1IKK7XRF3Tf/ZYffiyV
aimdnHTYRFNRD2M1BdwylFBoZvrwDKS7l4fglGmnohDBj3OkTZ+PUv2b2m46WMDj
3nYndw6CudRjZhE9w/ZfYz7cZ8BODNN/Wp205bRKgRqZSfbJQJE5pc9L+se7y8/F
GgF+JXic6pidnf/G6ihAex1IORr1lvV7Y6tlI935b5nMxjlh4wTs1cxaBkl/9Mq8
sG0a7BqCRY9UgI7xD1FHiWg1W7qOMxbNjSHANARW3Ao71tFo2QRzvnOiFFCiGXM4
/UX+55O4TI9smT044MOc+IIjSWBZxfa7YXOv7xrmisPzz2XYqmBzDtAhR7rezdLB
eY8ESMH3x3UOLsY/GFtpA1Q+rRoCQp11Qxp6j6B2/auECdm7wXi4pncrZW9Up4P/
WJisyW6HbhD2JE8qowYKzZns58Mj1s3PsjAQMo37xor6w3Mw14t4DAOhzd1HDQtz
8sh5vSRm96cxSwzYMjOtUQDscdT1LV5e1l7Sr9w4uOYMmBpf0bOy8cPSuLm0r9aE
b52nYTbBEMJuhKuXdzbU91/M7JDAiqahHZDM3XlJNx/mOuUhITNaxGL6jCDxFHNy
Zwrw2+G5+0HTHpUYcnCG+DK6xZExJY/kWYnRgQVPQKH1mrksfiHaO8uwrTo8IqWc
YnLIB0I658oRkf0S0Uyesa6LGfn4xFU5pKiMWEJ3FKFblVXQEdNHF0cKnl3Tu9BA
ldYjI3ycVLwON7eAhBn98lmmg0OhLNKzGF4IqYkskucQoDJhTkg/5S/nlNvVNz5B
2miL3uvHLz/E+Z4db/vn7IKSsjk9wOMNkxkAMlisrf3o6G0G/WZbLgJRf/A5MhSw
jyfnEtuK+yoT+6hhsqX7yosj51+xPyzHKDSxBFA4lMnYiBNRpWlsTFXtiW2Vmpso
ED3VppgjUTGTeIIOvDXMQbg9Ml3E/b3NcjD5sLTPDRf0b4mpgYQBqCuCfdBqHnrC
4sCvTvJixqBMul7D/b/6VcS9gWof0SSXxDHp9XAzmKW/7xY/iqgs0+p4E2yTNBGW
634vOd94ZHCL2JpRhJwB/yVf4gvlFRKDHxW7AF7VzQIteKdtYZ6iTx4Z14rvj9IQ
3uUFrgmsZ8X9l0wC7ycGHSHhEIk7Lxr1J/AbVA0UQsy3KeI3lMS6xTjahxuM0RHu
s+zbctG3gDmXo8yEJF/39WG+3iH1T8I1uLEju7x0/tZiqjRFLjyK3n2/fMoaoVil
vmF367+i6/ai+kaeTPlZJTIE7zwQ5Loo4Cw9F2Plm6LQaVSmAYuppikQTYFlfCqa
97MrZqAdUIPzNfCSh6lEQDA3Mof4HENzNbF2evzXV+G3kag+zgvC/0dUnhfXt/TX
8H39x/D/x+XFDzcXiVcG3J4WU0t/fOdRXzzGDVFGy3W23gJkgVoRZoWiApj+xYxK
FpbtaJBDVnZjC4CEcG39F1K+a8oBjC+6ndLQsYH0vmb2E8bOa1ihTIciBpUu1f9w
AAKEGxQICU03wxhTbGktUgbrJmw8DMVAWBEBQTNBMmJD+X4BQ/WQUqzowL4mz8a0
pgKUxo+49U03OoLx2NgirhX2X6FrBv0F5FoBlr9WD0F5nZMZqX7NqK9x/RT6zHbS
KXh8sI6rLpU8b8smEJBRIgiiYHIft/TukXlBvI94yijpQ7vRwvx3mgqKoX6gG2xW
U9dd+FUOnldsvltMKnnI7t4CdRJ7G+5v2LGoy6VvebOwl38VUSpmSVl54FA6IyW1
YLuWdPvKYcPGNiJF+B/gE0hL1SMtPOVRRP/XEvqbKpybdetwrek5X63od36tZVtp
u41l+JYIIateygx2qOWUsWRIeLnE0VzmsVp28FllldC9Bj8naybK+QOqBpblvXN0
xjWewSipozo4Pf5D+LqwXAN5gpmXgC+cDq54wl/HfBFykUYEMDKg4lx8QY1ITO3c
PAhbioGCWRwfmun2rCdzP7lRnvzI3SsXUondGQ9UGAFDtVjPoMA8R3+sApy0Urji
9SBL5yvYq88yTjPVuds1SodQOcxRtZOaUxKCeaEICIsAaf8gnzBpCFpf0yWiZrSR
5ZsTH8ePu3Tyuoix3tBRHmO0mF30KUBJNulzyIRr4bpaBmsCEU2z0DGkFHOCjTZL
WvUC6W7bnYLKU6/7QoSXOiF+wz8Gp+PcaMIJkGNr2i7bsJqnUH4975WvefGlUfMu
FumSBAj1P3h8TvsMgMZ5HfRaUphmUBwO/SahA9knGVdi9edwKJa78Oj96e8KSs2O
wUzd/F7Q2FzHisshkIMN28pHHvq/O7bCUveR/T4H/n0Eg2CmCIYMbvfhXYSPH12A
YBP8FTFp1xUW64VKsIVUQn2KpAOUiHSTuweEBCsRTvkiVUJhfZ3w2NN9PpKWsRtR
4f+JGSYkgjvngJs7QISI+LEPQZ6ChW5H4ggO05kFgy+TzFl5r/XdVxcAzCfkNCIF
zEWbUsFEtLZW6py9fceUZ4ttZG8+pOozFFF/XRJYDxLQlTg8c6oBY6QFr6n6VwaS
Wj6KZgDZcR9xLLnSTypMQQ3EetXuOhSJda5UheR2DwYRlHjM3kYlmVo60hOviBKT
xxWSMLophdc/Fok1j0s8tPvVMU46h7hO7tNcsZmD0HDIio/D6EWLfHCnslG/n4jY
b0xRDnc2OgEVF3JuYDiT3JHhIQUxC/6jVhnPy2WbVMe1KbwCDafOIOZgXUvfCDtV
fmnVXRSSGvkXve8fmUAnVV59SzsOaOzaG5bP/kVpHVI1i1yFrUoI50Fz71y4qDGk
7mMiiVZDybo2/JHZ7HLuKBpqweQT4rHKf9Zr6vsCDRTQPt3I4A2IpnH1vGNh/8Yx
amlLvH09ix+MWdueHK+RmelJducVTBx/ay4h8TERZaC/jbutvN6LKk0ZG/1bg/aE
ZW9HqrrCHnq5s5A/JeJ5rCWQovfOIqpyVGekQWEo2Y310OEmk5x766qfgb+hFMoa
Q9SjifL81cvWoLp5VvdWPvWolZ0Ld6SvEzndpdPrFq8/dcWW4HMIx/P3amNubdTh
ksBMUcMV+C0eTd4u1r9tAhMzNVieGjV/od+kYDesmu6zE34hYEJ/eGZx8y/NNE84
22xH/SapRCYrumAT/pwXI3D1vLB7lXX9Vl0a/9Zi+3ElqobOCpgPrKlkg3+vO6sl
sLTFVwSjlyobGxaoQZJV3QSy/BUI/VDo/2AJ/GbTJOKglpRqMDoQE5BbJvbPBZP+
1rfPmOFSm4p2q6v5tRdJWnxAumnTQMFxNiQrtcrmP7ZE/vblrPivoDdQC/GFQCdf
pIMr0KyzxMZtVW6OxBQlr5FiRVQ0jsPzYylKwpMQMWHsNPobk/uD+nK3OCDTU9w5
ydgfCOizTWTl+IaCoI+dMIjkETlQgZnBZFu4sscGSw9ZCaRNAXM9wx9eNbRPJdlG
u6Y+AaIKMxWoHChQU5jp1EVuhXo7KmH0SVsML2jlqs/MREq7K+fdgGWJj7zhLonT
YRDNIJZs0w76dF5SuQPWoTDv5jFyeeQNBRg8wJzrS8ECyBeWp+c5mKjkKfNvO8Z4
GDdaH64zFsaOhtwtQ+KyeOVlzE9WYem/4yJEv9OTJcRThYrHQuC23WoKvDlXXzO4
leNUIPkq+qQL/Cub+jB+XS2FLD49n0b6KrBmcfjglz/Gvw9X4WfORsEA09f1h+v/
VoBCBk+qGwlx/pvqBTE1MeFuAoyViaCIsq28c9BGa6XvSt9XIqOjSBkEa3SrKO/t
ph5cPhTNqZbb2vVnBgsx+dUAh6IwJF8aliO72q0isaKR9fvzk5zgveQZacL1Lghq
upPTU2k2gsiLIf2/Ro14pdzJzz8Ddb81aEhWV4BGltJvNF+uBJTJcsbAlhyxturO
iq9tVm4JvIcGlRpyi4EHPFsabMe2xFbq/T3TR2/6x15wPgbltYHuO6+tQpZF6IpG
A8grAkbLn9ETfmlNz6/5qXy24gXRJ7f1RqdwUCyL9LWFyAvtt3vTzpwM5Hfo2UZ9
N5nxzS8h1jV6CUSxOwROu/cUz+g2pk7XIVhyJgyNNq5UswsrAVDDDJTaK4hea0g6
BT4onHuwNnvCr8KmCY50eyFZ+CyuDtJmyGBDTQ6gRZS9jTSvRbmGNturRDRsAn/Z
N65J76YgjGVn2/9meuMhxknMpeytuF8iULMUEX5xr9CucKeRSPxBaw9BysmtBzKn
2oTcrCQGkDbCiNF+vwkkF5UeRECmiO2g/gNKG/QLeDcFYVS1MExtVRiAO0O2kjdX
tQxv+XIUtcCtWBmp6/s2r32J1gOGz2PYHCB8ncY5n7sBYOmhTxTABrxAAXy84SS0
LM8gZN0NLSYRwVKh7Mrbrh3x3veGUhvtzahbspx4CN3Zwwd5YoWRqcfhdpmYw7MI
Y9vE7cKTARKJJ8QyBT8KsqqRvy9bPShod272lMJytU+RehtG+E7MhZepuDECidZa
2kasc3YL3O484H6X3i0PvjhRvzWV6zAxTc+6lmnVnUGxATziI0abqIcudWIXKp1t
rEbgT50q/0II6Jhh2PX7A2Hzi563hnKlvezmwBawJIyouoEmHHsGxkg+haMqsNyz
aF0T4SoqihnrRVZlUidgfsaH3DeBwnO4FGxYRDr8ON6DI+FaSVJbyhTpq6GAt2ac
NGV4lAz37NslabUkZhHoLkzZ+8sU2ddMcsfchK0U0DU4vg0jfke6q+J6GShvc/0y
+iBHq6L0RAgugjNJTyFSM+E4hRpXF5CQTqXpDiY6cKSzmgv7J1t6yJKTdNo6TUuc
keoIJ4PUAjYHD2TOQoeClZb95IGAdBl76HBJh3Gnsibv7itUd7zZZeDyJHs8UFZU
Kj710yYA+v3c+CNUC0OqHQ49obkOGVtHdrUy0o+LcG33Pnckn7BnD8ZMsucWyvnO
0RtrSDn7xmBCcTyxvZg9dFmb55v3QAsyO8N83EVgsV6u+T2waMMoYtyigl3RXZBF
Jm/LuJyPzxjyqtkoJaSHx4y/nMqnm6Wc8UPoMat0lrYtrMvYw8SHvmlcRyoCc/7E
2AGLJn6wJqOTVv7AGsOMZUXH4+YArgTdiHUEt8yOV/t7tMEhT+ojdu2Ij5ds/whZ
FdHE7lFZj6Gz1gJ6xcT0E4WzROGk2IHg8lc+Sl5XeouW4NWpdU1k44iiPeMYi9w8
JEYHACetIbemg8eoXEmNEJqFqmoaKhzG4knXGAzOwFS2i3F/QjwamnYK7qRAuJEL
hyWlGur2Kkw3e8B7Vl6S1stTc4HgOG4cMk9VU7m7BgvqxghEENQ33NYZoDwE2NPR
a1RLKSynO9u5Pn1W6kFEsIcsNaitT5MEZuXlZpPz48ET8BshO9kthHCEmmpRUMEH
mO0kZrIKCRtwpJMwco/y6fED4Q/NWwRrk+fpQyw9Ds+QClWlnE4ggxecCQTkCPoZ
WUo+ngH5ZWa6uQRNACvgTeEM2g0BC9UDFm3rBUThy89k7FXC5MnvW7AcMAjXtf3g
sxvphQjtRzELfqr6XdDY+ILz8rSQCywGxf7eOLsU1W27u+5XfLzYRkDmdJgLYws6
3IVYqEHLXOoCS7lt3V1jt6Mv252rAiD06vtX7jzDcLCDtIBLc/Cqo6aIMSeuJysx
GRa/621TXQsQyx1QAA2t4PvklX/97DtrO7tcugyBhU8i1PukGpDbt5/BamrLF+Nc
j5/IedKxNPgwx4v/0B63hVmj8mRhRk9wELhAQ2gFH63UpOaoRn2jfcXTSYgVnnaO
qYPnqj+HOuoZyNQUYO082/nqG+iuYNxC1tDLHUYvoJar9dm+MnKF+qub48dGpTrf
aa7fTnZgQJBHFBP8Fl2jjiDYMnJvH6CKuTOGmNVT1pvwD2kDxkl/Ox70FG6Y+Q14
Qg8pQdYgFHKMSm9Q4kYuqacU+1GgVN2p6wCzkGIH/BNHJWQssPSRQGdv5tYrmMUM
FPGn9CjhBNcTMt3TNMtlI1J6DKz8A0DRf7kJolAfUUjkTKOupEzd0I4x0BpVmxY6
6vFMKO+6a0Mt+9V+Ia12yqMh8EGWkxuLe+wJRZQVscV+LO/TDi+Ds3LQUrA/b1wh
Hg9F6pN0OU9mI3rHcKHRGtNDTKRdxbE0zLQvIIYoLZQuchT+kwugHixbSNzfg+lU
byiEo4gs5xGSHtxzwhQn9dmye2GGJLTA3RRYz8YBArR2XKnrhlalBwHwhApVlG9x
lLHF7S3PNRAY61QoaH+2FAOZdI7YaumyJoOEqtg3igW5WqtGNtoGrQc//LisCvj2
Bid2eGpv2jdJIBgdXgM+ltISFXDOrT0t3IV3E0jSIyM0tZ82hkC4Y0i8WRqH0IaF
Pj0SQB2iCnsKSG/Rs+pmH1QqMUOxbmg3qMU2ImaqWYME2e/d8x4652uk0MxJ/fi9
Oejpb6bYJQqH+YrrI+qx53c+oy9l2qTtKYVWqZ2q+RNl8UBxf6x4qUrH3LXqP86j
hguRE6AF5JvNNL/egqpzoFDjazOwBbDF75JIiHoIOJRNO6teY98SgnvLuIP+zemL
LwXxWWfFRuZum9IJXH9i2Pc7sZ/WVJCqA3pzsRXBctuJ2B54Ak2Q0RmjTEksscVU
EteYvaTITPtfSPpU8mc44zhKDBqxGkrgzowzAkZ5pZlo0uFm8x8FNjvgib0glvyL
a9Zy7EBLJvqSbpH6d8fnSosAdcw3gPcrpXfUcUsagwwHwjvqADvcBmTaLipbd8BP
p0B5xq5hkkpenemOFnznQfLXCNcwUOyyGPQ8D3zFNBkcmMTBBlQ6W+HGUlAR/TG7
jQcVzpCTnm+ouBEjzB6u5bf5+iMEjKnJYEl1d1Iz0xvmFD2PAIJ17qds/xSt1yj0
k3J9t5YPM0HpnGoVcko6cyNTaEjmIB8X1uNn5jDYtN+mR31kzI0Tz83WuwAjrfLE
5YWAzMKcPXQx5bxCSCV3akkJP1kFpu7+erezcd/mkoHW8d1lAZS2jYUAf4WFmF1e
Ul0JlZyFAQHptf5PSGUii0MOoE7WoXOd6NW6m41E1T1uo3zAz1zc1H8vrvbDUzgz
T4X2BGSFTRAcVLbEkJyVnTeGbSwTRrCQPEdevrwghSHeIvCODMKMarp7N0H1px19
ClYebP3OMZj0BMvIlrK1X2FY4feDZYQynNiXJVKaLmJ1iBzMN/CBSv6UGucZqZ0V
dZFtFaPzeWS+Si482u7pxyj9nLlJByyxHvgX6sPDlK/3OszpKX1EtK1W6rGeN6WN
zBzQSADOBcTglCUHsHILWkGcXPmFz58sk3ntPDUGf7S/PIrLRR6VbrvhdFBAhPMR
zSEj1x/yfyMjhOKZ0Jm4yT/EibahizvtbXQpEawm1dmCcqlvHoOEUEQwE7tW2Cqz
5+p5UMNRS1INyQ2w4QaBGpzRhUQjJJr8nhJICjvanCId9s0jPC0lIKAbwiG2aeA/
xzuDsy2lNqLz/qNBweyBFPvkzBUIkrccFSC82Wg9Otzg0ImD5e7jRB2ZWR1LnIAT
6/3jOUzo6SIp9ZsM6oZHtLDtrKgsoUD608FqwowK4g5TTLbHtIiHWGKGRYhFB70i
3fZG3XMCc4RjF+89uL/x/nYvKF7uQKlus8TwVrlcNYJG223SkIOYZoNJv+AF7cpM
uBdNwf16SA1BoBj0wkc2hQospnR1nu/l6Ep3QS6Gl8xKtYHBMo1ZtPpP3YmEFScC
MwC/cgFGwHesAthstR9UuM/yidLEFgUkziSKY2646pB5aHMpY0VgCPf+6J/a+Dqo
4prRSrAOPTlU9y00MGgMcTFdEjiHhoZ09QeYdoHj6el/Pez2l7+8uMTffcq5t/mP
1rY6MnbCDRo5UGUD0+MWp1DwXAPqnGgQaIRlXueR6QpqQ7r8zWy+Bqt1yKLDnQnQ
eBeGYzrMuTcmezc4qPzn4y1EixWu29vrvvsBiSwobIYoKxp2JkttdS1yN8dGzHjc
NT+SGPi72o2xM9bEhYFG7c2PdkperexLsdbF7ZMXKx0SqMD+v3m+9qLbjohjS4u2
d/SjsWFZ75SuDOXxtd4oA6NdAKykX8pGi/scU2LveZkXDoXVGpP+V2PrZqpIMpsR
5p5B0bopFPW/V8PlOSlZS72zkAW7SlcTOOkrdCE52lRPAB1OXswc1BfI9dNqDyJJ
zMAf6YqXmsUvrOHI1lMIwaNkSNfM4pHwsYfnx8hBp+RSVHXeKRikWR4i124JCcYe
mmfk4wcMhrNGUTWS82T1BZ2a1V4yZBnLEZB05/0gRy19NURPiYQrEJh3VQr1Gbtg
8Sbr7W9wzMCxx893vzciDpgWMnDwHzpbwExJEroqUDJIEiA9kxnVdeVHaV+B+/ed
hGXAakLGB5lRpTb0ueCovvF8UuoGUcUHeRvT0H1kbzTqj6Q8a4v9dOh/aQnUVrbH
uHuzRzpn/h5L3obK1ZYII8yhG5+0ba9ZpSyWwbyidiAE18EM0kFQvBQqGnSWwUlc
aqTkvz65mAPQu1iojaGPQLmS/RVmHG1unkeYccOhvp8ZhF4G4C1q2QX2nHzuLhAf
HdxXX05kORYq8c3w92N5cJyWQgE24gKF3P3FZKtMpcmGXGgZyYVbC7eIvrG77Kal
AxsZ54DDUj6FEzliaSjo9vkSWzQQxQ2YP0ReLjc/oUXP5D8AMZfV6rsCB24GP0Sg
rTPS2CmL0UGrIzKnXU5hZhgGwpRigDjx/gW7CpA22kICYexG7/1F6c88qQzQjOes
OCh9/JGzV0LIXG2vhPRXW0P2+cNEwIlFcKGZXQbFwNSs9krrb1qa86M2tq4Yy+To
sGUiikL7DCmdz4uAgUkcU23Q8P5eV0J4EtImiZ+OtuD7F5IkxigvEAqDaq0ryxV3
wslGohSjarrT0zZbqJ3irtnXRvZ1vFfTbLP/pt039LLKMq11+waXZfUylrUSpOFr
aIhsEYBY51+FMM1SIX0HlBl4zfHrCu6DfYzTPYT1FdYjMru7o/CF31o09KX5J2Tf
6OV1JyfbfRxU4WheXjqpXmDRTz34xcRAGN8fem/wbeE/+rjjX7zKnA2Vf2iLFRft
Er7gk0X4ZgJ8eWkDNrHESNjqjDaaJVx9HPQWpOE+HdgoQT7aBX18wyPSh5jwPvRk
jH6cPHypo/TKDiRVN3wrnhoGtVTLQJx1QFH+t8lR6eUOh9lpxC5e12vHhZ1mJ0Dg
xZ0vnUsOVBW0GtJflI51Jw01Pmi4cx+OaX3+7NMldhCPtOfrwO+sRi6NNXOT6+gI
hR92vmwg8MFuXVIHQJuhXRP2Lv2i1lh38vUAhqrgCJdq18iRz+jCFS0BzlqSeCVJ
UYKoaNbbGhNQmoOlRUW1v+G7thcKwIRQHhVMZ6jcxHWfN8fPtpyC38QDwCW3XgHj
W23rf16ReBFe+aexI6LEKO0+L5VfFrgal0ArKkFXCjZovX/FCJ0VpmWICFjZ7bSL
lf+eJ5FO2qLn275c/uHFr53BlkKIdnh1eCH7k5drJQkmZ/Q7p/H74xtRuixXYc0B
dBMokQi4RM1nrb3KYzl8omnpX+2q8uaZxsRagMaiVSC4AJ8pLvTFc6d2cefrTz/g
C8Zr8p4k0vKkQfnqZE414E1nBKJRN4on8X0fivnBmQXnvUsk5k8OCIHig9UQcizc
8C2Us/HXtWVFVo/QEpJmZz8uvIaNOKW55FHKrg9JC4fERGRAp0c1n98JkeyLvdr4
bzFSq5jT7c0PUe8X2ML6t9d0ycvKkfaOAcu8sH/OegvOyqleVxjIH8+Vuy/hlB7g
+R19rZVZ0xzASHZXsa9X4Dew9ALXSzp2H/Qd/FHUd3cYUr8DYzdwiy9xYyZKFN2z
LfePoZz8Eik36qoKE9b22C7Rda6+x25IYJDN08bZNL0IV2UdlvH79wYrIW0wrWwP
zFM/dsOXznNJNLxwbLnftOBCo+HX6U8+2JTKKd/Sc03wcbDBg98I+YmTtuVIcitr
wuapGKhj/Ez3bHLfVMHa7tP1IJ/zBOh4gksRUt84dlAzqJ55GldqBJ5eR+SP/S9o
jGQFN02RiickES5HQW7+5X8wG49srTzZasRzEPKY93toZ1MoqGq74b9pkXRZfS4N
Sw02M7N6Nx6QNvk79vn9rhfJEs05dho0JfqmYjZ6IJzXI5gfWKD440JyHYWBbStO
OXlgJzZFxGTDOMKQAEMxqkfiVdwJlAy0TXz1yMq1IPM6kurid0gWzK+Ga3SfiL8E
qi4WJbdAyK9L1UC887N2mwH78dYT1d4L3hjD8NNZBVK9We3p8TNYNNZmwJkYKhnq
HWXioqQUdGawxLZEcxAEpXO2oO5WcxA5jXPDQapvN1VUzv5x4UEbjRFGcxZEFrPl
ftSYbE9utQPW5iu0mngGBPI1i7JbXC7dr7yXIROqVy+deLgFp1zOaUEpoHtyfojt
3PMzHYple12uqENTEkRal6fxF2eAKJOYp5NFGKCFdmifkrX2kIl1Ym1mvGK2y0TO
IQb0b5kDF7Kh4iho4rPb9wD1QNATduxOMhywctbKDDwiL83P569EYkzxnZ0eh78I
u9l3ksbMm9SBreH2rPlfTZOFpUD09x5tBVK8PRuh4VdkyuWOU3SJzb/17e3cE8Fk
32ISYwUsEfRN7wyoIzjaXyLmnWbOOo1G7SrTSgDi7ZHxAMGX3UTQYQAWiyzsoHWa
BeK14KatReSuyBCGFQw388QCkLL1k1neEZynzjGiK8m8AsZvnEJNksKH9UubLYW0
sYaTTtsJOWo8eHN4aGzA1vPp9iAlW2a3GgXZunNPcw0NWQ6Zo/ToWcRijoqupSfi
gWLxr9LaYrDo6Csp4B/yO3wl9OgBatsgE8VxaINOEPx68DoiP+cjpW6p6p/J2Vw/
bPrv8qbxfY+Xhdg8ECxuQB6X2+uGNMGakfJ7aZlicIHrPXACEudwmjajtG+hrRPE
YS2I1U7ycyGnL8qelNnwR8Pifwhg0oYIv6RDZp1CNCJoLVjTna+J98QR6nqSb/WG
zFV2pCQJToRuxAAYh0DscfY0dJTrA6wabTIwKrB3BsLGIyAkZj1mNQRz8D5E9AER
pb+JOGxP+BgGwh8IctzWac9B//APfmUGjHRIoWNSocqrnRGnI+Phgpf/02ohQO0T
Ke5zxSOB3Oi1orud3CJRuJwj2tNyekZmMpXfoefxb1C5eXYjHIReUX0IsVPSZoXL
prg7Pi+hbPSPkSqM2SLqW+Z334EoDVGK2o4GgTP+kSMxOFo3ntktH/+ZVxEwoyYx
lJVoFvOAFDwL1lNubv9szjvWY7tRql5oKjYZsL4VpKB4wsDMQoy0/1nc+5VZhgco
492h9+8NUMcK7xVxDPHF1cVckT24w7kZIbu7xDkX8a8YgwQNXhij5ULUmGCRDoXX
6nmdElgflwb+nxriTeORlwrP0DvxoJ8tzWJ+SO+UsQc1ovuJ7tM7U0AnNkL/JJq+
yM+lw61oQBdcSUoxQZJYeSp2SqkD6o/P67QODkfatX7WYEB80XBThsRdNXwgTDNP
fBdhCUldHPJz9Hu04+bni1mS704cBOPqyO6BhVvsrIhuogP9z02LFJjcnescdHLP
hJGlHqwiyUTdfSm8LbzQvDR1H7ntAkeYq69R8g57pcknoY6Z8RXiraa7uWL6k9NY
zG7i5d3XzPet8LI+dgWCMwz5X94a5gAc2BkxwiGqUsDx/zhMqW/1ELoDYKaV2xpb
mgkT2JrIHiTL/lMEIlDoeVtdA1tIjlGRZxvU0G9x9unfSHMYN4Qj/giWYYfpwP/+
Jl+Zj8aix0Rsna+GulaUvnHFKIHEY7N9mpoyOdWE6AW1d2LDsinDllOadYPhEyiZ
b9hinfyg6vkgXJkfQRS2HRiB9hhvaLQN82fkdVOVTMsfNpSMkeyQ7if5p+RHnsXi
Pbxfj9R/U4bVz9nvOJNcyCwPiggH/FLCL9OTOGtH/udGS5GR9dp+zxeJqc/MHMEW
1rW7/WLBATk9HygLoEkUqEv7ecHK6V5sdbv3iUQf5NoARxETHS8gE0aoV5SvzwpH
R5AYbtBNfrorvAOQmNlOZxZ4laVodrb/oBnytFKsmuY4Q+7+T4qFo3Y0Hk3WJk3N
fmg5plsIuyRlV+cv3V9jr4pMwcq6LeE65K2o8K1ItBMvnGC7QVSFwQcV7YuC06Tj
sVKUpPv4s1tZrxJA26GxTbkpHA+oI+ARo53CYPdN2s2tpOLEm+F36rgYEaTU9T3I
YCeLREKrALtYgdj+bwkpe5DMJ56VxDX7YMWDSOVaXNOl5b9+lIsmlehNx5itnTer
AYG9UQlnxlgmNnJY/zKHfCKwcFglx/mfSCxhHbEI+2XYYBbHOAH+8TE6b5i5U0L/
AV2Eo0JuGpDpUqxhNOjWYtmJXnJl+xGdLCpnXe9TkjgR9zrzM5JDX9+S4oTzzmLi
BJSV3d53ikHQjDl7gV5fYM/vtQD3w4DbNyA6HPvbvbzqNAejcA6PGLSLrmQafLFM
OJpfIrCp02RuxX66Dk2e5Ey+Tl895PE+d1XQoq+Z1xXPmdgPQm6Ux/kXdB0JFRUU
mBwxcAiiI+eMBxtbJ9YkT7QnKk4GmZa3oZs2XDWz0AMQb4yDKYsxCP6PrLWcm5QL
WaysafIl+joADrwC3yHHj+0gQb/CI7HFIn9EjwTSNVJRfKGkiAjfOI0lKL438tA6
KLt6KKB+hPB55WwJhm1dgWrKFEgLiKWJYtXig7qh93oPv9WhqQruQDtWj9+aTjP2
X3k5scbpTB1U1aVR5KFDdKRykBy5jMH2irh/oEHiCybEi0CC0Ascf1nmjWuPM1LK
rdF36m1nHdIZzf5A/Pn4OjwHI9B8Kh6WjRCwn2Cnzk3/LduMGB4X3crebnLjRrcV
5Tzvy4PRZEjldFTucw+bBlMM4PHMbIC80ouunwWmwkAqdwEbw0OQNqZy0mYiGE0+
Yxz7TEFuANCo2XDJ3IXP2OHE6vHuDvcN2UzMIsSvcrmtLigHaq9H6lh//UcJrh19
jKpXZLmieGNK9q72mWpn4efFrn14PxS5H+ddPRrZG8ravsa9n8oPJR/PJ5gPYWyT
95+nbF6v4RAFFYuAMAsoCszymJx0Zj4dy4faqHL4qKq/t85rmWOdleqmNEnKUldY
x1VvjgZXdIoAY7agjvwZKZcmubqrQaBfxmO82Ilu/LQVA1CehdUUy+fLiy3HfXXw
AdF2am5uB9lojpYlsJ18Zb+T0JwEcYGeQjhs+i4BXplGFVkHfcrn4rWBN6MZV2pG
SCtGSY25cx4k8UJtqAOGC58bLyFlo+R2JfL94jxqZ0ARRpbUiKiYJ9dPXOGsHPwO
gyEA5aD3qcJ3FVeUN+Qw4DEzsqr1AuQ0HzNQVLVG860dBgTJfHwmvY1rnjrqmgCk
E33sNps+CukSGafov0mE5OZ0g8h6cwlW1vIjIM4eO6rshvDkonlz3Y+S131I/fcH
x0+HU643+tODK14LA+MWjjDVJqtqZQW/7hig33IFhcQhcomOT6IKiuuD7fdddqJ8
LB5cYWT0sPZFKK6vHdmoz9y3Kfn+WMirGdROp6WlV0q0h0+BVGa9GieUwjY72g6m
ZeGEmEUrMPH9q7O3HE0uQ2KTku0oo6pxbVvGwKh1K/fhnvcPv1Ndoz/SfrBd1DfC
vu5ES8S0xZ06BmKjSfSZ3M+i4Jv/qupZn2fQat1OvAKXxb+886lsgjFkoSsvgIH4
vKiWPGNyiK6UIUMTDfVyZ2T6oJJdZcU2HrIcf1jXeWq1k89VXkPj1mbnW6amebEn
qCj1cdb+k0HaMXAw4+hByuLTkG4KibyEuY0ZI4N1rVpxqIyw0Ds4wXAemf++cdx3
7jtY5UflE+bJBm5LMRorpdbK3bpNG82NPBoAhBVafpvNjG3jVDUaU+FYGziqbFV4
RuD2fTBANsN1jvv8a7YQ+pwiaTE4Eb4wYhcGAI2XwvdFbke27LhrTRhqVuizJE1b
DKuMQPduhD4aB7vj5hf8DXI3U5+peXW1GFh4RUU978Dpc+0RiGsnG50JLgkIWB7x
xEwREf+Y2I7WH4rwunL9tsCGheo71oRFc2j5mIXfeaWsUkMWYqgErouo6Uz5qRSu
PkPStqehxPYNGMai3KnxZzaNwyIJfyL42SJMEyrCYVqThJBw5OglMLtJDoQs54Dk
FBEJe87xuFc7swCHC2ZVu3RuWKmJ7Cp2Kg0FkecKshtQl0+K/W5Pt/+mjZ5Dx65o
7fcFNdLXe1Y35wFDi9/U3dhYnMzMZ2V1iZHr7zd8UwmceU5WqI5x0buQl12IzzMx
hO1wCku6eM9zhE5h+vsIp6ggrI5qakg6itShm6vH7l83p/jQNIIgLiysabBQF2dg
E4yJIIGBmnIFz9XcwbKd0m0i2ua47NNmUIdm6bEJYdt6a6iQnGy7lSxVxrGwWkRp
kQXmS3d0ZZcy7FInVHLWJcQa+F8veu94TPXo4s/Q6z8nwBDBCzukkJVyi14HXVQu
xVCb5Qn11U4e3T5IBy112dp0pKcdV6W/u7E+lRU2itadmPh4UyTaHJny18VI8FSr
w3FxBMbNYB11bGVXWZmRvwzNjSW9R2hNtFmVqxYXYsFmdQr99c/tm7mJWpT90iqz
+AEghNl89TJ2hr/bzfMUfpHYYnSOvS0GhqNR06Whfu/coKTEyXuvbT5DlNg0/BX0
VZUPGN4cxz/4K7bcs3Dpo2zNEbWOSR/+cqeE/OkBWA0N5bjERRAlxop4xGWgbhIF
ysD2cZr1h8s4TkA/l7Y9CTp+t1/W4dyc+AvxTgUUFuXc1rptMoB4nZ+M7j+dFopg
nB8a8C/ptv458V+L+L5qKUqxuNyqRXMeJpT615yQR8ivuAsesxaJTbEV3hk5XUbE
hGqUqyTsxM1ZYY9zQPGd/jo/Vccs+JaiT6ev8c04S5S5PZL6IDzy9wvQClZEPsnB
N7FtV9/W1ODPdPwpLR1ksjWYBqLCaHsf7MrltFbGxNIxFmdHPFBe+h8MWbcRcKMc
gvFz3UEhTcps3PpYcZdObTJmH06rJ+W3kADHlAO19bLYJ/IlUjxzwUuN/A8SmP5p
chiFBY8M+RrfXx+CXMEZ7WosXXsHcFI5Hk6NvZH9KAatZmpi522Sm5/2LLTZqhSY
tGUtVYEg761WYP5CFF4IuNQ+/IY7CO3FKMm5S2XjNM7cPIpeyBW6vzLIBuNYRdnx
dnwYijdC1LHabPuZ45YstyygruFUa9YNiaNQWFa3fkAzlZLia9DXGKpwneSNRy0D
5SHTYuC+aMLq/+Ir03AV0pOtdgu2kgRQ/h6EctsACmL++Yc/lcfOdRk4P2R4xtQQ
ABqADA+Phkqc88MZls6md+K27F3txwqqwdvFCk2p/H0eoDCyFdLTC6OaATNkPefl
Va17PyhDY9P/GQ5p6S5TlGTziXDQWRdGiB2WPx+DMh8veAYFCRalgtJmvNOqWRW2
7tesP7s2E9ftqTChpIUJQursSifert86BBlr2u9d8ErkcpdlDUhc2jpuILLD2T9D
ENsSdpZQQU/m7t2aLZAoMyOTclk9vpNzhvaHxBBG0m8Qqn9wO4+RwCulkPdVYJgP
d3qCq5G5+cBKryv4sFIqDTkBR9BCVSd5ZwsnqGbToFHKTBNDVljgqEDRjG5eFp7X
pxlEdI/DeVGxifMBRG4mx7U9EVI/AL8OtNH2ZkHoiQ+iro1kxx9/TxCMefdSsDky
GHGHH89syy+EGsCUewEdSdSdDkSJUnX9uJRgxGfcczki43YC2/3Go72/wv77oAsn
OX1VT92V4omFS5fgc7Ft+FkS6J4WLzaaqWgnugqHFqD+mWvO2vf1BRTEEpntMnDD
T1H4MqGdyz/MSSB4x05AtwfMCYmuaksnJyEDcPQDaNc4fUJs0FRKexRRnUjADO6y
yKnuXibuPwn5ICjglwt1iqB9cnHph6rBK+gYsmrcEaFCxkeDoslrciuUTnRzrA+s
5RZslGV5TDC2GebREp1Qs+4FH/oafXPemRIiZkT+i9vcj44jjohKP3ROppTSqBg6
abMtvbTsVj00PS8Oda2Dm0BBjg4wjtG0bSfhKP/hqz0r8UrQspdh3C8R2pmaGbR7
co1Q5IM2gmdMM6dAQzsHNXAf9UVTwl33B9eIeeWU3HkgoLyp/lkzseuvqGIi7Csy
31nhFWTQotb74MDHqidNDr4rsQguKaTegPbvpgdsTP4yQ/Z9a4s8gABQx6CavaPk
O8E1s3WszgXa6RBmMN8hOWsCTeDpAA7kNnvs5lQMAWjMLUNL+OLt7b/hTVWtKVqs
nsPMLtYKk2XKkRjwefcPJvv9g1Xvbt7lDRNrzf+t8VbAV46hp6UyHKGw+HCcQVKI
JxR1CHsXE3CYOXkBbnTz1w/bolNqX+S9+iTUQV/oV3zlGIl3LFvjsRJcu5yfin4Q
ckjedBlaFe0ijOtrUwNlOtjrA20ufiuxKBVa3NvZC0o2mrqdmTcQ5Dwi2XQnugfz
LHS8XJ3pRd7//c2e2j2TZ6palP9vXvzSLV9k66piDxL9d4CdObjSLkvlsFf9H+bL
Wpi2yJpztXSPjZ86auetQbm1FtLQBL6AwJnJPOJy+jWKWkw9Y+e0hUW84YfY++Kr
4Ir5Eq+iGyBZcVX8+CQP2+CdFyDD9AmyF5TWI+AX1fuu85SK04z5ce+usWieatgG
dJeOpQPGVqqjBabhIKAEds+8bNarSV2GN5Lw8jK4LkuIWIuRSbfKP9GSw1L2wJFQ
t7n0D+3ac/IvC1iEmZWgBom+eNSa2FG6IBQDaxXNkqxwwuQauuPFQiwfqkCEwduw
lmGpOYx1yQXSze1hWkLQydacf1YjjHCiviXC2GG3UHrTUic4mqdxovXV+/mJIz4M
Q01UHpjfnRgND1fdPwHRvg7edSKSEDHbcapvtyb/Wasz1sOAKqpPYlUnDi0T/B/Z
bBCvNyXF3V3EgnKyapKr9wZ/N9J7x6uoDsx405eWY6UiPnh3iqeEE5uNys4U1RNr
xVPLguSe8TxB0HiWzy8AHuOehf0IM2YwRk18v55sWKq/r2cZlDMxdFOHoAYuFg7o
6a7Jl5KmPYRog6FVaMyDZtJT9TFfrKrQtshX8XJKGszyqZZOnTJb510MxrYlGMgk
NVd/bXaqeeb04+TiOMLR11Kl21vicxpYEpi7jJV0gb5ggiVpNFdOoI5t+OmLB2P7
ChyTXe/TVGeWGW5tRlourpa7hDC8UhQLFqML+SakyLWab5FinFQLD5Bjq897FiUn
sZ/lL1lNjmMJheiN3qiz1yNqu3ZdElRRy4geeTMnBAHqcXI14Dt3vBz4VD+sNyBk
nBMserFBpEyJtFNeYF2lYXQW2g09PrLeVvDDT1UsWTKwrjZtP9tAIfne2fELOxLv
L7UBzxV4Zd89hPWiw5VY7ucrarQXgqvu9SEjqNrDtfzUCC31gqwGDp14bUKmz1B7
3adOu4BE1aKPRa7hWDb7jj2GQQRakuO9aGhdgL/ylT2q97H6KxbZptjC7iOenBLe
v9wDkdIKvJSHOzBv8Co8EBcRL9efGmKWIX4NyPxtkZB5FCSR7KLn38u45p3Petek
dHP4lthvzLrZSdYg4TP5n5u1fZXFW9wiyAppTU/xfGUahtO55ZX1VctRZTKf8Uwi
nxNo2OO4djuSGuevvjAjmRW+RZfBPkRBjvtNG3Cw7eXbZiGNQpapCGUfl811e6C0
1j9TtSXYBmLCGoZ3tpX8Bjgl0kJS2CmWHP6o9lCu4fOLDoouU8LoOeUp7qrR3rIk
biK/+hynw55hA3q1SFzJ2czPTpYIVC4pph47Uhr4rVwzsDToN9OgqbM7Km4XkH93
JD8StAtt3NQdxQ8i6mT4Aq3UyOD6PKerd1ph7/wskOOE4CsjGSaKJh6Cg1cIsrO4
Jt1ftw4kGpX/E8ipG+hkLlgCsyWKjcR4SyaH8srTYhhs5WWfYQyeZqQMRFQQfKYc
xDvXPQtqge8Lu69oxgZ8x6N5dXx6ffflGZc1RbyoXYbE9zL7qoKoYHki9KLfTVLq
PC00RJBxnf0KFX8tD0XhHeOBTUh4x7tVBoGC75wOAYt+HWEsRSZnb2xDBXY/0+Rm
U5MyI/AzpFVMpd2WXjQRDLxZsI/oGSzRPHFU40T6C9TD9z1XQsboFtHMt2Z5WTiV
7WYM5qQCWfD/gW7bJAyw8huQ7OrPYBzLRmw8KdzwuiEIaeQPClvwHNaduu0/41vu
+5jhkwW5bUH+XSGqYmHTvYqz+n1TEs2G8fllRhM3s0I/3HOVOQt6QceQIqd8voc1
LhmMhnrBYlgFRKFrM2hpxdTyNMq8WLAhhx9lfif657rH2omFfvuuUInOnxeogwpD
cvtGOVfkuV5hRZB5mztoIJjrpuietpkkaVaFPN5c6/OIPM9JBVeQBCw6Sb1/dihz
F15I8Zk81a63DJmSgfQq4t1EqKsOyS2cRNoMUWQNQ2pNmjv5SGYCRcKALApBxGuj
6J/2HJe/TvkubBUtpHS7oLTAkBQTLi04FWQdmpD3SiSEYDzchlgEutDTwRRQdlZY
n+fTjCqW4sr3MwofxxwEkagO0CTAeJOseHzEyW0K42VcX81ZO6d70eJ3Ov4JgbYU
7VZFcGekAzkd8erRflPVdcj14IK1htDDTgQtWnjKWW1UoY9/FTBhbI5Nx1csPbig
GAzlTZRiRImFBlL9wDC42XvBkRRamuXWRUOeg3hkLmECZMRO5GOF0qskn2YnaV0T
E/mP3Qw7pSMk6+0vvqKW5kJL6nyCUl9/58pP2JtgL4J/BZCQxWsxznM1tYlqGTCs
nObwVKsiTd18lBUXPcXL7lTK9y3JknUkX8CK0YSSDV/gqKOigJf8RAbWuD2U+oQ6
c1RLCljCpyw809/3HnIMF34UfYLddndUNIuLGrYTYBaw7JsISxpOTDD2R8gxDCl6
QGO70fKXnLMssaxuOyW3zkpobuA+q+k4/PbQtvi1ABlrSQYAflU8w8yzCZxO1DWO
p/pyH6LSytYvMLvmK0/u3niXsqaKDoW/RzXVvMetTRmw9qc+Dcu2bAnPmOv83KI6
VpnSAMHiFtTQYDEmA/JUBtZ/QM2Ng4d6mrdkugtUWjIBwB/73XKO2KZjZgSBAnRR
Os0H9N+IT1sOPGxE9WcNP1av0bIHnxSiQYNwxBbuYdOtg3osLis01J1aiq+Zg+RH
QcObujlFkSL4rziQovUMSlmqIQYjGLiSmYAAskuO/wFHOwboTHAdzO8HJcVGvU4H
PhU6iPBIMip5ay3Vbn/fgKKiw63I1SMlcZ9xA8r7dKZtZ16Qi/Xde4KPS/0oyCNj
CPoV0sG5dFxmaoKoKUh1x6MgWyfZVrO/eF44ocXJYS8GNv00vZWtCGKKjV1Lv9xd
hOWb7CfNyXiMGmslyhkVQaC+GCFxcQbNHcN9FG7SqiTRpCMYCgcfcaliSXSmBFvS
Bj7iQDs/4JlRO4kJHwWTFBGFRoMkRnQtvbKNZtOIyzGZ4km+zHfcKKBWRSDe5gNZ
H3wPn/WgVByQymiFWUiy/hBkpDb4rCvyRPm4th9/ZxFYYvL3Hprh66aC5/KNPeqC
553eUc9d5sDTljd5T6HYuuJHjp825tvFV+s1BTRCPJRphsIUCxBwo0Gtny/cktwA
VV7WhAuJfzR5kf0fTOTAeQ1YQFQ1tTzeDNjvO5WFmk2qUpEUBB9AnV9wmeQFbf6D
0fl+3+XOxU+uaZ8yyA7pJ5yJiFI8cUCK4YNkf6wFIm/oHlX4AygYIZXsqg69jyLj
4oQZJ9W/MtnpaBW/rZGQotGw4ShBusejYoBmL0qiW+nd8gbvngG406veR4vmjNv9
zSwsiviz2sPSm9HjxXiCnynT8JA44raeOWLM0ukwGkN769vmJd+uvxfbXYuOnBPo
SCDSupTU5BoOrJsdwP+08YtWBbQz6YfyKFcqm2UC28Xn2R3G1RLyP2DyCkE+kXD9
nci9TX4YYM+kicQVTLW6B041kPMu72TC3DAt9soUyX1imzluir6x6PdnygGfULWM
6msWF6TbBefh5TVb9plEiF3eKKG8LMPXd8Lz4zO0M8kAEAZsz/cd9V8xvH71MS+1
yQ0ZIJ1w0kmqx0gHRps/kObmtuq81Meub5CdTtn/PeOWx8YG8oxJnfIcZpdWovit
D+NW4nsxZzuKEc4WxQ3/KMGdkVJo11YSX11UfbLwEEqG/R7X3okQ2B1mQycx4Pof
QtMggiGvYHIMY5YttIevfHBfIqI+4mC6g3Z5KuQHtG1DJEZ2mTlRcuDhuIa62JTB
prkTlGxOvBgqjERSNNJF3A9wkH/vGQM3pSwY566eWdNCw6J24MSCe8uen+o61XpA
+NG/p5JTX36qt75inDerErkR+kk1MZgUtY5k8B0AtME++fI9McEviRla9eq4teu8
SHchMS02L/mjMW2jgHdkvzicRqF+4Y7yk03FzTQXu5d9nVOprn9i7w9K3HqlyciB
3uLXpX6RF6R12Oh/2Wx95L0aiacjKo3ZQQv65OJ1/pJrNvGzGKkpgzc5fusevkxJ
/OpWZfuavPk9XTe8oSILwAuWP3vBiguckosMVzfQ/BE7cB9flpibpfNVtJm2KbDb
3+ic2WG2pIfk0eQJzsturuk5TgHSFSu4AAOXg5xphCns8QT4z1parcnL8bszYmNK
u6uXQut+G3smM24/08Cr81flSuYI71kX3Qr8jw6QLhSHlkPuIlciEalCf2IFB9su
cnGtcwz/wWFkgr1en//CYGY2N7wsCvvXViK9mF84PkT03kxDkqvx9IavO+65JZaf
PfjWMNpo9J4jhhJUBDJ+1l7cC1pOHxFjunlTEMIC3KTh3iD3B7OEcN1ZNsPDQF3U
IDSX16GRLX83RbV+4bUkQUdtrDu/nz8FNMozAxxHhkKmFQ1rOQU6ykQCwYgtoUIV
7bq+AzwDIPc7iI3C1D5+SC06Kv5xRBV90BTKlpXTcJ5JZMkSbSb5GUzsfS/ZfzeQ
RMRK61OG3YdVeVomszlPOJhohQwXeOuROMwfzU4z7tMSzOLKmJZ4IjmsBfjatml1
y+9S37m6GXugaImQ4x8r3ujchSnz9jyTKUE1iEL8VEdbSRXSNEpczgAMvjlkQD4S
L5yMLi7e3TDqOC8akIU6sVryoLzLG9w9NQrD3vm2ZG64crqAty3VtUELfRDlcN3P
TmYff1KpaZspm6lqeDsYmGsRnIZVji2FWxYEs7V6F8vy2nXPeuCeXnwzMAESsKMR
RscS98JyfzttlzwzAfvdi1JFPAckEbhYv0Nm5zaclqn9T1jVcnOznkyOrAEFXQUm
9JLk8bWeIG9YoJ2MY83lp/DhcLzV/lUmG1fWagnaQCFpWSkJVS3seuBJsbpnemp0
J8imjDaqcQpy6wTd3u/Z2n5d+vkUV5EE7hiyfCHWBA6Z7A+dRxSgaaqP72+Mj1CS
kwMLY2rwx4b+pZ7r0e8UjaCOPqdUCAtKbqN2yiOLHVJ4seyzVJeGhK21zEATq1NS
+syk1FJ8W+Vcpic/LBzqe/FrlRJhKaQjlLrs2uEXbUijNQzuibCGwJLiiVAXHoes
Le+XlKOriPLC6EKni1ttkMOY04MaVKGzqb3mnDP3YmAGcsuOPoCh6VM7OXSgAhj/
1lK572VJq76eEt0xgWZdr2uufH8UnDFu8H5+kKqbU40wz8zrC2yws3xd6/waW/aa
s2QQ63PhR97Gkwhw9YpzaLXYZl5gJM5MqiaALpSffgTi9GIBoEv8pd8b7/LW2Urc
E/C97h30ToQ1ZRoKB90iSu8QxCq9z47AbZkCI0zHSP7WduDqyQYf4Y2S6+pCTbF6
b9WOuYjbG0e2NGvc7gnS5XoFspEggIS5+O/3uFKix14TDWkVrj/cJRmCjLTimdi/
5+AMfrKa/7Bs38bbA8jhU1DeH6dB5nvuTo6WRBJVd2WKzYGnUa866npq0OJhDih9
6drynWUzwgMDyPlgVZrNVWFyuoebJJRCk1Wt+OtT0ft4yFEi35d2mm50+hPtVMvp
PAhCRdJL/h8rUbnWBZ151CEyuEwboLuJsbRQwC7WqBZM4iv4C9fLKB9+RvIJshdh
eSXqXtxJHHAlfNVWiDP5QcABnqeHrt5SD7xYCDXA1qS7fLBgxpw/nQmDfv+VSMdQ
zb+L8RdvJzqZl3dUbr4+mwdx6n9EXQZLXq77jzjb0koBn5kx0HGy9x9WmHtDIdMq
HBnzIQ1J4kPTarwogZRFtsV9C1kANtcl/pf9DPn5ZpzKxoHN5uapZEWuqbKzBWOf
NVMJbQcXaibhp2a3PSTAcNCjwQhSq0Ka+ILFMIyPThIBoqfSM+SeO6YsXZniEF9t
SlL3MSK2wOrGIiJdNdZtgyccB2q2iEXMsn+BeUj1mh8oodcO7R5FjAs4vnEzby39
aCOScp3oQ8aZ6NPMzFROlvl9eja/YeW3DxswSbC9sCzSPBnXCnetUc8gNXpRp+56
S5zD/LubO8w+perHeQzMXa0LbSNsmZP6Nfd7ADloNIx/QKtVEfvMMRvjXNEn11IY
Fcu9vIEH40iVsdojreSiCI+Fh8Lc1rmMz7qH1UO+9E8Vf/ZE3dnkL3Yjf2QEg7k7
x6/LoWFsbOC+Nm0ud6HxKKnIjHJr8e+KFUYHrWDsZiwqWpWzh22DKMy0uAMCs2i7
QXzep2RDxxEiqmyckUEQW4TZ0FIar2kW88B45cz+Uaitm07mw1JR4YJ196YO7XeK
tv7TTvH+ga8rwkWMnnUGidxQohObmSnGn61SgUTR35KHFoiDu5fIGuGE6ovRj6+m
Ge+y5kMFaEl73ttDjFvt+IPcqkY2MDrbw/6A8E1HIiZFK7iRuIKplxhll9qbkmNU
xNkGJ+WkUg8m/8Bl5PJctm0kavF+ufm6vsqnARA8aA+YbQBcW4kyalDMlhj9jdPC
fDqkYUV6ycdIX23uiQCTBKdX2YRb1W7o54Ir8fYx2kZi1avqs4PgMpRlRxYeMltL
ldites9jOaDAfaCG5ew+MqnLEWxP6l0rzD4SZCj6aB6ETgesuZZa6Zk3e9p3yEQ/
4TCWPT1ssancYqm1DmMrmVyky6a4f2HXywSkWL7zDreHKCtZz2GeZFy9V59h5IHx
bMrcu/3ih6MzKKCxTSp4a6zc2W059tHntQILWRb9MXqvhllH+tWG4O93WbIhXzWd
AtFCO0ZPq4uldmtQ9lGYqXQgEga49n0T7tGqCbJN/CHbPQqadcb9pmRNKEPFL2Xp
92FrFFVXI9zSa48eaioBnknUq89NG9jpJSVPJxZleYrYyIH+eRAqJhFqIzEFnQUG
o71LHWY74pF/d2VyQYeen2JwvPGQl61YWPT9RipJkYSzpesSxbvScFq1oXWy60MI
O7xFlIHiiPCkESonYPJiLBAl6Rr+1NNv5eYUJ1ys5YFTg5G9iKs+mNAQpaJLvGu8
6GtW5p9R2i1SojihhlCAVYsttwCjg12zZXPJujI9et8BHjdNPpZug6jFw945GhTd
opMZ5Xrh2BqvuwNfCuvry8s8ty7c8wsnq7SgcoNfyK/EAfJOsVrDkBRuiYW40xkT
misn+wOmk8EolngZkf1aBjFuVlHe2gqZGU/HntN/1BNvxGZomdybWd0OpfFpDTgW
Y/pFvZGLr7y6zAPlSKtiWR6MGObZcahm8ZAx6HSmc4frA2XnTkChEPHFP/IO9KKh
Xs4If19wPALUf9fKzYB4nfNZsdpGHRR4K2KMkAgdyvzAeQfofjGQ+4jXFC82wqfJ
s1LGK3gOu1o3Nan9nceO3r8aEmD2M/CwuJ/Y3w1fZ15/8mkMoH2XhNf6mkK971o9
LGShll7OM2DreiWtaObE62t0lowUjQUwSP6jv53q1UuWyY9S/8L+NuBa/KLN/vvk
DOeLjYkJXIxAXPKm2Xj1vL7xnqILuCnd69sCIB3UmG3EUc8pQvGPQsp5TyTYmmMI
mCdWCtuTYfwxMS8yXErL5UlmAEjamD2idMB9yHRDJIUNHz5LY91bVLVqN/nEH6lJ
WNZ2JVW62+8zuTqEX1IRG9VZ/hpMcDKHHUnB4K3uKLzys7Lc95qs9eTZqmq3vN2A
Gf3uRn6y9tdyrAsnXhin47uFIeHNwTJrDxFKxj9XfJeqz+lwvh5v3oVXCtkgWxqg
TeRphLSDk00En+moc8hZOxWk+dky9P2cb9dnM4cL7M8cqm1sHMU7giPstlKlSjJd
OPAevnSQo6Pflx/wyhzMgL5f2Ttajpa77UXLDkJI0CzpZYoVIeeziyNdcloCHqhc
LSWcRjAPyAhSWJ0lLstlyLosfQZ0apXv5HueTMJi9AUGBS95awAreg92c8T8M/Ci
8DVQNUZkzOiEGgxMSJ2fnXz5BzzQASlmCcGzXm4zUUd4DG/pUS7ma/UXvsyDQ62Z
kGPiNCCdlRMUsDXRahXqUJ/KdTjYlXnKxzNM2sM1gGOQntn3U20k9IuvfZapsN+z
NTaUC6BL8795EsyDKIw9TEcEd9xWAS+/N79jeUP6Cq372jSzfuHzFL56BYgThFij
U5Bn4VcJe7GT/OgSUPsz2qJQ0EQ3D47PF/HVjokf2kczEXDgqsVy1RYVZlfHxcMS
bQo2FeEvUUtqB0VCp8a/ceFRfKML2i8WUY56ntLOACOmPqyYHv70DX+QVAlkhazF
RzLEN6iBx2p5rdeb8UhYFbGnI/2Jxw3GY9ZahBcC4QxuXqqUi/uZvlwpm3JRfSK+
GpCJkvi2UBId8Z8yf9U90b0ff6DjavUTcl62vGc28yKyKLewUmUMCDkVUv3706eN
EQ3a0H89C445rhwDg6sMAgyXb9sP8CgCUG+HwIsE+PlKMYrhk+UhRj7HMB/HUNah
seiU0HPHH+nj/NixvcdQutYy4Q3CqefEDqjIc5dN+NgxXPr+NachgKMEEQvWImWT
L7/iqJFyJurWFYd+NbafYiUFlnKvfHI6YV0Ha5nAYM1GeVop1zzlogJoo1aIDmMl
qMBHjvQyvzQfbfSxG19grpBoI/aQ8FJnwBcC8qPymCFEe05v8tf23z0qEycJpoOO
qH7QSODgGAn209kLLfilmi9qmN2fMkYDd/admm6bE4Yq1mQquh3o/UUIL0xLvxxS
JNgDlegA934qJeNRdtOi4xWlW7PCce6NkRNaaa/5D6YgiomOlzovuoD7g4w/trs7
w+OqqsPWD0SfxB43xsqx7eE7vMrK9iysZqkifdAuWBdzwpUOZtaYlzzl9NrdEQMa
OYgAp/VNQNUugQoHMZeA6DdRSVpmjQ6TsN3Y67zG0O6cZybBVD0Pvd6R/bhQhQIL
exCAH7e/oDn0OxRYok5/AOwtA5jjtuZkBMlJuCuDVhi8qQwbkTvF4WoSlsCDfFaD
7YKQ7izC/cHbOFJYqpxkNKNNfedAT2lnP0+9ALTSFq3+QtXfASTjnAEn+Bvq+iMy
CPEEUXNojtSvFq0T27PZWCM2IvRVmLRA8ckyeYLzoK3yuQQkUBKARgRWiB5DP7Sa
DqsvQO9BepNeQBTipTiusAqGPMnxnORhUAE7MKZiBkt//v8RX+jzBMmhPcoqCJMZ
B7yabrI3l+yxyb1BN92L56qK3GFr8RfugvI2IiziO7UKneNwrbl46w7gRbejamQ7
prJZY5MOnzpqPyZ4CJcnfy/rqr3FaJaqEwlmHAYqVbE0rdIRyqyZiGp1+64x2+Nu
kPTWX3MxlkNMy2+E1LXL0w/ta+tisczg8wi+CPEoxJguqVmTraIEx18d+hfdhSx5
IOzimKg9mGll+PRCsfTMrKnWgUIwFBZbxPnsRJC9OFgFna0seePcWiRUI/zlLWry
pVD2gOTpThn0P8T0V1nBUnJrzZVPF8C0YPI+ifGr/QXyovKaafIXE/wbGAlO4Cmq
QlzvvqLb5QO54ejNIqlv1/cwgIdR0pYk59oUpgmtHQL32LZBCsnOQX5WbosdAAse
i/NRk4VU3VzfRUSgvy+E2Aw8DRuQPYxcGbsm8PkaRua/O5wDztYdXf7AlLtEM0ax
TCWsDZQOsGzRygXicF+lW4G8ebAC9Ek8JcqJ221I8Qah78gH7JTHzsx9KpxTFqSE
C/deJ/Q4PUDbvHNdJtAad1KvWx6CIWhvP7NHqYb19WiUjInBBmiHXSTXf8DJxb5x
ifj5ZzaLq3FIpkzJ8O+86UMka5aDijqn+UHKllW7pfEtmkHw/pNZZC6MO4O4HhDn
nUHGGZyuulrF1dd5vwhRHF7GiesBs0mtPjs4NKES7GSLW2xvLD1zYPyVcoKayDNO
Uo6W0D6jEa+B2t8PVOz6UVh3ZPnAMWV7kKyj3zpAJWMUaM8MeSDHADmOGQ/i2tpa
UbSDKpzh1/wVxTPENm0Qep6gh4XlRlsE4uHBgWg00XhTC/dhrkQqXBmba+K4z828
VhwfAQbx2WEwWXmAJo0gSiU0b6vGqttEykadFEufEiH64meYIB+nSy7tX1Kpmxpn
YR7ZBZf2LrDViQr/BjE5+psOvqq8fgsezLRETtyQOaB8/R40eBf6yzF5OFSsBZc9
UBNjodlcwuIwwbyY5Mur2pjIjLPOoNDoHWveypxUaScOVZOkWlIMldyLWJq7aZcE
R4bdjbu/3AyGLj/62hxDL/iIJAbN4+9BTwsUBZMN/GkUNUgg1UUhFeEP6yUC+vtv
XjpHJ+XaI6S6gN1wi/7touN6TaFdV8XjlsXvHuAPHtixD0G5asqO6rmM2KHjv80O
LEqnSSZ7H80E/kZuPXVOtBHLEZzUgAoqvALhFpUeqYULylCIfKW3eXspk2ls+kFd
ceSr3WDTVNUHrUbhAXjMWlhluo8Chgwkl0ou0/EhvVtkM/scMh1+4WLSVlLPK2+R
JZ/DiU8jPwRyC9jdLMUQJ/d7UhDWF6rWHDaI4F9vF0kXOkbKM0WoMYP7F/IHU/qx
jkGILjusOvGkgvsg5h/oZi+488IxBfZZtX1lZLSMVPmgREH/1lvykpz9Ew6iCvTj
7a4w9yqJxtTb+F0ArSujasaDKpV8wSoF+UM01MVt98cU5Kw/irQYrI5FbnQfIgYS
XWQ14aXmp+zlhSMWuYQRnwTKPEec+tVB9WW2nMECoC9r0vTGDrxmmkeUI0md4Qgn
bpbPVUVfOzwuRf2HnSUrg5c5Y6llW+RshIj2aXtB6e7uHgz8IFnRqiJvDLdc25G8
lveFViEjrAINQhbrfZEQRcjNKfrXDRWxJa63mgBYBApRsLuBRzO3iBOx99nwkfs1
2jSujwQMFFoI6R+SFWVogtE9D280H2nDy28shm1NjfqMTOGB2Lt9y2ACRoiJgAb/
W9nuBGY9/y7tnzKWegz1snGSn/d56skWToqrWg/+o08g2uZyuXwoYMYPur5m4+Dg
8wp0Pm4z/Kqm7UK46INZ5sZfwxPe371mr0IhqAuDNYlXXTPMpLMNGDa418f++W68
n27OGb+SyN1uO0IqqK+1GfgGxCa8BfgKqgVxVTBa0qT2bJmvbRKXyxIYQ7m4nmav
3tE+xkvGTHCVGJeScZkZkzTqmDqkJHhCUsopBFa7VHwZEMoDLZjC77etpK4zY1NR
LjCjR7vA66FfOrvD40xn684QMyIp9jeN+tWJJUZpxANiSKYcRP1MrhvH7x4RGGRQ
kHE0i9yndawf3wED+1O54Iti+VbM5HJJgUmUslw2dy9g5evYnF8/P37K6BZXTofP
VinJphihcgNqeLeI+QAkBYlIA+3r5p/F3e9otF5ptfz1t2ZT/wOOlszTI8J4iJWk
9dsrpjvM0P7n9Ie2OSGPsZbfMtZ1wxnz9sobkTa7m4lPmQZyMfDxsd+CjtqK6Cgx
4I7bYvcBokJQIFcrvJkk/uBzA+Uf21Gr8oU8jnKhl7RQqaI/fopSnyNMWVRwhT2d
nGd0u0pORsP09fqVTxBwG8MVGP/0L0zyJLrU8i0p6azRsjSZI7qBEupEodORKp9w
XHE3irCUcqCAavmTdyYoRxhJ6IsLSSgFTC5gsEI9t0PFskviQe3CtIDsAZBm0PQa
AuXP5a5mO/Ed/gvq2JwjwaV7PaMh+QZRSBlU7p1fSmMChFBcq3UwS51p8HR7nz3j
t2e7CKlUJoKIzBiaPXFOORLo9ekBl0rdQaMKVpYxi7TAKkjbAoYzo0i1nH0rxwgI
ViQEJZ4e6XnydH4IIqLoSL2M/6Kkuy340IXzMEH2BYVoDPK7w/ilufqkrB3IvC22
6w05JXlVvTbzhnZcv+g9gxHJck6PE3vEoIVVXynHdHKPq954p7h4InZSfK6Buu/x
FEHP5MbMSL3LeYzjFowoEOLZzRB0tkCIPWKSWgMYbodgj6OgOpBItk/NXtI9edTH
Ym+ueMYZUyAMVpOTBWLZbhdS5am3FiYPdYRnzcpnigN9v8grdHYtjxGyu3Hwgtdc
n/VGMPyWFlu0v2mZmJjYqmp2tCkiU3AoglL0LaomuadBDemI9OnUeASRVnxs9sTj
sTbvMvLdiomV0I6pZZGFhnvyJWxZAVmozQR/JgUUXBHhKMZ0JK9Sb1qeeBkq6X2d
sQlH5ANGtXPhHZPyzSe+nK0J7P0gOqGqVwUeDr0usiJypyVYQy9y/Qa5Vs701UEE
m2L4fVY4QFaFt7t/hxlEGbF3DKqsVbELN6Yg14NDIyZF+cl2Buy58BI7iWSN4Z/7
rkOMig30HaC1FwHfNyU3ej5/EmuBYmkkWE4PARl2UnGvZdJfWBIGnDUno1gRdsRY
WA6mpwXR/sBWNOi6knMDFBho0fnwChrAfW+ft82AmHHzbHGNr9AjKWz69YT/GD+Q
zclWSrNCeHLou/bQqy8vq/s6oSPw0qYBhm2QyaiMECP4OFRCCJkWjACVtTDtJru8
sBaboBcB2nI2UhfkOspxijJoTACOs4tQAr2/W59ZXPgfh7RHwevllu+Am+I0Is9w
Ra9FjR1lDfCcxcXp8k1p+GSGk5adxob5K2rbG+je8/RQaeE864iEcxAY2WKDmVyw
+ZMGTjFEs3sUBOOg040ZHhThMSNhZjFFzkFBxfKM43DZaM8NJ+fWbh9MafUSxV8I
7Yfdlk3KfM+j6kdINRtMan290F35iQ4OGkJxkauQOk/2Ba6cRRMHKIX4hOiYdf2j
ZjcjGtE/CMT4nj4eowp36A+kB32CcRatVBGiFODlavfb6WQxiPGBGShinasOf0XD
v9LsZ5VFkx7czryBZJX9Kree8Qm0wsJRCI/4c9cJeAYD4gDkx5vk7pIYZZ7ekwkR
LA800bCMwBjWuGVZvN0wQ2gDl9uEOgSj8uJLcxQw4lVl3PnfJ2uttVOsObroyDRp
WxmmNTUoFED+D2a5RpZIzSNd3seQc1RJ6Kpx6asxCJRuoIWpIGEDhbyLisDA09di
x4HFr6G+iYGl+G8duf3Z68PXRtRBEK4D3ny2YB0BEA1XUVYbxes2n1ZKR3YEWyJo
Ht4kMsYuecbEBCfo7+5Bmo/ThFZzW78M2cAlL7jVbg0rYRwMkGwfVIV9Pn4htldJ
ya+gWEMAllKwAM9WIel8NvzXpffbp5hXFZRI6f71suGJhSVW/1n3tMXf5m9s1Qbs
EVuUuO1/S5Po3q9GqX/Yb2qYsYPr/W7tqg03EpRaj+VA1ZCUQNOPYJVwXC3poVK8
hOQ5pcX8fLD/sfJCPdsavK8nSKowjcFGh+ERHG7Hpvd3WkEm3IiCRSqyGql5If7O
IjsQ/q7uIsYkHXyBtv0hqSXoe2yB40UIDoEOVsw1GgjIa7RyhQlzhtp0NWb0O5HH
2iaF+09ipyDM+PzLdIpAlKknEBKyFzA0ZggcWm9/gWRbwX8SjMWmwjISSH/jfNfx
f+sQeL8Z9+qqqzl69DRPbfg2mRi6EBQ7DD2yUhi3R/3Z7c1VqcB9hkEeg4i3nzWB
HG6aVgKWzIy4szxOXBy+F5BlPhO7RZIhuWwipUex5HuIk8Z1ohQpxmgR1cL8GRAX
pBOBo1ellTd/2PvPsPm2zjqhphc5RVudvDiVtFBPzWo+MacoXY7Xk0S3kP4uAudU
lbCXSmwpZId1QFfDAlxPOVauVDWPGggCGWnJ10h+hMh9oBo9UxdiZTO8NjRzMEDI
bIfzzZGWOPNAo/0Bq5XSlWVxl88oN/9abJCZBDziogo/bCAViJOpX3k63wLhCI9Z
m9x2htKaM5BOsZrG00ixpgWD3FK4LJ5N/LDAgQds6bXCp5krt86PQST1mopbB3OV
FqJm9NN3ESCQSwthhkL3Ft2aTb5g9wQPAO/v7yshfmfCrdFP334BiLKR6fhBrkld
BBEiTIAeNKfJNjNOAj//2sAU4/6NwyhHUPU5E7iRiW9MvuDH6V4wI4eFPqMMxPpa
PhBhFioUqGK5u+1O83EB0bsBQa+T2zGJldI7FbEBlhgmRup3Xi45On76L8by3MRx
P9Iw2wkAhlXpnuCMDdYMp5LsOXdAeL0to9gbcXg07LY54VMaGWndZKkWWn9FKQWh
f8vXUtC38AznkIWT62lC5bvUpZcMNHghgtEHe7Fa3XKRJLOfqNlVXN7vM2tM+j5R
lPSe0N3eEK9SxWQzo40V2Lgo2zoR2Nh5wuKqPyZWcTP8TM/hEJpAVEqoryiooSF1
kYn8aHpGoMkDFqbjFMcSca2yurqDLPa1p88C3Vzz8hhXmbcXo17yqAuEOCr9UmCb
VAjPhTtiLfLd8Xh/Xkw83lJCszdt0LFIPSowaiGyGFzg7E3Ly/fd7/9fWOYSxHaK
DK3krrt9USoED8dZ+N8xXH6ihJBlE9pPFSOwgCDMmttA4ysLVlcXyRSzO3M/ltGq
lQtJLS14oHJOsu0Xun1vc7IMEl4iT1sOkjRoG/YxXcF182/ttME6B5CqL9ZIBTXS
QKDvrGEKp1ibOUrLem1BhJ8+FtrD6KqCbbtdZFr2u+D64aJYv7dz1tijO4E/zvRj
sDsFBTx8pCnWE2+b0PyQ0TDtjcTchSBI8MK752jI4uDLERESEq1mOE+2bDn7verI
omB+UdQq5XIA2datakJcqJKgN8u6UlnbJrj2HPeBACYGEB2f1TgQuHHb8dsWKpsz
AchGMoLEFHixPy8BvVeAv6PV/4U8xn3JOsPkfa/u8GIxUYfgmD4jZmFDRLy4+AzK
veo+TujTpjMGkZAHlXc3fdghiwDoIMxIr7OmIUscxb/jk9WPA6uhxp6lJzpK8YbB
ndSi3CdGFrZl5MqqinfuoadH5Kh8jpYrsoKLl9wExQZhXxcPG4NFlu86vDji2OzK
KMK+GgvlgmZb39eHASkfNW7pJaBRD7mOXedWl0tRongXj2xUTD6uoIAdx1gPva3T
Hwl/iEohKxa5a86GDajlz/s0vbgaBCuw8u2uYTzFjGkWVgZhZS6ONkF9nYYMn1U5
ESETmVtMPMG9ECHAipC6zU38OzMVOZ4o1KrREQAxV7io9MAIHQRbHqdMi1QagF9j
iobiIDTCMx4tm0fnSs+XlhzD+RVphgD93WlF+SJGuo8e6eJKTq2oExzeMM0FcUa4
HaQgMo1ARrtL3HRqCjksIii001LbNJl7VFqjFNmYyeq87p6Q0PJ9dkbG5abBaVAr
75hcvPFhavF1Gt7fg4NhQOZf3jEByEeUd69DFRzxFr4KXAwg53EAKFOPv0a7i7y9
rEAoSeIrKtsZWhagZVSSbrGeRtmmV2S3PhU3vccPvH8PzE8BywmBB2u9ezr+kd/j
JUiu8/08Dfj8/TYuw+WQTxXHb7wv+E+RcSoiSHteU78UPXAb9bygvWSmq58xK17i
eW32DUuCzfZPQ0b8or9Za4E80H1ttuQpuPW6dh0N8LcfHJzqwmLiyxA9MupsEH2i
rNtChmDgoRCSDAfV2FqvZyIa5curuANou3YB0+uKGYtsE5bpJccUCbzladq57yOW
aXyJPu0aSCyKwfR2VrqitRnA/gJgHsHIeuk52mB2+DuYzPogZUflT+YFOxzW2SL7
ZgNixqLTwqYUPS6HBdO6PY+fj/zcBdkvKrZIxxcW2y9JYdslowR0MRWmZKqNzcMx
uunSBlPivhprq84sRgzD8zkxwunE/WhRjzgkjMEKQav+E6nBZhBL2H8SAeRdv2un
ghApg/F8EmUAltlUsqp2wcGhpP3ISpp1Pov/xtEVq7XQG00ovCtUOdPq8rEFennG
RtXf7uEQYLQLAWfQ4B3oGdSE/EuPkFmwrx6tl+LpfR6GvjTrS+Jgae4QslUMWi4h
HV/pr1PkgC0FiwmiAyGT8ZDETZjDzIE3Fi9AkYP0Fg7JO3bEYPG6QzBQ9ay6/gvj
xOPyd4SXP+ndJXoW6Ux81GmPU6Sv28ZqfXeqZgSLIjiY5x4U037HTL+IVte42kNB
oFVjT0klwDg+AHYk7t/ooEv9f0qLK+A8l0fRzpPio7rp3Bbg+YsEYIxT31LRVVeD
G2lFYdrrWFNh0xO8i3606AVGTZ9wdQAC+/GtZHTJLirXHpph5dEsusCOcXh84nIf
EUS60m3l4Msx+lRdSxOyDvbdq8X6svf6GSSMKdxD+sONgqqXwi3SxmPhMFSeUHP/
NcC9VGPyHm8UgSmCuB3d71WN6YyP16SiIQCkJjhuBb1cKl20+/549hHbu07B46Yh
WAPnGrbmiSbFprr73B0Qaw2Ph4QkldCqmG2/V5qUMBVQrqJhxiNKcw1e7PrFATLW
T3IEoGan/+GTXI4liuCadaLXpMjLowsoiygRmcThLnqXTwoo/CImPaToQFdlyNem
4XhH7p48CYgjF5KB0poGbj6gN8OMpG08PPQ9l5lktwaCwMQ0d31MwJwCfKuFwfz7
0TdeRhNA1URx5adkfUYCJzh6JXCn24rSxKqmgeib5uNoidyWKt+JB5RN3FpxvPXu
r2A1zdc7PPsXx0c5ZJIXwAMSbiVkig5DzkVw35taavdOef0DGl0v+HfSg7M3FGAl
7i7a4hp0ysrrazLGt5TMBtJ9jo44BUimTScCjYmd+dJthtNNvYROMN2FZcsq3+Qg
XRL2w9IE3A2Zl2owk4BDFg29r9sp2Wd72D4czY5gsm85rd9a3Ug97c4B02KBJnIX
cBfX+aapLJxCAEkH5OgqzG7k+W2UefXbIVRJxsc0MlEH7mGsGSMFdrVFauQefwms
Zc+N3GsqOjJ8KsUSyegxXL+Iur64ZvQkUShHqRI3w0o5/utIJYBxrLmou4hkZlQS
3alSs0CfLYJsfcWbuwxmME4tZ1F65QOQqtKh8tUr87ytOmBGxJWcshkvIBg5w3xa
OmDbVa21XdIk6MLj+kQApGB/ULIqGStuVMc6r7DZrV2GHK/8n6CTJehB5uZiO1Rh
bi2sYGf9ieMljjaX0xXwm5SrPEd6Jb7AnnFpnbQsXzaM9V7aHSUo6yjg91/erHxu
cjOSrL1fl6MArwJHL4agOi0G9/CgUF+1YSCw8c/wfmZvPiBbnaCSeEQo5qD7EgGe
oSg+SE7rhWW1QaHH7ZiCncaE+Gj7nbJBNZqqCMq+Q9ihtY7y3TreT1Qpk8bu/NzR
PTwZp56HrJPfJ331GQcNHv9imAcU02ETKzId69//qou7LbjYzQtisajXeDTjE5WI
qyUqqqEEc/ZANB+P1XxTpb5QF/8202sSvV97jS32OR9JxSUcuqfLa+dNhwqgs5qp
LEPbTLEuOvgGKt2qY2g6Bwc48omJaQaqTWi8VOZjpuo1jyo7/2vt+L97Sqfzc36t
JEb95igCiJ/xfBkrSjyXlA8uyYrPdeSVVUg1KQ39asCWvFVPjvx7sz1arRdHJq1P
bk5+zeRoVRfWniTH+WFXBrh6PQNX8SfDYVLECzJ4F5S6S8kDXh7KYQwO2xVJJ6Sf
431RNxrfU1LvPZZCV7EAUmqWTWuMGGjWY+LyL5mltyxFFzspiAJePMnsztemSkHJ
dbdqyVISXwVYPFkvW4xBHstTOsKRakgpSHOU5U/XU6RoML+wvG1jHpJ1A2Z+z11v
noAUpbwalgxg88CTI/gSoC0QvPHNug98f2Z2zVrfP4n6CulXe81nvxASD318dQmR
0cg5hKSFkDD5i45P3qixjcf9ueXKMGak0hbMQ2B2C8C7fbiacJX3+nSxUq307C62
gg7sP+0+J2Ba9vV5guzfo13HfLtckWh9+TwaOHPn5eoiDwRlLL0s4br2lbG+EZGe
WySzKeN7JjTUfll9LRFnFDdBrn/KqmnCxoM5bsh8ShoaBZmYfk/pMWSaQ2awL8cO
HM3G32WmXGMT2T0PV76h+fbbsvgrk77l+m2H2SWhIYPjLoVxWO13ebImUmo8RPR9
wrtdSL/gJ0A/IA+1fbHMTM7LY7C5ZV/Phg4vZ4ab91F2BIS/r8Xn5xLh/J+9JUr6
D8alK+PKt4gVIjKmdvg7rlZ10EFCT8ecO8e7fIzS/4WyEOM4UenOytH1XaFj9dIp
hwzOkAMmiQK+OomT9Pg0Kp8gVWE56Cz6HNMGGMacxVbuhBBCPqHNp2CRadcKa4Nj
kF20zro1Ezq5yhI+EMl9wa9/6nSi3o30d79bMvmXEcxbrcBQ7nbAx2JrdR93RD42
7PQuKBs+5Y591ghNHiDhYkAZsWodJtKx9hR9JRS1KpKPRUZhNwaEMsM9Wi7K6cK0
I3UUuR6JwK1wf2n7e69eI1jxWHXK6ZoqGY/H7D1nCLOSbgW/RaGZ6ikMJM39N5+w
fahgzG+1AtsEskGghaTSTys1ZRvJXMeYkBTfFb+y1iiJaPbuZwbqfxx8Mcr895ck
kfL95P4u7sSprlbrt4NUE2iI0zq46szj7V89ctfGRIQUSyK0Mdj4DMLWRGEIL3Ij
/XGveQD7I+74mQSlRiU6g1IwAaj94Wz5slU4q6OHASN0kZ8tLY3H3JfvU2cMSJRn
rCHb46SCLDrzXjY8z8wbEH3vWygf7QR49CGzxaWcahP+JtHvturfxGJUzuEL2Fov
2ExN6bmBZ0EQ3dey1zQ4QGHdX7Gi7rZFQzYwdI/I6yGsUBsvZr5wVMcgRCqLfPWS
6LmdtDXtvYOlGWEkfdynqTKArY4kQlnrAN8M0OssaKkiqcGtiYO7UH/t6OdcY5C2
Idl36Dz8az07VhaygJFQZHnrOvyXniZPNivEuM4pPZ+phlyvgXeaSfluKqmAYi1z
vLKl9YA5b9F4X4Q0gIxiH8PtNiguWBGLVyTvFr7m4VwZID/ZiFFf2WrmXdk0O0Sy
cCAKuRqrHOHVWDxLbcc8ZWUihsMBmXSJNF8ubv5krLuqIntfYtDDPihlWoSumNJo
DQgbSnRCBQmU4h/jmJZ7n/LD/1ZV/6y2YNK2dWBsh3B1zjl8TS3F70XRxISb+yfs
FUicaLKxkASrch42ZJYwNW7nsVbuy/pLzoliGtARFV+UpVI4t/gbRO0BSWHtV5dx
dXhNXBAYIsuyMZpRGODDmeRr9j0N/eSyJXR/IHdhGdkK9MoabYgJ1XqcH6pjwey8
NOJH6HSLU2DD96H2Cae8IRg1wkqG3CxukDwD3YrtRo8ZDoFyIdZXFCk5GcRV5KQy
L4dHvHB6IhwROjwLuSdYnQBjyB5qFYzXSawAW8nW1v70VPDgJrKfGv8ViiwpKYn8
aTgWxoERpegPIebIU40gyf2GD/tJ3CQHVUS1svPWhPai0kkalR/YMUfqlIqoVOr0
doabIxCpeftI8qFwfe0PhlFTzVsLWAtOIg32SsgPFN6r966QdzrDxA5qJEOelgk5
ccR1vodHFxvypJux0R3e5gpiP38xnwgIVscRbrvTHpk0B6fhzEtRHqMXtR0lx5xp
3+wqrg+G0Yg/GviI1ak2wQzSGfL14/t/Hr5oUHszsAQJ9nOLjmGhsfna9vck4P2b
enTlpmGX+pP2UHwjd+thx6W9fS/VckQRWGlWDwuEx3cdl0Uc6ZrGKmoTvjjirr9v
OnsrLGzePzgR7afF0sHnM+XuLctNaS3B/FvJ6rdcNNXj9oTvWrJ+HA0TmTtovffW
Hfgm1TsVPmTzGLlNT1j1sEApF7CaNmJqTxLs5VP1EQra8uZtEdhxOXTJupz1H4b+
KYcBQvZGFPPdD0yWOLhh12TmBclJU8lp6bPN6n4sXRL1pNSb7Gju60kivSSS02PI
N0/ERb78UYRwXfnOI/26XHu5RxMUDE+8wLFKuMnecd3x0q3hBquX/REeY+U2PI3n
FpK3Mcc6nz7YpxCxBZt9y0hmICdh3mK8ASpmq0DJUpuJeNCJJDibhEAVQ6On9RmC
Rp+w05LeKRmrVtshgdfhLWbcqtIOyok1RfHweNmHcuhWEiAL3/X4CO4LA5TYFyY0
/B79CiUtkd9VFdZQ5DFzSSK1ARupQ7pLfrdWDhZHVGCtYO4mIr6030pwVpDBxyo8
8YYnMZ3wvBMG1WQM+x8gG6u1ss7od+HNsbE7eTqd8BYC7PGXGyRoryjCdCRRQ/Rf
YJV3a+TbQdULE6UEdwrzddpUCByxpbTuvjO9H8oV8Am94TsumPKxnmtN5dVnVv94
rhsJNlbjSRDKnMON1VAwqy1F7MX2AdZlny4SMUYCvTBmMy5eKLAmsTwj/fwwxPpG
1o45w30BDpbwd1EeREUBUtWgZZMHhIJ5xsUAAj3ivMKqsp51lRxtac42k7bZnFph
MUJVuGwep+2LrgEdOw5wUvfQzVjbUPSD/VhHm3uckEKMD4ZhUT+B5jA31nSkLkf6
7foCgpWuPBqpNpK4PfcV00Yqmoc3WWeKXRPGFdbsP3VL5DIoDNLF1S3rvO9sk2uq
Ve9i6CR9DXVYPIzKhd3qLmsP9KXeSAgILyg+k9AjY0gZJzNCNt4uyS/HMSxZFbr+
KmLtPWmUg+Sj+Ofrh2T+C1wP8Nip80ZPb2sMQZcquqT9OXAhSjvnQCSwBcUZP1FA
ZiZXk5D2e6fqLwLo9hovIRMVlaE53aVFfuKXtaOixLPqyjZ90yqiNhZVa6jQD2de
B9gDgD5xvCrYQQAdzZd/V/VTK4JfGhPtgtVoC3wPTJiSkmLov3UeqcmFvDnigCRr
8uZ+9EEXJsDFLGuz1XgcQJoTtgGucXrQ3VQpxEOwFqbz/2V1bghEGxtjovsqgblH
aDkl+fc/twEUSpCzpGoJ8k9KLwWPrziVy1CKXN/afKMyKkQrNxz/rtOQD0O0RF2P
ZupkaLZMTfviMA16sWKIh0ABS9GqvbYhNBbbS8Uldb4eSVWAPSpCdy2xCAv+aeiQ
WIbgmfo0eYcTC+RX2BS6+E1WIrnPXnsioCx9RYlDYLZfJrUJVtJC5JA4ICht2Jwt
W9O5WyE8kwf+VUMhIyIPay24PGkPAcMH4CnjaGwaMJtbQ5BlcWH2GiZ6lJ2G2juM
jU0cMniSqH+ralKkTOgrPD4Jraq2/YQVeEgWkihzoSByA1ZexIsxuV3JCuuU1aDF
YZEu66IcAJRyT6C1d0c96BsF/PKMJ94cAuYQfcYEpDHCJyfKeygKopjtAG8IzHVp
0mR0iv8viB7AIEDNuFX33I/sqkPGZKvixgHfGzWKWUbJ7bxp5AYA+HTKGTV5YMJq
PUBquYJxNfrguSx6tq+uxGz5FG7h9F+XdyN0hTPX+GFXtdCVgDdpAFWe6uaNaEXY
jHCt+a1YniaejSmIXyNXUJw8NC85mSEHMq1XMouipukArJXuQuMs15cEWpA0QJWL
wZ1Rw4vEyQRKcr9Gf8BtPFSejG+BQLMdkh683+7oT5G5Ci83tpb7TTpuRF7Ia8yQ
R1iVbEH7rNPN9IiO83vv20WWn4jBI+FJWNHOskAWCH9DG+VVSR4U9pFbszuBXFB8
QfQWiN2fUxWjIrgAxPlYx60O6ffnsn/yA9FSE2sXwE7MxjPYbPBNkPSZ2q2cYqyi
1CxQYc58EAEAmsqEGmz1OfMkipMhPz6J4YtSrncM4pVS/3qqpKE3ljF7qbJqPyYS
W5WIL4NXaTKE5/Kk0QM/6lGU3vvQmDGJ6AfQeRodeujiShgfiNjOVqUFTh6Yxm6U
TMayMXEEzj0Y/UMa+L8ZtO/WHfKzvG39xS2KGA1kAOf75Ysk9dpoxFTdRo/CEb+u
zCacIzK0/FhzoWFj2A8+QcgS1vZw39oZGps3ElUQIAlpFz2fPuv0TRU/edxGKa43
btrKLAeDSkXcczcMnuNhlYUsp07duvMSqikZYY2XBdwpeJ9W3IbMH9H3TsBs6A5D
iRmu+Pz3A9f1YNhgZQUjOyGsXiDmyqjHfdCbBUhaRB2V9Gx8U2otPR5MRHqUqQAP
HMsXpdfaAIige7RC0baWjjkj3tLtXbka3BoBzMNbku0nWpUuwyjY5HZH8p8tSRsT
21ak+Qj0A5yEqEGOEBes48sY1Lv7DPbrjLMXAaGKF0+AxCjKqmlqxtHihNN97kYI
x/PQJULT2njXwJS82IyqdCzOpih8BWMRZM9uKUv36fblYWhHUZaU+zvfdoaOmwWN
FgpuKAu7f/oc4yDoNAYRq/tvNTYE112upZPRsTtw9ZU1euSqhMsWgef8w7D/tcvd
I/y0/6FfOFH/nYEXDlN4lijwc/cnoX74e1DcB46XGXUPdVGBTjKOPz8RDc+KnRsN
Tibl1xQGzz3OjZCMkV77CzrRbqlKVkznDNdvN6THHq31pm4BDQWKNGBi/FIfeUt+
vTrlE7AMrHOkq8kD0zYdouoROImDkcXLrCBg/leCFuGFnwxpladA3V2ofpjpAu7B
5O7lVMz0LbdiUseEzuut3KY2Bi5+3a/IVu7nij5x0MPm5eAoDTW0dNgdUu5QML9N
G+k9WLNt3gWqzdMroaUPPWdp3S+P/GDAerhj2fCcF9gulXkS51ylR96TK6+ufOS9
xx71wRwRod7MFAqRyudtxXVEVIciHeJ5AtyvSF/Ve9cK4DIQMUgBcy1HkYP6FoFa
NHnWqaCMaabsKNMxAKLe5Li+V6K3mvI4UTNb2IsOhBRhi+zVOev7cHBnKc/aYxLE
FIyihkrZhJgBDZ5vmTdLnm3ZGNRVF+fwLEDaD1WCGw9c/N5a9PbvhjhfJpTK9bhW
MELo+t/oMvGvaKRkS7UzGi2/Hqj3KpK/4/x1tYSlf9L0we5Ma68mt1i34SMCWfXs
eI1BSzAaFQPkCmdVMHNjGRyMyogYeTFAn0IKv7X4GL10t/I8U+P0FrgFsTwSs6OK
HKQvhDHuOTjk9KBo2eGSxlGLH9dMN6ayi+4UaDeczhUnsoYqTPF9Ye0/YT3m/VDT
5419QeCWe80s2KjVUeE1QUD+EeMb1ISkHCJ+tUxzY2tJ6qu2+//SC/9s/OtnLIMO
jM6smVr5f83d+T6cT/uIZ8oUYyJclbrE4nO90S9tG6aLddt4uBMcVsj15rpuM2ng
Ucj0cJHLfE5hNINWpTFBo4RXs0zDaV9BVQYnCkak8H1UwCU84X8nPOkMIFlMBf9A
bacNkQ4c/9F5dVK2/qwlYnZpbhEbzJP5q1eUtp86Ny1RItXlhqyAZ8+5hYbAOarY
aXdC2txhyAxj3mkmgs4gIY2fsXZ67JwUfMQDlfpOd2diYCSypplmwf62sp4NjSbx
LC+GO6UHxZirTw9uBa2uq5HUAf4rl4oXiRy97NGnLwY4qUQoludu0wY+FRowxFp3
E/Q8yJdkfE+y8A7VGK7XddlXT5702VZF2CpcEWui7gy/6TjT5jm4YfLdYe7Ys8m/
mi4jmgdptJ/Dn+usZwLSWH0aEsfb2Ezk9gK9eBU1n0hiw+j5SPJbAB1abRp4ulkO
ATRo19+WaDL+SZI9337c1inTBmPP3NY3mivLn3SUdROGDiFnGr/g+fpNagUz+tXq
Ev9wlrnZOdmli3q2v5Z0KP08wrs2SehrdIW8IS2lsoSqzUIAwd9kjyJIVPXiCgfr
k9DUQx/NVtuU4hpWrVChYbYi+UZs59UWeW4DMlPzkM1eydLCKIiwPkPpmUQwrTph
l4kpWq/cne66z1efUMwbW1J6NNC9rtmaX+OlXR1VHAhJmVovX5M1cgYoFhcrDO9Z
GbVEj9Sf7GB05HT2VVVvOcl1jjOwt//95IeD04s1NWTiziMjFUyl32+Meh5LWxXo
Jn74Ady1GNYpXj7p9JBuXZ6hRB5dm1eQ0V2ACIOo29DoXDawrZP2W4oGR2mzcboC
AhIhbfz5/9N2Y41zp+qg1CMKFwBDzLajlISZZoGPl9OCjt4B/ZJLNw9K9/mjSq5G
mexgIHpysc9DkEc0pL3Un8JhVcNH5IrPqxTPg6HPUCbGcBUkXVjss4I2n7LFdtJ6
Le364p/IA/zI5D10AiRzJ2JYm66e8MC60OjMKK/E5epKSka1+wm6NlOxICBIcqRr
IGUatTPvMWC5JldFHASUhy0b6ZXuji/Ru0vAwJudtJdpuL5cDwHgklNJgPSQooio
cL3DQ7TkCGQ2GxIjo6RQNLiJjJieHodbJPyk87XW1c7B0Dqcc/rHD64UivN2BtUJ
GsgbCEmIhzS6ATJ+aou+/fK6fYfbsoxZyVE7g6IEEiM93tml2dydlbImfAhs6mnG
hkIsywMVKoJ0Xw7bNM8fPoWW1sPlHAFENQ1dYoB173Xz7+gcWZ/FHX2DgitzqkvA
tTOyVboJHoPByZ9qDNJYX4/V/8nqxue8Pu/iHSFssEHwTaVUa0khPTqrbKV7/GAy
1NoL6UMmtvkGrz50FFzjC2p6ujckfudMcjWy9uZeUOw96f2FurJEZXSQUJ142W2S
E/B+7bIVeegcPVkl2wQnxC3XyPNKGon+bt42NerMs/qHqzu/MtzDHe8bECkCWHNX
W4s/J91hKjael0jnySNbGjhVUwnN4ZEbxL64zT+fFp1O0mcAW7iLmmLQl6yAsrbb
fPQlM56UF9zTvKGXXAUJpI6AexZ897O1EZCAl26GkaQ4CrBA2G3c/yE88M2R2kHk
KsviGRwavIWN+k7tV4T0nU+g6MdO5lWNFRShMb4UTIH7RApjL4LUaVAQTVF9Y+te
yYKs1YS57ymStn3e80urWPMy1r7W/rZsgEazAu9UCm5nSgS8KB7mJLoytWOpjGXK
PCfortScVLrHayf770brg4grCrw8JpfEBjBPzDaAAVHoNgw/utCNjGCIIaTWYUfG
35Im9l5m6ZB0J7CYNDmkHqQpeIRa7wMLP82lPAqdn8qOi5j/PsHrUBSpNoFfjFmp
9anzx3SoehiZrdu/9BPKuMrwuPkfYWgmOAJU6UcszCbT9H6SeaYrKA7JLTHhWHln
stPe0Nb4KU9yzOFEHqdWKCLYOuiL745DXw4mUqpwK2fY82379QBWWSp3bSXqRjvc
kuJ0Ldg1xRL71MRvjpzd82Olv1yDkuC29bU2PxVUVVmeYJF5N6Ld+k07uwUOZYXD
x+i4N9+ur37P9WJcPeHkipUpS6ogDjmVzg5H5VGLq1OzgH8Em60yeWyPKEMeeDhy
2veCQMfoUR8Y2HvK6xi/W0EhtCg9TJviADndtx/lp+RId4iz/hhxRDmMeDjdqahs
tpD6ztpfMJ4IMEMummPAzlhgzCEx6pJ3iEkhr7FhUdAbaV/xqDZZe6yqHm5IaUsP
TOln+v21z7fkdRBVy1Z/QLzvw9zpf3WLN5AstpcjxHgwNKrBo4SO7RPfV2Bd7sZW
3D9W0u/SI2XJPShlZModAgv7a3ChTzuZ6BvdJKgKFz8BswGIWKIfU8iZPj82EsGG
+GKc3k6Eb90mcBE6P1dgFar7fYd/l91XNXw4FbwbHXOzo30VqlabFoZo07JsD0d+
fHyJ/vbguYaiHr/kEpUMZekyZ+yi6pogQ4rNDOicv6OkNhQw+7Gn9l3POHh2gyJd
82RQ+vQrAg5rI+h00pLkRWJRSvuuwtM8KOVHSxc7cKSRHdXU1WWUZs62LkMO9RWJ
j09oIB6aSNcy5FiCKzjFTaPWXOI7hmTtuGQCIoBq6/tECtdgKI0lyXjU/EpAIJIl
Y2zSGD5iTcPn0R7tNR2CsPcKLSq3Cfx2BecNL7uUCMV4yMiwfWdsgQ9+zJ473h7/
bC/vzQqv1E/9xDb3v8tOtT+7F2cNAE6VhaYp9fp1pXmQ25krwB8C1XGV/shem7VN
pbh8Xfhsj7CYz6L+pL8/GKjutuzmrvOn5OROJd+nb5nk2SD7A9+PWVX3SbF8fR2Y
0OO/IT5p52x7hJKw8pu064D03h2qUrC5+4kO3ZTvLtdbSwLHlllNJZ0WcFQzAtjV
DVRwybFd7MK/kGmMaEnIj2z/yQJMedWEcutA47xcukzIU54pYxLxC8pcZjZCfVCS
P4LmcTpmvJztK+eQDkQScuIkslA++NUYByilMCjL6RCf/2yfVElq+C1sTLG3zfKb
iwxVANOzPBnI8XrWW8jdmZ+HJRr79ZKIeq2izKIEQeFA9aBgjONdi9ya1509WMWJ
l0CdNrw031/B36jbrkROGlPnIY7IsZNilI5Q21M/0ALTN06P+IBXjzWyOSFbqNAb
8tdGlLlbr2XE1qVWqwG5+BW6dq9K8i4xR02ylAFtCOWjoGjQgakKFdfM5xeIy5pL
vGKizorJfzmAYrh0F9ShUPhGrQX1+kfs+DGvnd46EvINyOnGC21aAcUrrqszaV4/
zOO7FRBonZ5yTQqlzi5JSpToBfWS47xnPPlkczkrHvU1H3eiVlp8alCLZs+w3Nxs
wJ1BV86ElytFirzu46EVymWeVIHcuUQ21XMLSAK496RBag2sqM2LBy1ZfHMit3vN
cFyQQhFfagRRHfVvfdJHyZmgtX8eZhaVfQOSWLRcdoUjtYmTgBkjK10dDHhq1aRb
3fmfV9PqmvV8lLT5ogQyVw8Z+nk0SvItbJttr+NlSulExQmylYrccuvQ5K4tSrFE
TigbVcB1boU4mJVRXf3ZEVgpc1O79gpwuTMO7jfCHZzmm0RL9gmcSAoo9faYt5Dy
BqNYFcj5kxk1SHkxCTe1G2/8PyvsRT0DvWn0wmh6omcTQm/hqRC3ixnq79dtaxim
Y0WzTf0iFBhFFRU7HAJeeOf/j4aalGNsKc0LfK7Y5U09IuI3s2htTh6CJAHEo7e9
831opxuVKkg5xEf3mb5a5vUhVMir5T5k5FMaGP5gM5AqgShwTqJnzD8SYd9gKo6f
iYKON41DiuQLTSc1TsU9WEgVeFI7paZ8iFuqCGOC0i9rCMkMLogG9sdrXk+aSh3u
7bAJd/enH86YgmBvIyi/DiCkMFIw5CMD/sCIY7DSVXmnjZD40xPicVLEJRCvZzHK
ldxmwXgs/1iOS5hQgFqNZ3GeevilvFek2J8Jq0MqQvc14quMdPWm1rbTdrUQHyVj
KHtVtkOCembrMuTI/wPNCp2FINwQ7tdGRQDJEgxvyWsvZIMrAApqYjuRTjMvD1fB
/xPF2+2/bK8sL//Euo9PEkGP9wWLuTmO/Z8iAwblih/pmgAx6SAzA94FFlM2NDO4
+By9hVHukbt9TM2hdj6Mn0vafnUw6qWCTAi+lEtoxCVQ4y6qKMBuRCKshx+4XvxX
3O/hcMxkDawtq92lKxI2toiQi5INs9DhdPDSFQ23iayO8FpWst/ii8Oqixc/jACO
mQg8RkTXZmNx03wG2StLgWjivLuLWZBHi2Ktae0wg3lm8ABgdIrI5ygLj0xYXmxl
DHMxRv7d2iGBYa0aq5S3jc/ZEPnUUkVG6TUeu9ySk10zW9Og7NCaJXhRbLbYilbX
bUtiTHLQuMaTIS1pouT2cXENBop5w5DPTAcK72BiVtq5R5dO3SJwkDKK74tRsSC5
L9xcEVOnRfMHZ23iAWb4/X1OkfH/G8vYY+R300vu8a+RS3wH/dvE0z1qWfAuJHU8
I66htV3fKSZpQ5008/7rpDKlFAgc+M9VHWMhU9mcotrC3WzFdeyaqmtAPNMU/xII
YWCjSs0FgL/rB6bhiXU3Fnvp+T9CzUzpKAe4MpF95QAwBn8duoM1eq5WgcGSXggP
un1D8C898oE3KSb4jKH7Ed3qQKenEOl8V+Do7Mgzqxuyv3n4nC6hfkXmUIXcukW2
6TMTVH6nQHHc6NYCgTloOiJ7UQIOebEFE2TT0IZP1GREFJ5CDMaUm/kqGRlH4avU
mx9wv6MPptvlZDoHprqT++4KuXTwEC/Ws5z6sffgWuY1cBe6NdZ9NQl1wCrS7a+M
6cs+0OwBBUqwoy8cSa0Eu43CxuXOR6ZSGzFV1XMZ3TdKFubhp8P9MpAUf3SUmsT2
Lu2QSFeDOneY2g0p3gMzjbE78usB8ZMnoI/J6r9HcWX8kjctSOC5MjsmhX4AA3FN
VLRa87TT/2dLnxqiAOHReoOhA2WVeLXJnfBQtb+OiFpFKCZZ47Lry6M5OHfJHr5m
3Klx8OXFyLT1dPo5GEAXA0Wk8XN8XejFZX/u3nfrqcHexid5RjIpZilIOmTemIrg
r/hov/9syetr6X7wPJu8QDeuX5HOPcvyQ/MZmtEk3ACj6MMiugrxl51YQAEM0zs3
gpWzrY0/M7hGci1kUamAJ1U5YlUke1WLxofJcypKUFjvPGI1Wm7Cy/i/8IT2NJQG
ejBsXkvHs5Vj0XsWBxv+Avef8LoEeckOLp6MkYyaydmYGdPwImpSGTkHMqJXMu5U
h04omWt0cI2g3suk19imZm90i9nc6D5aQzA9F5sucROx/OgNUAEE2UAUach8Y2lG
tsKYFzplgkmpACMdLFI2MGXSc7tP3gPI117D40NkheV/Q6CWeO022xCvhX31DP6l
hMNt0P9tgfxO6+w7ElUZOMGG5jfXNA0FiRQAl89ERTHs9L6f1SGRyQZjVjEFbQnZ
ZC6l3FvhhEpBQGxwlToNNXcV1Y8Wk9KuLoSqBhX/DWWiHEA4JcONlLjXYmMHonDo
kLCXGUDytgvG2mL0znmt9yDtY3AM5lk5ogK/+RWV8F0CZ3/pONXW4+ujP75qTXkd
eWAspMlVOE2+mlwJr2jOJMwVX0fxCDqxdSSebsZFFfZwn5lLC3dqxzGYsHl+R/+v
E3R0YVoacEbfOHtXz0vy8XE8so/m+Jb0xtsRmGBOmgGZVPneH6tDUrGvhD0dhwBj
/SMpcDTNeiaRkJ4suD4uo0FmdaesrNaeGgxNacDMqAdpj4Lt7ll+aHISg8smipO6
5yAQbVXgquXcsamvKrqeQRtC4CBX3dM8eDqp0dS/l6sw9oixfM17nCDu2/FWAQwN
g3DA/BrDjzvKiwSHsZmevNXRtJIy/AjCVA21t0nDDGyeYNmDC9c7KQjslpViqAlp
tls5Si/TkRnSrs9+F7b3/6TlZjDXF8pPASmzW3fUzvakLXlAL4V74/RSxQfWJ5KG
fcq+zHo8cceuwlgAxhHL8UBitBAXjfmitOnN1YiU4jD7NZtlXQI3T8Tp01Gelt4A
6fgDHFmrvJoPW+Fnro5KrUYiKc5k7AX0rMoot39XtDnjbNUmyfC/eixJJHm1JF+s
jm9y6yRwCljTL1R35uHqISgN+xgrYgGfVufh1h/een+OlzQfBI/zs4Od18ehcxBg
OU7myBxiNnYsefI6j9k31BzFW/VD6ygmE1hW1kEWyjGlgJD10dEoOQIsxeyKgRkI
hhzpMarcbUFSXsWTi7sG/aBQhmS+TKyyy1o4YPaLP1ZSrGfdtEWtvw3qRO7xH/2x
5xYFb6VjXKHJeKZmp5jvwC6STp1yW4xTfyDd/XEPusW8Dr+6Bt3O18dy63MDAuVo
zl5sMCQsqQeLipP2AOPOX5jgAon8RjyRDC1UqEsrUD+6FVSeBCRmaAgD4MkYCnMq
PjKxfb6mKllTLcdOKPm26P+lScKQH4Mr7YOu5vzSzcgrRWIIqFbi1vG5QK+SzYZT
Lrsi33oHv1R/du1uUrVnb1Ucp1BaZUPI97GNgqz6+/yBUggkyY1QdB96ZytmrCRC
8ry27GNeV11KB5VcRHXQImK2nPm1QgDC8DOr90eIwvdC2MRmPQTaKvxxqCRDMXjX
gQCPADbwgwLPTQTe+naWNHN3UKArddMnYpfmmmIlUlAy2Rr+jwQnm13NplZS+NiO
mwnPXkIn/yvWFWUCig+q4Q0ni5jvwIbkDdB7FzNK850lbadNZKuLYCuJRruDl+Hr
pEF+sIPSW6dyzsetYq1233IPAkSGm7bzfUqmTJ6bDl+7V6yDOWjAj1858sG6rowp
f5V/jHx2/PcaGsQxcXEglioVA5q9quxhrcrBc4OBtjJvOJxT5PMgr2X6cWiXLrhC
QA/8Yq6AsS2c5z67vTzv0iqa2xaTQ/INIAndvKb6EB0wdTDju+deZcCtQ9F8MVHO
wStAi5N94P1bHDaw5SdnvM6Pto8sdFAsiVWuRTquWPQCd/KmxzKK/hTs0BhiQkxM
G4Sa/+MSjFTgL2NBUevOWQYoMWCjFabKZd0PjLKNckqaRdGuX3R3sVjOvEPUKyg3
b0C5gixlmRdrQ2h4Qg8OUSH/FbfWF+K6xANBvwTcSFXZy9xRFMw/y3YF49uCpePL
y2kR5KxXuFjY2XfQAJ2ri4Or68X8wWbWMgoArMG0npi2lOdkRalLtrrLI4h2jd6X
SOyhuBhzEvsIsox5+IffGrdoqGrEDkuZM3GrFlfqTBAk9HagCXvnLiOj9EmmAnvj
Q8e515++6OUgwzbgilz5Ca0O/bcj8gioNTOHonEcGcX6ze9fZEjGXrtwmqgesqi4
lmNtPJqpNHXxuPAeqJIV1pfTVkbakhU8mKpTH4d7eswbCcCcf1AGMdiCBVhL9ptI
ftrBrcWNm6/qrI7GVNT6/HUNkWda6HtYtGilXDDYFLw4xCcN0taSYHLFRDoH7OM6
4Gti1vMdl86jM/CAnYp3JEawOtdEZdnCsEXsS+PNXTJ43cYcuqjFewTG3436lkQI
3w5htY1SlWKhr2JH8UvGp2ViXfvFUAeAKbsMJihM85GNETypXeFTcwFaivPCn3JX
CWVhjXc7Cubuv5kM/1AKSSGrOIkqJUxpdRhhp7QsZVuKj2mkHIzEM/GjP6MXX2qO
iWHIRs0fpRn61YBucpCHFjmfZPD0NRvhXxbOgpSRRoxx+aSaJT2uG9yqWaQgP85H
X3VBmOEOVZ71maosmUK1bxk+mXX2gMhghTWsrHXt0auVCKKknVGrWjROWIWGIZez
MHsCLOn5HNo7DxT+6h4E8OwWiThcvdoecENRZ95qQMBgFoOKqc9hyxA5SmMs4dZ6
utpaYNtsvrLiUAzb9gqV4yQIE3BKmEKLjHUBzDjZYfxzcx6BxUAqNQCtoCOJvH3F
zXw91gNSMIqkn0pAyTaShlVj/BbXOHanUMmvhV0VcaQIWiSuzi16oJCwuI3GfQog
Oop3YVk5mSZixfv+7wZggpqSnjH/nfYJUJTIr2JGB2yGDn+F2djbmCwVSHYAQar9
WVjnfJpxz9/YLTjw4TZBi2ZE+C2dJcMF58jZUSdvILXW8W5hNAr9ZQmY9ZX5oDuc
JsbjLvGXn3QmLyljM9Ml+cGYnxnr0sYxoQ73OKyHfFrbg5M2SlMEAmNJ9LaEBfg0
baCjjSNdRxO1UJBh3tlcGcgDL2G7IGEEQxRlEgpsoqIZwEUZnT7Fg/cSR0F76LzQ
eMygJAa2uQnJrEGT3VH+Ytjo5IPuGRtNpIk54CSkqP7nOBeWrDjUsumLzlyBaNZB
CBzxCdAlOQ5rqb0NkGfngoc7Lwm66NO3dCSorcBnpzkDCncgvqmQ+sYLzEFGCdbK
OxqTDz8R88PKYx+iSi90AErlyAezyu5cw9e3UDuOBA/1/QABJwtSC71a2Mwn/UVX
LFxIOl90ywL/LrXIFq4x5PCrHNXGPSsJPQcCJ49pt5nBtr/4CNwNrxZ0Uyw1Vx3v
10H8Iu7mRIAc7h8/thEjHoDnNnt3jZfcCvlQ2OZ7fXbET3hn5etYnI+4zFJu3u3O
1e8VbeZUjGX2BLZju2gStzWN8UF+TWP2rRb92ZJVHjhYoJ/jMeyN2h0bQxEjCQF/
F44B38pQ/LKMI5Z5xGOtDOR/vRnWwLlLMIRBIocqsslZbJ7DVP5iqFO2t9Vr1Btj
ZUSR3o/0BdF/bI7EJrpwKHL08ljR5Fn7/KT8uA5H2k7/aDIu1UnLrHQK+pt3aY/P
npucE9P7g9vN5E3hd8u50nPhK+IYtNwCABcniQ9N1CAC/m6Jycwg9fyJURKgGuTV
KGuAO88CJIHCAB4OSWwtk53yysDuklfUbFpUQCjRhLqfGykVfAxaNwiRr3o/rYus
bUTKEMXnO8EX5AgfO655xvjjr3xitgS01GlXlkQpBXWKVAKFMtgqTM7bHTYLimRa
EJz4G2V4btOzCM7zgN1uxcXZGb+D52zXUX4S1fOHstsQsbb1BUqNS5/hmrsppD3z
H1lDBcT7Zd8LGtguj0Izf17qg3CMWrBYghPIzgmrElVQaimz9l9+5AHKTUV1cDdi
33GirlftKXTzYKdyOSkPam4hHGI1ZPHnjecdeLFJE5YA4+rfdFkU702QLXlS1Heu
UqVs5Xt7NNULouDAohpWiWZymjdZQW4PtaM6WqZr5FuTmmAM3XgdiIzUpC1LxdC4
qwb+2SGD7Nsvn9hjJvEQn8MZVSotdr/eA5Q0XyKKlmd4x7VB5QKslFV19Xt+ls05
xUDUJDiiZnKk1zoq1OvCTnnIa/0vGwb5mHki0P+jBwy5e/KKlgU5didt4MZZX5Us
n/G6D8sZzQC7M9cpAj4b+gJYSaUe/dIKwNi/iMlnM1FOn8SSh9/v9WJWti5kPTRc
MFZmghXrX96tBPhNIIS5kuHxiwt6y4lIt7QpBnCVcq8PMeq6DY/zHQFixAuzxlzF
PhDpz6ftdXosSEXTOBVnn5XycPZXlkRCsb4vPYK3KK2uJjXZRyVqHS3xxgxT2NlK
UCagRR4GFvGTqV3HTCU2K9Lc989MK88gHVD2GjIbfhO6DOiceaQ202kS98Tnp71P
yANFJ5OmSy35jWOaLvS1xPUDe7KLdDSS7qh5YQ0uxiENXB9xGkSQ97h9gdVOf/GD
P58ah2Z7Ync7mqjHwYoNhwJOHe9AWBoDCF+D/1UC8CZUyIy5V8nU0CYpatDML49C
et/oSjDIyTjOV4s5TSu1gp9TsN8FPIM/AHY9U133M7sNLWsqfXH5no4xUupwH5eq
rldd+/52XqVPnWauLAbtYeSK8jSVwmMMjqb9vNPDiFHxujsp/DFReE+dqms8cKNO
F3fmygo0Tr92Pi8KgO8tuH6zC780JZjJNDXyOEPCDGNzEJ82ZAeft3i/jQ4A+JBJ
wB+oGW4ZtzMidfgOR4TUsEBLMKmby8Y1EBbTGitZuZnOpuCF+2fyuupd+lZe8On8
UsCOyJjVygOt1EMNHGPrE+ZhTAoP5pkUYWvgws0yvALYSwXULul7sy/bhulKobN6
xFkEkuFj+PMe+jNVSPdaczplgHb09hny8AQAQzAtfqKZFwotIvmUifKWaYNEBwKm
NZ/JxQx/pe5MCVTjZWAzO8bxeZyDcjf7laeBxSI7TFPJztSRtVkdcjuWopL/rVcd
xsCTyQE7VvpoW0Z4Je81p/fGH20wFG46wU+/5HjLj7dhDicYwI59UCynGGfQ2Cic
Ft3/dobi46r6Os2VgsgDgZKgcQIlFSsd/8j5QJUbezL6MZ0EKDB7deKSe3OQjL2i
7Up93Ct443iNvqlK155yz1R/8AnhY/su9+cPfNF+WSJXkpLXgi+s2M55vXV/bDfC
lp5q7bAUnahKn1t7RLcMWwSpBykDWWpFg4cUJU86BN1f3mUOxPsusd1Ev8TFZIp+
RRMM4BRAW0JG8UJZF3Tq+6F+upk4imyTS3Z50wuDtdhnqQB9FJZGYFAvRCJYPwF2
rIJIogXyn5HH0+9XPn9y5j3c//pMxWLDULFLxaYbH5TKUOT4SpK2uN6iVIG++ohu
lv7BrmzjMMxx2WI1qa8eTTEzPbZFru/nphWPwQqvyBSSYVys88zNqUrJFx7YQsTC
xhiT+fAka7qlMqPKYE1RylmfzH2O8DyDoWOnIQfqipKYZ6WZVqVUO0VjIbtY5f1Q
RA+rjKwblqELhJgj2erMBfIh0WLroTCVfSA8c8u4PZeXGsC/4cDVYzs4GptQnPjn
1TnWXmiNV+RL2KE41CBaj4SjjcaC5kF1va7H+f160V4GymIj/sjlNHaLPlMnchCu
eGu8Fzn4G78yff27EvU6WGOsbDLcrbnbWrDKqo/dtnKPCABVdHp8Dw+0kHNvTD8r
1Mpil3pygnBYVPtYvm6C5yAukzae8YXValLzvc8QTQvFeIszpcc7JdeNrXxkyNan
EHTK0FuJG8zfRvUt5MQFIbbh+Mu7rAA/nZcpmJPK23TvN/xy2cQi/KydnCLXq7oh
kH08Um7UTnYwRaqrvRyC288Q0x70UBZgMdfMf7gKKGaPenZIUipOAZ8fdDotzjHe
eYy5F5Wjx07CjYSRujoLII94B+N8IxAwtlbBMhC2m0hfAfj3b1PY3GYnETM/SgW2
mM/WguF21uwphpNR1yTLhAVgYjUEyCZ41NUCVLeBK7xuwGW2+7Eqbo5zWnxeJWJd
hYqOwjGEhAnBXocCqDmgabWvtqSdzdydfbY41k1jt/1PP4CxW2lLWAcGhuEoltYb
txv14jqsZx2nyv03nQWSAhGyShQE1xQ1+gZrbuYSnJNqZkyQcF+2hgkSYUKldN8o
47HNEeiB/5shvPu5elyGnmDyeEnzw/2B/nf7eR7AHqqfxnN64srfGPO1fWe6CnF6
r/kNbPf4XSLQM8tvsMpMzDO5Pn/kei8W02ea6hYYijTXJKvMnIlb6HxOKpezBqqk
jBLKwl0zVewMB6lai/8QW4KnBUdqfV99w2hxYYNQxFy3oDfkJbwQMSlrob5xXxuK
4Ln8pUEmKoDi4QVDQLu7hA4kwCbN+08VRMYBt9YBRe4HRQ+XO9sf1aNAJuCBMcLZ
ZCbEyap9HKz3rUobFlTgqja59HOmUISjpXAHh8n79llzu22BNfRl5SZE1dyRt6jY
i7HbTlxVk86yBly1fHaqgHR4jh/eON6C4henw4s7HWWfpUl6qT0u4nV759UXDagL
xP/hUHSqxNyX2L6t+EY5CNW7M78G9ITZEqwi6VX4m4tT4A7WlIvdY/psdgALj4Z7
oQOdcFH54UC//ip/VUMFI5xvOyxg56QBAHXkwCx1slgA9t9wMKzmnClf9hFpvpXg
K9R7iiOUig31C9li2ILnqK9q11FWRx6Xsp5zM0iC0r/v2iwBEU4/O5VUHjXsBqlx
rsKc+L2uaTJFED9ouysDUW7f7ONs82AzgxW2UIl2qS2zmkKhNob7XLuR5nF1w9NO
I6UKFfJBzma3DmPx5fNjbBFGnFonq24WvUPgF1ObVDpb3E4yDskKjlERofFvIfHn
wtjpWQDnKS/hj/bS5+fcvHJ7EOHsdiItCpTLq/6cSxv6wW/HAOExtExRWnQqnGjc
+0xuh0ISaCzzE7xSI19DyplmDk4ltAMs9vNiT3JAJrGyqljM3ROaLijrcj3W/VNg
hLJbDXTPsXrLP3Bixg58MIvfUAy7Tq98O2nV7gPR45sa3E27/SYto8/w78z5ssBl
+WIJgsOUOteDSBZV52a8L381omEy+WXt8oh1nRlPoR6irRnO+683r0u4bF+fejIS
A3DC/+39Y/94fu0DIa5OrhmqyH8yKuXur6DvhTFMLY/XnNSgRx5UyDq1E8TxRd9e
5cEFO63zjoEvA3mggk+13IxqsilEnC8kvwgd63kZKerNMDxKFnGT540gm+U/ug4w
pI4gQ0plvZW/RIm1nmku/ImSMGPZeNmUv3mZW/xFgKVNiheTkGR2DuPzDhhI68bb
hP2yu+dCBTndpa/8dPshmnGogl3HcpoMkumHWW7Mnp9GJsoIUY6M91bABNZ7BpYo
HR8AB4FpO9VwvWDHbPvJOkd3oPZf75+PeiuwuiAIu/rttkaNJ7IP/XJdLL2kFhnP
PI+GxypDNxkhVSHdGY73I4rbueWVSLL9nJ/ybItyleJFM1iurOpgGb6IWbaqDyuN
iAd6ODTOoSvcVo4DiUEI0Cav3KYVMSCd3d2VcBRHwAeJb80XAGL2JBAlly/CyihW
e/sFJ8W+SW3zv4ubeS5uvuygaeZnUf4oI8zcr/fygZbvsPKfnkPg1rla0Nw6icSb
GfZ/HsQ8LSE4/w1AiXO58GWXlkfyoDWTAIpjFc8g5foeCi5IJ3PzHPp+rUXwZrJ5
bEk6iK4I96BH1zhWTDewYOTBdWRgJOvBIoTW024VqnmKeRUtrvb7ypvJT0bIUnKj
4fZwlZ7wKXD1HV23upuAMXoyQwomDhZVqgmDmOKlUrL0LVlJP/w7BmJNVuZ6NaQW
7Sd5gpZhC0m0iUs1aJ5S1qTkE/X82O0Z0mtOCMmtzAlovEP3KEN7DicGfMDXHsld
4u2p1oc9rwydPBpQsngawtLypZX0RoG0PZCm4SyVJsyY55UNFLZjiH86CJwfKtZ+
A4zZe5SUZNqKxmZC/0eRtrrySM8LlpiCg7LS1cdzMhs1TRnyEIdxYVeZphvICSii
+V4rjAZGZYibFYG5HJUV3sti7/iMwqvMdq8R53ybM4x4lkL2r1xzgxlkXsU6QkV+
RnJiCp2VOWEyrXjpo0oeJLMCdvy5IHNyV3cn4SoIVw0rcpNdcd069nbONx/cAdB0
zofctpYbT+pL1YvzaCc2HKwMke/X1kWK68pJRjf5HQbTaxqMgSHVggNKEPFHGdu/
CPH+ZqS1nFJBiAw5hbqTkl94iFws+LRJYZGp0xEMo/wYIRcTumVj6rUtcNiR3Gk6
SqRGH2whp0Ipp/TFD6mkkIYyVgSVlQWANgff3nIkHNF30KN4X9/EEdCmJiFeqcgz
qO88lIlovCBHWmoPTJKprzG+5R/ZscxEj+jk0xf6YY6/MqpudaEjKsgeb+I8mIUB
xqQ/iGPJmzvhZtN4tWLgiDDANSg4TrlbCnb0rYmKIeXzPlGBloTrrHZ4yo5nxPPu
7mQI3qymimnM9fg9aGv3TNqhG4mF1aIh3PWmgZFYO6jUQmoHwU7C/zghuC/K6AwF
cYCDYlDXGkFuTQoqY+CWnOyy/P5PMUrKBb6F7RA3A6UsNHqJZfVJWUZPmnJD6Jpc
2DDdwtBnB73DuzIJ/K9mZ3Sg0kQjxP09pvDprDMNQjZK+90m8qA+jKhqbCdMmmYT
kx6YzusJiHRFP0WxS2gKjwXKN4hr7jLgLDcAkHQLwvI6PSb7Ld62nvCaFwr6FFYE
B+FO7hwhRPLqPKeem6Z45pd2RVjqS+kdCN/8C7F+r/u/qIXtJs1p+58tB1B47SSj
vpUyMZ8CmxsA5jHlFpauXVLsLEpptL24jJYXNAgjcgV6gF9yPbMaixIoEpz2c3N4
T3tQh8mxsUtehUP8yroK02dBdWn9gibPAi23uFqNEw+9dZd27gUs6VAXay6s7uMf
50TgP52HzAaJzFbDSRHt9NhXfpJLQ1XZE+qHElg4D4yNQ9DDs+F7+CZ5zWk0IU1b
Yp0eOKhjc+H8fkjpnLRqKVje0rRyuOe/m0CU3+Ao6pl0mJHqyRtYmuwrAEFuwAfC
okRk0CiQlNicYIy5dDGNT4iSz84demTnWy/RhMU0swonMM8p+l2SngKXg9zOeqfM
Kk7NNWi0QdEp6q3szlJ6LA9gan/pWAjMbkOsQMxwuei7aPSRUza5eSSsSdVfo3Is
1Ii5UVc72uonSyERp0atyB/Svg8FWQn9P8Ah1cDQyq434j1RWI9IClO/Yw8JdwV3
oz0IrtQpE0ESBoP6a+bemi27QbjloXxtbUMRjqT+F9tbcB2l7Jg/wsVgH2SOKUIZ
21j83YaVQBGx6H9S5PSGl8+E80ngVJsRw/QpqcYTOH/rFnjMcCEFxf8JW2+P5WOi
UYDMx4k58c5C2zssX8n3DOD6ay1ZBffayuOjYiqva8wbmveJkG2122aSzSwhFCmq
pg8ZpL+mn0PYGncuJDi2MSdIGFNTwrocazJoCu26shdyWWF24WFwuCdcnQrIUHfU
d2UwZVcTDw3g7/oAGazpVrjfxQ9i3V0YPVKCouMpfWqaZtd4FVMP5I/Ks+E4O//Q
oWQgVyqkEDmIZR9/f3ePThU2RUtvS/v6bAc/I7kslGmvKpfjn4AN4eQbMUvwKCGc
ftYRNlZaL3nzjfBovBoUIkWLA+QRjjo5Dw5pzYVmnaHOo6uW2IYTsG3UldRsMSwv
Mpra1A6220HToE+BJQ+YPysxwzL6Fw1+Ws79TE/GEGW6C6CeYA5RDcH14GEiKob3
CXSvQxgkigGkG/cRRAjwu35UA95XqUHDDP3HonO5iKoMqLBKoAKuWOAuU18ybJmS
22thgFkOGI1ugaHKtYp2xeDAUCjsOI2IGQpiqvJP8k9D2J/tIKF13c/VrFsR2Sza
ZD/SGMWDq0MWgNIKaaUHZUkyIhcSFOaiCdyXz+yipdqVXn8bLh8N/zjyF5kumRre
OeKm6z67a/2lWz2+GNHfgz/YCi1HVUuOuVOBQ5SOVGkraxRI75ewFCiv0j7EnCXn
B4kute25DdP9/wiJq/5pq0opBT6K5MDP4cD86yZUiOuL+lxkFcgriwcAzcclVgas
v9zo31MyBmQrBYt4/SuPsBV+jeHNIjLsbLWKutSXj1KKsXZZvcn+r7O74mTTqK7y
4q7SK3swzzYR88rUipoWPAGx8knalMx3HnQ0mPkX+kUQmxkWFD3wAZw7p57+8Li6
Q9CGAiGU33EUwH09mJ7GiD+HZuJKYWKOUjNKNTBBXgcKzrGM1LH8o/OfKAxn/Y0H
tQOcZ1eo8yKo8BNym/NGfE1RYQ9CJYoULj6iCSHLciKYOCiYFXSzQJgnMFVvkt2J
VaCiEIlqOGQUYqp7oTtjNckEbGf8CyMaQBWmf4tpAMGtzxcI/F4ApFpqyuVymlxD
5fZjHoNa/ykmpfe76jIsgtRcwwm73JmTiq+vLaCFyq6Y6UcPaaPYYio/MPw18Tp4
sxhUIEPju/k1p2VcQhcipyLOkX92epWg+Xt8TGqWusxFc1aheK0ViyXItpDxCYEY
QjOF6CKWJHo44QMWJMr8p/su8XDVU4dbg6IHGgxAKsM62c3jbSoyhWQvIoJknqpS
hQdnZQgmFVsro5zxJTZ0mUoB+Y0iihabRls9EVsPPoxUlCzQoPze2A0HZ2E8w8Dg
v/jwgQQl2p7nAsxwNKTzgrCij0PaJuKgmDkhtY77//pY+EUt0gciUwBYs7YrpXj2
/OFsZPoc/0xD16+7Xy+rnbwxmzFV7sWaQWbfULNGZSZm5ZdVINlIMqy9/DqKnRKp
BFgUqjCYUYV1GRngzi5vqdzU0tsLgVEyzXREAf67pQZf6wulxfvoxxeGjWUUtcjz
f6nna2Rp2hs25jGcELAt0h6curhOfhwur8TB1nWEKY4Y6g1TNBksRurwFhcmIb8q
CcTHkGLitif0deGsYGW0BrTqtjvNuaZGTU3je0SF0iwDTSbhA4o+QLDSvgRcEGJL
ud3wUqTowMYdjAcdJdqU5A6DFXpc2WSgCw8lYhhGpRpbiTxzo8N5MGLwrC0X2chN
HAARHY2EebtVLxT8DiuYetErbKbEqv/6LPA/gkfaah7+J0xhFC+gkw4WQ7zYCi9Q
Y44n4TGbMDonj6Ux3dQwp/skm/qfhsnQLPnlCoP5zFSyo7Gn6g7bR70HZIYwG4wY
xgbd1AtCmDORgA3QgjWYnNsK4lenADNrT6eD2wXbyqH/ys6xNHJ3h3kB+Fu83S2o
UbLCC99fUT8whLlZWpM10v6LCU3hk3AGs32usU5TLh1X699FMbdyeUcGd69jj/PM
LERjP3HgVR8A1M9vM04x5vWmUwX312RzO+8HisiteAXuiPdz3/HymyS4Jhtxsbl1
ymMkW59DG1oXe/nJWpN+8GmPLWBnkUCcJNxhND+x0NCXwGERQkbi9ipHmXo4BLAg
/KmqzyWGnl/L+syJ1R/xkfVHoKCfn/04YbCY47740g2UidWoIA0kUtE9K9Yes3nN
j6FgEVJ8uTYCjYgaH1QtojPMzwCmpY1MrPLZKk0XdtJiybuIHLB70dnvscuYU8UV
1trxqYFPvUEXHER/Z6B29S0+AwlgTG1PVLDTXx5BY2NsbrDeIPwUWa3C+Lijynmk
OxWfWPyr4hGQJU8oCfbruYuuYkw6nvgta+51D7XIkzpoOyw/tYkW5TU5Cd42bBhg
dspH6UK1OJBvV3nsQxdu/PhQzrJNzZKjhkKXnW/D8Aw86G+W943umWR12YH7u+Mc
Sf2UVEpEmdyqk+59m0MXD3o9STaqwXUGDVX1Bw82Nivb0qwDdBZ47PuvDbVf8PgN
GiBiNI82e6xZjnFH3Ane5b3VmpC0ecayXPS2PbbQV24JYvQHaf7DKJBbYjOxvPpu
ryMi1OxeWLrupmXK4ZBCtdmCztu+ExSYcaISq1UIAhTbozSCbx+L6O1mePU5/1uF
Tfa4MdVD2zIZy0FkkiOVhyQb1w4+pvlX1L1gGV5Bb9mQ1O0wYu5ocRO5w/fkB2x0
QwpS6Yjyq4SXpl6xqA24mgFms7bll156gCUmMVyYfIjlM3GHkz8iHL9b3mKa3QNA
UhqkmHaBYPE+XrDrvsvOHwvchGdbPEpMpVg+t+wBE0H6fvNic5JJrLS2xV9lMcbj
bs00SPfMKi9faf5N+GO3Tn9A9rtlcecjUIZqCaeZ4Fw7ZDi0A0gPwdhI938bDk4/
drPCzsKJIc8VCmf6goQi6zkedLc/3gZdvoZQDskV8o0MOr/1/ljdQTm0fENb7B7b
FkeHZMbTpTaMk+dvA6HS7oslQrlkxbCGsua+hz84WT9Q1jhZLwvR1bIgV1QSq6Y5
J+7SwnJZpIgTnqTOVi2CGwhBi9ty7T0JYPBgC+c3Dtgyc/A+mW4zva1dDwxy+3qt
YSyDpuZhi+RpVAEJ7xEAtF92+QmT4yqXIm0Z6as0tn6cHOm5fAameNPTHsaiKyWr
1vkrflxDyy0H/KOquHYrpOw9YfEKYaFXD68g99+DM8KalEb8nX6R48MhSVBP990o
7O1FJFvAkf2AGoC9c/OmVmeMuz1OgdfbC89SbrIvYyNj0Q+sTFUQx+8qDh3Sf1pY
VPT7SP+QvuTDzD41oOyywFKRRiy6V1a2W0eoeoJIbACmfR7JAynXK6f1nrivMhq/
bcr2M+FSydmS13630+WDPQECuNFhgOGDb9/7/1N22SQGswBXXS5btQ5AgyaHDJT4
5FRX/V9HkwZk8RBIpNU9E4rzYKng0joxYQAombJOrLkj4mM45n4EEI7wfc1tCek2
R7l0ne3uCn38rBV/oSHMLP7PsPeU1e+wNLDu735IS/uXr0sa/SLXNRaH0cAYJVHU
lc7b44UQNumX2tmIBNJlY09VTXa/OKdxIBhevljrWDmwLPxE3HHf7Z96yxVBDn0+
zPvXnBunF1eMSNMLAhe5UNGRUbdC14Kmj93iia6pnQLwouBF9vnIMXrl7mltnCo2
Vov7fRfm5p/yaneZElLnhJSpChmS2Ws2zFa7v81rloJuChAtbCabEgnWnm9/c+s5
3RlYBfTaCLVQgo2s+aO+348IeovTT+SZRUJMiF6k0c4lm+0sN2Jt4P5snMnSF1z4
Dk0xK2qFWgWkjD2swMbzg5+B20/xyJYlTzn39MT26XLoyBWdo2rldOcGoi8fDPVa
uyhzlJrNtHjtvcsBAphNj18Zji5G0kUMCpGzqZrsTDOI3Xvpdk2RSR/Y0m/2LTla
eJx4p/IWDdcoDTxoRhS7xeG9kCJGzOpLYHA6jeNPDEDxYamB0tBD0CqSbd3nMbt6
5rAJBZGE8G4Mmm44ZnkdTNJDBjcoTAAbOUydQ4faTu03mk2Rup/j5toJNcj6rt0o
ksGL76giSZj1HjrZ/Ab9gjk+csyqqo6N/0frAcI9HktHTmoiDncLIlZhIwqf0JDI
+XaQqXVbBCgddLl2qBw6srAZWmv5edrXt2AxbLI3fJqVU6diAcOv4gyrg0jJ3PEr
na7L00xCYhLByCiYJhWIRs8Ja8cH4CgbTFaKqwh9Jd7uEWKYAuOACC+XRB0OAeu6
8NAbE6iXd4NqTACBwwSvbyQanc6Rj96cAbZDSinpvxGXfyfu4K9jezaCmIoNZrBH
VEZLebTtsnc6sidFu9nj4CPJbNyaR91acgbovKN+FZP841gLPIbVx9bxBe99zHSC
xeVQagg6ExyMzMwmZ58bsuoKs9rzPpfqqHtF3yO3YxCPWnj47L4GXh/5T9MFphXw
Xh/UCFuRVBSRzxjDH1WKUU2wG3ofSWflYDO792GqOcXaPsBkmktie8baTWiYbLPd
aeY3IGx5ywfuuiBW6YsS/m28gqT7KChE9weaY8Y1Fb1JOOCQzICagjq2alKfAL6G
rsNyjMQWvEDpT6wz5lXb1cfQWknm1N/UhlFElY/jH3B1iEMF3RydWTDLoi3m5zcT
2skTAk0cQyC9hqrEJE0itVKA0oGY+AgUuXvWA7kXr4dgObd2AlX1fpkT7jYMzCe/
zBaxGAtYOyKA0dnpGgYXK7/yOe32X4HUH2GbETfTMduBQXs5+cN/glzybJiImRLq
1kK5qADTHSuNf9rLJUC0CuHkYRa+bLawEdYEvMuiJqtzGL/ivwM2l0iOxPK5Cv1U
Od4r/AGTSyeeadBN8bPKg2YXp4fj0hpQQP5V4S9G+xCf6BoXbD3YUKMDafoN9JPu
ovJp64qSOPsLOtcyI0EEejPf4rCuPxkNlgxrjjyUMXPyFehu7ffd1m1odM2WQaxB
xTlRp3EPM1sNCtt53RRAnCqu+rskUYCcqKohEAunOvvoaYenp6qL+b9WE3t5EzdI
qFa9Lmg+gYybn5foBmE77V/aDJS8igkV3SVeIIefKIyMpdWlph40WIH+z4tKKU1N
R28cz16lzxcMkRrzUcxc4trdBNtwrxxBOg9+nnryHB8TQz6HKj20sbcoCTZdRyzw
0B2pKJ4Ockn2DScH8wvv0NkdDMCx8E18qxej/lQ9PeOFEQwqd17/31Il1stI2emu
9FyI5FwKhuvRjkO1t7DfCx5S+UQoL+qCzZVBmOaqvcWMI3mFkLLV3J+p+yVa/tdI
LaC+fk3xQhbvMdDTZ3DJWTHy2GqhS7N2M/nwVaaHraLYGC3cT6dRqInA4+bon5RC
24VPNrc2Z1XYljs2YCKJFoSN4VIsxCLDQXPvzEWkXM/npwDCWSc9e3gcuWHoHp+3
jkl/II/EPHN/n1fBqU0Tk1o8oc2dmSFqSGAgkCg0PgzoFliPJVAXMTRILe1aCHuf
iFtI+rJAym54AVklNznmsunff0IKHhr++7mWT8hnnXFNUcquNfrJjTTMGwOUgVhp
lO1/vNvnwciDfRjitehde8eliJhYv+egYjc9Nqpv/xkBXDzpCsYiHZfBivexOt52
CdXXRGPU0qPDwmh1zKbPvFXBaeSTqoLgU6/u5eujH5eZSxY8URyt5d0oSRe9/ItG
Pe3sBfE5AZkKlfzmBd7Hudy9Kr7fCru1SFKrRNY8BY8YkdslJN5jFxfwsux+5trT
te9aSpWFyj/dhwbnTaihf0ushIDoAmMoXzdGwsBOM9vy20M37eHjOLMZIxPfdK0b
HBPj+zCZZfmgCP0UbCX7iFy60gTN7jURggqvqRkiT2nrYbwDdT8iK5fOoyg+1uTN
jorJS8BoRBblSh2FwbuKAciu0GW4CfUclqD3LXIvsisJ4jqKkSb89WVDWa1CpKT7
fXMMwO1Q2PZjRKy+sIBLhNmsWiQMs41QOxkFNGxb3sRdSgNqXVdV75MCWPrUcwFc
2xJafDb/tBmeRqi2/Qd/qUGoKxF+HZDSNpsmkkDyUpmh2XJpEkmsAIfsMXbaDLad
RBiQepsm0uvO2XUYhLWFKTTdYyhmSje1t/JJpqAtjgc2SjQU8ngempSZYp6+XcGH
ktrAoZtIQBGusvvYkyOXh3nLma46hYfQ/Sjf9FaxvlJ4Vg/RVqJ033985dBc3/jM
NpwocowVD32MBTErb/Y0vfzvbk1+5PBLNnGkGi9D0r7BZamGsNDAQlBmtmL3d5n2
X+tLjqFXxKuFD8pxgzzL8ZFtcBxJ5Y5KGImDCXuswlWthBackoe0sCH6scPJAL76
AbtalN73mvAoShA4afWyk45aglNJ4N4TqKlK0t8laeEisv2MjpMxMMXVTtT7r403
JhfMCUiIx8wA8khdScqtl75c/2ZxuG5Ne6ZK/n8QNkIP+nFgwgvmDJNEVowAYQbO
40hjw9kI9+rHeJRS14twdj40fWHEJ3aUJw3qTW4yEfR6lK7keo/aaSPwtUsS5Wfc
9LePwZUPiAJjgC0li5+1Vn6AqVaX7JiO9AKQj3Mqodp+6chGMpRg6kRZQZFmO0M6
4VuybvcHfnGTk1VkGMEPIdPwwwFUsATtRcbwi+DwsWkXdMloR6RTHN5BI7oQGJjX
hXAsFL3HC+5eMTBxjybQGLod0FZ6zwtE/BPHgJXNw+qFxN4YZXjQHnz0n0Ny0H2o
43BlfxD0ZJjpavnxvprilxDfpbey99VCssnjVrlthyKCpqi7Rr5eS1qmFfk2Nsqh
itHaGEcnVEplTRF5UhGdKVcvVhLtweaExAc83Rs9SEgBB0B3hHGJwAJfVb8rQtva
AVJWz+rkddVAZr9CuzecrBFNOkBPxxwvRxiTl2RuZSwlBbnLHxg0Mhf4lk/3Y0eW
UJaoAg8Mv8nOOuDOQax+hcpM4bGlpQAB4WviGfsH9571TZtFqbjj8/pBGiAK8g7M
Ngz54V6qvFj/0+7aVQ5MmAwQQT11ZFR8zrn51NIlTWlGXTTu4DjJnV+RoB9jzRtG
TP8OKM4Mf8Al6S9KcvbD4mz9H46N3Bt21iybF0AYVcBxunyvnoj6bK7GwIS1Q7b0
/hCm8wS0rK/iReF57gKVaQbYWx1Rv4lKfdFytr6yBRm3YqiZKNDVDQbrAfjb9y2b
MFT8ShzkLLKp/uYSy718r6/h+btpqpYMkT2nrMqyvoxyvKMvaOF57VApDul3r+kh
SuGMeIEOmDOFDvFQmtqW4W5XXxiKPi8dfdHgKXyspu0GqOdTH60udlkFyfTx+LCO
Ubn5QQUVhZtS4etbnTbX1Q/r8bxmaivf4ux3v09p64WBI7IHQP4qucPVZ/+JW0cQ
Jm6qYed15nf/um1P+9/BadmGV0fs9aZLtmmyQdfax1796SCEaMagg/klq7fOmm21
vfaVibE21Yh4RocJABcaEx8fvjwZi/9GEBtKSpc6ah550TTjGYwQNrNEGZq6JLkP
GH/wbUnBSj92eNnMbxIAHKDVOc4NZH59haZB9iJHfT6G+BJmB8XVOUilsLSbC2sZ
6JqI7sE+I32BUGrVuEZcCFx93chZdmKKr8STMbIt0UDlqpX154waeL3BBSuvqEWQ
p9CBJG0Z1T3hwXW5k4f7jKrPXNBd0oIaIe1yz+BwPkQArlJhQtoPqVdLrpR0mddU
zNWWOlyRon7f99FjEAlYG4QxElJMv5LQdKaqjXQKI/fXMpOI0sSN6VvwAhJ1WIW6
YP8ApRh0EuZcXF2Q7vQZ0S8AHDNRubqmmnRkBU5RCze2zzl8UMK9tbeJQn8x1m26
/DqlwDPAOaUU+yigXJ407ZmO8QT3kFwHcA7oBX2Z03qrRcznn6f0+s+OF94h3KzD
d4teCYJWwa6/+tP84oN92LUYxqYKjwbBo2+ze/XC4YVM6JFU2U2ftxGHnnkOFn2W
PEA+aEULYHEjp5wPnKykrj7P1YhGFE8WoDCxlv9esyZWyVLhKortgZXfh5ZanLqC
72/Vg6WJhyZuuKwErii3uyfF+aB7ILV91Zon8EXKukK4cJauNRXV5RJzfN1yMKHk
Mk4APEIX6yTGNspXKmfWXPTy9WCNcUmeKuIDlp+T+jArbbugknVVwH36jnVz6UgA
EmVW9QxWTNvZ+KDeb452emvsbTLlJ0Oe5Obast7AlGtjgMk5HTsUdvYgflTB1/6n
5nz/kao7XEi5HyY2XXYCFz1G1zmtMI+NFxe+ANUC6fPa7UZ0/5z676PC9UTEThRm
stxdDmMZO5oqb46WMgCaYt7tFlB96s5Zfnj31XymabRN7uybW91lGR+vTza56yoV
JJGiiz5ej1m/ktxxN3Mf65ODf/TrudZOwEbONtLJBjVCrwzFOZM8UYJMJZLivHrg
6/8DVeAWhYWkg4rfd7MOZD05v292gqCCI96tVAFTn5OXg3fbGKio5JWRpRYF6R1p
jtQSBJ/CXFWUFlWZMfyjHm/DZwD+c+JxkgO/33nAUeTUGE0gzE1N99ewCDFtIaUB
J8TkKB1BEk1+tAKXFHhWglBktTXfCtSObTg9u7bLm8eF/sDlqYN7tPBNOrBi6quX
3JhWla88mjkZavo09ZX25KC4veea6t3GwtR0A2J84GABI+y4iS64j/negNew02Q0
5OdYk6uK1ZHWvJn77vol5kbxFIAc/uJJUI26hhjRcVYcC9dBF7XhotiOl/UjuKlM
4cg16zX/iHFKnxV7kkxbKJD/j1nDgxiAg7lFkrJFAc1uJ1yK830IeVp1v0BcnWbk
gWIEUJF9Rj0e4gcV3N4iJMq6SMxZF1ZkDeVmLy+dHIzCaN1w/GQiXaPSibrln4mH
jSwGzwxIQxLAw5Dz1THLXM0JC1fF+CfUc3UHK0eQVavXMmK1OQfsPnxnsGhKU61Z
BbVvCWZSXlOm7uJ+zrN1J2Ta7w/XzoUS7Yy8xwStT8jw5UVJzfw63oMKsXROSD1c
Z+rjSdWScWy4OwIdMAmaZYBE0JIR25DjGJFymK49POcWXCbnnEc7c4tgEIkm7Jr9
RLi0VukRsuFQSiG/B2GRC4GYr7BNT+cyIVf452NhBDn81Ga++nJj2H1cdNeK0s+a
iKF4KTKP4Mv6AcK3gn77ViJekHfLNVTF19N/dzYIEyMkiLETYzJwNO0xDb24BFKx
17T0iedTMp1LuzKSclTi/LxL/ryqbldIKZRTPkbDtLPR0VX4+Y7nnJpxF7KTGx81
HB2Ii0x/bMDoGNIAsZFiFUHJTUlGO8mahRiQzzPEYdRdVqgPW8TuYjL+Y/kwQV0N
AXmlDf1jrXBD8i3gpek5gUeARMIoI1UiTMuMNsVHl/4jYBHimuuztskFTmGEnJfj
djw9UujMJQpF0Blf/36I9PAt8vJX13haSwkDejXKyOfPXQfOEVgtz8v6c3sVXtqB
PlzNFm0w+3NzHRyfgxyvEQwTaC/pbS3gFfFY/wGvakRlL+sO0kYYzZdSnV67R4iX
O4KsbCdY6HhpfTSv8Mt54eI1CjawrFSDuPJgUx/5pVwL2jWu6TPcIFzmFRAC+dvR
CFSZLp46pDczqG5Mk3DHRpt1JhmjTH7nsBUZxvTLyqyvMzNsnJOwbkdMKKu9+NDV
YYalz/dnjKgVHfdguHOpcPBbKudkg+586gYuu353ihGqBm3fWjLksUQEv99FECKo
ovRTPoi7oqLlLWSoaottFDITpZPaHED6e4f1hagHqjFv0e6Yv/PhqckcLPCB/sX0
Yts4qTpiP1QWFuc7oRqbPjajb0AayjIT7bMW2LvXb8MoTUzKzewER8VCvecVcLIR
/FW9VSnnqP829AMCI0qz719fLxgBS1/Y1l02ArZRKmlcelxXCDRdO8ZwfLkWE4PS
qH4eDAbgDELdYOrtB1HjxjawElwX8knkM2GTuDw1DWnHjIFTJ0iAc3EDuRu3XV4o
t+1DBqqD4sv+Zo3kavUF8BhBTJGc2rEcd71VdYmT9K7zcbO7O1SMREV5sffJtpMn
yw8h9o3Y6gYICUF5P+Pb7Yt7K+sOMoY7qQovcOPJAmN/xliSbWwFJTt8B/vBctDR
vmXmB8g+jJEAezHpXR7vE6z6EfJURhZrCC/o8X5Y8Kf1xfAYNVlVzBdzEfY37Rlj
R0Sv/z2s4DkZzqlOTR+vPaxNnv9qozZa/l6nIb5ISWl00I22UjborjLn5d05bPsW
IdSI4wqcGwZzut1AHhQaKJ7QjYN+5yQCVHOWH1i0d+6G6a5O7XhnHSajCj3G1Cvt
0ex0E3N7e/iTlFkgiaYntjZwKfnPKOqFjp1oPc+lQ/YmUzn7EuxuM34IwyNBA5bN
vR8Qd+kOYISCIKxAbQpuKwe019nEyxFOJMHI2KZG50yoFEw0hrXJDsNxMam6LUjf
ISarZQSVbNl1MemRSmavUZSnORjHJ9ifwEe6THlXNP7BdZm+Q2j1DGvSy0jPyCiA
BwxYFFKb5s/ADtY21tM6aD8UiJMxYfGb0hmp6w40Uec844VI3CNar1fEq8y/5Qxh
0o/TEbuSA3nxU9PpuYF6qawfDvKELsJBkCr4UBLrZBr1/jnWMAXV/SnQhtSEZcF3
RaJk7QFUFg5B8msLGgHGkMXloxhFlE2W0QWYYO2rgjXP5btFSobrEZv0vTf3dsFu
Y9gXthOIIdjh0tBH23wubg162ehkr2gEYG/P+1hIL0vjGSEMfeaFLA/+KGBCudri
7xzM90K7VMuHaKR8bY05fQDzo8yT+67Jas5rZbTNr3i+m9HmQqBkrvri7ZQchUcd
RT2finyNcx0iYi99k/rNBZ9ATC0Csp3nI1u0v92m3IQKzda2bUu2T/bymgKnMNO4
Qdk8Q6Iun7uTDT9N0W9vAE6LW+biJPuN2nLMzYTh+XwgyAwj3PBp39ctwd0p1kZe
oYVIKesenOzPr5B+MMyX6ZF0khkV7A+ukX5N4PlVRtMZ980nUOL4SBeyDtNxaQHW
Ol/UOVBRjBgxiTWVoAFPePx/9Ff8Qqqa8X0DLwltL/7suhimfphtwU+PiQhImS7a
+UBsijljnSxJ+iPgSv67E7NxVuesbEpF8o9B/ajq8Qvz4VAPMGjzMl09c5D+WPTf
aTQkvCm26F2UHXnQGDtzQFIR8ipacJDAX3cJQWvPfuA866DMMweB5oybKD6TNZLw
R6OXMZapWrleoqWtzk20/2uYXlZYdIecVapyqLQaXke5jhl+RfVO+xT2fZdBJhVm
OsUBFkG5hnDVr1EiNxHqX0DIRGCWXpxmdtk/OckIBKhd2gMFhV3eeuWjD4DeXGeb
4gFy4l0aN9dSUgD/zvm37nMCdmTyvZ3PWwxcbLvvZmMQjr0ihdmhFC7W3274sP3R
30KXy9eXPHNTQGmXMsUWF8Z8BaE7vYDF25e9kCWS+5lfAqLotG1ZsRwSbrqNDeqz
Uf4wiFK4HHs7A6+CV+bXou+FaoOBG9YC7occgTGtSYNtNe2g3kSAxAFI69QwVqcR
NnIR+J+0fI8Kqobt+N7AaWGnIwteeuxwcLd3E7LjMEi+m9leMR/URsl77MhPyWOs
GhD/sTuMRSMMWel1cj+FRLoXC1oKZVCrEtPKexGSr2wfhEEZWdM5lLfJvgCMS7OT
dEVgs1iBz7CNCrzFWjV7ISMhwtR54dnBfoW8myqbt9QF5w2Mo5NldlD2ulYQ3bxN
up9PAGbIW+8pnai9CHwC7+Bk3PAzxiWll5IzZma0dF2j+QtfTYs9E3pLMpVqzBvW
LsFn0ZIxOIJ/HTXRZKCt6Y+44uFh6KuKJNq2ozM5MI71yyoEu2m/iL9g7iXzkWjI
AhTXJC0fAemgFeUXoS/N1aqe5R3j6Tr9qz46b1kStG6jhzGT2I51gAPGgcEAmf3I
iXqiHZUzbK15nVHOaaf+e6uGfeEWV/g9YbxRysHu7qz8a510g3zTOJlG80plT5pV
vUAfg1sfJVYHvHMIuEg27O1JXq5wbFGOmFKqHuuEI4J3tj7QYdv74SvVsmMQHhpJ
Knd+7yY52vf8w2TLZkvkO/OZ+ulgo2bcCpba+vQq6MoNxLhFONFtrn6bJY7IMEsI
Idm4wpL1IhFYL69h789yycjAQE4YVj6ivoh3/0bsiqDUyTErkFScf39+DzcjNHZt
Q3BL9tnHDv/KkapSJeFv4o0bMRxqpBcVWLzwD3OExlp87+Ov9TJ54v8eW04/KOtX
p2f3V8UJmHoiwr2DjvIpwha7wA7VdrQVAcAz6oy+K1SJes/j1BtxqzdKNl+V3ZV6
+GMRcKvrU3oXxtZ8iyQfPCwpbiUn3LYc3vZ/ZY0vD/iwI0YQKJVL+vxtpScMskri
AmgSKTKc5TGin2dmq2mV2vn3qcCzHBku9fedQvxhmrzvX1BxdIUHvUU24l41tzS7
MLwQfEQfXCIOZSVv+AJRsgI7TIVQyDuerUx2jZwYKeBrd4b8GVu4bZdKs7ExKBH8
KMzzHkAnBtilrs1HKIqoAVNxON7PKg0y6344I+fozDxIfVOlMnX0oTXWN+v0Q9Zt
FZDjwhpR4KnVoOPkhcGAZGSGZfUJ9AH8u0LUV4uiC+rukEkI2e/fNcJaLgY1seDP
YIX3P6hBmlc6wmv2c9JgzJVDoqvrb0Qd0tqf9quCFYlOQ9Eo7aWG0rHSPKE+NrbV
YjXHV2Yjj/9/mkTTwXq1c0ts+FFlmOki7WsUI2+/u8fmaewC2O5SQqWAwC7jEF5E
8JaZYDwUJpWbrbi/bv5XLADtM73u8zk06it2v3hiRUv0rDC+Ks+IekHZvmVsWu2J
+x1Dp5kXojV7mQDw687g/DgvdoqfeePmu6OeYII1xbyb0Rg+qFFz5br6T6QCMatH
qV5GfxSet3eYbJ5q7cehFv27p4fbJFVpjgxea9IhX8agASiUtc7S43j7osXnJzJe
FofVULqjeEPRlhG9KzAQu4FHUQ3i9ETlxVhj50gmd/bjcWqcE66jbHBQOKG9hozD
MtmO8Sx8r3af1cG/k6EHU6bZ74w1xkxXwTiN53n9eqGH3DOpAUQjqy89yOGNIKs/
s7hawy0ZywLmHboYUV470n0PJ2KKDN220A7s0XR+XDULB8GgyAG/rsV76m13Vjjr
yvbZX8fXFVlDQ1orJRRNE69tEGZerdSKB37BgaDi4/fbnXUKjWxt0VTtvnY0Tk2n
9Ak4TAzFXehjdjISo0L4TiPhyQ1suLeJS2MuoA/lQEfZcqozBUJWA7p1bjyDWjoA
QxGKLcScmlDKxJj529QGDrPb2KB0UPV9sDa8b41PrsMsHpvp1aoe4VqNyTm6VFAs
Rhpn1CitioWE0jmK74k6OFfnVWo0hSy6hVFEDi0QfVy1E3vwoVol56MrbtO685SM
mxIMqD8OEgev0GFp++YrO46UVs35DDLmlnJbFPqEOF2HT3AB6R5HTzkl26H97txb
EQehCZ2pI9ApNwXQKiEF0k8H/l9Fc6/dB9nUnuI6VaYzLAxK/ynT3oWFrUHzgpEC
RFfgzx2YtAbB09B6obqoefiEB4mV701nu7N0m33VjkevxljJKaxahFzjVzRS5dQ1
bhjzi+uFx4hZ90/l4GektNR+93fmgvW9XpYyDGpu4D4gY01LVTjqTCpZXcmqf33z
bWqL9whrmEp+dqpSSIKiKpJ02CNTPsnxJMsryPMIpM4jN7wYApTAqjHAjS78RVY9
I72KJbydpI8Aw93s2geqCDPqCvN3fdHckw7lzYV2sGWnFb/vypCem6zaMYFxwR9D
gnqUoYwxmn6sqyWZWEMCHoruoFY6DW1LWOL5R+p0W5sEFko8XPma/So1mI3eE5dq
eWN1QDrtpFOleuexChWcMM0H9pmZenrrlPGP5/PblIJbekUoIZfjBIYCpIWSqqh7
yfMe0s7YdQRdlVUlzTjXn2TXQhMn5RP5xVbFHnG0Taq4CzciLt0BlrzExtHrW/oi
l82Qr6+MHiVsJzzqjey2mzcN6bShtEZIS7WzSInq5Vpzkr2+QELoUvuF4XQrBcVY
pXz2kCesA6SCTii56ZfstXFNdb7kaZGj63tEjYGtQFDvpMSdNqv2saKU8Aidttr4
P0VDLyajJW+REw0Y0iZvmLkeb5lQcVxHCNw7fUdLxijK5upLwss53gJGTaKdMeWV
d6saz6FTICzpGiNPYbBKRsBZ5fjQIbzKRPqyy6IUcSqlOHCw0rn2hz21AUevELFS
2SCrRuM357pIMYYQzEREzeeAb5HNEQmaLAfDsemsnqcxfTSiSIAc5mGYhETm5G0Z
MbGo5xKvcTpcodh2FFcq4jT5MX2j5vbwvqe3IIrv7mD910OCNdJ2CcHtn+gxUTax
w8aeAz7XxwpoH/1alWpsTQ9OfPXlx3KiAy8Lk/FnZS5OxVRp96M22qpetthb4rwW
2T86cmW+BLFAILs0cL9jZxy+y7Ai4aOD/aUfcLqgybit2zQVV8ZEaHWfI9sjNCjD
Rl7k93ww5JWnrhLVD26pLbmU9nFDUaE3rVDZIzC7vBsA6dP2Mm/XrdTWF8iK9O7C
tMyGmmvSOdl5B8ypTqbxBcjvBv6/MFYITZkezXrQxkoEuW2V7sKUBNKR1fXHnH/h
IDcCQ7klh+uYNI7mG1/tC82Vt9MXMyNTBLeirvelzTZZ7k5+ajeA4INwQgWDeVdo
J1jsM1k5m5HrvsJYh/+Quq8Zc7zwcP09dARduApN4SorJTSFgPo1v0g4/iOkAJ7E
jElG0keMt7Sh9ZDQJzqP5IORklMT3jCTdzyWHfEolQAn+xlKTEriBh0hW9/YAJvT
9f2E4bns5WTO0DH2m7rFVBBHqnVR6nv9brH0DQpmJFLo2DadXr7mfhQZGvq7g793
iSHaLgKeYn3kxJ6gzHN4nC+L34mIBI/NKOdDt9E+zsiltnsXFwtHr6+fNpRiW8Q9
J9cP+uJamLO3kv64OIaW/4CYAch7xHW9ukuI2vOC8ZLWS3M+ACRIzamqFxfpUdck
5ou0T8ye0kGbyBNoL0RaKQr7rIV9+4rO/qzWRNKtJzz2g0EZi0zSY0Y1ZJ+dseqN
PHc+NQH7bdOARfQqAlLTjOy9ERtVXt2NBcbbJPyNfsGR4NBvHuKCRx1WqvsdJiHY
WbCB80wgNTMCT2Z5Wy6llVlO/vGEbU4YzFBSIfeieJyc2d/MyuWkmNwlOcofJmqA
5Vg7pCv15LmbjBolxfjt8PXwksDvX8qhxBh0BkqrFJR3fAzegYcURXGXZsycWPr0
P4pHojMgyb4wnvXkI5oCuKdDPCTXCkuP7jWVY4udAVRNDMC/cfcJMkS15FLmv+ib
DIgQZ/8HKIUokyger/H/XpT58g3JdFVc7Ai8gnysipqGYtzSuziLdt2Ipg7FBCoi
UCBVrj7psM0p0sErQ46/XhDrkgxw4vX7C284bm+Ek1Qt2i7iLe5GWZB+L7GJITsq
y8xtKQNjTro1ozAtPGP+jM2Eys5wlD5k3e+1XQJkOyTbABRiyKKfm4UeW9B0bNkm
8JyzrrOCQj2EtvmgmPTc0oLO49MJw6oSfPlfrN35ZA8+jeT289xg+YqbSfxKLegd
iVgH1FhA1cd1T5/Cpvwyxq5j6nW3aDb/sOHNh5mNEQiJJ0u1ZiEimg6qpkq8qVdC
0HfEv9QKL42nj8bDkx9K36nMfvNKyT4kKRjwNIq+BjRMoo7Wbgg6/S22uEMMZJlw
MxoMEyJhPHnzPp9lHEfVtRdW/FnMV65bgnWfjUEKwP1xR5I0HIj+3PHxPFBBYNtE
J1EaEhuT2M/COp8Tc31V1aET0G2q32yRSgpFle7fKOk00I59splz/EVPc01FsanP
Zp4Y66lAM/Q06UqOPb2qCrtQyHJPWydqAE/wDhGmEvZUWUxTdZHGxu3qRQw90+NS
DU7rlgTLzehFVidzsv9GtU6njGNLWH8G6Eo/eknmTqVqk/vikt8qzp6f1U6zwyvR
0FyIEw/3fBiAcSRcDCEeEyJaEerVLkGJTw+AVTu+7vOJOS+kEnatmI1unT1HcI5z
qCy2u2VTr7fy1uuy3a5hzwsGLuyw4PYbghhw3xi9Wkd5szv9Y/OxTGyOosM7PqX9
ZAs8Uy1fVJT+BFV9Gb9IyVtlAOBtQ02toTGc5n2YUBrSUXnV/mBo8OsR9UxI6dMT
0XgJEqHYmoGxlVZiz55HkHrTiJ6vqX6za8buJG/I6Wlq/cX742T9yp+5AupW+HoM
BUt9pS452GlU495nUIFwNGQM4I37ej55IjP88cLFK7HbQSyBsjefUp0UUWTJcMpg
Pt7XMZtHqYP4VKKg6Pp2xNDp/m8U1B5bjzAa94svyD19IeJpTDg0FrWRPGBfjN8+
/zcEUxXSMiAoz+EGI0lGvHqcwE0y3wPSBljMK/quL8F3IWt25xYDLw0C9VSQspKE
HbCRn40uqwqXA0O2l5d5lYviyEirbmcqKBvwSv9PwHjdp0gArsZu+M6XQaIc3wNa
YZ8iFZkKuZuUMKYtupqo22zpw6e41QXumutXnVHFdYz2+wR/DNvFnK0do45p5Q3Z
aE3Lm6lNMJSCQ6CqcFU/DmAJ7vC6lkmdYlsXE5MGsYVcjLxnGuHv0gftDPfwWHwj
/25QdQDaJkh1wyNHsMGVXnPwgJp+TeGklsudV5wjukC2zRV2FPF38w3ESPjvmiu1
6+fRD9PGW1GgT8Iu0zA9DIrsEwannQDxuViovbYk0DqoiP17HTle9J4gd+5j10Bm
RaaksKxqE9YicLoHeVHE+d2xyCzH6m5/ATgLzCmu36f/WXIECsTuaVCOteqwuQ0A
eLYxPtmjyeKyGa5Eft/fwLbKVhWzJD0azmyGetb+qPubdQlgibU4wqOKj6hpAwv4
RzOdGgxSvmhkVTwXGb2FAsSLGF8XqM/Q0iKhySDoKxRXM+cLRlQq22uRGMHBoPpx
ZaaJTRzsv43QwlvIstYsCZl101iYghBab1Tg8InlswcNa2KawOeNbHiCSW8Cktuh
jXdZc/Hdc8bDfrlV2tQL072DTHcIV79ZjJebtzXBO5eyFTwidp/C1q1tp/yfJ0iQ
jekQXYmy83wtvfkllrPybs9uqESPojivS78nbKPjnzjmsQU1TnXRfXOj/JI0m5VI
dwVOC1uon5q8Ac2R2+/LtjNZW7FLAAsrNXpWglE4kEC8+xCN1K9zmXvf38qXumii
8+vn5897OcVx/w6/8XeTaaZ3Xy1FrOjo811mh6H02OAdrQdkXZBi0x2s1H/nn/cn
ia5k9SU9aKRssxDmfSodwHE7oUjfZDegmE0qvxBH2o7ChqHrYZC2h3gnHaw/pOf4
TtdlTCLTQM4BGvHp2ZIwtvVbfce4KJgkg82BRl+WjBAKv6tmhJkQB/J/RYwedNCg
vVOfzElpQdqITgyjuZlHlzz0jtVGUKBLEXjb7hxfcB30Zvabbqe1dMJdVwiuitlf
cfSaGR69tfvP3VKlTubFWpB+t0GBOQeaszRRcZUelcLOHSkJYT/E4zVlizsDJXZ+
VbDeyahXvreRspRi9LMAaHzDRX8+Oui1a4yAs5cA83ufaoWq9fJH1fYAawPs97tz
BHnElUmFdLmHK68DoX4eqOUFK9XZ15cqTiBA3oUFez/JKHgQ1I8iZsoJsCJJdxMo
sIxaLlV0d3Q0LnbnfLRaRp+hyCbz6pift05gQgAFDOw7Ur6UckjCVMqiCnsekkFR
zHgKPbFjAA5dOHYkffsGyD+0RIH/NweqLZGgC8AnEV6zPJ7x0merKSrDhMbHxBZW
bD5DIa4f5ZASJtnF879nmyTAMEaViD4zduHXQxtlgRQXtmoKiwATToP64kjyA54M
WD4ej07DAml15qSafYKh7vPJMavEPpE9+aKHbWqse4I7+oQkhKbl3c0Kn4cYgA6C
hqSI8wVyItnBlWGyvTrW0p2/0HhIg1BsFwsHhlxEnoNxQEUVhJ9Kpt55nqHX8Dkd
f1bXBP7Xd+mzv3mDn0/TRV8JQ+GFVTmCQ5KCRFuDglUKkx0eiOIFDbfVja1/rXbv
5SKvcShf3j2WQWeL2l1mJOFC2pnioUcDU1Ys8ZCJl9dXLhpBVlqRML2uGjzOw3D1
lYJBJHF53nifquCoDJYx0yo8OGzgiwPwzU4bc6liDjnvqcbAHoxlPa3ZVm4D7o7p
lMlB3APYgIqee+MrsjAuIaELPEzitEn51ueK/h2iVsUqpkmLR3iha3Y86tA7ZqLr
GZEXMv8bJUvqy1KjeMz9ImFZ/geP6RmDzIbPBw6CgZ7MeMcAX7O+EViGVfUHW+9I
FuBbJtPO4RrTzZ6uavsGBExc6dOjF60NIFj8g5fjsmmZs0XXaGCVBDVFWMZpi5Se
2lH6Dsyg7FCjz33qqeeiplVpCetT6xZlrWTZZejc6a3Ryhoct9NDmAPHKvbdJ6i+
Cuq6r76EYDotBySF2fcFBjHYNQhZrKr4zcNWt/pgvDau0O/0ns66s0K3o957LCSt
ES9nGolPB8b9Sr4jRREn1PfdOJwSHGh0qVoK2fy5ink8Eo8OxCgLzhudJJbzRGFG
VivnW2NSaUVnHIgERfNjEadD33GJ5lYjHTamctC5IsLjgB/ufAO5Ruass+D/HKbq
kUm4G4RceYldl926R8RGiJFLctDz0j8GhzIKTkPP8HL8H3ulplmUBr1m8H+BJ2ky
T/zSo2QcV2z+CSc3NaHn4CcXpjOWg+eWP5GUatOZCNIcWLPspERtK+b+uNNg4/e4
LYm9ZNVvVF2fgy/ifqXFqsd/fIUKmrP/RrEQ74/PTdItPs1L4XJNFTjXuz1jW+oS
X0AqxBBh5Viv0pPsS1p1H5xC79UaIRRNsj/AUImNAFjSuRW/c59yOXTTFf2XWxV1
+tPYhSNEqapU8nG40ElRxUpklNP92lKB5jvoyICjrZN0pTh2HnhJjv8o8cQDupGH
O6qt0YJZKheQaZhTVL5t8LGiyU4ECVnGoAi1eECZMOydWnVYU7Oz6tZLJw+SsV0V
33RKL95ZKshUSyYpu9GL0dO9SWItoYMFjl+xMJgU+2cU4U7t/G+btSzZ+UsrMrz9
PTxmzLHxweGvewktZ2xSSt51eb5LX7xQNa4VarNx3Sg/Vh2QagbC7BzXQk35U+XH
6TaLDHJYgEizTAov0xl6a8fyOCZ24j8PgseBHoKg1EEMlCU1x0K74RWAa8UWM9cX
ayJii7xE51fsEVtKZwMo8D3efZA4d43TQB9J9nZbnnl97nVjzdGTYABPXXxVp+Mn
Ue5AqO1yNBGvJvHXWUTZaHgb80VQ8DYR6++UcvqY5UjFOdWohucR0vVJDR5L3mdx
eKC2m6/5x8l6QH7SNrRowi9lpPjbShhzqqfaFoImPKjye8w75DpVhK1lzpcgbdMu
J2IdGsZr8chz92FGBw3+BtBkXWu0Z6PvkYBGyeQIOVMZjpprrKdwIcDikixJ295j
/u4XDtiwcSj3Z5VFtiTgxJvRimCEy++PRzXcQaj/eU+JAt9Xur6VsTtrq0NowsN+
cHevqlxVDxScy6kpniy4aW1Sx172L6UtVCCOjLgyd0TzfbM7Ty8sG68gsdbNsxWB
MyWfBfMcaj33DqUsqcR+2hMsx0BPSBHV1nDwpoPjJx1dXWoT9CS1kC83US9E8YP9
vgfacCmRSe8FgUBWHbMmdUYwDxx7Snj/K5cDRPn95F0iSE3Mty55/wR9iUTYdgr2
XK40JW87nv9NagxXGY3Ud4mKvM/d/9pCiCIbKz3dTQqEZr7G29eV+fwcmbafri4T
zoidq/2bm39dctnIXGzOlRO9KJmtcBfryvRoBZ/ItFfHZkebRab/PgH78nCf430E
GIWypritLIZw+rBFVfEWlj4l6kSP7lFvDv4Ao61Xrulmd3EJ2QQqBwoPPMmjzrKt
L09EivpT+qV+YkbIOrUWtDVJiMx++x99mXGFLsLpESr3h7k0UDm2CvcjJ26vXlgz
KbMZ5cMhXciFMJGDTkQDSlw8h4SZFLIBnR1khmwf3dL3bYqKuB83LEevzIQufySA
Sc+j4NGgYtAtVgBBQjxC1JA3E8PNPlmJMMKOG2bOkjlxkW5siQ73giAgSsDKe8vz
qreIJ8A+ljQCkuveiZWvUn3FhAc9h6uK8Ofy4fBfHyPD6ksE5QzCn01+pi30M4Ay
ScgttPgLxOL8q4EUUmgl+BGYg8Jwo6d9e0+FSXR+j1llOZqwPg8jc1u6nPLyss3/
e0cnD2nYSPjfnbhIfYYqQpMRioR7TbhsVYJ4NdSJut8qa8XfEJ1zb5A7tQMGKJLh
U52Ia15bQO/2jse2KHcp1zMaXXlsx0OVOpylg49aaPK2djxVRy5D4rwJFrjk0WKm
BiDwjH9aaXBb/LyxVMKtkCkXJsLmKxESD4d9h9WR3ojDn1UnUJObeaVe1PTBrdUI
45RgTIpqcD8yReIo2RYkVO+5mPJySvDeS/bE/YYDHlLRaepY/mRoRojlQSRR/WKN
lRqmobdgqomWmoA48gu33EbChgxNLaLZkCQ8X33IZd1ZLWBLQGyyzsyOQ8jzC54U
ZiIHHfva/XoqucUWTHcy0dumsPjJVhE2oPktNfZQ/Qv1thHdI//a2CZHYHq52QDO
A5j+rMyIrARHbfFTrCwGmisbMaXQkpjVmRJD6ajSYrmsYDR9xx+VVddcY+3U6T+G
+epE9ssFONrjCO0VOPrwnHl/nLvm+GJ3BNjWhzqgaHe72mVrhGF/l0x5k9VlcG6d
l5DzigIJHCvQGLnpId/1tyQ72tr8km6VnqYj8n6z4K8kQ95FJb0+nvTqJ+dcx9II
uUmIG8miTaD5nvJkYm455tPc8PlOrZG0EdfhmfocMP9pfzECFcKtamp2QrjVNKk6
QRQSz0XJWKqHSwpnCd4Utz9sb6AIOZ3zjG+d9dkFz8VqtsDyso36wEEBQaWGmB25
mEflFTkwh8G4IqBShOB6bZviePCGhJRVfUYKHBmAp7TIYGQqyzv+dN8x3mzNiaub
FP9eai/RDpSJHZcjrfD/pYC5L/WUvDpXYZY40h+/NJhckEtZPUKoEcUP22atZmpf
symz+u9HlAhn0aZVvMdA1Cbke5tDjFu+T8AZcUJWl5Z7IRhe2ABHJmtk8zxGTduw
D6Hq5mOy3b3W1LP9QBtH7LZ4xXs7+cK+Gf5c0jDaQZe5HgTpEW+z6Joh9Ufz91cA
jVYeBK12eMUIMEWXUTLYJLSyTGrjGjEPeKPROuHgtli55WLWwbgITeOeytAigoNC
9bkmakKMW0zhmtBgPvjgRYlTbEmp37qGOT1EWUnSkaTAsKbLL1q2zJWB3OJWGFpK
/xQxakj9nb9r1rWHVXz0AQTjFqQDCpJn9ku/BXGYKZePtHYXDw3osisGXPZm38cZ
1sSne80yEXFX6/qq6TG8UQtAUeFzQPcL5pePxE1tVeohevkTtPcyL9BA85fYIdF/
FadKWn4KtpFv9S6V0pqPeUy2u6V6CzsQp02TUr8ChYf8oCh6Mn/prXlMIxvNaEw2
5RW4qum1LOuVNQxIfKiqeaTnXF1a+0/a0XhgRTeEkQtxhq6Qrg3wGlgCqh2cNBvg
RJAKHeY8FAYwJe/+tWj9/z1zO8L3Syef7K6vAzMt8Bklt3CTsFU8WkUeNhnP96dk
k9RH4RSQ/vO/A8NE3t0IpBQ/0PLrVjUUChCZzhKdGBPxrQstaDJYVEyBgL+uFm6T
ClsPJcrbgMBZsgUU2PKDAglAwHcLkkeRIW7sC6QHTTTzTGQ8g2qfoX6Z1CcN1w34
RxoEoP6ndv8if6aI1W9aj2ftS6z33pCbn+fu2JsKfI/Jt2GGZCOtFa4e1iLJpVk5
LUolJiXVLGmTDer1e+PnkYqt3Tp9YFotytF72MymTWMT1U2A0p3TChKxUF1BuPv3
SVRyPE3UuAGTLbz/uYQkdoDjz6U0RuUSHtRs7q93rBf2O+TBawMTfvaxw/w6ICpV
dwrKnlpMxFXmmhNqmbVOHCNmjepW1XjnGxMaaRxXSAvYbMD/3LnYx3HYZ4ub3GpH
3SJr01Ez2He2KYGPogMPG43eBkd9LB9u8y6ukXKY/06jTnC1/lFlGv+PgQhhzQ6w
b38iaA3fiDwCNr5VWivgwiiEM/ggYOMgL9xmNx5nA5k3FCLTkUxSjqqhrOILNPwN
SQFmr1nrD1ZNk0j3KDPPWGZSqGKxfHikORGLR+ptbrXmhyO3+fggGZM43FfmwpZh
LTziZ/Z14lMrlE3ztHK9kk9klJWCXyHrUQctdrJIXXBu5aQ8ZchTwjUkdrF3uX+n
NDQVhaqiLlphRfkuJe63rqVCBmU5S9yUCH5ogHqN/HcXJG23IF0f503CIHRbPV1/
gm+sF+PpTDdQlUPhWnPcTLkkWgYUw2SdJ1/JK6u8gZXsVpj5nMO79g8dwUXNCZt4
fRGZjkBCliPBZFMPDR5ns5tKNGo1K4CLkVFaBTq4TnfeQg0iJaHUXUBDPqDkYBxY
e9dck2ePVAO2kt7m+Pw7IQRX4IBwk4dwI6JVSoqqkI9B9DBC3oxwxRiIm5cKQTRl
OX5oDr9RTiZbO8HoPeL1CQqPYtmdxJwVep/CE+5StU6ptsm/OlycXO3UlyOlRqPT
i7wm2uVl8FPs1pastwAHw8t1gLQYHlVfNviJysg7+GEOueShCRyWVjYGo73RKBqL
9fV7jy2dG2Wn52IzSR2JHMYuOG/DW2vOMjP5dI2IukQ2acUlHVlmCPgu74fUuSxe
GZxT+H4rw8m9UmUgenhr/7O6zki4jvC2bbafPgLn6Kd0BeXm4NVHD9O0rMSF4AeB
8V3L+BTvPK2OG6qCKPLbn5Mvcb1sGwHTmgvkgvAZjkaCnKpDAuZODzN2BTD+UvkW
/q0fVTWXOwsOL9atOQwgey2wA1C6ocKZ3zNQ1QE78ebbn20s6gjR5ziSLeWeL+RR
ecA9nPzxQ5Z8/FWjL05ZEeS+uEHsA4ZkpJhxeJYihEdt7JOB6V+uwDoQ5+a83WXF
3cZGqX79gK4rJbz2z2Mn++jGytpzua7u/crHD5YVP4lbThZB0WOATz/oiWzlcHeX
dKF7WfFOb1CmnwaChFc+IQGAg/4slv3wTgm00ZrolZnAJXojSCc+VvC3uy8E7Y5w
CVVFsqb1RVS7MYvEVImgWKbOrrtqN/uw/I5WXJblts5WeFqLtJ1Cwe0WSG/0ohlm
ovLdDZWlgKMVxItlkdrYbXPjOteoMV40l/8bDmBcjLCyPfJ0aeqnwmby0PIZyq1l
t9kGVht9CiGiJFBC7W9ap72LdJQfVaN85Cd/H+8hZl69ARyTu8xqXZk5LmQQztQd
hf/1nGnKetTd+9c3qDq3NZrSQMJtDcHm1fKEQCD1mqy/ZzvZygI5ZngNIiFaUsLN
KlR1/3rsyu2xP1Snx1wkcEOtDd21grOypGqO6JPHk269GLtQrBEW2qh+N150qUKJ
4lPorxcdWYTKE7a31sjAw4QhiuMdPo2q7VI7PRrfFi9g1b5kyiARXSKrdQ+xTt8t
xXLC6qTqinYafKN4J9ZKnj8k0ONwvs6rk1byPY2PvkaF0gn7JEwxuRJB8ARw2MsZ
xqjKvJO1IHcYWjrma5NYAAx1OOTulIp0sBCwaccwtkseEwXcxgLhNOtTkwVYoeEf
zb5oYydm6KAQojplIx8yhVkd5iRmBjQLfA00BxYuFTosLkRGklwdeQNUo/pOBL3J
0TYTVZ5tsqJq5iDxzGEaOzi0hyWO6BpHACE2a0abfpqnC/0r+iUU2tvQEaCsYGgY
Cb/dpgHbCufwl6sACAzDR2GnRVU194jVymo9WvZP0Wp+OJod4U8PU98EHuI62fnJ
fUy+QA6sOugcsLTVdrUOpOe0H08+3Y+w/i2cHDAH3lq+2LpfSpR8c5asc1kXYPdL
zuSdlW0GUUNGUHlcusj/AUQeNilg/dkpOVC2ADwpkALLgwIjH9nxshjZRXkkSo5D
hFs/UKWoXsfsJM+phLOmYHezQ2UwF9HZImkNvtJ3UxLTdBHnGu7I3B/kPPvC7rL1
VKYwbAYgfhq7LuyejaazPpBe+bNwQIB1E5Ht+gBDovu0mmMrBYSmvepSTwhhydt4
hWIy8bO6u92TgSxfLjgSUbes8zJrLSR80hsoFftab8CxsLFKxNT4W6F0qBwyVUv4
034t+mXNSEDruZ8LpgNutf4GGplm6z4lL8PlrIJzFgjHZmU6kmZGLSS7QYQzD++L
ryyxoIYT4WZGRGxUhIrtSHM/bsdZjCFK3lWANH6P0Cl0ejfFdrp/VoWsxgfNJ9p4
OKmM7qfttut2naI7+lL/NPcHl12JXooRoSqqtJUFf0neiTvs7DdG/XaGGEqjsvdJ
PRXJ5qq0cPqv2zo8zjEr3k3b33+z5VBdEqIwVsU/Qf51+CkKcKuvRK+WnE/8k7+0
kgdabA8o4UsgjPs6C11Kg70BK+dcc5ouzaz6PEJiC8k1tUeNrvm2L+Jc+2S2dduf
Z/SPne4Fgs7/igYr+mwkSHV9vMTxk6kgkgM49cR7O4unb3oRu+q1yG7ocb8MiWI/
ElRezPqgkHLmOZFUgObDtqnruCyrYHJCCR1xU6dctbDuwUQTdnYn67IlrMWemaD7
wx7Fb/VhstHeCNKR7yQPeULy6T7IDFsi9vr01r9iQ2yTuYUsM/1rQIjCExb+mT1t
/W4A9IBp2a8LK+wPs5d7uKyKJ34WJNaQcELjxMM9WTb170GJpZr1kv8FbP5NkVQ9
pq6+97u/fnjWvfqUWoD9ugQIX+vyqdrs863KlB1DzzWVuaWDC6OfY0GyT0bv34Rr
ackEOIVCn/lFlKnS+4ue8aOeO2YRjB8e+6o3hQjJ04L1JMb9o0HtOcTkpsK8KdaJ
dC0eb2KEePj9eGN9DBMc+iU3Dmd3fP0AtgIgedunzzqTCQq5kZ0d/139sTWtJPf3
9+QTfT2nXZ1uW6Ub5WEzInHUVYmbB4lMko8QShUZ4suJ1oaoTuxFmBhafua/vNCe
jBOUz6ueQD/nCZqJc7RTqOCAFyVZqyyPfLq5XRujjyTTKYu7SeL34OpO5OJ59YhI
qRIxRDdQg9csQ60SvwtpN9zkMwBb+KHSGy9YEkd4QPX4lHIFdnfqT3TPekYkrZlI
Hrtn+EMod5faKpAspuVbNATN7GDDzCYIEe357Y4sJftULYWbV1lt2UNsy6ma75Ek
sohztJ8+kihzv3uXFBUqsnuVnrfgSwP4wMTGi8GbshSsaZ+HOKbCYtVOMptBk5SV
sbTvxyFbfWZ8sStfdVfJnnPE0xvQfylUrEBuM5bBQh2kkEwI1HXxt5rgru3pUy7K
PyE+684lS7OuQWlVsD6pHdlD+QOgHbHVcs7zvkJ8sSpNXBXeN4kW9OOY2NUEB5uf
epTg+tMnGfJZaQ7W19wjtps2OkdIMMApmY1ulAO/9ASe2D747OEc60gaCimggCre
VCJKmo/yFBvD94zYYeXW/ZQkrHs9W1phcHb50kofGv6yxtA9gdVtF8JO450BkWQb
u6GzcK9Gr3k7AHW0LqEcQYXFQPWCKHU5I9ZYThtdZsadxLeoQuFHI3rWQq1mIB8T
AmYXYqii4opvMKbhcHsJT6KmqIep8Pbs5BjUN3AQJfF+HbKrmRHx3b4RKjS4oUrN
kwpV3WfusY964l2MZ7sSXNgHVhN4nmCZF3DeAJ8CQhQQaeLYEEongrheOrcoLq/u
O/BBc8MajzXySZZ0zW17j6Z0mAahjNllZPXQhDm2BxNmWRCjUf1PZm6rpNBpJ090
N7gSUiYSA6mxZligXVjI7XK0rjaHOZ9agP8La454vU1X9rCghkTUWvH+rjbGomHv
KMIus00bakG5hT3IZsGL14AxkKwOyjPj+WLIRTeuUctVmSfzxB6vwlFut7ckBvhc
259+lB10bF3XhZJMjrEvHC9grmZ+FrEwswbj0Aku0i6zfSTGTt5LuUOFzc53LHS3
Wp8dGhQb6tUOv5ZGNXn2oG+mBiyLxPOHdPtiRaGqVVOPzpw6QalVAw64fIlW8V1s
HXjk3uGN0c/wmpSnX5tM4iFYg64D/pp3hz0pO+jEzu1stzC/8BvR9NJjrOMzpxHP
l6MgdcduVaPke+bURo0QC75K0QvGa7g3oq3d9npFEx8maNMkQVq2Oy12Fh+YkGdM
TgoJDpKba2yQA0rN+izJP2BBrz0z7XI1PlSA3Z2W1RC89PGig443+1P2INgpPRaM
ukkjBbAC9iC+eQEl8OLbySChqqo9SjtJpfMWn4GuqyrAZg7s6bD9O129RtXNJALB
yh8kQ1FnH8kGqdX+F4FAzncmQnFHRbw5nHd1yovD83FT2E7C3bldxQjBVZYnwmmr
4vSANBX73lZSHKj9foUhIIu5rI1frGAZvfx4YuOpW3ftoLKBRUW21It5bM/Miyux
GKe0MSDlxtSpJuUIhnSGCXUbYpZx9f7M5muEYEMudB19QTxgrZY4kQTrjRjpdsQ+
JIQr3X8HBHd6K5mXu2Eq3xoqlTYrQy4qxQiPM7GlZrQ2UrgjUoZjYbukHO4nzK04
zKLUs+OUmxuNEXFYDMDkxpPm1WwB8lWo32zNT+cV2dJll3ko8URTOvw71IuAn2CI
dYenS82vXm/+Ko0yezN9udC9x0MLYoDD/EUAVjNXR4bedTKiDbS1vxsr0g+HjQFE
DFudImx0R9LPe3XrLDgNKto6eRSUbPC28jIJdrfUugj2oiDluf86pesqH3zdGspk
69o8U76OeS0oFnAYKfAw4Jw4DmNWS+mJHTnZHBx1Xk4xKejmRWI3PMVLk7Hizrop
uh1qks/h8pEbHa5UJLX93REsz4aVK3tzefcN42hQXB8fR/jgOOg2fghhyx9FXE6x
F+KLM2xCaJGP2/ScP3G70rVssfQbGP9gkHSSRzdD1wClEDdJvHxmcmXwTCPm9D9P
tSRHtjCd3QmbdKg8H53151F+Z/Yr3702loajJeClZ3AefbDwTktE+n3nslrVB9eT
kEM7j7YTIf/Ko4o+K6PeSywsxi+A5sD4EBB9hRcrAo2Y2aCsJBI6g9MG602yGkZe
TmaGIIbhZrwSwgF5dO24Fy2+fFyqigO41XcxvCur1wVqyxSXfx50DrjLD/AzJxim
TTW+gtfZXwF2V/j9Jl+drecxj2RqTJ2IcmTscjQd6IZIlvLwakPeaey9/3B2je2P
5DxXDhGOaTS/8yzLRUNWh7ziPTZQXS+ktu8TZddO42o9YX+cMDnsV4QGWhKISZtY
DYlgvox6a5xNqqwayHQRjAbFUiYr1DLAcWWX6O9HsohfyYEtpWpQy2x8s9d3ybOT
fajgSrV7uyLBOgqX/5OsMBzeWfaJuSNAff2Qv7Dcxl+HFNL/gsl1UklEn6YZT7vL
GDBMXm12F3fDosjEzNgFJT1dxIWnsVo7t8uL+7VPuQM8W8nL9Yz17ugRR5qYSXlk
2NoQjcVhwZXHvfJ/cMtK9Z/gSMGIyTXjSCCyMe3QPfwzj1O9DfuEpGrwz1uN+wPU
ZcF07YAqFHNUHT1Iy/SJmEIVA1M5UjmhPcECJZnOIHXC3esrR4ZuQKIw9IIk6c4G
gq51Wh8S3oSrGLV/+WbDkWMUsegjm8sx64wxxAoeX9fBDlNjZjHJkgUdAXvxpkhJ
b1PMAe0+TdRYjLEwRp5zNsyfJBLGaxpdyAc4O1sbKcd0T5u7T6EtjKyXjzaoku1f
VBHLoFBxnLGQvsW6u//pAdNNpOLEG5gnpd5rjQzGyFF747AYhlEux0dyHA+wk6Yk
HGJNN+SN+joYVsXspdAdSb4BtbOCFo8S0TlZ2f6NhmDPS5NDAzg4SBblE4OOxCbD
LDzrQJPDyxJ5h51SU429F3fE6ulG2pDOMqNGZaYPPpMXunRiXvAqhpo54jwJdEXM
pbm4aV4QHF6S7yIg/nExzKMQTppe208JoxU5JYHxnGXdMryRpbgZKl8bNa/HOdkV
YdXioxfYvukCGALCvxJGILDJKbt9enQAaM5wYidopcwGBuTxWNRoL6lKPN+dujED
I9yWHrFxgqH/bxL6GMf0lMEikmJZdAOY3E1Lk/nqb6s09AGuzfb9rUUcrxjUbsJE
vsl0jhX9MFhxDV3aEf2emqnF26qaM1zH4V4g9HnTKWZnI0pcxw1ZN0PcS9DKqpAl
6KxwG+MS8iHYgYUj1T09PDtjVy/iX06SUPi8Ag0GjsnUIOt6sIEzqgqQYjYrm9qc
pOGUwqgtbKRg/pZVBU6NbiNreHo5yBNrStohjCGEHKma6SBJApfystO9rcNvup+o
+O1uy0xH3qZ0KPDRWnsxJs6j7uxZTN+9sxHYDiXBZjJlD9yfxtsBz1smJrzNqvXq
4OgmaayNcFfYCE5vSONH6ksQCteHh/x7zPR1hZkvATdGO3f/5ZwYwjx9OyJReDYN
9xkW1KBxq2aoqTz6R6MIhY6+yrEMatdj/H41KT3X2Bo7Exr/YfyqL6kqKpQwt3aq
52m/AjiSKsKOHvccJ4STxmtc3xn/l+UwQV+r/bgTfPB8c1SSqOqlbq1h25y272hC
ecJOhMGPxbamXhA1VwOAu4tMcX157+mVkiznYDuMBEc84qEgoIIeveSqQMdRnmXn
lCgSJSrkwUJuqF+JGiH+PhWGOspps3sI1ij/mmXXjQzXco+r0nNnXN0G1hKOvmD0
EJy10CZoxPGu2la6Yqtq833WVSnqKjF6xCZiKpGHGSrLdmVyti+cnTc9WikWEpIj
YEIDOe5EuSrytI+kTXupzh09FN0KGJXfAdnQs4tNPF8lPrIrBZ91sQeLcr02geL2
K4Vo+gaF0gb7ezC0caSv3m3f/vS2Bh9sCKRHvdf1LDzxviDQnJUoLYeE5CjWs9Rs
+7YYTUaQHtvpwWkkmly7RNGDkFmrKP/50ehAvLcZF983FTNrvsz2tkMviTIrFIAc
3/nrgclv6FBkVjqJ2VN9NcbuGZrN250QpNPi8qxTj0ivzMlDKyVdlb0wdLvnZcjf
+uj0mr2opwrxxZRMdjSB6j73es7iykEjxc2/GqY9N80cePvDRtRu3fvISS+7lJVF
Ry8LKGi0ioHDG7FaXDrqMHwE5PLQ+UahK5fXE5UrhYg10EAQW6E3BDYMiJ2vYrPt
ZltfWl4f4JnTPUO8dePYrZbqg2ZDMxWq9hhfb/WgT9b+Fa83sbOSHR19JRjP97xq
QLDt5lwcdWLsNws3lLlEjI9UTm15hxIJnmkoAdz+Xt6eFgDtnqIx4dhUDPC1rBIJ
hRW2RHXwG6xG2EZlRfRqCWJnbvdaCcg5yRFMJmW4q9jvoZLXAABbA+CvwjA9bkLN
9+J91WIjUdJMqeEToC6gvdT3tJt0d1iMwaKLc042Ax2QDwNfoVmY+HM3bSX2QBmZ
S/rVZBmKuIY/VdHfMfC1cVssJ4JzqlUhbGMni/4L721c951S4DnNJCDXOwZIHKs6
6ee3Bzh/9wEGCirDroQA9S9U6KLlujHZvuop4ceL6eTJaodQqFNrohSAvbYVFWIe
qVU2rlXNypNHNtAjQ0IdDQPGHfzzJ6VaR+55uDvTAB6kUneI4ebJEkNnPf20hMJu
jnfmNy0mraOFDELlKIsRq0kh/1pbtj3ELs7oSZVaWSmloutoC3V7iCF08EuT7Tod
WdbWSGRPEfl+C2zBFL7JGPN+mO1QkPKRDSJA5co39qwqvo1ug5v3/MNPdyASUPBg
CAc1XEJhnBAN97mHzBLxpgpH9t2wyMaqhU9nF0iB2f2ba0qWjeOjt5mB5c9BKTLz
fyaKDPDdJ61KeFtNjbEsJ8HYCeJTV8/I540Ji0vC22VL5Dajf4BMVutAi7UqCQzF
b45L6R0PHxigmPPSsksb+pow5VQ1NHKMS5Ih/zlo4B4RFTQnoGopQGKfuRdRwwIW
GfNni+KCZyG2gRNRNFsWTWD2jt6VGbiW7IAJxAxoA8E2/cDCaRRTaTxj4xhxX6Iy
97GLWoU0JEctG3J4thBs6oLhn2vbyC0LMmP7coULw/YTbiHpBsuaSrK7r1DZXpqS
7ALWUCoyUJrkkUbjYp8A0r4VDJQp4bWw0iWp/ODOLQ4n3RmCuscKPhMy3Mcbkbc2
yYfnWqIeComcSt43+yj2rIr79+Ybw/deGSLRI/KSu1jw8hsT4OFUL07r0zO02EV6
mDSfttJ+jxnn0tnGIdUSfOhSgk8ekIAbGywreLadoLYq+CzQFUnEGdrdEG7RJ4pW
8KLI5WP3AqJbMBXYss7HpAnHgMgO64citySjUwW7CnDU2ww5RoPbckeLZYii5mJx
N0IbtwfHl1kJ3bX4aSzxb1ZtZD/bvNiss3iXPZdhr4wlwnewwGLCkcI9+JYsjc4b
7UiTLroPOGc5h+sKcNDkQlLqKsGm+105l4h9cx43vD1/vpVv0OgYOE7BRyLW+sfK
E7IAmxYFv5kQOq4rsmgSED5HRQbDPnTQRwyF1mdxeJ5pdnAFb+0P4t0Uk2nGcvyM
Qer3wHpORzjolpcTVojhqWgvUC+DUJwru9WWZzjdAg9+cZ6nc9LA8496EtqF2N0/
OVI5QdMZTX3lZwrWgtVXmku/m+QCm42jRLleSlMZh8Qwzi1DsR6iClxPBYrOYxZ/
4T2cMAYRdOVN4dGr6eIieC/Y2RFzPKqKHZCn/jI7qkKprPfa/W768CJ1lkI63YWb
/su7Wnx+Qh93I4GpbIzSjqBiIhO7ayvetueLlQ24JTS3G0FWqItbKyoGLMP2/9X7
O0v4z3KccKvzk1VPvE0xz0i9KzY+m9Sgq4iEwuv1QuRnp3FkzNoqqRqpPPDGDZUp
NcF6nCgV3d4HBqspsKg0chCzgedVsh6vVIbWvtO42nRhe2Z0jNGoScqiBlfoRzKO
jty6cH9sRSrS6fzo53NvcrnTrUYhe+TPM9Ysx39Kdft8nsO6iX4uakiFTJ69zRuI
AVEPLCICIyxvO0rT+9ujBbq1nnKItu7I5c+w/iS7qPzALY11ICSSiEgdYn9zANTk
IRxBduRHpvhcHUENriwDS7COZboT/+GNx83ukGYHyiDUcZQgRsOx9uDfZGCr/AgY
BDEJhagvKOpPeLZd9XB6IguMJkXBdRNXfhUPPHRd81/N2IS6q/S3BOWw44DZeOFC
Btm6+ktxDStasSuaxvMizbDGqW2azAiruNaNnpR8esXWLV8StqjFZ1WlQ60qp0Un
LDOt6KPczik3ElAb40vlGOxKLe44H/UBwAknKvbiFlOz/+7g1ezTeEzUKEFUA0Z6
tmG3YJgtSXna/f3B/2E/X+F6Jq3jrhU2De3DLZl8numyCDS0zMsOQHooin2PXpSb
v9U6svn3+Gqi48DrG0E3FUYGtbIQcS//phjlBP2tQvXJHcu1/VWuuvvZBhoInY9S
Y1/1ulYuO33nh0kPxGOGZvpaC5b86iao1jXj3wsoeLX+vRryrwBEGELPrqjCv0nw
0NeHSB598mikzOk5taOnVNgLr2HTf+gLxYF8CoR9Uf4upqE9YAtyS0YBwtn0Pn9a
x380AG5ROgLIDXH6BSYdcLqQmkb2/ZN6BZGZ5rr7I+2qhB7PMhXr+4SXos4hs+eM
BA/G83r26tq/9559o7rp5P+KOlynfAFJ26dOZavZqLXHBuIY2y+vQnxR3teLzrp5
wXC0fQiJdjzZCh+n8Br4Lvq4yrck8OHgaAqyTn54xOt3hr7lAFXyL8WSz+jBq0FG
50RlJE/0rHWGL5yoRZESK8+ny4pF8ASUOSmFKy9lk5wDYmeE8fkxC+ypi3DHCQBb
zwqZAZaATOK0zqpo07z+4V+swvd+qGvVkdB7FM5NFbjanCui1JqWHoghDaY+8Uik
5eVZGcVWhUm8rGjnQ7usoVCYbaTsRsXLAIK8VdIsPOyMjILz4QwUHNA9vgHDqV35
zV+a57R9nwiN4zrOT0Hk6u3S7uUC7oQZQz9nC5JlWQBIS7hGg7MZdlEGRTveUdXe
ZPV7otMTEzTclUa4eC+jXyQxci8P+z6HqJlj9r9E5tG5PxfKnCyBGv8gkxxIbYj9
KnxDAjI1t+KN6ambeovaBkR+r+9CmcLOI38n+0JXACRKqMJqhndKOmV7NvsPlZqH
+WnGUv51IRGZ6ljh48j9AVr8CLqKmiEej2Nq1vdBOc/Vpmp2CuEjuUSidyrmlbX9
qJoRerdMUcRRCPUCp3CevWiMLhs7Oj7/CSDrtdKgLYbdCl4ccWWEkNRPNAfUbn4c
qbJ4p2gXPMBMorVhD7x+26Q5ytCJqJnjMjRIGsmn3SockstTv3cO9d6F91Zc28E3
BGY1wBKN/8B26+w6a1GfpQJpo3r+/V2uM0j7LBU2mI8WbrVx4Sl7cxhi5zzN4gFq
+tqbR/bd5JRadfpM4GEHzpD+ZUMbp8d9wPMaPbLWgjCr7iBn3kMI5K8e1a+7PZk9
yTRh+zcYCN+rnPPEjuCtQIqVVGfLF8IHUv9dM8h5KpYQGshtdOuU+HNnXD8495fd
BPdBlUZyYpYLz2PQ3PKCnJKYILkPjdyEkYHbUXXO0ExZJn4aHH/IXGYfE06QOQdW
5maYzwcCy1SklB9AEVBJzTU/Y1Q8EWns8aG8qBRCwMqOTFyi23jpAa1Uaa2hTn9G
r7b0id/9SdZ6tzsfHj4bPD8reoS1EUJ60uu9E8+D2LzcTHkJTP4CVf0QkXRJlh+i
r3lqpoFEIh4z6YE/j9xAcMIsEEeO3soGGGho3p482Z9brqgbN7rUVJ6eFcXjngO/
6a0PTdrBWUOfEJ00r1qs1YQPeRlI5z6AZweFNsZPXqIQfz7MLShTYhOq+ys6+rQw
E+tO5NygtKMIaM6Y6ZjsBU0KfDVf6q4fYXoeCmBd48N7Jh3AjMD3jOao2MEN3nDF
4N/O382edzi2WowwbQwaP3Z6HUnHiVkgocLazsZhB6afrVjujx/bzOTkkAEVLUvb
xRhOjKVvbnRbml1SfUmABYnhGVplf6HfPyWeg2alk6wlf1ujxfROC/96K1FzwgyM
oC6vXn7daFt2ATJAzv+VnxxIq+HfFNP5e7KuTc11jDOBywKj5jF9iMrPBoGLd9d9
v2Hug9adAtLs1peSS3I7PdjsFo/utPvnUJ8hXgIuXpxKOxIk6RX1eVy4fLIvnW2V
Pbv57j3soRweTNli9SrPwJu6Dm9+zA3jHWAvSVVr2A5NXu6SdHFVfmxcRMsymQM4
aL2M3jYDoRqnFL2y9VD6LjZkbDFWXbtr5WP0miy8Sd5ywqXvwATpQxMV86EnbzAQ
Htl5e60xLX+tQtcf/ji2uzuChvIRbqVPmNAsSbcFg4fO79ld/cxZD8la1wJbwu3O
XrdjkyKy7MY1CD4iGpNJetWYOBqMUBOVgmrD3NLSVHw3M1uVPs6fZ1NVc2VXAcED
QhCzVnFm3l+wEdpQ5Hp0cv0Ztrnytnzc5h+oeHFh7Or+pDjwEems+iagyPk0CiCU
dO4nAXr5+jtU4u92iRlmmXLL00Akrva8FgxBXlxALOLc4veQGLX9BPcT38BUsLqk
z2EE/VfGX+LFF3JWnS1lEr8rdpJjdFIFJmxqZvezQNcavj10Wrv7aHYnAGOpYMYW
bFWs7JSdFBFG7Dd3saoXVA4uvOiYP9VoOy8sQFWJHtQOyBto+ADtIUX53dle1yRJ
Hnldx9oeEbTZ0f366FXy73lnj3qmkWji5H34OuqG8RnRUJO6ltjuvNjvjBKT2N9b
NUqWlLL/nabABiIF4FhkpEKEmn/rOJYmL5Cz4UiBf/FsJN/FSqam4AyvbPEz3gMP
52qm916DlE7paKFG/t64e7YydKFo9eBkIu3kLTSZklQXPFifIEbWkkaDebGsTDR4
tfM7tFYES9kV2E/WMzZGs52fZLl03vN0JrMhpQnNjFT8Spiqyd6OBVJqdtk+epFB
azYpZwGC1UPl9Js5nOb5qRRGCzvxHBOTh+ARzOjiUox4J6X0i9h6MUoWIsZw0+sv
8LnbbehgaI/FBybkAnk1jL5/1F8ak7nIkbOFkmRB45nvC6rAVQyBKcBxa05QDsxs
6ts+fI2/OIr602c2hjb/QMHeTl7BSOqyVlEtq4xr8YMgozGU80grw2FwRtbbRFWT
KGkSVc4KuRLWMVgrhw6RuDbw8Q/ukFCKJZH1jSE4kbnoMJOb8fYMgeGVy90szv0J
f8ckejXspUiP51Ai3g9DLEBwgOpG5C2o5oQDDhaJl4glVoyvsmkNp+ZHoOMXHS7b
BWgdlvmTM6snO5288AUcbViR++GgMpTIMFAPxC5bGgJjOtQNdl2oD0X6mM+2pfXU
OhM8UU8g+v8/Tw48DqngH6ep0cEU48MrnZh0brEmBMdqALMZ+jq3HFf2Exv76hbt
sy4sW9AQJitbFbXnbPYwt+BQ+NJGEf7Evi0xkQIh+ltQZ64YJzhhzNQgjzhiyWHl
o1YncMCicW0Il3X6H/5tWtj9DCvWwhUfzHOlPAyf4cqoV6p/FDq3ScRvJb9AyDhP
XdYzqatkaH1Amj5ofN4eVEUydR6cipmGUQ8QHG8FwvteJ/qyDZN2mKJp1GvrPkkz
+J7ByQcJEnG6vMd7ip1J4bVzwqMCH/iPcXdboCvRq82gLsx3O4sagrtrfQMO9S4A
A3fFp/d5RjteJTGlf8bbo0VZqgSHv7v2U+CU4vY85+7xvUzrqJTnKUhOJjvminTY
mVpaGr5e87nn2sEwkco6u9ZGvfoOP8VOcU4+jYTfiVZVcW3tinbgWhHafV16K3SG
tWeiiTiJSi4vdClznMt4HpuS/Eg6fq0pSgZDsUP6zo/YRPu2f1b2Zh2vS9zKx/To
T5P5BlMExwwLtOYx03sadNciev2spEeFsepW9n7HbfVkrAoLAStlUEDVEocFagjD
CkttqaP6MzVP8l+i2t//m2zHsosPJUmLwG61x6UAbfurLmounThPtMbXfmDMGVi2
rve1EXIcR9A98uS2WMqxhyNHqUaKMrcW4JeH/udkR/5D2YXh1vxLHGNRmEbfMxx0
+ptAcHcSXfv0165Azx+6wFU91FP6xdF5v7//b+V2ytZZhwF0+8eXOjhUEkX9MXFK
OvGPLdZEeXyl/p4tjGo56k02UMpBGTfA0nlKqkoPhLatZPprfYIxGsFcpWLXRlgA
Y9yDHoeGqmbarJ9bRUl5IINaYtc6wQjv6G+e9bTH4V0LsTTNocjttf+dFFHPUv4E
zLgH/Mcz+2xFATH5W51A5d6/KGp67IQddXSS3J8f3WW5fu4glZySNsHk7mHiix63
PyMkGWobjNAPTl0aNPKR4M7415GpKkgyfGiMlN4Rl/PEWCp4jXIRPIAdEfyfT5LV
6/atkF7JSYPvAAZrC3og6C4hTzquL2+j4MyIWkhZ8YNceYOsQIfrPhDftPWN66/e
6m2BVMC4b0Q+xSjdMshjT8klFzYJrL7OYa8JrTRNwurbRwNLpoMxphe7tRTGLAh4
8p9vQfqdu6ClYZL5ZSMSXneW2wzQ+tbYadDtJyId8saqVxMBVJ9JxMkeyAo/q9HX
jgNQik127M1JfWpHuU1rbfypmfwcXWmRW1TrZ+yod2GRjYyZhsGlomMscvQV2Bm3
HRlYfV4CoxCCEseyvhOolR2VHtYfeVx/xBVZL/91/tZYeyBV348U6vZnDic+Ts1U
E2LOTcexP8wBr8mLMyWJo7CSybrlgNdaZhd6Dgm3E07RnmoqGBM/wnm0VC//13O9
qxhB5r92q3GaD65VK0x1L9eySN5nbAqzsarm7eFD6LMxd3cJ6vf0B7InybFWr78N
tMC8docHbGbgCrzhY0mgwEROaotHb8TvIFkLoYiKsQBbpGET221KfTHqm47KTYnX
YUWwTeDzHBq4U3J3sSAun3ZoG5aXcGiWedkX/kSO0Q/3xILH/DBN2Cjyd8FlssqJ
iYA8nuY114ZGy44sGA/Z6FGbVTcv1RP/EGURob9Vdprj+vPZh5L2PB0INndpTfjy
W4W7Vgq3ZWOU1Omxio5vdSiUzudmgEgMnwcyYYx8e6nwePyQhlzvm6hg67v5iGBd
wFBl8SwKGvQu2VK4NSHhTLXfQeD6T0bLh38q+vVBNgWIZq6nKyYGoV9eJsTtScyY
Cs4DQTZTkjkhYfQpwq2wHRhsT50jwjdJECihIUybi7pxYEdf/ndXvIVn89X2gfNj
QZoHANaKfA5eegGkhvQmvkHdkvXBOfMG9dBFoDP1tRTsi9CkiYXjfWv3EMiYErM1
XLuMBbTd7k52ACjfJwMxnvKibyylYAfezyB7nNNjHD/r9HjxETC2ydiFWHxXmXgE
aCeb5iHEyA4usKFCwqY/U5ooCQF3nTcrgr8h21TghMplkXAdbt5wclqoi8H61CD+
1g3L8RcJeXQu5fOsqQX0AwfbSbHgcoKmLnEY6eU8qU3z30mbfpqxB1/hXRYzYjBG
0vf3LObWUDelVpm7Zk+IuRbaLQoWhcZEJv1SMtHgwQyvGvoQFP/uvK/Lh4BuLYzj
BgypHI1gjuf4NDriMnCizbYfDoZKRlGs7ghi3CYrRrsoxAIGqk/L7XF/HM99BlWV
0G5jc35mFFnL0YLg0R04ar+hEA5no/p4A0zAJaxQyM08qyridCwxzHYnRSNubpYv
bGtQ8wZGz/QYZnpCz0dnn1BsNetC8GEAxMIC4sZSp7nMV14TX+TKK97V2yD1rTDE
8MOb4muBq+W3P8eqrU498Ql8vkg6Pi6nz/zAknGe1C+nrbnLjFP/JEeJiLbtNi3r
LKqQwu0G3wOnoabVAkNXkjKZivNHTHCWcuYPr1VjgsVZ75q7MSh7Z8CaUOwXQSmL
yrdpmh6fYaf4z1w0uJQhA2YDAjn0wLJ8XnAQskySeLkXp9JdgOPzCozGKLafE/ho
+Zii0SPAh3jElerurOp0S/LtG8LUrOogfKMmzDTuf+b+XV5p5BqMl8B5Dsry6VUi
ddRbK7NNmhnibVdkiAlmyeH1C3R+k1aKUjhuuQ6e7RF9ASgeMtlLP+DnkpN6audA
317BLDF54+QbNxTByRjCWlcrtIk8gD4+yIUqDt+0qpnhYZIUNmdC6B15/rOyCbwD
cZ6CskTK0w1Q6SwtQWBDc/LIjJeoH2XbbATDM48Hdpm338NoHpwO6EW4DoZoynvv
3fSo5wpq702u1xJFo3+r0L8Qs560W5jMuDQETDN2k2CoXtmTJy4EoBPxkF+FDFVc
HgDD5UiV1aduE1SL7A0+HkkW4TOG7OuK642/tLm5yEvsz12OAivUnvaipgHr+KK7
i6wPMUeYf5JAEGIvsL9u1KpaEPM4bh2amvDyWZC8SURPJXF6NzHSI4ltjjf5vE9a
GiRfxGvPPB2AaJrHK9TAj/r0YlbSvQ0aNiC9nJyj9zIwDO1y/NXTC2uL0nd6Vl6M
OrINylwqNiTrAaBqmlRG/4FQu5SNDTxbnVcrsu4K0uzOi+0gnYq/GrZrE9VHPM1i
3Q1VdOQKFQj4F6J4hkbsr9d1NpdP8yGIYJOsO/SnRjZiKCCrOfNf9F2va313AVvf
h7AujqgaXNcWV6fnxy0B82eFQ6Td0uowhvtuCllZf0uaNBC4df3ulsV5YCcA8D/b
w77+zgF3T5j8mroSBNMxT4Op96h7tQJWOxrFBAf5CU+/ZmtwFnrRJI22G8Zg/74w
2LisQc2wKRwjrLTpG8/QbiDac3de2iOQ8b/lu83+VHdPuTTM+LNe05rDTujw4Pgi
6Ole2ifgJiEuZ5cUW9n2qz/oKBk4XdoNbLF7lLOYNYQITjTGFRVMyBNZQD8/C3Zj
vxXY0jkJPHov+3cjir6IaI+GjpjNzdlYdRJoBECwmqYccyZLX2nm6kyNgIOQhC6a
2WvqNBIm2Nm8w+P0qkgNrFFXfeNH9/5Yw9+8uQfmW/FjPZEkjmH4G38BL0HN3sWJ
xjj6drnfqSVmer35mMr6VnEZFxjbCG7CZ83IzESIWAfLgJ3ImfuOXFWn/STO/E3X
fYLPj+F0o5LM5ihY5F1Ohfteu/fOT8unN43OIDQ5PnSkgE+cB+2NEfpjNzMCCVur
rvHMHflg4aOu7ZTTufg3EClp3E5M7WDIATFep39VfMmL1njXHipY495IKOZVw9Qk
xdLJO4Qw7VJo8ATloeET3VhMwNYeTZ4klKSWOL5xAr6y1VbOoQxW1nw5RFlOMiQG
HFxGFjSke0Cy84FSa5O1XsxSjhx651svUAU6y1i0XY3NrawViMNoziERevvzmtuq
BMM7L+mE8hFS9csmko9zImlmjnjd3+NUiHmKDCVwsMlwtiqBrttx7tLHNYWemPtN
6MIi7uWn//B4btoB6afs9OqIppOXv3QpWf343O1FhYyKEQ2aUQj5v36D1FOMZbAY
lIpmp2LYkXql9ASmai76hlDJYykqzyH8zn9HW1342WPieZVPN5cvY8uFx9YSpyhi
RF9hZBnNifYTHBLgYOXkeSorHE91qoIHjniqnDb8EI2fZUgDyz0LG8bHmtyzIuhA
SQphdf4KVDbsS4KuMARXc3rASFR7I/8aqrw192hU06GbOFtkCHQEAqosAxqNttbO
C0l9qC98o48bvUUt30gFllNUJLWbWoNHjATrdeFR2M5NEU9Kqj9qzRbKtl98ZQcT
V08UwVRlWCVctIg0OWxcGAAtElnqpjf93lRbWLyU5JIBA7xZh9Rn5eGvMzEwDE6D
u+AwIY3/9fwxQzxg7P2jqTlT4lmoxBYF9QArQPe43tIuLSra4ZCSXP1xuqK3R1uL
bWXxrBivCv4wU6ULA4jfqyR7Z/6ysTHD7HjFKH7mUqM3SzD7+BRdTOHRsCV63dHn
ETCRCb3AiRPwSFuT6D4eYeT2ny3mWp5pJp2jcPFRhzKeMnnR2P+6SYoe6GtP43gx
Elxvf8m+6K+d6HssjXurY0zwCOXgkA/yQv9g/lonxeq72DAIof132ATTi2EfIIyK
7TyKPyQoTRkeNoW03aG5ugeLjb5wwejiprQ5QmyCM2T3nmzhz5nz0m0aS3TpBUv8
XQiDFEmuczNZeeWF3SmteU6R7jJjrkbLf7QNpLXJdD2+3rounhWd26Q4oxUALtIk
DpxGUaptg3FYoJ4qv2mb2x74iRoZb8vtpkL6U/vvlW2zXTp4W9dAI7Ro/rK8TUUA
hbWX34GKW6xWLz8qa1gKKsEH+qAbDfOewEePiNlnmQeeF46vefIBJJ+R6s6ZmUdp
JiiR8RDHCV4xN9RCgASei4nWGsB+mUNqAbAMm6Fus4A1InJ7dSoL1ONbkeX3ksgc
Y3kyc8MhrbWHRMU3BqIYFmZ61QbVJkySfju8F5RrGeq5WUXRBcH/36HCaluJc/dk
xbgev9WwoosObSl3OBuh05bPabdhOQPaXmqyZN1Mg+4YjYE+Edk4nSRHT6kwfF8+
NOkrBK1PACdo24PsrRHmCGy1ltq4daufQgRqS6g1P6+ZTXiBARL1OjstPfnq+l35
HRgeh+nKhtyEuO00Y6eiuGyQ9vZ3u/I8uINHJnfBgYZdYJdaLcpwIckip5VmtoQ/
f/MBUyus/tuOPoIkaf17NBtGRwvBN9dNfbc3jjvw3R1amTBcaqqcUlw28oneBOpf
O/PkrE+9su7BeB2LqFne5F+Hp4ezKHR922Aqb7Gcr6hzyY0RGANjwC/unyW87SKa
t6eCkttWnT4Rqe388UhVvUjLvQ/9FWUyPOMuxMHzG2MDLwsAZSfTbPHQG5JYHwIi
dZpQZRR5Qz7TCKWo0JpDDRaNP4sBKhtnsXVmUNZw27ACCKx3jjb/2H3O6qPB7nwI
ssEyCk2DnKyZknGxjI2sYxQWped2HgeR52cuoz/m+90gCAXZ5I+EIRPcjoAzJowU
KTU1qmScltV7C0TXKWdcHFMqcA3TInTiGoXCrhv9EIj4BhhAPnP+LevbNm+ZWO5a
gdFQYLsv4ewDxzUtp5bHf4ZvSa3xwtfE32KwtBadreprHu+Vni4RRJGr+bv4laTs
XTvnBZdDkPivgLsaGbcLAFIn6QU6jAjwy2PgTGOyFWPebZZm8WN0rLHMgyolaxk1
vB9nCERrUQieHV5C8L6O6nsBh6IWtT0wdmcVPnySnlQ1HZ5N/OU6R4qwU/JpLD90
GAqBI/kEdUsfCo1HVgPUNoR2s3cMNA7C6TDm2UvZc07C7obM6Sy7tZ9RYmU6Q5XR
HA6lxmPKdX9aKPtlVDzesdCGiZwQOHu+BhJsKNWcCDLovXNv5seQSgOd7COv44dH
0d8I/H6q3XfbalGu/P37lmfGXUsP1bMSaF1wfYAHlbrhC3trlZ47T74tBp+RwkBS
eS7OJYadn4BlwtWozD72xE1AjnQ4rjR/J4KyHQrDklsvqJ76JMjlavK3g5QmXb36
xgETtBEr16kphTC8ktoyJuTPLvmjxvF3hmhzWLVLXx7l+ork9WE8DvkEHOCzLyCB
tgqev4RQ607ZIHbntooYo797OZhgx39FegFVYzKMJM/C7+6JdvQCh1/BvpSNsV+B
TPgZxr46efg4qNcvF3kDMxE0w2VFRtAg+vd2mTSki2BnNMPIDlhwePpiyrAXWnLG
Pth+F2hKwYw3H2h+bY90HK4TUrhlr1hqzbl75cBC9zFfoLExrXoHDvcSI1VnUHQm
6x4s2uCZoJ/9+2zYEl9KC16rqHv3mtq1nfvSCF5bjRrwsmO6WbEQVyH4r6fVutvX
6/HA61BPGhcXgkZg8I6Q+LrvRBpvG0fS8Jm2J9FMyFQXEHJrvUrN8lTroxZZgSQd
c047LPgp990+KFJDrqalqbWaT10JJO9xR78Qvlhla5DE7syHtz6oNKC4eRfSZeFP
0dgszazAyUoRuO1Snd5oSi+NxM+JCbG0HmoS1TFvevQo3PR8RDTug930QiSzcvjb
MR76WGsL4GfGIw4M+Ne1MQ0/nZOTXRNDsKiC3umITA3+Q283qMmofXsj0seEwd1x
d2PHV1a8C2vICZ0S5vKY6F3QlLM3wYv7q46p1y3Xg+mFPr5fXOO1ZutkDFag/qIB
PXRKCVIFepA7+G9+2G0/93Vfq8QjGloXtw+WS5rmu10cp3PRkQ4kwj+oo5KL1hJK
eNUZL6EBCMmZ4BQvK5+mVTPJyOJQHeGwbl/6NEcopvySJJjF07y1Pn46CaWDV8e/
Mkk0+PWwTp6l9ErN1koaCP6mWtNh8fUCleNuK+1CVD9RkxMSPg0OBGAIhhbagj3M
UE86UvB4egsBv+tZykkFaPV/OAvaqxcIcDOVmC2tHBgN2Vr+hHcxHdc2yFV3biH0
T9JC8+rW8fjog4OF0/mDqfhwICbHJe/gHuXAVbj6S6xy+hB7T9dz0kE2wq/OatGX
URn4mvHJPtoLJh8+evrJ0h7VfDj/uBQqp7N7Vhko6OM5Xh8RbuE9NAHciNpem4rp
v0u6Ii4ZyfhOqVBoJSN69neGqn3h8P1Uq6zTtOVvEqlj3sQtpvQWzigO1lyzF3SB
X7bJaD61CxAUy1SBgKFH0GR7M+mESF/9fpetbwr+SAXWcZJViseIYy7qJEvXXvYW
K65+5yOQO8H4odYek3ecek/rPOo2YQ4umiN9awhAQB0jdFm9r71v+cX3WY8Ybu/T
ckKi3B2p0UpSgnSd/eDjq3/rMq6Ou6ydVaLzJQuQ8SUCWiNPZjnEu6rA4sZGONdB
WDz49Xruhj6p4FvfEpmuOpmqWFUf81yN5IavJLwEA0LKLjzxYMRjZBNLNVbTlMmS
3VGkZ1WbSOrW7cSs7fREtZgIv77JUnlyxSRrrcYhbzVnSvM8IQw30KrtznHCapPy
ocSrYd2S7LqtikAgkr8tgR/rGAsXn5qsGTKzfT9CIco+GujxdcOrEYf0EPilmTW7
ONjxZZ51U6LzeRUJBG4nXh+KOymbWB2HCuxZqtYrFfqC3FHu86XAerP/Zihxc73N
M7cJNu7rk0iqGmicHBjKywwEC5xreICCH2abAhzp3vBX3fwyEUk23s38+wjQXVCi
CzVunGvmDG673IaMSv4veAelAsKroNLI+n2OpNV8uRLTmbZauNmy7vHKxvwB/Ncl
nOJ7y2HcqoBRB03mM9E7TPJDeqfofBdFJ0viuCBy/fl+pxgsfjoxQIM8/egp2qwY
5ZfRPIgBFDVn98NmX6xuUNBBs2xKLrKAG8HOVH6OynXRC2XUNoK22l+qZbkX+7VW
svYbpwZiAZKv79bNHeIAoz8Vfr6G76vVaAoXOBNJ+s/UELSbX4E6/PlRTJDqO2BI
pQfEgGsUxRiW2F8MrHX6/gsTV6llzDG3OQTmJ2bsp10UF3giK8M4o89SsxcpqaIG
tidqT9affxwCHw76Rf1YoqyFEV2Ljbp/S2md4W+7x1cz5sLRhCNgvvjbSH9bU8Bc
wP1ww2C2lCR71Z9jndvjPx/q4KGUsfAA/DxtEZsU9Uvgiix36pRQYUumCd3a1PbJ
PaoLcWg4VEkC76AIt7+hQRr8h5c/rjPPPhOKCyt08xwXtZVn9DF56EGkUOsOrawK
dC+0iPZt+04hGE5+LRysSGtiGFaImfbE/wDRItSTrTmls9gP56hFIa1+DMreAoRc
65m+REw9z2KbF4RPGcZIqo+dkrNXpbS9247H4MP+GiWlcZ+/UbVo2CvgoJP7K1vY
0j8bUcC2QGDsl5Tqkkt+uDDoFNv9qgbXgwIRy6Bb/csdjkbZyODjQMxrne49ujR6
Wr8f+xcDU9WODIiaubOpFnPcyWZv93F+jXc9kReqhM1gpixQqq7+8KaZhNyno9WH
vQuy+K7jWqqaqNeW1bKF0K9j/nuotQ+XjnP2lQkYOfQrCNg6Dw0hoEjSkdmJxe6E
LFRLnEZ6YRR/KpThimZG36NeU/PSz8sy2x1C2Psyqoe1v/JXkAOO7jlstba+wBXC
ckV12JzYRuNqniz/ElxBBTKv16SFy1vlSafY62isHoX49eJWySslVpJefGjUhcES
XDffWyGEXhhl1ddkSL6JUdVKyRoyn/m7ga7mf+xcj5G7lJBVY4j+qpBTOXrsl/nU
kKAiSXvcS73+OHmkAos/32og48SZmbEdeNgTwboDFMJ562LHYPsGwmK7LygcBX/M
XUl6mIt/Bg1Lr3swvQALcOyCld50k6EOZUp222uQ6E61zVDQCE42RizAQRU+aVb9
y4Iu4I5VIzuapTPWKLwdz1ebS9AWdlqwbfxoYlRvOxY67mwfWvQzM+fMZyV8CVce
45JQvbewK1uX5jZI2ifU7XjSjQ1/JzdSbOBfESMtn/J+6dK0cSmN4fVQVQCFcIyE
DSAs1s3ib2ZI+WMapy3sE1W3z3EBuWOdoMPesql8ruj5+FBotJHMJpHGfd8yrB/D
9m06DPX9dXfkhoYiBwMN4/4mufqPfPmcCHiuGMC7VuGAA4B5Gmo5LSBwGiVIHPtb
kWy/dyFyBjWekp+sXCWqh8HlYwe8EDnzkaf6VpbRrNXnAsQ2/XNg/hQbjmOiNN/R
QHDaPwzaDtUIB8NOcsz59Dd0CUZIuPg6nBI23yTpPtprQidXnaWO4g28Nnl8iBYC
X/9AWrnt6ADjemYYuAKo7o0JhDWVCRNPc9uM3t4NZ8yvg0r6PXpYZV8rSsOpQzi6
fg83pQdLphQpyCViZi0VRX1GmgaMuN2VcR4JQv11qooHBUixbFMZ9WUFGsErG034
nTIH64ehl9Aws82W3hyDgCQ0Rb50s9n7+B5XVKcwXBHcfvkE3+o1YxgjnSxxXgbO
FAC55c/2WsQX0a5o/jua422CNUZNB7qplQrRHiwybGw8117rwyRohdeeP4Mca+oc
lu2D6KgLNAqQLHzWRWWMGMr4thPA/xYP/zJn6/NCh29VEQr87h2zhljaMpKSKHGP
ztEyp6HT20uZwDYK3Jq0feakUm2kU/q1moAcTkb1LHW3lDvLS24QZR6jH+LrjpOQ
tVnHdNyD06XBeweHoNwBqT1szsH/2vI5NkyvJthCO1CJv2rAwT7JFOj/Wyo5akqR
375GZvQoopA4SboLmmcVOl8lESaU6iWtuQp13EC3YBrKBuk/GpI8nDje6saEtj4l
js/Ru2zzOikcdlf5y/WCUz8V9ohZcTmeAUHwgL4XPpup8KoKqezJOfg2ERuRvEkx
OWRhq3XK6tP0NzS1WhzBk9yMLPDpAk29pXkwKsy8I912RhKT/ue1t6WydkG2CZ1A
wZJHF2JCK1OuMXIQUxpbXQ6+gEUB6TibVbk3f+xGGoDHvqSCYeCSsIA3kx9UDyFs
2fGf9gstbnlSilFzJtSpYYBQqw3bY9aI4ntdEks7dWoElfSuOM9AwegtDuIL6OGu
BwwhMfxGrgAWUDEHQDmfCX7cwJKw/83wJUStuxWMQaDV44m7vCnuW9z6VXoQXaKs
7jUqRnqzDFksRwMPb6IYT/LOpILcUd4d9Nvo31Xp4FMoaMWVlIyP6S0OqrS1rOG2
/G3qvoovlDS1/cXlNU2stbjkMW7ZEAFF5Fv/HbSEuCqX4yzza2A9J7wgjP4Rgkip
ZIYKK69p73miJl31iEAzonOZp+3eWpKN2ZKGZPBi8witk7LhiVlKz0haUFNmi90o
xX7Pa34iWVC+fYzUBz47G7rEMFaZ1BpW/fAr9/Fl353nxf7nkmeu19zc1T3n3JDU
xAGyyhRsiQqVoucayrTq8g3NIG3v7wf+eW20mddBEymL2fytMqz/BlivtWOXDnDs
gt6KB7uQpIwY2ZmRt+y980K3YMcRuWRQUpzHntTtW72TGux3AhaB6xWVnF95cay+
pDQ11s7lIRwQZink0cSg/QHF0/I5EQGvzdnykzWLH+0wb1G2sDTAdT87czQ1QJe7
rIHdlTisYmcHU8LblrqIIULmjR3HVzMg8E6PPVTvzwYDJP4sUx18RhPdhII5H+aY
XyDHmoCGZKBHwVmfmvdut9J8PspYWIAjH5QFV3rSBvDAPZRNAxvTb/hHc9WYNC8w
GJGYZGPTa3Q9zW1Eodf+G1NNO7KxW1ltWfB7R0pzh0ioJoxpsf0pzTT9vABZNZ1y
yhPJ8jIooL2ROvDyRexjXU2UJ7/J/oC9SQvS0neLf3d4P3mZ7ujM9M0PJs8oGSpd
CDDPdyjo01jB5JnVxLx4qEbjGxrXNqQPlOFvbtoGQrKSnwg7sZS/ba8HqfcqPjdF
Uq0YMCFaj4DeW6uPVUji5ILtBQGpeFGOjD/cwmfkQFMRQz4dR11is5X7v2k8y2zk
sNPVfXvefIxcKIvJudFgOOYWNTdpy6q3C3wscxDiLWs8y7vJbDcq+jpEN0qubw0R
v7jZCvFoLekcfs/AMmFm3FU5ecJ61DMA0UOwwxgPYZOc74kbTabUocrHepmL4qkf
VQ3lqaocS3EdHl7I8T3YoKx4VaYbPSW8uNy4zk43DBNuIwBeMwuRIceEriF+q9yb
3iRiu83BMNPWpCJEprcrMaq6eef3BDNrjX+wbx7dZQGbGTEp4EjwL8YgtzbusmL/
DteHULz6NSvZcUnEXJHskOmeayNUn7ZnsRQs1ZhWYbkO3bx3gztfZ7n2WyEgL8Sc
uyvzNxajeP5npTHPe4c7HROjOXoGdlNnyZWIfu8kV4dswZ3/R/+pruv9+Uf+PvzK
fVPyTS5IgzI8Kg6Z22BpVmORVdIYFOj4EILIvCgx/uhzR19Ml0BMWxoXeGN5S3ck
hGBESPJLgCKiktpUPFHnB+l2r3DEZVT+9izlEl8aYuZ6FzSCZ69hvKEAsTiIHH1c
OcK6fIXKjPVgN9Juz3gYueURzeRj7ojgZeoSD2+Yvpojs9/ZGdXA1MxdpSWLzooA
q6np5FM8Cd0Tz9uWMvA7S9Q1IvitiIDqza48ZNLutmm45dQmXgy6yKUTmPiCqxIk
lp4ZWWXje+UT+3bbSgAFlFURVN6M73KzNDlcAZaj9Rru0JRL/+w7avMTcGpS65FY
UwSL5k2lunqYtfBhzvSdrBh/1VYeikrxhitspX2/ZAiJqi9YNkNlZ8bpl49hotG4
zd9o6qFVaF4Pj4KNciWP/qIz/t8sJ3gZhC+bzoHIdYGFs+34S1/Fw0UHEpOcVwON
134i4/okvoalz25vQmc0pKTLz2QfqopTNMsRycbOegaJRxMDHciCaG6OIQeu/jNC
mDodjyk5HNlSlPEIOedBygXZ68jodOZZQmoHvnbU7g5HQE+dcbDT3AVrj+h1z+SN
Genu3Po0wX16PsJuIRZdqJhTNrkbHZm7KqYdmGJ7kFPHdbPh/Fkrfw+TwoQaKRl5
eizpacW02hCeHrWbuURHGP8u6WEQbdyIDby0Rs07ikFw1LFtSdL2BVBWgj4UL95e
pFNuZxmQl0UOPn+LpOBk2U9RKH/SOId76AdWFwJ1HE/8rauhQM0gGU+4iRktqu5J
SOd0tbTaavlR12E5jvb8RB2bUnBTHxEQO8WX5TjmoOmb82w01osw9badkjcmyBTp
saFqbK/N+45lWbE7JhJcs4Hc3AEQJ1cvh6DeQRfgI9GFLjjP44rxsp39jlPAHdEP
D7F17YlqvXQkLNBRVNdGJdzfsBZA+sdztN3ZLrTJHcNz1DqHCVCbo5Zzq+VdEUrh
NdNYDuZqUwHx1gCM0Jo3/1n35BVX8Zk8f8f9iABxXJtieBTb/ZSipQ7Mn8B8uoUI
KWWXiSMsy3Gq9HxzpA7Dq5LT4cXtdz6E5Y2re4dtqDTV37hvmb1UXQ47xJINoDYj
j8FM8MpCWx+BqU6hEW63e7bWtGhz+wgwcYP5CL76WGHmRE8SbDhq0qKD5yyZVWS/
ToX8o8d5sXRUhUbteG7qOMjASHoBxuXQPJmwPY9Q9PDhqCmRs85Da13k2qSuE7dY
KzgFBlVAUuPspmfbh9ad31d75INL3f3GP2YFLrgyRBFVNAF3Axd3VxnbMdjeoPCy
4ANk5FiU/NLFkJYRjkd0bpfe97cONfdE1+9WPmSh1+fQKgvdrJxw66o/KMT1ya8b
AuOuWcEVzyJ+4FzGYnysj35lVai3E78lRvjeQnlqyPK01EuYsKMvj1+4TarFZAMj
GLCRv0FWM4nGtTloNzyOTfwKMOsv3ZlfXfXELUvYx1PbLOLrRYIB4Lu5QzqWdkFI
JsAf/jKklsIAZgIKlwWlLaznPdlthK/YaYI6pLabuDi5XmVjBuxPtDDUnxBw2M+j
A4jgp4ZrSclWPdXQtrOlnLSGqpIg5R3PvvjQaUDPZhf/2pHn9r8lL861bUg9H7gh
MdahnftdyhW7cpP6AePNJQt4d2qDp9SY6PHpBza/IlfsVvhi/i9hoOfen4wpqVmA
zhMxGMFThuK45koJ+L9Ln1JkkAumnSeDz5BN0CiqaT9MR38j/xzPDwGLfq07LXu5
5qtBc/4X5damg/7SzCTxHstzW+04shGOWrdN4On1kEhW9aAIRsd06wnxnDdyHEB+
ksjo1b9Ul7bSA+jRdwMcem5gMSN+nUcwQ8u+SqhiOCmS1mNDRZyTn3taSamaDQ83
52t95TPdx+9qC0rWGR/gmqQi8IYW4NPiPOCCWe4cc+QQzdQO60dozBcyHiYZNG3K
MzKK1lb8bZTNSR3N9LUhe60Y7un3Y49s/Rsee27U4UkZ2cN8DYSzO/hGS0VJX0RP
TsPOUetDP5NPzr8sXRx0jOGS43pM6lnAUqT9bMQjZVFi2Nq/2xcYmTzr0t3nyXP4
TjLO58RFr/oz5ecxewXnG0p0DIMddBEzirdNt29rL5gHtlbEF8Vklk4xwGT0xvIj
FWmv6B3ke4JYcIJo6XV3Cu5xrJo3KSiiEJ0fXD4SDgjUwONmlgaiCf8jEB52IsBW
FTsqw+oG8ilbXxRWhNYGUMS6wY9HUAQ8ruDVQPs5Nzhc7AKbG5ZI9eDmtH3LnZ5j
NPCaP3DhbwegysUmAwXytq28FpS8qZTZsoraaEiByPsh+YxVE50gubi0nwXiFyH1
P9HsLf9grjRExY519a9rixKj3pKJ/l7xEgaXGQwZHMyIiJnc1Gve9pn+QDpKNZdC
ADjNWZwogFKpB8VAfyqiU0XZWApW8CWULiodA2RWxf4n/ndpWp0+jU7IgClD33Sn
55cZ3j4649HCVIjYO1hWPK1PfAX/fVKu4w1cXWJ3O2LJNmip1lhmx6nR+ESYswLw
1hBI0uWGi7DQHB8JeoL4GluiI8QjwZpwux8yk9e3/CsxJ+USWtV9TIz/f2W8/dM4
YQIVGeU95Y8+6GqJ4pgWy6WlxPhwabXxe7mSNm8JAw3/7SXNJBnuBuZm0JFcuo6I
/1FtRQM/OuwbCJNPcYfTty5OuOzmw5X3HPS+hRWjZ97nvZ6hTp+SU9wuuarkjMJu
ob8yyumey0VaxJ11zffHbugnLtBQvu5lZU6mSqcFScmDz/+H8zJKpOheLEXp31xz
hNwCdRIQZxAOO7YW/X7Lc21bOUTY6xMG4YHAoAQV7PeLv2q6oFeyiydLa3GuXblz
PgaFsuUiCWkS0gLsAJzsP2PyMGZXI72kOzzn+XuKE3Gm3QCOZ7lTTUeVWfnb7zUW
q/gNc5nM8BFvFbiILZ7+jNFuppgYNzkmqkM/rkqVpJ0DGcoIIdehjlMup0JeJJHa
v41F3GtNZ2tPkOGBdBHUOagJD+iaAau2q3pU/zceY3OuvgSh5qZqpD6Zxz1uEnEn
sTHn5rKHw9GTNSwPwQPQdLLlSiemwEqLhOtTHufFDfM+C1c4Y6S/UnVUlj5Rnn2l
dpxCu8OnaaNckPWOp8z5eeE2CAJIuTnFrElko+ItAScbAwduvHw9gKQx88EEI2pw
RyaEjCOPekdEUTZsxxid60+Yu7/SO8+qgVEdz81EP/8auHBh1F95Hdoy5111JeBl
x9azwSaNyUoSEkjxarJOa03Ryxc4vBvkLOU9PvbGoyBw9eE8D5CtImniJ5FAIyOa
NsexNNgjuB0YfEjcWa4BILL40890Qd7wteQZDVwuLHwXJE8eh2dq5mX7U38nvmgq
FPInFHnTrozydyRfZCeY2dhlDzoZ0kd1bbWJlfxQs+cm2msiAEx47qxip2rDfuam
aLBfBwy+iNmUpi5vg/HCXTreCGXX5hZohrw++UBRC3wIjxbBRIimuDt1BnasClNv
YoIFchXTTjSMCSHvMrOQ0F9Yk1Tm4oxK+VfL6RS2m7/Ozih65pj/q1bZQ6/mrjlP
NGEzi22+NWHwt6CW2HsyeJkxB4Ff/triSGaowQNNw2FV1j4l5yaGsDDHGntKPDjS
+Y3dzEajGwGM5eq0dTMikOkCxZdyY/lpHoZLCUJKqUY1DdK8TarmIqTPe4ylMPef
i8cNzmLXAJRFUKLhDNhzKdXNB1O85mIZy1LOxL3V07UMqrbHBsD1rX7DHHH5dkG/
T69/gDzV51nyc0W7dEDoIBvcJlN3f77xlp/gdRjiLtI3PyvoQ13yCj53eo3KshpH
MramDxGGsOvNFViRYro6KrYIUzU0eaQFTVkS6cHqFg9zWMrWJJKjW8C3MB7bwPsu
rIuENSb5E3ebOOaUI2nVcOs//SDdpHYepl6IqPDqpATYGglwha2Zag4UipPKe12A
+4LcCMauJMJaf5rOSDQE7W0w7qkoq0s+4P/ZQPhup1mFUT6FnjCEjTNnfNDnMzYk
nxCSeiCtSuyh2flcbUM7MTwL9aHM5mnrgWmtodIU+RJ0d8NKv0FYqa3Rz4AHkR2g
jocK+4LrpqUxi8Ly1novESGNesBkFdDCPniaOaONhFGXfHjTf+mYudVeTkpczAth
CnGHiRFT7zmMN8fFHshH65ByokkqdgEMpJYJR5DKmfrAHuW18r+lo2gnSDSCZ7vS
8wF24yz/l/uDu5MguIzfI6CEEImOUWTsLYEmcg2tgoZMDVDJJLO3e44qYWoWCWC8
dP/+EeN+B5aWcDU906qKoTBGUdn5H+p80I9HEVKmrmnkaS4b05wVPxMTvKdkzupB
XR3itvHLL9mWcoNl5W8XrgXMo65fYaL18wUHu15V0N/B+2UOSoHx36+SkSJD37uE
Gqhc5Qj21hyhKxOF2cLpBTrA+LMyr31ttlsWP5XgaB5FjEG7/mSByuco9KugzsML
BkxsE8WzfB2WLJJ8k2fId1lOrADPq+GFU1RnizZmNmVx0k3Y3ERvZXeUU/wpsHna
V7Uz85rg3P+2SXGghsOaqfvdUOeeSO5RPg8ZbEhoaJqmOJwH0wpyx+bE/wGZB1wF
wYxM+aomnwa1Llt5bRPKSQZnO2akjIwizPIUFx7mpd3GzY6XUNgOgUn42MunwFFk
pzF2QDTIIxuw2Nqx4UidKuE4JkP6hh8JnV05XZ4ZatWq9endnaBmTMpxZAeQt1qO
TMTKZtibJyu0rW8reFqBPMyXTxpx4NgSJtvpRazHlZoPCJlE5+hNYpeBO6WjLflA
dlrQMl5fzvqSkwHJiQodkA1jeTbd+WRGbkrieV91PIrIdvLbB1+FVDXK76MC91rR
t8+Qk/8m5scJbsji2LyTWgi4x+sHh6//fQPM7hnuvKPbqz2H9ZOEjSZYPkMqWmwE
PLX/seEQcjdMgoiMlOCVGB4jH+wUJBuF67RdnWAqwceeY1Rkz/OlNyrIpCdwDgtM
3mgbs7Er1jAoapcTSFV73MhqQ/B2nploUcLUJDyCxJb4yhHnjfzx4oMgRJfw3EH1
A7RKgGsP0CM18zvkNgt61zd0LkCYccILeRFuu11P6BEHwy1h3pxPHYkg5PdfOmZn
O5VE5z66XHkaQLY+vqTLHSkwtGX5KZ2pKW+9UTGGIFvc+svQxvhEPG9DKcWQxzZb
MYmu6VPqoZS2FU5qZ/BC1S+vOHhX28iO4TuQRSgLtXTIHwAfO4KNh9Ccmof1nfU6
NowxweqBdJKBcfZW2oB/RaUgPEa17fEhPJ22EUHbxROIpVWnoqc8SoNEm+Hmkfyl
1d4DvdAWVBXkFse4q/ecuXBuiA2SXfCwArf4hVYZGm3KxVQ5ivE96cNhpaiYSFtG
DczsPfMb7WpmmP5osJ01QRMfmfuOYIABnuH9weBi/kt9WL6eT+nVfARGLDHahS2t
7W/+Z7nwTwJ074zeJEWVik/2Y26McdM+xEUBM42XRg7TXa42xNThp1ro6gbOuepv
QfcowdfrvsirITTbick9HUdrXu9I4mZg8Bkg4ZII5F/x8Nejbw1ccuLkMcWuodsa
w31+Q6yFvdcfNwGcfobzdRvtzNTwm+hSpr0opfIm616IiDYpIZ3TAUM4IGs6knq0
LIGrB3dfCEwYeTvTJxECZiWe9aVlt6fdmwSvu4IS6xrb57JePTwumuYUpi2q/+GR
x94fbqrgVbijuK0EYJv6xeQlgl+epnwD5N70T3+9MF/8meuK5dnGpS3nTMIDzXeb
ZmXWNCo4u9Zp1z8MT0PPX6fh0Ob2aJKwJ2VUK1M081N7LEyjsaBJ10pKl8IBk2cP
Pt2h+zTQZnAjMjP7wP/1mDlZh2n32dbMFWNlrzLDN8HPtrOwGFnlc+aPvOmbQzh8
a27GnNXxuZYGR+ppK5ZV50TtCrtIXkavgZ3aa2iSyTNz3Q7bDEHQ+5y7iqh4poJ5
DTfNk0+B8wQfw35KDJbP6SlT4FH6Y0jqr/cImyCenph6NQx4pc+FlfWfejqLOTK3
qE8CuPsBcDDZEk3cf6Cs6W0zD+zsRoyp0YOCsTL+72HHgM30UnKljCq6yoKtb+ig
7I9RlBuplwuJOiUKLhZ97wslHTEycfoXTx7wf6KM02Ki4sZ+Rwjz1UJk1DBZ2aLF
67abgtEH00xfQUxCh0bPzFET+MtR4wv6NHHyG+NZEQmIsBCIFARKWJjz/RDGIW/V
E3w2Wz9JQB5y3H+sKlptr+MYrrauYmTAsJBUNOKVYD4Vypu67C6h+ujmEnAiNvzM
B/m6GnW1g3eRxW6gUvBSHzxJ9Wc6EkI49vBmSB1/oxdFMbiYzro35uZIi3BB5UNx
+shgMi3DuFeBGov9lmY54VFbJkPcuMvnsuSsU+/+qy42Im2zTJYm1qH7DnInrDJo
rPts0kiu1pEZkw0OVBGik5UWE90otwXHSJKq7+C69vFgSfxzMJ+6ffNILECf/oKq
AcvlmrK8zMlUwQxtp8NJC6Tbt//YUU9ynIe9tauoVP3tS0wlMDonfCHPrKYfUvOZ
GGbxPWqmsaSF4XsQFAktnhB/II0jL2J9obzzEVq4IaLJE28PRTU8JBH1jS0TKYO7
wCTE7mL8LnzNwVF0v5o7d049UiFyKBAwXXhUc7J3XprIppLWMvqlvcD8nAtEwaNJ
yp9ednDpgGc/HKTxX1rE8/Sgz9vVvdy8EI2yXP3v4TUGTEqH/ZzAUuKwBr+Va6+0
RsAf41yWXWQcI49qUP/ttggT5Fcls9X+CQYbbn7mymTG2zcZGlxrz29NqFUWhLow
v4ULTdCZyC1h7k7mhs6619VE1KwOB8440A1JC/JPbXz6B69Sq5Wz6Pzi7DWs4NOA
t2M5MzMJSpmbyh7icIyfkY2zeN5JdJWJgKqzJ6DzeSbboocARFYVMiAH9X4xH6iK
GKOEbftS3ZJtM07YrXh+9dESSnPVnuZ5QvFX40cha24MvyHoXG6WfNKFQCIpbsET
lqe+D59MdHW+vwaR4VUnGnT2kQ/uoAQgNMBuo2aRRzAD06n0DbHv1Ab9XZR3KvE6
Ud1Eabvf7IVx/ElOMWuHFg4R4UK3jpFg7JBEwMAOyTE3y6TUfEWjzxbul4N2cNO9
+aGzr/dOlS5//p+9HCYdSQkC6SYVcbmGyNW/+zYuHnqCdJp/vpyuUG30uak2QlOz
0Ngw5PIEpLKEv6N5vA9YdOHmJ+RFuw7GXPwHcvbLzMUY+r/F5084u4AB9yZuMSd+
rgb9GsHsO6bV7Rkas8Xi/liYY7oXWHGOn7YmeXoTGiRdPbVyOqx7WWNbb9L6/5il
t//xdffw73tctWl3/2cXsa6rKS8XgkuDBIplyQf/x90l1s50AHt/2By+pk5dxwA6
R2PV6fQg5BKU2z+Qb1lLiQ5PA1e+ycsXNi7yKKVhH67Nnf4VsXntqOwvYGRfT12l
YcCJkJyVQ9FXAxGgj2zpu/QiG5qFvcOequscGGkNdoShMRFM06Jf5AAS0nvVaVU5
0z7RTZUMIeZXFK10Ew8bzsgaQX746Mm6zkXa3jvuxK4ALdPmLsj0zGUkyQDT+snq
uQ0I0Q3oTfkInxz+eNQ8CZ8ANoNi5mdF74Q6Dyekb5gTV26gS1DyYlU4F/o6b56j
zuaW0w5oEFtB+ubC2lp+fzwO2t1OAXk3KWR97sy+ZlgLk/wdjC1allfk4JEMGbuY
YYHOqkTTWaAjpJeiTb6E6GkVB3gwSLCrasFlEMHpt+zFRnGdxi2AglLi2mPaqzrG
EJfLHGWg6mcIx9FoAejcdeqDc2USbUl6RsbX+v2/znKTMFMIYG48jJeYlUiOtwlU
iVk+iw49E60liNjiKgG/iRp6LAygdychTQPdfUEdLf7N5+HnJKTowG3C4kqTKuU0
YZeaVq+IpJhjDlA58lvlP9/nuODzE7HbC8n84AnT/k7pCUKDCbABJQ6NPLWj5TPs
al3/5fJTpzL1jxdaaahDpmveBXpRp+eR++bkV1dZJOYGfBlOTFsHNSU8ccLeyC+6
9xIp9O/2T0ZAzRTLTWOJSKjiLp9JiUTbZZ6lNW4ZexuvksySHttbxD4iPoXQlWqo
Pa06iML2pwY1r/crc5ay1IYSMJCA03YN3LR4kprKcCJJj5SrbW0e8rO8ygf3OXda
YUJpb43RPz3kUjbn/xxjZqk0nUl1bT+wB/zhTJSiPZxyPAmIqg5KBgkJljFIEl7V
BGXe8BDkZK5fh+x0mVX2ZcfY97PCT6ktSrvzrIKRjTaIx857tDtyjaQzj5CL6nqt
+M4DPU99QwF0wlEURr5tVukKixMYO5ND1GCZR+o/w57d3uMBvEU2eHKZ16pOTK7L
iiPN0cA7xkzJSiAImVn6ssNZJElgM5UexQYSweJYW8DpxOu0raPvK1I/CIW0lrG1
TSqR//6AsNl1Udraz0priHaR1Bz6lKm8RuLvSdFmWrzJAhQ/wBpG7HDIA8Z21Ilr
0WoFOKMHQsAcHPfOKAjsHQjcVGx1YRK6MjIF+eYtim6/zThJGFRtFNg80Y6m6/MS
Aflz3S1LS3sss13UiIR+zt0sHtvm5snf70Aj7p92MuCEiYbkNEt04lgQcLHqKySG
SpMRaJl0BzKursBy/w75taPWEoHTi7o9hV8KV786ppJM4Pj23JsjjvPoOzuq35UO
srNj4T3uLJfQTYfg/Dm2fEBch1RBonYPiS/ZCWqGLd+KencJcl7q8h06rlXZOoHa
vLVD9HQEmDJleL7iTmN5TfB2k+MePn1T+BmxeFAdvGld4w7jN6a3tK5OVtFvctic
zePA0bfZ+QnWZUv4026TwTaMU0pw5p3sradmbBetOD76m5rg7nCEVO6UAtuH6E7B
+KqhlGWIhM21XaO3TN3EAYZbOYPn99P4KRjetE/WLpW13E7coxeuV5dYomz7+J3r
Kgtxa99BPj5YlxGJFG8mJpBfikSH482Pk47kNw5B6kbeubm3r8H2fwV0gnV1H+RU
RuKQN2EifxOW4gT5mXZjd4kPbqbFWgmRYGLS/4WxYmz/jhw5wDylK+xYw6axyCW0
yyAzROhnPtxBs8gKfk5XUQhL/Fo3I2YAICm//mNPd1uDkP/SMkjFs2kUQKzuQfOz
/JDS0xxPK8303vF0y5x4gx6tUIXc/SZyiJoFCWeLfg6+1vQOedXeEMC1rOARatZH
5246Zj1y+NoPfYtlTu2+n+S3FYui5ZzeoiCZGS+OoAOP0sjdKyAQVC4jUOmPTJ3W
asJisKIip1g7Gc0RJFLeq7pEmo4kVxIBr3JBqVKe5wtWONo5JlHbuQUCHVvTfYIZ
UmysumGPubyqZP0A0Vqe8XRULZC3lv8S7kvpQU+e35K1mgC/6Dc0N7FuYtsi2oTG
vaQunl6mYlRhELCSVTGKd8iHqAg0SH/1LOAQJeW+dOYHFADoR2bEYgVBcsTUwEPg
gifRu687JeEkonMUOyYJn2+C4swtcOnWkUgxg/qjsM6TRkOn7mDqaA+TI8DSY+LH
m9ogCog8rAdm2fF9ZC+7eA+cdsT3RZRjtr4pKQBhUU2BvaoniN4ittaUaok2KgY+
vL8JsQuZEXpJ2hMDrk07Irs/8ajPlKSKAGJRjHTPPHil/GlS5DNe4yXL692lNwbY
Kj0+M+ctEQWeRbGAGm0a79phjsPHK+xWx4qL9hjJ7+tee+/nYNO2zckznxf4q4TH
KadoMBRKPC9XicceenCOGgeUoSxcVtH3UrfskIyV7Eo64xl9eO5J5CuirR+kyW2T
nntNWu7yfURo+TrOdFvoDrZUKxPYZYK8VvkPf7AquHj4YAbDdYXS+QyHAO1F0nJc
CYZigInBrT9oD5i/3pwAwGS3GSxmkv4WJ62aVZuWZiNRI0W/kXrfWmdSS73yI+Dh
uKw5JC31dZAGoSArwUyJPQVA5cUoHFRE7/2GoanFzLY3JcNacaGcjqig+Et5tRGI
vEoiq9NL1U6BCHmiJSUrawyFHXvSqhjGCSddF5qCKfFNN3SEljazB+6jnWuj93mq
0dnidTAyE75/bSErONMd/IIWOc/CtP/puWHiyebQV6+qtXoRYkfuNX2KN0PFQW/7
PXwAM0tnPSeCMfO0EwqxD5J1Id0ficRsctCQ5ThFVQuymev6XOmzt0BYU8DskU1g
Lbh+pPbPogkSpmf3t5hd9Bi9YkLL2rL5Wc/fyOng0o2GY4waIPSLKd0sWEc4XnlJ
0lJPAKRhdT7WpUUQoT9gad6Oa0sTA2X2lBSnoUQeb1XEw+x30aYTpkruRkyAcIRS
ED+xwupnB0AU+HNdMdOntjHCxpPcYKOYdlp5/TIgbL2nw61Tw9TRDWViipWzNxyd
9ErUaTq63HAehkpoz69jA7pO1Lt3wFF3cGSfex8xiha/tqAmEfh89dHg7AYstLVP
jyI+iUnR1CPbj73Zo6N72K8Cy+0u8xpgciLbfgW3HAMds0AHDxXlIOyPz9H9yGIl
9JYxL6dsDPFkf4oUuARlImeUn0UIKvx9rFQTTN+42g6j0e2LOW6Hv/slZw42+FnG
nQuOT+SUMme1/vZRU6PRW0arpdLhuh0I7UiH2xzy23NxfkqiFsq7qykVSov2KS+9
cbBAy79cvumYUYyH8eDVqmH8kerF6BPvVgMC+z5G1PSXH/5+1tVpOoDez98/DtUo
QD3xAgnzjx/4BVEgiAmlItXWvRAb7rGybapcNcAmLUOkrXMStQridT32PxPdGjAz
9iYElWIfy8oISdbDBDDamsylO/I4g4Z5swK5LoS1h/i4HyIec5b5r9PGmphF/0OL
7ZeiXzd6xmQmAz57oyM6UWdGO5pFxV2xP9xievjfEKvpDhX9PTAtufmf2OraJcsK
0Rv6KJugHyE8BSVCIEh2SNiFbYw21h7Z3jFM5CSoBllPrwMOrTj3ht8lULRdZb8U
HowD/lawbtjmI1w8jIX4rsWcdJB4SoTV+aK3VeqbnBugCn/45tbZ9vCEmQIQ+jNg
1ttvYcXMD4BcKPc786TX2tR+QcATVjhDFrai3bwy39qfH1QPEnX8vFqI09PiAUiL
0ftA2mmUlPZcWeDPn0Aa36NGdE98ZPtzvPJ9HY/jrJAwSLANEl1GNnladBHZdVFk
9UrwkJv+tkfYBs880RxkUdKxV5MjZg9pk7aG/CZmQuLK6a5+m20wITrEEuEcVZAB
H1jOWxChSBBZ/+KG1wPdlTbZZkDGhK0qDMyvtDzyUI8cSgw/qoQh225HsAuJc5+o
F3LQQVd8x14pfo2LUavrFpmW8iZNM4XJ/Va1gLSlo2t1GYPcm0DYwiNa6ncO07A/
9oilWnTkIrZ0qs881iLcA5evwKocZPcmQ0xn3sacp6kkUI9WmVYow6V5kGTeOjH0
RRsSdpMLM0ZtxULKHRYjS8N5Akbl2U7o1EWIKaqzAC4fslYtoCB/YaH6YIf2/gVi
qOavyevO+j6n3Ja/i5tCv1o54DFkEbt9jR470wImVHIVpJeqYxwpqS9BBjwnqA5o
9ai7LhFukDvnCrj0rmhaMO/oeQbtr3kxdVZ7TMo6sdwLpZYUNIAVFwShBIc1rX4z
VvqHqoETZjAWfGNstwr98pJYyEcnWESJP8uj1If6T2/fEPXc0Z7Lo+PWVPhD3KsP
BRK0zRd5mEfoJROir/9eNmBvW49hMuM0QR/VhJitohvSBmjSCs6IfGPx3u5R8T/e
ye3udYBaYy7t0U0ae0M2LkAhYwxE42X3N31CI34FcC3dQemAWA7UTwElzK2jB7BG
+V9zChLKHPYomU0PLuYmKHVkdhJpTxUooIC19YKg3Di7lvOFh2WLCMuWiG9i1SU0
HDw7cKuOiJcDPIfekXjK5RWJclbwIjK44g8rXJKjlhpxPO9jguL91/2eGG54mOLg
cDDhqnNKs+zDrh85FZHsAZfTq9Um812bj1HQpo1RuNCcDBBE+ASyRDxduOf47E4J
//i1hEgj4CQxZHlw0X+ho1WJvXCDeF4HxwZyTM9m14uIl9wIt6yLbXUoJp8Rk4Rk
3Ea9CikafoHo+anaq2comsvrVAs7ZB8Ndjdgsf4usj72GwpWGXE9l09NQS/3oBwH
rBAGw2mKe14FKMjUJH27qN3xnR0roIrZjBi3S8Rxo+jjK9Eu2JClAaUP3RogQdJ7
wGh4nafQtpPgFb7FJL7v7izzXazZFjGnOjjsRKc7rOauozCfBJHXjCgFViN71o9K
sFfxRcWdbs/G6jnHUfb7R7cNKOrSeTpqnvgi6bZl72v2uGaFvNqyodGyLMoxB8Zj
KnLcQvYsf6CxwJhrFoHRRCjep4FhTQBQTi+2EPmg1Du2irdkZ6bSfOYVhCvk09bN
fkgrdnk7ZT/tzyQcphTiOFrX00i7kaYCvJ5cGhU4ClHmsUTZbOvA64IOv4CtTELs
r91zhGrJcfsKb22xT4qmQjULplYASnQUkOJha4JPfLjx0aO9Pfe+6T11ZFAsNLwN
rcBGk9NuWG10nOJQNa6t9pMQDZ5OI5h2qcMzh0PLgq4P1tH5/QXn8IGtX4BlGHlb
SAaI4IKrKCL8k8n/mDEoW/IcKDerO1c4G6AejEwhVSPhApj1kT53iFb4SNctVYSn
8NDXTKr9lifkLg8WPnJM0BB+jOyRNY/jemDXvxyQ6ZSeEMU6BKiUnwZGk5AZHANn
RQAMjnKVtjPCsbd+AOLfEPwifX7FwBPCuGm+P3hQrC2Rs9TaGrg41moIF9tTe1J5
KPiluqegdOuGuEZuOAidkwdHdvB/hja5oBxLn6owV2KuD2VYNYs9ZQ+Wyx3btFvY
xRmPB+Yx/ka5VvU7C/stSLcaoJgPoF/w7/rFUS5H70NGxQfkNba4rJ+LXCBW5P5c
8sXJ2jTaCdXYLZZZCA1HdW7/pNiHZdbmEB3TZK9X/ZXfVuNLaXuoRXfa6muiz+gp
1U3jmUt2JFVzEpKwf91rsDTKE4ljwM68xOM4LTR8afZPkxBWa9o++iAKxU0RII0L
1xEFQk6IYCNwyR9MlA1C+knzrmwlnf4CnUttut6p0KyzK5XREJOVLyzMfqdEKPOc
qhohFTKK3VDIMEU6s0VccEyavSS5J2YB7rQVtJwPOhvYXyIMAIlBP7Ljw9sjFUCv
5dyop8RQn30N+VneCbGKvG2JGn21zmD55eQmhw4pH16jNAWsB4ZqBwSQZocrbhf2
mYMrr2aV9JWAkNihoiqXaUXFBy5LrGYCOCZatSRyNHa3X2G+NutEmS7vkiIsCwqU
AJP1/sd9Df51rnbVPOY3+/r93wK/3rL9ZcCpFn8NuIJz2Xv5nbB2+LcnhvpzQMgY
9sf9reNMxI213oUIuIYSt8HwYLeMFcgetJzz6YewKdi7L+f+0ggVw9wEbfq4zqCI
0oXyfBUvjX4gJnhGJCccuUTaKL3VNuoWj0RhIB/MCjsETPG4iGM+Tk6ja4+tZEGq
edoBGFY+h1GA3XWk75tXDEE4n8Ynnz0jpejY3sO3F03iRabeTM6VkDBBkeZAf2Rf
iqndrOSOuPVuKKnUokoHoKZTJn1SIQScSUz9vlUWSxJcnCrpDPbQJ8nZTiRWR0TO
Vf13HMixTRW/2LmA7vrgxfXJw3862ZR9c6S9C/NmX03QqG+1RFzVPkpWeHpQYTVn
yo0jUjo0NgAlHgCTrnF2eMQYivgv+jygQ89VXjHxz72HEk94ElxPkJJmShRs7gkR
0b3F1IX+EjD0wwbcbsfst1W034v4q2DcjLn1mDrWvP2L03LFwZ2F5lrYOnCZeqwF
xl/X1fYq1eFoPegEMzn7sPw5873Unji2ZipxgrNTzAeemXMp5kkDdPyYXrDlxQXn
CAI+Eip2xh5k5L+N610ty6d+AgipkGK/+jRx5j5yois9TU9JajUJKqikhj12H901
spIryNi0CYIS125+jxC3WH6BnVevhXWbq4f+9cClylbkB9VAwDhdJusdbAkVzgSZ
vwScithfx7iXQ7k7wf3yUfOAHvQH/BuA5At8OssLa7iNL3gcXxHXIdiquLvetiRc
AiyLnYcPJGWqQhJxu7L8wjt84Bt4jkTeeeUKLWl3f4PaLEJaq8bQ5ci8bIN0cDiu
5hQvkjf2Kiqe+0bNm8hJzsXs3czLFM4PQ8/oX4m3JWH9GrSyhIJyiZa7ydcgD9+2
Q49sBSd6PhXujvxJcTmfH8rbyrRFErw7E3XcMZBnC5aQYmx4ngmpJRq4eUNg68gr
Ngw+dId6DnuU77zAXdADQLoBTB7WcwyWLymxBcJDAuevUnOsL7gQoKcfsdfGY7lj
GQIdLmACt3rMS0o7Yr+rI3Yk0Yij2OFOVy74yKbcjneCNdE+hyjDg6w+/oaQxUue
YBJZ9vC6WN1GAa02ESX/ZhMRoIm78TBqkuq4YOG1DqstUIkwJibbCVdYciRKdI/d
xBBAZ4/GxOKxRJXhBCtGTGtlYq3YNu+MxAxkT5YPLWGzDwyVbc3X8qZEqsAmAxE/
dby5D2XjqpSus4mAq+7HPNfUPa66AhcrqXb3fp93qALF9Murtw96hYkKihBBYg6V
6InmK9EtavGCcNjQ/8ASqu7jIpepLNAzlqyi/cvE1NPdmQq6VzjVyakpaNP10VYa
4+4BBjFme6Db0QxLI/jgpBLxpi/e+qCLF/YsN6HQjS1XLJ8z7ymUCv+TVpAtuwll
4H453acvC7fRThTq9UvKng/tBpp7tlVgy2YoR/A9pqckXPkgAqydgr79UPSXS4+2
TheYI8VJsIbvZbbTXHi9sXp5CkAI821A7rJIj0r2Nwzr6xrTd9vUGhUI1dBiin03
gPtkEVpQNqsIpsSwAB1R2rP++EWH1ZisOSA0y3npfhaeHsZhADjtq2QVe9QlcYEG
1Gay2OLJ3htv36lLqKOu3UKp6P4k8pKtV6GiL46HE/6sAds6D4Kgqo5ZvSkMrzHf
8JzLnIStDzdCQhvweg+c/CA6+gc2EYQigSDZyt3rVHUFGq/IkWzR7/VAD1jIbFHL
NRvfiZiMpwx7oqr2b0oPkNItNALoNCxPJcBmwTJg5KdgwtDRLzZupkbLHjQBiN1u
5sXAb8LpQo0Yu70gnT6pnR+cy6S44MGvu2YppRtz6Bkuw42P9IrMyiY7azVSRUED
0ouQhZ78tChaXW1toil1fbgP7wcDk7bsABHwZ60GIY2Xje3LX3q7kKwCo7bod7VJ
qaq3ZibMxI5r62lWk5yRxWvLcFMtp11N9pMOsYnSuDenZd2EmvpxOW/00jVXpexJ
lE6DumfnSMKZFoVThlUuzd+WYumBl2OoOd731hxLmuVyMhEwppXy3N3X2DLaNXrc
x88j8+Sro7Exgwu5+zNdnKEnY27QzS1eaGGHETJ+Ve+3+kbSkTXPwTWUxglxLewi
wy4veZTuOB/eslKUCdFp+IbCNtgdj4lQWPiv6nTrogZb741KfZpc0IVgk1AeFwaM
/peLiATDFPXugt5phEg0nz5KexdGVjDpggzIk1HVzlrsEUYpbWNQTu/re0qRDpJD
NkJaZLWcqUGqsfAVPKXotu2GI8cQOAIFZKFwZiRiudSR8jQ/oNIp1aUDIclX7wCD
T6uU22a53RiTDlNQQ8Be8xIPgCpno5j2ExWyfpEoVQiwMKlmd2QWxGu/LGEbZxVt
GgrzxA67BWmHlABmACC57enau2TV3O70r+QEMglQrVILNNczhdcJHo5jhwz6OHaP
ZANcuB8TGTyENyF6HD5fpjR5ObH7E6G3zhNXXg+cNuKq7RDoDhSkjfWUucAnl6Fr
IoGoGvuAczNEkJyCzyZNXDQoLp0LavjcUxGg1cYHyUuu8293lhUms0nsCOc0S2qP
1iGEIic6rq510nhscnlLdiJqtJBO0chNQENHCSVx9zYxH+As9UuDh3b2JOHGfSgJ
n1JsVLkjKzcABCSU/lU6drgPTaStuhbxnky0092nYmDVhSOfZoaYzTUDmG/qd9Yz
Jd0EmXOTXIjErKJolIOMkCq5zvrKdrxRNHOJL5XHXILo/PaVh1kgdMWTFMhaHgP+
28ZVoseeTzZbeCvcVy/1n39sSme6lTj8b5DOrTFftp6Cu/gtMITHtZPR5oGhBim9
fnOn/qXLKN6qh6FY1WI5lko94giT4sJaY0BE8SwesYgzMiNoED4MyFwPgruUz9hI
cGfUmVBE2J/Fxe2z+bDYQNWnLpFrJjmrTo8NRRcQltBiDGmgGAG2vWGbqfHmr6/N
OGYXhmZeWs8Q5bVEgcN8FijW+fC8emtQicHBz137im2wzg2NlBCUnS0rUTUZuirb
bYZRrV33v0XERhNQ4eGN5hTtZ2i9vqz8CwfPrZBnOqNcRyPhEua2pJrDHsQyFUrJ
ODiJplUWSCNL37HGOe8PHNY+tnTzVO1nNab6zf2sixZId6yzNZ+NxMYdg78pb4yw
woWF7kpGO2fIV32shIAjtcctXErqf8wXNyt5tYizC9b6gRsHrDMA0xiR8bpYXWxr
S+hCWyWEFgrv2zi2NMUat1mN0dzWd5s9WsRTZGTeRU/AK100aY/9gAym9vtqbmPh
+KP3B0eiqmn+3KC6Ur5YW/yjccvWDDkWw65iGf9gNhlWzy/hkDvGW4aTlYrJ4/Fs
EzaZeczjRhEinoamPGtd4ApFlXugyQufs0PS4HMQEOfappgf08tgAO1M6fzIr4gA
mnogA/rz+ki+N0fIvfJ6WGA9B7WawQwsP3bmC/bF0N7cJGDSjyOxr5gAXy5lEOtJ
dnLW2LsbXYEN2afhaVwRazAMIQL89nB1KqY6jOCbUcwrtGuZ03qf1PAAzuilb2hM
tfaxncX5BcK/zxP1KJU1tSdbUiUyxw+JcKUuxGraIyNdMB1tSvo+258KSa1uHYHK
XA63w4fWWXBPOecVkTy5KsqrtWNjh69V2pak4yhgzi5vVs0m+Nl7AxyDX7c8Fm2m
AeqcajORMRUWOIr82nen06Y+jPibftaNOBw1niTFUvjjRr+FuqXYKj8Fo2HZlrHK
3rucyA5Ty48yaRXQv62FUPkCWF6VxasTv327kCAYSCVTnKNf4wOz86gJazNkX2va
SngFNj7xOlg+nBSIm4nGd3zOXN1wBU6XpuP+xxQMYLvgm7BRV1RlsEGj8f0Y7o6o
3JgxGeEriT85AaA2d7bbvyauqUOpKInGJmxodE/+7T00zoSky86zmkE9DXyQNvjK
p7R38RRvynHLlCUmdbOO/C4VsY5N7vEbiqKjN+0dBTuh401hMLK817KmalcuYIMo
+Xw7UaQO/qo1T95AzjXGL72DlVzjwqD9bqKkSIouiOszmX7thzGDVSX/g8w8s4sv
ZVfpOnlkw2AWTByIFWsCz8A0VIQBRz/hxxaKUXK8VryPoIQK7+rtfsrzOSjTnBYE
qU2iwbF07nB5p/j6tTFN7vy7Tjs6GTLKaM2WpDv8q+fB1a0KyD2H1u2a9WLEp2aT
wQKveWY/mrcbY0mG8387FSCkBAo45RAOB+mgem8a2edxm7cxYN7Em6PZtg+8YYIE
uysO4ZErUwuD73TR+O7WRCincg5pVmwAbE/R94EW9kZSmhJFAb7iZWC/w0JISxZ+
CeMClxOcxlwkX7/CYMc1uZCLTzjjIvDB7QF2nA+VW1wtSyPiK+8zmGqvsYhnuua2
Wn+LMrnwkqtd0SqTuiWqGM8ujDEm7CL3F42pjFvGoRexq3YYCWEwzez7f5/VjDKc
p4m9ZQCat2ghn0IEnLp8Na4v2iIk8OoZAZ8M/P5vigEVhJA+91DNU0FcRVVVd+iq
1PzuFr+ZQaKBnpC7IUKmCRB1qprNJm0vvt+SebgHbT2PdmEMoI9BjEHJYRw3bXGO
mIbwSbWMz+b9Nh9+zlIIPd78klxCyCgiPn73JAzLWeXieOWHRO565mN4IAZZepV3
DOnYRgowU9OBJc7jyxGcyh1XnmIDWLYfIfI89I8RMBgXvG3kYlGbWbnbxVA6BdRZ
tHoUpn20u8egwkL+HUwYb+R+c4R6yRRwJF93+LBvvWiNo0H12HRnV23fk7wizyoT
zCq5zlX6Oa3jLE/6FbqmHj+iqETw/wyZrwHO1MXP4M8yGE9imAuzQB+79QDrFrZE
nVmrSTo8eDA1Zq9VbL6rjohPtsHj0DxxcfwdmBX25cuHbYC67zCWz7ny79J6vTvu
YqnFoUbtfymYR7p/GlCff12XOWpopJCwiO48KF8xQsV4+1aKY+KQm1VqL+Mi1Pfm
ptzfL0Je0kF1LQJjhFqNFXdcFNgbII1GZw1CpoWOVJ0iXL4euZlME2Bj9JM6G0F6
+0llBogroE757cXmmP0a3VJAp3vGqojCWzA0i01vnJJpNP3oG/4GKUl+KfkWXTkl
SHoV8B5qzBGFzihKBHqgKJGc+FMm/bUx+oB6A3nV5SUUl7K4FxwQgGotLSlXxxfd
NPs9UIpU8OLHm5HIfpQOH7+xTETuf6Nm0Z2rImICZhGF7Q2eg2V4Y9GSpDSOCkHy
2/UKi/1MT5pGiItr09dIIx8+TGYL+rqmQB7rLtC+FTL5dL6guMwBkZ2IzVOdBL0C
eX8kMIO+/Dz/0x5Asa7GBdoLlkIxFfUqJkbDRsbGWxDACFfOz01VuwK9TFbHAdLb
NFFJrHRpKjTp9XUocAJmd3Vp4C97arpDZP1AiyaCZ/2e3s+sAIYjI6wFL/TAvDMH
SXWaoThcnnQpaS8jhkmNxTy//HytvOHwgmFxhZdMFViCyC79/OJxrL8lY97X6oyK
nSEC4td8Cz508qn8x4LwO362b1Rl3LSB0G6hPFQj/NIXSVZXqHp9OX2OlGP5UZow
KhwK6/z1b+zmdnAZ4w66o75w/2q/A015WXg+8I+qDsujcY9CgTyN13ttKNAYvpd8
I8PaCBln9OpXZ0+/xQ8Otw4HVOR1Y5f1kfnv7oF6LTwg6B6Tf/wv1BK4yvY0VhjA
Ywoudihgrf2pX/zJNKQrAVXRYmW1kW1h6L1G9x7SGvU5UN+h+ls8xqTMnX3olRUM
zNf+rK1ZRfScZhla+j3PF9ddqLeiSK0SQLaZgnjZ2/1A5/cbH/yafEKKTJePrDrZ
mGqGZjYU6yD/2W/1qCfimFRDQ0tE/+Jhw6agnd4bAyazO7paasUlJxxR0HOqea/A
GnIgdLGeAsjRBy/Yfh7xvDRuJHyvCnLwK1VqL5n1hWDsCCgMDJi29E2s3lo4Dd7j
e0ueQQCC92A6ZHbDtjRZYbHtRaFxusgRffYoCIV3L2FuQ/uHvdMftPsC0KEncUUy
cpWxZmXPw5lLyA8wWY27ToFoj97cWO4/rS+HsTlqC+qTElrWViM3+Sjp/4GSlWsm
lcGG1bBHM+JG6OwtsqcUE3xhukHTKgw9lZQ/2bIR6DosetAq57y1FbTi9QnoS0Gv
bvt18hOpY4jaD6JsfZN+9BzOI22bJCH2NGjTZI+K/W7qMt3hlHBqmx3OgHsYcy7v
fb4LnPyKQUEnk/HQeDGws0ybaxLzKL2CE/vbhv/lbb2aHUkNZ7jmcXlxLNpXs4PE
vXxTIeR9lxzvTHYabOuapyybBHJrSUDueCJaufhSzCo+af1xra/qxcopBA1izrqp
DR568yk0fUOj9Fld3WcOHQpRkGUnLqquZQ3+Z3C2YIhVVPqO/hjIaRup6KZDLgpd
VdBRRKGEUqiPTpPaxMnZOt8dGwiH2gJzxeQEl1sd+HViJPZJy5l81T0wiBKyW51d
naRGCS4kUzJXG+r0Mj3q8FrV1dmDvzGZ0crxnwVwfLOE/3jOsmm5Ur/eZ77DU0af
P3QcYvU7Q4QExChpUnguue84coSYmjMIwnewIowdwpfwqQsdI2rHxecfOk5yf1YW
L4sX7Afsa5ny6gpjKmh/Dm6jCE5bTq7WfV46GaZQAPGxoXoB2b8fDYyhKlTbNaqD
0Q8wl5fPV9aI4lpzAY+Qed2qEgv/jpkN5KYDPi6wwjjfo+hDk6IacjUJjWsAQ0Jc
9IH3Ymf7T/LtL/CvlMwcxkRyQCCyCWb/WvBVIwk/JG1IQt4tetfddU0E3BPLPHDp
3q9PMTUvk/hhCr1p/9ZCPSQ5x4WxGC/cSWWgAqJJNfIZGfTvpjUK8xWElCb1bGnB
v0KKvh2DowDylZYMkrax9oX8kkC5lCubGzPYjX9cMYyTfthI8G8gdGWx0j8QyEjy
mvnp/7w0qzMIO5FNa2NKmuuIOgZaBQghAat1qOGqal5Y1D1z27gX0Lr2Rrp/5pzp
YV9v21lEmUqhk8q/2q/demIpNVAHGzJKEbnJD/cOcx0x2NjlKfp52YDlQ6ag0B9c
Ik2RZxmJ7Ri7xQ/LDMXEjXYskHsssTFJ4HAvJOSojjCQXt1GIbFrMA4B+XGHG6Db
PwU2DmhJCSx22aOwEPuPKJPVyXKwvBPMAjyJ1cW16lGB9rnt46FPdgcTBpjYnkQw
OZ2RESN692VqR9KjKUMDumtHTTjMy9bqzYUJfFe8VvW1eN0uzid+oWIMkkTF7ITK
lE/p5ZS1EYaXjz9DcpqN6X8MRssnylxGNO0MrXIXmGfik9qUs44UFhYF+zBllHHQ
5fJ6SG7N0l/sdZ1R54P7Rj/rE67O6QIlgnJ5DWJkigxf5wo60XveaWJ0Ga5d/E4q
4ts2sB6ypcrxies2GhD1u5Eg1d6dYhde5D0VbkKtxZqZGSo7gvsa5uCZsfcH+yff
IZ+VrK7Oijzy2g8SIZYavbAKLIYpjL3Nto0J1JZqe6AU6Eec53nwaGPqal2loMst
yQ0cyHVeeiN7jfQNRKd9BLmmWKlhXeW5gvZy+mQVyBdUi5Oy3Qu1E3ESdjKwga85
hb5jFc+0FBDFYpTK9LTSIXo7D8eM/wfurLtkaT56eXejavYIQ1SvM4C42gKcMHuV
Z9LQ5BwZjhN0zk4f4+da+pI5lHCaF+HId1/BelBwa1kAVxEkt5gdYKmS1Qy6GeHS
+xBIoRK1AGERYJQGW5R2+iRg4dlQyM0SHtMdUav5eHhLN+vf5NFQMTs7P0YuWNhf
YR70+G7RrSN8kwOeKzDd35TbShI8xN9qNqfXM6qwLTATRvV80FJUy/+KsY2KRwnO
AapstMjnQqCTsi4NE8rcp/02C7+WG5YBnFcRSpxm1lbldNAsPsx8Oi4HyiD3Ep/Z
Vkv/O8CCKgBaxFxMC6n9ZSIkGQo7MEuCOErl9is3IJibeJqo18n/NkWVZFUHJBY+
tOkj9dGngs6+K1+dbuAACw1cGh350zkae0uklqOq7YJZ31IfIIes07iJxtgWiDJ1
s5EiGAmF5MvTI3U9xU6ijawkC1E2tAaYQXVOMU7hualzR+Trmy+o8H4k0V68gyol
twbXNUyt1LwdUo2BEcxp6IQJWTsHBdLnIaDiTG/xFmYzH/qQTtlGIpuu+jMWP/1Q
YXidOcEorggM3bibdUnypHtIFwYQHWBNcYiYVCZzupHMD0QEjaj5oKdWUpu16Dof
em41F0ZDyLHHYOXPnqCphj3ke+kkPYiMXy2FHFFdoAdQtlLjCiFsF1AsF9GYTlfg
ZJqzvWDffGqAzYz0VsFJnn8y6n0h6QAbQIKrONiGkTB2VlwHgIBf4RExI/So0Y7j
ha9gm4aBvxp6RBk9ubWiVzN/9lqwtc6r6fIry6lM+iLR8Elugac7wM7VbxkoTH4a
kRtgIAIzQ1XQ1U6c0u7EDKTPK9MwObIUO3I4iu93ohkWJR9vD8H1ilvv0X2DDfK5
dSQYqLiEYhYMQz8m8FP5RVLngDDoke5+Vb6NLv36aCxGRYiIj2HjjyYDqPgXQRBA
qqtmXPyg5gmXd1RiB7vyaCSr7B+HSEZmdz1L+/c5Zrwe0chs6HPS8F9LnCUkT6SM
XCtEqesf+BfnPnj5wZ8zzw522Sgi5h7JmmUkCdyteA+60PMqpXNv8yyIJAYzRHlF
hOKfZs/PKCL4QM6zPD9/t6HSH+ek5fWRIJk1E5aBEXVx+hgMls8LDhT+AlWiGze0
1hJMqGkCw6sYu/+U6iwp0QgNumuQCn2qTOgMleKLErJPhDaut1Mz3GCSVdwodHd9
RG1MP1xs+YJO2fijdMnKLTPo+EUGuOB1GxojKDw+830yHebd2ZYBgZiIolQbT6+T
zJmFKIBdD6bMl2Pdba970QJ/myJzsQ4pQQv6xK0o++L43rqwoZD+7W5Xucjd+du/
Chj0uJVKCpvzT6BIct9XIF/VgoVw3Y2hChFz2liRi9cxo8qzUv7h0Y8IyBfJ6E3K
QQqS30bEckTIfwDf/hYVgx8KsKNoXtO3yqSoFUqZlHUDEog2ifPPMKOZoqtHf7c0
K04VDj1GP+dKJ3RpKZUEqW8Hbkso+LN+kLOb3rCNaF/deQLzPRR0CCFr2zGrfwfL
qgNtmOJpaaNn/KzwbDCjU1/JqZtPZDpFWXWhedXPhYCGbKRbElliwFFfvYAwEx/c
5DLguw7TjIWjUetmO7fC0c0DH8j9MtWOBbe7ADmlvfNgWGJaL0gNTGgfTLCRFvzM
DMO658EDS1YFvLfttfCVzYWD6nw+QetbJYu+PuHH8dkz0mWH4KOBhRuBzcIVPYw0
CvUY1NuZ5Jzcv9REEkA++y8wNfy8pgxBI2SUzkWThtsygRvlv0y2IWxOgQEqqXC0
o32P5E3qT/KNc6ZwCHW/jWM1KHCZg1YZcwCrPObJK9u7ZNh3Nx2LZ+FdnKCTxSDS
kTPZsNu+GhR3tC2kHdazT1nECqHdA5A8/OKp6fn9a92H0Dz0uvZG/smhN6UvrJXc
hB2U9i+9vmi8sj0Vy0YvpE0dzeqVlSZlFW+68jYmkzW3LNpV01XwP/fgPQ3xsGqY
iJNihNdFUC5XaR8RGY8hAPAXxX3ZuPnNGMMTJ4VrctmLAIcaXVxjgQ2R+GonU/X0
ABAUP+Z8n76IP91nhG8jzgQMJhn9hujapYo91XlWw367ofnXEAJTp6O2O5kk5ZwB
y6BNZJFAlgO9Wz3W9zqkaXtjmIeCdQNw8V93zjc8D/y4GIiPZFbzztOi/10ez+Ok
53Cfp4K5K5wJvGXeB96mqHQbzpiBrVomQU3dsuPQ1Jr8g6Rpz8DSsN4nnspTcreq
3paMoa8hvo3azKEGLs9Rd2IWQP5uxbXOgcAble8sAt4B7dobrQokZLiA5kFygwoP
IHpnf36D3t5Nj4wwEkApWcG6c5IW06PG8/VNB7pU5g7LQaX1Hulfnh4ygzhv/nY2
UwdN+cloQx3UYjFVPHpOfKgIM/tT9C3vKepb9Q4vhuhFeSmNPFEtHOlYVcNOWYL8
FX6AdjrmuMflG9mZ6G1eNmUK+RhsEwFoKbXKkiZrBWyx/wBvhF2oDnHwdl+d/N66
zV+g4hCg6QBORdF4nde/T6O8oMR5j2Mkig7O24CZXL3g6PWRadsHEyatR/J6hTfo
RyRPmPrvmB2SDBDylvhBLkpP6Vj3//PmI70cyb9Hr6nXeMx4hFXNDhLc2EsIbBGB
o0Kbgqci5XzaJbioC9yIMjOQKPYp0AoJvbxU1uRd/V3KsIJ+izHooCnsQ8Semey0
jvuqKdBQTkfUpBsznVFqasHatIlVAprgdNYpOn5Hm6UMjmQhf26kD/7dqHLGhxbu
p0gDUXob5ADSh7BbBSskVTKnkBf9WUQsEmq/V1ApAjjanAg4fOQ7nRM39WI9knx2
a5s4UY/f3E3O0pj508+OhaT+G78RuzHlVmeBHPHLVGXVYFUm5QzV+wBGsRmAjpof
57MZcHBNnLSQG9g2VT2+QeBtupEGZPocEiMlZ0DUn1199dmw5ySviAXR44yU+/Fy
w2gdcpMRvZ1dQEd+c+PCzgokp6/MB9CFSuFKUwC8IC4ITYbdGvlI8v+LiUGCJKtA
210zhmLOCO3wo3PjF/XRQmNjDpWwPpWw6/xjM8QjVzHr7mY+26DAc/nrvQTJrTnJ
mVclCuX7dVb/MpoqSpNzQ4vLjGcSGaVz8CwFwqp3IGeozgmxKjaA2fQr4SBxmpiw
oy/WzLKBvfnGidoQ+G1OptReZvdSssXtc3bpjdI+hekE/vmV8IAIU0phDIN0OP2r
ShSdLADLVXK8uSMc0/xtss+wWb4rP1ph4pHexplIY+jGGukjFa9RvNmJXRSUDveP
uIVuqmbUJUs0DxN5WeD1ikhYL5f7c47B7Yj2Aqz0bOcNy9FD5KRKcMG4Rim11wPC
03LIr2KFuRYZrLs7wEt/EmyyTKmrKoyB3k7GpN9RCt1lU7p9J1AfyH5IGekovg2H
ZLn4eLndwvzoz6wn2g5XWK/5X0Iry5BUFgwUR1h+dK9tEThNWEMyrO3L7AZO1YHl
4abaFl8NqsYLJVhxbjr34JTGXMqVzXy7pdJQWSy1xSGO3LQVe24fTaFBAdwbPwLm
OE0MJRoYbtStvbOkCcU+6fSRYFgQAnDkCuZGKwGQupPdZjDHta9vp80EPPxRbWPA
GBuo23/+SJmfyp/u7JRV94AwZbSUnoCJBCTM7+NrVbTagVtw1b+vx3E+q+n+TLs9
rE4HPT4bh5iYLNP7fwldgOrfZ3go6cDabomEylOiiwyPBI6NftvV5fOozXt9/rlS
yep9sH1OU15dgfRieWi56JhZNBuUs+WjfoK0HPc8LWlgP2LQAHJHJg7CN3aFI/yn
jsK1+dDz9AKxqpW+L+JlPgS2Bp9kRu/lcUuqU+MG1Bdh7A8FH1WC13aW5hBngSNF
KU5hW4jMlRmIa4qOpvzzYm5KTQvLDg5e7yYZoCzwn9VQplgNA1fKYdRvMslt9YTX
KgL8o28EAKomF65c1cyNqwZiCyoc4EIEck9wre2mB8pFzHFJ5673KoaK2iCTesyf
q778yHuDFWsUhfvEn1u12G3vaS7m1iG/z8+927QV7mXtTmUBjPPoI3eqt+a/sFMX
gHDSpLYteEFBd+fIpQw+QEeD6Egw6q51f8o1mPs/thdDipK8VZl8HlVnItDr4jZ/
oHBjHgPxmU3DOdndVTWI1XVxryFzdTDBZKkUnowYyRGps4gSmaKFZ7baXDMvrnd+
hjMM2afaNBu6U0J7hP48SWnNudVgJws6RaPz+wjqcWADG3dwfQ9DN+tdPwZMKlg4
k6nUaXOSaP4RvBOgejSx2MupOuFCGEByTK3XsV00OwrkTCTjB2zALwgmUJm9vCxT
NqYtZsFBidUc75dDOB5mBw1azLyz6aBghQ8jwIeBfn3Wi8DRX+PlYKijQP0iR065
K2eKZpxKR9Bzo5daLoikRKHRPcYm9hI83lw/ceJGRsDzz+Qz/oDGujTfWAO7N/T5
/94anMqI+IdLanYIm50okvKYMFzymlywF3tvl3+4KFBH9ntcPn4CEjt1SsMj28tx
9TuqwK9I3qBv2o1ximJgTjVbphQTePdf1yvVAlubMv3DLn7ks0eUnvlmImaUbrqz
K5N72PQBuCvS52uWgF73roCjGNevEOFMTXKIM9Xh95ur9fQf6tjynXWMJfnfb3c5
qD38qZ6JgAbZ+p7OPRzUakZ13aGBMU1scH0FpaJvZjJwfY8DJedjdyY1a5r448zT
DB+Fqm85jgZKP0VQ6e2yuPFl59MYN4N7Mm5DRYNlf7RBB/FphIP8mTw5oWlUvpZ0
/SlQXOSufwDsumt9zz5etp8JbhM9lzchHl3lPga5PsP9eAx7Sx27KBXvQEg34OuI
opSGwezg0v1DKQRRhSckxA98t6gCtTEBh02XHbfy5uYWTivY4nAF3CaLyRXChav3
cmVy06YlivMnJEi/IP22ZP4zGsGMYsj8t2as1xi0kG/GdbR070lDGA0dPqY/FGc/
vytCak2XS1JyRK8rnJkmae67BVAA4I3FeG6uql/XV/Ac89dlR8pi31GfB9Cgo0SL
p4viDs7beAgHKlCh1ktn8LgZf6HL63sqttdpfjHHH7bMewdomwilpkxNF/k793x9
ZrixBLPOxLcS7OZrnYSux9DebKWXWNpmQtX96t2UIt3jFmUC1Wx94C+9Ny6PpZcT
yESuHoruaxw1xAWt4vvT1B7ZnWvYKdDCI+jUqXif/Ip4qdkmgKVbZVnbMKyE4l5x
3cOXYoSBALaRMDJ1E090UquRlp4NVT++vY4VhAH73QLeItbo6TnQTTqRK7rRiI8q
42xuBvj2lykMxpmAIworDKPCvVbQtJaaAch3g0h0fM90gXdsqgdciDE6b3LrY8+o
5I87Q7MPAh326ebJ1734fxKg6zpX2POq+uM/UUY5YmdOdAdLWBXOJdIUIKADbjg5
ST0ePS7UUWJflpzwIINq+JF9aoaJ/QhABxXF0lsVZqmkfYP0E3mmBXcPxkAodHzn
dtVJJS9HG9OZ2IBXH7aarJgOwtxcyVYNCOcrnl7xS8iLHfaHpdo/yG+kNOEOasPK
Si7RkFc1GpnN6NJTzk0/Q6eVsh3MfFrS0OMhSuhBg5pZZqbkfLPuRCUUTQfYi7H3
rAmn6nKmYQ1lfOtQsZ0QgEtpI6CNbuVdRD2rrBnzigQ0jUX/L4pgzJ06uXJF2Fup
GvxyB9m0bYWKoubsjgM6yb4ovoHOzfDk0BVqhyqek4OTYoZBYqbLr/bOSefM3MaG
znfSopcgJIGAZkAiokgSDNTmQg5YDsVDmIjXShXIGLhWrTLTL+aeMNVUMRqkDecx
WEMw14dU5/rIcx/8IMi8RUgrUZ1376ljFQedq/zFkeDhRGXGiXOrfHYccwCdepnC
lMWkYfKDa7GPqhPh2IaB4WDHmu/KHDXpa1RhuJpUxTPXCa0t2UnjlZYF8TUwGjxn
uukNLR4CDuyBK3/IFgpYxktdQQcQEJ44YXPPcy9M6viX1Deg3JQ1Em1JSFa/QMGq
eUyeoftoh9snce3XCDTdhBhsPgZPzWDx1afqKd+zOJhPXTE//EcCwC3q+Mg6V4se
vR8sabchFjGnbtFBef092j7nkj2fQ+qwiTYAkBEdrnD8ZatGmDNLlmZNJ+IFZtB6
yicy6NVXEjJ6uNYrCphiznHRbmyZWXOI6Jp8m5n+pHDOaEXD1jgyNmQwd4c95tM7
TnzTF6LblZpdq8i6nogAwzB0dQvdhE5MoWR381XUP0eWTFAyB2Vz/4r+Qxt9Ug3e
e6dnrhed0JKepxDFXCKe7syQaXZKzcrjbE3dSoKZ/QWpQy0Zr4B1jjnTUh77VYVN
/ZFgP1N/qHWX9FTKzvAU9uzSIaCo8sAnTgfMPuUSOOCUwBp5oSCE2IPyvVIY60jQ
aTCgGoeWJwpXdQzSiamhVU0/dIIDARYL2hcF6Zc1CErPhw6V4rSz6wDVCnbceZyM
tsRAdhFLbJtHVAlE7n6Sn1qRYD3UC/KKe8h7BFiheictJkGgvG099ltBU9QLZ4HB
4R5Zxv0d5vjGMfACXQLO3WjNIlfyjnyJ9NgiQYmVgrTyGXqt7bRanT/7IdZJZAuu
HIkSNs0ETH5bOMgPxg29v1m6AOb1ESwc6Fnttg1QYMX2hBtDnUEUqFm2Tz2zjIlZ
wPLK7fYugyub7BOJWoNVZa7ZNL90oOImm3b2NwVPCQCM/6w8h8nI4l9MWTzm8cKn
Pny0x7PdVl2tHRbygqfnzsPCzOMfl511/iVf3s6K31///nMa3e2zlJxDsvC7rfaO
b1zRBGF66ei2vLwu0nCucNaJAomsg6TBTw5lj1z/oLvU7J903mbYbAxnJLlFyZCj
8SBcG86T0rXR9FHXUPhLwB5Wr33h8cnm46Fn80KPGpgvWXkYwDfiwc8/Z1ZmxLPq
yYBmtq5e62Ju2y5hdvD0lr3NOGQNQzNR0tHlYjhJzUEQbjTNooShRBrd5kivmt3G
b0rNe0L4bXrud0p+xt3t9p4/iFSHymrxsXGxs6Bn3k00xFiHTsGtiVgYHEIcypNH
3QFjQDAETAqIFoqqTcjcdd+JhBClA/i8SrFg2EMMiO0x8OLy0UkBtOyHng0xcN4M
/ku9RtGzZA+0Nfu/X1+gbYK2ALzkMcX50oNFaxYZaKkke+2tR4JqsW6B0pXN1n5X
e92pUWCzndPQ+SlCm9upLSok60n+IwSAfEkhAAJzbB4ULn36YHDvw5x3eoe1bGO2
GWWdDj0xN16TTB/nVB3EYh8Y4AFMD9y8lAAnu/kQGtAt3E1TDxNWzOH0+kZARdfr
WRQaLvXYjApCGSFWirT2iyMrBMz4D/ENUrMyPdY54bUasJBcv3Qr1K+WEkIOc370
ptCj51NP624b7KMYcS0kp/jINsXmKL0CBx9eZxl7eg++yCCzx9PB4gIV5rTLJ+Ob
YJ8w24xAt8UxD3ggn+VpWBgEe93CEg6W+DohzvOIWk1F0naptUGopXiKv63ASpc2
0DIJya3vtSdGmt7teSrRfZSkJlYqBoXMBbU7TOlULGofXXuEfMMYWq9JkT1aDQPY
CiceA5I3lWp2vzO8vypmYIb4vfOhd3XayuI+O7c1G0sNqdDTuQe5q0g3jtRYg8bn
HccMpH07YKsTufubLNO9hUAf0ve4Dl6DauVSa/0Kd1ERJwd5VlbUU/gHcOJTT2t/
2EXihcGIv9RJf5mvD5SgWJkvixQp96Ni4FxAa8h6fYQgVskFby5F3t8oSt2Ypw3T
2YCBZdu6klMUDGxTbSHRfKPczVgyi/j0K4+gYX68bMyvtoSBwa4WVEa7IkC7d2aM
/MZ4CGqx0LXz10VQgCc2+UJj5idT8wmD6tW2KMyL4iDc2eOdJkJUQwBloeu4AKsx
0ELX/YWQFeQnFZWRtF4cBnOfy9lBoGxGa5jVxPXqJlHPOKVaS61HqwhJmVvmbqlA
KkY7twI5v2dqiEr3P7UsRtbdLxz8wSxlmSB97LxaGTRz8neW5j7uAEJ5toDSd16G
vJ9fYoYQY/IQY0oz0MZQu4hi+qHwr6uv4kFK0O2VAMWnbD5wfEI7aFfrKmAEsRpn
Q/g1PxBd0BSqTHsrBh/FZNf/8e6TH11zvh0xso5DxdqYYRz3A9N4/RlIuwZOGJdc
DfKFljau18upX/45hIOIAVd8oyevjp1fOq0ehVnJx3G2P/TSp769XF5vYFtTfpzb
lVm9hHQVEIGsSCOkMPXdgyFym1YEwOKCsy30DGmqFvgaEHQ4hybUE9Jzl1NYMq/2
LRkLkH3rDbl0hZwelOrU6so81586wYYpd3tF2l16xsdcqBqo8xs63zo7ywgnWRaJ
8ZtI5Ueq2bSVpdx7QW0DYn1c2tMTEtI/1hRwpsBpol9dlOnjUYgZxtjoDqzxFOvU
1hWtOJ8xKG3AeLhhnZzDxI2AGhksVZlClkrPN4MA/SQ/wCNisMt2SsOrUF6+S2Xj
9wXfNZ6jDbDzHrCs2KmNxE1/DLhBzLiZjfidynJbxFwlV8QE6NLVelzd+/7xzHBg
kfsukKtZqDXzVZdpBtkpeSSXVlEo7LEGUQTEntWmOyMARyY8whtHxy60EIkvJ7+o
ZSD9jiRgZ8Z+ojfNM91y1NfsmYg2o/Uf54sFMlWwXtnUKzF8hqXMIXEniEMwZZ9y
yTcNLbYE4IdjAZK0rw0fRJrWiEITwdB/NopX5x3bM9+lMuVUqHsvR/G3aI8/gZFa
6ek1NlYSOfPnaJF9xr2saZUKkMzoLGVuEYgaIxJHn8vnRcCjsCESjDYK+KQedMRS
VqiBrDkrIydkGvXG97hAy9kLHz47PL6mMcPalD0bD1IMhMYGSz874TzR43JIhZUv
tnYSdk4HN/k7wNKc8lH9ULtRRdzOcb6m1aOffdoA4eGCnKg2sevRyMOC8Qc6L0We
ne16TISMkey6fPKhNv7zkAq8URp1ricy31wn323BH2TEAlQGrIq4ZKpjkcx/zb6Y
PM+Do+73/XZEtemotCkPIGqRT4q7aAOzvZFEcKIu+VT0EOCq+CzB2xNsUMeZA2r+
0wYNmzf3klnRkziS/3h6J1ijoSVYhT1i1kF6QbKEdVAgTlCPaXo62BzwxCovRiL7
kC37chba9a23pku+NpGCNCUMkbXTSr8GwPf064JnVS3BU1Wr71r+fYYE6F9KUdcR
sN6/OLkZRzzOxzaeyY42eIJ+vR88NMllc/CCla7sXVh8YwJOSQetXKgmDsMNYqle
zFkQR48odMX9KbpOF27jaiIbuPfmkdLUobhYfbw/5jJCOIqlkKcNShmn2KYIQqr5
y4UZhQHAk7yeDzraaZPqkO0WL5KP8AfGj5RhI3+B3q9CI0cdXlxGfEF0CVKfaBRW
xJX/vb7ZGWnn254xBHbT/0ZNGhQc9KC8e16UhsdYKhYfZfgJrUUzE++jGvJbtst7
cGqNZeA1Z/U6ftLE97rkWrH1/ePmVbMWkvVsu8cT++8J+BO4tukceUmsIxUH5sQf
Pjbrnf/gT0BnE5usY71twzGynboq2ipyQRaboLUnDj+ubd9RGrOBMYRN6tyvsw8K
FOVkbmIJM7OIe4Wyuj7hp7A0AdjHdi27A4Ud8RblEnDS2AbyMgVXgA9PnKut/ROG
VbE29mu/v5EpFux6UYKCEsn0sD+TgXgewPqNVuh31/cOhQH0RhHikbeIRI7bBhX1
psalChIHjUHHlRNnvdNebvArOjoOOw6quZ89zG1CS7IcknZasWSjf2yx8olDA2Rw
gyCMiLTA8q4G2RNidYfc4xKF+NEgZsc2WijwRwedup1IgKbr1DJZyWRtLkJC+lk5
BGBY5fCUkv2obrAxACGm/XeMZoRB/8PRa6+ePcTi5fVRB8yFIkf0ChW9sswAlMvZ
Z3E3hd6/n4EufxwlPauKJPoF5I3vYaENmX4rnJJoJBrOtOUzlWSVwqw3bL6tf7No
fumjv6Rv1JwzluK8HKfQ4YB07LMjmVo6C8xZGgJkpa6qVaEZBQQFG8sNdtF55AVd
gfrQvh87aiprVaI6ruMZQ6ZUvZ+TI4NwUccdF/ZmjNrDHDR9a54Qtiw5mFfiF/oj
9v/aGPCcwABM/NF8BUz1lxKUnRwuWc5xk6p69GeRoASg2LxwrOoQwhsD7/Z2+gb7
MiPnyR4gd/uHDJaHuhNW7DkgKcVAX1HFHlheSSzCiAFLhf3s4TzAGFGignWazP3I
t20Q2mMZ1+I+V/jVXpFjvD/ZVUsmQDOjDgUcBM5f7tx4zpuu/MYlwv4TLSVcxwy0
VusLLdv1gMxK9X+r77LThf380H9fH38+65t9AN2KWd+DaRkGx24ZqCFMy2jFNVzp
1VBZ/skMpcpYfn3lICykbUQCYW0CpW0lr+j8gqo3duiYq8w2D9KMPz5Lu34kWRiG
Zug+m+vTeQpJlep7Uz7QCcbJhvUsg8TZ2UrqagEPf2e0o+JvKeBVGcFl0oPxyIPV
59ATzE/l8A/3wgqAkdHv7CXDcOK5kZeZNoR9sWia1pt7B6E4IoOzOD/cvz9Rvdbp
TYzyArAJ29hc0Kr5tM/9/7D09KPly1DN/awzHMRSCF0ayhjJIMUzI2n2eL6gRn9Y
OKHfokk4L4NYuPkc7WMctiBINqDHtEc6rU17XybhwIsYLQ3EzfJ/Cc+1Fp7CiP77
t12d63F6FUGlEu7SBPsfqJDk+EnmLqZuAsHUBqaCRMg8N3SAnXjRy/MtpovockAv
B4sk5E44d8oTwdhvh/kifYTe+Mffx6ZLR45H52G86uIqQuaiKtiIGNMNnm1wcDCF
JxYXH65TgRNAcAnTKYiJ5PAUV/DX+T3GaDaCFO1XXFUx+JV1Pwkj/dXR46IQekgl
PidIOz6grqB6z80Hwv0CUoJaeMD5QWYPUuwH0PGPyap4mswmicIkUdk8Hz+iMRSO
3zi6xf6tsg+IJ6lcYgP6G7Q3evP3/R70cm9JcYZV70LaYnY+KpKD6jv+KRuEb3Ey
2uKL4JN/3g4q1PDwvBnKEQGdr/hiXPlHAsXE1FkYgYKXWpWad1M3nQ3xAgRKH7DQ
rXBKAm+cLx07haeDC6/VmHdF34bum7DvZsb/sY8LYLWh2ooPF2JU7Ske6csB9ARO
HcwOmhWsgPNyPYxsGmFjJot+GhTwkwz4+Y5FljWWxueXHQQVxK6lYwopZUqK7563
/ulE+oGlJpCCrE8ELofNtA2qdGn6M4HJpk6FrD29HvTWUr6RHp8ecB6mkqs8JqnO
3GNNfZqID0lBIK7RVDCt22haoiHx2KwQydOs3ONl8RKYfhSAPKrcj17nEOpYpN75
OkLfiUP3+rcMZZTs8sj0loOmcP/LSEHXiPoL8tefq4Y/+ICRvR/stH9xW91s/teB
mPOGx11ojF9X9Hy8zscCYuUU0mKw8Atve+fE1afRNDtjluqR4h2fDaMkv88DQ9Ra
VhmYpg+Oyti2euBBrE65prt1o/XNn46jwunpQy7+Wjfa4YSZyg55P/7K73bP7oXS
6GoGVpV7e9d7NoCUn4oNzPgW6rCjDlwfG/XLRY2Fn49WmLU/9pph1BAfXEdEqTcm
T4qni58Rb4tRhfri+IMKLEHXHzQuiicI9msj6XyFC312LSET25meVVoA/DMXOVvT
QF/1P4a6WLBQ+clC/uIty0iHKrkcNTwRSDd66QNxy4asiSwb64nVsxdEFMuW5jGc
YLLGzItkeGc1QQVSQIpBf6NdiaLCeCUVzqdabuYJmkjPSP+KGwGCDSbRUzOiVXaD
e9sxijd1DWDP5kFaEhRMy236j82mal1q7T8GKnNIP3+JwfIPjz7EL5bLVb5r7Sg1
56ehxxEWfwt/Q0or1CpxRax4G7kVDQWeiYEPFEkZBjAQJ141vzrG3AsqA5Bi92t0
2dCvC6ksWiFbFUHY7I0PV3IR0t21AP9JXtfpwpd4XyLJn5QjLbwO3Au3qQVL2P59
yBr9z8xBEP9UwBWjiT95u+mzG4LajP9YY9nR/jOhnyllsJUl8+h/nvrQ90j8FWX7
8Za/blNE3Uz/cqsh9SLZAWwExsyH59v0HcInfc/VmBOVhiBY+GnGkJ4RMvtOYEgf
DlKHvfk61DtplCveNe7hNARJE0DyDxO9OzROn5ykt+8mOhRbNsZtrrmURiKpWcMA
oHWTl3dxCstwyAfmCBse+3eZ1SJHv9WIeCH2PsaVN2HPRQMAbWfnHWTnm1orhBVf
GJ9TtNP9XDKuWpeI4OBdUvVw1qNzteOTIz2pHiON/Nd+Nmv43uznspnGfa8pjCs4
W7EDT8sXF4oP6UJRS5MDixhigm9LGnZqbHX5y5U4GoZfzLzroXiOUJVU4Nyu/Lez
FBxOsdZLqCSKozZ1RX8K2Gjgl6993HOHB8WEpTrnT/o/c6jBqBTdo60uNUJyVVgp
Vx7uyGe/9wRlBhLPDpaZuM9jsFo8y/G5pg17URlAKgmLRCNaWiOTobJZO2zgiBnS
6nqgFrpL5t/K1uJY9fMPEkfoGeOx39LVEY3wIvg6g/wjSWM9mLmqWtvPHp2mr36Z
VkFOT2LSXbYbwzYhHJFcgaxfuqzVJQrMaJQ45G9eIGDhFwwPe3hC4TG4ty85EZs0
BPRwopqd/neLnJ2MIPC8ODkS7zh4p5sn+Z/TUwT0eAGy0wNKMCbPEfgU7D0oMt2Y
74jTu0lWqQEMmvkk5VRphNeVd8JyzS4ltba/+21XJ34oj3FmypL3Zbg+nFCXJKgi
sb2Uaa8Sh23Z2UfiOReo95SSwuuuhEKT6Oq4pZhnHGXmmzMIah5S6isaAJFImXLP
kxaPa12e/N+SrFmjDsjxuoDLpJYS/H0FUKIQi4iYTZ4jAc9orcVil72Qv3EyzvZC
3WyvByT3ZgAeFaDG/XwWW+Glel2uhzDxMj9KXNnw/FJhX9eItfXV0fQHianuWJ1Q
lZ5BPNJOJEpwxFXU0KUKcpnivOTybVT1iOpEn2768H/m1G+qZYzKTShcEDT0X4sj
jZVMOEwQiFWtyyKbIYigHIW8HeWx6HF+sg0SRBAHmtBnavIjAwG8mMm2bXZOkJ0e
m+LW32DPz3LnrRtVm6+NOUFbldjzcNX55GgV8HA/U8tiXu5Y/esWjkaZk6kda4sV
97tnTxjxLCkRJHtNk2t7cxwEyQWDfaPZmwu0k/Hd14U3Fr53HX721mc1xi/v95yB
85TBEAnCUYQN9tJJhS16p4cfxvZpc46jvFaxpDHhgk7IQHq7U2gytFsnVRRhUl3z
N9OJediJgvQRdcemQg2TnmeVE9pflayyhiL/PQstmsGyBCy8l7WPhTaKj1EwJE3Z
eKsjNRYuUgYWk+j94aBSgIzXhGncfJ21h0cIaaaBmOj6GLWZcpH7JM8J/3oc+AO8
2Lehg0mWZs9fooRdFoS4nLa1EU87u741XKpbMzmCRWIzuYUqtSizqKzinSvCW8TB
2DwgcAXedBSl1hoV8tONqjptz/vCcvxpMta4Lr76nGAiFGyBeD5hQwNj0zvwFdpd
C84wAmzCSk9xdIUBffPhXtAerUKfRZ7as6hXBHOa/t8Yz+4UFSfRaE0FuHKJvBIV
cJkb2+uy0HUO+keYME9V/KSWsWuhW4+D3WANfhYRjtz2F8ZIvoFQ78kzqJJjEcia
8JDV2RskvX+TbcBoU56afUFIGNeT8t1bV0Lo1iJxZRzo8r5Cky2CmyzSfKRR/03d
ES3aHvPEYBij6g6XMXZKOvzj0ijC9olBXBuvylH1HvtQeu4JgbptK6AtsT1DzZYI
a+BIjXTxwtaa5M0I+mtj54iAPJ7HzlrCOwJWgKRONveAEOA1YjBoGKpOrLFmcmOM
XusjYzQKnaYdLEKXI4DrnHyOBh/py/gORI/afBcNnisSPlvFJx2bw6cEc0vOe0u9
LqvJR55h6H8YdlgNVeh32T/EexonoSm4LSEpjRAHyLfT6IUJFAA8uYgIkaTCzVSN
tmOmJ670vNxgKztjQqRrdE+3ZfqExe2A96/1tvWHKkTYDlHkdR2SpJXLSRwL0VtZ
dVEAvRTDgnKNdJR1MdfaLjIqiSbT5AE6Hzrr4r8oUvWQLp2+ResoIrKNw9yFfR4H
DYgAHUKtkqKBSVEn+U7E9ktnAp2lcgZcPD4vg9KLa6s8tuctxMVt9FD371zxOkXk
8HPKWMT9FYfNvFfKR4ZaB4P9jnJQnpnfwyBoeQpcYaT0bj21Pw3qhRvKiU1B9mli
6gwHmWRlJdr+5zf/PRnrzZtC1zrJv2At8oa9mDT6aLJkd2+Nn5VRJUtBksPuBhCG
hKakrlxzkABcQ2UPQkGkaspK0uSiFfUPBOJjzO++EGWtW2jn3K3n3nBsu1FKQLV6
matjAIYnql9TlGkkef42k1rkt6gRJ152otYbKeWnZCWS+gsb+kB3or1g90QuwS/i
+0okPXdE2tMvA46Xc3MRUx0bRKX/+WPq37lhrDJgOujXlr12ot+t06CSoYgRZpWY
RLeN/zPuwR/tUD4y3eQUKFhT88pwikKTRC+gE1qL8eJ3jetm1USrlJRLGUbUXWKd
qFHYMWQ6tu2a8RQYAl9Ij+zP8wp9I48yq8SwsZnG2tTeK0nryRmTgagF27flLrhC
O3CPLbRBwX2JnXObmcMVCHxpgy+CwpQ4h3v/21RdL8sN2gA7aUFFhvVz1qh+pX1F
tftmTNBZQYv9Jvw/sbHW7lEyYDbwx4+f4yYsNGvoBHWxI7z4OFyqlir1D+823XE+
OONdcvl2TztnRZpC/8hZWKHcWqXGGWe7SOypmCiQZYtDkPnT0qGDfQI/tMungUBt
E/lZPHNvuI8+bLM0aEVAuVbB3s1aHuZA51vFD0cudX9NMcEYoFM8MM57dZPKhofR
g8oYAdYTTbGbbqrsMWBbA4OtROEHIaJ6h4QdWgniU0IHhx1FfMCvp9eS/1s9ZTRF
5NumgEsGWTsmI36XvW3oGsIWLHp8722gJNTTwL3Fi24/TfbvzEksphbuIOGZRp4t
eFWrKC1W2sLVslXlTTxueecdwdI7T1h1rvweNu4+r/0uXg9kZ5tXhPNGjiHdAUtk
dCkwU+zA6/25JrpT9ujgHvwYZmAAt9URR9ZPZ+8BGrkiNba+qRVhoPkDyFtPrw4S
GEs2Kvjny8ClNoHOZfgluQWcfBc1XIPyJZCSfZD9tMNM0g9p6MOySTFvEiy7Xqt6
PS4IXvw9ujCgcRrdbC2RR+/52ajP0SCph8WnPt9UpKlWTehfC/kiAgkXg5iBqg5p
cQ3VPTkOhYoF3cmVWIdasZmdpb9BPHmFDZjUfPUhBn+Ru93e0V5Qr7yt7Kv0HHHb
kgLnriEIK/+nNbTXU0sh8Wiey8MrhgcoRAS7Z5Ay527stC9eEnRG/zfWSisiloUi
HYF1gwJjhfhixNa3XKMPMRBilV/kuOoucvb2uLCtvy4a6CBV8bpeNWdFxQNvpWrL
tGZojHZyaSOWiB7xG4EuEzOK92rvaJr2WfveA10efMT/6686p57m5rX55RM+D69o
C6T4uEPBnQ2EBqeYMFxnc7G1Ag/YBkbTOZHzvtHIPx3Zmvb+urM4lUhkga/ArcBc
Xd6rbvFwVL9pryVWAf3N2sPMGVzpw9K6EdOIXDhJwYuCsQfqGCfR3tqnKORw65ab
3g7WXMVPIs4/qVSH35FQnEHsXa5TKeYH2mbhLh6eEUaRn+lmYh9dt42wKEI/mG6i
ihOL76Fp8bScT17SQUZe3wyKNhsTo3iP+MMzqil0zLLnxfAyYS+jPoosgL+ex2kj
feRYy+yVUqDqt8UfizdG7Qlz54/nl1a3d2u86K5vwa8RYu8Bfv2WT9qTGloUx0Xl
TiEsTpkTe54x5kYP4fiazYt/UAJScCsSUbriPu53Vj053KVn1ASW6p9eotBjGRgD
wLKlyhNGG9dua6fKWyYGqMDutH8VN6VXlJ0ps7td5RK4o9qTJ8mE9VJAe66L8ONE
EvzWtBiZ7YI/GH0lw8+E25e5P++GeQWZ73MYfB5ZOXHXVa9+dSXoMXRvNcWFSTke
GmXypSxkkFKHs4snTgPz+PSKhJuGT3fRKALpmfe4CIfjTb/nB/CcP3lhbKsIttM5
Sgl3WKddhPSgLE5e3DHXq3xoD7bFaqEug6z55BsHzqR2/0SadKMgN/Rb8fw+sZ/d
FmmXVfRMtSVENznDgEFx/ogKSSq3lN6ibzmh4w+HLmJxHeOb5VACuwLinQjtY0a4
vnWuwmfabvemkNf/WB5Dh8oyKUaGoReYOhsl0wKzJ4/AfdwMbY997N/sF+xCxBNZ
8pVhhmmEGlPNpe2ppFLdFbWlBrKr1PelVtnplr4WbX0IcP6kHd4kibjyGKEIYLEK
WUyXtDIlr1JVsR+5X8MJ6XivkEHLxASW6bQqZb7yNxUAUL//iAIpsjYLBm3T7hi/
KK/gXUo7VTC7krwpuNlhfD443z8iVl1V+rqmZLvuhJ5fs0oo1b6NtvzH78hZZiVa
IX7V8aJUoyMOGRyt4lWHHwaC1K5bwNuBEz02XQ9u7gmv+R53JFKlziLvjUzv+wd1
AIb5rdFy+bMB9xIELsBsW7GU32xKKoFDo9BvfAzSN8xMtA+Mk49T+gEMhfgX5bjP
orOJs1PQ1czbV6RAAnuKQ8DqGRNomT/Z7smi4Bc9Crx2Ipm+QjqB1gb0FB+mLEcF
K7FSs0rLnkbawapobZh8TzZLvWrrCd5RY5RKqtbmNQyIZaZuqsPgXp9g4JegW+/H
kM71clRaQg7p5lDauoFiK94nqvV8FvRg2+4EgD6JJ7gV1wF7CFQBo6MOfOmUo2qg
ZYVzyk4c8V2NWmfy/snUs9BR5XORbyFg35dIriVwszuWjAq+A1oQxeLdZ7uXhZLL
0KPXp1a+h7HNiGwYvI0Y1UnWJiENdGRHwzNKqxu2ON+z4kzBU7or75CZeyD4YhS3
R3gHt7ixcemYY2BopDS7JjGV/3ETOz50y8hJ87qlZ20QrgIAJ/J3dp2elWDW5+as
6Z5rChx7z2fBJd7PX8vRcPxXbDic1q5e2Y055b/lHYjFnMJL6jB5Noct24NM+cNA
AY/a+i+Y38rnm7PpcIXyjoAy1VSK9Le9xSB3HL1EAOCXRXK8ycu89eJsvaSSNael
x91Wts2kOkP3eJMMbmlvWMFgXfecGP1eHCZxpdT0xNCUxNIKZTVDFrjWStPAOz6G
j4kQ3tQe03PiJqONvbD1IDQgIDr2v3oUwuVYbpXJM/c+Lxtw/FHt2F5ZWqtUIQZh
QoTktflGc9PbsKMxOwe7CrVp1kbBb4DtfoZqvc655woWFv5chz4b1YB8GMaMBQOQ
8dR0k4g1PJtkcS0wjICd/59wyRsdfpA0h/h+t65KO05t9WqWJ6azMzDcVIzRRlVU
HZNbDZCP6OHcGbpNYO6p4XdqZSH0FO0QF3zlez2mcKRhgf37MFSya3U18O7BcLXj
s/RFIS5dfzog9BG/meIm+t3QK+8h0VtnwACQ6annQM09/bGKVK5adQuguHYtPm+8
+UeSxGkdjHD9uosYL1KZy7Tg6rYOsr33QVuIJv2UNFd4MCYDY2KQjSWIkn2az3Vs
5GZQxvAARFnzU6h80pPzQuCMcoroQV2Zw+8H1GjS9AC0Sof4iUJJGfUadvOfutHS
ddaz+QGXR+6f4TZuiR6l5oOYGeZbKWCeyDql2RTt0iOjSR1QdjAYOG+pi31BmMIN
+LrYDY3NRV72It3bIZU39U5140xDJ34gzIzlFi9kpaFDVtnhND0eZ9em203ZjXxU
JkBhbMCng+fw7vTHnFFsTaXwDmN5fB1cgCQL3p4HmCR7Z5s96sIELBVIaDP/RNkD
Jy6+l5Fry/+0A1nACE12DmdqxVMv2H/vSQunxnMGOywhC4P8n82UunOuCOqNXhBR
cwiCuvmtDhWTmUdfQZg+ZGXMq6kFWd9n1e3VPtt8PIwQX48NDZbypMFCLm/HEkn+
zcKU/5Y5oI6L8G6QX37u1hG28VfGa2TB1s78iVonGaahXrMTBR+htn25c2PkA8eP
m6syb6UK4ZRMVqGYB8bgf2H5UXDEp3XYgY2B8XukxWxVTgLeEu05leAXPXuDqW5E
U8NnywleLnnuwK+TV9dZ7MqhDVxN6vDhyDar1zeYRVXCXahww7m1Nwf0Hys+jXTP
nOEYTJSvSquPD51co7vNyIIR148sJH0kCMScowgUyXo2l5Iz+dv0dmEkEi3VAXZq
EEPO5oWGGIp53FMXuKaXVDKOpYTzonSsyILyULbTzeFpbJ9P/GDPWmz5f1hkSfd4
/l+ftMPMSDSemCvPBY18oGycDeJmKe5xOGsmEs9FN3Z3qtdfqYNS5lBPNtobU5XK
RLjlOFAoPnEJljDTFRAih4IX2b2yJ+O0jJ4cbPxgp6BZPnI29IKdvcQTLrZAa6Ig
fNMxKXsLzQjV1cDwD+FfouglzWra9ATveyOyGaYMeHp+JvrL95w8d+Q0ZuSK0Pjs
htIMVHy/p/Ly3SsBrLvXdGrJs591CFtW243OHy6KPMUDY+oyplqMp6iv5XW6N7HT
orRhmbVDKdUl8haM0R6GIyGcUMCI0Wy6HA2uW6nBOPx6AVEMBsL79fyAUS44yCET
/ChJnO7GPFsRRcgtQE2LqiOLWYGOVvjKHV9xzCed22+BTjqu2lg32OqkMNUmmCbc
HmpMSr2rAExjGBHeT7/WLv0Bw2IsjNMxBHgxG+++laL5yxVEqqYEBLdzs2HsDVyg
X/DcE+L4iZV23KMyxoIxjAYT+oLBsSqI/qW0+/RHH6EaU/zmYOCVVgCbpsiDlyf5
UWOhw2ujz+098kCKR7H5CCMRSuIxup/TnokCTBJUuv9ENQCNaJtH4LN2FxpQ2imY
/MQ6xPmg8K5TsDoegYx/P9C4vbU3ONa04upr3WHQzzHpwe5Zvkm8S4usuJ0tcQXw
xwO3ecspd2N0Vmg6an1sghZwq3W28+q+RwTRujjSsSEzGoCAp6HH7suUwzGGdYju
Qpr55iLDeehKUNwKRRIIYzo3JxET008kaAYVBy76GHVkwWaAWTsE7MP1K7a94Q5W
rIv+MSm4Iu2HDSXCn/krF2ALj2UYwZA65Inztzw0Sl9aRECZe5s1XjM7rTXKYT9g
ylctLjHv5YfO6YIWbdigpgxL9dLg7/kP4jwOZe7MzSkb6e42bJDvvyt7xlFynmV5
vrti6ikNJ/EvHyBOTdJgtsWCnjB72OP3yM1httGztZ5OohTMqvDbImCjhA6WGpZO
qvM0LfDIilSApDxFJtn5gInT1uXXQ5TbUXYPN7/uxVidB50F9jyjrTydXkpTGIQ4
DH5tt5Z9i+FOEhkfprZZYzu6K4SMwLzE5tpVmKtzI3UMLkA+fA9xc7zI//HAT9qq
Gm2tzYCVEA5B5q+T4CIFRHpf0WVjKJfuMfSmktn1ydP2ZU8YLjqzVlPo/uZK/6Ax
29P3RNUyg5/NzQZVkjJGbGzz8Hsf/VwZGazPph1ffDs0xUYymblkpjMuvTZqQB1P
BLKAzVu/CgwYizcOtf1diDFPPR7zaBRTKqe2XaI3kdTDly74hFUz2237ZFAxJwOo
lZsxICEXY3reeN2ogAEw9dv7HNEuSKxAz37KZlxefeMeoeQEcUKQpgXfgv1mb5Z+
sc9efzDmcwBFpUiGUYPSNUL92fiSk9sILFEzg6TaKVnrTyP3PsaUQpxk+u/EoaJI
1/trRyuMUIPe4WyG1+VupU1fsy/kvt+YRrAUO4fhwVyeqcgkJrZr2+N2G0UYcwgw
TQVlj3aOujX93vQI9D1hcan4AGxdrf4tXIBzOJCfFwXzFdXgRAGc8HVouYRsPXR6
75bvp054gkN5wtkwpU2fqhFqU+5fscJlD3H3+Mjn+vxmmcTTeVn+hCRoSJ0KVXUs
7aFh1XWsaFZPz5uwHeVIYv3Ki6bdMuvQr+qOyAM7RcPjnkAbQOTj8q0TBYkSnlxB
n7WKKhO0+N5aM0pvVQ/tC0thQ7LaNDKQDUvy/i46CFq9YoHIs+9YSBy5qaME18YX
0XqDE9QHTl0qaedujmohnufzVXuuYWH/PgCX1Ez6CsxVR6G4CjQkubeaucrHfO9E
whHRssGP6h4SNDEtB2ov1f1af7GKa1wFcrHmoDWBFvpnWKATjMz/umeDT1C8MdqA
E0wJLtGRf3DZYlvP4XbmUdhEdkPKqfxvttvpPZjb7blXDkkFrd7rWtXmfCcwkG1c
9g4rH9ZwQY8/PIlbhjJTboETkqaR0bryXMxBSu81DEdC7q4lDtioKxDnIH/LlNHK
JNp2mTj7ZaPVljRm2ynAARFU+6adTpyKhRqZJwiAvYneE9afdQf3SWbv2PyKfnbZ
TMZ4ED/MhWeSbaE7DTYMoNNcmta8MLAn/qwHcfWwSfAkzMvcIU9pLfU2nVMBCBtE
4RLlbuPPvz7oR4J3iZSXVHMvEhaqWtfjU8oBPuf9X6eBAP1vBsGlZ6TQA7mS+Y5p
cCcig1eBxmxYgAs2hYa/M1BM964XJRdVsHf9h1PEqgxlwZPBejTnQE/8wO8GiwuO
OgEChWG4vP/L5EYG7oSPzj/jPVWVkM2ApjVkkUeMejk4slMNJ9hN3FEidx9Esk9N
DMrwLG2P8BlNMAwG7/Ygygq3ylauFdQVoOp/9aMAvQPBPLHdcX5OrPxUtv0e/yeR
j06JB3ed6GB61jxWInZ0QHueg1c/Joib4dJAhnD9cYLPRIuGKIDkgm7JynAfQE3u
xNlVXWtzkcWjAN6fcGzzXbfbLk5PKKEmVSqK//jxwGisU3ODZCVZmBNcXEB8ERBA
vnFt54/OsGiBStl+q3EnjOe7INDQ4b9vcZwuBD+KuAG8+HD614+b/fEusTpf91zn
knljQBpt8fZiKIRVCIDi6kDI271btioIhd00XmdVMMuK86W65jAPiVQLSdQUnkj8
q+5/+L09QntcpiuEKGfb+z/LOcHCT8yZrn4BBe/TuSklWKYRJQfVFMsZ3BxG8+ST
Qj2eCDego8Pj1Ci0Aq3GbTj2WHWNROjp+PRWSNKiSQrs0NWnM9eEjtUFO7WlkINq
S+KnJeGvyogpubHFPj+0xFCbVRmvJb1Q/YbCTrLgHL9fh/YOAu/qBntvZeS49klg
qJ1NRQ0zByl5URDwJ9ByB5zHNA9+xEXIXd5aDaNDkvh2GvvSCqfh6gvsMMPkKy/Z
NSzbjvl9sjRmhrov9uYS6m5DlNzPKl0oxAEQnP9xHtTWmTuhKZcKnTJ6SlPdMiDN
XFKFpserv7CewfkjpIHxzV7pjLAVC/SX2mokjAg2932IgPmKlX8TNHoiGVVfyOSX
ZuHhTpLyPTtwi6AI6D6tMpI6XpeYmFA68KuA9xhTVvbm2OTk8/2OrK1Vo0NSI6Cx
EY0o6DJ8jb+l1wqnINJhBnSUY9rCQHXCzjjyvDMNRNVbfX2hO0qkyEd1D2tvWWUE
Svf3zsZxJ2xCsJB+LJhMIxfZENETqMBKKzCmD0grT2tcqCjBzQURtvuhsj6gqm4P
iB7Ap9cBWTVOPY4mlVHFhcEQZzuRrElcVxZ6UHVxym824wIB2yRK0Epr7Gll+fl+
h+zhwXbp0YQ2yuJH2aaV5pHpA/6CM6GpTbIEqDZvDhEy4B5HY/RNgYye/IapxjDN
6pKtDZmYAeTnQl++fI3SdfoSO6uLGZp9EnAGBr8MC3o/pg0M5zmkaNtD400bJmUj
0KkRfiGsseHp1NkaUOQ50TNYrCMqHBjl0iokVe6gT3z3K5m2B9ieYHGoXRLDCTnc
Ab/5et+AAVQ/X1w2gAUihljSaTXoRSMtQ/RHgeZ6jGCTkavU80kJ35JELiTC93p1
qBNW2v0SK6HvMMCYHTCKXrxn0tG0x9/LneovfGOKBaqPQMOMRc9tZy7D+fSpMCqJ
+sScAIzl6Xv5tgAc0xWh5cO1YkIqQIFhlFIQF11zkSffkKioiFx3/fXiO2wJmkZ8
j2scpIBTErA4/ptmXQK/Dlz/wGqW3IRmwlNBjM++EFfcAv4XjZyr1e+lYYEXNmCQ
3m57t385Uc87q603t7QCbklRhSsiIzUnw5pQVuMyd1JAiOQHgDlocnlSBigScPxZ
ZPbiarXTOEAuzR2iLOnFAM80fDavqh1/XML3AegjMz2FQc7uUc/uMUyEmrFkDBZZ
s1TaTHBkIiGonPttrBC5sUfwrA7o1gvyeXGBqRq7XF/yaMJXQ9aHmcS9Ezhq8KJb
mR92vtxIzlzX+y52XjJxMUVoO+AqxEEFYL+SaNK224KotcEU8FT0j6y49RrYIAh+
BwGs30rJblbt5n2XyC1SXO/o//oreifE/hLxOKuotz1osr92Dle0BuPsZBbgGFyc
/Vx5+g0bWhDSHUluQH2skfEa713NmRffZXNLlb2s7bAt+kly0Ef6ZdvVwDuwUsHM
pLxeQjl5wlvGrJcPkHosNLWSfQERtE0hfzfbLp2Thg1Ss02a2UR+Ex2o8mN39vE2
Vwa7+4RcaDsHjMwdtt2qmvyBJFVXKANc9EePZ9VLZ6oSHNLFYgNkGEcHhp9LDaMf
DKtMkBEhBn4C0mJOXoQL1iiiV71LKQ9lNoM2U5ftnBt5qHP1bsqvsk8ShJRATdDa
gMm6SPS/RUPI7aIiZfs0sr+d/J0nmjMIJBLRQrwnHOGWyyp6eNxdcRA6dSRsb8Mj
tnU6z9EcxSRS3TDiWjfzwFZoiPUnjZWKxHhIi9b/y23nqYR7zgGp0hZ2M/6k1Xkb
5goEfs3DtnzL7ZKlm+ezhrQANBRlH8nNWaWD9b5OuEl823ITQChu/bV3/5rjUX2K
MY/cspmjviYvzqQq0ZiLuxZ0pYS03CG/DQbihSgLwtikBmm9Ek1vfBfw9pHYvW2l
YIMqkaAZUUAV3MSz3PNrDu426cE32YVgTG6LQSUvGUdQJbj715Sk3/mJbm+k5ajM
U9dedpvHW9a5SAeynAZZ3kBJNn0z/2+7SQJdlzhoRqjh+GO/2tW4HUWbBz3XJRaL
WM9VR8TWLuW204p3U0yATrsZySY3pjVAf0Nz5wSHEfWjVKNZGEW99zEd3euliPAQ
7g0Qjo5PzUH8iXMz3uFLRmrWgImOxcVdPrGNjNhmYB2cb10XPCEMaoBRTH1dCMAj
SLvaXu+jLjkqeLwIgu/zGTGTfTGopCfsI9V/ceXSa6kNXjlNeFVJROk7L12Snryi
Tgj6Zvakmuj9Lan1Z8eBWuHuWLqRaqkjxJkt6MsR/XPY2++8/SkPKHZojTQEfgVt
sLTAORqW95GwEH6YYsQq3dzvB4/Na2W/Psd0jHACxnywISzqjce5o6sKWlDLeBWu
ZGdeTT9nuUxsn4zI0WKCPZ6rJDkde7bclKuTNeVt4qJpfunsUn9BhCLqe/1UBJqE
A0W3lGEszeLUUIMH4Ccw3MPB0zceaVFWeHy1+dsS/OnshpfSru4+MmFU3Zzifk4K
DFDyNcBMhln3hwHQc0kG3PhSNR7uuREVgYKbgVlEqYbo8FE0bzkEugQ/bHQfUw7W
8C4i14AZ2s2t0JrlsDd14UWvasoNW4prkvkDehHNOqlOMnTAbbfXpaOvIFKPhK1L
26awULqhRt0uVgUdiukScE2pbs6aEvV5a7igVhByXC7hfcSvSwKoFuRVxFFbMu/e
aY61GMtQqZMTmbA1C1MIo3CdRYD8xdosY1TvFOpicE/Llh6yrhPKHRBNBh0sXKx4
UkTuB6vpZxlypIp8sj1XBTHfvXeh8C6ADIWc3N7+B1CneJUvRwe/fNakF6GAN3pN
tT21Se2a93fZKWpxPaRJ4Vo/In3n/cl0ppP4b9eu9eGU5mKuH51XHFiTSDLls5qw
SAvg5BJH65OUNMzB0qdlA6RVEIqjo4XFBCNge8HflXtAwx53dICD+isCQQVK4Wvs
DL0Ai+0SaFy0FoCV1n/UxeW3OJx+T00Eqh2PigtcUdPAdx/i3XzS/AjfdCMJsP+1
il8lB2uXwZ8gIuWu1Px4sg4rBbsEFPzM4gv7OWue9sb3gmkEhI3Vl19mVdc7cnm1
u/jSOSFc6UBKdi4PFx0yVjXWZhKYVwlxbFl13t5BILq41578J8RBxmkDJkK8s1NT
rgJ7nBu6sdhIcm3+8ou2itfU930yQ0kQalZb86uWUsx+6avGobayA0zMqKXeMNk+
VYQjThnRZB+5tw5RMGSZXFJQmUo0r3whTfDw8/0xn9OT3sixT1b+AESyvGQ1P5O9
YzS0bq/4Z+daRKo5+2GFr9m8C1pWaP/r+d7GFkgi3P6N174NIn+YzJyCY5QB1IQ6
Rae5GEj4mHGmslGqOdfk8NTkdSA4Pf/6hBgHGSdonHcDvrc9AR2aU/zLhpxmPZIN
2wn9C9AVi7b8R45R/3Hkui5bOymGHq1tcrCYVjkytmC8Xpbkr+BaYrg1kn8w7+FR
zrYK6ZhVbBh/K2bxuw5YF914CvDjTSdf7Tc7FYknbGOSHhow9vp9gFS1dctFXNDk
OoVa9aGVA+JNyYUk6/v0b9u8xXQOCOwNSdIn9lLaJk2bAlzW2C8SYDy5A5uxK1Ds
Y9AdT9AWqquEqYpkxF2r3+CPT+AerZYXW2qVjBuelYQKTubZtNhKmdTmpNBwsB0G
nJKkHvpcpvdAN/Sh3tZ50jt72e5uuf3perUfToV8Ug0OqXO5zzInSSNpTuygY88a
O0iHmOsG+5A2Q4YC2JenT8df0EDwtZ+FBk8JHjMebScl5k8wm4cGsZD1WyzDxpK3
nHCVsDPOnV9dkOW2k+rgbBDSP9tSHA8mY+dL2WOn9nEtpd68sErjf9qvf+HONM5+
OQwUAWCz04LGzEllrruf6+toZMveanKSfDQb+jRvdoiF+sMnKAFNFlNYk5ePiLvw
bfZ+eNK3HlRouMKNq1uX522VnCKjfFFUqY6pGsNOmORJd8mlYmz9oGASJdwHZFEk
IfXrey2N/8cSydV7w18R5o0ePLNM7MT9o/TAo6+b52VR7Qyr2xXyfgZIU1sW+HWd
2W4vCZgvrZg2vqnXFIDnGtpvORZAN6yk3e33FFqmjLpWHq9fflUpuy64K1LafqIE
AOQJoMTuUJ6hQsZIZGrAGR1OQGjqisTZeTPXHne5aLmnvO6afr7ACfEHwUclCPVW
DAw6opaUqmScdduH94jhtcjaBpe+S9JHdy1qQ7hSQZKK9duptXRWdd5Esb9BgJkL
WHoF8MCpmA4tJpEgZH3rOMYEXbiuwoDt1OXG/P0cfW2eRhkRb8Zb8s5nFfX4PlIe
uONahVQ1AxHraSrUnUvGQI7mWLSjZVaB/T7ZdhtmDgJp85ZdbS61VedGnyET3CaS
bQTVEjua6CcLQUNBbAbwjQl+9Jpowci7N8MQ+zGKSrFkT37GR9+8lHdJxg1XzAhd
VfEMxx23EkQxLKj2QobjOCWDhRGmPCrmval6kRBLVl363cNmwI0VZgiOWJHNDy1u
gtAk3BQ5B1LTczoElo5PTcsfYqR1QUkfiWhrnQoGze7KR74F5dB+bkmp4tnceoK7
x1Ty03oKqm9csjVzmR5VvFM+/qZHfQlQLWwf+FZFlS/ltGbDp9jX86WZ0Ae4TD9W
4K45zcXNLzATWv7m7F3buKjvSe/YlL9xY2apNKO6lTGtBMzlAalJbSUmYsrJUkUD
p1a/RdrCWT3SrFBIvBrS0Kci6RO3bkcijex3EHrf8kIKhpRC28LCQreunLtLaKh2
whpQSSPwNPvZ1NT+aW3J5hBmUHqPn+x+atVVzBeuFmL7GrWXQ07cxW6nk0nEHQRQ
2KvweEAITY/XiHKiTd+gUP7DrXhNwfY526K3EUxlh1UP/QZo/6bUBpGDpawWNRJb
TFdQU5+AZON0RRIf6b6o45exDey7lsoQdNC5mAh86eVF0Cxzhk5yUdpYJEoq9n5T
mdt8TJh8t5B7kPzorFja2vYq5OFOrKJoMeW7/2QoYF8yNvNcHDVY36x7XmDdnhYk
M0DbJIxKGkK5FJHF8t7XCqq2gkdZzKrn7OR70JRFVDYbPnRQeFfjn3Hjlz+IKVDm
O9ckU/cJSeQylFmObKLPk6byQG8x7Uh3BU4Ji9j6bVtW+KZ2EzK1ReKa5utf4TjF
XAu4gQ7G2VmyRI92K25LbVDn4H/xMw/k0YUWT0DqjgqNMSH1RCGVUszMTclU7O06
u7LNA9VEcGE0zReD2XOMRmtnFzQ4/9qpyRc0ZPblIBUX/xCmQdlMrTC++A9AlTWe
641u8igUKWlzJt9gsKcjufLTRpwlPKjDL5l0r/lvW7ZY9sg1XoQAhGLsJcdGmeYC
BuBPkcvK5KWcq6Q9VvBxocKKDCjF2ZeD791lFbh4GuIzjWadfLkuhe1XCZpd3sdc
fkv5xwhVNVfiBEvjStstXDF0WtaGvc7pPltFawnxni3sLEt78K2sAyjQWFPt0uUf
h4a+x8DeGJRaJFL1XYoQbd9Apkf3EwFXwapSwJT+YuKx+OoCCT9DziocYIuOD+xd
T77I0fWjQta7BGo3Gk57KiYO33EoPm2uuJOcqMYS8NNxSndGkev0BHQslAMDCbkR
o/M3kkJzeMxJEflhOLadxl1SosIb/gfz3Q+MAzf/bHVJ/TObfSvANDVrjaz4R6c5
FI00WQfIbm8qLmIrq7MM5OBXzVmCmaM2whrswuL75gmF18rY+PfBRq8gA2g++07U
bFwqWVtB/HV2kA1yZjJtERqMh5gAHoh+te3BEbeG4oVKLBWNRZNTTEdFDTop52Ev
JjpkpAwxEdtNWhIo9CWKMD+gUP1pjrZXTUHBsy0TLCJbQBZ0jteK29HGUmBgTWNL
WUoJRl7y7iAsATCLjWwpHY3pUqtjYi8UbtOnOmUChV++GitQehM6kBKLeRWceMVR
8xt9yOGhdBzTEvH6BOXNLhTYeKPOvgmr+QLeih4dv7hpv3sG99ycn4X7OmHj+sBs
MZkHT8KfGd92PToLDX68vAt3B+LAFRNkvuB31eq0toV2IIlflQHJnLdlVteHgOzw
5MERdbeLrS3Qso9fu6K6v1FIZjboV47ESGc5cumWL81fTQGYrhPGqIuXdulLozA3
VO1DGzq54HvAehHI0g/qcYhOwCHdo5aJoAylqbTyzYQuoyNIjLoScIwfntI4iPFq
w/8+jZ6AytiZZjxQK8mGrDzqHhJ6711tPWSmryXUJjImPnSQSVpDrrjajJlMNFIL
hksL2o2Q8PWCgAB5pdVDgw90+tthiZDJQcL+6AmyRoG5xQDRfeksxg1M/wPQsEh0
TiXO2ZfgecKaUdNgQTu1Bf2PkmiQFDfQtW1VebTFJyB2y2PTq1izTJBr/vwdwPpa
C4uWulVt3Qk/0nb2lwMGp8BT5bh7NIiyQDSbmJdv/53Ew6SKRLXRYBsjYkH2bkpB
6FWvHjdnD029U+E/lugMVcohqhATaLxNHvCXn9X+pAZ9JHwShYQ5es22QDsTVh69
OviBAkdAkMYsT2bp/Jlt5F6Lyu/r8gNbIzzr6FvSSKIcwZlqcwJHoA5dFdsYTdXD
/3TDAn5LEN/ZglQVuuhvHbmc6BhXnvTVRY1TOvvorRnD2Qt9U8o3HZFQVxoXZXi7
WH3IhL3LQBXWbN7dziWlKLTc8Qj1Gx79NM0u/DR+oARIjsQu5oGdFF1pJa5KtLWC
XKyfBi6pHXwnRRLZA1WYHAsO/CFsJx2x6J28immYjiDdrl2eHpSvdfYzBbEJQQKy
79kVV/OxjP4NoX8ubCOLcBt1171xS9mPV7S6H+KjOYRY2f4r3sepyhqrTs22N4TP
uwsw01OqKLRIoL+AybeLwzA8yEojwwOfcpBWOvaJ+XhjOKEuEYUPjpnNjET6bKTo
Etse67/Nmur/k/55vL9dzgLEwJ8/kXrsWG5DafNTmkt/y86Lp8dFXlHWUus04B7S
AKFL2Hf3NDP6kT8HFEpteGIT4leqLYxfw2Um/BHNbQZvByYbrC4kun5QnLxW6BMB
tu2U8r9YRxqn5SJ3YTbuAB5gzFyTniw9kQelnJaDSvsdfFMEJuYMlHz/Vg4ZTJZZ
BT76DJTv8IoKiF8bTDg81BoccfWzrVez32HUm9P+klfCVf7Z8aKUUf1EJ0VLZwzS
sdDMe1/R1kUsOcHApiVIiqkHPXYr7TpCUBlsPUo8Q8KJEwJGnzwWqRwmq3RW2MBD
w90JvMSsGAy+wA3mxo+CxHa9e3S9QKfbtmr625KJ2H7vldtx+VolpSxHYHS1cA4K
68p9YmtmsHzQmd8oC53FRD2nBpw6Z6/2yx1Yta4xJ6N8XDnGghpBW6Rx5oaUh7nv
2i8/xYNVF9qC6GXpnUjZ5O/P4/UVGtcAJaM6cJ2M4zjXwgmJTjHs5MmIyu+LizhQ
6VqSifP53SBQebw8xt0yGR6E3bYDHeAWfoGfHLYtbf5sHVMuscE01wb8LpdrOT3q
tesPqONyasHJJo4iZ2f4GHmjglRHk9WV1zcN9HUtkbnsMRJsKx1OUo3x3s+uJbmo
yGicmXdfO6Qj2JG//6d9B7l5YYztu+2Ssw2vJrq4/PV4RdN41B4SFFNFNZpFAdoJ
l3nsutwm0RCCcskHBIf0g7zqkDzEnzgVHDfvun1F7nOB2MHGzwruEdcCrrw02FUh
TMZrkCbQpXM3OFtMETVweGExr0BpJgThQN8Y7xhFf8fmvxnw78ded1MkWas0aile
SF53ackGYJQjMhNbGnvkcJvQaU5zoDyhVI+HBLFC3Di7zd0iX/gc0mVIQcbTj0j7
oYiqGqAhhiFZDhr07sHXZOimsSFQT7mW/ZgmteE1SSFdfFuhINTxyFEMVbGGC3gK
7ovvkZWUx7nnrI34ILYtcYcPNAcq55h+0CftDlqfMzjbq02xdIhu7gU5b90v39iq
ibtrMInDkqyxU7DG8oA+cdBqJO7e7mc/O+M/2NkFvMuyUFnionW8bAoAzDnoqy2r
yCCs33/PL6Q5jJ0U7VW55u5bSeSpEDuJlnHr8XTwh9GTsiue39uuNNA98bwCXa7m
rJC0CSmHIdWrmnWCb1ILqzs3Hy845/GMkuIxuGzy2wLglzYBVcl0K7hjvb48jEeG
vDtpEJwWjvtEBd1C/0G+lDMjYhtyzVhhmJdtf4bL9mr21qxyAM48yHvzwQ0xXwql
Hkp7uWjhGVnBECXUGe9ayPCDsSrR1ItUxRI2t6FgPDBWyM/fXIG8wGQGv0vsHjwK
WTZXeSe31S/1dW7XMSfgesyFrpKJ44YvZy+Y/USY2j421amlnoXCCXX80V+lymbu
uXJjdX7fSMl228CFGz2paGQjqnv9gOFfEfGQWK+MqT8wHlaF4HERBHW71W4EsB7O
v+tLkoXCyVcEa4NRS6tKNUKGed5tz0yUh9+EIc+pvO8BEbcaKaeBp3/jSxw2Bl7m
ueLLg46Rn/XHSHugiIZCxQprZNF5ZxJA14nDpFQtJaTG3frcAypRnzQa5Nll4bLE
UO089WbcgG/J6voRlIdJSGnX66wnd0wxTjwaLKyJDorDYIqG84Z2h+80NKZcWUNO
ratFUeEq6L8cZzz4AAddhZrgyCh+deJJW1Wh88Fe5bi2O9CqSEW1AZCqnVNsxGRN
2cvLHaA2jhuMiojVZCJEVakQG1cTlfT51xZXwLCKNJqD+jOjPOtdghOpFnVHdGZ1
aSsrBYOdHIktDB9bdJvM/d9Hj3z74/QNcAVrUd4a0EhHkc+R6qU1JHSnup3Ujd+g
9ypYwLDbdNJbJ8Qf5ID5GpPuZkQGuhwtLZUsfKkzfC60U7s2aoLVyyeGvLKbuPmu
tCez3+AOkj2Z91QgxiJuIuMLDUR00MLjZoKi8yKIDYl1X74tzuQ7+B6tozjYGXYK
pk/9EwrljHD0dxjd7GNDwGn2TTdYHUgm/wtjxYiLPaTV7VLuP9W+eVEgnnXegKh2
UUw8Ce7J25sgQkKYGCyW89fXPtedyMn6D8iyEBij5gtQN0xvS4P6pInpmqK/U017
FJkGDrecFTqCxarsCiR1ifO7P89MLgcbECHe92zqTVWkeE7bPMJ77pNFgt4KdG29
IMQye+Ul7iWbx4K7n85l0nNtt6x+3LndChQvMlqHl4euLBGF/e+SOuRycqE3aLFv
c6BeSbRYMrqYhkKRtiH6X0kkofI6T0CKDncuD4+vEougxvIdu3cQOuSB90OZWOUU
uAozclODa9VVgrfRKVhwzfS3NtjP5UvW6RkXjUipTZ3PwEyJnKJvIaifvxV/V7vu
gkXhMBNgg4k7/Ns49jLwJu9PkBtwBL1sv+4tyB1Q5S4zcbNIhoQtQyDNMHixwfsn
mXRRCqydDfRdme240r4cVofuhSU+NRK7z8ASa0wMOiiXHMOx/JXZPP6hq1/sNqmq
7Opwxn61eYWTqXZlILly303dnfErDIKiqmp5SyHVsIVYtI/Z3V5dQMnOV7bV/IrQ
op/czC+jLn4LQcVYcj9G7ThvlUP3UIc79BuEfev945UB5Xztk4vIZLVPpiYu/rN6
pC0/U+NrwhPMOkPAKyMOpwXCHU13pqhzvcktF0m+aRIAgEWVJ7pkZNVmM3znFRH4
4Y30xFzZ0/VH/Er+F8d2OFjQ8rPC+3y3/riyyUWDrdxEHEemPQgG7BhaTjUCKk1v
hFsmu06c5ryvfHNZOYtBBRSEfJ1lhB7MoQzZdzZfOmW6mfIF4rY2JLAenS0CwYUW
Bk/6dyTI4q2iMc1gBt9wbzmYMJZueenFjcpTysUMs47ySVXndd+pLO9Lo5inJdWd
HFAmfP2aNGs5C9oKpI2xZ+IdlXyOo+SORkIO1Zdm5KSNBGWr+ovMNcW0NdNC8hox
cweazNpBxnuPx5EKB9MPQvGl5O9uE3e0KMcnzskZcZXYbr9R1PIAsy/R1QvGuu9e
uW28h/siPF4g5dDpZ9iHIW+ByowXzGeLbV5anWh4kXtIksKzgtoPNV2xRssiwlOy
dK5vOmi9Dhu3af2OvIUr/o0uY4sbJ/hT2c0V0lFbN0Ej0sosl5ZJhqwUOyLNSzLO
hU1mZpRmxGbYF4S7+o3s+fOv2qLRZyWx9ULo4J7GKFOUj+mCZEFu2luYWIbg06ij
gsq8q4WD0Qf9YHYxbhfV/dzzNk0N5oHAMo5iiy9c8lvgZMVJRJtNWGtYiRfpkQr/
8dk77zNOlU+0f7h9dlUh/Xp3e8KINbVRm+ylJ+ZdobYK1tYkOYz+6f+w1V1ErPS1
WMiKMsBtV6xWxFqady6sk8ON6Rjk0r9G9w+7k6xqaP0xzNViFjyzZHaNtLlJncLN
lQUWazlAJTZX0Fd0v7B+ahKSmuD2kjzIOTpHjvOLpSNOjtgKed9d1tC/THxJ+edi
TEe41DcAql3IS7IGU2Os02lKIUgfNfUJuxN69BuKdKbu+QvqjPmdaYpw8aUfHNYC
nlGRdCrtv1bL8vdPuYOJ6w/Syi51qeXossltClp6GAiGAVYwWy7CrxLwc3E8P7br
7MG2dnU78Y3wgSt1MlBTu3okpSKRZe3hTonppL+LOLvYjyJKQNCPJ+lPSUlCB4l8
Am9HuQaLpXZ1svk2NFKZWng1ktUkETesPUPKzS8NhOgWKIMRqkxOF4L5dm1nkwxO
EMLC0l2yG6sOjziRcaSnu37bEo7AMqqrMr3Z+QPPZSnSUS+vIbX0q/sKtmg9z4fK
L0kM19RiVeLwslwUt1xqu+O4sVNl09hlMv8FR5n0VIstEKswrUHt1gn8Jw4hleV3
dxQIqrSt4ekFyQfQc72Pv/G/nzNG4W7wYRghuHDYXFlISS3HB9oJsbt2gy6BTB1O
QIs9ymP6XZkA3Py3iQTJ9f4AwQdP6+EbDq03XhDFxdgQ1AnUZoPRwecrtaw4youp
kSWqL0AUnnvR/wg7yZIO6AYinDFTo9dkOx64fIhA6ipjsxegirV2sjH3EY+elM0K
s/l1yV7BOHEy2ejmYL/lTz5/vw5FVfeWSC1z23UuxWBZ1Z6vOTLP+ZfuYRY+oz1X
GCUw2QTw38QJ9JA/2hWpAhiXr2PMpy5LflgFGDVjVxAPBdA7F1CA1ab4ZpjaCSRD
tr+pCpnwvK7cnr/Hp+qdTWs25yuNYdSxr/2IXwlM2v1C1yFYgmgu0DzzSfkSbZyC
Jo1avFFrTtz16u1/2J8DHtX4mSUw4hGz7RP58ejd2Lxa4IJ6nEHCC/BudvYz9Hgd
4CZgq5IrXf1bjLjlNjStES8tmdxcNW02LsTopNOmimCgh5qefqw5P/w4/Q6GOEOZ
q/ceXz17yGOLsDYFuzZDgzi/uHHVvB/QPACWv0Y2/JPARdWxUF6YtuaSgd7RCAIi
uKZW1mItqCsIWJJcWnje3FgRGaOLYFf8t5VYsk7tehyqLB91D+CrMLLOvsFKI3vT
6LSgQy0ATuMElD0FoezRqye2ROvpPP4yLhbqtd8AQukhuqFmH/QwXkKk8ZSsUCGA
a4F9iH4GG/50E9VnOYl0WJxon/fuL36qwkWDDgamfqEBcBh9XCBqHmZj+Z0+Vv6u
g5IAlKP8eHS/wjPXo89RvVY9xAtWGFZARaPIdeNVN1CTSuqmaSlguqJdUdYzWINQ
K04iYHxxp2vJd4MDDt9JbHpBj1Glle2Gj1HXoVm80bACM8qhnLs1GXSmWF91q1bS
BbtLiMrkwuFRGk+VPcd1+60y+495dSFfi2lFRWlT4gljVGBiLs9hQ67LEiMkF3Lr
5Y735ZfqFwa3jX2i5UtfKVY/yj4QxcqWBR+afygCnGcAQgBd1AnY70KeFiZ9ueSb
cz8K0u8vNbjwJMK7CIPcba+sHtYk8ybjUB9HqEto8EeDOuv/wW8L3Y37FsOovqZU
jX/7aDcM8Qlyl10Chclmiv/SLokP0UORxx1zRTaCqW9ceAjfV7vMK2a1BhcfZXJ3
mvvj3SHLJjhJJxLXlpDgkpx9lZkkpviXcI+nXu53rtV5zKj7KexhM3R4+Z8Ih5uw
iJMT5TlY8hzXj58NyCSTcIQamdQYfodh+ldeWKfBWSMXdJCGAkt7X/inKWRqQpj4
19xrh7HWtFtXKLAG4CbTGwv3dy7YfIHiLsN5S0LKqeMjlHkabJvOMxnmoqnSXuoK
vGx5ZW1+Jvt0uyaGM59sjF1hpzS2XpvpEFaCa1HerYUd+lP5S6ZZ0IhhqyvmJFx7
vf1hqZkrM5qvnK8db/UswMjbNy/77y/ZAhlVeHg5t0H1eqB14yZnf9flqM7BFclm
LogZv0Xjc+Td/a3hVk0HHw70Y4l3LBPyi31LthYnfSnI8S878og7KRpXcdL5mBPZ
sPAuCxRLeJ85Fs4EEiAfcC47mzti6NqrkEy9ZdAwDeOcBp+d8rx3aNFrUiF2IObn
C4Hoezc1Q06DeWNHCAau6b1EHEdEqwg8dFBT0GUDFjfwWiUhEpRtBLVaaGOHSJm2
ZOIv4HBClbbfS4fguYqxrRvdrKEwa1VFRlIrMmJuauvTE3nNvvP7+/LpqtCB8Jy7
1EAXtZkzJvYFuavYRZVBovfDlL/zTXTEblLLujS/vMDX3k0UElIDGEXkP6kDMR2G
gvhVuCSa/SpG+UqDN9HnUawnMicgd7mdvmD7KUNw8Npk2XvF5zZIRd5v7QTvuXQB
xSdWeBm0js3OeL2Ygd9Tqlnyn9KcgossJzKEae/DXfX1CVocf2Sm68yePXmH6EYF
r1VNTseqTaHRarTztSwOy/usWwt/Dd59JU5rtD3XyyVIF4nxwom4ghP4PRX37BgL
T/riUFSUC48vXp91MZcc9A5tee/19bYi5rmYINMcC8G6USuWtk7FC397JZZkFiex
HHyUzV8rH7mFG4VK7xYdIY2Qy1XAQRmo+eKgTVZWPFu9NN4SYiZtjG8427+m+5vV
8lSTuFlDV9/WD+Oca9FfaaycJqCRYinaDJNtrCuIjQWsvMnDl5siOSWo8t88Abmg
kRIbmSByUxZ+eX0b7r/Jwq9vEnUbN7++lSNDBnkYgXRrZ84H8U6T0tdk2IC57X2r
f2CLqaSw5cJrOKRjflrbNLqcIKQke/m4XXGDj6+Ui7n6VIncIiIId17d6K7DsS+l
yQWhdUGSl3sT+chKBpTHrMphq6KOQcWKAjmkuCa+K85ZhxP0/UzEaNwCCvx+BwpU
9gnT0VBpR5ACPOibrVlQ1AhoUpcPeixUsrbSXFYsaBkeNESkOGZnk1kVP8Btignn
RWI0A8NtVgkno/HQGF39AB4dM/KMrTyhLRTx/Kz5OBzo1EeWnQp23kCTp5e+/u40
EZeioE9KiAqcVjGpn0ZRI7uDkgQqeBSWF1GofkwBTuBlWKoqSoxDX7tPw1YXTcfJ
30Uac1XKxDo7Ibw3LzQtXuuhT0bHTwYovCf9oCFQ5Pcsu/t1SD9fBmCFzvYJ0CKi
PUSZzbcT/BTZJ0p0JXyF4NQQ0Oc+k1tHecne7aCJRZd02IDZsK6ArwzdE3vfkt4S
jBkL6Txh+37c26dz5GNYmMsrZPhj5NkDidmP0TxTvvu51jrR+Sa13CWhkgFWK5Dm
Pt2fBzOWnGGYLR8ZhntcrBdRiZIqGZbOdJWEboPXxaHxybncXxavYkgecctL20Rk
y/F8qtXzqtUw+5l3qkXp0BGGucatZl8CPNL3kuAQRmnY4onJA0JK/+GxiKqNyeJB
6pyZN1NayaeCiXZLTwLK+ypSzZdXfNfqvvmRyUTEk9/YoF6jlbRmqO2vwM41pqQ/
mMngvdlf8JSJAP9kN+DFn+uTLe3HX5Yk6w+njRIwA5uyBST8vWBvZEvAmcBr8lqp
tuk9mmcSdUIxrfbmfXiInlJQSuEdiZJ40xNZ2bbtZg9qZ21Txv91/ohMIEdP4f0t
1BKXDWOmXJGkadOOzD+Wa5lcLETTmmelke6VXMPhIwyZ1qqB7erpafM3D5o0YLq5
15IiBsjHIsafFP0jM3G6oI/XTM6Gu4WKArKNbe39RYfF0SOaPz2SE6xH8n9481zr
wYAX69yTHlQsmyxBxFWI0r4sJTgfAMOXyr4scNqsebpU0k7lV6px6QqO/R0o92kB
2pSRVss63dre5+YeEe8izVfWnI8ZD9vXogFAFo+mDYqaN7CWIUyjZ8PX8ANXul7X
DJWRVIJ0LT+KfbE7PFUgDHiQCn3OfomxkHVyx3oWFc+9N6mlSS0OYwJTGj2cNtNp
d4hNwDdrlqJ4tm/DCOeetbcj+HikzCw6BX/e8hQsc1IGJIBX6EUc0Ha8A9miiIFq
L3fzJY4xkPj+f/xNPiE7qJIgxaHrKSOFj96czIejwZ8eORmwqiGy6kdtqiPJ6EV+
5NdDW69K1HVTrNvs6EOjyqjYf0H1yJNyTuc35VS70kbvL0wXk1DOR/cCajFY17mH
1KcgRyBvB7cHZAF+jq1tnyKFNnLWpnmR3u0PiWVQxdBYYNttOwzUush+XHHq13zq
oNDQDdU8M93JbP82YOzRESQVG+xMBFwHli0HiztB/hfEvHV8MIWuVsuHabgO44A3
v8fQLwhqoBvkuDNIhTsVdLt/g5T6m01jif1BPvMcgy3amwqFZ112OPvkKglH8Vpy
5LRBoxPh+xXlVUM1/Q7W1cPRLOmkNcmLBCK/jly0olbSdvDbyIBYXhuGURiaTkv+
e+3Do7idbX/PLFtdhAVA/H6ck4F2AphQNQDmhLtYW7yBZrpKpjRROJrGcf7EN5aa
5/mAEZBNdwulN7tTAXz3nXcnR0NGrF7BpyILLQV74V7iAgzzGBYbzyav64HmCz9i
YMgFSTmtFQs9EzKY908hl/m5z8juWgR45vixKxOqy/r8UmlRiL5pUD0dG8UCOxlD
cEM8XEiQiE/S0j3DuHb91+J9xV7cq6ycm7jvK48TFSWSZPT2xAElKg+t6DCLjs4v
88EpfegPDfeh3OiSPpPwfwDaxt0onMnImmNv3jIYAkieQ92MzNvuOeTbTpSv+tt/
THNAV8d3GdtX8Y1vZ53FYjBAeO5oZ+LQZN5zWQNvYCeWkzjZO26u9J+ByU0jGdUF
7SKPhMqypf406MTqIEXk7C219i4S0Mga7rpvRWlH4X7lv+qMam+HFA+oRJA6Epm8
o7YgcXSgrI67XW1dN4H7LU7EOSkCyxGicPLDA5BQQW4gnOJMRdiMfgKnf/k1e3LW
3tk0FAhU7QxYf4tazhQPAhfObBtcqUv/UluG7TI2SgdKbbbBimTE7SWZJqztJ9Ml
5fuHfETq3Vp/qMS75fbZ4L1f0f17mShw98XZ5UbVg6QrF93/ELaW5SUAYornLXp6
91O8rbKKvZpV8z5ntsuSNj3DFFl7ZtqJ4qrRz4RLDgn/lfyyoPogR7czEQLmn1sf
NWC0061GJZ5l+V5QG0Imw58+rmrf8pWp3J1wIkfer/7o0hfPh39qXRmiKf7/7aID
7aZwsoPEn+L2+/H192YUMaJeb3adewIuLU4yULkSyOh/SRozVuu0dgOE0jKez/3+
rWcrqeMN29GTbjxwq/Q0HzyHQvLe9C8r/ib6PgD9LoFslX23I1rroKfrd+wA/68W
/AgEc+3NVkU+9EicLoT6ot6pN14cp4nYP7rWsY165YRJNlELH6oGC+8uVbqK+ELA
RI8YJWFNJPZeWL5QYDgbCjCVXY0mNyBROx43tOyuX6aid0J14aaUayWfhfpJDf6Y
+WZbpZDMlEydLct0hp4+WZpOrEt4qw2zVHZ9DrniC62Rx7UKYI5lj5GFegLPfCJc
uyAZFzZ96ZsvzJ85xm+ulj3X38h4rSeUvsfOaYr3bQg4/1QY+ZnxI9B7mYeYN0jT
/4v+SXlgkX74b5nuytosLsT2b2ZzEofGq4mqwGmm7TjoiE9kaXICx3KdRV9vu030
aSQpAOhYVGUMRMvYF8E4ZfdHQG6fCQAQ/ux4zowHE8CkWlcwz4wkUSA6hqJmY88Z
zeIbULXsYaPnVyz6y3NFRn954YxP6I/tU4g8ggBkyKp35vhRv9HPdMuh0WeUcoV/
OV4zvGwSHwqHe+c8Kq4tEuZSHxNsk7OwUce+au3gB3RY4vw2DnYicsHfPpg8l7xM
QeHqnjL6UoVcdlmbSXSiscWIEF6lsvXcsoLh7l1TXyGosagJ9VhxCtZd2VMlmX0O
fBdqvuSDvILBuXS8nxw/k9MgImRq9T/+i5v9WPnIi9RvBdebIdREilKLPMHtT1ck
YuzUI2J4hfJdr9um+9Z8XREDu6dv0j2Dk0IeJTATNSJeaOWRMvW/tFYIxwy7iG0a
RQKEJoZs7lIpXq/Zx8eacAH2XfHK5SxwsWRrgljxZV21k6QYueD32YZQXBLzPPhr
ZlxJkGcTFOd/WIpn+HWcz36v2uvo6W3x/uwBprxMXgE2bHISrjlnRiCAJcw+Cpkw
DswDsDlJVWVPwQFK7aK1ZDBXJ3PhN0mi+6QIEqLFyY76S9ZSL7iJuW6HOBmjitMG
DCiUwpF3uR+tgc3K5PEdXYAMLhi2wyEHON+k4j+QaiyGD083lIFQR2tn4ppqUg3I
Af6uizvNeGzoslCebScTQMeubT3ePJlVNNOAUbqKTk97m6iozfjTdDhUPW8uJVd6
DpoLtlXd5fFQKUE0oHP3b/k1lQG10mZe+lwZD6ergydIWEOAo9t3Hby+CvkCs74c
eRy0ZbAi/fiWQqfo5evJ+ojCud0Z97iXiSn1E5uwSLaWHsfFhaaPWA8++LrAUT1U
9B1LUH9kK1Hi7Sggi8EglDhmKihsBOFD6pXEYIF3Bekyex1KaZzToSb3mVdYfGcO
bMJtuQWa9Dq2yOwWEOEQMWL1HL8cgt8fBRWx+wXEG9NqHyTejC7QE3mYIYzTweTS
F/BnHP93vKrtAKvO/3Gnj1szUUgqqTcjoCsjDyGeT4MJFDzmLM5kznKHtikKyE+E
zDNC7ll78Na65kCRWYmmn2OwcEFWJFB84C5AIYHYEJ49haDm3hDNnCBJOGOlLVCQ
yps8pNcOQs9GAtp2jqfObSJ+fWJ5HthxEQkDt07eo5MkZ3U4CRAxnHAtOu811FBQ
wi+/e/9rNDK9BOvRGKjW2Df1OO46i4cO0bBoJ3nP2M8NUBv8i7c3e/t+FT2dAQLh
NgvGxrK6ZldaXM2a/pkOCp2yNEQzbw1Jj10dGRdE/UcsODCHy9RyTWXqiax6is+M
zVHhVviFbpexx/F0ok3LByiNfE8rNkxBjybqHLOYPDNOLHE83JbzgGJ6roSC7KT7
ZyfExZmtuCNFliKRr7OEBjZSr1TcnzE7v8RTtze1xAsmnZmMD7OD09etTUTsWxZ8
N9k/MmNzSfUcP4Xq2swPfyTFaZ9/LN0QQQtiXCZdoIgsyIFf/ZpGmOawImf/VH+M
1sm1Spc7JwFV/fTabCdgyBJx75P17wxodYSjwGu6zSjLv5p6EGx8hXJr1Ww1KI7A
mOODeW63bkcl3YkOeTE9WbR0OYiuc7MX7pMJb727+Os+aZvjhwDFQEBmj/KfNTpI
IIySEbLChW8sc5ahP8JzTxmOZWtWq6StoDVhlgefFNejVNksf2XTlwzDAPGCaMpW
JtsklqAVvYiRCx5wjubDaijVN+B6eGAY/7VF14H45O9X+ep/tqYRR0KGTrU3i6Ma
Le1unNImJzwkOhTRFDz0KAhO2V/f9+m3CUKrIG4wfAndubtf/zBOIlq+dHKm68o0
rEomX+jvbsAbUSqvbLKJfuyvK7ab/FxUT08vkPu56psVBhsIeRFo0/GgFR3wzAkY
52CF4whWJOfW03mhgw2NCj8eWJMJKs53SzaVHCf98DkrYuvk5nYyj/+2Vt5PkKN+
jRJLufbnesf+dUWJmnBUrMA0b65NqYB5N2XFiFPVTJR21zX4TdpZTRKhXDUeTbjm
r7oxGYoEjJ2JQqPYm3DJN5d1bFjVU4lqYSI77RJqsyGkgU0uf5jfWgfoGVOTnVUY
zUIqpl7cFwvd8vkPsqGDJqd06MAvDHwlvuyrWKePPKcrQwnahU4nhssWFYnNdhaU
Y7bQ/i2bVBUDasdz28dyASXDNNZgDcv1Psqg7+ODRWCFD+h5Rt3YBHCY5mszBsAZ
93E253WMbAXgqDm/u9H2lODxKddimNtb5PeCraqt/NkHkSYgfp8p+ceq+DEtBgMJ
vgS91yl+Alh8aJuFJAzgVBGPnbJxsLPcKYub5yIVM+CgY4aJUMg3nRgjl+69BLIy
+K8xagmezTR5uuCJoUd/jGPFRYLKDwbOJVH+aE/qG/B2XKQUe8uUMrdOXjFk4JBS
vIropYjE7H8mu652nXM8eLYK81+tIk0d7YWJ+IOB3gQfaxH9AY+GoncM2pbz+plY
NNB68WpRvmST//gvlg8WRNFWUBnt4dfFqKTg5tzAoqJgz1s/tDt9JZ0BkDModuuf
r5CwzpWT0NErIqgfuNq9wQNiJ1pGhyO9nNTpeYos8METNTNf7vpBMp8hsl53qBJC
K5jpgLtU7yyTAUYL4V55dqb9C9YBqvJV6VLquf2/cg46feo+ZsjPBVcPHwtWU39P
NnH8tOTslhg55/MxB/UizoNEGPeE5ipE+1OHWT/oqL0VlRf3Fe/Ckq961G33Pg9J
1dZl7V0ihGjESVUpHwp/OTo4BNxeSpOT3gMkDJdj8thWagPSwEa3WOLeeia79naY
/FrHYq8ek3t57Ps81b192JnrH8Bc7mLOW+u6Msl6pcXKUkEO0Aae90jxaZoSia55
kaIsTJ6UTPITuiZI3tkXruNS8YQB3Xoky4/pDauG+9l1TcypBcYPJ/j5qZpZR7Z+
r0ycS0h1KCIHSXRkWi6Z5eC/FNAFKQT3+LwX3rpLIxu6I4BMY/aq8wq04eLyzDzo
GC0Y6+dvw5/70708iSuJVLix+PIwmHLcLIqfyPraFpIxNswlVjWeXcsOIS7PNXvZ
j0r93Tb0oqZRDnDD7BnLNE3/JzyVf37akbcwk6noJz3avBrynogdpK9b1Nhg/PCB
JGRXF+/JJ4uR4KpOuZ4BFGMOvKKYhfIHoxPt59LYZN2Ar/n2qyXsFPOBV6XRhwp9
W8YsGSeVlVxNwgcXuLx0avIcwBflt2kL6/cHH7UeIGLJ4xKELbyKNV9nX9TD+SK4
slKqCjRc320E8IgtusT2nK33DlQlOGijEolkgwKpac7LYuUUFWOR3CDXruacp5Fo
unKXohDV3nLHxVuK/vDflN4r8WnsiRl6MMjYaxZo+JnRCuN3tx5CORKKqxncH78Q
/gJjgKBJwM/s01EulKXVnJryDV6ne7imekXXPVccwWf+NA2Z1iT3ARt7lkT7DbUf
xNPyNIXS8OMFUEmUP0shzUpkU87/neXrokPKgtKEFv6ZNKgitdVc89ew+kvM5fVb
JXKbBkAtjxjltBO8h6W3XBan90D2I4j9qrn6JBkDJz52z3J3XEIIAu/6ARU6gTvD
Mfze55zDfmPELq8c9Sq1iNTJ3hJg+nuLDSqN0y8Zk6rMfqsivyBIobsliSWljfH8
QQCNbV4FP955hXq+5pjAB2cY/u81mygnbJdvRcaMC30U+wIe2Q3ydM2ogUlAsQ26
cXeR/IXks+x8sY/m8xVMaLmybYeD+hQ3MNGdIwuuQQthJPtaXCHcyB7KKJTTMCU8
hD9Q5o2rQtvqv4cjnPGD+CBh3TfrpX58TCzcUBrgUW7cyqf/Za3vZhP+lNFLU3Jq
7nXlOAMpdMnOvvCz07Nx1LlZ3OxA4A3IivDOMLnjXAkobJ3jmAUycfa8pnCTWXU7
stNtg1Ky1rj+rFUXhio+jQzyZ/f/8UIxhpplWX2w7oFPKw8oR54r9gOb8CYEiCYq
P791CN+p23qGV8nHoeIKRAdy7AldTwHwFgrjzun/QWbRsnXSEgLFROeDf5tXHBOl
B78M/4F62AdHwTI+JsHsJapvPT/8IkH4TYcezeobvDSmwpZ7kxYm9IRqKrXF9bHp
y59ZoQSeAJOSNget/zSWTOetn3bBq04fp1kZf3Jqh3YP5ciBafruJwRsoLr/Bl2+
OWN250057+ZddJf+SIiUiLQZcjsl2qJZ9J+qcr+PV7Zb6WdmYlB3gHCKX6cdQcQ1
zFcmInkSLhNBiz+pUuq9zOit88whpK2bEWOOYgSlifG+VaeYk/Wd2XsLwv/3c/0R
2WqTA8dBoY6o0/QAoyoBMdLgTo/B6XDG7HKQvXgH3JxhuwiA7CsTkSMXPu647uGW
pCzyxtxCJG7jo1cj2teGdYf64zsGGxVwqXdr6pDa4/wxxv8k3PiSNwiVkLyVh17u
qRwMFYHOV4tYZkX3QT4JnHVrUewzyFCLt0fIBVo+FOgjP8L5yztXUM8cH7fq6iCP
HrO8Fvi/+cJVZ9/DtIq5MZz08L/lc++iX0oXxB67ignzSy6tbGPnNFObv2XNk4sn
DvUv4r61VK6ImwOkWT2lF5wMiLF13NL/s+fIrZD5eEjlc9Q05Bv8kGMW95K7TgxY
XFQGgcngo4BeUv8Dlkh1xZAYq+AsMyG9Ev5PPhVVOvooWi1e6hXiReDMoNsOT2ph
DNVFmDjkl/EvuM9XjVj5tFW9/kkxZQlMzGPb/9nW9f0B31/65OCaj3Gg0gAY6gAZ
vWxrDjWQErmJ/utl/AuCQJfJh9l/wnmZOoEiMp+9dtbN2gsHhgucQMZzh8wz1JHj
Ln4xV3WpYqGcnvoeq2oQ2q/FY6a/7BtPF7vMZXPTttPJsKXbQpRU/LIpEia1eCsZ
IfD7yFZE4PQPv2K6asf+MILriuo6m+AVLpUz3NXcg3QQjuzXgell2pGzWOV5KUAY
xyaLBAXSc+fLuufPKw64AQ2b1FpsnG9fbkMYWxNNwp8neMXG8c1b9NH6w3qicXYd
wDGl7WudjBgw/7m3zeCL4HUSCpbP4d7PF0EI2y5VxZZgRKfPl1ZZjWesAHkL7N0V
hWyWUfNL2lzdpPCcg193QIwReypdxNgk3DmVMTyRf5hf43aiHKphieHt1cxlGHm+
E39ziFKnKjh9HdSc9dJpl8IBXnBzXThJ5gsEA1rz82gqFfCFg4FkxotOtgQz2Mfw
lgJqWp7uXinp/VHPvmvFT+HDpuEA+FzS72BeOp+LNFiRzDHwSykj+L+avANS9LVw
yubAIvk05nfYRLLnI7tPRjAH4GOuJ/Ps6YfdZqB9Poa6SmZ4Uo+zFsPKsJcNkcp0
wbar3us6INn8pAlJodwUl0BD/tTFJp6xDc37koiZPLUS+gye9iCZk6Yrx2pDiMjH
QsEVhOBOQfTW9y5Zv1RCQL606aHTyCL7wgJvQoGbxCW5qVqaJOyXnSuOZB+z/7R4
r60W/YCIYY0iAxfadhD8g9lNqf0ZmiAwH/ELWkuGeku2i0cB+rX5NFlQZWhao/sM
9eaNwNx4nbtvd5yiRb850wZfLXPKr7w+0Rs3vrLK2j415L2pUsrtEwQgkdozJxEM
WJYhFqtTSgZsbOB7u38PcuRDFPMxBzCHE3MzyhPATwKXkpFR418CvyeTC6N8yJAb
VKIPD8QrXgQvlT9zfxlnOsP21hFubOXZxNShI67CIu9k2KRqpWelvvU3Yn+iWCQi
19LgM9pr+deP46qJzrY3yqkmraLSut3J26tB2YsyQ6Iw6wzUTALockHvM6bg5Koy
Hug2NZGUlbDNEgLhGWjzUqAMS2qpJejJKTi7Y/5SlHTFBs1ZrFlMBF700LGSEp8Y
HQ9ZZLRXHtlsSGzLyeYAg+H62ffk8L12lPNeZ2uNQ2hGs/z9EZXUElZ6aNPIYw8p
s+TchtTa4VWCKW5MQUPKgH+XAoU5M8u2b7TXIAGnJu4Rfbmh7baqvXyUOkzsRQLB
nHK5l4WpLhFJmpnafq9QGnXBEedwxEH6FwmY0lrEJ6bGfO2YxtEsZjgodKqF0e5E
fB600c+FfX/JcipeKVm4/4Dl4lgJiuR9wBcEcYYXino8QFCxT7BzaoACAIrhcgdz
mSbdmYpNknNhPMHxh4tT8PH91q3XQ0OUviJTT9gCq16Q86WVhXhodYTU0S6KjHnS
Bo0USKxaiQp7xxWBgg3+uN1a3jd7jhhXpzHYEuWvJAOVl11OBMZA0E2ifCmBTa0K
GnO8hQK4OwvzhN0BwC49dNcc7qkkGZJc61UHv/EkiFpOsQaWbkc1Ii3t+kYERGNP
WoFePP+JK31vztUpq22Jm/E68LBcBsN222OiSY+u6wMjsTyAxSeq7AYD3ywe61j7
G+cu7BywVKf/L4/DW/Jua3aQeLPOMxFV73j2kVQ1EC/pFEZQAf5qyO0FBjX+0buD
FzEaVnvLkuzZflGP0jTJtqrEgatVDkjvdfGLWocKFFp6n/wUs8Fsgb6wb0fLxl9F
idxGEzCiUZkDPjf0Nql1tATU5f6oE6BT6w+OxQ+Q3CacCJj2/Bwxa+cDJhn38/He
HjAkmJc37Fax3GFaSzLR9R+wLgeJqj72ACNkwvIWCuxDe8HYWSBWE2f4uWx4ULq4
OlqBIkxLG96xPDpGP9xzPziwz2XyfIYTGgoMkO1nvLdpCqSp5W/2nFW6rYtnMX9T
B5Gy9H1s+3qo0TiTvZR34nkhgevbWBAwya4F0HSGb7todlrf7i0k7XVwoHHRiFwk
7DzS0pzcO3wNqDyw/4fUd2+4OXkk/N/f7laInJMbNn26Eujxjm2lI2f3cYy0RDGU
ZlWZTzFTiitIXvlRpdhaqIuCX1Rvjlzt5MJeQrqfql60AE6ePh7zHZb4hzfL5clp
qGMWl59kphCAw049ItzshTuu639R+C3V3eRsjLCeTIyPxG8+ked2BNLePWDIG94I
awBt79MXew+2wO9UZZIuih3irtBUUi/Y/zL1og6/WTFGVTiufRkUyGj4NCLQ/0Co
vn/7kqpOFTOq8u6ibu6ISFTLva8JHBi6uXUcV0weOpTflYLLtNxRxQok1DbGokEP
Ic4bOsKppZ1ZSV2AlL9X8z6kpj31N9yGgo4JblkRqFt8r3k7RfVitcW3Vs+Utb7P
l8xprxCj8sFH7PWLhVNAJcy3HfZw0l9QKDaslpIr1AB3Alj2R4KOkwZDRS6hCjZM
QxL1AIOody93Hb+6J1oR4JW4BNE4C7dDAn+dpkwmxHarwSBGB3XaZwlJ2rReseRX
qwKEgxu7q30bD2ttJapy6HVNhGg2Dd60y1ZUpJfiCtpVz75yprL+1EI4oGCR9FTm
oe97+xLfDgO78izGENp9F0f5ccnsnyQJh0YAC+w/tbYjdR2qEpVSWlSvUBA8ieMt
fSBvKwgVrCRwKg5FnekfZHr6iOwacevkH6tOXTKwLD36tw9XogORNdI4v0Dr2IXX
b8ghxJr2STER10blkSehOULhW96j4IaYwbwhvwPLImJgMdd+Gp81KDz14xl+Kv9X
/AqH/5vn0oXjyW3SswIR+NoO2UfmsPQbsUX6snCk0s8RMgHLcPVesJ8nOMcvN+Bb
X/JZB5/rM16ahpW8wSBFHqvsJ33u7Xqbr+7hy+DL9DyN4PDxOI3FbimnCy4Erxkr
2y7NFkkBYEdKT6lUE42Vgyy9qD0OtWdHWfMmb9s6h9dME3K0vUyWSANDE1BMrJu+
aSL/DQSO8N89O8JLx5An6gDagrIe3O5gxiHu8/g5PLgYQj+5fuGk7iTE9w8sNaBx
IKc3tHYoIGshfFlcnOcPBNMeKKGGSz21erdd1ARn42JKLfTUV9hX56lvTNXy6JUo
giJkkV+NpRaQAwOC/LKhQiQHaB2Xejd8ZFylVHgBTsFPyGcu3ecr8XPxQIq+LOv9
IMcpAVr1iNtYHe3ueENEYhe/M07J9z1NW2UwDFO39DQP2grPp+6I6Gy5zmZSuwtP
wfU6EDpdEfhu4zQbaiYyqOLeAv2IMGM19k+Uj/1m4Lf9fL95tjfKqlT/dv2RWE7O
ZBxGdSqjxtrRLb+l+2qPPLv2zoVh+jC+SNoxR94OKw2Km120ab5nscB8uQVxHnZH
Z80pW7nPYPm+HIYtO+Oer4GvcxU6iLTUsKSmkiRrVwClgHVDqH0TIjldxBoVgGmn
5gVR8wqFJr+1NvLZ0c3cC3QkRCgwfV0yV6NgK84X4ZVMyxIDfOP2UK/5g9k8Lhkb
WZm/UGvH5/nONFUaeeDx0gBkVANVsBEw9mSBHLwlZFlED9OKwPi8hE3Y+c3YcGBw
SF5y/EhC0s1ufEv+6QVMaFnsFAOVtt7QBzslVSJ0UB4JSHbnX5rNOTb0FVy4XgtE
YjATkTYUg78G+xlaAuH7zHdEho0zLoZqSlBjX9FbDVWZy6xAvR/olOluKho92iCS
6DAyPd6P5CJ9BTjh81QUJEkknXKpXw1mth8s/W1Yd6mQbEo5sjSlhk9PyEc3eCL7
zK546+QGsa2pIOU4LjRRQ6qh9gxCze99pYBeiKpGzjvsTBb8ZrOslx3vbKI1BrOt
MLR6Oweqar7TL5q4FyMrp5S6SNFwHw7zCGNW3Ek/LS7D+u5ixiFnq5tgDZCtNzib
G4rO/Zn0q2bIZuIX0dssAdwE75lQpEup39/22Ib1sds/JfHv6Jr//tcnFGl8yuUJ
cSg0U9KAa+6HFaFdzkWW5UTDLI+N01ESphTkxPVcx5IVWouTM7hB8MUo3XNh5ou3
dvuzsVSMB9YDnD/uqOE0odebmuEgDGlAhQvuycxkBOBJTteldN4Nw3wWxPJrC+Z4
B/CQdLWRA8yMCvEIdbTQtW6Rle1jveGXR6QLqAh220EupV9hvGJQAntl3K8XuGFq
3XfSv35CEQ0SNtRyg35MtKSVOkH9axWTvXy9dunswd7Rb9WBeZI2hTIVBjITkRrU
V5yflNlugSdZi/4ijAMxAPfIEbMtVmDEs1N4qSAb/iDi5LM2neisAKrAwSafiKI/
UEEVhJ8lW4JasWWYScqwmXssrGWtL279nYLEPep5NrIc85ASVyLQQStJzfU132Fv
XHEYOHmggcXG4G1Np7x969kMLlHWmsU9T4Xq3w0DnR1GKKXRcBPIiuRsGTI44hBP
Wwz05qxWFPFGmxquV7xQY4dGlxPtaN3PqA+gpJSxDwvTaUkJtDH1hitl/NvUIQMS
UzaK0583/a1x1Qoc+DcLkhIi9Ok7z6KmPdEiJ3VSUKLo3thjVQm7mHoFRJ3erJML
quxEu55rmcuSN9L9rn0/wEGX/dHNYts/uy4FzwrglUS70sTIXDjq7LhfmUxnmQh8
eVTvCjpDzREf/2GZAK4Ohj7q7NH3JRmgXnfa/9ciWjGfuwiZP7ZU56i1pXcQJ1rI
AS0A3wpUhDR62eZRbhMza9a1doMd4tUP301Yj5ZBQnaPBK9iTskITsRw+fY7PwoX
lxoGhqWzXgOiN9jMmp66YLJAnZTce238mZy8sEjo7H54crUaTTXZ3v+7WoDzT39d
sfJJxbPDz1JvYSxWWf+FT/ttPWi2VfI0clBzIQSEa/vN3VWS/4V2/3CEulCifjkv
rj2jQilPp5LpQ3sDvLz8YmkGX5flSZWLyedcbwJ4nxQebfGv9RyMWt4DGdg9u2cA
+L6KScmqJMziLcD+nYBM6lxjupXRLwdkobx0RgFNY2ipJhxBWmvYhLLfsMOOp7Ha
Hexb4ZjFwhBCpmtRGMSpfdq8zYteozUQHpmamZVildCWPs6UJlsTvzAHlIuVf60n
07oukxuQtPxjajyJLd1OD47Lz7PGeh9Z/C8O7UW45T75pXhfyR0tgHqdyuO/pwfZ
YuXQ755tEJ9CqoUM09xBEf9ITLrEG5mOarbvgkd+ttRLRkPHw7btfL70/jsm7KEZ
rKq10wo5/gbwdBh8w7MPqTvc4NBLaeZjLCSrWNhOlRRG4AKC5JWFEwLNfmg8pGig
/x+ALzRBFCEQZaIWwLN64z5gUVf+Gq5Cyd9sku6wdju5NCY1dlLfHDIzKLr1FH5K
qpR8S19btiG6y9d0PYxayCT54XQYHYpl829ZEkS8QhBSIJYOHNyBYZEWUVweI8uJ
RyUQ/qSI5wYxcga+752wao7htrCQcxFYuH0sp5J5Lw8E9HzKZlcVNFcn9sOGs7Ta
jxZKNQPRQ+136TyaPxP2IeS8Dt95Jahae8pquqEByDhef+s3LV6MIAPGmjNaZHWP
FcvRXln36WU+tnvYMwsUe+lVt84NJmL3pLXIcQN1Wdj8tHucDmOek/OKFBW4vHg0
eR32Uk7DbGSdTs2dkqrdAulKuIEY6OVHPGUbzTev5iF6AovuIYqi3uA/sKXM1103
EupGQljXZVrbWCJAx8qibtkMQrkaZZn5l6v7dxh+IxIFzGjsb+F7X7h3kpwIg0AR
nZIvq1xPCrpC1HXF6XDxHXt+Uf2dQUPTeMUPplqDtGsUH+kc8eV+GV6CyL5mcvxo
DLty//uRIV4EJbXn55SsbJnTKVqja05UrDvuObLRj7uDUkA5AaJletVQsG69q5QL
zgOx0P8+jp5C0fGV8EstPTdG7cJ8lCdvSxC3N8w5BPr8jTrLZ4Q4jK35zrFU8LWA
gaWsgRKytSOWM5GH6WMETzND67vRpsPBhhjNMkXxcmeIJ5olEHSH15Uy2ZO0Qgck
g3/y/oyEcyWaIxaXjmtAi1tXFWkqMaGo+rvNZhdXRKcMpdeG45Wz+tK7SZTd0Gvi
BseIrjwxK9JDP7JI9wIK13NiQi8o9M/tLA2a7VlFmknRYN2QO7Cu6MOQ7sDgEPnC
/JIOqVgTwwyNniINr4CCB7fXXdccUGH/4El31MkFWH8OMyaP4odixJX30Pco8r+W
fqbIWn51Ry2XxDS8SrLI4l/V9Es41l5DCUiIP5SSpLCzTmp0SA6GcbUdLrNNL4Kr
9aKc6n3TE2M2lC+DiZ83mse6ofIhxnhL+hoGThz5rDpzORcVm/427gByJcPTtCsr
fy+8jaRQP0eV+lDqXhYCBinn8ZWcmu9dub8uKrQdVEApR9EGv6QPcmdxfy3lzI9o
+TrnPE0YUe9eGyMLAe+6WCmcCQq7x2eVyOXLxhq0fZ0L0fPJD0bBIC1xzbNd+0Yf
yA1+5S094JI/IZo+BBAFON24pNaq12Z1Xh/cBgkjCT61Rx3V5hTUMkCJQFPJnePt
1sRIvSKsDFjoyLfI0TGTdE+YsA+FqiNt7bNPAQdsHyecMyX2h+taBA2KwzHlvmIQ
eJNFaBi+b3TNgky9X9U508d7uB8EPs4zMMlHwPaRMS8uqsgD9nESjkCA7qiZHSfi
pd4HRPC1XznB7JZ6ivcwhsfQ5GUDcCc7g5J3I2beGpfJtCsrhcjt8GLDzmxLrbZH
k9T/CKkI6/HZZ+zXEY/aCaVssCrh5d6X9xMvQqgRf/GmVDYOLMhC8nQCo2CLXo1d
XhpzOuS/HqCDD1myPCVr/rtVzruMuhA/asZEUG+w0HbTPCd0x2izSlZ0dipRHsBS
OKtmyUFnmgZSri3v9H0+m3XBFX3bif2/FCwtbuMm53MCN3z1m3UGWihYPZjQVJWv
9WYVgW/512Ch2IVnK7tMeNEvtEV3PUQ0qlmsUNOmOaT2FS90VA4liOHQXRL6ZyYV
dM5+K64YS3EZ7o988r87z2WhoUcdrbfY8fn75BZ/Y4me7aKclmPk4yxTpyNX4p/X
Wn8lCJe+i3a8bSN0FgL5awpsEaJcDlq8CntBB/Kzq/jfoIkbrt4/qezVf/bYHIAs
J7BvqTs42Oszx+ys7hiId5144hmQbsc5+tYGInmkowjp8NJsxlrcYdhkkzkh+XZo
r90FTOeK4PcssoYHuKdugneJyKnDtE8TfzdKy74kiFQekoYd5fqr0KBTW0OWjvHY
WHpkHzOGznrxEK2krpaBf9DZxUcAmwnAETGcWrhXe5mbQqvppVgIUckyKrC/0eoK
WMS8zpchvmyLZndmQSRZTphJWQdM4B0QfgD5dXy1iZragw3MoTdpoBwhJkC7HMdH
7PVNd+XPoXdipu8C7KqQ/thIMm9WtQAn9tZjYdc7yRL2+lEPTu949+9iF6hK72xW
X+ruoWxxT8szLfIlqduKpjHgr8y3XSyfUP/d4z5FN5454i9zUXirIbWnon780HO5
V7jXk/AwtZeK7lxryBjBf3Yi6yse2UolMse7OZ7hyGUbpnbfMiD1bze54+VrCFpT
wej7SPwtZl7Cv99UkV0kVEQCPklzo1izk038DrQFCOdy0CrPfpOSXFe30SQ0kZtU
L+tH4jciER2uxqIA6GKNF8ogYO2sqhTTwMvVsJwC11mA2qx/UnQG4zz7M7ahPIV5
F01dk0R82nKzeeKP8nOaE0g6inx2tc83YW7y00PdA1fzOwf20iy7VjyWK5WLxZS2
9rnE09R0uqfiizhQl8h5f9HSXRuUwwWUvAwd6Yj+OfuoXIBJt+rEVELNrrFm3Wuq
dM/isFPbOYXlB2PoYJ4xtaJsuKunDrXwSSxW6nD38yGdsJbkhFLC4N/GYJNJa06T
LmHL4YF06L0SYJRGlSc8CbRQwStiBpwI6t2fz3RT/JbSPbaDbZmkLBPIcKAtEhgI
ruOJo3vij94fGfYLRf40jrmopaEBxyT3I2xLNs3GaXknneASvTZaBKCq/J/vKyXx
2VWnBtyC+VLgm7IJnS+GNuIR5FggFw7FU6UlMdlzf2G5L548rXQYVOIdDDp6NGgc
t8LQu1eiPpKLhUaYpYqwNu7xpl5Yy7CzX8oU7l1GABTIaAezJZ1gEDZiP2ZWK0IQ
5lk23jXbppMEcOhth+dT7CmF6t5CODO2mpW3rkSL8UrxLS0aG5pgyjE9XXqx17lP
4URRcVKXCaam+/9ftFjHa/jjf5O+zFQeXxARDsNoHgWKN92Nob0nrtmTA+Uy1NYJ
leUcU/AqOQna6q3REwe6X4CrJrfaRxhvLVaciBJQoZfg4KfYrbhAJyv14CGxtKQB
B8hwXKf5QM+j98hi78ogxQu2Yj3SQIQvKUxOOMRqP6LghUM+mABpIOXGzOpF1i3m
bsQ2JesGVr5kvHYlDsxNym0lFTuPmuk1rxpf+dZjv5lxh/7mKKOwsstwI49yWrC0
6j3nxHYc7dY7vRqjIWa0L9/t7jmAUvEb/Thft3w2eXYT5HfqMAs5Puf5l7eR2vkQ
5cD7pnsnV+3BpJEHKnDFShkOldgwUS3TeoIBEB/vdLprjkAPZn6mmALQsMXDz+LE
smHL0Zrp2YLQh3XvVAf8HBB4xIKfen4pDw16aU7wpnpgs/Wt3xKJfZAXJtrIviP1
tb+NvArgfcLS0A4vF+mFWR+0g/nRO/NYnFmkb3H38ocpvEPxXleY5O+pLahVk3vm
fQl1DXvXC1I3/efYRyQGvOedefi1GFopL+mZhYqExzeA0GgX+P5KLThRUdQe54S5
hX0DWfmQEEAdinhoqY/cxurYDOKYB/2WJKcD7wo07EiZMjnz+9K6dwuIMuebyT15
mdK9n4BY5lmsTkue9mV7tYWmvKtUbOC+z2TlztA5dN1uLgFlq/dvIm5m6fp86WXK
1CKjHewuLJ9KBfu7foLhZysCSp5oCDEgmsb44d7kyvQQq+bczOZQcaeBKv7WH+2k
GP6Fanq9RxqIK/a3GhQNzyajyU+Qgb1UeG3WpHoVP8xR5Su0rBEIsjsNAuyL88M/
RMYn76WC/esaR18KtlmeQGVf2dDyVyJfKl4BMEeG8Gg/lIaXtikN0aLss44ZHi20
VDxcpxka2m17aoFBbWLDvV5gDzIVRiATBnzQZ9C7npwAS8dyWJTXUWxNwYTYW34k
vYL5YvBAF2n7zg9vZP8agPcG1Imkxu1EgzQdw+YP/m/efXLUr1IWo50oJXjy9OeM
ind+9g1MVhyLQ+JfwofyI3lamsoWYmVqfftE2fJ90icT+L3cSOykY3C2EsuUpPvq
ynkYv/b9XMN9qPuSpnrUNbQptQJmBHVsbP30GHMND9s9DGUc/V8xZWZINM/pItye
CfaICKpH6xsvr419iYWEKjRB+xLd7i2CgF5ut1CPxKYAQNibpsdtYoA5cSDcAkrb
yP5kTaSeRb3ealWz0yMNYkBJod6yNHvJcdx1xNmpvA1xAzynlWGIPyRdLQkjvkYj
FVil8FyOypzFvadR2dqgGsnp+O5Wtlo2Ca3naJ9mZmZhyo9YBa8CBslLJHwslyfx
UxRcviM8DOXgbfTu9CJR0FyxNOZat2bFlQBpjaQJ9/2zA3kQuwalUzJCWoEeqBAy
KqBh7NVOHahh5C7Gvohx7jy8SXQYKBnoeR/c7n5Gl0h7P96+sTB0zRTmWNHI0FXR
/5cGeYbG3tQja2r39XeBiDPFAL9LQOZogqXMgwag5Ud0dIJT/4wMbJxFGrMp1gEw
akBeOQCQFgvmfVwhAmS4zjbb4WHr9FH1Fi0b//8Q1MZtBm5WDowUFuUwRLU9Y7fP
Mkunk6FxQgjIbWht16/xwdgzcgY+JoT7uo5UldFJ4Mc9t17Qnf0Yd2rGsM0C10B+
JWHXsQDsY2RXkHUVw9YZRlevVERZpiqCjbsqCIXI/R14FAMRG5Q6R7iaYrQnUZA5
4HrCnDVp+mVyaVqsdEtAi6Y8LaiqC++/WNTZPFqD3mYZe9aqQafp5hpXVJ+sMAx2
YVMCyyIvSvljKXfPiavZfo4Y9RUlH0Mi5H7WR7gKMPQsgNMVSwgpjkFWfJ88Eokz
Yj91FzRMPetVuqT8HwyKsV+5Tz2yw4Ua2WtXYfLl+ADBDq0ufHo2Krtg1Ke9yj/2
K0xe8LG7TitW3c5AEy7uRz6w3PKwaEnAztx6xWI4O+BJS8VRfcgXuoKIP1ivf1WQ
gqv601mV1nExe3Ze7q7TryzFIIrJ4eMyRJNkYmPqL0+KxcC+qAbgbzd2gI/cYHAi
YCETc47e4+qRqYO3T6kwDty/rTXicYp8OlDm2nCUf6o8xITXplzllw5l3qDxZW1N
MrzZkBz1KXN0kM8XGgN/tXdI8f4zFg9XoOh7ZM3b+6SzFxtXMAdA89ymDbsVjhbf
ywxviSik6YqfeLtXKybiqjGvUOSRVTKUcQXY2U+c3ymzRAKhp74hY+6Gqpa+U1uV
Vo0SXuGVYxsnRVaVMopbEUF+rZ6Z5qi6zhFUo/xdJ3T0kKz+u9KgiTYv5IrUCKvn
za8Zn6GWYRw539vCGpYfmx7oSks2yJtnQ/DrsT1Tv2oLmVmE0yhlHShGk7cj2jfC
ZKxSegxy58WXUmnUIq8vSF7CkeGNUb8K3fVcYE2H01e+HtJvq3JNWcMAx6LJ8V4c
b79B5m35HwDFfGqbej2CCJx6qPyYJGVrGkTJBJneYoPjjSG/258AD/WWHYF/A0aB
eQlD/w7M4chOQiiTS65P9MHiuZ9VDRKPqIwjjkfIZiiRHEYjQbiy9e6+2KGoCLIW
COtPqaY0NkhrlX7T//HtBpjqhCzbW52+vcftvr7CqKLLOy+15PX4cEpcbH9izAw2
Q0yHicQI4GHeMyvqnQItixQajq9/sgQxnCr98+uE3ogHkn3MAAp3nrQVHfqaHxP8
uWWRcxJKv87lE3H9+wg8zBQWiprYfZIka+ur0reoAflc+t8rjYT4KUPlh6CWPyBw
MvkGHJn+MNKy2OzdF1fdRKKoMrRlLxDlYp34TSxVNj2hEThWOGObiqsTmCz/foqm
DY+xg3SB3QoDcWtuVI/TqOTxduzknvnyIvX89cdpoyXwA/KKt7JAkM1fj+TJQwIQ
Gx2hPIy+4OQIHYhlXa8iZOMmX6etSuP8QzbdGK1XMTcb/NhRtby48qFJU9iaS4YN
3t5MXPUCRKfUMtOb9n7ZDfBqfcqhR5gt6hlf156yeqf4b8ctHXpmzBBYKiKnRpoL
c/sTxzs2nGzHkwJM5T0P324lr/PuTQ7eFhOLMlvLcUUgCellAuuRFVGOvn4Wk1/Q
2kF5M3SeJhegdrGjK5pqrxouO2QjlzBaD/N1v5/yOxJUOOF0wO8MeVJ/N1SDATxx
TTPeTufwMJbdd2N/npMxzefFNIJ9acb2P5dEpehhEJeNq3okbYn+tgHpeQvfUbjx
alrHlmYRey7rDihzMFDjU6lVBKTNTeFVd3RcCDlqQ5SAiN0IdTxHndsoEYQUXytl
38f72NSrarf+tosXUOAAi4UV5mAr/HLeHIQcwjuW4NZR04mrvE4Xwm7bWkl6mTMH
p2XI8h1A9xmMxk+qndjg3PfE4GL6N7Kh6rWKNwIY6g+izb0baYAjz7bLBoy/7Qvh
3GEjWUMX2g77qIeypkmJhnSZMsy+IA7yDqBLLXtdbRs2jUGsh8xtiD3go3G6rido
ripMXzCz81hEkYG75fwxKYvWnQUU3AoQiuopmhb+GwVFxxTTXNkwIPId86hMHrho
2kcRhwMMdbHnTWaBXacyK5BURV7vvR2Fy2rwQIPGcsUl1DxZ0rcaLePvzVC/VOs4
Qi0qvgLc//+Uvwh4Q3M/1EE+Hr3YKbFWkhjOASCdJse1ZRm2jPabsUzaxVbxHR85
1wUL7ULF7FDseVeOU0kWejzFMeXC7ti91OntRJvc7ThAimDH6vM2BEJGl3+56m4W
3RzmYRFFMwNcAaGi8eho3m1PhrnB+zNTA9M1soDCfnrTrLFx4Cc+5ZH5KJsEsUCK
OE/AG8Oz7z00F7e0mChvyVHIzOPE7yDasQufQlboGUekdMw5M5QnUUeGqZehaIwI
GBs3/N+oOJSsq5GnnUGUo+YLs7MvBjn616ZllcCcRwsluouff1We05UfYjkjVtg5
w4DdSBzAmQLgRD7pDPRAI/RVfFxdZbGJ37A6fSnAhnmqerldVcNbIaqT8s3WDXcF
V7BIt/9NaPdpkDGPGZl6N1bl5KhR+AvTxGlCNfupI3oQm658prYrVB43849YWLaP
lPoMyzo1XRal0dMWkY465K2RUqWq8LSBCFrgBrEuf1BLao/iG7yXb6J4fwt+txnF
O1mjbJOGIm6kvEL2oWoHUBTHwxhhf33MORJeqjT+0HasThkMEJuis9AsQuSVxnFh
miW6IBk9JD4tbimAgM28rB7zMLbqK31oax0URK2Gk5HksLHLsEBYuomXk7KZaexX
twSy96OEleskiZRBbXz/GoBDXxDtqyfHOecjPWsFqpIqMRkaDScwud7Q+zKX80og
aX47S/eYdi6cguEO0ReCXUjpD4+1IL2+zqSYSm28OsO6ADI8YUilcJkipoHDqNe4
etMErCu0w4j80VAfoIZae5IEpOruxeOkPpmxGDJ+lR1O6err1ODBjf4w6LskGxpg
ZGchLwCpQDUXFEL7VfkASFHQCz6naV47qZW340HIF8MmzERsnJol0H4vZWFeXbSq
jzjbYPcsGJi0Tv/rWYC7UdOvK1VlcziGbwKXJh4eOnrFvSUVuNqe/QAd0cugyVE0
vVDp2W9afVtKOsY30vhb0AG9hG+UHSMBwQ9cm666WUmIoHKrg6E9oaybwtHYHhUb
TQHNs+Nx/6wMb+MUPx5t6k3FsJI1hy91DOrwZHKzMmWzXJrT2RcWsjf7hosIQwFS
42Jl23enJRjzNRf1DSD9WiTu8DvRieOumoE1vVzvg9wd6aCXTMg29gch/Xl1jhSP
zPDJScCn5IB8Om5X+EJ5NYTb0My/vUaiGmc0x2PcCHSPk5Ypawc2RUIndRrnZjoe
4pnPJy7t+ysIHst9MRCP4G5m3Y/HxWHas5ri0sPkVmNp5H/CDbwbWjfS4OoWThSK
O0iVtdeZIjApjBYCkZvO5oVeJ2FToj29b9/bAYLYgJAkMg2/FQjDwZV0j6zvVB0S
Aw9ngg+i2aASgw2OlRwXDrSVVDQ/P51r+eZRvCWOdbpqYdBQmj0X+vxK3JR/uE80
FM2oEtwTXT4rZE/JC4Zu7zqUv77e71Qv87/M8yp3cl7wpROmTvrn9Wve6zAa/LP/
cXPADV5DVur3RpZ1oOSI2/t1lZOdn2uUkX0k6UAuRlXdKKLJSP/6ZZ17mTgFax+4
jjtksCnqIg/lRiw9TSAMBdiFDZLg3hZ+fs9M6wJhUpJ/MJLt5D3GT3c3/ZtAZJA2
AMM2nAEw2nVFyfYGEu7nIdeY2a1omjwAw4Pg4c/7YJ9KPRU0KlPB7W25dmzn5pu8
AeDm4Pcapu7tj/i11BfkJhESWNGfUya7LsNuFywP3D+gXJ+RlP46u4eXnsI441Xo
ByR8KVa8AksqR3+d4V5diFhXJr/yKiDY3+fes3qpYja/QLqpdWt9zrdTs6kutEC8
mkeTA5IINBCLXOg69twD/ZR+TRvCi/2TT913uVGyVkErdDpCJdz2Y3xm+0i/abbS
QrL6fw9z4AJTvtUSiKkv3PTD/IiqvM/69YyrR1RlvU10PcCrgOaW+0X/MKpSDtAa
0JAJzg0HhyvasHFb0NuolTXg3erKsWyWf0Fe5txOwE4G5QwDwCrRltNVtf4FUD2m
NGXnMIkYyPwMLhJAlJlZZtqAiYvu8TXsKlC1Z5HLQv3o2rlB48nPBQsRhL7tsiEc
eQBY7oHARsudOPZ9TLSyCAK6rgryEFtDZbuyllKrGGN3LHF0KGxTMn6d/Ao6HPUM
JmMAsa2fEwO2KeNPYNhRppZ3Ro5YyMC2YNXoj4GZa+bXMJD4y3oMsxEQVqcMYccY
kG0g5vAuuAs7ZDAjI4aqL1hzmh0OhvWxIvun6YECDS8+tIjeXweTr6XDmiAnjtRJ
1LGZgNkX7smNsKCNU3gZtVK8Y+vio0heTFC1xTjQrIrazBqw8o8n0nJ30qKnhJhf
4l0HEaYvfOxnRIhiFpFVXcSkLwSn0aoB2EdrFbACwP5tycGusr8HRH8IL1JQBZ3i
nGdq8oIw6CoT717mbOYj1bRRyEdHGX0EU9R06Xx2ODsr/6b2IyIuBZt+Y8WRnUgv
g3SGgUk8kNN+3jPd73F8+DZd7KqQblndcJ7xPAlKd5veFnFJ3SZZnLspBAVg9wVx
A5AJ9rMFO1UW9g8EXxy6/EKZJxamdojQuVIcOzY7DIULLeFUWPlvUmVAO1I9Omz7
S/CykDBsojLSMEesS3yJydL2Mi6anff5rcmWlWSA+b0JP6Fi/hWfl3woCpygVxkE
+J9O3KuKPetGqarZMXWbViF8BZXHgAlhIvHyDGcbD5IhGEaFOGwGItVWqtBipt1M
QmpPFruvzuqV6zFcjIdQddNGD2pRzxqoLMY+YlVI2hkqnshWPBB31Q8SO8XlD29a
rvanNZArCKR8z/xucPmfjXgHofa9/4kF9UYTDdMazVCGxuwbcd2XjgHKDMEdXhya
/xtyDzfkxtrgA6817ni/hyDEGah3S+gNRRaz9crzdYxHfFsGvZm2Oehq9pYPDLTz
QHi8ON8c/EPzaRMH6aVX2gOV1vVMag+FgzEMNh85EQWh5Fhooo0Rwol4HAjKq7HA
oUK9xzKyTN3Rtug6k8Aj58I+iRoXuKxIRXCOikCa9aStio2JuZ5XPWmm38JCEykq
DSwvabaZ2iUNovXnXzD7iUe8wnBy4d8fQfliU/w8djOooa9j8zMjRhXbbjSdjHPS
KRnap0sKUUShlF0fl5NwuonkTDMxzmb2Llsh9Yg+PDs8Mf9gb2iU1SVIR9Q1Z5+M
oD7M3OjmkrOLdEl+npbN7W5gdj+grUrGupMSII7m6A/WhKTZ1RqxNPFhvtfyPSEY
ptsfeibmg9JgN09z/TWo/I7RUVgRRgxPXkf9QEzq3bk1zPawlE0Nm1FOKM3QoWGH
XgekY5pBC5K2hqn32ZqoWtUBc2YWPVcz/x1HY2WYEZ4i3+MzXRsTyZsEmw/HEDLi
BguxyQUiBf2rUB8UCHXlGEJf1rApix882dzJIEZyD+6/V9TmjOaOgE2w8XMw7rsE
0I4t4Xq+JJO+mrJhyFi89ux8IyIq4Ve5NyptDmJYZOie7unzRXyoNJGKUoxzsQmP
tUPZEea6CKg100mxXD+PTi0FQ8LWNyze+mibSKoG1+8o5TWp2WRW0mOCMqznkO5j
gpyJ572SmqB+Fl8Hcg4pw+vTsMgKiNxHhZOGYQNFOmV98UrSMkIxkBTFR2ld7Pue
dhz22VjWRdLfX1hn1/xoe94yR4tis6E6pZfVBpwBzogRxrvrbCtI3iJ529QW8zoe
6Jp+N7CCGsbSjnFnlX+4+MQwMFskOIGmYFB1THnCECddBTSUcdBFHEMYUhNFnEaU
PRCya2+Edqjwviiaem6BPVy+IQueCyKq0ukJcbmgxOmF3F6bQ5vqv8W9Dbflyw2w
DqNW9VSuPp0Wt4TVEJe3mtoLatU8LXQKxWgXJlOzNXGXDbdvpPUCjy4q/k7sQ64s
0v90O77q06Pe38mVXH80c+G1f46e5prGTztbdN/fcKeEFGSEA9/cxj53BqQjWX0p
ZoPiy2++1maYYO7b2VK+mrFiHD5Qwbev3W47MMmg5GuA1orNKm6jVF8MsnUj9Lg7
29PBEpoHg4CaeJYl+LOQeUlyDLPV3OowiEeA48VWsR0oDuo+gOEi7atc80yLObaO
iV5D4Ua51bDYiiqxCDbJ1Ty58mttfPjaOtn6aZItdVcfn6WJfu+uGitjW01Ui5T8
I5+3Zl54pTzh4aNzujrIZfl+Q5PM4kNcDDM5FsQT6ahVt4PPIw94yj0Fw1S/thSJ
xiZSj+VmUDmlEFK7MOMawxkuHEBWia28l8fk+TitR0TADQigPX7fNhU988IZaSz2
1NCEND3ukVxztEJDFoqhEf3hNuiqQalN1LnwZHwhTFLKkZNbXPmrzmRcVFI/7jBW
zF8DscjuMK0JhFZKhceiT1IZeOI9dSrvD1tJDSjei3DwUaaMS3xEnQAbHK6FiuPL
e6Va0YyTdZFrPFBTIf0ZxwKQiVmukAPj0l4q+lJ84GAUKZyJmdYHQ0eiJe2fuLea
D0IRdNhbBg5pkJ8iofoh4O1Uf423xgNV4f2F4vdn0hfQ+0QVqzRiMhSpzgCgTOZj
0UqMXJ2fhEX/VcwokVN9yYTApYLIFO++mPXyMJgR0PU1UKmx70/zFpWUed99y6t+
b8TqhxinOreg8HCnfqjzFBPV4nJc/RNH5XTLhknMsBNjUq5FgmNkN84fad0nUD8G
yrm4MaKh8rab5jjjlXoWcgWJZeRPp+v52MHnsj2jzrcQAUb6xLoVzPEt8aQ07ds3
biK4NfFcCZDuSHKr5g3w6vExIFUFHpeXoJ7JWSkXWztzPMQ/MFDjEURkkk/xqeBS
G0mR3IuepO1d9QxEBWq/Pr68sG3FT3q0YW+ghDQiJvWIubsMgtelNWB1sMsjn72M
r9Dj/Kf969FHpLTrJg4QpwHobZ4GP/7dwKwMkZgTFOzL4IRq7yS3zxBilcGJ3SgM
0o8OLXVllz2bsXrscig5C/IBlEjp3LlyliQ6SuNALDV/E9hxlI+NAFjGdme1O+x4
EGc2oijFVB05G6LHgqK0jJRfwY+nfiUCzajY2oVC/ZNjvm1W3k89RYFzUgJWKZVi
JaKpFSqx5+fCZsWuwgw14bThGXBLWIGdl3L8DGd5buFi083FgCVs3ElZ1AI4nCnG
Q9Qco+3ajFfQ4Ah1xPeV5NWomPkTUQr6szd102TAQLFCZXNZpMgyorvdSxTNggez
GApZosrL9ENCvw6cwsKVSeb1Ybsca12KN9BUHGMFRZOO8AsxPAI3fLeixWTTUDrO
cSAsoqJX1XHJt+TVol7eYNeGslcCMYNsNzNagS/n1cGgdzuz/9IwE19E+noBww6z
lsnOuBAxgFvLRi/Fh+Vhn3PS2qU7qpqBIWY2m/0k++q1pgFwVcm63hQZXM+kyh/g
8sSBlk4anTQXKNoeiFdPbwff0dmS7WPiXhf1JkPZfYU+0xsJ3xxRceYxJFkSSUcQ
g0nekn8sZoUQ1h4Ucsu9q2diQ8nCqEar6wgNoQMxOeqWIzM45QRcpAdMgrVf6/Rq
tfWRcIJsKkyIX1uyLCxHeX8M2juDUUm7D9HGWMYISmxmyJ84zs98jyZtwLRgXQ1L
wZoCyxcJtRS7pQMhQNDFhFDI54mkpmsbKFb4ZPK8Et51IJWw+lJx5PooCb+kSZOc
77u34ZbDunfnuJcSvKbeYT3MVhMUtX8cCTgzH9s6o3Hsm/3Y1oi/of1fXhKT++Pa
gj/2fTsHIwiD7WjahWsnNpefc/u5acM6leY3KmqXIkPFGLAldcsuW/P1R11kmIsw
iL068VwTit3HhP0r44+Xxh3PAOSZQiHohgRiXOsNoZpE2U+pf1/7NmLH4emsBHl2
tda8NjpH63kYPkFSju17BD76WcxBrzKg8FjUjQ6HSUI76Whu3JmGv2lbI3uP70yE
NNC+3Gg2B9akr/6DLz1LlfE2vZ9HyRAQZPBL/GiC5Yzm/NLqc11xjNiBadDMWXt/
paGi3HJAu9jE2R8CTWEP3jwJo9wBo4ubJIIlXwHRO/5h+DTftWeDVsiHWiayr4dg
YQkWOemXSGAb+OVwXrpqmSM0ydw5Ez+k/Up+HegGar3o4LGE/UbMZ8kbxLMah/sb
WEeAVktYQXU/eauBarnEjWq0+mNr1ZqmacFUcE/IDMx1iDM2YdOlLAk9GlVfWi9K
bXVTVGLxlucRzecE/nbCteqoKUfj7nPhTJA8J82P66vsqn1+LhbbztxJVpqya1rz
GxBGkhWy3/g0zlgL1em8ImJmVB24zMaEiwWD5qGABK3UiElWDG8RRY3VwAw2egvi
X8PH7yJLDGu/+RvgtRAftNGpxhNb5MlI+0WSo+Ck/BvTFliGfqweLoaShHEs6MLY
cLgCuQWmBCQLCLAQiv+To1oJbRMlPX2bYjHr+yg23SfJJQjRjfGVzuHApWWmBUE+
Ziv4b4sYzSC+L7C5ZOkxt8OywZKoxxr4PDqJMaJAqQWUr43C1KmLovyTQLOpxzZ3
f/qVpx2R70kWKkYwyltRb0DbrUYjP8NuFfo0ByAikiG7YM3OMIBrZpemSQW9Ij5P
hUflkFuljE303K5qiM2YKIVov6R9r8a6a/V8loxe3lNaQJTPFQ1EYmqObjJyEnsM
QpWqNF5JYKC9BzBzSTVYBPdst8rU2aN3lW0B1a4coqgc4datZpMnQeCX17luMLD9
N9FGmK3ZiiB+HWrlwCqMIuht7vJPgUeCM+wcOO7LOGqBE0DWlI4t2/42MMW4dtuL
hDejX9dv+kpn8rz/eAsnLHsCE931+3I+wtmBRj+beeOxwpIjPYvlSmR0G3Xdofq1
Mls5OoFF6H3ePKb+j5OauXc28sKM62Pq/6BnjtJ5AdFljt45FGSz0kgUGQlnWTCi
ybOnhd7vB2O01TTITHh2N6HDfFh9N/dtvuPX0s6dmKo/mTIkdNMZtnSDQv7BLOeB
E2C5t/5xhVvc082whcvtllt1zzKJinzry0j3fEi0IujYVHnGuxhycLzrueUtleVx
LlJ4KeNmJfvd8Waaony/Pg2NMRlbSlkGdGbyUn4ZhK/xydqEnVkIaQxRdr/3ViZT
O6C1rCqKEVEmYP0yMngZBv8yUGmH2YvCny+qgerXhqjzVisr8AfHT/fwDA5KkVK0
fbbOYvFGRtWl+am4n91pba1WYAKpunefHG59DK3JmdZGdEInM4Wj4FHosU6Jp/vN
WV14Oqd2lHvFD8HxdFzTmxv3cQAU6FE4bcLShk8O7x5D1L79Dv0UmY4WBQfeynTh
xD+yhG28vMvwv4hp1JWOcULjQyH46gsR1vfzeUzMixsRHBnvAo2kvYfOtIclgk9p
QiihEC4vMYUvMxvM2hyakoXr6ZTM++w44UfrKRhU1t4gqzmrGT4/lvRq0aRQ1mQ1
dnNHrS4DBZBGuJ6mojh8XXT13W6Yi+bIbsDbTa7r43q8nQM0lKf5qIXS7HPi20+T
Nj7UGVySGtPToLGCtGeyJZXWXoQT/26U8vZIA5FLSzufRlZMzi25UA43vBDDx2QJ
HIEXbpbIqNAE2m0+DQURR7nfU2px23ijTD4utV+Q9+lKTP0tYRPfjUY6XW4+pOqY
ewn8AX4ghw/0eapozttYcylj/Degu/chfH8pdsFTStDmr8k7uW73z+Huupns2mH9
l5XwRQl+Soc9TAB6zbkSPWWmlGl438jR8YYz9Z3d7x8XhxhyiVshYFZEKkx+eWL7
xp3aAuORdKT9d7gptH0HdWchub16x1nMT8WVpzjJEkIAlVEPxiOjMaFQdgmYC+3S
U49gZancd5kYcOxwQQPeiW0h52tSbNcSrWdBYYsfl6C/kgbmwMfOZ1+wIL53bWeb
rBrG3LcgXH4jyQS97C6tS7ATpdEH7AmMMd+OpVyoqaqJe8QWuSdc4ZSphsfCyeuV
AlQ2uoBTFbNHe8fe6gUwKMB7EegBMZtCjMdcQ1ag4ioJArV7OXwZwQx2s7pMqbKB
5xXD+vMQYOMbaHYnFPSrLPJEfyx24e7ZGLz5mDSW3gakiZbD+KGGaDM9FOD+jWdr
3cLjUaakdavN+bRoZsfbvm+UOfMK0xYGHKjEyXaGvmq0taxmc7+kntL7QCytZpIm
pHhp8t3X6nGw5QrGswLOTw7C1hGVXU/ARZ6Sw/QoPK3Apqsu9sKY1cD6bCrUE65C
76vsAsiaEdEATmJnBXJRfuw8EmnMWGsNoir36vk9o2AQq+bpUOSiDffrH0Sxq/Bv
OFDGB9nYsAXSnIptIklt7Em1LEwiNC7Y0L53RLfRlV/gb9UfpGTMT9wrQPsbNExr
xz3gQqJt2fStx+fZW8fWEahYEl+sP9M+G4pOURVBskpZHc5LY2XpHdIpIaQkI4Sz
CEFMuUXlcT2Zd4ih76UwOWPJCZGfNP9zA0eyGTapD7owwyDpUAGaJHoW4n27hzb2
s+FKJwqSjwXC1N61TuaQEEkO1Kp4GdNWbw8hukry8w/A38XNLtt9GR9EVw4V3iET
3dhzzNsfA9bHqn+w3D/bvAZ6PYLKFhWN42r4TIusfTfRS0UeCTB7lEORHNKps1ab
x83Oa/AsB1QqZ/O2MT+BDDGqDUrFHPO19ENIPkHaJ/Fuw5lr2D/z1RAh9Qn+UiD3
25HA8fkmkvfyA/jryIBRe3I3rhD9o2AKjjj4ZXHN9mhTFXvJ0prIyJ4TdORi739i
KzjKRfczD3tZCUPIQfXlyhQZ1mS3pk+8ohRAB1F2/KaXis5Kjf9U30VCst8WuYzc
7HlnZkAAerru8j2KZoyoqfeGt16OFDFbtjWwRairpQejNn6mKZZY1AmSyGLLGwc2
v865lPrmu2a+pWZYP9WZzgO2n6Mlg8ugvoGfTseAOr61Wq7khmgt9ybtCFNfjMkw
XcBQy3MkO19TnpUDMRkpx2hf6MaVrjw2aVfj+Mnoa8bRzS4QqmZyb7l3jLSpMWpb
a1ju01yPCF8lPk3NqaMe9VXi1NnZuj8UfMu26DddNjN+dOkgBfub9Ks1CD/TYOKC
DTykaTWFrnv+MvspHWYw0Y4ETgPAHoVS/92z+95t2bcWIEdw83A9jZ5jX7hJFAxh
M0obK9mSJrWtMYwX8Hwpo6IJGZ1cvp583AAvnAzNXpJPrqWUojiDaqsr1qZAsv3k
D5wV+1kuDZ/FszvXJwmlalixkZ8J95XTT9m/z+Cdmd4+V0JJYnbf87ZYOPTsBFe/
HnnHLEUw4qRC9NgKdzybgvkn1ZdlgT2L4MhqYPZxsguqyelLqAP2aLmaYa4vdJJS
WMSYo+Fr7Z0hJeevCVRqQ7KeDdaAjDqltlmyXcTJZ7hlbicCVWGXT3KNY3OUdd3l
B+9kyeK59ygmBa/tJff9or5YLNXlPdB0WW3miQd49hw9hVoue0Jgea6sUU4zSgQf
8zi2q2rnqYFFtdK/vT6cSIDdIpY2d2WZenz1fDflQ3kkPNc6sRWJQjB/jwOjyXYj
G9vwqJXBIqv87wWNfxYcH01crqmw/J/QQGzsxC6WF2SbX9qr2NqKQl8M5KY4zMP1
sp0l5V8ykufUF9/XEC0AqMDGvuiyQAf/Aq5dktQCa2PoazSXwrhwbm8Oj3GbI9yM
X66ofajE9VSbTLpMpORXsXhX4Ejh2isNIhrz6DbyTZC+CB8K0pKeE+XBtDPJcVuF
1Gsuv3nxMbQxw46tejA+1uGARrH46FKvSBmiXq7Spsca8lU+7RUY1Lid3MkURu3i
adipdpjcrTv8u8Z0IUisrRQv89f4MXW3OENQlrvMejznMRlBSInuTgNxJn7gX8a2
H7vn0LCV+GrkiUray3gjRRJQlBWJaaAVOZKuLkdg9YvjWczMb+Qof3A7n7mlmmAS
+KyMenhF811vpMDDMpz/kQF3gUhBk2R4imuXkYd0/o9DpsxHWSEaLaSdiQltstTc
19nt1xEbZRW3GmOttaSZrbKds0gGrZZqLTu8qhnGZ/qmAz/EEGLkTBNTbC3NfGTj
Fv/PMFTTDow25yXI5iWItve0c+6QltV3i/2E+IEtTHjQ1Xe5sSWN+xzKEvTnlX5A
KZCSZHhLJRROL2f45SQUE59qTurWbEiTscfn1xpCdTifTCECy+7oBsJi/YJI9lml
zuGEQu1UbK0Hsf07W38MJw2f3gb02512n7xFtB0phg61Ks+Sym82vjFq58e6GFaZ
d6Nzz1gtzwniHPp9BBUw/tMpdJedNEmqF9T/NP4u7MSlIn0mX0QOPpAWQTrEGT/4
JhQ0cR9mZkC0LZb6Y72Ez9g7DYgeaBFcMkWB8mZUkMGARvPqa9jj/Gg4zbAYMMtD
xCZOLaJHt8eBx3KbuGcZj6xK0uB3NebVozKdAXmMDNuJUuCSVVd9EVtDUef3jYgh
FZDpZl7+rydHdZJZNAVEpxokVYgSVK5Xt8I/GIUWpapSAJ0e3Hn4nIoipNrScszE
OibXZIqbtcqyogfE5tIsYhypsZkGj1mxL7G45GJbgHi/q9NYgupvVjV1p10LpVgm
+F7HNGKx3ouHbBkDeKGasKaRoC72od9cLehoKeRA5aZJ32ZIyonLdD5suV+uxmOc
Ac7AqM6JorAXbDnP7+KR4k3TxZnpIO59EhmuGsHpi+a3fFAlOTXkCM+iU9gelMJP
TlAS+RkN25AjnRILg4QCQ+wbZksMIlahd8VY1Ze3an8/dvehQcC/T9xp6NNRldmI
Arltw8QpgFOSQUpiUrXAB2J0rA3XAH0Kn62pMlNabaOb8Evwd+l5VsgAKG9xc0Ek
E4rn5lxOAULEV7M+PThty6KCfvvxJtTaznJkleMRMdtvFr3mOCgTcw7PEbFppGoY
tSjoSMB11WGBqucYicjT9s08lWl2+3WX/A1ijOmmIafhsP0eaNaspkS3iMzrSEMZ
F9fuaSHzM6cVzdoF/oNRYYmUtwEE1NTZP/UF5zIy7wWSqUo6ZZ8b/mX6EyfNTEHG
IveDDROg7SKiWbMv/cbdH6WLKMiWQu9LA2QjAbsshlf0ECIbjJz1qGtMTGRAtEgY
rHp6ioMye38ttiOE6t8HKDv2tnflkjX0XQvVdmC0mM+UE2H8wdA9E4C8EvbFGtaY
O+ZtUiINvNDw5wa6+ovyaCzwgz49neIf7JXMt7KgM2hUgdpOlcAty60h2ov+VwP0
ZUW+ET7PcnFIqDFJW4MlDp6Af8N/swijUmK7dotJ1xvOndh2FPN8G/bmpasAU0+d
HwrAN/eIpY7ts+wkUcQcMwy3qcyWmFLOqd3/wbJiqvl/4fVtvknkdmNWWd1LwMy9
5fm57Au56PLUlqoDGF9ZQQIwKscS0jrI0IBStRPirDJSfyxebnJ9wvYwyxMErD0m
61tCz/3g7UzOc918z0sFFbsjOZQACSL/uEE9FoJCOVmrMd3v3g8J5azz0OTkNDKX
/UmnEWxfFRtC0swOkK3+ji5iF7u/retMLfBitkIEIbQVjYkka2jru2eQ9F9ZTYXZ
J/GnTtsPdAxTk5NYA2TJOC8NWPpQI8SotqCVmNH2Gl8DyNsmhMPmBYCQx+PIE7NK
X/r3UOWsxmnN+nC/lMk1vZLeexgOCvJDgGAS0Wk5kI3N4Y7AlrwFrPtvsUVr3NmV
16Ble9Uo+8lc3Vy3aG5Iz8K0nvi/Pc1ELcv+tuz1wTW4Ge422TacP52VUUQaG3N3
Opb+pNRzoITClIJGaGSSl4LU4HEJRVCvd0vEe2aT3zv7SUUoAovN8DPQyLz43TwI
kJ+j1t/sn7pTNtPT6ASh+sjnm3MRgAoawZwoLMo5I6qS+RSqjpFSoUmUjIV9qmyz
D+fV9/EKTU3gQv6nEbMJ3/L5jbgAcy1Rb06+vtaqEkEnwnV/XsuyUfYB5hgX7Ik0
4r9IJEquq9hB18fUYfD4wTg+nL+f8OaPDiA0mVza7Jpcqpc1gRahis8/KVVohCGV
the4QSyyKAfRj0kk/bz9O/LEc6XT80G/UfIC1LRrZz4EMbC4E1DLECgDQ+Oi52GC
BMvGs5pSrFzVolXy591P58XAZFe6sN9iXhJ/4mWu00ZeSqgcEh38/as60DKt+H9h
yNJ9Teryr959oq3A24ut8IYhQhbpGWIpf+X252whV8/q/32OPGTy2LetPStx2VmV
oypzuHyyWcZmfXVIYMke4yoiBb0gK3/ovNboj8acIYdk3x0XiTryUO2p0MeGM4eC
QUmHUQLbM3WJieKkPJkbsGY4+Xt7nSq9Ei8o2WF9PEWj40jZ7yuVheKeoaJ0ZaR6
EwVqQ/ZkR7uESR5Sp7ShQCiflK/rR0kR3iiJm1TGoxYMUNAaJoqKHR8pGIU28ccG
PMFu81sTY/yn7kQmA6qN9FimYFg6Rmr1sfDsl2IAwhwZaCcDEhwVZqGrKLueysAQ
m4HxJVxZFhpOyxwO/t1xdl0Ouzeypt+6kgGMXqLWu3Rxty9ZJnQPnPkCIGWebggH
kq4iAt7NPodZGwt/qN7xIwNkWQBSsC0vDiZzlo5PHZkGNmuIXnZRekK8cesaecXx
W5QD8u0FpCkzLSuvpXXhaJFQjOWzViXj66MWrZi9uwOAvGILTKaRrtIX97ee/j/M
VryCFi/e//czQBK5N0wlZgfJIZIWc8955e60qNkDPTef0oTv5dKvqiJqQJhUHRTD
+i6RJVYdS4lyPbzv3amyFdZHafHvdwHBL7LOkZfv3xxi+Mw+HUAA8vSqjU8ri5Yi
4BfjvzEuvmYcCvNOvMPydcShWwu2t84srr4rCQBarHnvi+GJeI5ZQ97K2YzMjK+i
2ytkcc7qUJasC4djRr33FeTnDblaKsNe/6sZpyGPAzk6uCo9S7UvV3vrgElID7mg
/xN9sHof85k04SjxX4nZlmwvlmal17PSi4rmORuW1PiGD4cwDRAKWHXdB+q93Bw0
f6V0tmPpamR8sI5PMN0s63BJSfZDLqJisxGrhXhrKNAnZW4t80v2PdbaO7Glw+wH
XzjhOD0Sn/YPraC50whjltZLMr9Z60hZZtywHBDfVBUMia3PJa5BmvPWC4XydAsV
ILIzJNRnBiqz53UKi/YET0tC432g8zpLAvcsAAdbQTXBtBjgBOOPqq+CNPk2tpBr
KDpTfFv13BqPlf0qXH9NcO/nL1J9favrAPGPOP8bUSJXj714rO+W6xgpqBDOYGCo
wFIUso+AweVNiqqVVLnTwOQSNG0929nRelnESFzI+BpFbbOJX2LL/kUrRIk+UwBY
cTAoPCZNbJGDLqnkxCL9ikz9tRfxCK7xgvT742idZ0nKGjj5pxEzR4twoIJg7JsZ
me2Ik6hmMdie7XdNHy640SycvP7stLfWTlwpdT4DdyAr6Na/xgBtbrK9p29t5XDO
3HjUEJPhRKqSdvdbzdXuAj4pK+71Lf7IBDXk5CfraP6A5QzrZkgJmjK0EGqfWxOh
2/w2zxWmSt0BRwLvgJp6AZ1+aXRidpt4fWg7Ed33448C5dzjRZCTianXDLjzXa2O
ZH11BYUMmug38hO/pLH8mlHxs/3m38gXYcvZuYWpgxLwBrYlbEZNrGQwXerhJkGJ
HA6U+YLtl88qVGI7ifmKeFUow0HgWC/5bhTpJDZlwMUc5NXfLrKWBLGDEAvrK7Nx
gBYT65t8/0bqdonpDZyCbUGOqJ2lhLgUGIUYOBgx57iGYLH95MTfVBc1IiUb0/sJ
f588bDgf26b06c9P4W2/zY0qUz7bXKpKDL8dBUfpsl7LU5/nSP06gjvOIxF9nWvo
c+1hx4jcj4V+f42/uW54EyzVwqMRcpRVozl1h510Jyb49y7LmmiZ3Fjb5axkFlGY
eKPoSluGKQEF6f6KH3QC9X4RKunNAocT5r9/buwjvdjRCciRfvhgi38avfOsPb0A
o7lsTqbqHnd1PJ2sRrtdGsu3tlIrkjVZHW/bQnZVVvGx20ddqNCcb+KxJBN21/eR
d5kKcbs5Hl58n6aOnBAEaUar69tmqSHjEGKbta5chf6qfMgdTuCN5/Mtdy+gAwEz
6wH5wlq5y3xQsMdTUblHMJtYVjmZopmv3eTh9GyOSQZYUj9gQx1FC8QrJmUOVFf1
HueXZrR9ytP5H3CKPodckrRzxa18v55/UHrZfPxAz/sUjb4W85GLjd8n7YTepJQQ
RDF1JbvupYgUKCZqi9cjAgDZGWTsgX7Yv6rog50Z7qfPFpeA9Xjg6o+3j1Zfluds
VPaGpDnjUwrMZgzMPLQ4xaQQLqnf/kB+2wWK5ZdvQi1zlrym9CII5GL39GeVumd6
clpSIkI+3ECGfKGJCGQZLmxhCDmLBc3e7lwQuTAwpKAZeN7vaSFHI5lNDJYZHSN8
sFFBIdc4dbU3N5qkAzPPn4op368/2A+RNzcceXJjaVeaw0QMdzuUQYOiiNVcBWP6
6M0i7dtQdpbL6zK7ElxPDQz1akJDS3338EuxspzaMLTwJ3wM0jAtz2F9H1AaRs9U
GDgtkkKJtnonCWiKr5FGvsh/RZN/krJ+MlwXAg6N1weZq6yR3fJSB5cswmhsI8VK
h6hgXt/QfW6HhiDFr1aSgGWGXqid89ThG8tBjOuCA1Z3xlupNOtd+biEE6/O/ldo
xNTPO/OHUVYPTOg7ChE6XYxJ+7nYB90vT28UBZNIiaCWJGcceJiCJZmvb30nJQW4
dYFFfwtO7kO8aa6JQlUtsWNZixtFJ1H3KBlDrI8gcK9b3P6aYp2CfeJWeuipgRh1
JVp3WuYrbsVW7dDG82jQ/FPnV9yoXYQP66jcH+pve/HDTBMSzPg+A1f5KAz4lOdj
X51ellQXzfP2oUHwrqzVYwYx/z4Tv24yLBU9Di92PwcCSYEmx2KC2B48C36EtUFZ
KTCN4SAmtOK1iy4cXtMKEciSfXE7I0cTN8g/j1fwdPOIhR7/nKb2Pf5fgzczvTYK
n9sR/3Oloz3MMHMDYL0Do08GmfbZcS+nxdV13j7H2sJ13KZP0sAjdABQhUtdOfnN
X5kZS+5wD0eBNCbaIEchHvtR+L8WPS0k2GF1JzAQX/q6mgycE3aWh50FtMmGZ5sO
w5Irx0GDGgJQcxsNBYE3/XNjSQKJDMVU8DdgD250ljRhS5a2E2paP0tw7vUzQzA/
/dOa84BWIr3VX5gcACKFbkBu9PkqQfde9dI8uQHyykdM64rBTgkW08ixx6Ohu5CN
YprgepDB4xIEyPT8bwQguOt9GMimfMNUDI8wjcmSlmIaCHNL9DChT8LBbYlDYpkF
o7JwiHz5kqSHV0SeOuv+F/U0ltZUUlQbXv1+FepzzV+dQmLyp+7RUKE3pQsJya/L
s9dMluetYwhBjcieZBwnXpvvgHNpmC4VeMRNHpxjvX7UyoUEFaetgPmPCacrkHYv
xj5ZYUlCsggpxa22N0lHzfGdEKzUYGA2psw2lkUKW36k/ypFXj3b0TzLRaKcq0li
nHZTuXnq4qtiEZezsxcseFV/q1t/2NfE5Hi2YKN/clpcI0QPJGVKLgPv7ZIP3DqD
iIyTwwyAAJPuzAp45PQMnDFCluk4oJK5rr0ht+AiIIwXEKhqXkNBzgE7Brkq5/hd
QuLQuwrbK1LgVfi0PK74Yq6r5rZ7zkKTjjDv1XwswUJ4Eay6pBVZDZYE/MzIDkL/
T+8vjt4DXJ8CnTZ6WZ9hDvN4jiKK7CzDmEXfMgC83xuh3GH/ilghn3ck+IF0mYUW
vQE3DdTfbrPQJSS9Yk966bve+uydO0vlaSI46bHIYTr6BIEo4ujMP6seCK354Hl0
wso5uPVEEOCC+0j0LQjSFYPrbGTU/1cHGB4o5aeMdYMIrS14/bucnRawpi9Cytpz
cRwKvk1vzfu5Iy1yPJRMZYGkpAUC23Wv77fVK2rh/BP+0qEbMsi133rIwLmsRhRw
QHMgEXA5w1hNvjlCzqkE4qG9Jks2J39BL6jrh1CQW99Orw0/0w/rt79+fyFBrnHh
oTseqqmcxiHcNpcFKkLMFPrN8O4lxz2eCP+vjYzpV6ovRJK1VwqL0MaVpQQWFpZO
RiT3+HlvTtIrPOPdIyZqjIisBczxg6AN4irsWvMyzFtqnEYHs3RsBR53Y757JB15
Z8uQ9FPlXHpHfkjrWTELNP3htc5Vx8D7fwt25hLcn7kMfgzG2lguB2FgsOrkziQy
aO833QKnIW202AiBLrVVImcb/JfIi5jdlC4HK2nsZOpoVN482TEEYk6hqDJqkQ4Z
nyRCh/kqT4BeQx7B4OtT2vvm7YybXbdbtHWNLhkbiGRqjeK3rKvo3raBd9Fs+a/L
XYksRr6T4V8UO7b4RbTc26pIfDv4F4g2e1ZNV4wXphdK8miCHCJMUzYjnrr5s0SW
gPrKeUB1pY+yqN/8yM2GIJJQQwQ+oQEfmMKbD8Sz1FstXCokWgczOHqoIBEVN3nh
6KrVHikItqfu+wmDy/HATKS2Pm8X82uSDIdLjsTX/+hFBp1jRFY5c/A0krqfmMZL
IW5T7CSKPeMkHp5I7kGoTu+/gOhjj8RGGjEZYHB00Y3UCLLUlTthC5USr5vKtcNl
jov8RSElmqfhUpjzIBWScCIXD+TqIuJn0+BFM+6uiQzmGfkf336Sqioctsr5lSt5
pRG6/68MWMMFB3PWy2O7Ojv+9FtrcZi4Gp14ZY++Z/DDKoT7Zch/WpAQU3+Zx+4q
YwjxbWylGNNOSgbJe2KK+zVhFcER63cWB8b0NkAvd/YilYl79RDf+V0tluPlcVCQ
zwWdu/NJ5R2k8OSEQlemKK80GocbkZtZ8gs8PHv6AVErq7gu1D7zQyjB7QRiwIRd
C088qJYPbgFVfjdc2iqonxVb3BC1zXHezsPGUnBi3UngBmLZU2tAgEu7puthx6mh
xTYYfkpqe7lPsP7oolCXiaBkLGppGaZtq13q7Agaop3N5DSHxFWzlJcZCwVn/Cmn
hO2VMr9TEcKQKNhmXpvAJWQi4Nnu4vVK4K8ztSLCbfbdZIGHtwtdg2+CjAeTXlkJ
NGdkJadBedoN33EF0Np2cMRZGwLsxPwytgeVg3nmGadILjvWjwkJu63TpkaaYx01
jBbdjlvvC+03vYM2r1HFVh9F4GUl+uL0GEXMiKl7cZOPRrC0S36ddbT1GNu+gC6V
EklIcHzr7xIz+HXR2p01YkcTEi7SpOssTRWcR6e/cYWHMz9lWaE7iiM1QHyhRDfq
RgZIFpgUBZbB122aRGbiZ9313S0TTy6xHOje5Mnw9ooGPWHURyTcLTwI34NUMWIg
990+scfnZnO0DT9bD4syaoPG9VqlPk+yjAn76pUd27cAdglYLnE/a4brak8s1Hqm
EZ4iAPjuq+rrlcW7bFmZUtHc5lcCJYkJz6w87Gw6UQ6AHei4UlZHO0Bm1Tds7ePN
9gyyJXXxtUQ9NW43OWNXmk+aiLigqk97//QMSqs/qhgDnXz75TqthIh1n8RnvVOF
GJscORqNqHxJIgnNg3O7JTXAK9QPu6ZypFtNvLJ0N2T23/pQ+RbHw+ZAxc0HiQcZ
3mYVyt0sZ4yb66GYf6LLAbA17F3PdP4p7kVPQXQAHACLI1xO3JytgcQxXe5QCwu0
ExCGGbrViGt+meoEbr/uFIaThKjx9x2VUUt+dsMBBNMdesWqUEkEhIwrQvu36H7L
rem+lJuRxIvgY8SdByQpv4IOZ69brDygO0GU3Xr9UMfOy5tusHR9ZvPjBNKxYa8b
UE+WvzGrmPhdfoVEuKhUuawSVvAkIljMcAtXp/lOJt0And74Cx621O9ptmceIkKa
2exGNp5e0qzF2bVyCleVL3jeJj3QKn51IUjcbG5zijil9dbFyfYQecWiWc4ojrdy
qnFNg1agvRkFMZG3p+WKUatQ4zK5XB/ZbxOYnV3QpocrrRWCUnPxTl+/wv6D1dRC
mUMXZxCk+9VeWrIybZw4k43r9I9S9C0zng2AVStO6Ig326oVZedBOGwEcjz5zbP4
/5G3K40a7OmYZ8LZacsIKDi/DzbnTXJ2OVWMSHvfXIg+vyYXQRF6ECk//+PcWURZ
3LIhCqnlwKlCGzEhcdxUPuc1bXW7JlcpE4ZrchNBC7cC9CC2lB8h70oWNCYmES6T
JzHlK1VlgMHQJnTQL4juqN0a73NKnotzGw9GsthQplfklUTfOCC4WIV0oeCPMwgS
GifbthqlDGsn3t1ecJmNAQyfxYBF0FP/2ctE49bs53XIIJpPcBp93sn+iE66nbGn
0XqsHLhkZxDRObXOQHEDQp/Qc3TWbQ4qyVjOGtI5pW1buTnHT3tryjZPzWddpSHr
Bsv+ZyGrZ8DlVIF7tyT9TchQOWsW6wYuR9qS3a24Nu7w2usrfrKb9yiBOnr5D6x+
Rf4Hp5EHQjyUAzyc9vKguuAg2w+HzafjOvkUXboifPkJLp8wKN15gUpjYQvCCsA4
ShNmeZJFlBmqR1/llR7ewBoqZc9pjIh2vCK2pwWshEpBrg20pPODHTHpxtsiC1Rs
OUpMJx0Xn+bLrxaxcoxQBBqVmc5GgAomH120RP0gCaukt3C3lPyr3AXOlJpkyfex
E+E91JSS1ZoPRXVfivXL8Q83+hLL5yorD2MxHjFZGJ0YO1U4OUzmDmOq7rUbUcLz
vyHNr9W3raWko8h2ITiM+OJ8Ziwyl75xMhLLEGtnUeo06lnagOI2NUErU7juVE7X
JtfgXSCWhkqiGmbKFkeOuzCpyEldO2HS6Yh8NNyTgjRaiV5BtbKDGkddjeawDklt
LlaRxGU5QKUCVp0UNeyGrpIhlUbeuOiButUakKzNTEmzyKzexI7gffSrnqj4uhd5
hSOcR6ogydhzEIRvUFUAU4Um9Ql6hYM8WeP6QSW9Bd2HQFum66L6z45omKJPsMR8
y2Fb7Xswblw4N6ZnJhf1detEPXvz3MtaVOjhcqhTFatK47TL3RGvVrjSOKGtZKRm
0Ef09maK7WOtqFO6DYxK+EgxdnG0WWzgZMlcbfLVo3FLsc6CQlDeiBjPJuZfnSGd
5BQckup8ZAqf+vEE1K81f/PnUNHhugVmoYAPPmyWysveNHXjfHw+EXdxI1UPhsgS
+rT2x93+TeqFAKMHV0rDQIzNterpooofIZzEIvWDI5CLqSOtubAQ7kS+GkswCPqq
kcu8gOlJyaDYYKDJ1cSFnEjDe1jtKLLaVP/1vK5FenemNH2Jmy/7TR2dih4dGzwR
oKHRFhZ2HKhR0abmtz3yKJlNKHE7N6LFCH5/i563e8K/BbqO+9EzIQSaDsFVdGeD
46qoo7lhrgcIeLNogPIUBzijDYmTyPx2AVAbSQAqKOEdUY1qY8SAuX+d0bC0JSPP
jlVl3BODciJDtyKAjka25ziYYRoj8diyuY1iIoYtO+QtZ7N5lgM+XR/EWRbl2+4b
bbLee/p0kx2TXyXXPrJ76KMWL1TBe9DhJwnp9I7Rts4ZyTSKx3fmQRZHXTyu+g9g
cnKIyfx5VipEtUJSrc7zVc15tKGFLOnOEuOZCgOSSNWrzmSoWXx3FdvepeektLLQ
5c8MWIieyLwz2lKuU7Hw+UFfRozPKCDw+k/T9w12FU8W64Qn3rhvGWDMYEO+F0uw
0ut74SqYPUulCJJlR3/IohI17kVr3yHWxlPyRiqpWjDY6PJrbyLrqlmBZjvw10oH
e/+Y+FRxeUHRYOMoTCGX6QOXn2AOYAd3bLcZczaNb11KU28dLxuO4AqyA7ZWXV7/
JWyTNgkbcNPQIonTHsFqKaAIOJydz8Ho+ioNMGQaj99F1hTmbOZ+rl3h31IffcT2
NFh/FJyX8r8CT/wzmJnLukYmjnxWVlpd2eIZIYn6rhCOgUCr8JT5FPErS2jvmBXI
V7j8GoNOvRNm6IyUlebsrFk2ovis1FNfb8VuQFZOK+GIfWoCMXlAsOPrqrSGyRte
PkCBFvI4dWuLFmlKLaabHGavMb+xFPxb4ku3oRk862j77Vy1DOO05g6rrm6Xn9GM
yUvYK95z8hAXQpQzMvhuUjhbEsMCJOQyyGOpx7NUdCPABZsoP265vJNKiadLdeuX
Y18eUwvJhOndwwLn8cLiIJRvxSqnlOhl41EKIWXTBqcMyts/KCvlt/21HkIpKOCQ
i6MA8EJT9HOBAQLzXDFzBge84rDu27rY6pB0BZlDg4Iq9vMHELIuSN3bSbXhz/mw
aWz5JLXr4zuEOeTmtSMemVWhAsCH8/DDdNNV7MfT11fQP6xmsZemPjopaAmTQ2d/
UAtO40OeBNGuTSjIr9RLQT7XtmoND3Wjv6cCAzZS1l6wZR2o5yKUgC+oDF7CdUe5
wbE9LIwG74wwFtmirXEl3ffsNbsfQy63oRFb7xexlrbTTqjXKEu4Bx7lvHRXUCWd
epaVm+95hUj0G369k/1o9HIcpszTdqKQ5EBmK61ZLIn44K/qX71hj0SPn33e8YN2
Qu7oLFL2I7YQiJaNuetB+7lD7nEYgxclTTfNIvT72WH3RszpMrhWjRQlx4KYgq0e
0MZ/g/E2xV8+oHZQfB6HO6hCV/AEh/+yfaNHB6lUFJOJyrEVaxbin91HXvhKOuQr
KWDtVvo9BF63F/T//rCcSuRwxhRZ1AQvWVGbCFlcvBFX9Yo1BSw3oOjwuUWuR8px
o6sGZVoHE2GenDz5fBpFmOtHeHqRAJixhzaNWncAoHd5tlhZE/KqJkYkz5MflRt/
2Zmooo2BfpAzbyTVIX2BH/0n3yN/hTly2G5WpHWFR5+tyFrBGdDh0Oo4iEYXv+LJ
OIMWA1Si4bv0F1SOsM6oN+9DJUw9LNb94a5BGTuMHgT02HkksOUIgRLQXEWZz3ty
+4pczj4p/ToQdHSPXG2X62AtJIb/1L1wsiZZQ9Z2XZoGEjm63diAnOf/UvHhnSvS
julVE36a+r4VCPdNix4BoQCQuCdTNSwS7SUjRg8EOj6dD/ban/nFRnhhI1iykkDR
lZXSLN3q+RR/dkGmPvMMrRO311STA55RVt9fi1cCgzqEk0E/d2/Ja6Elg0X+cMje
lbml93dAyxKUqYAz/qEQ1pzHDnmNUK/5cXWV6wOdN2iI1VVbK5GVES47w5RDxfBJ
xDxQweoy5YLugTs+Uy8X2bM6V22HyaJmmNOFf90nxnHvKD+F7EjoEyFxplj6kclO
ggWHvA1/QeQc1mrApxYCFGJFo/DH4yb59LmBqgSeEkQbruyghNZzql0XqbGKLeHw
2REhQgbejTRUkvanbgIO0Z8ZG9a3zc1eSg1dug7oN08zV75it1sy6FtZ6sfYa7p0
32mL2vQJUOLBwPMuPIKu7ey2xDZBlWI0bSNHa6+HZ5h0pKhCB+66gsv7FV1HN78p
Wr0CYqzw78aARIQxEJpiDUJZ3R0zhyu0zx7EgieQAeaGMrvOWA4ZBNbjJQiBz0JC
pJcwFLCIfIMwLpvbeuo8KQVJp6glRjZ8K8O06zs8cPwxxQilG9ZId5WFyiTJsej/
lBnOGXuuW5J/SqafMhXiiRW2cetDA9hIKpAZjg/YmPSfcqWnP+7+F1N6DrbmogyP
MeoWY1FgV4B7u3HoonWatRINcRoeqFE377oFItt99FG0DqVBrmi53qukTYgYj2fd
fgfirWk/ACdQ0cC0+M5LKQqwQicmEItIkbm/RVL94+FKDOENCOk4MlwYpFAFwDH2
n8ExoUEOvSCctH6EllCDjFsS0lOOnIIaYUal5LlCqU7yh+RxRs/XM+aG/JEgLEo9
tsdyQ4+FPD8XdIDcPsf+pdOanqCR9cTqJKmtlBs16rNCj2B4I/XglJs3e2DrZt0L
ByPaulyxpK2u2VrC81FUAk4WOjpFQMIttvFNMC+ESHcOO5uYkhCz6Hfp2s5XK+4I
vdwsb7a4k93i61HV12XoIl2e0dB2OeFcM2nzl+zDuvvRoTZlVIWkwTDQCZUxoHwK
4muPVC+M3DPWUWm6Zrz1CdDxUOdWxDdZ5DNc7iYph5tsqPYwV81c0mpWyS0oVS11
75I8+CZ9a7EtxCa1fNkHWH4JEo5t9hz5svm3vyMGusOolfit1oyl7hGqrCpTYHPz
W0o3uM06HUYDFbWbBge6b1iE8U1N3K5/ePujpQLFd8uFBx7vAksnZ0LgteN22JKJ
xn/Jbh3tiJwEYp23akbPMuuzYpBrtgcYxA8sxc90aQqPGo+ICH/bXsFdOMeUABwY
HtCmYchnSocnm6pTTMqr7ML3+GmZymXAjQTjEQUYcdyPoDOVw3/1q3iSHSlzTEk8
oth8pCWTkW4EfOhKa+drqAHNC0p40/328CoNrY50JvyxULueNiGI0r1tOlDI7glN
kdXfFRaN99SL1SL2b0r0RhM7OoSqZIBsyJzFimL4Dt7kwxtcROVKv8eF0J70zZNu
Zcz98tXztxk0+UC/VIr/R9a06SsTMwKxC8ySI89/JveavmuPoXC/CwBKqGWUPqzI
dwKf9t5fujcTxGN/3tvwK9z+WE5SKFuHNCHtO9SW2D8iLcadfJTUJNDY3Cv3ns7j
qQlWNdk8CIQkcj7xXk4+vVAyWI34oFwsOnIUmSDyh55vZ2kzQJyIw9SDlS0S/EqD
Ykbt/YYvxxK+COBFL/fAhQv56V9MU8Gn6IC5uIBnr5U/+dHrMq/IeRTZ/9kID/7v
XmWJw/rYG4RabL5DSUWG4UCbstrHM8QMRIgrn16SZRy0FFg9nuhFKTZs3ZnSbTIr
+NNWfHsUNqsjU5skGbWCMd12eB6vIWlqlxblczWqYC5cEHlZN+xXzF5Vty+j9h+/
N93W1VDPRyVzytmGoFA8Fz+7vktifkqlGfiwefLeG/rjuDPXPUL/YRuI0A8OAAXR
bCjE8xTyaZg4MtgI6khoRU0dXH5/fgiRHJHDLMsrLxit/6pjOQNb5rEV+MnNsCfy
xvkjQDQz8wrvJBzbL9FiEsO4YgJLRaCNG9XODPn/77Y8Yx3eyg5VEZ3yfEq2LmZm
6OQNh2wQ/I+pVtUqh8MDhEGsW5hdl7ELgdAs2H6Ww3oyGLMQuLEabZ58h9fNjvFG
ujny++oBZ1s5iDw2jyeiNXN14EdDAXdg3Wb/5p5ZwEqauNrWVH1OHRJ1dWoLrqBd
CaPtXBzWqQwV9mH01qlox+7STwPUsY6Y8W+XsTDuPwl6sPt8u7Tek5OukaLGa8Zo
Xv/+qeK9Zp4BfP+cnjjeYND6FCPc3y5WK00QifXcXmvT1nx2rS8jyGwhCoO4LUNY
cenqvilgdr5CYDKrGYZLl1ezwmZxsQf/8H4TjXL6ymOItK28USiLUo5kjCgDhjM8
2W2ydf8hDVPmU3ZIn3q4Gzasv0j2kUEOvzpDk/G8J5dBcPhAatyI/IpehOa7cnzv
pZLVmdH4LY0yPFq/GH4Neq+rPSHufhBB1Rou7Q+QAj4ijkaJKoyLvBDCdGoWfy7O
NmY0gBbTCCnXYPP5psITIYmQmDMTpHJmhwZqIg2ssHUD99gbj4vfffWAgzHe4vgF
fCO9JKCNyN/YLyPTki1KoJb6xzwaMKAB5IEI4FJ8vuVYhuq0CtalXsmOgzDsGqFJ
KAN4eUTAwZewsrgR4K6I39NHSBfnBBI4iUaB+TFov9WKwoIhPyfnX9ez7YNFmXx8
X0+cIS8NaNSYenrZOgI2hkFl8NiHKyBDyPPVzFixU3uW0NM6eOtktSWceTogba+N
dQN5ziJ0FdOPX55bssdT/VBlJaXTQ2rSmuqfsWUiP9fT5UpDEt+r6liNgYFbX3fB
tbeQ6xiskYQWSfgeOQYBYRoeUNPEG0GriiahHNe6SntBvKgliNenPmzc7+/G1Pmk
lPfQKkX06MRF5XdxTy3/ars9d7C6xMxdpgR3aXG4oHzV8g/gLOLNxIbeB8nSfUVc
xsbInd+7W7slGBg9Wd10DG9ebAkjX/mRbRdgX6Xsn7fb3g3JC5PSpkHnf0qg/Fil
WqziCE4wd2xn5uyJYkehmATk95Bb/Df0gW4InX8dcLwE7pzaxGGCsakQfHDenKXW
RNtZp5exL6mRUcs2aeOGfaoknN3dEZ3dJ3BYkEp+L5x3XKhjDXOLFi9smqZ80Y/n
9x1BeekK1FUKH7sNf69J5NtozHfCP2dGgfuyf4tCrWaI7nry8D8T1cJtTYAT8Mvy
WKAoBXD7cMSstl0SzqurhTNUmXg3CGX7ksQUGT2Iuaf8WwHmhCgj1v0bQkSqL98D
wg2NgCWSq6hPBmse8J0Qpc/pLZRA7hbGr4V21MBcys3ECpXu9vLM/TU+GQuwVNi+
fZ6sWJwDMAaPvCTp1NtAqmNwtKH1EzjzkiEN/JwPjm04Xaxzn7cYa+1tTcV8nrRQ
0h+nruMPwPQjxL568I76JwmpNX6TV5atSFhzr6JY/vrLkTUGkqaUZBzoZo+4n/M6
fNVwiLdy5qpr7gAMj6p+pImAjXUOnj9YR8UfyWdJVIM+5eKWdNMx0uYqN4UrHj+f
vt7YMmTQsysLlBmwIJrAUVrbYPbVNz0g+eFRhL7sxjXrntAVNrWFnKoNdAwm1Ns0
k2kB1GuU5paIofSXiTcgrNZl8U7gA7a9Sk/WxCy5OBRoiC9MLh4orSQpF3tcbhuX
jBOWFoT2YjHkr27F8oEf7V5yYn0x4FhnPP/62RBopKmb97nZ0PLbkmlgVGst9cmn
R4ItWzVW/UPVIVh8aaoxbteUv5hQEhDQyOkgbwyS2DJmKwl3DOFJ25mUg8REJvIt
tZ0nBtsLdzDFbJgF+LQ2lwBP9nRIJIbueYEwq4ObFPUfTFGLYYsMVDd0uGPH6w8w
aA0xMWO51cAGLJmVwE4ScG4Jbs7+SIif4KSgGlaHFtwF0Az+0Czoryep7ohzI4B1
zCYo20M/2B1AfE1FxFIv6LlcE/e6EWSno3/RnlwQVqjiQGMf4UR8vR7rqX421ZZa
/olqlXqWHgMryAufNnZNor12ULw+YbepgvMh/P3Bj1z0pzS6hWanu+VkNga1sUo4
lkpLAAkB42ldoTLARy0hkYe9dyFXi62WsAymPCWoUG3YRXi+s0MIisXAmJeukfC8
z9sypazy5bK2GlPxKyIBXXlOhlqBu1+IBswCrLLaOwXkrh10oq7vfEBWlHLMPguD
WZawGZ5xtOa4ZPHb7YD0s3nUidYqEXVVNwAy6rjVUD4BeUaJGloZ+9sWdUZD+YNu
Dc/UiOkBPpLSALvOvz3eoDFXh7FERXQdM0FdZJ/kNJSfLZ4ocuIu/wVMKMCTQ66W
76XEE5MAIgSb+o1iLATw34ZVMwWEmdZMW9iIddA6Bcw7vLVc+iYW6yf4Jy16zXqz
Yhp6IcFLwPGd4QFL5xMrATpIkqJLtpOlQqxZkFPX11+eniORtAFE9+Shrlyd2Tnj
kR3dGQXoDpjyahnPoG85p2Ft8PAeffPIpyl6DlCiEF+Fi5wjvwCR81h9KDkDyKe+
MmLK/sstlY5w/YlaKlXKF4EnCfuzLgAOblRtQx7mkuByNkVGLJjAA7Bv2XbEWq22
a/SITHBRweOBZXtXxTbF4ySqTYDcBBv/mJE3e1dwm+3h4pzIr49fULd6mt8udshC
wI3oH7i/NyWOqvMo6XJKzERSIU6j1nWJznV+qXxaJM9efqheoofSB3Rcblu0CH5f
HGbMWDVE8CzuxMqUBIsMc/ynOBwYdw30i3tc72E5YcYAbzuiMDXQl0vqQs5tY3oh
YLVNO1fAj0tBrBJTQNPHA8zZpG0df7vdcRRwK0VFIq34O3AIOUSZFl+3ho9KI4id
knscEAbCI2Pato42q6nq4WrsDftEaJenG0BloPkvmPvpr2tiv9IkymdBCOlwyv4F
NwhwlsF95hPLUJ7qxuH5fCW4MGUrTI42oCvobHOyZuk4DeSUQvt2/MkZWQ+WNNWF
PLay0mFG12+B4fu4VKek7JGqMayGiF9DY+Capnrp+TOvlAxVJ+JpuTQBcRJ4zIaT
ayDo1fISByMAbW4C8FgoJkp4ns/SSXWmfI3KY9oT8Hr78cz4L5QxxlUfYvc027FY
wCsoYmAKGXeeDCS3ua7uI3J1Z4psZ1tILlChlz8pxneQ8Xzvd2cl3MPg8SRH4Gvn
4qwtGeAAZgJPXrGFvL77+tgUdcromN7QaU8aSh6DN5cbJJvHUpJkyzjXZ8HBHjmR
m9xWEbY4iSRROeD8UTpAhwdH8HXxTH/RIETkkKtL21p/ioAFUIDXKDqoKBKg/Yth
c0bH003Q1wHLuOVSMrNeEjGgvqq3Kur/VXsEdQmvKci9kXUnxpfrkpxpjKgm+J5w
Tr65JVWfQDqVzi1UxE7SXM92u7yEnfAYuyTWK51cHT8FOUGl7thv0hzE6BEEEL79
wUGgJHFK3QEjA4bB9mMOqKEzJN5H43RUj6BUF/jbPtxT0j8VrZzxRJqJ0eAht/vJ
BOVJzss+dhKb1m2GzJ557s5Qe1NOQqgz+WpMlLE1phk3u/uC7zEIvEFbPrc1tKTP
nvy+8zhGB2f4i9GQA/dPgNHG5zKuJMq/xpOs6YPENh51ivIdPwpYEHpFqQvcpwIB
L/M2yylRMRL9p8bwk9RXx5QrQ7+1l3LBYGPfAhuIBy8JXjr1TXYyJUIi7xiBzKX2
AqKoSEdvI1gkmUZCFxED3TmyJGZpCVKgTWK9UzfzgdXxunbU7Q2mLXuTcnW88MiS
M0kNi9yM+McCP6lnPFIdYssG7IpD9ukCPuhIcmNJ8Yp7FoXIjhNe7bDVXB+78zu+
Gs4C4+Z/6SliUT6lM2vH/YRZMOgHW6qovpd6W6Z04Y9XG1ljkhyAOyh16PACyROv
A2GC/tUZMmzmL2lp1jhptYvDXEhispAHebbTsA2RFEVF/gqkGLl7g4s9uQfYqHHG
/BYi4PrcPFepUd6DDgvVJJH5i2AXdCNK7r4zlfj9H8roOEZbf/nngcDk1SQl+u1Z
0bCoENpkf47C2irKUuT4/v4sppNF8Z61upucuI8xZxd1vAMqjPTekNholw5QYDQ2
JNZBEfKj2wNvoIOOzNCv8z3WqCfhYjFvW93h54sDsaIzQa+yE0GH6pbS0fXiFlm0
MJrhz8k+gIAlL+07+EcgciYFSBdo+Slabu8RYKeYkanCpyb/mWlfLK4mQ+aKHXp7
AQvZknXVT6rkW2G9aWpanUNe/PIFfs4b8RIFYOkaGGXTYMIATstZigdFEpKMWcS0
yJu4CxHlTCK+udbl25OaRNHB6YyEb6wFjA7oLR131njQzPGtZ789imBi0N7G2tC2
IcJnlr0UN3Ds61aVNHDZj6JRNx9xN8/cKR0jhwnPL0c1s0R1TiavamYNc/O3rejQ
0kc8qWFN4SGAmDbWS0I1IcuM94L3ZL14ThGbESBR705TXfDk+kNB/61ShID2DqRr
ZHeAxDhvgfOA6t3M+wuwYzXN1pmJgyFi0cZFeemWgnUnAxEmtl9xC+uNCw7uICcx
bS3vZIQ/89tgTeYYPgatDtu4uRzhulr/Rsv7qnmf318/dlKBRyjsAyJMtnzxZNKT
SyTtOd9TGbioxMZm9+DFRu/eYa2BGpgszLk3he+MsWCZENBox1J+VZ9Asq20AkKz
3d56/+WMs7FXAqRhgIxF1Z9mUD9LeK+TFmhbjTVj/H13Nu+D6ti8iqucrkshudwt
1r5bIYa3KcBmmKQpYnW6kzfZF6AfpoLXDw93MECdpmp6pUB4k9jKQDzT+I1F/8m5
DLRAZAVjRmGNjiV/SU6uY6cSwHjxO89d7j/R1saSFiXVad5vzKguZYlEJAHjia+P
4f4jXof41tqD7BIsK+Qi1QL+WLQPhZfpyXVqeSrfqJWu++Cdkjj+JFAnp71uqW8/
5tgQo1haC0xqwqn6zNblcYRdKRQJxpXJDxLOMzoLx4KUuO+vxVTGnE/IkxZUb4ZC
i4LqhO3vKLIsQhdxBAtjpyfcISPKBjPNL95oRJFc2Q48vMUY7xj2YCsOf2h6TZ9O
DQyI20V0DECx2Bm+hIcfiA7mjQQZiAuK+RYEdoVI3qdGkU0RcWVl8gTz4Z/RN/nz
Kk3oUwSxT8DPyCuGKcU8LhgW+WelfY1sB5LqWVdZdVoqXaepb2CCOUVdaZvmKXpF
mIynDBGCfhLaqzUWFexCeJ0NXSo6sJ7jJzf11nZ8tdoUemV/nClAPew0WFij+TMJ
jcOy++WHFHca+7Bkp7ETYREfuQrDdl2/WFNRNEGcujBTD0+aseG+7i3EZO7u5vgy
ghctXqdxswK7mR5OD0RAtCOENkxrBAMKSbgRZ0vb5io9DSOcgyH1HxE4dqrIgRnF
+LoDRll6FSQ4e95Go+VM34AKAJG1TX1CmN8bpHdSmwdI4f/Z4XRuIDaJSHlYDiyt
A65y/tGBwn6cMV8ISn6d9PEUn5wzrw26BJsBKLVOiGPHJGcZCk59CUdf8rQftMEj
bddWpEPRuxfuYpLPbmYw+icYj9ypqj3rZtX3ztxAjB75OCFqd1mto/excmXycRQf
N9QmhV7jl7KyB43hJO2m/vPUtQcdZQTNW/rvSujxjEKn776iSbXlb8hn6sAbRsh5
bH1FZpwJ500gxRKijxiTReUAe5LnHRSt8m7zT86noxVYkb1rYJJTt+XFVufZU9j1
eXqTJk+SLc0PTCB8TmdT99s9sH9U+pzTUmePASx4BIWEbHOdXLI+Gb5p/JsNienV
efB2OzBmcMwZsmies0nSWuOEAy3m0EQK8nqI/6y2bt6fZqiC5Q54Hqj37a+9wZUQ
iUtuPg7dJ6gdMEFrwKQZaC5JotKbyqZcnCwOeoOQgnxo9/Nm8u+/ZT56OV00O5tD
vcA2SdhPtW1ZhHdJFIxKw5JUTImdLS8kWGSKFLZm2BbYKzkMRr7OBkIQ35FPPWcu
tXbr5x6lIZoGlr1cB+5h2oHhqTaqr4rOX4PJmJ8v5Zl/8ndq2x2PvaZnAzqANa9q
8IPJejpRn07jQ+SEktrCkjVqFqpOfFEgwg5mIhvrZ3UnfOwfA91CfdHc+n80FZ54
3EM9P9SDQh8Noaag7wBkxIRDzZvB34MovQKxmvOBI+aFQqtm/w95IZWEjNbvf930
tyLQMHcGtQqFNuzh1bxuZbdXSoH56j5YNzJybGjir265+fTH7Yy9kWmnVMV24m5A
KC+q+f2pLZP+fgko0wV6il9DajAVYv/Eadrh19/9SkmFZvuNFY3ctYNFVMdQQnmQ
6Nm2yrNfzYN6w5xQ1YrU3PHYYUKUPg08tShBmvvZs43cG5sGpMSe+2EEvQLHvscu
qbus85OCEV2cfJ4eO0sFwc2+X0+GyOcZ99v2iZ+Qn5lL3dHd/7fvIm95mf3BZoZL
2Zw1Dd+PkRhYOgDnAiFL2o9qqS0z6r9pE/9oBsvO80tPVuNG6cyCvVV+oKzjBaLM
ZJJ2htaXm1QnrvnNquQUJjTGi1iYT1mfSBT6u5ZfxblrCEMcKGQTXFSgvRW//dl4
DCll6Uj4l89HkJfV8dd0Cb7NDu16oARJrgRoQkN4gJBRcEM24pcL4qqRDVQSQQ4K
EeZ5rxnEMUvNvYsdoMNKEDN6Y1C0MUgTNx3A3ExO0coIp+H/sjsNwJEOn2Fl+4XT
n9WSx8Gv2BIEFQrNwYUAoJeWNXG1fkN3kOErD1SdplB4C4KhlaV0IFI7uRp8lPuU
InDTp7ad+Xaq5oGtdT3eqSoziVtvl996OAR4EQXwkMpyANDCT6HCLtIqGZfq+syF
7S66Tii41Zjd7+lLbyL/7+seUAc8MlryLeqhtzWRZH847e7ccof6pAmbK/5q08c5
LTvsAa4KYIgKqlkZI/24Wl6c/6YPgoNMuOYjWEcTg46eyst1fFU0EdtASc6djZcc
bgar8IDH3Q8JQCW81QTKoXlDo0QmA3hHW+xeHuSrxK59SrSr0nz5R9TZrYs+mu94
qiLBePPnXOsh1rJULtgMaVwwFh69YltiLc9JZwfewgPpewgtogqVkg2QxCzNXNPX
PCmiIPzUw19Q1ku8/6qofUtsDWULmdD/CcRGirSVmg8Kw5yev88hV1aMX2/yrDfG
Mky7trwZQYmum3hdYi7nDKR6KPvQ6z5NWTbVC6FeQBq4QyWl54vj5YWXoS7HMIw2
uxWnLBGdH8UJfKlf9fAWCEJgoNvW3eOQAHdRT48h8vN0YR3NZEbU1KGaY2Zd0QoV
DpjG6Mqayw0CDAhMK4N6+dlawxVEHj2UcLI2cnTaTmjG8Pc5HS7EQLkSpXHejtOk
pRDtg3LGdvEu68tdwXnZ9m4t8hbVWVFE6jFxoJbulvxOhU3ttdrE0H02FonbajI5
dhV+ONhwIVCOtX7LLbApwmTKqCo+CvlThMgQyAbwRimLPvFClzFQDJICHHBaC0v+
wJtThYWhw3gSrOr5Kus9KWIShcchHid+d05uBjZcybwWnSQ32oFLOiuSKfSP2LGZ
yeoZLTHKFpl6PR6ug0QcBszD1J3B+CWbvqliEkmI6D9CWrS11WhwgUH7+of5Zyxg
r4HTeHuMKfrusszVWw6oVGemVKPdg1rNTb3SgWfrn4dax0RHLN5u7HgmMaSRZymq
Sm1e4M/HEidPvGnFJr2i/yR28PwSsyflXmQiUwikmI1Mpq8z01Kbu8d/EErA83aT
OxWpS8r4dxWDThHpisoECHN5g2PQKW2QnvSDInnEdZ+fmtaRc3OsNnX73tdtAo5H
W+GaPR6UGGXcOurBaKLbSCV7A864AjNnfG41+UL/OC/PnaipK3JpYzTrH0u0D3hq
Uut8wVkSuHv8YDY+mXf14ioZZ968lAAwIQOPvCnFuiEWaTgkUspHLjL99EYD0+Gt
jcMRZlsnmZ+v7RDyWAkPHrsnE9DJ78voqmRUM/eC0Cq+I42VWwDQDwyl6OIpywRx
5cLYfsqInIcQ8Tc28kNsY9uvwt+nS4xMPVvhEJBDyzvLIW2v3UbokiUr7wf+VyRP
YbQL7AJzDpQs6qDsxtPgX9Lhv20FkddotyXvrvNOHlx+YU831wohSDgd4J51RObM
yvlWlsl4YJEXirQa41KLXn8gvY8461daQPBAWmA9uvRNTHYGSr1qfDXs9iUBHiCH
oL2d+4LWZFyD0tBu5I1HuEPJZlBQNAPCnFZHfTnamNV8j6PXAZcqe2s+9WJTmMPt
6sQM3Tt2pVNZUM4fVTzKzNJg7NZs/IXmLT+LIyqZYk8KsJ1o5FGUg6u7f4DHlxVd
sG3+aWmnGP1WSycIzxFb/e+7Me8mJQrmVBaNc8bk+03V5qXWIQmUqn3WOhoQmXZu
ZCnDIG99OX4cw0HMjkMcOAImPGpU+o3Yw39NYwW1K+nDl15NYHvem8W00fpHaVVS
E+o+lUnsv2zlKw/WpIdEo2oiSXaSKQoLUEMnMHez8cZ527X7OiaRXfybtup7nVMS
0dnD/Z+9Ty0tjM6+fKqVfGiIAEWMyJvVsDUrdrvjmvBUTDiZO+2ae+iMkYiypP4M
QufEYtk79EawlcbcrOiZg8JV9osBwzSc2Uwl9qKle7+ds/qk4qzV08wlgk015ivw
KH2VMgMkssHbubLaCRCqrcfJwqcRR09JWTzY8pVW5wwjHq0kuxchumNP6PPmvDrP
Wugo3s84h8km48ZKJ7ryrxrulNAdFPOOJfalBQHufKz+1lUNppLA2RYAnptL8huf
Tt9x2RuSQaFTZ5Cpo5X+rxDKVmiOmw8AIxZOMaebkydTu+aQ2neSfc2mS5T4G54M
tPQlnL/fYNcIisf0nUaENqHWkkELkmMfIptDbK4PCXQKgNQZvAbfWjsPjyF2yIOv
aNS1lDA1W/c1HN99ZaKboTjfJ0WtZETEUZqfbcPLo4Ciq7+6zYLWliIFuBkKTHJx
2NecXrsBOEgCSlOZvu8YRBLS/HVs3X/GrHzAtbjR7CEDg7ZOrwLMhYliCOVV0zh2
fxiwl4Y6L13xbZsLkGuKkqXgXWetlfdgHXdteUPABD/2ADiyGErlPUclkd6+eOgE
NJQJ7O9QnrcF8I4+7hEhxzX+1RR1NOD88gCWv/3MScv2zhkwKa3kWL/2lWjFy/Ls
Vmq9ZiPl2N/9URt4Jo/3+/wkro2jh+APDGrHlwd6tN0WcrDiXkyHAfNzdjJ+ijZ0
ZtGKShH7q5aGfgHw4g3EoWSXZkg4HEhtKMFzXVjVmUabnRLBYIal8XfRaVlOl7UD
ZerPTWZnW+hIAoS523ndad33XRMhm0adN23Qnk1u/H9pz+JqV/K0fjqX1gm/8gLz
YE/akS2P+dkQ7FOGBlov2R2eyEcmgySkPMF0q6TfiSAQCgDQru37YZQey7WNt0SM
YMNBom8tMdxAOgapPxTW14KeZPtYys9tVcTTHbxwg7Hp2nD51bqYAMxBZNqOSMjF
xTqAeppn8wnWGPz4fKSuMpN5mFqfAUGXY5ytwSs5HNI2BkWAmrS5akxH9WwR5c0n
KxXwm1iEap7jpFxWgb0T+aV4Im4v/jEeUKa3ERcTvZicvyOzSbIqeYEpYZceUSBM
kzQoJ040rmglO8k8liE5+Xfnj/O87ZhIKCf4FMgMGwrOoKH2Yovd4pF1MltcsgLV
Ova5pYfr6ioWOfHhmgUVSYLfd7ULgsf6cFcVhAh/WPTE/UZEg+h7joAMev5RJhew
MGcN2hKVfJm+IfgWuuiTBpIKvD3r4oa3EDS8louPgWJZwgIcapjCMKVI6a0IdUF6
QI5AjDGOn8ehRUwyVglqDtoCN+JtERy3hYdB+QYBnOVLbFjg4YA1LAEiOg9x6PVy
pgqWXtjm6O+LI0SqGpQ9+GI/elXKrpjzJ84i5LrbcAghAxdI3UnyJ9gAqHMsu8xk
ctGYZh6xFDABNQeaxa9dQY008SMklgT2HZ6Gmktzxv5MJsVb113OwCOzjQ1dE/7X
iPWlVMBu6f7BfzZk6/uAryA5MUEJOOmEnZ4c0nsyMK+HolduGKZgoXPsYpjRbCcY
XihfcgjPKN8ARZWvk+oYJvzZkkwzF3jkR32zoq9QJgE9VY1AlCZk+DR2hSGr6Udp
Y19QHPa8+Re2kZM3REV1cNmpV/MA6kdSa3Kl3CjhBSbh82nsNSLWKocpFvz1oiT8
DfZgULkiSBs4bi01qE5MiQwM1Tdlz2Af9+4UD5c8qJTV8oWL3Np/oVtrePTIIidq
xlfPX1JzOelW/X+QGt9XZmDHed0ATJ515rBWyowGLhRGROugwKATbN2+dYC1Kui8
hvnFJ//qBGcs6fyaS/jsTZGTqTuofs4rSEtyaCumJcjmAiyGNe9pHonUWEoOrMoZ
lHurWIm6KZjVzSFMm1uLM20jfFO+a5oTDD/gwhk/Bsw1SG8yGgfiarHxQDHAXpCi
q/7DwUAUri/XNhSf+To0qHdqP5QEgvNva+6Yab9UGcpl5YCgoxk0LQsxgCzBL6ms
3aEYqQY6W6wBk0oANwfP8+4cuUW5coYnJZJtWoWRYLKU4JVqurTqstPwzXUsf2Uc
rHgHRqGYz9/b4/xvnZUBVJRr4O77GQYQJ6FujNAC1tBJ+7S5SNlzRCwYj7tPEwSW
X1Xlkx6q+qu6Fs2hOGOrR7rVu+PGkmKwSERhYhtI/ONcJXc73eAB4t2cAVdXjVh1
eO6qHo4luYNBVw1JzeWkFFMvt61w78zLNH3u2od5rsKRZci2/89ounixWHHsdNM5
3lXmKRhi9dRRH7CHmaEwYTIal8RGmXI7q6obbGvmRhkQwNpWc5Ro4wdvUwe0zPd3
sP7Wc6gqrYqde3iGLNGkT18+/ETHJGoMp/nBySOnZT5/hBFN4V0o1fRN7sT3jWHG
lkTxfdX0tClJ26Mm1o42n5k8YjQSJ5hoeYNbHBDWFiK1Q6uwsFz7rRJ2CTjpaVP4
NEKba0+A5CFH4ETJ7CB5OxHyb3rJyfjRNAyxuAdTOwnqWLHYlTnmrHXj61XyfvgC
2pWSEswV9UhOHY6C5pMmQgnzgh5Qq2K7SJlK74ZVvefepuUFAt8XhEMz9pB5as74
KMj7KxcO8NJs3PiTuKUcDgkVRhHCVlveKKajCV6U2Wd1m0qx6Nl+wlrflApPZb+h
iDONZRA4+x1bcQx/DM8ZF+MIc+8sFihTR80vR2liz0wMk9BgRL/uEp4L+D8JVIJ0
IAsAswA+B86hlZZV2Y8upMmmJhcX5guWeS12RcIa6UdljtZgcWJHf/YLeXqw4Tzq
jXGxz6SyT49OmyaEa4esoYhm/ZjKvAoURzX4Qz3UgWhLESNiFEIDPIeuDUW9ENuT
tuBufAdY0wighfgOL30Co3fc0kCb1TijYUODn51ILUkGcPV2tOCd4toCdXOuq28L
TcUBYRWZfAQKXQKg7liUtT6xAqiaZqA3QyA8id4URpTbkClHuYfE0s3/Mx5XruW9
GjcT0ORXklPHjVmrMrSZTS9zU4liqIRJjKfWbydNftwpubqw8dlrkwg4Hzjtm3uC
/U8lJRn8rGcpPmxE57d+dI//6VPunrJPGI7OhY1FD9hKj0d/6BOc1knk6HiRBtOw
0f2kXXmCrNj8rwO95N3sotoR+zMdIYVzPwm4IaJpNBosSbNaAFUP/mPm5CehVCYQ
9K3+V5N6Oe522yJVKy7R9asM2T7v80VRKRgxjnt0DO6tpnvP8ikypaCgx20ftK83
6iwomOuQxx2omMtDHCKE3+tk9QRFdbDSkM0zQP4kSJkESrVdFz7knYtDBj8ta8k8
HlPTp0QtFTlOEfJm0AVoT2nahpAPSz04VIWRQIWqWlZDzsSyGMFAQ0wQKkjsHjdT
RisP/KEOaOAWrvZOOqHKrcyQb+3umhV4rjvsqhc23fdQodb898hj6DDIcoYD+U9A
ZEozmugjgptkeFX0IZfzH+lLDw+G8kmtZc+JbbHvyCjeHZnjXdsqOMbPhaCIxBRg
SlrC4U5aAunPKCyz5wo2q0iG4KQYDOcXNR8Zg4L+58laJ2n0KQim6aGiuZd2p6oR
L8sjIl59L1x/JXAdDgPEESrE6VWz0kIc9ky2cCBugAtAF50uVzEOKCVMA4jvcbjT
Qk5kZtVG7veDVG8PpmUoUSWk631XlfH7iRPUR314U1lfn2SmdCnPVXFBGjvNq0fH
8MEvrlwZdyjbqXnF1LAQaY7QrsJgykGCuAZ4oXZGbMRQet+AbGdJ/0cAt4H+Jag1
FoyZOhGxGIdhyeAjs34NCLEohP96boV9xRNUiGdy4ol3Nd+65txp2qYrtuzikSVo
C9uLaOJQNbfJckY9vmhzbJMCabg+68eivZ5wUVQ8ZnrmOLENCkQwpYns6EerWuqp
WcvoAxstLe9Jn45OTiH8mXw3jjRT1wkUM8AT5zKRQsuLrq10AA71Kz3Vn+SFnG69
z45z076i383QUP6GbZsrnkeM0itwgfWWHxlwG1Fd+gkSVNEkTh3HSx0be0n5E9vo
COlGzo6XunKUfGOC17JG1uaL+pFeXUDphiO72l+eDPhEMtlNttkXtCpYmAWUJ645
Spz2aIPehWzdVN0OY/42ldyQ4ihTnTVfvtURpA2BKs9qqecZ8/bGTY1FNsrPAAgu
09LnWPT7VVTBpXSf8ixMVieDv3VWxpnt9ejMGURs3zgxw+RJkQTjlJSzxRNoSznG
Ity9/Kk3bE/kT+H8Zbp3vKgflUiaBvaH2GsCv7g5z/NaewQJR0rCzQAIJ3z293UH
nK/qlEZhQxFdYK19CUT/ktcuDkBxjBOWzMyDEmDAyIVs7kdCq9PYRpONrUVdG1v4
3r41aEhe9I+/KIuvyxWW6tMg/Cbuzyiciic4Om67bUBWbUenMwvStr+Ip6Mgt/Rj
4/xcSYetXyZ2yE1LPsHHqmQ4kyWKdVXniTqw5xvO9juBFCDf9oUIZOMbuGLDCTo3
fLCUg1xBNw0ZZuQgLGF3cMpWGM6bF0ILlIaiYW3UXn5k20mSZvf8UcEMJvgI7kZL
V+1O187VvAkr/hyiZH7TDqCIJ587MWfi76CBTdF2T5blgRu77X+0W9wKdSsVydou
3pzmqpUXdSX7DcfKha10n1K2Pi6VMgmWWEFfS4TiCH5zy+4anzB04U53Amx1pb0S
mbtDQIfNhjUjB6x55IyGsCA89sgjpa8W8TZvs4gAzJVQwTQCtWpJbXDQRUK9dFmq
yXaBG9pTOAMVKa5rQGgXm7vFv4HGGUu/997fQcOcq0xjsT5R8cbR2fY0vTofFJt9
xYpbwvtTjpKqY4CMpMzP5+uBXmiRRFJ3715BdHW1xemzoFb3GvgiMypw/+qDTANm
gjOPuPunCL2v9fpa2vh9V4hFduHAiFMzoQRh9qc5os/qIa0z37/pwTBkLd9qKgC/
8xlUSn1oViyqxfO4iS5qOcOcu1G1fr3RNEuGFTg4EwfE2BPc095eFaJnQyttHZse
rS2l+bELWvDviPUqET5K6XS7n10UJGHx09OiVSpEJV+4bhwP7KzyWSEqww6LgjIh
jXlUlyOyWfFjyZpB1qbcEvpSwf8LN8MZ6YEGRhYtBa/tpMAjCAiQSQb/LiJgBPTd
6vNIN0oWd6WnADFZl+qJqMpc1EicShxBWEllhLznW98lJGpbHzZYMBUX0vUkvq+x
DOGYpE7lpa26nAh97Jt7Q7SqvpidtPOIkbEssNwl4Zr/wUIg2b55bGIBwpkLmjf4
QTF3kbAfHv8lq+QKWdChwBoD4iNl3l3AdftnkaJo6++QTEOb8Ijyl95HmgjQDUVJ
DEn2VJZq27cmlp+qTIJLt8ix3Q6WeMI93f1DJSv0Fvbybt0y6Ok+ow/ZlSRkYCYv
q7b4/WOs6JhTr1G6pIisecyLXXjUTzRw5MiIgjFmAhhk2/FgOA4Mhx9syNaSIhKu
IpzZDbKpTMBnx/HztHl+Uex7Af0Qcz8k5yPRSgRECOWmGD0GWoQ7kEKScJMpG5Vl
avfXKwlqwdDVNQ/rvc7N7YXq0azSiZ77nwSv9dqt7yhbWcKX70IMXApeolbTexg7
QkxMUEvqoniGUoG1WE2tSylC52cHTpdW+KpAgo5sSznqOTPc8+t58+tvFH6zQGRQ
5fc8K7Si2kfkK3dbztgYHzxvygpYt4kXonyXgYt5UuRYU34N6Eok2Y/Zik+uxvjn
9NhkyydEZK8PfuY8J+3LNwgATe3Q6wncY/DQ3m7ih6CQXxEB9/Bc3mP1Mb0X3l32
5nZEqGe3WpgXC5Ggll8HROzjGIksrx70EqpGVDADivPEVk2fmLM7R3aD3WDG2goL
1EEfOzG1+LnEg1Rib6KJQNCizMqLnaKcnD5fRDOu95hsTPB7/v1bHxT2Sna01ylJ
dOTemRY6kUxzd1iybVa5aYbQh62UwsxWYSOpF0L/+qSDeAbWNYV+YxBGCuCzShCc
FxW2iFoC9O8FEfkt2wHfI0VOtAV2A7wCh5IeT8AWvQIeNT6sOcUXmm2iIZUhxvIW
LbBMUR+2PcOHxrqLxvlP0QDRKGZbURGEtK92RPLXZX2CVt6OB53pLGw/OQP8XLz1
pb2mJaQgG8nrQ1zvn5R9Rc6wnnxEMUt8j71TTabjO/oqr0SECxZdt279213hyhfD
JNHAA7NNiwnDPX2MFYMGGbyRy4gvzkDFicNZ2cKZ35CjSyKEIX2NhyqM3IchpAmA
gmrqMSq3U+mECsTtDQGxYGJII6btcpTyuUmb1g6oB2UxGiCRyznXwDshxOEWUMSE
4LlBGTGrGgPRswefLkwGMdgtqu84NKV9kXvoyDE08zI13NBy8Ze7NM56avHrIlrB
ntTS6d8vqCUCDQUV05RCgLplQTKmrT8qBgicovlX3QsAGQqUXFo+ByykLJveViiX
Izr3vnQMXOtG8/sKtioydb2J66Tfw4bwZMzBTtd+WkyqFpIM+W97xGXWHzdAQk4x
78f6OzlBT+DuixlDOYtMa6VBevYBFyhqmS1HHixzp0VkwXD5363uK3Tnlv4WqDQ8
kxYEFlqIpuqzvACqiRHa5jOt6MbnwP+VmuZygbLqfI+dWENVh6Sl4gGuzBUt3/vu
Rkp1rf0ai6uWZb7KZkwwtcbKPIlV0YJjSYDpdNHoDE67PHD5CXQckEpPE1fK237w
80aMkx+A6+hZp0U+NXd+mYprQE+DFB4gwIJkwuhrOS1zHhLRQk2ma0hwDBQtpEvc
Sv9a6JPhWyJ6KnD5W7/z256Qq35tLdtedsQypJPg2OJHK254guZcnY7xzNesaMzE
BLAzbRPjTw3FG9+p17AqWGXmX8yDo8i581F3B0oVtz0/RpE8727LgBnoZnCXpasP
Jqc2SJ5Tu2NisZzXjKA0as0eKl49fRawbpAFLrbYZJHqHJE4Ze0JXWqfZCi/tx00
6EHCmioyeEi7P2fXR1A1YEaDsalX+Jq83CRjoVoield/HgiqC4Kzk1ux/g1KmOZs
O8wz5x3H0rqgNwgwc6oMov0r+6CDBAsArRMY9L9iBqI3mrOHkb3+P65w0p7atxhc
fzIKGjC8MfQ7zpUR9bdAvo0rR66s3q3iuYXNBNWjc/sjohkN/Lri6hAYEJdWdl1G
4yvbo62ZDgJ0lL2Hucll6++vA7gmrW/cId2LL5iLLHUAF+gOIXnD2/eq43qbDj3u
MNvWXG/8+yFlvQJBN9CrjuV8L+kAQmvoOjRxbGOTFR24dnIByopDhvsSjwvMThWD
C5MphrSEvJyzOs284yipwHmcrP8mMsGHgZROaFyQdQlF2oDk2zEyxVZE0kDR47TC
iR8ZiF8ftwUCy9m2ugQa46CMRcOYemJiF5kuAl6vD9YaSFaBLXz1LmZFntlGDVJH
k+2sgVe4FgnK8A6qd53TuEmfFQvONZ6jSlyL+AvcSDkvsKncMvBIjt1wA/49Wrdn
5efaYB7qCp9BNAEAtYB0/FdLTqTPXkJX2a3yL2lRsPqKnme48pwqc8fgJ2EwME3Y
8bIlEiUtAzhYrf2JPrKntEg2SIESeU2fPbXX94L4IzYdx7ogx9HSY0ikoMDU86io
YXciMvA0uZ1ZDXthRdM+RWINd/OQUrmKAJ0CZHAeSf98YPjBQ44yKvqE/ky5UfFK
AbIN9QarDN/6QAhjfV899TLLwPP25BLSb5+FuVdUd2qEPm+cCuNk5NKNbq9J3NL/
k+1gMPD1LVf58sFJDWnxF5jH1W0mjsSS1l9eO5T3u0enC8UApuSrZbS0sHz5Mwdr
DW5HaJxMxJqOeBq2r+tOFwOLNFSsfp4mLAq1XWqdSLw4TwBMKo4QEvxR4EcWX8S2
Pyn8zF4udL/PO4qV+8OQsQkyf6cchDt6VSGX5yIEja8/v6E7+KVGqnv/Mf+2QvFa
+L1wmLl9YnRdw+fZ4t3JIOerR/RGyJVUlX6I3gnz1rteYCvrl06oNxNTyGGd+3cW
hdhfA5dWgItKce5zojyXFpjtQPXKPg7x5MePa6h/Bl1+8wu/SvbodCTdsRr7w3mS
E4xmMby1yKJQetR32gZoJo2zLRgexTp+9QiJjbkdM7smhFsJNCiDzmvj01KMPKbO
oQCO0BzVvcoVATef/jH39E912UR5Cw9FCBrBWz9mn97fcZTtMfh5IW7/gOlhUOdY
bYMUjFoSz0Z7aPP4HqvLPk0DgyJctbTLTCap4HhGZxDPzk+dN/7YjxtgjG5O9VVp
SFFvCqvcm5HQ92wzxQMilXXFv8jFVhpzZiX3zVa1rsFKpdLKT7BrdAWb8MSudV2l
oEByTE5LppKDTSMZ2ucxnfvEnztlp3Z9k8Dyqvl9lkEHRhqsUI4GEFxOikJLyP7n
6LVPsOqbdjAHet06Cf7B09uynYDz5Zq5f1i7GZhl1dZDol/vNV1P42B5XCKli6n6
r627SCAFqRX0l86ffbpE/g6lCYZc+JJUj+DL+FMPeKHSQcbf7KxYGr88hxuMRf7e
SEpTzid1oFr0EBr0IAdJG5ERCE3cGzUelI/65eevKsk2rrasvI73npIUvREp4kGy
ARVHOXdhmOxpCENFJlyofXMKitD/DBXC04n7Xjaf2GlMzwqf350aCRlnshN5Ih7R
KN1fePQl4+bYv+o7g+j671asd23uimP4nDOozdCIXu1BXYhTrO8CZDSRZA4VU+qW
E+3uXLhU2pYz/D71XhAt7eUj1Uc6XNMAm1rx8N6OWw54MrrvmTwxwxE5D+XCf77N
9Y/ZmEpRgZ5uI4OqY2HchYvTqu5k4eI9fYQs68P0oDEWXELXeVWFO6Lx0+NUS+WY
HfJ00MpsKcAuswZl3w/Df8qR0u1h3hHVxhjuP5uTpFXhQ0j38LGbaBU4a549STGK
b2klKUhOgRImmSyvQ6wTupBKUfeR2zXRQrvewNkMMGqXByVBYzEi9MDQn9kErGSz
xrqjmXjfeGYOD/sj58iwXqbvXBz59odMZnBM498b/s4wLWJoCW4k/x9BQ36RMWdC
4m6WfeneXcK+harMjQ5kNCPhqticQne58RkK1B+QCmFCt7jh2RdlKIv4KyxtB+o9
p3cU5Jdk9IxbZgyS5E1GJwouizIWcWajOQeQ5QPYplU0lIT/iOZY6M+atB9ckEYk
zj313w0UZ8ZECtj0RiaWQ2lERTtqUz/gg/OUy1aV8LE57G0fPJOa6yYSgMB91hFa
z7XX6hVRUtfSgO8TleJR9kqczCC4WMNrudqNCTdX5Njjyyk5NkWDHiUUFW7ABsJM
6UfOGNbRvIiDZ1zuJCpnNqf0QcP4MJUbN4CixT2wuyjaHc/9qThxW2i3CayC67o4
BFCugBOLc1lsq7yacP/F/1Zc3//fh1khJgr3Jwt460WAJ50GyFxULNhPaXwtKsaG
Gesvt5ic7t2ky1u9XsRRv0V2a4k2xxipiVzXJ0w7b/JUNm7lES+GuwZOdR/724Ru
/U1fD/2dtxOnl3YxVOa1Fwdjba2F3dzTfTVNPRwzZKKDhjHLYVC7c/fMsAnAo2z6
huUogcP1pRe/UQ/XkG+EEUgqiiaV0T6ku0260u9mK+Tg5ljij0YVz8Hl9SyJ8jP1
bDuRUC5t25UDgS6JQ2w0TQkrNI3eCExHpweVo6e1kCYIXbAID63BudlqRVE5i6gw
j0MyvFzaGtElpuEoOt4MAt7WaXbaZ8uxHrxNkPA3lyVoqmHQQPUURC9tCbn4zM8K
uhDhA3O6M5geV7DGumznrp3jwPvxpxKld+LbE1oDlN3wpxBrmUtGWdETk1dgokad
ozIWjXC72Z1SBfyCFwBoova0sQEfErq4XPCQZ5CchPOUoAKUSKyeLQ3CONWLGTXt
e1GXzNtLuVhBpXZqqIDaJ/YzhbkB5u3sZws+iAnsfIO8hUfhH+YK7b/ftTzR6+8V
tWC6Oq/1fnsb3CO+Tv0CVN0c3RAAND5vsTRWJOf5GyLwn5fSgpDC7iqOttjrEWFB
AdzsEIJiGqYQ0cAKZybETxExhqFYDbs+zksi2m1oCLrqij5MRQP0qwafyirPumwo
l2NbELYj9n2BgRTu4nem79b/+kXJFzCiv6Z9WqAM5FE/iEzQob3jlAi8yaRHVvYF
8WumcSMGDgW6pGsoWvGXU2gN0/hyqf2R2u48FNVevOFuFb0O2/KXDyBsEIB1Lx+r
iiv3bI81qJ6bTwJUYGyBGkmyrCeTx1+ppBwfXKmS2+wzieJht7DatNOfE/VBnY/J
EDivkHZQ/89kWjW3PSlN7fl8Ji/qChGtedL5AZHP/YsRO/NhJDlRmABS6OeTNJ5y
VCuar5zf1QJeurh1Ag7r1HCaUhSU8AwJb/fk32RarkEGwM33SOqq+Q5RLS4WMK0M
n7jU/MTsdPmbMe6TfTV3iulQvRlMe1z6JCbiaM6xrWZhys4c/jWRxFjMfwoGDSnK
HfT8u1rN8NTY3a1KAIzD2tgyU0l6IEjG8tCnamR9ro+0Ro+rk5nbADViSPRHM4mK
0T6yzZOpYx2uGzUNee7F8FP+EG9evAvevXsGvjtgUZS5Xmdj6616S8v+UpGWpVFu
52+mYpISZxYoTac97ssyyCgk8hO7ojHMzKxtCVyNXNvT3i4AW02Q6FSAGo671w8o
SRghm9T8KVJwVS6b6blv3q+udYsIV0tD3pDo+0EkH6KKr6VnSPujDjUwDXvDBdyZ
Kap+zUwZJu/X5B2h4CEpL5fGWok4KfP+mo+CGzUmPgfGE3moS4QFj20198+l9uSY
W8sVNOf5C1h9JcNUjpsGY4SM3hYhdlYc7zHBobECljU7s+RmzfeDKsi/LxrVL0BN
sZFN062+FGfqIlk1pJsD8nbDESYGbpf8lbwH3CFEh3mHaPynCnWI52ajwUbYmeKM
CIdPQjY/2+KNh8D1ZTTNTYSJI1VZlF3IHkOEedzWhYRhEIgIUsReNSUaO4jOQ9Is
qa7NJO/L4c8EJRl5SfqPvIRJYMJvT5bh6DhTJgAm8BgV6LvmPJkiDDJiAXAy7X4x
lJf1xyDWV1AiW3Yz0RXugGZV30CS1og7K1bW8PC9sA3QgjHNaHeZ5twJLpu4PxEs
CRtQ0iJIjuHj6M8RauEpPkAceOyx18n0m7/we+4a8jxWBk2JORFwxu2SvGWAcDml
6Aw0vp9TEZ1NbUQBvkpThSaii/do9P55Xcq+2v1M/Es67kBsqgGXbYQmUUL0UDgh
xgCIpKeRyJ+QYxmf4MjrXyJdDclPFTE1yx2tFMdX7OXoX3IwhbFPFAkJXKFKUmql
uqlCsLAqveJD8fi+wr0tlXPLOjx/pLNsdwOOyH/zOHBSrnfexpuP07oEZ5sQyTtG
4HPZ5E/TC+OwCRNkB3n78xe46ej03KbDxVkYtL77s5mFZ/TWeORFsQKB/w4HH50R
wzwE67KrT450D0S2kiW/U8sO25x/5/RL7vcqZlNvT3Uz22j26iSNmYsuqhIAxZCx
Jnxdxqcfqb06ys+YetgDveTQkAXNQhUs4FID/BwFEZsbXCeMEnuxTwcIoLqtHz9Q
dEE64QzilKjA9DbukMIkxcmVC/p6Dgkm6hnhK6MBzelI9AnjJKtZp6Ed2vCcMzd3
LzOpu01RhzWKmszq4b11wJPaig6/knHyJiBSfMKfnypGtiTVRlPsDWUH+dft6M1U
iTzvYt0z0eCZO5zXv6vFnu9CORSOVCrLfoIlHtenene8f1Qd7Mmkd/cw6zuTs6PU
7uWE/tDkZQbMTLRfERruw6Mjel4W7rbIi0Sfm/zgKGTFvUWw/t0d3u2UGHZlYura
FyhrwCKCrtx8xndg1zjUv58ALZmpruIx41WJjHHyiKa2Uwu/Rzrek7GJami14H3T
VHZ4cQrlmZNry/y05qeAnYx3IKGR5oNn6eSJejbEhicDKEs+mhvAGml4ilV3d0Nl
1RhPNg4UnanxkmC5Y+2vLZAJMxOLkPlbd+30eYDy2dtm2KihfYISgmwyta1ohgpo
Yjh6O7g405bYSoHqArVCKCA+8txNUgNxmmp6Pcao9h8+545gLoz9WqE3XKl81NS7
oP0pvK38ltB//l8JHTd7sb8ukxYT5JFU+QriyN6ufFc9QPjYwyXn8nV0ReY26OXN
37Mt4ENnaKU6PkclheC1QTFqpRBEJTSZqEof9QvlZrq/lnhBsOoKvbNJmt37wkiR
ncigatWIIJWnWUabVD3SCnMCJqeNcPPMYluAmhrwoKwJp0849NgV4Vizx7lKmeNc
et/XppTGOA+pjSh1++tEFxw/sg3a7/JXrnNEqXRf/UXFgK01aOt3QO1E5S5z7fER
27JfAgNchQowljk1qsUDYUEy9+I8vIr+6sKFB8Ej1jZJ5hGf20dLHDWGZqmQ8Ksp
7rwcHMhDVlWqkHSgyHItEixfuQuK9KAnLIHTYfbYbjT01g5eowuPb006lKa5BLmv
AnS1DCuhv0x3aiDmvSvb1mYTjn4VFtjWqLiHqGTwWMsxGEwvkZQfTix8gX484Aso
r7/U6i098xjMmYvuQcgJAluTOUUlHS7XzYZDXSEUXq6bM0xHy8eGeCS2U+oE2kgu
8CCII4+9Ti9D2AkpbBf19H/eKLim3hvixRZucmnPKkTB883+pEb8xe4/U/7JkJUZ
WpIAGE4Gotdjg3VLShkI955MJl0nRe4uygxIkSU5N7WQzM3PiYqEVH0YH4zek4u8
SrUUeRlvZ21jsQXHIKzadrgv21yR8l6LBaIZ6pLSkYLYeyajdG36VpLgj8rZijYl
OIkUMIbZNeOg26oTw0OjA6/umngXOXp6hoCUMk90eYd4fTifzPZDTrxpDZnBMGR+
UuWzFkUBRp9LnWJkgxOgBthI148bZcjTI0DyJnCiLDTASTDIaf9rif5YGVkmxI0I
vEKsdj8+L4tQ+630gttIVIW9mgw23//r2SWzb8fkT73zIrTqLE9oO+ZYr6cGJByQ
hc1XmxrJa/0iEPKsdtxNwVNlqLom6iO42a4ULiJBsvk+kkoljuZq12dTpXlrJlux
SpJeZIBt5aEC3MAyhSsHdb2rABM/435IxzUrXoyhRr/A/FAn2SCKrJKqv3iBQYWF
HkxtXv2xZqYhzEtFpg+77RzLFlV50msEE0XRafbSFQZnfU5tQvQHjTkH3n+KmgNa
llQK+VGfAm7tXNIoK7JFXf8nICvXNQweFXkJpAOpyrFhWd9UZxACFlkuSbU+onJs
512wSW9DBjSqd8fdIqDOEkfyMd+3wSrzfDfTVpBZfptEV2apiDOvxRTGg/45prq0
g1m9HPFVLZfZaH16rhLH9/ugBW1rqUsZeubTILsNRW4i5lxCxwH8ZLVdDfbvmQBz
Z9o6iS8EzNMmyd59GCRMTvEpFVzW1ZNeMf6D5MPFiTv0i4N94xN1sYPL1U1OR5HO
MV0UlN5SFA7BzOb+nKzhAsA/6pDYx2h8uYEVC9aJOcGYuyZ+FtXY0bdlmGpG8llo
eArdOHBwVgVaPt0ctCVPAMJ3y03ddJoF3ikLQBG1xck6DYtRFWv0T3zWncelLN9b
uSp0KETxnvn+KUIdLdbnnYL+HPaBoX4XVcIJPZm+SOScYFIlDWO3a0L5oLHvdpsM
xMP99W7HAVdIeaP1mfHlNt7xAN7diacvlDx+RAR4UQ4R8golA2r6hyJO5AcYHlL0
zCeRsz64VxFo+J5no5wrWLlIb4q+gDuyoLSxz3RfjcsCDiOufvHDe/osJ47xQBPe
ElnUtZ7asvDrZWyynQ93QLPsSHZuI/SsuzjROv9orpqA1SEUgTnwCQwFSdliTNiq
9Emjv4CuIMYz7aFXnyV5swcnLq1Vq4KQVNHlddhsbhW3aAhOvINul/H6QG1k371J
uCI58eFCMexhiiL+c9+mL28JS0JBbu8wNnjxeOQNOitIZxLZnbxGaUTnzYkpvy4l
0b5/dN3S7y57lP5/r5nsZ76Jrf2BqEMyKF53ZL+5uNakvRoFsmidZdBbv1JdhOAn
BFwkvz/kW1zjGgIj//QkoLAlTo6QIhV6afOdYDr3wOh5LeKwXpZYUhUmSrdNPFKh
YbMZ1drEijDp3cUz62yogd6/5to3pI/OEx0cdLxJM69wn/AUl5jPAIu/Si11I8L5
t7phJccdAsHms35GxJIKsfifQbhd+a4EF1ZS5DfKLWL5Mib46f7PxYsrEJqQkSAR
x5rT1dLKmy76/mcY0L6KVIWiDv1MbLnr+aHu5KTMa8cofcD24Gl6GiRR6Psk2ke5
6f7Ckg8Vc388ymhI4rDVmPj66yAmajHMPECjYI+2Nd2ZTIDVkcV0ia1S2Jzw5vMV
G5u0hyYw2Vdv9fpPlUUNv8H9lP5EVoK27Vr+EozBoyAVofNv6h6N+PRQ5vePF3et
8WTdFgFo8HYyyfs2KwwHbevEnBznr+iPxAI1UbkDCs4KMivhxFnauJNjwnu8fp/b
9WRmEcsnXvDhk0fiBx4ieGx36U7fN87apZKykswgAlmP6d7v0WWGoFgBO19XaXlj
Aq3gxhKKGk4ePb5WrSLpLy1xqr1mygN6W5js2WasD3iDc/sElILUFW2y25hFrWhF
SKGLAgV04U8EriZ5lWOar2LQD1Ew6WXlZqItVJjuI2XhxTzCaXHIVvqfWfM5ZRYj
Un1pzpu6dtvzITWVr5vGKf8EXg8vZiTpnF6ko3h5OrYnMgoy2h+we8ipwMa3QGuK
aIHu5sPtHeq6z4e/fDaqrNtwVnAmtKAyZuManCYzvYcCWP1rMFwD+O25853jh+IU
yPcHm/9v5YkxnmGt+1Ac0NWqNR2MuF67juOawAH96l4knN5oY/OC15w/UQ/hkpU8
ZCHW2cH47x4n+dNbNz6tvAkfjI2u356Bw9ak2kVW7t7yjW2d9w4YZDeEhgtoYwIP
6z0awHSWk5Yc3a0iOztmhqDn5WP3vwjHXEKOs6ZzlG+bvEA+WsKxfZd1gsn3FZIK
PBR/v0ZsGwBOWF7GlWJYYC4TfYdtmJSlZLoneQMl6vr8by4s/GrtXUFWJU4Hru7/
EjyvlTmkDuygNVB4kKNU92Kcd8LGjavuu9PS4yLjvE0nZJB8hRB9IRvI0gj/+qer
YfMM41FfQ7X6ow78ymAyr8iAjPV72kAqCm7dzRdfMn5tjdOVo/9If9INKRb3vYCJ
nCOvoxtR1fc6l54quHEwQIqfk9t+vGKOBnvaXDOxuKUY8oe2tVRBGAamATOtcKuZ
iOE3QlK7Q/p7UcVNGyhUsMDxtkUMf/O7B3z8liVE+ddTgmsZH1fLqtl3Xun9OsOK
a6+nD5t9J1sNs+6xsJoAwsF5K5ZjMITkAbSDTI62lkHJLIi3A+vuJeB/pJ/kgsds
qHKjlfRK7lmcF671pNh62CpE/41JTjQtc9cgBxa28Ogu0UhFt8/ps/iyuFbS3VW2
AGkzW1tgi7n62CiGviYGhaTeocGB/AVUkZXWr1DiNUqJqHWXgPaYxIHlZ0xecp3u
onIFK7VH7J1Qxc9+oa8ZcYTdV+HNofbb1EOs2MyR/WxXvb2uC11dJnLY5iZVbwou
8wS0oq1UE3BaM7QOijDPhk0TkRkp6TWIhPCsrcckua40qVEvY0qvZNrUEtrX7LNE
WXf6zNmT3hXp+O2MO7X65XTaQRHJK/6A6KSlPmQ6YniLXC3BrJb951I96A6Nl2OW
XwgVv8cF5jIKVRd7qRpusJk7Qv6fQqz3UKiVPF1PgYiiqB4Eg7StyeGqBHbzRHXo
Y3DQ2dsYniaH4oHpDMZcW5eapwYw5RWPQAgkrrJmOfSHR7e1XWw15wkGedBh7hrG
hFdV0ITBvKnIMxwJIgvEUQK/wHZlrO2Kfm2LhpxB9dLSZRzF/oxeuWcjE7hfVFXk
RBrcckNOWx04KlAeGJ5M2elpUtu0geDgI0EI32Du3u4tZgaK4PqbYKJ6RQ4+aGpl
VPZmrpd2zPsfWqdRgCskDbbymFwTZ8/QwShsx4fWtz07ku8je+7ivZr8cgr65xGi
Yz1Ohxorzr78N5AAIxY+BVu5YMdCYXxDxWUCjrXMYWa/2r1U5ysjnEg2NdwYA8xM
koXRhoaayrJD6IsKiALGooh9KYZZ4n+FD8b9R00pzXxNQPUgxLyfzg1DikjG+oXI
qY4/J0HVlQsglWuwRxaRq9cAysWpP3ApJV7rhc9jFneavlUEWsDO+ufzlinH1IsS
fp7dVF0xvGy1iYDjGhhMy7xoJVHuwcVqonTHXgIbPBk+vWoWhNOrreovshxbOP7R
44QJBO7uQKYYcQoUvs7FNtfjsukvTY0MRQn12yFsF01TIkBfxd3mhGVRi2jeKE88
IIMPoq6ZoYTay0jMvtKQ2JXrAR4zviozqGTD42RQ7K+fOLfByAS1pXxR+7xRbJzZ
iAqMXLJR4Tde2fLJ/BjwJLZ5JV/yiHe0TRW1+q0SSa6NO44XQgMPYppKYhcJnvOH
8eoAov5q8GghWUhgJB0DJXJqJt5nwqPKLRlcU+wawrZ6g6yAPQZ7ZE1dILlxfA+z
JX8XLlj9dohho2dfMmqyT2l4AviZNbU3jtcvljdMQmn4kTT87Vmzf66HUJyuprpQ
EWdfgj66JjUWMG6TK3rnEn8J2MQss9rlWrX/XLElnLcz0DCKwV/NXOlgSGS5zVpR
hUCmhGFcmLvIsvoiGB251Z/tmWp0zx3kv/yv3mecXiIUiXqODibddRvBAYmp6p/Q
KCaovvHhCE33tDHaXXzOEgW+gGZYVYFF+FM3gJz+r61nBFLu+RWM1NtTHOGUKWDd
AH3p60XjXKi6kSerafoJtqFAxD1JqH2Wnmka8LBE7mNuHQSW3dG3GeauJZMbhybA
CO737WHF4WWAD+6fq5+jOULOGrytP2j7gQHWes1XHHAONRXgGQ42LWb/0fQ3DlqU
RqLCKmjxejbKJpJsi4S+1D54aPSl83/kOLUg6ueAGwiEDbr4MpX38aAEyY7Og84a
V2QR/u4Jv0peCX1VAikU+GeFME9bIQ4aTvLW0xOQPIeuseTB6S9KCES8HklEYVvz
iNeXt6U08SBwWU42UfilMX/37beQlFi5jFj5rUETuIYc+77naH2Bzb3KPoY1zZlu
G/GybM2QYj/uRS5pxOPDI0874VvXxAfb5fg57js8TTbXERXhwwGlo00Zrv+NPnVC
engAcgm/fWfXNbE+laXifIPQgADzdh/6YXbxB8zIZy7MOFkEOEZ5p1FNkV5jIMVv
YpkcHOQJz1JMFpOjxRnYiB9+utRDnQLEY0D38QT7ZJZ4u9wVYrh4Ghsq9BA85+2y
yHN3/eTSy0mGB8c/usbcYuyfvRaVF7yTUrnqH8pLdHZc6pl0tLJi41ZUBpyA2Lmw
nV5Etyzra82naK0N0M3CGyH/ygEzSdgArzU41Qu5F+fcZjEu5v/MPgjUgDEQBuWR
M8nNShKxJbUavxkoy4r0fv7pqSIIwsZF0+sfEDeaZRBvGjO6mejDhoIe017Hn6GD
J2x7jlfrGrEqPvKx9RFNJM7hGUejnqaPu2AE4HemyqUdBMyQ2sqPWMdyK4FcyoQz
VZuFW9icLb+7/Ka/sOssC8sJSrgWECY6qFbYkm8NZOPx1DRYuiaj468FzS5bKQ4d
9HRrVhRp4gauGfXETLHVDVkXiuKhstkm2n7NQBdhaBwzgH5NdlnsnkUxWsO0nU3f
2/s+QmUiOyP4B24Vrck09yHdUP2RYud+gilqiju1yJL9OR9xat0vOLMAvAEw8Oyv
9JfOQw6FaiuHS6AwAxqIjStJOcAmxxiuNa0nHb+/kk56+LTGLhQVhEucxtzEhWEH
QVwp+GRNCAxOBSBL2qLPasPlbOrxHhbQJqvh48Ix/beMCWX2m8jXy545FTyAfmHc
QDE9nYxjEG4nv1lLeygAF2AWMzqd76oK2mpwwCvUsurjpOrjd/F8jcilDQsaUHrY
77OuP5z3E8Zz0KAmb3nzzVH2zMcMUuQ6Zpm8wkGglRL0/BKRyPjpsPEyTvrdyAlV
lpyNHCEPb2fCWyVfvJcFULQZCJo2S9xAxw26o6XEWwys7MYqDx6xJu07lWBarQj3
cKZUg5Za1ZktLVhtIQ2ufxnk6sXEX7RbhIjd2b1gi4MNawWVyMlER5dUWh7Q5djN
lZkL3zqoMNbseEfrX13aMCpZZirPjMAqwSbhYCtCqdU7gmibFx3dr+erfBwFbS04
zHgNiEAlYNAkBEjAZqfIq5lkFyQj77zsqdtT4f0L8qhMF0xd07cfioq/78FBiOfD
7Wi8BnqCQJbgDkr5yILv6RWH8qUBFWE3RpIJKZyNFzCjIhsc5Ui9d8DzCH4bz64T
gMTzfRTwDsJPNzVg+0YoUarPWRWiILBxQFYdREXpHvPK5uzLbQPIhWuS/CcV2u87
1DovWuFKBnGxwC7772ZAsIEq5Z40ln47TObroPxppjCFLR7ks4OCfq9ua32DZyQZ
MPFrwffxPfdfQDkw9u5L+F+8qIx/FGp4xnAf4uBi2JQ8AVrdnYa0WSOuRxL4Vguo
G4sQVlmiASkogxSQr2kPk3hQp8LojsKCO9EHY+o3EiWW+lfLUKlvLHWQmQ7hvB8L
47HMT0KiLDik99BOgYbRyHgpunp6z3SJRptPcUka+alZVG6MY/Hxnny9AHmmN+2V
ft6hogVrEOm9O95PpuuppVAuHIhf8d75GxxBa92c4YPSgHDi2qVAOwd/rTxo/uFu
lsScg9Z92C5+Aqw3e/3yUfXNe5J5YSVL6m1rdx464ym7A/v1pFb7CTGe4flEBOX1
2da65MC5uHbiFPUOYRgwgIH9VAkqNi/HjC6+nOaIHqS/2mNT03Siu27gyEf2OXH0
jWEj84b6rZ9FXLTzI3HXsjpmKTqTj/kZXjDfzyfwouswIzud/sf+8HrhN5gxVFdT
jpbr45HWAVv7GRgx3ZXzyfhc1Y2Bmml6TeFbUPYc3soNKx4Vpl29AHCt4XPdj1ge
kpWDUH8CGbLIYScyRf4DI3Q8HDCmTVEN4xP8hS/4ES8yhKX4aHgx30sYanOXqlpi
jA2tus8Oezav57OGGEOII43XyM4SFgf0CKg3GmUc/+VZ//+G8SI9sWeBiAmGuZ7B
n5GgNbIq+XwZUAJIP3STwwSiS9MkAbs1yzYLEPOjTaBS79oqvA3Sb7VbsKNhv0a1
Vo1T0ad+OSqKJv/5oPJcAvjitUW8cgLEv/dXZq1W5pmx8yGWunaV8JrMKq9OJV0M
PEbi2xQIuQ71Pn3fK93sYRsP6PiC6211GGAakVr704GgpfdtAs7ZomfUTtkVETRM
vfhdVWz7flW3B23xXISamuDJK5d9VD7YO6KFV1wUz/BYSwqOxTvEgF7Rp8v/D3Y8
Hl2/Vmv84N3HNqEp6DdxDI+t2yny1Qf/WUWbhdHJhZu7vd/mv8CN/tFju1a/Ufe9
By9grMDBEadj4iYFw2UpSu9yzA8Ps0OyrErGJD5eFJvBe/N12alI8YyZt+GuN3Az
8yLjscIuZZSBgFC1oG79RrxurjyLfp8z5GoAakYBkNvqMpMCCnHWlb0On4mOpxO0
I1haJ1XOUuhhTJBsL+zfkwYdE+eOLXjmKZomOvbwr12bXuflvw2Ku8OG4mryxpm8
6S8GmXJcCLBwPT4YthYIFob9uhMLo0pLbgNtNACAzry/yTWUzV6QOoXS1hTP9sBM
YFQC0O5OmSgMuLkKoMeKuTRTC88eM+s0Qyh4amb9TsHybl0MxNaInYMLz1ohR/1O
PgDeEgoi5YcCsY8cDQ/6253N8JaV9QV2iyCT0QFhyIkQbyKHcmy2K8eHRVdiZIdO
VgM6Rt4ExtMZHHhIkfOmowdPMOkoKnsgeHZ4ye/iwPwIVCViGD6VM+rqYj+868IT
6KB98vNmHPCCJVP+37fPyrb1vi9vW38YIlCCnSk5uFxCgCx0YCWZ3H8RNnm8zmS8
QlP0xTSAu3EcdIwo7U262gwa1AXecNwsmCHR2vKys20UmTGDvf/r78dJaOyP329c
lj5ApF0xdzsidm1Cy6uSC/UGYm+SnYSosjVaVt2waPt9jSp1rscaMG30GCvwOaqC
GBCgVYhEfGktQC/zO3AYs6E+LhMJWGVG3YDz9foWt0qKLaJN6EmpH4oqwz1QdBA5
jyR5htbwObzTGO4BoqD6WBgz6bPDxvSf4yi384n+v4+vV19kQjHX6BUdG9y43RnC
xoiHWI9ef5f5pQ08Eh16RaYO+MAZEmZidkw7b6wXJpyXFMxl4OLU2yBtBhZ/BHbc
WY1ZDs48VPOQrNyvA9/ty7FM4blYzoYDHaizCjs1Nq+Z1wSgtksoQSiZKS4Dc/KF
QTXVEsdSO/iYlS5mTC+xSjCPJ3zoOARE34k/jW2aBaqRrvI3DnIBxra4Wo1S5vyy
63X7+QDSmKJSYrTu2Px1t0ZWgMgKs0HEHBCQteaA2LMC0cnKbjuF1udvnFhup4UO
nl8z5ybl+Gpt2ABwai908k5agQfZjG+xX1pYq6pBFr/UrfwK7yd7We+0242DJpb+
Xd+0uVCPMB4xM2LlR8lBdt5Wsjo4P9GnJB8US06SGVV2fwpj7a5twnlj3xLha7ZP
MAKrjCKebbEqw8EpZSCADYFLe6KGLIspTKv+FH6b74Q645/KySa1Vt0+NEOUIp3N
syPIdNcMT+m9Hkpd94iZC0wzvho6wL7iUYauQ31iO8tmMLaPZsgCG6AAdkj+O7NA
apQTaXsJp6a7owvdXo94C4LdHYnKTLHTn0Vhmqgzs0tIbUSBj2oJ1qMJsYpKedKC
b6hO+xW1p66510kZN4V8BdVbRHUTAnX7+IsOrZNDjLniTfMmVjC8XwcF4ITqkUxn
MUbg/rFLvqYLOBgk6areKCknWuWkVqWuhrGKv4uEK0mOprEmN1QoNbBLZEsCGS3F
73l7hBmILwAse6cP5rtt2Ap73MSojBLPuwx3KEA8leufpYABjGvwQ5vsIWvrco1u
/dbn7V7UkgON1GJZXUFWSXfZscG9At9d4mYAScBBTupgqoLnKH+s0UdcNS93+Eh9
uUJxtYmvzLwcqPY1h8GNTlLn+XFYg3RCFw3/YL2jN491PEUSFCIO8yunaz5Hk6Zz
giBpD3N6MUmO2Mza33q1HpMvzu0W4E5brNMY2FFdGf5O63KyI2ra1/VpPvYOXdxl
aIYOwlvN8IudlJHf9VAz2rGcW0MRtXSGhktyhRZjlJH8vu9DIYeltV54jDqyBs+3
D67Qpo2BkphE41KP7ZVCQc24WYQOwVprC3z0hJVt9Hb8t48gFuFcbAqeaqK6bwNS
J7xEpsnX1V1Cz/QaMnWwpBabiPIs3bPOT1JvFlibi7GCEgFWhpuRVhdasmVBisZN
23UYNsSknBk9mb0BoVOwnQJZ8kKqyieNoJi60JQphnGK8maIC+V1HHVAE+SO6sUU
T7KCzgZ/UTHm2OdISJajskpalCNTV8EiUgroN0jmt8zGHAVnU5IcMrZqbLKI5K1v
wJBTKE9GkAvCO9Ao6Q3no/oGtk2BO6El7/jx2IF+vWx/OCc7ai2Xrbf41lxo5QD0
/seYMWOuXANLqqovhWeXzhoiTMnz6aZIZeR9jC/owrW6oaxK9SCRhNqG4LclLij/
HSZNNWxVVFSvAQ+rdf5pdRNpSUJ4z8QkJK3COnue8FMcmSR7J/nZZ6HVkxNZAYMH
0Ea6C7np/l7mSZAf39VSXyPiEkI8vu05am58OjZB/0jexbPPuVMEs5FY7krpHpCA
sUEA2IdTfepPp6+bbfWLo2WuH9TpHVJnDky84Z6N4IrgteaKh8QJxG55Th9yXfWy
3u5qctHASUc1yFvwLFFokZVKuG/jPdin7aQw/EisoZPBA/ziAUGzb1zYrEnfA3eB
Gxu4r+HqCXP3GahlAy5LsMRkpN9c4qYQUGV+2oX0Gg5MfZpKMfHY3iuaYJUQ1kjQ
6uc/2r4OrjQZpSBHnHFF2gRilsATiUXOd0OLj4N0+jDv/Dh4uZEvc6ZK3fqljb3V
vj/N9bsooro/Jz3QLwD04rlt/DzhFJ+Mbh6+2oZyk9kBUvAomauz+u79sIBFgkKs
Fl0f6ztK19El3p+x+bGHS6/804IxV7SYsVRHVkZyox9tqvXFi+40XyGWE7xGf9TH
XKcJBonpRBkAHQx9p+FkGqEoLTNHo03iqm+Q7nGIWmPjlXviSWxvAYngEkF/mRvO
hDLlUGCUppr/5hl1PSM3BoxUZis0ZwlKE5ulmGOwWyRE2nhBJs5hEXk9a7smGwd0
8VIZ+qjpWTB43E3ffmv2V9LFeqApb/AP5Ce5+6JzcFHD7kP3qKuzZ1toMfHAJ3LD
owYhulKAQYeGmct4q5tfEuw5VY/NPYNu9vDEQXhx+uSiCOTppb0jmhzSbMuz8zxn
FvNtUo657KVr0RKBsecEBnLoPoB9E1wQcHCK0OaIr0t43HPgySMBD/DNNfbjQ45m
2YCSLu3ExWDTlz1S8T6tWq60+/Uj09dbSZJAPxO0Nlfuif+4dIv9SpGm+lD04x/d
r2V9q/8jNzJFrpfOFAkf90wLox25W15jbecSBtRPVJLHFIu6ZiD/4J9fKEgc6Wxj
c3l7eLoU6iQkQLUg5gcvAxUIkKXaexuBIdAkMyzwPFVHvTkqqNjlMasut4ULEBy0
Da2QiGrA8zchn3S4OWQAd4iuXtdWocDY+bqA4ktvF8DJsjYB2OvngwM7h18BUrhS
PJFC88c7b2R8u/qXmCWRsMpif7jje8ZvGTdxBgKKzDPFpcxtKONYuk3jmQyPOVXK
lp/DQdEOeIqgwLnkgKco68VQ8D9Q2JPp16VB5KWeH5H2kBAOimeOdeevXJ5sNDxH
qrhONvMtQJ+WPTY4H9apScV/9TfYQA0DgYb1rWku23mp3rPBUPiQPK/6S/3bTgnK
LZqegNhUYTtyKckM5LtO3SfkNkJ0daK+pt2MWVPMXEbLnV9ZDWg3MUWfizPJWPvC
V589HH0Noa4dLszuFyidmcwNjHhlBvJ759Q5RrRX9fd6khEbJkKX3jK995/STEHU
ahnf3GdVVN0NV53r4nu/sjdBFXNPlIXcpUs0dUdtKfvIBQ8Mz98dpZ6oI4B42+eQ
ZHOUc43LQxH1jt1EvoxoWXQlaCUwpBFr8OHgSQPY9AcqzVjE85o4gdyTUz/4WY+9
8afnIHdcREtv6nP+/v7YB5f1FGXkp6J8CnAd34xSed6UiljYAeUA2xW0maHaC1dm
yFJZnUhnYETjJqObG7QW//FBU0Cfou5H2XFdFanMZypnbkf2+E68Mrcsjf+GRHFw
/g25AUH7df67zmz857gJ7jyiSdzqNb166HywK02rqeH2+r/lzLx03PGkXzPAQ0GZ
WNA6JdlKfzqDXe8O2Ske/bJsrfaZyDdsnai5wT1eq/x3biARKMvjyAPLLtoe3j97
+KPqk0q+bCgwxir2Q2JAeq61jswnW6L/IMFl9hmbf4irTCzDVqB5oVKxJjRt108X
0INHOBff2eICWVjlHc6tGbiXjJLaMp2Tt9/2naLnw/0Iq21zbv6jdNOvODzJXGm+
WuxunqaFlfq/c5cTSqQrRB9B7jGoXXcFlRBDhpAnSRIneMJBzreGN2LvzEI3T+XJ
EWzYEsn0t/8tQOTUjVK6kjCqEIxq7QWJ/4VOOzuDglErusDnZ4Tbb5d+ZF8BdXCB
Nyf2QqCnIjCQUxakd1pl8OLizmBH/Ma+uQWTLuejri3HmHh5nKQmGrMRdQ1wgAUJ
pgXkOAL5mBTQdLO8JQjtItYoE+YpSfP4H9GRGieZknsrRT5q1esf+eWBc0zPpPK1
empq3HHtpwjs/TEQAS0t8f97anK5t/m55aLFPoNcpnngcWrMOr4oCAy4SDwsaEMn
kT21ugrDYPgNluheFcspbhp8w4+09leMAtkk6Ed5UUypy2hE8GcuAmwHx5l26PaR
KqkrXmGdtDyzL4TsC4iXf8mreL9YAPsoySWFVQyMJ9jcvsPzLzZ3V6BDcg2Ty4DE
MU4fZusxz0OcZjE1H+WUgdbpXXX5WVC7R7OZ/n4zhBSM9OMtw40dmEhh99whFa3x
NDZMcPaQVJrnLeCdK3pyiWzyQ7XGxjwOO3U8/erXhzY7dKwR6b+jV68WuHxaouST
jTWIOJW3sNFuqo2BB688W2ie8YFoE4cFc7w57qUrNBwojJXAzxahB8Pp3CxCLDRy
T5SW6o8IP4WpxywlOB6WGdSxUItzs1vMoouLqrUbi01SHVmL1VLS+1uslNOF303Z
ATpsH3QZ5flh5lhwnO74ado2wjqW6FXAnVdE1RA3U8BdopNLjDnSta8xFS1WVwXU
nbZMJN9rQLfuO6ngxU7tHaY5GCpcSW9TFEMn2VkXUy0OtmgrAOVkTjvQmCBzFRdl
TSbUsDJVNwt5VN7ls5KctLDvQ9k+tmuYU9OmYSSQnTcTkyPnXS+0rID57s358uUe
2pncoyksWzTybtPWUOFbZrBEgSN2zTz7/89sPUaKHmX7OxiTptzjDbaXB/ph2P7S
RueZFTYg2Eq0p24qN/uXmLg05jUYI5AlcbryACaSpGJJHL2gtp/IlTwO1hnsqg11
0GsViFgJmOutUW4jugObHeW9k7dOPZf0jpIetMZpUEbJrcqHXkgPiKQYXnEaKYAS
t8bcpsnBYR80mgvpn0Uef+nDz28PrNgN3baMss/1fhhlVewRCeuCmKA1aoD09OiW
R9AUUHF9DsE3pee9dlpJ91wnETr+3q60vTnLOjJk/FsPAP9XBSSTuhWniGQboJlx
3E3sQjo/e9968qvux9v/kAqC4eGXT1BZ4JNdF1x7z3h41kZnoXIUqgxUrYFGgMU6
9/bQNVzibF2xO8bXsBKcu/BTpgwk3VBo9SVluC+Ax6wDzudFmYHTFXX1kZ1LSDsE
g2Qw2dPS9Ws9ZCq0V/9ADsOkD+rCaOIrtl6Xq27kIBZ+9RALJndDsUQyHu3sQHgF
LIvgc2xoFzVKJOx25RWwY7HzPsR1UDTszSpuK2uBcRfXSJKL32gLrNheGwAkmhRn
W58qPqLqGf1FQpPS6zjp7Plw89CnMsGTnKH1HHizV2tHzlX11EoPfH67W6u2Gws9
THi+nsKwo/ry6Nmy7F0vVQd7welzvI0E0WBzLRtCD02H8dvR7lBAIu7S0jxb+8K1
7JWhjtEjYQvpwtQOGH2jrsXZO6PDCq1QR6NDcnW1FxagnCJmSd1EpsP3lwnxVFg3
xFIOZANaI7lNsDD4rby15+2P2NZyrvtPwLSGCazBVmgVDqpPf94466ZYS/3q1kNm
MnwJ9JP07EUeIZDtuKSKg7K+EAAwwi3shyPTAQRyZQd5rf6VsKbQfAVQdZQPJ+LA
kDj9VTQRGuhI86TkpfKw4UBLnC9BMVH0qb1zsEaS/I3QN7j7cPut/6mcoe5VkMbU
rAitUgWVqpu77f9MIovzH5AeALQ470rh/pXrAqBK2d72TxUbvcu8bgErZs4V6GiD
5rSxAgB+fuhQQeylqQ2vGndoTSMMXd4FoT06jqsn9KNaKOilEatvELV6pOdiajyB
+0OnErWJaabuO/AdGKbqZjUEBOWPojQ8m+dvmCvZYOBW4xfMp81Sw/xNwsgrWONe
gORXJllWHr/XElmpd4icfFmizeGOVlT2iiclxgBE440m0ZKQzQ7DCAmu/bYoYxq/
om0x8KjNSwb+HQ9PIJBBwouB80LqDDC8W323yXo8wkWErrlRpVxE3Jc0jMx2S677
LQzJV4MPQG54yireOC777yo3Dk544AM9yn1DxZniJyn8wBB1346xJisvLOaBdwos
yo2PGc6uddG4ISc14Umn1tDnDM9x6txuAFBHmlTx9saJ6iEn9+XRgpRKzTWdETyI
GvTJOv4aRPgi6b2n7GgI15sZeV7itFh/jdeU1HKs1yjajBFV28RBjd966fiNoBQd
z99FBCflegOBTBs/JTC+QJkslY1kDpODxZNwXWJM+HcXRrJ5T8jPcab7y8OJQJiz
c+Ok7q8aohS8B4rFsUAxKr5yTFFzdP27RGUl4rejBA7clGOhfQkfV+58N3BqY4+h
xDC6W+PqRkcxgt1Ym+QyVy86sZwqMGUJ56VlRpy3EQxTYQ+NaDkZeHYsnD+SLtUh
RN4Q3LaSwOV4E5g58nDeX0zWG6JMmhXGk+q5EwNpHSuXTd9BgwlFncXr2EGEov/S
SGnwkO8bjw042cBC5dRUabcGi6PIa1pDOuCVLGbhmyPLI0XtyOAwEo3afOzPzpvi
jzuFrb1vQcN90lcB26qRIQsp0eayICUfit97xdVRiAMqD6XUIxWoogoUw/7JarzL
4ddu269HMwMEXIAq+nTe7UD6TQOTGiKmFtlGz9/geBe2rGkJQur8RbJwLEabnMdD
w72VTLEpndXRg5UsOo8QXUKb6YKln56u8BfVHtLiq+9tJ449rBtLFRrCnw2FVc+i
hKYG+xKWsvb3xDSsM9IdmNok4ZSjN90yerMEbgHZSHjWriFXiBoMTV5QqZs2yAWe
snwyvX+S4ae9QJhqzubFkTZohhWcKaX77tdjonK3lroWZCeSnDA+JQXLEYon3cp0
9X8fZIZyjVlwcU52RJNwLA9RMIj3l/2VWStcBr1dgXhhJ5zKkg8Oj0xI5kVAwGmW
t8T86uotEo9Y/udA/ieMY8ujrcBNQfEnkadm4/zmECL9SZ0+PSCiagZFSaCb6fzB
Hqi+VakHdMj66zmh6ievrRTlj3p5DxBRyiTqOIycjCyd1wJ9ocJyPJZiw8DLLDZW
3q+YMh6PXUppUSO1gtOC1U1RjZLoyWd8telcectPWdr613j4v68TDyoBUHQ+qM6N
T11FvPuGFqxsE+66h0EwbrpaEn8OSw+0JLOEVLfx/hF+e8tqQgf9E78Zl1i50csk
AoNZkYegeKnSKd2CaR8CsJLZU+8St/IanBdrzZ1OYfWYZouw82nMcr2NNd0Y6/Un
pzkp3mxSaT+cJ6iQZPbrS0IAzGW21xcXGFv7xdpI0wV28LtPA49HyCVtgI5ujN1v
Nq0qzHGmTT+/CaygBQHFkD2WYCbWt5I8msNgJKmc2Cu2AZhjkqbdvGI/6r/QukqS
zk9B5/ZUDdeZSLSr0dv2Qi352kgABXoIiytFp7xVjRtnBWRpsU3lszc+FE+5hpxV
afqBZA7PO6HYEw7riWOa3YBP/qkU1ERYJVGsfDQuu26gXKS8VJ2mPuGeVspUfJqw
1jfYLW8EgSD/v0G+njyYIujn33FOfLL+oAVf9SiIyyI9vPUTWeSb4nH87PVO15mx
13+YMi64M60Z8Kg/oH3wjmIuKKXwQn08SY45FzOb7sAmjtKrZdT77iKfYig/EPrJ
PdlETv8d/oPvJJ/OqUHENbn+L4P+ibFNF6C+wfO4E6gceLCnMiwaLQIwv/Fztdhz
YHkPU/zV8Ggd27eqor53f3hZ+tLPgRgwAxs+C9VZWtVVttgKN6QK0slzGLcG1qYG
szrRR5f+SqitrLdLv++dqWoP1rSQ/vfWGO/czqTgRI+8sB1fEF8iqlh+CuIxM1+v
X1m2BaVAlrG5zWhK3Woxh7V8fpZ5W3ClBv+Mk5geZEEpdbb7AKmdlbqyB+p2XOSe
ElMcqYKjwVewiZa65nQF6UAAJIbDNxF5E94MxZ9JphUKCxelVdASk5wtNme+7WVS
b6RmS29g4AepBmUks4Frkqr45Z6wz9hbgzBLCzCOUmmT4C5r1FHkUNgk7A/UfKiC
I4WXlQZgAQ70EALipkbEB0VsnoupLmaWm5T/Jgsj+UAnrGysaVp2DUzv5Tk/4uM0
UO40SeAqlsIAqXTnPereRqp83wKLx7vuuATMjWOnXTilh0tKFKmHKHO9Ie4CxZxU
Nm/jJwvKi3G2sfXj0hUW6ZveJopjx/0O1k0aqd466GWQSG9uggUS2JdNJ/3nwKGN
HRgq7VqzCT0d31bpyBdn6pz5r6WYMe29LnD6WqUqig12/KhLCQCdCP7RQa6Phku5
9p+73Dhk/NrqD/utm1XGcC3aWmK7URVM0ZF3JH7BY/tElSkZq4TIVFgzYUBqCbkF
UhQ3N6fLs9ZdCYgjckgZF1zzvinFzhMpLzHwnQadUWCwtrkCBeEpWpzEh472Qa4d
Cm+ztOrez+CmrbuW2FdfAY8HhP82Rehm5QeovwLmA+uS7v7GUr82R5so7qcIZwUV
PiGQyeCc4IkWgF91M6s5nntPrg2oFyKmXiY9Nt8p6kU68xqUC6f0glHOTvhrJd16
Ew2DajAUMzPqyiabX8n4OEVK0MFOO98kBiQqcV5DKb8PeZ7l4+sm2Z+JFO3I+grm
7eNLqfLguz2S5m+x98vzhCp5iQlNSfw9287VL8n4s1WyF/G9n7coPlIgx/9AAcW4
+jh4DYfSHr8O9YSpONdt6qf6WX5GNxuSsLL/7uioR0n1hIkOLMW4ctacHIS8TCAF
sxeBwSN6LwmZgfX9NePW9CHco5g6Ttp+3zfEX8tGnH2VAS9bFPnpolC4MmFbo9hz
rHUi8d7UYEmPsOSdfBl6BZMioW0tGzWUNUbZO9HTpiRnbzVEd1lRdlcY8mGi6gr+
B1gcuiLnscAZBSuVCed/BHnmjG2p6XjHV9Od+s49Ty4WP464SgnQhjEh99cOXJdr
MEKUplp/FUwOP9VB1GGaubq4Kk8ARHGJfxj3j7GzbO3zztU3jv2xlc4vZlTL1PM1
v9cfducHneD/hmzbcvCWf55waxnw0ZM8Qo+YHnr1W8GkAh11zaKrFx7vALJj2/Ps
/TneqwApSJdfAAadlVuzkhY5NtiaE0XIQY88pzbSgpnmvmQr7PY8hJcXBJt5yBSh
rClasoefpNKqclzqrTW9u3EhycwjcHiXXQSGzobESuHpkAXqcArkwksSwhAZBlry
k/vyz1osXUWUfPvyQiw1MmLRYGs6uiNMR9OKOsaxJ87/RONvcuNQU6X149j1RWmt
ysKdbuJJPlh9w6yJ5Ld1WH2kFvyV7P0xpEn1fqgOEs9mbPsJP84Y08rfeLnPefX8
GYlwOsK5l39OwMxbWCxUp2MKEj9agXGXQmKcQ9+8bEz1JrQISEBAKrW0ByedSg1z
5CH6whYzUmMNX5Bmav9WGI8dASFGiM1jeaY1vrGVgfSJF8EiLJ+8CzdoaKKvOY+a
K99TUgtJirpXXVY7dMmqPqk08LMqlXnpyG9z68Mlaten/AX0dc9f0ILcCMQYMry5
KjbYmhr2CMs80Jy6FXMfYVXkAG5bnuZBaXpQPXf3TAnKeQKWa9VIK39BAT6BDPCJ
imPrfn9yVCEcGLBPkjubt/h+ubEB18VLLqPBnfkCm+1VWDWFV3J/gMtyve97aqKA
I9K+kW5nqJ8cKmNCdcqUk9OaYnhHfzv1bzDuIo0hIzLI0H7vlxMe7w4M6xttkHT9
e1DSyIb7nvpmAEKM+gl0mlxmS3sF3cujOvCuqXwTOSk7LyKRG1jmpAKa0pWIdlXD
lhf9juBq+gpfHcDT5StLHfE6ahMaNx240F0MreK1SXceFbvdnnplac4kYwy+PEtD
KCS6BhZ3kQGNY+hm9w5cAjcZ5GdSQo7kOlPpGbv3xp4K0IyXzFYB52YPFK4vnWUE
Tbbd0gjUEWc85HM5VFTuWZMk/tcuQgswuDKzk8HePZQXLw0UqG9tvYna01x3+anF
T3WNfM5yWePJnNfz8UDBXjV/mVch1MQOvxKoOUUWgY4QLGaGVVnW92vwbN0Ip8SN
89+IV+tTqad3XljY/q4tY+kXYPGjCyoPUHKcAe/kytNwfuzLQtR+ZfRHDvYMZMDY
YURN783tCqcE4ejYRHhi464uLN9Aby7ptPzojqzFx8yh+5Z6kBG71WDn0TWXGcYC
lVjbmBbzUkQ94lGDsFewHJGmD1PtaeYYJVIzJPc7Gfmmz2bSAVUOGaACCyK++M9A
Iqtv9wQXseHALD0zGt2VQWRu1kHzLZAr0sQ7EE7DaSIrthMXTQJP7SeCEkDjxEwR
K8AMzLjDUmBR12UH9E6Gv/xqZnCQ9I+q3FC5YHzD/DGzKNbrw/+lfmuDItLJQj5H
0qszUZMW8xM+piyDq1aiOor+e5c6Ky46VqXqI2fkGOlgKwfAQ2ypI25dXz5tmGdX
huWYc+aI2GpebfbaYSQ3LzOBauRDv3GtFgnj0JptuM/aQ7Rns8RB8rEdRyBgith1
/uE6gQQBkpDAice22wbAYZMEx7zSxyIZ2jThiWCIRkFTowo+bcsODaxCZhQElK+5
0yzBl6oIiLw0HXVARaFSNFTgNjFPZWShcMePGOLaG5p4PSXyC1JRBDEqgfVj4mMo
8VmXzdAiuTmONJcc6iOF5Nj4BGPlqnTkYJhaK5GrrUePnE9QOTiTGd7TyTKTU1jA
BNLdsg8MnlGy1bSYNc9wUL5npJ+XZLRVYssWjO1wKsL05uwD1DQbgvi2x164c6ys
h5xTa6ecDwrGL5sUxDBMyVPjPU2JjA68Ld9j0xUxZ3fqFWGjOAh4LXLjKyaGgvnx
5pBF+6WwtyPLvi3vamUoRb22u+GLnmpCgpxOr0yhI2G2S9rKZwS/RsS69mZ9pX/E
3X2qL9D+UWcH8X7D9rWmz3DhSoI5cw7dRqeS75yUt2Wb1WRsHEK2aSLW3K2tqE8r
rZ081MD518GKUj003Ztvq+7piSouKWa8/3I3fVTi0uyIWGoYMOXPBzQRrDmLFNYb
3NXoHCrC2AGaTwgC7SMkbquOOr5J12huXcigX6UDKR9medKhZEe/cXbY/Odi+ArT
vejg+eLhCYattvEw+JS9H7ADYtPpVkiUKPiIIYIl616LciIFXtNXMpxygPyWX8aN
7j2j2/Bwkc8Qo1QjiSAawBtjGwA8XVdIGng6lK+/KKJ9xlMDu0D+OmVkp6MWOshw
btoYiHF53ciKsKaFeUEXUNd/gR7NPBF2lDg6KGEjnOuaPKoKOa72N3cyGM963aIn
oW2KkMw6xz3PCwO4aRmVH9xBxatIIsWIlxMFpzJ6F2SRsaLGQA50O5i75F/dFPuI
N5F8P0Jh8lfYYlKvDaPfpQ9BT8SWYfUX2Et/mxkeEr531JlFNbU2/Bwc0Qo+h0qo
1HUDaZ519roJ8x4AKQOXyqh767Dw5bS+VjaASxUF2KOCD9hsdy+IHIqfc81GcSc4
B3kiMhJww11hgfqJ/qW36YN+whKWwkERvj9EGas8asNquPp0YdiTDWSKb7ET2Gaf
FlCel1b05Lczf3f5Gs+fHqM95KVp3l4iglxHQXjUPcgkSPciqNVPDnHZiurDF/pb
Ps+9ARMBLBYKlPAa4+31LGEFS+GtcFN5tg+rv/0JzyhZdBQMVghLHwBJD6C8K3x/
GtoIBla243ZZ8bqmOu+Vya4IIkLF1hRtGyW/jy92nkHGCLqN7Kxfmxs5nLGESfbL
NUnHTT8M/3x8gk/7ReBYuM3w6hOn6YzOicFxi5BtVo5z+L+Vfmx6HDb8+31Xm7nI
53q+HdfwyNj3YNfdy4dS9f72lG0Vfof0SB6RRXdUAT9v3eTj3Vx3hxb1Em8gSLJo
jAB8kfWgZPMQ87cskf1GlK1qcIUyRXqy/6UbAhCsCajBYParyX/Hsr1KBYCcAeHR
quA5slO/Y/w+0/FS0gzziaLSH5wKqOITBWxd99gK3xBZz22ymVxeoodJWPn77QpR
ALJ6mtE+snpdiWvhGxxWTU3ZkUVzyET21bGGc9W0N6bTkeBpcjC+Wox8fuYRyDY6
ZG/7pbbV2AHPpM921wlxYzYDtG6Cb+/OZJQ99AAhRp4nfzTfU17qUHcC2IMgfJHd
GpGN88s//1ONhUQ3sp6XOLWdlLX26usdYZbaOXINpOcxM52+mb9LYW3quAEz/blT
Ul+hUJfT9UPaLPE+53/QIbMulZqL/kpqv3lj4JxzRDZmAuA0nIvZI9cThh0l92oa
0n9yReXChd4sqk/fubgmhjfjzfjfYZX6Gh/FrEAeJYWfLj7bwx4mGtkJ5mZrwZkw
n/trWRVUwZ9kYCFxYkV2oWgNecG+8Px7A+s26A5ljRiJYCUbiOeTYRAn3Vqo2Hnf
BExwfQgHgw0Ezst8cNB60QAIHwg+MD2e8Ukpbu5VNtSUCnAVRduzkbMS5MCZNt2m
bARlwmDJ0J5mNRRNWGs1IEFgOY+eCYPH23oueXrSoJqKBaUujPsJK7npOAjzcQ2N
mqePVFNESx6lPA9cuepxWBexzHs7lr8OiORhzuQ64Hke9N0iqA6G/xrUTSn9qaer
CoE7xvEECCUatcecQP8iENej+x6XNa67qMeBG5kBidrAZITS1NfZYDqXQHFZYj3i
CkjvnLCVxkkSzDV+Mbba9D8eJwmGKtX5Heb4oiN922jeh3WfWM6ita3qVDGaAlrc
lzfnChAFUGByq+hCfzpLmRMNpOJA/MPg/fBji9PtzF3kGOnBTa6lXzeTGP0B+4of
JSb00k4FBR3dxJzc7bIJLA56oASjEHQFPA7i076dGgjI4Vr5Lj6m1b0kuSOY/LM/
tpeuIYNsj/iJfNWgmvbo1ky/nzCFpth1uYZZ2U5VYXx35901LU2lb55UbkjD5ZNR
9eAEFTJJIC+g28t5zFDLoHGD2hOFZ9TcbZMteA+7E6IUCRhB4OPb17n2kNDyXhdG
ZEM+TAifkZPc8EsykW/krVq8/O5uwT5Uffrzd72XOn9m/MUOo9eYZbjHqcr3GsDT
itlojaSlD0KLpbySagT+pETf3zzB2rdQuxNzJRZbGgqfc1BmwhVmsXyUPNdT0gna
B9mDfQi+SvsXfwBLPP1CiXc7on2GVGy9Oaxdz56u+Wwr6W1615ZBqotNYSWt4IlT
0EeVCd6pFkwj4xFACRSj0gjSyEwEsNluFpTA9MF1GYbV61nZl9xuKzF/6eTom1td
RoEXlPj6/17zFSMqbbsgfcg7ojp0V/T2liaTAZ8PSlq+0+Clc7/TthIBXFsFrx3j
sekKhUmRWAXfaAbvl6rSydo7Q8OxmzWRCbYpsVBJSe2/LTuYbqJfkPBmL8W8QzWZ
YJzMyawpXPyLTVeDX9yCxfAyVYWqNt0AX9uAWTp7alMJmbBNPaEyeUpAc4IkIuFb
GB+rOL+sCodf7mYXeRrF81rFCpTQqvynr/0HmaD+q4f0AsJH0NQiGkVl+nNURjvA
cmg9r05ISHFDYn9CnTloUHhRvxWZNJ0W0XUU6HJ1wmXY7sbNjwvo1IeOV+kkyIGV
3xe0Jo7BIoAZ8p9COFkAAeC5ayYwULXH90PSHSn7f2pejLHHumauYQyIhwu7TOBY
hKCkuqaWHEadNupS9xW70UhHamO2VrtAjy9qktccRNOmJLlDWJUsWKT8CAjoF1+s
Il66aOqRsuQhCc9Lp/IN6czJY/B6pusLKV2QfJLa52YuK2vlPbcfGS3x74zoEpa8
jnHPJmFz+eUJapVDO67dC1DsPfqs2qUUQovP87infWT1SqWmyqLXQJgZQ2M0pNJ5
WhRIgAT87ByVwos5XYFlQHQ5ZdNc+9Lx0M1H8kmw3AnL106d6PeOrPuEy3vGs7Aa
qpbZ0qKawRn7ZurguMOOxyuQ3Hzg9mJ24lCUJmUv+4JHdwW7qPTksIFFdfJgT/4O
B2EXTeB/q/Yn3XBDq1Yq3Uhan23z1a+Q3M2ceZt76pEUx19DAItv3jimjoYfXnxj
18QWAItYgSMPlTMDKxH6a3Mimta2NbnyjKIVkxae3cXl4BOyrxFgMyV4C93jxDIC
OYdFeRebDsFKCPWG4baSmJMjgWQ6dlT8t9593IKlcst7w4RO41Uzq+hLx1Xc+aoC
k2QfofGwNhLk3YSNOeWKvFp09l4hhjZCf21kJ6Cf5HzGpi8hPWZpNYYKIAIoG0hw
QxeGy5T7dqn8PHD/o6V/JYZZwTnBsae6t4d3Ake9xflCCmjUaqCwCarjgAm1QXIl
fGkUMFgwf0M3fczBA9HMIKWI0FwFsmhMhNhELIFDQDM1GnjNXx8XN8UylbcmGamx
DBMfAjppRpVWtJ5SWkKO84v2Fi9FrVbogxleDzCXub05OENx6FCY0fSFYE6/b2Xz
CfINgzVP2CRVG2QrCA5kt0iEr2m864Ni2uTZigDWgsTM0T1pK+YXIiaiiye/a8Yf
Rxjx8UTwymbFWP134FmcSY6Uq12Kte42dG/H0fIGVYo6f14zdX/ZNGPPqjLlvUCJ
6pjcrpptKcSc9UtADdl8UcouRuR5+yiE1Wv+FOg8ROofz4v+Z6U8oUUH7Y9N1Shh
tSz6P68h/v8iIfxvXbWsPd42IGcbyDmLkDNd07XXt0YHRFHjP7CAsY4OihYdGjie
x1U30L22vemhWzRaMADkAy8fxNnDN3MWg+y51QupHmQhzylPVpUNEVBy5mN5hTn/
FJaiZf/aNRq82AAnwXqwjy4hPIR4SlVf+l2EelDZOrrsSXcRYb1Nx9gpU4KfpB4L
okcE2FGIweropEeu98vDqF/dkElO/9cFEvcxMLxBHvtcXPvBDlnPYSV+ceyNohNs
feFjsksAgFjkqrOjyuj5BaE1NTNBQC7z5Vr7e3OYu1De0CRPkowd4oRJ/tgb/pM3
3OgyDnLLix43UKxc5RssiTKwVzYGH8KGUc5tYB/cfWenhl/2mm6jJu6diS4OY1MY
lrVwId2hfAa9E6rc5/OLN9YKsMhp7KP0CCWclPEmZ3V0DPhse5YVW8kRd1uCXR3P
rzbYQmbRf9709sAi9JExyVE33z1gzXTUGUlhX6xNyx969ykUSlUfW0HBkXdPHqrW
UvvdtqIsJAV2aPAH9UPA0BrESb42fg+vXda2cGAD2xt2P0OEe4mbRc27TBcPy73g
2xS+jzc05tn67ZFzmdFinJ4OfATls5v1QywdTbNNsWNxfwipax2t7x0eMhfOALsL
ubosoSWMtP3QrX/NQTl0iedqQSP0RUh7K6hq711bhsi2KpgIB0BGf2EgeuL0+Lhj
vY5qO7U5EaUiYQTXGgMxNgjTLZsr8+LYe8vfpTGdNUGUuSxCscDFUP7Fth68gC/x
wxLS2eX4SbqG5MRvxeF+x/S4urt6P+EO4GRAoMRO/MghL4EYFxnmxKRL+duYL5uj
1M0rfqn6x+B91H8Cl8V3uff8mGw20OHzGStEFSaokT5Hv7uQ1udOHUWRJPWF1Iwt
1ksyQHB73DfyXwV/SE4qu88qATCaG3ol/3LkupuqWOGR26W9emPblIJNYyLmW1q5
lkTCK3PHnr+p6zoj9XKKtUPZkwiPLnXS0kg/HvJIxknQZKNO9bfZroKksP6ptL7X
KaNCPMq0xuN9L+M4+sNbYKnU+c1f5QkZSFlKlo93vguG3nQfSqRQThHsYuJ8oBr2
1LDEG1VCitTTfKCk7FnJJ6kU+dra8DkFOAb3DuvU0YMSzSf8m0aq9nSD1mEQIrEp
v/uAjvAteo5OVVohScBKL8QnuYhsniOIOau7WIYrZP5+wBEnDAGpp0ln2vA8waLU
z9NjDqbXd1Rbgz996udEH0fq+YE/YZEgizeNA5nDsC3PC5sUiETRUa+CfZfyMJJ9
QjhKHenenbt6LjVLL8T8fjXPJ/8lz8l0pqA59dYzi25Gmp+wY9x2RVyh7wDp2SrK
LFS32h3XjJg2F5U8200g/85kCvmlYVFiiGacqQn4Xhio0uS/AyYoGgCMaRzmyY5m
3LiyjvmUY8i8xDnqnjAIUWUpbKKea5slc3zkUHjVy0ljjChSY1J3KNuADCXKIzQi
wJzVnocxQYizLTgXj1xhSKNHGyZbwUk7YF3MGLhkbNr+hAZA18Mxrm1PPuv/JaOr
fVJ4beSRyQEfW3gGgWTBRqcZo6wu0Shl8Ffm3/cbUKfwLhzJcbngUpg/FrQosfRL
uDIM/M2oGk14PjljZtCgCjapvHBS/uT5xtkWXezaaWgaQ4EhMe6lvCtywhmKQByd
+pTTV6QPOuW7kVjUG6mEbLIpWSMGnn/3jqoJ5/AERGPsvM+JUjQjPE2mElkObZg/
AMAyfG+1i9zLHiloSpgg9bsOHcdS4suR4q5s5LSjUcRxi1VyGaFTFBZmZ6vhVudQ
3AwBm1qhuaZwD1Izbjm4/Cv2smMlhaH2ZK45guPkmJq4wehqkDpwXqJPmuI34hJm
8zATEap6cZw0dOmlq+rzqeL94hGjHJw6+bJ9Bdu+RtNfM08432S3WQQCa/uixYPH
b2tFUn+zynLRYTJcIA9FEKaJ2JutY86DmZGILmGn+pN0N+Uc+G0OJ16O3rVwnjBq
J4mXCnFJgfg3Lg6f4ZeNPejh1Xc1iOH7VOI/sbgiDMy9J07I97ZTi9fmdtH5KX4I
a3LX6nyvv96fUZMWnBXbFO4SavIHZrQdyegYAhHiCC0mr5ioFdfz8o/0FzOHPH6C
GqfUUHsgT5VRQw4ehlUTvYaeCNTV44hMK2EK5o1kerv+6DULOhnoymuaxmZimsWA
zAiJz9W4kjrw6YeAEt87b8MfXw+c/2I67g6mu/Bt3ge7QDtbFEbhhA87F/9IeDQO
+rjQVSbvNjC0nxYZOBPg+kmeAncqpqyfVGt6yYAFqEwzHvYt3IVEa/pcuM9AEGpe
srT+9N1s6RdESi7yW8hTrsgnJm1f6f5sRvq4kvYmcm6IAxEJtdoVXVdck/z3kH15
fWN7XnBD2lR9cSDl+vE2uC504dvXrJTxGHqIDm0DNUw8WigDXZf/Gy/lq6DMUC9R
F4u0vTWv9LXF+aM3Y9bquSgSYqoF5KOA+mYZOvSvrvW4j+mxZezMQr6kJD/ozZT+
eFl3ZZ3V3jAgNRLjveyzMMxP8b/uDtSmquc0RpWnt1nYgSX292yLxnoSLqB4bhcC
pLIPBR5GSBNqh+FlrU9ibK8KrhibowYg/o88nx8opNW6caXPbnjjhEY+Us3b2ZDj
NekWI/tf0MaBx1KN58rO/p/0d2vLjw+mfB5zwO8gIZu0k8+EoYS/CBIVWni+J4H8
yftqSQ/pOBLlUTLeK92ZJHbx6Ida+xg4XJL2xCN0TYHK+zO5gLpn5ybL0Vqu/QzT
/R88yHoNSztV0zcKWpGCd72eLtiWxXSwyEKdPiZh/7BbTJb+g6C5Qq7hRo2S425Z
WhhieP2tmbUS5NwtavgI/b+pzbTk1m+VyblXvhGq+tnpmpnEw2LFzB7VGdvMgbaL
mOpwGG8TaZWpRPdvP7+6TAbPd4fxso5u7EPN6FhivrJ6EBiFQwmDZa9HFU9vaapc
jbWs7ku8CFbq91VAQBSpmOkU/2Mzx75pK2IbJE4MlWJfR0Wd+3OQ/XPHhttVqTRX
KzDklUqsP3nC2ol87xzDKUfhdZoZqjLrzO+oLuugTP6thBez4cyYEIABEIMVxXZ1
4oQ/iGy4KA/pRSESSIN16P/ceXub6jyXAmCs1Wp4EuAHYI79Irsn5uBknCmPuuj7
odpJBjaaDFKTrGbAJb1LmpDfrukReXh7DhmJK550N0iBqT1FiPBKgYVidLRoUkGa
bXY1eTVSFf+8ODjnUpip4IoGYWNO9IqCUPFcnYwl636630xZ22wWzdtJVOlLXv4G
tjEhfKTBz3sIV9zaBhppMuKr3UObWrXy5BC+jS1zikEw0cINP+wy8ccpxxg8Yql0
7ZzRMc0L1A6KVQ9u1YF/OTZUfCXnx3RU9ll0aFSSOc5yRY3htLx2e9ODbX3cBioM
DhqIe0F/1AEEYRJmBfPHRXyLQTLhloMei3simi8bwu6T526cXuadC4a12+0c7Hkv
ASyfpoM+0xZW/vnv8vob5YvOiSh0jeIWvG/wWYt0xP1hlRLyFeX4MRwNZ6dE/7/U
aHYhraOaG8A1vlSmbJT3dU0cLrxvgoMiFh/ezLiXXlmSqminErTs2NOKKiI4hF9D
AKPu0QrA8x7aHyK7DftblMZMatRt2OgTtef46Iw+4aC5gx3XFqTnFVDik0g/MiG1
GbcNL5tEqPSU2NKRO6GfxPXBSWbSZ8DMeftM59p/qhMMwJUqI3mYS/4vCSjmCyQe
Kkit2iiPRBPk+yxaLuQKwJyUjjVLil6W/Txw6T7HxsblmMtFchuIeckhENbkKmlK
xYLKwXEjC8ONNpngAcI5r8n4U/mls7oRn5VO6+S2j5mhliCIMZwgcZg9ooveOSsj
FX3ZdvbFFJeph4Wc0WI9GzCXfoGA7aFvvteMUeDmw1G7VRTOILWi4sjYh/yPhDqK
nry4DttnF0H98TsT9tyORskbLkcasC5QfruSHMPC9wO957Fk6JORsvmEN13KKcCk
b7HK2X96SFtmq2avemfj1gScZVmESCzzKvrtFwzZT7XtwRbfwcyj/u8WiiPD7X9f
EOa2tpmjNS8d7o4Oi4/pNFALXMFSALEYl8QPYrppNCAZB4A1WfJrNrJMauizUG07
2q32kJ1INJd41wNTeB54ICQIJBLbgjxBbXZ2nJWMD/8bl3vgnOgOe88liyLByVcq
xcKGy8tVOqajk2eql2G3jjko7+tpcNc25f9QbFa2XoMbEO9aBPk5i0rag0EFniu8
RhWufQwKoxqDit0QkgCUVZ+b5QkrcZI4SVaqZh2IuzoUcxVEjPf2gctHGWx2V4T1
YB6slVV7TaNDMKZMJofSatTzXE51bXYBknzVh7501xIOfNG+hfWhJQE1uYJ+NyJy
ddCp98Ov/UM35gZqfJMDj9mzKmUmxJPewzkkjJ7jCYx+ZZdXxCLbZXHk86Q6J280
UrmlYBIASBbBG8KBKdVzLv9PtAZhmDMXova1+yWa7IPYWjugpjzLBbY6xMItHrRB
wo+YO19KKLoO9DZYnuCq245E006mV+lv46YhizzqR2CLo+btZyqSL4qpHO+ph1Qf
8YSDRY9csUBqyol1Rx27unYdVLIXh1a7bp4GmzCrYqMevlj+xpjjXKi0ObQQL5z4
mpR/DwkDSO0PG0H6kruVYdKLJoQB9kfgEhqAohkjtqhXGr9c+x4UQ500uuluyiCA
tMV0KCsmMrZMffRhh4Ebh9Fd7yTvRwOyQ2Hg9E4i5V9lI3qSDqUr+WJW2HA/xLq+
5RZ1+qQRMzPXdtQxSLDgF8giz5+Or/uzCggxo4+3eZ4HvsCIpTj6T2sIUT5Fj1YK
lPB3Enf6r/xIaJyBJtf/GWrgniDLZ8ZWV/exMs9PKHUWmKzjH4P4ICXio5dsCkgT
Iybo/VRkkCtwsIfk0hI6YfMrCWyBJau+tKFkeeEWjk4pWGSUbMUtbbX3rrpAphjV
ExpGLft6SYZjEFwdo4p9itvLh+nyMdZIyJEvB9BhtVXh4YPZnXXXacOAMQuv4JgK
oU/pMc5g6qAobUdLXtHbHfG+YghJ7/lVjVtNyZbqTw1r2oEWiZ6jU4gwRNSh+bKW
J90D9nIq244BVTSkAwSkjtcYePxZ2WYkO7xdjMpO6CNkzz1ONIBe7PYXNtjj53Fe
M+YqTSdyKq705JWc81fdVrRX0i8XCizeec72tuh1IG5GeSdUA8m2i/zI/akKWiOW
pwP1DIIJqaSOqV8GcJ4qXJlRA0Erfa09vg27iL4VD+euR1WLYa7DPnSJpCxiQ9TT
/ViL3ZbC+l8xjCda1WwFrVpZSkA0mb6bRy+gROcbr/Rncrrz7szBn6Vz9GD2+wxS
XOD+NJfksQqKomjNasnKaRxt4O/545STaf6DTdIWESSQNwj21/c0r5zxKmi3L+HJ
iqNGMHoiyzt7wEy26NyCnuz+08im6Zr7vqbcRcQFQyBXx1/sn0mKrd+g1URzqejP
ygP7oqhTBGhoO/q31Yj54mLhXews4J/XXEicCwmvuX0Ha+QrZDriRU4GUSMhKOUC
BWX3uRSO+eNF52rvv16NMsq4PuL+zzSp7mwQ58lMjCIaJdCrFvsrBzq8S60Po16Y
TtrrMIeCSqiMtzwE/3H3d4bfwACQ+a6lt/yVXkTPu3L1E0N2fXQEbU7fBq4M4HZs
cgfqS2S4GRGRftYGE/iigVwNNjt1x/DYleFpd7Nnrz6jpAQTSUS7Rpr6KrTN+tGL
z4b7mf9A45ne0QaG+od3KibipWOHTAkuZEx7UWOV1QTcglKOYB24fg9mFvG9uuIy
Qv+2PCxypyDGp1M6iwtJSVUQXpXxIOkmqxWYK3dvJv1KQAUShhYa4rQRGgtvOH5K
9dzPsTuDoxTHCsifhfTT5/9Ufzr4M4jVKa7nELCwYCjqYGhQyUgll/QnMc0I9yqC
83JD2n7O9lXHk3wzX23K8eDxLDTZoffD7wSGf5dUvSg7RbcVJCiqkz8q1oUb6142
5iqhQPCwdDSDwl/j4RJK+KaGpLG55QgotQQNp6oIdgBeeJNbMhWC6blfgSw+j/JW
nWOJTSjYNtJ/eMkWvSnb2jMoE3WuDTf5UZf3+StwNFV8TGOLzY9fIlv2kg9sQJdy
mKIOcF+xNVZlGLWcg0PfceTw04txQ4Vm1/FuoJgy38lHO586XnvRd5xQQWUdwYqP
HB6DuG1kQHfuT/syihZVQXQ2/o781zy3Jaty1eruBNesgbKqHLzpz40G0Uq7Z6Yz
hhjuGMBg3np98aX3N0bE+o23udin8Fo7Aaz20DbstDCFQbfbpXqQbKBQo0wzbTIz
oDWzzmiio+QLpzwU5IZx04wYu5snOeFDy1MfS9OJbPCRpxYzRJZHP9IwYoN3XVWH
PSyI2NScBjq4vo1nvKr0Bao70nKIdh9s5RR5MO/5z+kiTTQE3EYCv+q2d0BhcFNl
AlX9gFjfJFxwRRpbjv6RwCwp5HgbkXbcDjJGfLTC+eDB3/W1t5WwNI5ht/Y54s4s
/VEfpmKkn89fbshw0wMnS46k/eQZiG2hKLZdWDEyrL+v3M/ryOie/JZGGjs0D9Tr
NRmnBPgRqXs5SPAFFDQhX61qDegVUCXi27LHSxQXRStlY8LnEDeU7hThW+T3QJmo
z2Daiu71I5ROl1jozRjtbTzd3WMzsTWcxYDDz0h6oEkzwThQckEig/F6omvK0cGg
rjRVFHkKf58oKD7mr9FS5C3IEW64IHdQq1qrB9uqmOAQhQ3KctZccFPqHGwIJbdq
kckUXdqP+vVlj9wLRgkovfP9Cm3jhJ46d1saUAmzxAjYTdcCCAWa4nofh6T3Z8Aj
HWECB4bUcsMl87vqXVRNbfTMHnATudTCVONJlt5ro6T0eCXK6zREPgn7L5n0esAZ
digaXLEDQHeqWb8Yvrz+Y5oiUDiogWjTXoVZYBFM8zTBHK6MHBaBHg/Ueu4VtKJ8
qaGg5C5o+MKL1M4PetW05gBvfYq/m9KJmrYzfujYPIjHYGtXnaLLjoLc7pxxlvQj
d5jbFcmaX5C7Q3tIFgv0yr9HFiNxfk5gHjSoJiR1XROnDS0iQH4qqxw9RIOO3PWw
7F6UHZX3IF/4E+1+1K+yYuFiF236CoB6/8UZNXLulqkV5e/fbRlI2ZErNqfAilrw
foPmH1w7DcSFFaVaJM8srFjbbn9jmv50a2xG+FTQyHwU4NzUcCvAfjlopaMGX0Ca
bjurR1etTMANH+4RZMMx3wse3ORZmFyOVGcYYGhzfXDEP2EaDEMQ5B1O+Mh7rzkW
JIWy1QuHKDLW0ufrmBa8+PQKeAZWDjxJ2cs46zySea2/Z7Dh/FZK5ep4pqfhrBfV
nubV6Zmcw+v0467mH+4up4rQoyxVSE3gKxblR9fQhLBgu6xVUPqfJkxoDeoFFw/T
PXks5KiR7ra9DAliUNMk3pyE5imDF17DZ3eJuoDrMsns+9gX2ePqCvPBoO0Yfvm8
aDFoBgUsV8wMjgXyD2icwNDuIYbMD6Ml6T7CQJevGQC8uzsQD3eWfFbI7w+AxB51
8kKT2mf0l/bNAMrG/FpAiGb1hw6/VPJamP1OzWu9VkML3CkTmo1wFZj4ybb0pbOq
NYxCJ1gjheMkWfKMcSNyZ8OyRnIL8rG6XV71rrKhCa/UoqxHMXqSUzPSVAoSIP7B
Y3VINMMIEW5NUBliYO/5k9Bm6l5oo3oC58UC0EiAsj4x6yGoBfTHjmFr6LJGRpsP
OrKKhFrZzpq9l7tEliQbgvx5sHGypxwemLL0vwLTGao/w3cWYpxMxozF+UfnPZB9
GZ+H5luGgU+NwPEuU6YJ9KSVGKF+//5u01SRU/72q5M5DXCpZO2pOXSQ1TO90FSO
P/HCHEjmlumKMchGE9fNj/c3iPxjaqhyO2cKDHVNu7FRdrnL2ZQQ9FJ+lUs7mA2o
9PdpGn3XgvsSjg/KCGmLsw6XGKV8Hfgtx8UuD2d2JxAjnE5SVxy91qRwT9/312zX
5VvnmT940c1RPUde3sJ0DM45P7w/DuX2tujT+41zRiA8we3auh+GxaTlhEJ0EDTj
bzHwcZwu3I2M02Z/Z+cfncQ1dGCKNUcOWs0pUYWUpGK4xZHIRFRNaEZP8Z3Xym8T
hAnapHJ1rQvAhUJZU5W5Qvx5/CI7yhu6PsCyR3z9tU1JWwP+EbU1IzJoXj2biCKW
p32Aj/ItEveUiwkz3vL0Qi2U+CRan1WKLYX/uNtWRXcumXn4f2hwKCDrqgDH5viw
COGlGYTGo6+Q/+4CzKq+tg+/3Rt3B59tJUJRnXYattZhAA2bUKjT7/XRJllciN6w
eSp/B7ZfLSkwVb8Mbf36lpPC9Ru2Jyp1LREbzqF43nWF4x2bVHebQaZ5SFqaFMyl
65s8C4ofRPdHY5IOEFZ2oOkUcHRInsbdaZ6IYLKoEI9omqemNfu0X7yW7dwshWuc
Jlxc+/xwhWNq5RpIQwOrTIvhWYTOkjbE2tb8//h+ocTawuFWhw22mT3bZXZJDlkM
HViDwUscepbLvY+OqJtOSjn1gc7aGXq4rr38+JCUNxQzwq9ysO9FVWwKxGxbRrb2
tNHMs6uN8p1lig85Fa8VqcUwj9MkU9cqLPHgOkov++Xz2lMQcYHNNfciPXQN5TSZ
X7UXaKrYBJlNO6GE5fEk57gTylKg7Lklko53zgVJNnRbbtebU7Ad4Vs9jVvNdp1T
zTQYVABIHfit7qgFhEijidlM9/7iSLbWGVt+uOLN+03CUiMIryT6RHULrI79eRfS
0fytBCwfbkkF3wliJtJU/ySS+qsn0RyPWI3JUfzsFHCQKNibsXaCATa3Fkk6uUUq
EyVAa1iyWtpBiGMhW3qaMQFWFMJAY5rQrT3K+YMBu+dpFMNCwrwHM8slSDZClai0
Zm818FM7RtfObY7hUn0pmCvh+kJuiwshN581wl2gklVAtjwJbStFjmwbPG4UfIcL
h2blHNYV4eegA+ozssckfrAEG0WNWeq1DBRsb3lQFrGJqQb65ZmHv6flSnr1pRXV
vWf9NND4lD8jdvMgqvbGBCqxqhQr0vrPQ+9HcM0YXkMd96tLkN51hL+pQqb33l6m
xoFeVo2XIjPotuodli4klO7vxYBRPjwCZ7Wl2BOq/2FUDrH9dNZ0TeukEkgJnhWk
fVJTcQpTyJ2pfQxo1dV4aLPevewiUtCTN+GfIOg31skmF985m3SKciTCOO95Qtnq
D7SxEbK6C8aCaK6F8kmhxZbcSfFxOiBa+MiTxQQhNvhBVm2PpdCzw7AJoZK1T/R6
rzIfO1QQXAVO60r8cimMYw24BTf2cw7S7Uez1oJejfCQ6JPz07ys1qKiwHGQH0qp
Ej9y7Ekx/FgebGwNqeL2asUFZkG6ZU/hPRU9yzq6S2eW+d94u4LLtwctiw5prQSF
26wsjLpc0c1VXXULc/Nh5Oz4cB183sBldq3NR+OrHl0Nmp3Vg8T9liADD1nOd45b
6gu2o6QGe/cIA9sR+ze3TZREzn1vGqJsfdndwahAP8YTaC3SKr8rOL/AkLJlxIMu
YtZDshGzJDXtxbkVmUXxPydZUONj5HExcuFyocEyLGBLvOMl1a+fEvphN2dVEdVf
inZMXBBd9RriNC98IJHW1gN3A+fvpbjEDhHKv6lATTpMd9pS1UJZXEiqP9elhIJ5
QyGRCR9IGn6NchtG90wCjuqSezYjy+zTGxuU4rYGEQrJTkuxVPI5tW0/YWDz5ezU
HX2NK9BoMCpV6Mq/7eJipCQmZY1dn3tER9QJ/nvOrDfqLYAupLOZ8r4nTTn1tVy/
0fAeevjRbFOFi7cNxn1FoBmt6FI3S1cWCNNvAp1oY0Y7sAZfxlbV/754lbtewe39
OCmWVzGh6rMsEOfhsMGNGbF00n2NikJzrYLQh8sFL6biA0WXtXZ8tLpkFEFt8yU/
odBejvcVqmanHa7gd9aXepfO2uX+QO3DIT1sWGfvYGPvY08UwciA7M87kKFwpzOb
m5QIEODOvgJIXkZDKKwe+YkGES9YthmP9rwdhs3qXZAnb2jtL7QTK0GwuESd0F2G
vrokrx5QoILX7B8Hf+3k7cdjT3DfIP4qkMYDtJuGDD3aUmJQfZV/e/hBCSPdU0HV
R6I7/Fq4O8ojaZyTnBoBU6t8mgjs+/TPP0i8kui2fLJxXsVSGulaTwlBUaMSGGZ6
5O0H669mfiTV56a7hmONgiV5uYOURZhK3UET+KSdp+9vZ5SL4jOm6lEjRq9/6r07
3+HXvGZMs6++tWPydLTvuadBXENnv+gJYjCFxxPjFHCeL6Jeb7RH0bTla2YhakmH
jYA9QicQgXF7l+fk2aZuFyfdpB2v3eFEFayonRs2ohDol9QzihCtriYt+4xOn9sc
rbw80FdNEIPjKRPf84GgF9i89beJegWKkTPuooR8R4/A3zP39QkyXaJ3kVpKcmCN
BuZVi0WHvYB2VJJ9en9aLZ3YwcsCO2IwOxEdxO3nfjx0tyR9AezInNBKbvagMHTr
p7lIigZTcczi6JjlbUOBFdWqtS6Dqw2oxN3Kui5vQ7UjBCtXo6an3FH0QDtYaumU
00JX0AD1m649CB9cQpiB7LD8qYIijP2wKQyEWLGFtK9mNRq1KwBSBsE/b1kZarUn
RLNscR989wAAybOrY3m1MBo6FIA62SHWvIBfwG/8/Jb1secmSanlFpygowSXh4Ro
0rL/DoQAd5A17wBVDgu8WyJnCkzk4wF3f47yxeDrq4OZsIvKxnX+8bFZEBipZDOF
ywfQmKNBtDtiMT+QO26J5BleR6zJLaIFxV06+NdWckPZ36rKIanzIGzHNdlcDr4R
oaD+YIBdeJscUn7OFsRa7yS58amuhctTQHh15xK9ggSNzLz2eYlEgnktPAijvg/I
02vfpoCmw0y2EapNI6X4M71kK4wm65znIDaHMvuqmIZIrQdk3n/QN1snLIqWT9nC
Wa+xC6B1xRnW7QX4ch18MzDecDJsG+eVIR+8Cn2ke1DFfNtSWP8EzY47fiw9+EUm
LT1zGh+3OhZGEhlW6x4JmDwv4nXW2ea2NkJQrpkJc3+TX/hx2VXyoxLespS3ixLI
BD7Lh4vInx+vZd0s2cgL/AWx8rSUBo70sqWvR814y7kg/lh/V6WJXvGaz9hViY1a
mBVO+wI3WG1Id0yN+zB/sywMT6WFdZFy/HEpKqMmQ/z6d1AdaWktp8O4HsEhJ7Qa
WZi3iltfJN8Jo2XOshu5owyrjmADbNo02sm81SWW7Lm6IHRusZyhdaxNEFcBcMOn
L0zKXMjFirUY1863e6MjtKtcXQCyh/982kPCkmGS8isG92g5inpT5ddOcC/gUaQw
OHNqtobyLqmqEzXCYFj2d7sKitPOKLRr50JkhkMvnhy7jtf8qACHFzCflfbtkVOP
yspMogLET70PjevjJ8Cd3TCXuX8uUGaBC4EaKjDSg4HkXeHtorexH5Gr86Hvyi07
cFpKf1sfOgloP44KEOSEzlYoG0X7VrQqZ4Oykq4AH5EwNEHvyd6B/xnH0BJVQ+jQ
0+il2zsKZsALxmtCoxcQ2/WZq2N+kCo3TXP8e/3G7m6Nau5NnUiUk0AXXBBHLd73
k/XKsA0oqsanD8j8XwMIuyQBERqxxvEnRQzwfOkF27pHOEnzQoJ48+k20jfhiStX
QdGq40HoULPJatFVrvfqNLftuTt30M6JcmZX0de8sAfL48FNRKFOYLwKMTtNoKak
FD0tHbvazDGQiBAINP5DTSB35FQgiME/sBI6bTAWycUJw+3CuBPU0DL5Mmh+YHOk
MnVjARAGpO5brY+OP1YYc5cvyjvPYKWYScDUpr2uQg1wxj+OSB7/AeAw/QSp0Ewo
5rqafNDs59ITgyGoOX4m4g+HdAYlf53IcYYqzNR/tjXFNf3haYMqQegHAUJdMka1
o4Qb4o/tMyYYRbwMxQ4ecpzcsxGkOJ/8xhenmWVC8jSxS71zXlDLidw2XVqNjgkH
rZ3qBis8+kEv3VA0/hAufoYeqDIKcvgLRcTeIwK11bO+qXNZD1JddkpmzBT8kTNe
l60DBqxTEg/mu4/cMvvnstJG7lH666ljoG+tT7Sd4b6eilfi1FNk8AII/uvDOr4o
Goq9zUjbjsekxzobJSVewK9YWXw+BYIeYTzaF1RUV/iCyyyQhc5h9bqcvHqy/2Z8
OVhaCghAiGV7x+BgU5HvHIpxn6OuP4EXcsQCJo0ZXPF+XrSD1U0Fas3nUUbzRj2i
RS3dlEMmkRQKDopBEq3EXFfS8tC8stOH4+p0D8m8diEzlKPzaVDRMYxI5CysNzqN
ymlgr28NESCoDE3y4fjFCMVG89Uy4plat9qVzBIP+ZxBfwh2gobtkTjqg4nUxNCb
x+2D+OBd2cUHEDeCM9VdlRa55M8ynfNjK+S87yvKeYGXttuCfWzky9znRmOjMD+h
ZE0QC4WFLxlf+1qmBXLG0Y2BWFU0b+LiT3jvBlgJaZ7g09IabDIH2jooWkWkRq7V
8BT/0FCOjbeobbmLFKe7aBmFVHYQXmG7WufmaF3DIS1NndEhpVOaxjUWAfbCwIo1
3SZPwa6rWAepAHfPGyEzOWUxmYucerV6xLTfsOdM7rng/X1rxsnB1NTlo0ZFwM1O
3wVu14jFTEKl6SqWswxaqgqTnPxDjWo3BKA0hgUJhdJiAruZSY6mvYEJwzkaZh7S
u0fOAzZWzxdAl325QzV/fJ9/Fs5p6noONo8iiiMhDXWAiul1Qe3D0EwkrTcHGnFX
lpoI9VV7xGHq4rgcOVNAGneCANQPQ0XsmKVSNawP03q1yXe8E7FXdH9IMwXCnqsa
oObGJQq+QbbpMMkQ77RS6VMimmy4EvFweZiHJu5Ijnt2OlnZA1AaaxQDA29xNf4e
ZRNDlG4GMleXg8wsPuOQVa2XOASpRVA4jfvV6EUkCS2AidR9DvnNflFrhMBT1Ghs
LF2kT2aoC3ucxuh2Q6U/cDjw4rAEvO5bSMjiywvcwtuVoPkZcDgf9VrPx54bT0t5
nJYGwZkimaWsYyNg3SQfK8rr5mvcZ4PYWbK5lckRKhfg3a5mun4rg2Xp7U+Q4K1w
Nqrhi4Pva/+xy4bVrBHVPTZZl9RvtcAPyEatsePGvpXD0CMGceory0lYnUzfwxnO
Y4yNhrPkvkB62vN6zG4IJwhltLnntkZMLqsK7ShAJ15xtGwTNIojmGpWIkvWDFpc
WSPTJwXay9xuit3o0r+PmLcSQleZUybTjrhBfjkjAJ8vxO5laVtbC185/vq+w0Px
u83taWdivoyfV5B5T59Q7BM6U5vWqKnmdM7GVlnJEy0MU+S6wapp8lXLgeTGtWTg
dLlaTtpXzEnjF9cYYJr8pTMpkX4WXhwsC9pYwywCU0mFk1r0cIfdXUurGcnjFfDs
bSgKR93UrvmCAV4N44LhgaqodGUfB81a03RIhmrLOFodTrnQ7y2eLDFrqlKJaR7o
qjl9d2Z8JwH9naaLyKjiO/KQRaT4EdfsfwGNexvboBMJv24w/D/VaqgfbAUL8jXb
fog1D8qQYWuQZUc9miSQ7llQjOwK8BTdNYhNU2xFc9LJcst/5y71mIEAMyS4uKlH
7G5hALgmQwGKMy07BQXtyqw6O6AaHws+a8uWlWhOyu0hD0pZWj8LlY82cXn7iXYq
LrjGEnEKzsxdu7qEgwkmAUz8YHX6sk1EuAm2CBPUGqH965kPW+iG+ny2OJ8UL/r8
II+SZLZpDSnD1QtQgYpK8DZwAEs4nJtn8MsMR/NUKis34FEOUEYtzInGzaTUiKjt
STxrJ8hb1WpexgzXzg028ALAde18J5RtJXTfffHZsWHYz9qQTEAhfN/csKNYjgx+
qIQ02YaIeAawMwgPfarSk/uQqF4cGEzDbRlqcKGXde3boAVTEdfavX5Uh6z0xnpj
8HY+ODxMZCNvjtazGBOr4CEMqKuxi8UOXvVZ1ufD61E3zz9nsTVArcIjlrDZu+Pz
A8XTLlRnvCv5xy7cH3u5II0Exb9pdJF1sWsQ8a59pySaEhI391SumtJsY9XF8G9Y
EobSiiGFlSugL5wWTEcU1p6hidjYNNK3UGM0b8grE+9532lN/z1PGu7rOTJbkTYz
uwj2RcEehQlBPbDTHP91/t5NoeT1c5QjQ9AuGmEZGaHHVEkwPLZRWcbFpMjcjOTb
RIQtMW01eWlbNKbTRmGFe0XXb0glDWAEcuMWPWPY1k9HTGoL5JLFddzBdnIm+vD4
FOZR3CkQd3gQuJIjVQgfAvLKCKQgj+aqcKK8bIU0cx32yBnsnYkqTR90IeCmKfzp
KuUsyUC8kC/jkQKiV/+PyjUJrv50WSdSEE0rtuJtyqDWIt1xn6szupcAAhgvh7Wj
uN4zb5Q78jwIRUHE2p4kEgvHi9gEbYUXpYAmMlp3bsSBYu2//MuRxTsoQuWmU/l/
zs5qhHrnRg9p2UTppj2KPYZNpxAjVBc7fmQ8aACCzEz8aEL1PSobkkyHKLMGWWRB
JjwxvhQxDS/qcwxnFqQ6+ltUVuHBriiFiPw8T9LsJDRIGDRHHtpzPI0rydo4YL9C
ud0nA5d0Fq9I2RmVKPhS2oL/HX6eLpfKG8OUz8vsa0wAvQuebOR1slg9fsC3/eoU
dFEizU4qFXVQxk4LbmU4jv/fM3qXdM3Zj0Ki/oKsm/1IOg6ahNk6pnEjIxpqZnYC
nY1FwZ/0iSeW/GIdoMxIz8aw3W9fVSS3hQgHhx+2SUCKoNLqvDsOErtwwh3cNqTy
3fXCllrc2M87cRM2mdRoEiXumH9T1QZjZWTmpW3UdnyVZe4XoGTVJXUo2gFToaGP
xCpDF1HGICexIvNtVW3D2SgmbN/Gq7oyok1B1WF8xK7DQN3TYEpbwrUQTxf1UVvU
5VRVWspHgFEGx/qgJegClZp2kJeyXbfuh+8SHbOEh6djb0bwZEp1NTYlTxUQNG9P
gHizGJMOsaVVxJQW8dNVHFIYchQkAUxiMxmCAL8DMgOXEam4FccLyUfEZ49Vaj2v
uIyFTjnSvNfs656pDUCZehSarg0VaOO1pd1heaTG8+5RMi4ZbaoXpRfKAwItlmtL
RMVtmfUgA6c+5B7mjRoFvg4DQa4y5Iap3ZrFwJVid4x3MIYsxuNObu/FG/aGb0uz
nIwrLBb1zHfPQAEcfFw8YBKkFE/XmmmO4NjphoHe+BQ0GqYCM2W/IyxHWbOfAo35
E3opAOWHbssp6v5YhCpmr/dOsOMkPnLJJAdwfUmiDex6ULZ/Jy5mmMk+/Ow565Sr
IX5fSRJGt5QWkOZ49NbVeKOp6zaXisr5y1FosNB1F1pRnT4oNWORcBhgAu1ahXEu
U7Q/UvDfp48TZ6Uye59Y6aiuZ5UUSw4UNqSdJ0rax5wCAwxGDrg+B186gV7GdXBO
SPG0CgQjL8ad7GLl1EQE6GUH7C0oYg52jpLR/IBfkB1YqDOzqLTfm9mthQcbxMjm
n/4RHHtZTqdCwTG+W0luSB7WA3RZzByXg3ogh7sj8l+lnbnL4sLLw1WNKeUtGk1S
8Cj8Fi8YEGiummQ/ZtY7bx+zN5OnxUT3eEiuWgnw/Mo2pW7aOgFb1X2wKoVy2HQP
4wa9Wppv6eutX36najI4lktVcQpd221MeIyrbogq7N8+73RlW8bZE7aeZ/qhB4co
v/XTFKD7Www+qW0Zn4LunC4+fQJ9DOXxG1BKd7WF4Pc3pk+FTRnxb9T1RdR1lTwh
+Yo3dHIiLs/M1aL7b8TF9foNJedLkZwDwqTV1BcjK82A42CM1cvm0qrRxDgeDqCE
VDyUuI9vOmZY9XtHv4eNU7csViSgmqCG9NshZg51Z+ZMwP5kEkTzFDTuZfr05y8i
e3nnDMFoKlNJzhVSpCxG2scTp8ElOTBUkRI2nRwTD/M/rlFMxHRnMYUo6pzjGaDJ
wPoR52DxQGgY5gT0eTvslCVqZHhTuVCPbsMaHZxVE+ugPDwukwN3wT/83cAXTVxB
j7IiEqZC0c/pFD47zvanI7XfQqNkVZPtkdVATwpPG+/VM90vYjM1IePkFP0/U32/
2vqE+CnLYkLv1VEtHYJ/9C4xbBe/BrQueT7+khUzspVdgm6+N42QLnEtlKUZsyfp
BWbu8xgkCeMXULCvjZJK22Td8qpjdhMd/byTVqn2c7C2OTgw5sP/mBbDowUQdqCD
fTeLoLAYB4M4AFBSzzl0VHqMeYEBshwBcUM1U/9K2kcmhpIQ3es/wpzShswYjL2a
NpjKfDXxFUntEGePVkRobtIBlQvAe0IR3bM3xs9p8V0FX6p/WKS8SapmeK+wECRO
Afr7GSTv/hoDxtn0c+xMaFEsLzk7Tj5ANDa21yjZ8cwFwNPyOUnKvzKHAEBLvvIN
U+uAm3/6Zo9D82xvBIQ+qcBegB43dxSDkgLKL1U/2iT1E7pdecxXerAqtnAXvqhT
R4Y0eXQo+jptRLA9+y3MR3Km1wsNnjwtSE894IZzzuKcTEeSbaPIa2gp1xSLHsLr
mRl4t7hNprzVikpsPQL4E5gXFmBGJkinKn0BTsnWoWEXM/EqlpgxU1bu8cjw7Xfb
yNb/Z/Dj/oQhn7I0MV7O9B35tSdw+t4q8Sys5X8ZD2ZDu/0MwdE6y9tQNE9FhyU0
WRWVuyFC/CtsgyRe5LzNrCTAuxxIkxuA2lQi4Dxo0qkzqe55cxUWOiRhJrdBkz3S
q6oob1EEHB6eW/NIp5bBuN5vug8HdAmyfkBgp8hWJGbEx/oe7gBr39/cBcM2pxRJ
3g12/4Uw064Y8E3WG8jpXPBrRr2iaVczIHA/4bA9FeAgOwFOgdzNeGl4Cwat65Br
h6lSl0CxGyB7lxnGTM6TsLh/6XCXcHX+CRaCRbwkWeDzW9EABzay50HBZvnFT8Rj
cf6rtC8RR+BptpWFYIiBjqYtuAkub6mFUB7B27otyFb5JRFX0iZlZNofpZLRlbIw
VCBvcfomJQ8yPTkPZoKbzXY1my3MuZbXWCrir4UzzeJv+6B8TGm48QAEHvsmegD+
1zEMhWlHhg6QNev9IRlMNHDKzgBUzH3rxJ5pP9sO+WCNkinXXbNCAG8Kc6LSAn+I
Jsl4KeQyqQOdd01FAhuzBq1SU3QR+P2Scpp/rTUbZUyXaYlnAV7jdADlBpu441n2
W/rYl+rUW4a+AX7R+TmhApFox406C2iwN1Dr5W+g5WYOmtKuAZrCLBushwmJPKXS
fZTSPlRBnkfx8ndw/eqHs/VjggEY0XosXO+KF3QOpl/z9vOZ7IabVAUZ+vnJRx+K
nDRhSVs/p7XbBBufjuG8sYkptNp3JAicZQ0uLjHSD+cJ6FAZtyns6UPH+MFdxmDi
03Ngwm5ikRIRmWBsi11foyRCE1PB0sxR/LcIFaQGLyRNUHdHmAb2eHKMkIG1CQmR
8ZqAgtYYUx2Pjqimykz/VjSxPgUigxqBxSCLEL0BNGSjjqX4J/fKfxy/yaf5qvpz
cgsqWAGObNvwY2N3gqdlrb1bsIBcR722Z1cAXjjiINoNJy//8NH/zY5ky+K1+DjY
otCKtQ25IyklufVHiIYcDCWHs2duZxP3/x8Axow1XgnXjfftbqaLLenervDReRLm
p0m3CwBJAJ+FLmwyfX7l+rCLeaMQFlFZ50ar86dGuozs1oZQCfWSyCujPl+wYec7
yLZyPwNz7yMIo5uPsl+kJVRhd8G1j8nMK+6QSIrY8rMJb1/ebHh/3jKBIyWFH2Kb
F8e49IOxGkV4ySZ6R/jo/4uMSS8kSlSmvqwW1F5jcQR2uL7FdEHooQxhcRO6ty+c
GEHPXjReoF5HSXsleIbOdJGEwci6Ek8+dSVooy/W+mp3Jxr/PQ2Ci04F8POjp5Ef
k0WAXUAALy/HSYX4oovbsMgtXbGcR5EDBoJ7byHkSlfYpWMm8PJ6OSLBVLH0gHcV
ySw/s09TN2T8NtKCVi/Ktg0JA74tyQzJc3EkN6mVvj7UWd6T+SdGCCUbpaQ3/g5i
fFW87LX29p16u9/Bue4l2OrJEFrjyU5hiIHIwQJ6B6qOWOPDJXC2aKxEMJbx+lwI
ED8n8CqSRSjdFDnb5x/LUDgguQ7L+bav6XVVvuzdgI77wSqSbAvk8kjbIGnn9KYA
jGJw1yUAmiG2MMATOiQxlxTbxYNeLFA7LIBEcIEMpwokywet0wRfCZ3RINs336B3
w67jtw9nGgECfWfhg1BdUQ0pxpxOVJJ+ElG312y3qhySH1gZMGZADiq9Ci8P932x
M6wjmPUCO99DsVxD7ZD07JUvAZiYiMak+4nN4+rn1vxffAiC9WPHo9DkUPqkd3iO
P98ZiHz10cEPVgLOKYB45Gk8CvroXXoJiBPXHWJxhk0I9f05CiOnYagRPCDmMklp
LB1Xc+mhg2jWpgSOzyeo3WU2L27wuOhBNlUBr4xcW6sZusHDn0L3IUKxcX7Fvwa0
g2xPQ4a8eFQ/GTWjgKeiJPtmeDet4h+llaKC88alqPn08puyEeNnBGxikF8vOUtE
LyFyJNLiKErbPyi2OKEpir03n7UmJX5wBjUWFfE2kKGf3MpTOcKjCvInLcO5f9WO
ih0P1tfZzSe8jirDeg5N9P2U9jJaKQye6D9sgKHYtCMBmsOd9y/rFSdidqZunOKQ
fcu/BBscCRcmatIfWOVLtUNcSMUvZ+pZFpPYa6de1/z8zmTio0P7QZZ1qUI8XHrQ
saWk2EOGamBN0ZehroCrEpeDVB3BFOZWzaSBy97h1GyUX0hEp1UOUsuDZzJ0rrDX
FMRiTbFTaAjrVgGjv6fmzO9HAUvn/vDzdETecRmJ5rZi+XM170J2b/+aqUJUIsDK
e/G7pdhH8Cxt7q4SMLgWuqsFpOXojOs+tK+faTw+p1AIixw+lE2mEL2SyP6WSqzT
mHGG2qWUy5D6BK9VkZmgc/pYL5XvJ/3xzGSAamvX6GZvgef5/TvJrHfCV+oO76tV
SJiXOSM/KKEXQKgIxY+NBpcP9Q1OdA8h5xCesq+1sMZcoGAFv4/M20KHMA0ezEYO
fqXc2AKj3+/mkUWPxAHtqgfcQjAUO3C5Un/AAIbFNNmEdDZuF04ywsXQ4mknB8xF
QPWiBoeYsEoOpKS9dxYyhai+HGYz1NFZsMuNli9V6YNyunIcv3pT3QraGaayzSvq
pNF/jhatLqecZTmL+HBieC3QYi+O2I7+l6lDev638Nq/T+KDNaVWGHfp1rBx5a1t
iAsEjuWJ0o3+/MeNhq26r2VzdFL9gvHqHbNp633LSPVagbRQnqmvw+esGxltsHP2
ZBppI514/EXOMsvxB0y/BW/QgqgQQdk/4Bpnux7Ur2/Hv8ZgyUY5JNI+DGWZV6gl
odZtbak78110z+5EeTB+KDTKglwoqoE/Efo7wmiV1fmT5EvCiV0IPQ6a9Hmrgo6S
GfDhYU8mhAhDdZ3+xIA/GJdM2OF3pyIooAnzYggV3w6CA5R8x86XSQ280Q2Rx19e
g8WM1bC09B0Pj/1df8N3p6G6cABa6Uf9VKycb92uGh6pApua5NdYZSjkQxQDH1x7
P0200oovE3y1SI8Nyha9TI42N0RC5SkoP/xQ5P+1UJJbsA+SH741YIGQ/xmvXce3
8pQwZMhGNL18xEMyafJ9z3JUvf5a6lfioKqFA/r6lNG9Sgrf5CYU5rUHD/TDAiK4
dTiRJ9rsJlr1RKjFQ1g9Zb2Xcfw2WWK/9ET2ho5Xva/O60HbflTpQJXaGHvLJ0lS
Vyz92I1UKfqs7m7zAtB7DtiiNi7OkOCMvvMuUwHcC0vv7/afsmQYo+soLbnWPy89
MKSx29uMa7cARNEGtMGZdIJDpSDJNfE8IEacJxF6DVnIrb0kdeQeX47RhlWoNQL3
YiBdn9P1i6AhmwK4YpVIoTPFxohAtOLFK6acNNpuB1gzBR+mLabblyXnarbx1OjI
nkRaWerUZKl0fzcmdlpeHC6I/w6Mt5GwtQY0c9Fyz9mRVzi3YlPd7jstFZBqrBMt
+dzfZ5LTGpAoLTDhF1DTtzvwzrZHdUOGaQwBBv6YDwtm3nJN5aacTUiDHUjXjHU5
fKjikXrBN0k1BjSXWQFghL4fiEFiHjTPTn77AaBEZycQClmMtUag3fL6usKUcbK9
3WoibG9ZSiLg6VbdqMakrvH2bv7JFf2grfbHJlqDOTYP1Yy+Tt7kK0J7iGwEkf05
h+dcibcECjLkjdf0zop7viA3cRNRuPZANxCp+w3bW+DtdQuw2rLf1dgxWSpI7yFJ
XYHjpbPmB2QpxC0v2BLHZFP2R2cCzuIQF0EitN6BqwN6rWaCtqVp6SYfxwxiAxOS
crWYnEefdUf0CdeoVvghTPTnTxP3XADrE+WXNVxukfSmPGZeIkO/CFuSeopZ7wst
xllgs701Yzh610E24N9K/OaW8IlVjrE9poJlb4HMqWOW8Di9PAzcdLww8raAsoxQ
0ip92sr1otleuwsNTMyed0XP18vsTgk4ny4cis0d/UYEx9IVPjhDj2lFTxNI51fZ
YclFbmOtXmbARvWP7HOxE33cLZmViguhr4RYHTvEsg9/5Xv2S7Q9s75LMet1ioMV
+5BEDK1PmTr/TabAfN1/emtVV9ts44X6GO+LDZsFXFRbWBtvjaHVfBEzg8KHj1Xz
vMtX9ms9V/lUcMuqTAhMBWiksp3ia3S6O+6s1QqcBOEeC9tfm4oRHAqCvJOOFWyr
pNAvumNrHXdmQCNNqf3CZxpr3eBPNbJ9AfaJ4/F1AeHGbxK4m8jxB5FZHXYNmEoS
Fmmn9BBJ0jiS+2NFFavxCrVm3o29xePqUKcnu2kb2Ux7laAOfpGqhQQB7CYLOd+w
IRVTORxwALkjZp+SeLVIth5yqcZbDTneMla3JBnDA4cfYi1VE4PHqAdwRcqiSwPY
WiCR5969TdxscXwfpRqimm7FLE22BBOsYz3+6pexpaN/VSHTvuPyPYGKBB8VqkGT
Dp8Cugvc6A7Wot09TQS/Jgjog065AViQKgD0lIveSLioKXk2f03PgyTVXmLtwCFE
QojUIjGciGWBMDontaXvzuOvNiUBj8MZPbpvbYANopQ1Zz/7vbSlFFJ/dj7AT3gh
7zDVfslu8oTLpBClurYxba2tXeuE25c5uPjzmN6/SBV1sFycwUxFkYhqlCknW28y
hLwzb0mw76qKdDVQ/zrLfQKu3MSiM3g86zUdEklia4gZiOBJG/uGvhS3xPJb8egS
glsK3xYT3J+uIf0T5NZz6ncIpWz4g2m3vWFgIm4tcbDyrcDab+ZUx0rgkOssLbQ8
I14hlhRT50AmMw1HLBNqj47+2yfyRBLhs7JI0VjGGQVZRDLXzrb0exhHOmWjnvyu
HcecYcdmx33upLWtzZCw4FCL3J6zCWEfBv07ibazZViwObC8bJ/fmoxmqniOt0MZ
FmK4R92cJRja48JRqcOI4dHW53g2wpD26QbR8cax6EzR7h8cgwFzS5UJMDv4XTHM
cM/KLtkrz4vrKZLhcBBLJd80AwBcf3DiliPSVdObX3VwaECn6Iv7Vplaf41QCECB
SJA1r1yW2lS7aDWGjpqG9FXahUsgrmdPp/hHK3A/GSjC7nTi4ENfA07kOhtBCJY8
yBOngkm0WTPwpY0cpMpQ829Vx3T0DXbeq8kAxEjIlQ/hXNmeIHnkg7jfFZJ+tI5r
R69RA3ZQ8rRr5pMCrMbimEp8hRzCExgQ7hriU1rs8d5t1uME6QSkS882DPBr5O+Q
gv3M6j2/7h/eiZLU/pUbGB46f2FUK3EQ7/stK/2w5EtHAMqV8ciHPNLNhtyNOhPw
XirAvlj8e/5wafW4bSHt5fE043IimAwmKUl/I3V82loDBfmPjSGYzhmIASGrEUYs
0GRg4RdwN4nzXPxzWNWdhLiyunQLKIXMMhb5uUVf01KLabNs1rd9y/o91HCSt1Be
ebd7jkrAbHNpPtE2M7P2gyR6ThaS/6yLqvMQ2ViJT0RijeptLQ5BvjhFn5IM0Bv7
ZWRLDDk71GixLeWUliREpmE76WsGVpr6iKXrCnqNoMca7VvbFcwzsWrosL6C2JJx
9Xq99dMujvNPcKegZwsM0lqaXp3MpBp6V3rjTgyiUmGPCyuvRvJoooCgYlYGY2Ra
5uaA8JAQi7PwLylf9v7coWAgs2CsBx2UVddZo3a4IsSfUFMvcQMivWNlr/9IJHvi
JMwxsQIeLuoHy+0sSLSm/ANUR+Xcf4c/Pr1u+T/jPVlVlYs9+q3cfo+No3m7IZEr
ChyqzrFEy5VVf7ycuinPUrJ990QR75/6SLxzrr12Vkcs9bcIHh/NVCS/6qsjhRkD
CZGld9GJiRrfFbYAf5+CXTY/YukGCwyRQ53cak9Gei2HY1/J9E17aaUDozCkHY0E
t2KKS/baOGxAN5Ae0FAJ9l4V1mY36AbFLR8E6QTChsHEMuZ1jA8FOetgYD4xrvfz
O2NODzZjeXomqNxJMmI0PE2HYIB53PyigPjgyvOev22clHLzqQg+zS+0mnD7nTdK
gHrbYiuYO2YmGdh5Kw4Zrac5TUwnvaZSNNM5VePaWrjv6GQotHIwrfT3OZzLiQhf
iEndaT3cSyYY6bJizf4HTXsNAYFSi3TbUf0+5ZX5i59oytjNrJ9TNjrvQpQK+2Zc
4iyw10MryO8L+O3e9/e/us/CBsNWrWoUUw/6Fxxjuhe1grN7lb0aX2AKK/n6d3ga
3Aoka3cQ6AjIetcXKpySmvwbq1tiYEBN5fkeHVOWAmGmqcv+is79Nw2ok0bXMmVc
0gCoannNIPG7pUqcRVAuvBwfhu/AR0CLopVCsDX3y5QP8ZmmgAuLb0YGIS5WGtCz
6kcb6F2nOWxaMvZTJ4WNj65wPccRNuvRrN3Cf+jkV4FyVEjV/Z5eX9zPQz/ynfaE
mfk2Rf4HAdTyDGZv5WUwlbR3SxIyDVaw+IouCOa4SL4DDQUKsssKUdIhZAlvzCp0
HRuN28WrTQ9UdzVg6NKMw6QWSWCUMaJm1h4KnYJ08Xv8yYriVmgdIy+OrhabgiBY
cE2BP7XT35m8yzImNkDtnbiyyut1xh4UTh98nump2wWfT4fnSU5AGa3KGiTt/Goj
uG8Ii0FvCIgE4a6geoU7eYqhnD97NdsyhfQC7DSgKMU0UI6DavG83JMK5gmoXjrk
MPvkbZNr3RfWMMdKxz4BXI2kwwbfDAfqf+Y6aWjSIQYXFQI3Qmbh3eomGFrqhvtU
uVt/qhi6l1NJKF4Zw20ScEFSCJ0bhDQXQmFeTwN/u2gHBHqLK5NKO2tf+Vim9Lq/
afUMwoYfXQGiY16YE2vyaEj3AL70fzoK4+rept5rWnxad/M2sRCN8p8WcLYiyThC
EbuxRSvr2Muku7Ah2hQCna5KeKOQcpuCikS8HTm/ZhPm7Hn+OaYdxoHL9FlO1x2C
xuNbgZiJRAFxGGD23g2ooSjcFdX+pZEUdTsPwn1qPEkQHIhCQBPf61IusgPq2Z0G
QhjL8U+oFPjC1MGR1enUIbzcoSAOFcVAQotaf/XLzf4XCW2+/+q+XxUu/eGibtE7
ZUa5TRcGDmgPM6qofPPTaxneO6ejIXhb6BYzDi16HWuBixxMY/lY9YVPBYjLOcSD
mbrvKmb71Mvd5O/S9netAVw0+NrBJ9cFVvaAq42mpdrCCVVVUnraoAwlc+wrOu1f
5OqsQA0opQi/f+lE3D0cfMhtsUi2V0kMsvuQ30f1wukkBWvdjHnq6EWs8ebJw4x6
PftyyyXfayw47t8sLxZZhMITJg7Tr9K6c4Zi+Wtl+E2F20+18GbAS2wDpGyvl5BJ
CNw3vD2ajLGEUIZyM7u02I5JIm3GUTm7UGOu5mOiC2DYozlpPTRmkTC/fM5AJrSh
ayjaiWL23NnBK45YfM2V7W/keYHEnn2cXSVvM+jRjzQSzymVimB4mmEEuzE6IapJ
YegB+tq/2JAFC/aiXSWASOh0F2ya3q6WD54AH4RGZ0n23f2gYJgB2sFDMM3tX7xl
f7Pt8E7w2Mx+Sa8pnEdkLgkZ5kxZRzeBLY6FTw/yVQIUjQX1Orm4i8mR4lIvSdIo
dMnaQbdJtnDE/2ftrazg8OtpLDqzWfwwkpmNLxAXYetwYRoeqaWxDnl49fV9WXwD
wHUq1o5kLlO8wdJBM3m5YSvyOHoWsHb9NH3DjAoxNVNA3YuhYm9eBc/BUN5uwYIr
VF5pdPNbyuJJSXX6igruhcwK/wEZUNxan5Y+eoO+A645x/efsAmBdugdk8Fh9dZV
HAxQV5j0UyB2V17cSxZxGC+fpIpP6KTzAvx0ojHBHYE4PIxeCGRV8lsq36ovG+d1
t0xbt3cgJSoTuo6bN+cLKSI7W/xIsnCpbq6RUbvlM9LKibMAP1qISkbnV4NnCYvb
9B/4UTtkFvitOTJ9v39zB/32vtsHYn2lCmmwdk07BAz/UpphNB3kixtN+oUlKPWU
WZkIhAiZRN8GweyYbWiC7WPpA+uDBripr8ZMWfGPFXWgfaU9dSyd19OSLHry6D6A
tZyWs4ZyhHTSOkuzMNqqmLdgkfB0XGA8Fg3iPN/z61w/EdYvpB2wQb8C3Fmf2/mi
m/dHYGOWhNrMGrhWHGI68pqgZbOnm7Ocidkf5xvg+D7sh5DevOUIC2XpncbN0pZP
Ja5aIE9CxjzcAzTQmwd6Mjvz6R+dh2nrhLJR5LiSk9NXeGNHe1kFK3ipvKXSWBVN
xsO5EuHu/sKesLtDYwwUxfUyEZsOReBfsq0bNp0jsbb5/JoWEE7NVHPPFh3MiH3t
YLBB8YY/At+etQRq8g8b7w7wDzmMwcLze+uBSN6JfAsiAA1tFBihoHYusKVX5wXR
rg9PTSL65zsL6qcPwy7XiakGQrnOMI1FZ25+vPhYvO6g73VPs/MWyf4YtbY57lmo
FA1/Grz4o2BRXnM8ISxLca1iFgEKBEYQzVTucBPNFb+amTiR8JCOaTtqet8xqOVz
jXUFvdH9HzGFxK5qixafiTjniRhhGRPQ8o7RsJCWWLK+YxusAKazpezu0b01b01O
pbnwM/NUCaj/eh0mqa6g+5OxdULbO9nVpvCymn6kDwGuWe1aZddo/2ogiPOoAnH5
Q4Lva5jUXcCjb6ritaicgalLrhKOiPRzEuP3YX40RbZnXHMkvtxwy6nOPeiARlWC
Lgb5iGD/IF1Aq0OqSYpmQY8xEcNv9yhQYRpy7z2C3Itvz6+fIEse/KlW11VRxob4
qocKXVndRPwJsIRPhPLhfcciVKJWKz6SPQTTVXsNdT8UER1L5XLTB+xIXwf+ZHpG
l9jCqvtIaL4hahRAg40/qPRM5yFwAAw3auuLu6ziMMl249zhrSXAdWvk1PTJsfbf
qkVt0eWJ+/xLtYITW6S5PZaY+uwJ6yf30QxI/nn168+cgfNftPv+TPN36KXYikPT
xQRswpU9gHt8T/06MMZhHIaAI+vmXOF3/x/gemroGIEr01wlbh2IcvozrD/7cunm
j9UyPkN3vnEZN1wRURE9N0BC+8m9rZHskgNd2y4/PU35K9hC1MvhamLvF494VtBO
QJjI9kvwDp3Oo+DhS9Ey2OBCkbRiOadeyJQnZyog9equEX03+nkARepmSeOgK6tg
4MB26E4QwLcHmmw6B/qLq8CyeeeVt/b1QB55tARPOOUBvohZpUF7VudWVa5V4D5I
LVqnGuoIviYFAmyNgJw5DBvA9JgxEU5+1GWBL6KFQzb9Te62j7V3Be8k2opIBLGg
rKdDxtdwbNB5lYbbZ5fFhXogPks2oQxCH6L0cidoRuMTZFxkBOFBoHPZyqy516Ui
RYfIhmf+YA/054MvCyGcW5OQAL1arzqNYhLR37IUzUapXt0Hciz2AASdQc5ExhVU
V6dKNYaixIYZz1Nlr3XoIqvXwJ0NCYkXE3ZhqTD738Fk+GEB+4BSjD6CudUjeOyR
z8wemLx5S6q25Z2Fi6LAllddYjPRHiS8cGR30OHZhT/QEqSrL5jrk3Nrbne3lVtq
U0OtxFfjNF6dWBzifWQ3BUSzfkFAdHq/asQC3A8u9NYb0W6AmZ22Tt0cRUQo4Xar
S2Ho8igGucCBVA15ZRuH1Niqj8CVoGZfD3T6psltUoKsrbBPZUGggB2tmJu+LMec
amRpAhg8r9vTK6LPmdftQ0oa/zcFSz+KumkjKbC6YYMrGQV4qgE6TFAzuNaANCQr
U4NSKBk0i+i5NBH5RpPihFgkBiuQFOgynzV55YSChOflX07nxsX205Qe2T6x6kHl
5HNQjiXPgH2Eos1OedhE/JWLHglC6UICoHe4LAMmjy2Ca0MiA8/nbu6mSKh0iHY+
Ay6wAbY1ONwt7g1ZNxc6YYCjTjFdAEMGLQXC44TVmiZ9PF18aBjIzYgRt4S7eYjF
WSX4VQmIqa/0oYK9LoFi6DHF3qGAw9HY/3WjRrdnFMs3vLFc8QaWUbKF+mtxjn9F
eTH/Z5OxEfDuU/XFVWRuUs7Hg+SYUbAuq9liL6K+DWPIL1XbffGOvDwnCHU4tt0B
AEZVaudJdiILXAZwUphWzVy+XIozKol79SU7VsO+wVCyFxsuVvceZu3FuNjo/sFM
oi8xXlwQHcz4ft17hAFeUaZubFFdwB4rs69mLaQpgZDhK5U9xIP7P+SXciv7wBTd
cyM5RGVzNd8Vd2UkJoPd+KOKYr/MJhkfmVXZRt+Dg3wShmZtjmk1f/ZIaruysFJe
nbujWowEf4OpcyqvHOEkznkzeUMIBBWIMKLs9myHxTbNbtFyCWlS8yyi9PUx0z3i
91rHhRx2fFyrBzdHfvqMH0TR7oDef5vOYQKhTMQHYXgCJrhhqwQnJ+8hmrDIMUTa
aahMasi/ThqofL9/e1/CD4a3Zl5BHGq1wQXd5RTaZC3peEZAo22rx3zCzqkoeNpa
s/eNjlHgBCFjjW9Sm0qnl2LvZfYqFJXV7CljpAGgneNdTkOaHHG6uLINPculnFXt
X8A/zRjpWA7G76O+mayrukNuQyGEVA0O6vBJNnTwfMdsrkLv9iPNe327S1W6FyrQ
IrILO1OjFl9XQfu0vinTP15zu2+INvZnyg6RkUvgKhQlUWnMLNhYvdRTlTvztwWh
qpKtmdND/jbd/HZhnlY+PsOStUVyLXQ54DprQwlfuthx66/ZO/rTjr9OYq7NUwJE
O2rByR7tsTJiBqQLxGcVzv8xIeFWkmMAiwE6CdX4Lsu/P0Q+iAOOoNdUWVlgKyW1
qNx3JiEMcbJlvttkAZzOugxdmLOJsTpcFPaBX5lYzP29Fgz4/RVjeFbQqVD1hP3F
Z3Vo3JZHIG3oQgWnU4Saunko5FtuBEw+S+eKGTGi+M7NvC2Kz+aqvW6+W2HBaQtR
xynnc70PUOZd8ztjk5FUKapMOgKaJpPG08jogSBwKIoVPHIH+odUwlefmdhvaq2r
iyvuZ/djj2Kpe1R4MZmDA9hBHLk1aqn8f+7Ja1shNGe/RD1ypXvBcJIzYWrtm5FI
dsrh8sGOFhKH06mKxT5sQd9kIkHj4T/DF330h5Ot0FbhuDjCUoS+TI4vKbJPN5F4
f3kylQz5EqSBHSniB6s6te5zprL8HJtMKC5O8bCPMaWfuDB75wPQV5GHRb31ICOm
eWM6a8qjnpL5IsWlYnmChodxmN0/NnrhdH4AK9zuwN9AcAK9OZ+61aRrF1PtIUj8
0LQa8Q5wtSYdNeswlpODnM5qPyQk3U1Nk8ofWSAlVxIMEhXS+O4ZlDV4JLe2iCP6
5/3aSN5Y4fsGaAtJrCngE+CDLFE+LnBj1iNhmj4re8nKVhcpaBl/lfI5b3wzkMCI
srflcEJF0ZdMeAug76sTQEFglHbRc977F147o9dTRHFP6ztCiODOAyQueF/2G5Ko
MRJG/sX886BdlSA0gdPSynTAQXgFaexqweSNq2WYEusaFwlVx4DxztIo4fOFa6dG
b99aCut4jiyeOHVLEDrnVZDpwHDY1VbHvwICIYwiDNmrLql3WrgqN1YNXKcjNRQk
ApeoVOqEy7o0IOpsSPfsXMNcDt0+zduPAHPKqSaRAG62YYsdyJz3b4JjpIVOLAqX
R41cHCl1fjCAfI/3PEw/IZrd6s1p8i/kR5kuItIskpCLfXRTManA0Pq0+IugasVw
BQ/ZxM98XWApEDvu5bM/HtMb4/3eVY/u/yoVVW2TKWuDmSbWaSKP4yJs3znwF7HJ
xQN7nB2d8S07PTmjzVmgHedwt0eDER37Ww2j9tbDfL2LgemAiiD2NRcaODOBERfv
XLUbcJwJdkmnWrd42UJRETbn6iMthSg/pa3nEE3LBuaOQB0urfCaBm+OtQyaLYk5
hIl2h9lJFVRRPqCIKnGKDscuwCqROW8Fm/8CCjM/yltZj8A5R6rz5jinTUeIR5ix
Z63SO0QR5zGeM4d6PzIka/YrY5Ysj4dzJ30yy9PXRMefVzgg4bYRgraz96YOrPaq
+SGwE9lmZQUFU3t8EOnRq7hiJJSIByjvqNsUBgU4Sbe8Fr+Eg4oHmk8IuPt9l3+b
jmySL1tpGy7EZ+tHKy+IBmOch/k5fgsZWTTyqmkN7yAJhA2kjm2BQ4LbNQE7qnjT
fnG4jzCHkInnfeR3cWX918BE+TkS2hoPHZAYZj3h2yd8aEGlJg+ANc4qUwnSIFQr
nrWsSMmYcGkNfpeMdk583s8qqbH/HvtmLvyEs+9PznreOyS6Eyjx1MF5rSF8Mbo0
mcXirOce+Tyxqspy+q86rjStuYD00P+/1ofYvVeId+GiUNK4DGBecez/HKnek222
SlZS8F4M69GLI+n1lTG4+/ZnxRL6+9Rr6ZK/65f+qulHcrCZVKJenyuXMnQ176nU
ysYRfWzue7BoFW68wWlbgEjk3B6+8n6FRZv0MmYTa0uoGVqxeCRaJ4APw7+eVzvB
u5hZz8hmPzQxCzHKRmfBZuqNvjHSaHoJzThvedJ7gmKGPO1JCqm2A2XJb0VJ9nMC
HuRxP+whniaEgvNKl4p7vZFIDqt+i28tT2aUI5VWnlNzGhOUEgkxiHt4Crbohd29
1vX5fbjjLr02rzy7dBkwVSABF/Ho6ptxDwJQ3ze2M+2odH4mb22n8XLp/EAbjpsN
2mwZtq1Vf1Mjv96gkvIEO8GzC4DKzve7wK8n9cOZ8fFt8AYQyh/7oiMBthW0vDhY
9LiAfuPRDxogKvvZvpYwkWopYHPN+3onwimk/qW1g4wiJybi1Bsl4hO7LB2+VLHY
WjVxVtMA9hSfVVzFIVuj5c9AfrnZjrQOx4Fg9rV5HyyYsO8q0Rq96MgoKbh+Q+0s
KvYTKbPCLwtKrLxP+OI5d8fvjtr65hEUIDBM7N3PL81JdKh35vdldvWmFKzFXQ5N
tPWZIo/VTxd2yq6PWDZrz0hNHgXnz7T3j7yfO6F0lhiubjJQsEqPXGZ1li1FdrzX
NsK/8OF/mdnyyCePPHH2CrYkxQL9sZa90dbLDLwGlfRBSjEka1pMI28x+N5520UC
6juo72O2rRHF7D8K9wlr1XXIbKZXmklnbpM0ZPJtsVJ/OxBUePaGd+gYX2HwaT6S
MbwAa+Q5yRtX4q6NnD+RLUT8lMRR7AJmDN7xzrbJuCOqmQrXANKiWrv9ZSsoAd3u
o98dB+hxM661LD/NOIbUF/CCaAA4DPptSB18XDxaCXDxRlr/+bakbWDKmZWvSJdf
xyaQiNDLOl014iUiXjkjfXFGN9sWGhcQbryJcUj0ydwN0ixB24Pt0+8fVR8UVkIg
x+POZpPekjzEmvo719xFDFKOQ1Xs83ZzeBpNiAaAfIm+CszsOfXS2+gGv6lE3Goa
2Fng9lEAkfzyoJMPAz0k9Zt+38o/eAA1S/69YBoTaN4zJEKHHpGAkB7kUmpMFsiu
hKJb64k1ipUxd4Z673Tka9GEyPXRI7Vadarww3lffwkKqLVIU97l7YKZtGF7bh1L
2jTtvG3O+a40V3on3+71GIvJQqxdwNgHlLUwJeJRt+eZqCvZ4Qct55U7MhgEksXa
R4EZa7Hboq7bE0cKtpA2Zlee9Se7/EQt2WTaJC0pvuRJpujmK8se/D/fTdnW77cK
pW6p0yxu9D65klJ/Yqj3WJpamWTUkubAjYthoJ618XZOEkaydn9we/4qa9I7L7BI
g12DSQbqIjC+rq3FzECv63zgeF3heqAmrbaTFex06+OJ3+PsMDGgYaT9l++BlVx1
djEIaAdDdA7EhlHDHlTlC+T9dTkcTE+hZQ9Nx8TEoZZoiCNH9eDFWNixl71xdpjK
oaSjueXRPJGHioyRgKW+9GMhU5WcIYyFCkuhpxVyeNHXNY+vzG6donFBc0L+7AH7
XzhuzBwMHLMxPjAphowiYdepoXo+cImGl5DpCjoB+r8nb5xwSlAVcG7onoO0miyz
DbQcYPhuta81aEh6Hf6oOVs/Dg/ltAD9dKNCjKB2VLQbyY3nFH+FCpTDPTk5brVV
2MRbBktAHjOdh5Ne21trwovzRGrzKpsG4u2oMISY8LbY56BONYXOYMV1hYhrQPRf
39b/V2QBZLbFlXZERORScqmpTrPoLU+h5sLBFOmPmQbQa7sLxEVm4L0VEW6WMraU
YNvy0TizUIVYpJptL2oybg0OW9zhgu/cBkIA6uYbYKyHXUgDOL3UfqoFXn/f5ibS
43tf8Bzg+24XYAPKQ8oB+tI3qFjWrNADXspe8v72AYr0iH+gex0AAOCP4RAIfBF6
pdioxQSAha2NCPqKNDicg0LUZJHoGwFLvPOx1xfWP9bz7Nep/VKI+Bl/KpWWEBWZ
dCLXexFS5RlZkOJTiDa5v2eX+kyEHx9vmOt4Y15XRa9n6W8SdH0xi7HoJ6tsLcpn
Vpt0tzXFOzid+hAo0k75nBzvK2iFb1XEJ/zXakkTuRliXEgl2BYemsOqOB0003Af
+vMR7YpQP0iB+e/oZUPpn9KZu1Qkf1VHpOKARdXViqttiNUSJJHgNBPq9MBZlvn1
0PA2PbJ6zrP/7//qo/V44ZFE6pfFuhXnwoEc6WYs0PVfYsRNm0Ega8S4lyE3Jrmx
4R1364hiosRAqoRgrYhsTP+qee7O2bHk5UFzAS0DAEFcJJXgytQ9/WQvnHN0bbKn
VJBMjNO+Fz+7RQxykVKMQw2ybdn/eBIrALdKuBmpHEzCDTJGTmnvtYyL3/zXpfmS
aXsmK15dkU4sE8MEYdpQo2KXMQlTCqrxdpJkQQ0bdmiBBsZjXLJN4y9XqIx+K69+
i72SN6392bGFGxJCRIyp41IQSrQn7dSxD2dp2NreQMkePLtNuyGtmQPx3bx5MwBK
Jcsk0aPIKO+afeQwYsLIQc7PPH/WYdIa6hbZlPFw98fzWpUUUs4Rop1Jjxcr0aTG
itAxAl6UI/UNBBWhpUEZ49BYFINYg16ZISNJYKgYCa+DrXVGpR2uomIrxE48qhLT
hAVSYnyL5wkfKwlvKj+NWqBxbkXeAuxijbnLMwz4hKlUt0Obt+IMTyyRtVjjQ9j/
1Bb2oo0XE1mBaSBgXxB8hD+eUxRDkf4/6SdVGcGx3u06A96Usu04A0ShLRFVEkrS
hl9t2hyyvyw0B2na7bDZacNDRk5+U4dP5EkMEA2mPqAKe8vKb2Pgb3WUARg/L+9b
5f1VuxOyHHFT+RrXRv/T7fPI3fSbAoRe3DJIkRq7mcM9VpE12a1DZuCOK3xvGwK4
4e9fFVpk5ZClOM45BrPem2cIWrn/+Vm1R4lOaOPi1Xqz+jZhz5TRyMpklPwvTpbH
zpd0yN6HvdcBIb4fklcybcEVntH6eN6zRu2JRXnNggj5bfcnfksb+Bti+s+1ygc7
YIwxX+z1KfAflr0RoLL76luqZUB/JbzXdGBJdZy1baV19gDBV5xEUOpGI7vvh0lw
P5Z+SeNDyp7Uiimo8Ve3RMS93cxFUKBiWTHpRnYS4QP3iHmUaqzp/iUsNqrunDYk
+OGBoIdBSdA97/z4sh2ko9IT5Bxl7ZDTZ80z5fmqYXcVpYYw5uk5z5joXdVqcDip
AqKAtpyCabWBbVYEn1jF/osqeYPn4PtU9hIbdlNHIuwT3xtP3p0qwq5ye2UWvwyd
Mzv0pWwDLsdABN8J+Rivvnzzv8iOzkv2RQZDvuPJPRjIf3S/St/h1Foh06M3hWoO
HMp/xQ1bRQT+aAlTCkUaBLV6O9wU04YqVSSpj5XpcNFVj64QheQKBhYTb5bNBw5/
fnK4S7TsKGvVu8Lv+oGfAiQhgiYAk8T4fpVti2IXFl5pxGOKmUFkQwL3MzMJOVJ+
HxBcY5str7CN4vmhrBd7Fvw/JSf/5Ew9qyT6kBtAJjH0xjSEL55aETyMSEuMqI6k
RZXwjIeZM9gVR6bKD20fqpf5+/ejreq/MXEvn0JZmqAuQYwV8pSI1RxXcaTk0WHb
nlYMfv05oOUfYF8G1Rc1cKlPVi+CtqMO5mqV6Baer0DGa1Ag6Mgx36G0cQ8KF5lj
eEvwtzjVScmDkIhuCPIpMjZhcWWb3xbE0cdLwl6buTtkyrjfrmgX31TPYPWbFPP3
Bruxtnc5IZnmnqtbInfp+A4+75R1nlvJS06laMqEo3W8ox7Cusfh8Z5eOitwJmpC
Uqw3kdQ10kzAzWUkjqEnCj0G5EUS6QorwCEUWe4N/Q8bgySg7gM3d99wRKU/I6ve
colKn9mjJJjZPAVC3cr5S1VZJKmKa2dfipHT/lBkEPf7yKLQZ6qR051ZumA1w+t2
Hiul29bmAiEGIxzR80mkZBNCID1/XQN98+ISksCCc1cBdaval+7DdFwjad4N2wm0
SGeGz8hZbV6U98yTtAgZhOiICIMlb8mf5EI18oMRkBIr3dp0p6TD7kFWdxV+1TTM
4Vee8DiFm4Z8ZznznX7NmGfbeXd+5DORDzwzDK56KlQK3kn/Px4RSb40B1Dh6Vf8
31cK2s2S09IiNGWCZGbedJXbacyLP61rY6D/0xn+INXMFW/Rlv/Q6UXTfB8bebSy
MhDiSS4V19Y6CH6VS965FrPXDmExECN25ChRRZDQzwOVTglO9Z8t/lzp6anO3nbt
X+/V6hE/jxMDyvPHpB5TBs5JNZWPH+8rn/USwIc6RhCx/jnNDYVT+BGMfdYbmYPD
ErIHgIDPV5wWi0e0bxBDBemCIXd5EDmATPzFt187ME1yBEhHz/ZBIUYs6Vjas03d
tJE3ox/hd807A3BiqtRuN0hUtBUX60t4m73ZSLVEbXU0Y2HzuIwUsE+F85myHIuV
9pU6CxxRJMWLFeUbzDQlOH4fc3jtQ8M5p2ARC3GRD3ai0WWejDoeMRREkSG2fSFM
N2yCnPzVJJsJmqTAkOuWyKjeOE6MHgA0YZvEVRZKQvDmfqcmMMgOwsEhg4+Fr1O6
ctUzhUYr9hk8IGsKtIHc4PE6AKByHI1hAleSxSTZXowOKBK2VUoSAMcIn2g/DXT3
ze+RU+TR0RRKIGivbgMsL8EXLFacqN7KCGYC/gHpXS0pSFsP+uIx3wg3K3pC/D2G
ElLBPVyniR5gpnxzBgkGt7WGsqgRlwkaIGCiGmqqsZtco5HUyGqqAqImw1XzuCZ+
EFtcrOWLJoWk1PRVPqzF1pkRT1HpG78afjxcDtJh9s0ceimut29QqHVCflIfCv+N
8pFOkoj2Spjr71lR37JczRX+pZN9Mm290LbCrUq6zXMkLNEqO0MJQckv5m9M2qB3
xsl9seh8Sf0KPySKQCE+Vxp1DRh4W12TIoFpD3jWcSQEBDPnUAQjg1QHwvZSfaqG
bpg1TCgNqsNHjZ0nXcaISzCBcQl34PtG1zvq3wMb7j4OmlAFj0vBNexXSGJmcT/J
wrWXPxMecnmHgssaFyBNAMbIo9uoNKZKo8SRSstRTLCpln7TMM+jx7McLdjGwz4S
Hm1xm65sV7016FDDkqFtZYWLxGHhKXVon3lgZc4OEiR5GtSb8nkYq7/rfR9qlh6n
LNJGBmz0qHJLn+qFv29HJ3Mk9Ri66wRxs765JhVS3K4icyj2iuiPxleWrwex1MLe
o0HA/8fecYU8IeJrBXcIqL8ZfsAmr/buNIFn//pYVgkB+mwk78R2xIUgNt55pFOF
ElYpXRHZy8y1tu1s6Yq+jMDbwAAqhOuzC9opNkdiP6nN3N6TfgSS4G8dROg3u6IT
63WMtIYKujdh/bVykxN/GMuetX8/wCzdum/kj3Jssk8uh6h+ROe+KR2W7V54n7A8
vR7vngMDPL+CWjEdJziL+UoVTFjhkvTylvtWqBqjx4uOR/xtXtzZ0aTcNKSMhPnq
bmS08xrMmmtTlk2FEzyxJj8eBcllos9XH+cwrwJ/WKfbS5gxLV5/Q6mPSXD/rmio
pp90zxdPWO9rXyHUYOYImb0lgKUacwM5lUmPwhyusDapkiwY2JsCGBZLK+IpZoUR
BXTpkmdWNU5CBGBuOnvoFnQZJBUclsgXJK2M6kzgVXyVdt2Jm/aNb067wlr2828l
qfQtVIOIMyvb7lZ2XulsGSil2wjI3WV2cx5uVl5j93wEQqqBIw2+i3Yprs3jlo6y
qsmZQh2eAErYUxlqMgCIq7M+gvIpE2zW4mjyPslKL9TY1GUUhrlMdjzwAJpoGsPP
31sCATP7OIxudqHCwsINIufPjA4pyDDbOhebD6dOVEerRu2UOepahJHVJqD2ge0a
cv+LL5222JL1wKDSa9oFBuuChkm0hGVUIDN9x3ZGjKoK5+a/pmXAIaJqNNhLCc4R
XGMqZDayXq5WSESEueVzGIuza/b7lcGgA1CEiQUUD+uL52uNn8yTFSUpC1gEaktm
6NihkmEb55BQ9OfvHyRDEua0BswmoqYqns00M6Wba/CtgrjQQrAQzEu6u/MQUThu
FJVg9VqxKk4bTSTiLffF7ui9xMAuZnJ6ViLgP6ged6wyaSx1pOPcO3msfYHLEYJx
keeWkCPX5B0TfA+ALMXP8BT9UG4l6Pi8LCilgVQcBzQg2d0Z6X5j8fxyCp0C1NPc
8PkAcsvaM6DlItPNNyVJWEgaPYn07GW0PfVNJCI5aMAQFW06zLfzdqEP4Di+EUxS
KappF/hgCOb2j1R+El2svj3GeWU8QyN5lshVmOFLM6gcINzDsSenyga5TMBn9iGy
UefIz1SEtsM2BEOAIs88+DW/FyyvIDtVsnI5SMmwRm5UEJcVWzUmKK2F3o6/5ZCJ
71OxhHkYkHUXKjj07pEYF7vzBmZ7+pEKVua8FlosRIXUkkFq8DyoG/Nw8eBAa7dg
O2SFLxeY7OV8cSM6BoD5zPHulO/54QkU7oSNUm3gYKsIdhD5p7JKgns9uqt8lLk3
Tfs3jaRX1WgxFbUpCi6+472fePZCMxusI8BpUoDlTpAuY1lFJNxoKbyyqJXgVNEG
1PI47tha36JSZlXSXr/xHv0VP1T6kcK550vhzizbMoPO3iBhTJAg5XZ/rkPMljYe
GOVRrOJrhuXWLklY47O2CNIEzeXYUT4yBHtTf7NoVNBqtSsbI6tniI8jsKf2luaS
euXuKGfwpszd6TzaenMHGctBiq+SIlE3Nj/dxp+WVXtzmCmY9NDqTnxiYXrmeJpt
Jwku2UVyhtu8YdKKaW1IzVUiWduySrWxoWq/dNZ5zYXtoJwVaSpve7E3oWqW9Scn
60xQKtIfyB9CVWjxsaO08tB2ZzCPXOEV68VZPQ9XImhkG81205Iz0i7ISuwow9+P
UEzKMYbpPr1eobB58hJ0nK2VVGu4lDy7WA3/4MMvkmfOSkUbw18BDGQHagWeQjWs
3Hg/JUvmsyxYwGpZspaf8gwyCKkW0d+TDlPsEEPwyubWfUoO9PqgSRPESLe2aHvv
/r7/H2JIcwDEeyXxzFYxidOHFM58plLPHB8rYSNXG2tD3acALUh1YOTAFmb5qiGQ
DXmUYp+FA/a/Rc6AMoDsJyozZqehwS8cbGWKNUtG5oMP1U8GVcPuth05wXgXiDeT
d4DglEZJe3r5QtfdRV3WsSmP9Jk9MeIrfbSQPoXe1RaoWSWcGddBEL/75MVcmD8A
3nsmYjae5omfNLLpPsbW4nVBLcmeyBuWuCTDah25iSVUaQqa52xYvROzaI9lou4n
znZscy02co0FNVuagRZdGJd/mwZzuQ7TITgHhGwozr1Nb0JoGdbBUlmxqxgLgxUq
iv/SFZlCTD+lm+QUnTDVChYtVWR5XyOqhKDWnYhxoWWnkJBaN5cf6ViaQHCL065w
3wHn5ypFOH79Y3JfId3M+pXV6f4AOo2bfa1G1F91XWHpQIIPWsFIuyDJMmlIXCgF
n/GZ41ve4wNc6dpQZGnC2gu7pCeq2GX2uZFnrb+CC19YCqfSiPCZUqkNxMeg2Hwh
dGkQo1x5hQJC2NYPOJIJfE7zrL3DxOUsSNhjIvYTJrllyE+dY/sqE+m8rHm9HAvU
gX9xSTmOc/ozwck293Ptl4JHvhVWXI2SJF5Q+C2/BEfeN6wduLwDGhlpMpbt5hJR
XLkpczHh3bDIb1Ljx88NIP2Uri0PPfbSNwF2eKZnVKyLsXSALdt0NGKxYdF/W4oe
AZUVFXTE2lsZEAGIQzFEYnVJhg49s12TeHFY/fYzJVAyUIWRIGV1etJhrfSTM27Z
0WaSENWIng6CiCMlmnXjn5XtyoNXZuUOY50ghYYEYjAyv9OQLJEtIqjv5EuDe045
bKUjOpGmy44fp1q1E+fwJEhO2LZECaOU2m/VZKpWvYI9m9DJHeEhjWg9hA657VJd
otS2tSk8JwKGK+xqLdGhg0v5WMhmHP9Cl2Tr754rUSNea2Ccv2NKt1bphl9p+r7p
HotqKJMlqi4XGC0hC3+2mEN9Gnez+AZQIP1UB/NwjLqMnMDUcFs7C6FCBrFB/r4m
nr0bxmMo/9mefyMEfL9iCjq5JeIKd7/HGbWWoRFI9iqZOTaKjLnZXP8X5S4/KtMc
yt9kaUx4cTVWwcbqoLBwkR4Jse1M9+XR+1VzVoA7LoFPqLmPdKScnex4UCGKjaQR
V/JNLpr8m63/jg6hcbn+dGnBScXhjh/Mr7Y29UFZzA2FSJR1/QtBrnPdL4WAcVlZ
nDEe/8tgl08zoEfvYDloe3lAACCmPSWN17HykceMsBnfkTSETvq678x8KU3+eMHm
6a4dq3LACjEepAMwBlTAxoo99wJVg76wrXwHiufzrog4QUUy10r7QtLPH7TFTdvD
kp4ufSz7+UmqYODOjj8ozI5Mg/l+p1aR+cSVHRfq2Jt54DbgektOCH1xdLzCKivb
sTcXMUTX+8sReHg1bXq4ArpbDf/j506qSv2KQy9SeP4j4hldJrn6iWq7029pR/xx
Z1U+041B28D6KHroduJcDhaS26K3/Ujd4FfU6NlXM+PzSAW/a4AvY1HQKAb3/nTz
lTrO5HXgojfseOcEqXZM2fg4MHq+maZtE0gt+SgPrvTRnn5voDbMjfSglTKoD/F3
LI2aygE0MK875dBJbpxTHNrw+SUVrW2PGKMyvKospBBbSF/SGIOuSOuLIdhI/ooH
0OQXRKlKxzNKAFjjWuYP8LWAekafI1p12DLWlHVYGpJqHru68tyJlTRmk8TpxC4N
H8EGYmj9SdkvFs+pDxFpupcvioDz4k7K3UdoPD3ebJC38aI8blMJV21k8zVJpFKL
ZSuoztjWi9xxjG1D5FP9KIs5xXYSOVPbfE9HOfPQQueGvXzY86vilsnL+iWGNEhn
lAeuMPalU65nqfg369W69hlEA3V2xkBSoisTp8Wh/TX53yhRUqVT3K6HdSuXKYSQ
K8b804Tw2kdhN9wNqbRoBf6PfKrP3aklEc5P8S0vuuIcyB1WBN6ExklMxsNpzSDL
writ45mNv2cwBzOh4B8om21n+/ZTeSLda7/FgJF1hTVr879iwYK/IPzPG3zCkvxo
24liZdO+/j5+nIvJ8PHKCTeece/1fYuu1wbfYj3ESCrwlig0p7it7db410kc7iA1
zDobkAx0nPydul74np3yYJ7GNRBCrZ8nmaaYP2X/dp5hQSUNz36sbgR+xnaTe1Cw
N56xOgxIHLjYTlHCqh6yTWUsxueSVqYCCt+Ox5ZMRjWClOcgQrQyxblZ5k+hd38x
UpqKUKiK7869T/+xguo5jxKOO0iQp8QgBYlgesVKOQtOdlJuvC22YUBKs2pRLVOa
Wl9AltdqMO1CvuJn1JZlLSYsjdRmKwi0SPuj1T9RtKwpNiFVRiGTTuFk3n60YjKS
FZLNuK3/wvDYsbNXogwdbGD8WWi43emeIS6+QzjuGHFxQH210kp6qgpAbXjFjoGK
cmrCRCOd3Y64m412B2HutE02FqiozvFzht83jHF17DjBuCaw1xuFNcJvuRzuvGf6
lXXI3R2pOGIjvpQeIJnsRUixwzhL2tLZbPZf71oojPLQ8tMKOG1rCY4f7Uwz+Oe4
T2NUAM9Wux9NqO5SEzWQC7ov/VQhJMoVBAiXQVTfU5Du/60lDuuBf+xPcLibGYQH
nCjsHxv490OfvmIVyJGAS5ZFiMU4TVzuFXgJx377rhRIrtQlFxm8xB85RM5dF/PN
T6UZ78gXEJZ/ljPUNh0oqScF63tN0m7Rcqa18E3gjkzN/bLLMa3PqrWBYAtg09DN
vnrwQMXn5cMXK67h8fQ0Q6AsdwiSucHw+w24hAX3nFIaS4EHFu/g4lUMc79jYUUS
+SEE6NnfDticzTmPqK9BLJZxdSyc0qwOJEH7X0epb/zHBSSRISOqZI/19zgaLPOW
xsbN4ZoxKKYM4jJhQc0RC60uASN0rnc/j6Y4SLznLDa3wa9bai3tnokeMK7TiHCY
QVU4T+sXLrQ5Cv4cOtEdubMBMFNc1Ac4tvJGpieTL27AJdydIv3MgIoTRqPZkJfh
gL4cPk+b/MIy9oEvgWHsJndiaj7sH0xCfQjMoItVE/5G8bGxSNE9jM3lSfnyjSSo
H+V/oYF0MWl+6k1Yyv9s2gFaFV37QB2QLwDKPge3P1l3RQglTNMfDsCTJc+gW9WB
eV+UxKyMUEXYUB8E2oIWC6oUh2Dobbx1uC4brox9J0UYNcgDuY2mEGOtHWfHyTiZ
C5gV8A9xN8kE1BJH0XWek4LLJHoQbgfBtuRkHZI5GGPqSEusY+jYNmokaUFg+GH/
nkSkj08qU7HDHednZcMU4r15CW9JgWGnx9lzYSJFinJaTUsP1ermam37p/mt+gRw
YM6Jg8mlv1ursMJhXiAHqWv3/+POXLpncJ2ugdlF3CursuasQbxN94SSYDEEv6A6
YaFM6u8uX3CC1ClmSZDKix8HSMlAsbz6Ed6XYylo3K3cehyZFtYVFSgAieeVd6/7
KA+MBzWgG0SnWBdexuGlSFK+M2/1/APlfh7QqLq6bNvJFytUsGQ9Q6rXURb9Htmu
mS5+TTahv5D9jBu4sbdgsQwX4PPPAVtzDHrLIUJvlOHY8df1ZW3c8v3YX7QBodfZ
4IMBkDM0Wk1Zpy/B4WBTxpF354Z0msAAwIYf7+ApapcO30Ld/F3I5FE+OgOGwFOZ
eepVzsh8cI6h5cwHv8Ui66v86xwrZtEML+xTlA3tzbtXZUPgCeCF9VfWJh5+Dn3b
mNsd8Lzes7nuhEle8Y7Txe/IFh8VlHZL7RGQhfLLM0/j/j3i4ZEOE7hxvdOSelNZ
CXM5dZrqLjxuetMTBA58Cs+tnYhsl9BMpirzZ6zer+GvJZrnvnrKFAkoatCdAabq
ns+qdNznb9qHDo39bjt67Y1+OZVH7E1B1nvKYvsJnJEElg9RBdTXvaKfo6fFnRdN
YT5gzAiop66soUpE/BfwMqNeeptR6mYIepJJk26J7Vj55oyLPQ7b2zMcFpw/9Nue
6FOEiEFR+2G4cJJRtGH17TH20NHhTG7ekSJ1hO+34eC0ulmqBdGTe6e/SsZuObGv
hFe1t9pmL7CjbyZlOhfQcRDLsxOr6W1PdHS1Dx7HiAc9pyZPeZDHYoDVO/5ixjyH
Yf6Cn5cyFdUaUSmD+jw3bX7AHRYmf+sTf31NiDuV51IDkJl3rBi7IuIyLtRscb0x
Gpcbqhmg1evGm21e489vph0wSQFVwum58BhVVU3dMczNBkqXSnbyVN8IOO4dDl9z
/FqOvxVmVc1LRC9mZzDjZbqYd6go+qohaRRBtu7+3xkwd3gw4PUYL4dN+JT0zXPh
pmsm+WqY734lDE6itk/k1UyMApj2BNXwx/DPBwDBiWhwhdOnvrbCRX1RgOXcPy5Z
eAmafzKyhE3nLb8a/sDgxJo8y4+bCWmwW2/jgXdixnOLUu6pZLX1NQyp3KeRO6/u
hhchMCzkAtPUdYeCjftoruoeNHR6PVd+/6tu3lgfM8hZTOUQuqF0TTILQCYXBTIf
QAuXcVFglr5b4pNGlhq6c3qAi05YwcTUSVUMdElx1MxlbCRDnPD4Gzd+JMaWkPMA
DxdSG9nP5gpTwxGwwr1aLDQv5S6vIQEfu+56o9Nv5k698uinpaLKQBTYoD54NUV+
lzTXtmWeJqosaQYgdfmUQHeQ+T/EkyF47aWentjsUi/HtJVItDpRC9G75Vmwx9Ng
eoCeudwb1vRLB2niEW0rtzmR1JY8ofKA+XSVmo8Wu15/29x53Ph6xeibt5ZTJwC7
49wmAOnpY2BUvwaxIbmmk96zFxBRq5mfWHV9nFrcf1mh+nnW7fzkXJ4lEdzfY919
JJoqybgHyzrAgDQZANnVGWSAPsvsGt2E1T0WfB4Uk4iSrGDieBWBbKHBq2UZ5S+X
LUnyP2EBFaFiYzF48vk6uvq8R10yvZEkfGfooQehcB7OWlrzTj3UPZzqUB7mAnRg
8AvbIb7IDjKSxUVxvlxnTzWUXyUVaa1Ntgvg60hD8YKQ+9rY5XpRDlpKubUNJSJr
AeAe48RGurPaAtiqFzK95Md69xWkkUwIIwRDfzBli3eCJkQ/jGtgowlLa7lT2dUk
bTuzN9/2o0V4mwXnxEVszycInggNAjsgRiDWKdtTuxcZh9Png2DrsmrA0VvC5V8x
gt3y78wz3p1XWeFIuPaAdysN8RcrL9ZoACzS5vNu1wwIlmnZh5Og08BgzqNwivw5
vYK1la0wi4T7RhUm2UMdK+Hce+BXM6DjzqRs5rXv2nwoBndxOeMuP8F1abDaJjBo
PIpaWRas/gVmU2/TYAqXzghyxiYbUiLSda9Kk4OA51ELrgGZyCT5B4iCS6JxONSC
aa4QmRiWnAmTSQ+t6H1fJGkpm6RPHEB0PBBrk75AaRWUBSnPQq94T125Ua1M2tmC
vgU/jJxXmSwridnYiiLOSgQ6Iy9YGOnOytMaW4V7crFxaz4QBJ9KXkJDUg8DTX28
60wlLRDGZLAjgovlxySQZJ1nTcO0/wEbqBKQE5MK8BFcl5CsYrhynnLdeIbY/hZT
dogihF1jhTplCiCtQpV4A0QP4C45kgl8MCHQDH0MH1jmrKBGdj55/8E2Sz6scdQu
yqkfGAdbBxFNZ2Sfmr4GRJ/ipTVLR8j7Nw04NFNjs1lLdooSBsL+7nUgJ0xHUOwK
BHlmNotFm5TFFQWI4PTJlsLemf3L/CzMZIe0QljKlTp5JOcbFx2u786e8WQHKpIm
NqqJ+Fna+pCUoqWJ55nifHgdVvTovhauQlGYGWbT//r36h0QXiaFqrEmaRItH4lD
vu3vwKroedH9rT5q2mLE31h2AX/sJmFfpDU61OzGckXYQVu1L/QPqrHxkTS3Fg/8
c550yofSwIY0KXjjt9X1cLjtuW/9jAG+41IUYywBTBF7mcuURPqLS+B9D/YQ2kFX
ktfei1JZNuX3gZNAbaGvApKjnjvEarqioTPGwtstDvGTu9rpfXRxWQcugV5hTrOx
zz7su48QD8RZFJ85HI+diPmcDk1SEYsF5bSoJy4zwAY+KX3c7uEltSnLS/4My4HG
GNYRyw3eAV3r4CIlO3y3/p7DqtYEps8YYSUuucsj+pvcNe0KiRMOR7aaFxqBoJws
WynqvKCoQTgTGmBUlyzAcNFxhyg+8/s9gUiCPekCBmKOv7XHSCxXSUbkZj4Z3PnI
51uCmVLV62MN/g54zsW3OWNgAhxc/y4Sb6WwHunDH6No258rG/fQhIENRgJbCKz1
dM+4uywrB8oIo21tEHilOcnRrQ8vW4IwCkkMUMQsyTRzkoDzF7KIKn9cMFZ/+ZuV
NBspxh88O+EA2xtjx4naEm5SC+Jijd6eN5JYZuCDlgBWTTVGP9cRF+nJxC2enmeT
hU+lUsgn5lEo1J7GLBiEzImonVPqmZjybs98afPmnW3+hKPDT8b3aHS4dBuXQzk6
jomP+/7z4PfUT6T5PxcLZq6rUVLWWeeHXRsjSY55PlUiL+qKllIlbCy7FmXBzBqL
D9KOTVuUT+oFeKFI/n13kYh5dmkixJ7vXxWDybzaXF9CvHPdQJ3NVleTXGqLqg86
ylikOl0aSe8mkaUf6VdxpFw8tRfWJey8qpujx04MvZvL/ZMPbHZ5pwikuuGtCyWR
G1otVS9Uwt/uuyius2cFRO2lbSMxj/fahRpKmeNCHj1GzW1OcPzJD0YpUoukd83/
lqLUaoj8XfeS+2zqRcadAG/i15w28VhhOaB5YfahO56+3+7lut6azfazdQrDB8EM
9G/V40h9MveoSvgcnwS1EIdNiyAmNbyU5XOD05QNi7A7dBfz3tt+ubo88OznAjWC
bn6AUX/GAbzWNphX4EM0qSYoT0BWTD6LcyMNNbsWVGsDv0sOhsUARgi/kmey5UsT
B4b1K1iYEZcLFMaHXsViQwgzv9jb7gwgaltzyKrhelr0zbG+g5bvjPaPy1t96alx
1/H1wYnUWe3ftn9q3F+73xK3T2DlaLBEAZvtWy6YGTnvQcO3Z5aUMp84o0Sxj8cy
RNSyHqCrUl2LwqDk1mXrKJwYtl2Uud9mzha0wxf6WhKwARMwY78gbew68uX9G4EM
lfwRINfYh3bxOifvqnbgTS8q7V6DrTbjs4nGUjwkaA2OxOfFTaGOeP13BczpAe+R
qcp51SxhKrHnikt5gi5FlAfVsX+CHHjB7ZreF5K5gQ9LIX/HQZO587jdI2UeNXvV
CZ1V4hFm6S1Aga0zONWQ9Rkl29EtsWEEbBLoIebzXQHEReC7uXyEz94ztg0YRshi
7Ag65AebeXy7LREg0ED+GHkOKIsxrpOzCnK0TPVpnPZ6MOvPOvB858xlxCNN40NF
jGHci38RgODudQ7kquPsfsa7fcMVif7o4u7A37I9lXOvJfD/dIZaVYqDClggRlaU
nrYlYdPPtZ1YIXMSlPfLEP/sEnQ/xd16BPFiVIHC+ild+doTuikLYnRXjP16M5Ly
84XrMxtcflw/XHL6QLm4s6/+OgTw2I9Hc4B+6CN4E8sAx5BNyhPc3IvtIGT+k+Xh
0k8iKb8bLsYuZ9unoUjAtzIFTuH4L2C99kYTzZGUNeZ/FdKFnnp6VNY4+G9MEw9r
dnXuXCkQEMJH8+OEZ+jCSJvuZuMPB88DrSzUHQyMjDwQG8NUFC9v5G7DpA7ZbXfK
3+kpKpQqNCEONvxEHSuTrqFqlHpW2He+BVCbIiQN/kjLbGDTr8LD836ijH1ovQuN
6hdeEaKDn3fBOTDwOllFC6YRmDxthRhH/FSWw0F2cTNGzptj75xEwNghmAb5ihrX
MOeMyliOlQWPQy/EXv+d6f8tINoBYjjRWPTQgckBBU/WwK/P9AzrEO3IKLJ0Siq8
OMiRL5kbqQVE1+7Msc3qioOdVped9ffKeajqvJ3Tk+C7sguo2sUoDyNPLDvEU1a2
nedJluO+pL/Wh2+by/5cj1MjBYZGXnqGo+J8bP8XAvqs/6tr64xGTHobHlIQJDTM
MltDMl1bUle/C95P3vIQXX8tTr+WDZa7HvgKaFl3lQrCEsM86VfydTgJEYZzTLUc
5k0iNEltrgTejPZNf2l9xjbxadusTEvRpToBPiGq+RRkUVLstt5X0DW8X8Fmw2FW
H3/XfJRqEJ+GzbNdRkeE67YVt1CIQF7b3ozUzMRKMWlEP/Ju1NxBtm9cgNgHgl8f
5jBLlFhGbhhStfJr8ZwBhXaDP7w9qF1pcpUlg04XnwYQkVvo79LhSmOIWMS2dwvy
TGcF+xsEI3lDiOYdRSjvMhXoWSF3FtTTGUt2XrMlyk9uAQkTlfkIsKgNJJ3WL1Hq
1KukroWm0pacPDAAipozyl0a5n/X8p87C9ehysSV9uXoU8yBRYkTHDF3kAXthMUk
Bi2JoN5+jQYjGYO+HyfqzZ5vhMY2gqAyEzvFumIk3dquLe1BKzSPL1wwYgK5mjum
CkezJdgPTn1BH2fQ4B+Na3qYZY2CqsfqELrPSrOUhb3tRnFLUO8i+2QY1Ds5VWhh
b8+NtsFsIIpk/avoXfCVINeG3BD21IThzHTMNy1ODSwAsUeGYLYPGEQTSlnRRv3i
D4oyCNQt8XqzgREdlyAIS5NjKG0ZLnug+2a5ABRqpWp4S9Wkzt36rO6KswNF6u0L
xneP7kShs8doAZE6h6JgCS/cbv85RPrGbvZs5GN8sktoz6Do9/KXxJH2v80JMByK
kebRTszZzkKVJNMnocxm71cljgzczCiXqjNtBrTCH4lTlNn1fDKb8hjvenCQ/T/p
IruW2W2iB1GW/d2j7AwejsNuj2IpzRNHsS3ITg/R5Bx1TiONTqHUPavrW6VsMgmb
ufHgWY1NuK4LGA5fNrwS7aeVcl9gTUGKmnU8gPSRcWQNLt6odQvS095/JT6jq4ai
G6c4gMn4oKn9QFg3xinikQQIOxVly1eEFRIrrhvgmMR1uaRO148QX4brFNQo79ra
Lq/ykEfCy5wE2aPui4z4rK1E6bfc2Q58yvYNhpS/S36ybi9WaCss0LtIrxSaXWu+
K0ae1snqgyx/1q00aArbIZ+Z2f1YN6eWt6oFs2jXZER1qLrZUnWYNkbgRMgV+eFS
zfeNBU/aReGOe/T67vbQgMQnb9BqGUa2h3E0CtqEXlVb9pS7IKpdpBUHJWYYwclV
4+XHqWeRRBpMQAFohKKtrDixV/xkSMSXFajatyRME0qs/6Uk1w8y30PHtKS6IatI
RVD1Sjc0a183xbkLUKV4sTCx9+S7gz84o2/dV7hUSIU7CrqPu06ffNdhmHn24q/o
T+KApJCDihgm1LE1qpZbkVsySjzOr7rclOdRqrOKhMKOWt6tiiNlruBitE/50F6m
tjcxvKuXm7EunwS5UfwIyitDzK3MlbQev93gKW+ly3Td0A3mtKWB6ALWYdFbsA9F
J++IXkYiXKSymA2oFzqfQM7pnaWUrLlKvw4ldO73gdOIN4kk85XzEJ8KJn9Jh7eh
p2YyvQrHcmueJ8pGbNRmm9yp+t4aprra8knz66+xCkfNybBl4iBXJy23LJj7RPLP
L85Fnc+eaWaUIa+LS2GQ+KUqTai9qUXrmXvUI3pdJEPPO5nwUV5CRhQM2T5s67Wt
sePlatXU8QkSQvSfQFGipQAIrduAyGrgqu8xQQ8BfFV48LhjoMazVomysuSy0t4R
a2lTrNYYQGt/mWMqoyrSGH4ZzIxylhEdOW6x3Bp7q9yKsml3tv6CL+OVSOtqHJ2e
cktEd71aK+5+K/GpK9yN3Yd2vAi7nJtOQL0Zrzg3dljHliEsaK6rngNvdhlYv7x1
1EYaXUaFR7PpPJazIqPBNkS2fgmGM8FU5JoLvh56XoUsTlWfO6nNmiMGX8tN3Gaw
YY8PAQrXOK5XciaPtWpjVdyJhymJAamfsiUkvfZqI1lC6Xfa2/AiR0OorcY7XGrw
bYQfRotWNr6GdvBbaAEci7XqsKM26aDVsL0ygVaF6GftyCtArTnEvViidN4M19o/
BTDR/ncAITQ3d+tkGpa5o/VlU+XRatghyvtGcr7FCnokupqhC0HGeyjpJom94Nry
t0qrL1jmky/6/NKRuDirGQwkUUP7bhAGVnjIEz/L7HlQZTsT9XAIa+CEQfO0sMUi
s7fXCV2CMKxcaqZxLkkpuLPDNdRwnNUeuRyJizeGgxT4BagNqDTBmGHdcEh5V0Yh
eafBWd93qL6W2yiT6FJBKCyQFS4QVC26G30KfVP50+j8LnNF5AzeWqJ+F72HsyY4
dPZ5G6Ti7IfEdUKiZFxZfVkt8GxVZt9tLeAFDLpOoQyPOR2mxzyNmAFpg5BLro/u
ueDQJZaIYkq7swLkBkPdVXzZobop2XjXo1hFm0cA/OnNXUznUj4p9J4VkaxMjiQF
Yhwnh08zQx49M2jrN7Pf+zIN5if8p4howtlEcdIrG+x2MdDgPOKhZKa8AIEhyAeF
15HZPBhyNe3WmPiExPgXgGIEXpuBEQholHqJjeIWBifoPM9lLHS6CeFRb8xXAAmR
KXFkYRwNZ2+jp4D62qWiAagylIB6DA7ZgB9A/OM1U83kvArHmBtOcZULflNRG8FG
2JsLK+Na+tHYh0K78QjYtl/Kh13P2siVdy1OI7uvwKzNpQ0GPU8JQsbJpC3g0QU2
wLtYHn0v5WgfcnnKHrs19KiPi5IdJwuba5DdOhF2oXBXF4hbp273yQiZXo6ov4Fy
hS7Cgmk+PHU4OoxWC/2pWI962IiqH6qJyclA2T5ggMvQo5jSW/VG9wY6/+sbY4rS
bJO7qpw25hGtLd0VmlNB88vlSDpU1eZUvUq0nZPMo850yaUpgy6IwS7G9W3qbgVW
WClCQmcU90S3lRAfE0Kk6j6AJR19SvwdCVeHgO+VjdxFXJLbFnWdxXIkz/CYK3Gh
L2kuEWq6nqo79w2FhAUK2VFIdxpfPEaT8mtin++ppgkSwA3f6DqhXuFIKNIlK53E
YMreLOzItHPahaEQKKyRwlF3jKn23wk8LShdBQm8oRA9AWpf+2Kn6/SOBBlzhvFA
I0qV/kVN9eUE+iBJqYl48PAYMEEHzL0hMWAfE+osXwyBMVpFEv2uWLP9/iqDRHp2
KQdWELwT+D5+7/Pkh2OcqG9+beFuzoz9mwjdjaalBPH/0POcnMxjCHywhToSVTfk
BNoj1U5W/XsCQ3JAnS8Iu0FryFlNJuTyQupFFSlMKsfSst9+QmaQh5aHt/1WzcAH
GZKRpYaM/vEK8QjeTq/T8WXSHsIzFgh0TsvgfBJ83WYA1PxCJR4HxI7WMwEb2kO5
bxAroITvm0XFhIv0gltNjusXe/otacDzfXLzw5TbXcIIi/2BHa/Yu30PZu09llx2
kU2t22fL1fexUeq5KUQp1h+Uj9Hky8XgAyQHnL7B2nNlNtXyLLkgD7b2eKvoOySn
boDDiAzLbAOC8H4/ekdU7NO63nsUSZPsD3MMpU5B8/PVnAb59Ax7OymqHELYyKWo
mUUn6Tmc4TODsSh5aAAD3oiYOdGR/mFAvQ313eLgU5bu1rB6yqwXBaExJpuZZY0u
C16zEj8h6cZ8ozHAPahDVz7MrGtp/VqFct3vY/HkoaUsNUc3iiE1b5tdMhgYvI+6
6niZ6hK0UhF9CrmTb+tdN+97t/L2NPQQuu5I8CwJhpQyPSzWyeZhCwpR2W8S3SyP
eoxTbH2U+yQLwWkneBU5FCge1orR2N4pSnTB1MJBlt8MI5Z0lo27HV8BQu8e3ejF
oe2kj7Mbi0dTE0XmI6DKHt+4p6wbI/OnDwOjz4bfN3tmDXqi4QWGwW++3PtMVO+U
mQhvvt/IYjklmy20bhX5qX2uaiUq5gjOnWjjkteHVIEQSKbDX36x9A+jdmLNZ/cg
mTC5RUaJbIQ6AMrC19QDJjDNqq6NjdJvWY2dOY5+1t412lCcZse9Rnvb7M1gE2hP
D4NWZelVDomsSt+ZFsJuQVxy8fW4sib6Fs+i9hDx8nnhy5ujTUpJvlbMzBsOyM0n
LQIrvTT27GSTV4WhO75cZH1/10Oy7g8xx7+YSbe/J1SIVFpzAj3qwnljzUCDSeYP
xPZg+2d1ywW0UrY+zhNI/QAw/Hj2LjMJ5nbJ0N5e/zHAOISueSQ61kvKBB8YYg8I
gMEJXqtJq3C+x/B+vkytWC2j2IjNJ3bCl3zCtGLwNzL8vibzV+LtHl7uU8OQoQJX
PloCPPhVcjjzqQf6Zx+Uf95m87q503kyODilmlXRzizPNUqhmr+v7inlr0IiFOE8
wFsJQDccydOx2LpT/3WfIbo62Aw7QYPxPmTVS4jlWf5Vw1FYt5FUP+nXvHj4V+82
6MTtsnk7NKAzFsh2kZIeHfSYYdmuT3qLCyn7H8HOjEaNb5tXaw/C54wc1JNwxnoV
La7/MpSCxgWq22QZGLMfYMcqDdbfWcUIMKPl+ZL5aJjyqsW8Y1K61qZAdxZmoQHr
shLvKVKilQAprIL6okL5OwOn9XYNTAXYboy4FcNwCxivxB6XG/QlJEBh4qwwTkuA
xzVLbWMCFO410LasJJqa/42arxNqSIODUyxNokQ3t5/RLKWuEs3gLnNfD4eKLdZK
UTh0PEyP8LLc5GkeyAffUJ7x/WH0qUYQ7QzGr2GQQJhgiNRUkh3Djfevticc4jM7
Yy72WID9eZw+ZRAqLDrHimMgN+1SUnRF4PYvC+v6sttWU8nHZ+hbHGIg4k7x9XCS
rOB8+VP1ErHXv2vo1GpTSgpgIZbMzcnkNydN2H1IpIx6+RSxs0lAGHg+XL9V8jOa
wiOT20qtS5dBRd1qxU+KiOU+ulKsjxRqxcLVx7xMdJw2uN8EJIjICJAAP6TvrDF2
bT73kA0gQ/SlgObhPqTxcwUEVIgEQRRLdgvNBB3i6bxhjji6C/dCuruisB7mh3NQ
i9vmlBHGIKLqkSXe/RfxShhbwQAXHsK1tduNp1rhkxhYBn/by9c6+xu//dBHLUGQ
Qx5O1urtNWlbGfeut5B1EvjzI1f3rFnayMt413OMupQ5BzXX0sFQjsxZA8OWtEox
Pq2c+HNQLgt0POzFQFnPpd3PW3Spa06LmD6QB9aM56woUB1AmKrF4+be6XVrRi1s
1BESel4h4iCT/fKcKgGL5hkkoqdfrVFDQ1hElOttQ3v9/q+2X66zHDq1rNkW5xPC
kNkmdnkgGJy0/QBzxdesKGBMOhw9fFJVmXnwtW9U8E3vpv9QoLtwV9st0nLwS9UJ
+lS3DkbcmMyheI3w/ydf6inwgBxRQDgiji8b7a+Q3eMhB7l5ENnsoilgnAfkUd7d
R+CxgPHgamQYaxiIGxZH6AqQDF9dV8b4TMrBCtCWq89GzSIPM4oGnwRwOA0/ukvJ
XtyucVrszi3UcRk/VQ607iFdNo9eXWl2bRUmQtGG2iaGxGMKeXYy1neOLJ1CmW4M
RJAaFso74H2hXg/eRUGC5pRcAeHGL5DmqdqRlMTC40E7Jt1YbAzM1Cstyy2vxyqG
1+eh/NzWZDOfEEd+fiHw7/iSKSkVThzAVkxUElimvKgCDebS//OMN2GgQtR4DvLW
ZP20AkyeRi6nduCiE/UuseftbH68C5m22KrICTdXg6zDHPtXBOA6opmt54MrWwpD
vh36kOwaCZ0MUUQaTK+iJGAZtOV90J2Dq+VaksuXdEXebY/aLNnUBGQRMcxhIIP3
N8Jx2Cv2k3VyusMCHPAz1F9NoTOORpzbNXRsze6IClBHgG6orcNyAstylV9FVL9i
sCKxW8734Q0oUvhxTKMCm7Xq/D0chhA6rL57anNa/o200AWNB6SYCU24dEVj01M6
/oWSzxPW0OE8Xz6wOeeBk6faYOOHvdsuKs+klynf6L0z52pWH6S1kcAxgppXwXpE
x0/DSq+HGHNCvkRNTcxabnSQFymYFsIZkt8aoGTIw8QyUIv23roFKRfxtZeGojWR
2+3UeltA/jwyyjgJfpSnmyyGToGvOZS7AteyDtBO2EuHTa6sH4UQx7mMSFgdHNvM
FK8LmYQnB5DYDxmSSKi/bucsuAIvHyLIEplvRYtBQCKXMXbYsHgHMOMZlDjnU+0h
71xtpRU7o1COqwrD028d5Suib2fjxH5yZVddQa4wZ5jOsF0njZsy7SVR+cth5FX0
fx5FYfEcIU8VmruLYQOclM8aBF/i3hkw2Ps3WcVJJYJcgkvxQncTFCoNEcKFldDS
KfJOOqCLslwEVGwt4xgzIFKxTb0rnlk+GlADLkmWVJPJsJlIUCIouFrBIQn6xqAd
B9sOD75igcXqm+R0/iha8zaf82A8WDd/vreQ+WYANPEBBwryOpK3vj7xFGKaKPkB
r+ogH2Bc//s38fYLIihi2XGd5i9NSUzBvtu6BfGQweiBQfqnLMLcHHR9UWI4gcdY
U22wk4xCKhNSWIPEcMWt4ChscdJygYokPvAaOH8hI+OsNNu0WJT6tRmcHMezIMgy
8SERNIcgR13ot0MdMdWheGbIcvDDRE4PmwUe2YiO/+fEIt25vrdjQWrveSWG8hWi
Cin6Nke4+zC4PO9Wb9pX0wJfyNhqz6fzPzpHqHXMw+X0dFYanR6MlsqRcb/pIbBr
8mK9AMzr59NUvxWrJVGoBlwSMUSd6ullx67rWljp2hT7eEXQYwcvwspVVrLv3IaY
Q0od2/f8dGAnIaEY3e+/Or10pO7ka16/spyi9gyAwB1RCjmaOeq9iMflxfnMm4GJ
lj9PNvtQBtxp0syngTyzSWVYiCWgdHuvNernOrXIpzLQcpLEu7f4lgR6uTmv/i3d
eWhzUuQr1a7hdCJw+soy9mgP8rzAe8LGCiUBxxT7iRvlClrUbQrKSLr98W5V7dDX
lzQz7LV8tr0CJ+eoXIMIHUiyhYtVgw/METVo6IPXkHpq5jq77hHy3Mmztetg+kx5
VPbmd4NMZV2D2XkgXY0g2ROWV8ak5u4VBJQsgn8kcRulEbd7Uho6y0hNBQZWdbAB
oGfxsjPRW3VJ/Wp5CMvPL5jYF8t8Qgx1rTaREiSPSl/c1WRVqFNrCjgP/e1+vPFx
j4t+usoPAGQNsqhxpLqFQeOOcY8s0YPcPUeheHAea6uEIM04Gz7S/dK1W/m4leq9
82xR/0uthIlWqDVJLxXJxzNULQVtoYkKsZmpGRByxB+MsuJIHyPgSgeQRp8XEOxc
yCKZasnOQA4LuiwNvhan9cWCt14gs8I68wjIwLAsOEQtNTSi3TCTGtKndDpllM7U
4ys/5uRabT3E6FMwphATg2lzza4ZUriStHisXsI/S030U+ZCFFe+NEiwzejPgU+u
xHBTk3wqvBeSHowTdB5mVvPFZM7lEh8hNprwbyU0bmVQ/opJVJsORiSyua+YcSMF
N83q5zr+aKMjbJtDuS2v5DZrMLOgSQYL+RMuA9g1AuesBIK3SH0jlhrz24TkzAz1
zzONP/0dNJT91F0q2yq0b/bbQQvp3eR14R8BO5P3+FPfwK1Sn+7jBu+UX/A0Pscw
RM2ffEaelXN7CHqlyAvTQQV1BhHwst0BntJfdaDODJJ+771DVCLkA+NaSw8E/4vX
OwW37NVXVxOw9cIKbfc0WLbCVFwkKSG6/zz3IJ6MIOhnDlwy9s9rI+uKWC5kLe7A
PUnjaPGm/jG3An5hFl30PHlzQoDm5wIIAgIP+JOmRY43blvKHOxgwfIOUoA8WOE9
miDJptqY7zJxmNTMOUqii0llQaZOUg7+JQP955euQ4wxGrzFser4m1oEOVcrZUOD
KNTSR4wRSXp5mQDGNmk6YREvMyZrWWQaSRCKY6ksRruc6NZjogH//IqAtQU8WcKR
ZPAUMFHBCXgJL8T4XQNLwIQEj/V0IBvJth4vqGJ7jEVZL9GpUvam5eWbijzreT95
p6U7PO2zG6NAcqRSzI850uuuzaz2TP5Dqd1ZZnNMD03m4wXhLsMdw/zQjTf/p0K3
LU2dqLfuTOfq/vfFYLyeVlfU7OnKp2qzgnPiAIm4+HZ31YluTyFxO0Mglc/QG5/A
CiYyL/DncfvSjblB/xK7OiF34+hMN3J8zdzx0CakXIm54JVqrDAaHJzy8FYtwzvp
VgG99tr+/xKohVc081HAo68DZe0BsKOov3m/IrNUM3cm0aViw7jbCnCUgv4lfkR/
AW5Iioan+ubD1oRgAWJy8+kXp0sRchg1uqvcfKEZPQmkr8JzV1lk8mi5BCdCQUbo
FWfMwTYeOPqk1XZ9VQZQsEPf2svVdRW13yLbWIxylUjWq8ft8/5F1WZ5+ud3KQnY
t5i74eFJYSaYauGEH1gpaLDyWga/BqRzUbe53WUaTSzTE1cijKQlp5ZkRvXpemp4
oyVy6qtzj+lmVO2n8W+/b9P26UX1zH6gKgaKse9VLTHB1YvWIB2x7PiUlvKLMVtf
+3htLPuGnsc26Tii1SjNHAbjj++3gpSXWjnJmO/kpJrVy5OH3Z+zGofCoL3lrnus
Zyk2iFLhG0DZRfl3nMTR7uyJdfyMsafr7I2aAhYXpODnAc0TooO+re/UM4bNnBPD
19bMJ2X/S/QxG7z7CFN8V1sfw7w4eFFSkduEVACgQ+qam2Q8qQZD3Ipb7Gt3Kss4
XB97YEFshqyIFq4mxlM0yZg07naK4frOOKvb3SPl3ktFseZ0UbsncDNJjy93HGE1
81OpdIE7ODWCA5LH9t271NuP1FhsIfAwOhno4V4NGfGJB9ZYqJnHCd2OFXqX5MzH
1y01n4noilZPPAX5yF63XYTV7SY7zHRsqjD+foxvBaiwrB0utW2NjPaMizcHZIJX
p7gpgL6FAyLzVVS3DcA18FjnYnK5Nn7jQGW4KB49ty7jNLlF+TUeYTvRzwf0SUgx
ocQQ0Yp2NiDGCprYedOxOy9KAFn9NjZZ+zuR5Toy6RW6W1Ll6GsLCx2hE7AHrFiA
BQ+l2zoaavcILhYhiVRd6+QiU4j0M8OljxgVkkBW/UaVMpYR/vNcrCu2k+n2xaV1
FtU57MdJPz4SoXARUKDQ7oCWHBjFGC9Wsrp5qpfF4hBe/S+8IC37FTogLNcW6o7F
kfbeBhQ+9m9NdVQnLaFv/M4/L2x9NdKZcDi/DJcZdA3MGDZ2KDdSC7spoHd94o12
2cTMZEwC/w7wiGGzLmRaDWq4T1r5QndDevXObctlP19IFiMvbybe0mdlU01cVUvl
A94nsCNtCchdSR1DDH05p/7s5OJDr1fFjahYk8FfWRGn6g9SH2Hz+tQ2Ov0OSf9m
VnGNZ1oB63o5VglMzMUwno9JyW52Q1h71S76MTy4LKSc4ALp4GtFMEjb+31WjibF
JVAMdGwpC4fHvXr6eUAHNpulTHXUDPtAJS2hfQPPuiKJT1eYnIS45CRorl3ih7D7
3/qapb4ys31ppKNcO2pS9RnUeRrp0UaESZSAF7jj4LzDbRTpq/DcsT0z4PQr39J9
lmmBKHZwcuw4j+QiIugBHQ7O9FH3LhE5iNNIrwefjaJq5o2x4BOA1EYrQAfESqb1
nPtOCV3J+cr2WY3071wqjjqc6VGuoKxkCwdFPdBRhnHmrtTer4tNktEnomMXteiH
+CYbYCWBUyh9+lkIxd1AESdMX+spBz06kRX5BgaY2EESR0icPXoy28P6qxvnZIo1
/CefF+9mV3kzyvFjvzj7wcULSN+YqtHMUjkvKrzfo5OnR4+euu/vJuqcuFvf5KBW
xXcnQiviBKvQa/7A1LLH2AoGsQKeAQhYlUTaGA6OUrmNnnDbem5n1RszTZxAgEyp
cmf/IPiLWjXiRwPQ69aUvKQ723nHUNae9Jqgzp6/5kj0YsaStCXakeMcXRgBTar7
LfmYXEuAQphrGIHHDwoXKi0ZXAjpO96E+wE3tzqdBeRzOXVki8M79RlIrxv9F2Za
hs4THm5MrtzQ6aptCJa+PWb++P/3f6dQjAEZ0tL+gb1Dnh4zcPp7B10TiZWjvyC4
wvwtwcDhiGekk0MNogX0xfVfkXhkyjeE2omB71oYnc4WPauEiERYzXGCCgCfOYVQ
HY3C2CxY/y3rLSWCmUndGUo9dmUhur1bTprJ1XrwzZkK+37Uq9cxpZVGChbzNHXt
nfupH3ipUDs9tbkV8Xqh8E/8R+01Z4J9AYfiFpjGp84vOi4/n3GUpNzzt5sf1DiZ
8hkhyKGb2yM1+ZKOTCCysG0xGokVQCzo/QrxxvWEX7kju/uqABFTYsTpsHZNfHBr
qeKVOij6+cVrUzfQHFXELS19UFo/uNeVldUFO/gct3h7XOp6TgVRkk7PgwH46kMB
bzwckxqUc+sca2lpVCnqnvkwOLqFYST28i/xHy1Bc/lv/+CLDBH6rJ2mmY40tYop
XB/aFa9tZ4eQexVZSw7WZ0RHWo8LOpAliZKHaM/mSlqXNao1b+qI19yXwaBYEaWA
G9YfXOwerBE3OXffmzL7hg3sFy34h/ISCH0VuLXuon+Y0D3qy9u/3ttN4VkBmekf
ao8uU9uW016jIeNSkArQdjV/rbUt6k4F4TrBE6TdkDzMwH/yhz+RHkyz1oQaJ8pQ
aBpVd/fZN2ee3UGLFyqqEgDO5GQq2ZDVrSgYNYCnKTOqCJfNH523TYzPEL6h/POv
gU01ef07rR40URuKSZ7rHgLswrnqJyfHVRT6DqNhgYjmpvxTI1PVCN0QI+Al/ttA
kb0q3wqKkDdBNFzt5ark0gQ4IFmIzHJe2WC967tue2jE6re6ddkehnRSY3Aw1ekm
eDrf5lxE/SyKmRE0TAT/KgqFBMWfF/pHt3TbcwMDx0e9wZUb6R13zypxaNvIO1LG
rmXNpUgokjUMAPwhdBx7PZWmMPmDP81pfzA79t7eoBvAZNM3S6EK/WG7mory+F/T
9OYgb6orJeI/6Pt8rGTdatYOsaIdigrVYjiVhsRRTZfVS6KJL5vW/kV7PV0MWvWg
NKkhoUlrIexz4adOViHTS/1M9WyljJpDg2/RVOoEa/5ygPdMPqdAFKvDmyPGUsso
pUjFKb+onJl4q2HFdz4+c78e5ZjKTHC6y//76gp4Nc500tCxSqQ8KaFUsVwZyTDa
xQ8ZM0U8TNuwW6BRuykbwa8qovUDUst8Bdw9m1KveFctva6pQUG3wtRp8Tbg0asy
o5scwq8UdUp2eHxo9cHVXLnuos5JC3IrNsMpWUCWumgr0mbx+HxF10CkW25uXgGz
cL4HpDhdKZqUGsekeK00QaKka2FxGSVpX2rUJeLgjzSZ818KHDqlqnF3X1OX8yI3
5CeM3RlETAHezNKoy1k6BrJCSV/qLW3tndmh0Bs/j8qqxdxlQbidqh1dl/+dxY1H
31BrOi2GgA52UQDUXa3UKEm1j874I+smsZBhszcFlG9Ius6pnE26FfXn69wRR/Qz
Ggg/rQHw/k8XO5hUjLbIDJAvzqobbbdAzIWAINjmanhO7fInSqQwW6TkNBKz3oDI
LTQgE57SqOzdlWOxL5EAkamAwXd+pbSpSLr29zeJsaLy44OaDMoCbv8Y7RHA/pLg
JAchmYqmQ3+1a8drrMdGXnU1/gKus8bPl1QsoBe82T95LdrDu0ru0aitHVbZYQ2L
azAG8DK4CYr4Os5pvAD0m8VNOCqtHtYSL25e4fTLhzPE03sABu8K6qjeDIHcRoZZ
SD0hTawyiK0/HNSbmbTaRBxQd/vZtRzuD7BENsAHJgjq/9gCA3FJLo2V+3Qf/EQ1
Ubba1P3ApK7YZSLts2DE7g4+1AFRKkK6CqZQ7yBs/ZMhTnxenjBnXv4gHKTkP7gV
nYTrNLigtlReiJIQ1s9lbR38Srz3WfJc/ooilbhgaeXcM3fvgTM2qSR2+34IDyuD
HTzxyBfFXTkNOUSeEZJS1xDFAxbzlpyaUIRQ1ZKXQMQL1hRxafS2LEqp/wAXo6Vh
g5jjjIRyI6EOxeqxs2UeVhbOSSW2Dp2OE3kYzyWr+WKMdsmQl4LglqZY1q51mNfW
rQmO9vH804v3Hkxk15CdSzkfDD/9qjd5McxGuN68Y2Wd68bQhfzP3VDDlCx90eS9
vZNqXelTDyGkLYtVNjeiyQWOEA+Ph1seru88X8oGRyWs5OLhD3YJExR3MkqASLF4
l7nPh4kjxnIVO3olslIJOljhwIRtSjW8l7luuxaOhC+WjbonF9GRA4Cz5dxYY3Sb
H0kKgSfs9dXuNd2SMTBYyFCj8u83Ey6Z0sQ9OCqvmrGyv9RbzSVZcQqNXICZQM5y
RSq1oKeZNu/Gkiv/OcTWnuzuJVWR9blGOGzVm5G+U9bu+5it8hD8IL5YfrdjOEbs
SoJ4iMy3cTINL60zqTS1CUP6dRJ080eI7Kr8H3TsEZl/bapMaOE+rzVE7cJQdfA9
oaKfHCHDgsfmk5F7yxdS28ftaFMU2p6iPlv4j3rFLY5/JnhAfhMBi9Ij30zG5ppg
qABvVXLKzAEXnHIvzCHh+1R0P1dC66O9IBjhQC2OfjUF3Xi+nBi/WcFoksVXkoGZ
PkhFzjFeuDgRkALj0n3ewoFDfdQz4iKi/7CN3DG13U4o0foOqHMOF7JL8OREE/kC
vALNLehZuF4H/Vak6W38ojsqAwkQTXtPrsb/r1Cnx+vvGukBeAgeyde49xD3jlSA
qU4Pw71tjbRJ0zhbV2PPac7az0xxyaN9xLOld9NhktGKO49giJzzr9ytBvP7uipJ
zh2RdMxWmcwwTkuxptCWqQ7PTcG5AJTlQ0jLlvF+U91d5kmwqetgoCU6R+v/5gKt
6D+Qz5DLmEQ00hPZ703/G3IPEO27PrDRwbJuL3rrg9iPuJjwDuRHXSeTnrOExAFz
rC4x06ywVkggkkmhzfvSCVq6n9UxNTswI18mAUv26DMC1WSp344PnJr2QwwVfADI
IrDl1TKhsWoN2a7t11EXeMU1gn/LzlrFew81tNZMdTkZxJYad/eOBVUqCQp0t9N8
l0djU3ca7u9O8JCkIxrOF6wIVNrfwidO3CqafvAfSgXeQqdi7X6lGLPC3BTafJp2
PQJiwriMsF9BBy1aUK/7xzZ19H4YBsywxZmBKxKqvbchHsbo97bCTCk8XKsuwcih
WNwdZyzOI5W4rb+Qot4kvQkookynRxsHQaML5Vmfa4VnHGbj9yu0S5zoiBURipjp
ayN+m0LIZV052FflBnoneMImN/6Hu9Ev1Vgc3eF/bCA4hT9hvELZs7i+ZADoJE5q
UFxbq0YGqSTqUX3J9ENpNqb7BAxSkTU2PI1Sk6CttgdeNVB9i/XLWwld93DlpxHx
0UcJ8iEgEA/iQg5K/fuAYbWwbGMcZf8JFBJ2Lh5NqQyFE8sWf8SJtQMsFDCg6qK9
2Q/wgjTRb0HHe6jeWjGr879FsxdXZZO5iWlj987ayQx7Phq53TmY7JFcT4NmFvky
hljYbLqxL/qLew0NA1HX5u9r0+LJrsGdujTKUkrAbqY0ix2EZoOta8JZSPJELK0F
ql8gkM1Je/IH/zKSzNTWRzYWOuOB5D8mAw/A1x8TTJ+Sw/2gq8PxsvoDXbrIvQhj
+lYBRKnuofTG/i6QqTZbUPpRSDXV9+LfLZ7O8vCNHo7o3m+dfC0lnvADndlf2HEr
IJg6hjE0k3mhQXPNg5uycX56t+8zd7IMaBzsaMINja5kzg/MgPEP86bZqkPpqHr1
+yMcKtml0Tgugx6QcHm6Ow6z3WzhOR1jx05tL4iX+rdYYhni/5WucSZL/2fUnjDB
/ro3IAA1Q5IFdtt7lUNdOPPsnjN+lfMAiZAlpZ+UN1xLuF+5LLHt5KpAKj9fpBOE
2IZaJNrp46d1AoXBcWdrxFtizhvBl3ZAe6YqU84r35KHX1qNybH5nfxJytjp2ujk
zwCGNQ7MdKmp2wkoIUjzVXhRUcht0tSwhDEPihXLFcsWFT2p6tw5qBC2QcDSlBdh
JE6cbMURZoxpj7kDEm643V4x7Kn79r1zjzlAdGgFdTbzgEr5wII3W8j0GqmJ9UDs
LiN4L1XqP/Z0HVGvJCB3Say2WQ57fgJaSVT+s2689aza2XxojyxF207UKsQ/+a8C
s5naCXTRz1gmZ+UL0bJqQXY0x8BJyxSrwv3836G4XVqj0NhWYPb/wZzoKtx6UQKl
YbMfzF336CtaH8U+GjvA1rBqmptoPkznJKtrO5zS+Uffnooz+MSBOmO2/RYCMqfa
x94hK06VuyR3iC6csa8zkandE0uvsWLFsIj8Dipyl6UnkcZo7Wl7sGyL069UIm9r
pKMAxSuHsb0oBzdMl0xs68Yz70PMLtieMtIogo8eOkxJpySQfaQz9yaIsdJWJT38
xasLNkTAPUCDyOMtQ/cioQODipDJMIuLFrLl/d+II7nCfpy/VtuZojSd4b+32lI3
F60ddkEzmFV/6du3ATAM16eTnptMLLsOr6AoM2x5hm1DKMc6SPB+ILDmZ5IEkp6M
bnx8QpPl32pF3949NRMXKg7wDVqFOZWxjnlNwmfkxhGyGRTodMEMgGi7QaJgOxcP
hDRxOXSz6ZTFM6BSbwWVOaOlxSPnSG7iJhZeCxjNaLmrJXaLI2Q4Kc/b2+GxS2aV
seKq/ueqW8X5Ac2+l7UDZ9BjrS+rsPlRvisUlUtjCgdscyuGYdt3x+ifnR/ic6eq
19gfiA8h9WH1KwkK0OpMb++Mv22cOeyiAIOsEw8JLmLhecEpEOj7RNyls9TvQ7L8
k8jGbpKwhftrKrV1oL/Ed5ZlCRHfAzbCpooAiqptSXSp2uZNRG+OiKkSimwqvnaX
Pgd6bK2Y3Ui+83+JFH48bu2pGVkRWw7XXJ49yRwkoNDSpD71yUDTWul+ftBSSETa
PVM5iA5Zg5jZCYKh+8FhxiE72DfIBEAWvM+7BLKA/TES1Rru5lfu8pWmLBi8oubj
ROUACjSBaYYbivCnvJtSIjdQVtbgMCYkzKqnhK37uQwWr6OQhCgBCMyDJp+ZhF/q
sI1vhmAjgYWRU9/EmKPlim8GkNRbR9ecQsS/pVYs0DGfc6//ghzt8VxaRatlLGhd
AqBpg8yWTcUcfOmRAw9UADGRCvXSvu8yODWPY64TNiDMxws5HMTPttBQUQ6fbjyH
69Bn0/KVMQN7pl6DTsl2DW2/GgO/43HCG2lBAzMN5cZbXEaWpVPUzthLDhB1RGk0
OjRbfPrsSGJVA4frM5YjqAJiDjgux75sFzTR57Q+nBp6isIbPLBPukkrHtOnlW3R
1NicS+yvAmhiCsOqb+/kstBQdjrEa1Nk5CCSpDahULRGWi7KZrGWHvUS7z5uvNyW
rWKGf5gtJa1suKejhz+yZIT2Lt84kNadyiRW8rQU0H7/0ta8hkI4jR+QnEbdF3n/
PCBbu0IMdhCSlOXb0ZvubmV0alwQmZzGpV9jICFysnzTtdkx3Ixl1CqruVmynp9R
KiWxvEqeUbCDVEYS0FPutgJz5651XvWo5Lw5txd0Nc/2mxafYkLR+Q7e8L/kgJDq
n365TBqaoC9i2+ZktoKJqoGoLo/UDrvnjLBRnO8jW7kR7/iLvzPGQk6OId+tBgXn
Lwvma03U61fcpQBlgi2ezg6CCcd4fKCXZj1aaE68F7nSLhAPFep14jNIyXTBulo9
svoaMS3/quP+GkU+ns4TF7t7j00NaogLxCEoCgGhHGdhLnkZaSjw54mwzmCa1g/1
BexgSND5UvsT6xLo5oXq0eTAX99cBh/8W9uu/Lx94cAF8Kfon6bKt/rUSlmDC5Fk
h1Y6BtBo3ndbYMt2iHrqSodfBt3GFQaTMVhLNlZF2wqdM3mzHFYZXDrTadm1mWvN
i/DUN/iW96U5wecj+oaFoi21EuhWYwViwZ1P4LiLu+knV0VIuEBmijMVGC9PsQUa
3Uv4xi2VPQ6lDqcwSMCMh026ebfXhBihdEq2ny+fBy9UndSKNH6zWRyO1gVLMF19
drfyHU6A8vRhB9xfsxUvbqWVhlVrEtEoG979vyAtqNA/yUgKU1ekBO6I58Z5dsmL
gpnwUk9st6cxAMh8zP6J/fjnua+3589TPXhF8XCN0PN5hrOlPyT/K15KMyG8kGgL
V2fZihbTdyF0PjB8dkkuZb3/mhXkkPclOpbu6qzltmfBL5ANTiWkQqGWpqvro6SN
FGcE4HVE9ahZ+1ZntRRR8+Va6LffWbh9xqAK1wdBQQbbwgtqqab+AyjVY1v+khWG
C4L9kwdAf38H25gVE778bUlmB+FbyKpmM4C/qNlUjJW0lMC5iKiLgduB6BkXabRl
kFN19o6gPTNOFPbYWpjcbRBf109B+mwOmeIE+dBNrJVmPOKauTKymb0uShzI2LQz
mDoloXqIzYNtRNiKKC9XkIHUoEagdZRHAaLpbpVh/c8FNAjj/rXqqIP1CC4m0oCT
JXYGv7dYg4pAnHQQqcp6r9JUVGmidfpDVKdX29chRm5VqtDt9cK+TJv3WwKfCz2U
dbmJmnj1+HEqPztcXATv4YvsMkZu4LwIy3ApGgsYq2WXdTJDv4Jrn6c5NjaJKNDi
1j0M9f3A3DbjbWbrSxvT/Ce7LgqdCe1BMtb9VOtyZuOdzNWIPHh92jChL0yo49dc
t3S7vfEAgRIeKxexsyADVG05/abe3CcXBtLhiPn/jP4DmpGhrqWCCUX7772U54YQ
E/fhIe31wug1aUuFjvNjcm62NPZ2GSh7OpZVr0kR/U9EHZ3dZ8TPbX6aK8kYoeGd
qxZW7F3yo8h20TngHVIjy9bgpGbWxIXMcX/Xz0g8h04XgOPf/P4EfpgN4orMz84h
9WKFRgaVD27YljxqCSN1c/se23ScjbmWQuKSv9uA2xyou994siarsTtG6ovP0yWS
9hvMKNcrGembff8s1A2j1vKOE7dU7pkXRxwWU4BKiih7fsqzsjwOMaIhUFTcizvZ
bwH76ZbZs2awQYnbWE8TSpVRXiT4QSswMxO2FHWxTOAtd6AN+o2VGswehPaj55DO
uPi3U8+FKK+O90eCjw8PSpQUPd/2L8ZMVtKmkIvszJt0UcMvt/caDJqWkeAIKP5R
2fQ0L22ulRL9zhqydeQcOUPk3/w5LYD40CwN60b6JfxAt/MoixNGQafgTjmBQEX5
/O5ZJjlkU0QTpGhU5sMjamSHsIR8SlmMUP7y45fbZto2usamcmSZE0tj+x5Ogyib
7q3EGl0m1bnBo5d4EWP0b4hbCqO7rZxBC4agLAw1LOzi+jFmV8zUBRsfZK9AHHaN
p6efBD/af4++ZCDKNbClGWQB7gtoFQOyLFpGua21Gu0c92KInj9FKNk0iJR6V4XU
WgdddFGks5kVobLcNuodufez12bgej3K/etz1+D9dL+/XM0Kg31AVLDD31hFrost
ZnwxTuLyYBWFrsCKC0AOBg5CZB1+RECPgLZqXDJf/2F2/Q+/z4gTY2k+hxSGv25E
GM4lrlemWT3wBG8B2LgvRQBXZBewZrQKRKSs5nzHnkti6J43/W8k9PZalh9gNMIK
F6dlCPLSnX3j/I1eoIcM+eoMGQFAXTTDwEsOJMt0aTYeIlCdSomt9PrP37oCJq8e
Y5IK46Od9O4GH7yikkGDpQo1tg3wmXscLcrQ/wODCltVrQs/0/z6J7PVK1NVSmk8
E9ygyY36Vz+5GspGcZ7UJ+KPId14lXddCE0NsycNqwCl714Vf0NJLjaLCfyTvNLh
V2pm7hJBuCPE6RaEar3fk5JJ8GAzE7sAVRpuC6StRLViNOY3CcTRnSN2DstVNNOr
KycR5bx2lIFlTbIT8zwYcAT2ZdCxRLfIIi8i+BOmxZd5n0ivAsaBlX9TboiFjxPz
bzG5dIwvmdlm/f7YXv+DsigNS5q8x86dOLygtYbApyX3YKKCj/BeSoQOS4ATovTd
HrYVKrJokKmpimnMlNkH/Wx8za9rFtbctZ5G/rxhd4kA+jvoMRagptYhFvkKg1Yx
E6bfaHLJCNwAMRU9PZTEV1NM+tWLpoit4RcmEVwLGzAT7TWGLhzclj1w3yEpj3ar
YxgfZ1/S6rg4N76zqPDdBC7jtr5wcUpkR6tIJarYAfhTB6flsLS3GosZEBnAG957
LsBmg8qs3RngVzqiOwHRpDcjrtcY74DGSe0MdqkmChTCJmOZkI0/EA3HVdUrzOK5
DFxg26BvkMryTybVSjpK/kEF5YaZnoY+EnZT7hf1lXc3TzF7VtY31hqRDO75SOmc
7CY8ozX/CxwRATNyRsOU0mWgLftm7FygK370QkT/KCla0AiKDhorfKivpRGC6wQr
vFQ2v/SL101q1M5PotTi0gnessgEgC47bGbZC5F11NZ3rb9GIBSOEimx59cHR9Qy
uTCy2UOzYWEl9vOrdaxQ+ppUXfuKkXmZLxLo1V7Bi37FPCG2IxYMB/63g90iK4KZ
lk64y+lHzxE4t7WWcaBg0B+Z62bHMP3TJCjwo4kAhpo8G0B/FRJ5g3b0XeNXlaN0
izO7nzH6Ql5Chj08LtPaL2tDMUgPVHf+767Bx5CnkY0Toxsy3WofGSw/qofuEsCP
kW/s+I1R95mbZMcbsYJGrkrDxlOpUAkM93T/o/7/tSs3icldKyltlAzBjll664SI
OcE1Edvtl+/Z6F7ejQU7xIPbj5U1A33aKXV2Ax2ThknghjBxV1BGNw1qIrBKv1vw
HPuL/jQePmfFjJN0B2wNzra2+3epeaLP6MOKN1ykpGzanhlkVHVHM734F/kzxTIn
KM7UKR6AyVmuft6dGVAkUMAtQBR6IzImsdEJB4RFwriRmtzwE0ok6Pp7hJyH/3qS
XRPbIRhgwlnQJMv+V/NP+DkuWghHr4reAKDdgY2ksO9KJJBx1MaQ0tp6tt5jv6D8
12Lu8fxQgceZxAInSJYYHWv/xHOHBEihvpmwkaC1vhEM/+E4u+a65rox55iuEP/Y
olW946XmyutJFmNoywUpapevY3xr7smu3paAEdeDsQUrOaDo/c9QCC6L5LO8ZIHc
sRweeCwv3Ci+YmUzaoIQaZseMUcDj+L5PVlVa0huuBJ1u+dPS+VAYuz1Hv6riM5b
PsUYg/3K5Apf46v74euQMqE+4OJmfww7EGLqVcmdskeiugqSkpkYb6/GNoGrLnrU
H0nk94Gm3Abd5b36RtKECvvodZMJgbaLlj1MGoFMbyn/hI2dL03zGQFrEqZm8u/R
zJzZWCdsnxHKpT68ickFrKx0TWG8VEHUoMREkZKCxLMOpY4TIBjeodnq/MmTyIAY
bBoLYtSDZXHbxqwkOOnaXk24N6/Pbb7fac/m2jahaJsLf6NL+Qzm8C9DQvnRww0c
FqXz6VIyUMzBXaRfVioOLdNcJIfjqFDEfCJXistHYVpbsD4xdVV2Dh68h4IgBdon
CjGUE+wCMbFanTiTApJoESh6phqiJ4YKd5kL/w5vX+4EVF3gPyaDikbJUiU927iJ
LKBTfuThUcMnrybxP6EHqME9Vz0FyzjIGaB2Hs8ldPi7OoEa4dItqeiDrLOi3XnP
oG27UhVSLNnRt8j1nAe6iTuNlsFCQtNTGx1NLDWXXU2N4ZZovZP67bmkpTJHsw3e
+IkaPF+TIDKt8iP8UAL92j7LWtSqkixAHwy+jOrYo6BDILxCK4vJ7jiwPtQpZdhZ
7LIfK3X3S2oaMEteeovi06xt/mznBxdtiR6HO8H4Y+immN6zoq+b8ZxnxmK7ZFM1
HIBmVB/i/smNdw5Dv/k1r/CBLmBMQx8wgINZ0HgrBd1sXGGmzmzO+8Uu5WBW23mm
3gturN9QnR975Oz9VHUSni8lcfrGBfKU/Zill4XzefX/EaTklreW8zKf2UCXLSi6
Y9c3TLqsQN1a8s/+5f6Khrd7XyfUoGVhnpPIHCDfEXI6oc2b1IHF3U3az4abEz9t
eWFqumD4UK2WL4jY5WMvhcxe+eDFsXt66dvtnA6G0ztkJDw+yB1imCZ1mK6nsu3S
1unHHdSaAcx+OqShuWUSfY0u/58ui46uSdnVTFJKe4O9TNWA9h9k6NUdpvfsZ9xj
CXqnPotymbfkueRrfeabVx+AT0FNUFnW1Vnk4MJT4tOUjDzaWFWqPO6lWtFZUt+M
sYMl8tnXX1y0m0OQMMWsBWlVzLVWI0PYwCsC6GlYHqz/AUZhFxWAqQVSXHiIA+/1
BkXCh3PJyo51OuOWbNO+mhhXh8XzHUYbn4pTe9pkm9aK7t9GWV3S5METL5Nq9Eky
NTnfTX9UnR1ch9GpOYGMBd9Pd4r2D52RXcnSi2yXaUgZQke3jNkylrOk5tP+1vbP
29TqHf1U62KzEJkcENsNA705t03+E0jGLl7+9uY1n3eJBJT+xKT12xmvaIvyqeUk
XUe7Vi+vueMEbAqtWfCQEP2G7BfEklNB3dAYzHrVA2IVEbgjL9fdYAFKIjYWBeUY
VPF6zOIEzw0JASXQpOuRAEXB5XLyXAZjCxQg8vArv2Us1zIO+mMBjinxGIXi61mK
e6c260sAzi+8UY4CPiKGxMaeRi6G4CHDQG/znl2V/dJjXwls2JFCin1o0vL7thIX
1pjuo8cVeizZQp65zll8fRlbQp4weCGrVF3GIFJPJqlq1TloyFDVmLKHtQdWTE3A
3w4OI0quW3CX+vGxOfUq3zQBRw5aZNlIyPnsN7qxIhFw8L7WgTYXtBeWv7+R9wWD
55x1w9nsxAWS/DybBPA1wHsuKG5VbSR/g4MH/9Xo6OAeV+++FRHOY9csnJi2am/7
wmMm0zAjAB2x/LoxEz9WsvPkea0jjccDOB/xtHMTgjEQO7Ca6ruCKaJFc/toYhAL
mVzUszTJcQYVaP1cBb3jHzVNeTfwQrCLlku+OstQSV2JdPvuqvrNThvjTpg5z8pD
z15fydCFp0bxFrnsX9cPBc9N2XYU+qD+CVDiPB98lrMJWX/Ltn2QQchr01XfZwmP
UMA1jK2mcZCa6NsP1b5SvaHa3HchM2W2Hzwitgsg3v9tJnt1N/6UFBT7yEZNkuHJ
b1uvWQ8mt6KwkNpUVjlb/QU7Uoix6dtG6qQUeGKSg/g6DX1JtBFyZ6YXd+tq+o4T
FdtkfjXUeDJR1N1gHJpALqlEyS2TMmjgrngD412g5k7+Jl4j5sxfoyquGhyUtSoy
PZQsnYxxuc0QCXyRBhqtFaFSOGDEQvUObC0tpWInaZCYu7zh2IX5R/p/2rN2v1kP
4wQje5R11oshFBBhajpfsIdEarABRlLEdO3XQnIT03M0iGvW6GCxKFjDii6xEVRi
ZhNKoRwVC+2UPENE4vwuyo0k/pjdWm3wosDphy2iCWetZbCJ0MCVn6zLWg4GnJYz
KC5izeVjwd/MDI8K9p7u7gF/VmDHFZeNrSSSnsTFnJG1+ucCoPcOPp265RatsEK/
gc25Y0Qy6t50F3wKsdrlIsNJA+B/vKsiPtvnqofl8HKo0YOmfQItanTnJXzaQ8Wq
LnX2f8J3YQ3rA6N8tjGyM9OBkDqS1EIApSQbkrAdMqwUDqqsJ18IDc7ZVpYU0ic7
Xyoz4H1jKrOyXGGFWZ2///1HrDY2+Iuc4pj50OHuN3v4cDdwpHISJk3u0ql7zlvQ
VxnO2Vw3M0TM2vAsArBe6kfbfo11nwOZ1Ogq5GQDsKLgeXotZipaaMg9HAHnnY4R
eJLFtdS9fmXkolcXu9hjMQmzMnz1fW/bdBnWU0fHuXp3RXeMRhUEsCBL5mSqpmqG
jT63AWG95rpVfSlnJ3VhPDYyj1SeW6Tlnq8Bx3FNrNdrj/NGUAKOJ4H9JYWpYHeI
yQS53RoG60D0EF2cnb3cTcKyFntfKOXOq0Haw9R3gKkjoWETytvz5TGlIMyIgCfS
yIZXMPrihSqmScOFFucwxmesEeYD9fXfqbdSFte/mszFDscqadg8jEGaq9ewY2Un
bTWitSisVVkCyorchsbHv0ny0WnDp7HvV+2jH6K2xPY/TNAPpOruLjQpIHO9Br4e
/Xr4EwnHmMhk1mt50/70FjrIv6CmBgPGspCQQZLIA4HKS5vt9iO3QSCTkC2jVhQq
w1S01eKRBh6B+6NEDVMf0VMZ7C/bO5J/EUnkcSO9MyeU59jqe70IZC8UTtMKVQ36
GzlqKmh3J+B0fYjq2MIyL+f1UVngbzAPlKaDoXbg4ZxqPzPbzkDDvwnxt5SwhhDh
GYfLrvvlNVv0XwMC77Yj1A53SRrcOWexelgxXbgSo28FtAKkha1nlu7igfHV2WLe
ja1ymZj41VsA5HVhaKHsdeFMqWaDxviCQrm8r+M6s5x3+aJL8oSh9uWqocyjChWT
N0qZU0ei9hCPmQniZwNNZQCPf5R9hNkSdXJxth7/wcgXJRPEyrKAIIdWwGnVRarx
1o3OIyQ6fCE3jr+2G9N5PduL2Iohvb++uP7QthzXayauwis/VPGPH6Dt2N2gw5oa
LG1Xel6k8Xrc/JvHFwSGRjU+Hn5+aH0Qb8JLi1fYNdjqFIGBSpl3fSlqmilfUJ95
Q7TkQOPdPwZL8qP5PyjoFIKuEBYdpRoKYW4I4LShaIRyNtEuTm1PrXPuKVvMOmZY
CBfOE2PdiP3qNwdpGjRYBgn2bZnQJ65GPK1NbxXSZlqkl4hThv1LM4Dij41krZBm
CxSMgTA9OBVNh9PzadOIoPWuJ6HwOQ59318KSPvxBr9GjGd6qJ+SlH6bWhG/4dOW
ygZosc8gTl8ihkIaRaeS8dpYthGpeSf5CVSBRQI/UUoUqxbF5NRvFeVmfo5O/0Hi
XF7vkLCB3n+yGPy4dKVKuYeVOYvCIj3hzV/zR1n+jwr6zn95RxO3E8Rcdo03nXmC
DQRBHr4P2/4I0MJ116mzCFgYu9dEQeT5BQHOnChMo5j8tK76+91Fcr2zxnpwJ22Q
1GpFqdY4RigXlSwgyD0KldMukXJTVDLMIprzjC+XuTq95jNbHuKGS5N8UTNB8PvH
tKyGJ9Wh2FMlcTFPhMxxQMx7YPiuWF7ovrs51VXpaw1zN0vb4KuSl+hiRXjsSwYb
QahAgrrUVXsYpM6aTe+1u71ehqozinIufiT10ZCie0WlBpTAkBzQcIq2JixFLcP0
LpE0b2sXCGIJkKC/uj8xAO177Ehg8hH74DcYZuvMxxuEDB6UuaVk6grGbOKe+Nn2
SuucS4Ih/BEC2x0UTfYfGfbkqka/xqxS7C4UOWLVMBjQvXfKyBGVPzEMvbV8rAtl
vecXsUSlNvCaiN/GX86jpwlZfjAdks2rqcd410zm/RIZh7EkOAddKLdhd2rDbeB+
VLVLPOwNNMPe81DHM62pd+gMRxg+/wFKnI+qxhAsyA1yPJFZjT3tfy8jcZZJvO8Z
vuCG5ABSFVoAreos+P4ZRalM5LN6qRu/RQzrsEWcgkBcr7IgGIpeLsU8MhUNbNOq
SJD28k0pbJEGpJNTEIdv6fusCWHtkFihR+iUIjTVxM7bP2XNUJx+qE/mRXXw/kpS
6OBEUhUJd92plfgk7vs/jAUuNgi5Cyb1S3nbEu5VMU9smYaBQPX6+36SFBJ2PdzX
hTrbhkWPUOOJH+Js+RK1Yx9ucWedAkXTYpQAr+IUSiTe01kHFF20f8SdHB1Q7rE6
5WkggMK+3/q9mKc/DTIyYR97WLGccAeH7LD2HMerFSyJt2L7HmaPLKk69SYNQftP
lEDsaGrwSa8c9B+qeWpM/t6c3YUQLcjaYaAnEGSyXwThQcAG8dG7yNjo6m6z0y7U
UMepE61L1O21EgYb4yu2Zag7CmNB/XDezSIuDdv4zcdX6kKEaCsQL09/dPM6bsrx
cP0CYOhS+2Cbqki3tBdH+KfRp4wWbMB8OZlMnUNwEscDVO/4n3H8xKD3vKq5zNEl
oYUnF5zLL7L58NSSzPL3sDUM65Selypfi4N7RMMim7/XbRSYSogvCAiwK9mFNP5U
2uW0voFr8JIJdtiUBNdXxmdo1PQY/UjoSdVWXrH519d9HDbki3nzGxDwDBj5Kt4U
o+xor7JoyIcnXWBFCnufmmxKvWO2k/mz0PNr8vsOWKi4JuPTYr2T82EDXZrCsL+P
7mrMuDgx9iRCjiKYIYYs8qGdRQlgDLwiV4tuDhWB9GmzisV1ze+52WdA1pykfJbT
b8GEbKJ6AjQgsboHUs3+2E8niWvIXJDGdjpk/SdMlSAvwO3xOGu9TWX6IsF/sIJc
8+WQaKHOpypT/5jJJA+ZXXLVNmN631XCGPRkKt81RiuGm48Dl9dNRpM67eJTMwBg
J2p76SoRptttj8fMMtFipPZnxlH16WkZ3KEG/4KWXj2ovY9oGO5YIela2xU6ITAf
GQikYKlCG7UFszIeTa8bLVo4cIEn+eb+Q0tQXqfMij8eoAx+O5C7BZIVAnRpElax
deJmha446piADUUySTHqBuhXWcokV82y9XIhNmVHEIISrRlVkuZWZchtoJ7r7WP3
j/+9U4XmzX7OxSAIN8AKhxY1fK0KM9LXzjW8XpJwp4KmkjSF7UpzfBUZHe3V+hqi
PUwu+b8XNQ7lr6aV9MNkBwp9XSF35sM/5sWaVBby5Wp8mPRLE/sHvDZuh7xagJIk
/6cRSYNP2FYJvjJYEAHK5u+ddqOZzyTlgwVPpyIa1cZbam3u3CjXuo7hxf4mGOeT
K0NmmOVJj3n4EIkMpGb4Ej+eitrntJzoP/ZpsNOio5eOE2lhemvRw90GCCElQMHD
ggLkdGnHKuuSBXuRiryChw+oYIycJOZAV57+uPvcPCWNVrL1/0enoBG1lj5HSfVw
FfF4Ajl0mCfQ7oRTaGVq+7hDKPce4KnCbWe23wo5vQjRyOc5P9dc2xvmB++gNfAm
O2mwiQJmoCriON3PoVIUMgnbDSOnUk0aGha0dmaXWV8GS7wSjnOuP4R8N1m5t9PH
m/TtN/ZTBDwkjGRzRh5TKtmKrFiV8kLx0nJb7Efpxi9vU7tRIKeOo5V0Uy6YWRSE
7PLhOvnhpKuzsd/nFl6EPyzWvFqq1DYOlb2eAX1HHtKigox4MC0Zqgrr9sbqWqsY
z4/+xsFxNq0n75AY5VSe96ZYdkzaMro/iQS2rbXjJBMqGpxkUBtRGI6JiD6km8DA
uBQa644rpMIkII18tmimlhorXFf9MfjQiWKQQSzRYhqRAQTRQ/FK7TqYUGVv+7eM
24GoKe1YZp4NDj/KO72UG9SrGBFvdKiNTXmM2eA38LtansXM1eG7dOqRIGxXYb3G
e81d3mxlZ/55F8lBeiJ0ntw7u6HBATyTHmJvtdCzvKqOSY84r1RtUSAA1Hxi7lHQ
FEklxPfPI7N9zAasHr9bcM2VbtHH5Kzfa7d6epreyMqt67tfg2FsE4AGZ0Feo3qo
Zc1QY9sMXvz8j8BNXT+50XRkv5vEEE/+HSeb+sOJWOdf1yRJhsu4/Ie7TFDbdhIF
grKMi64h/2yiLvkrmZkXMVPauWjv3tjZC0Lxz1kM8kNUbIHHEDSDcUVdfAHDUH5J
kLvyFa/PeTXyp8KJHEyyKswf4j0kcQKXx3lU2Ue8MafJEpbaCCsGhoBv1uUPcOJX
mPaKsv4pKT4Z4aSvGR4LhsjGwDpL+4gx03OoZBoMvSeK+x2hrHJKSWyCvR03gNAd
W1lHYpSjjguqaKIhgnneUR4p3QBZCKjcoRonN/p7JfGzrs+hEN7sP1w2kcTFCYw3
x8sDXRhLIErW3QU4nS+f2QqXJoLmTMJ5lRqId6oRh4lz/ox9m6XBDsEl6WvfCEyC
1UdJV/0c1Vz7MIIT2/6LsXjM5iC6gw9MseOqghHFg9xSrKqLPtsp2Qu7EBICEvoW
z5gZXtjMTZeBdESjdOXKmcp+AWlEyHfgj0LthO9Ze1PXPQld8OTXLr543BjFwmCJ
geKRe8y35JoxZF4G65aaubTYXujHsyaIehsn2gHOv2Y9Sl6YpcKn7BLqQBjqAHY0
kHd3sVrTnqT5zUDlElpGCFiCVr9SghhNtn5YmM6FhB1SVF/hW3iCAeu22jsvP9Mq
szxJG8mlytdcHvS1WmSeEWKC42RxyCPmD0eLNP2YPtvS2Z7p07rWwuYPhruJbMuZ
s6twNUF2r3j9fCLqVAiiySZBSy6osZKqqmQ5qWVDXbdwft5qJaSTKCUsCXA9QnoN
9/Vjo2Uo4knOvsoG5V54etKzSRQSsGWBsK2zpWae+o2ACetGnANS9esKBelZjytf
I3uHsAab/gb3xvM08SwxCV5mtwNvrIu/46JiUaEXvUKyU0N9tV2aiqabGEwDikIk
ELZ6VsV8lVYBW8iXxKnfh/COxb5rt06YmTWlYwmuotNTP4ucLlP2T5xx7jhIWZaC
6c6LIM6L8Xg3Bjk4hVjfYzMzEXWXU5hzYJPFRWceLcxGUe2nhk6N43FJ9scDJhHA
fEog8giJ6Ck04x8/25VFESdKYoNTyl/VljLjxIx/zEZR3eYxA0knquVJSoYDKrfh
XM7O7aDMaiPNoZkLEGIwHCOf9IC9ch7Lz8X0XKPF5iR6g+2fv2DT52t3OQzgpZc8
+B7OomyMGtQLdrxcYoHt1+kSj8AqOhHXQK/7ORC8dPLXSpVVefoGm4AFq/2Nyx/o
QhXxt6Gv3uq/+HPcZVVds3C4ij9DG3XJdWA9Q4R5Sp/nElWc7NQqKvMYSM5mDMB3
V5fdSuxKUeTfE2IQ+Yl1GOP/rl8la6lbLpScmUcWHOmTS4d+iH94awAVd/XckEIP
+/JgI+etQnmw9SP15WL7efwgBOHZvNj+AWQdKDcKTOXG8V7ry9w92PfyOPkYns5Y
K0M3uTSMvxdEv9tGGq3nQeHr+L8SKd8harVBZL//Uw2FrAuXERvfUSq1NMgF/Zfm
08fvdZQIdIKT7ovbOwfkm/yyb2dlTsXcL0/9JxvJElJLKzK70r8rIW0mIcNTpf+g
JYVk5Zxy87Id08sU2DpgLtFjCfFNJQcV1qh6ZO7HSjufMXa+zQ3kOLYdAdCV3ThQ
SPEoxeivs74nsSWbTYcJDUwdy3O8tv/Phn7V462vmBff/ao/N98KvI8599r46UYt
tv67Pe0B1eGC4qsMNFkjR05bDn1YvdoeCV0eFKfTYsXGQW/d0o1ZXNVmPkXwUZDN
dzZExDsFHzoYQieH7xoof2Lh2NJRpVfNio43G3tW5d5LOUh4SuWSQCcQMrTxZPL6
ym0yAYy4QUyTen383TcvIsQHKFXA71xxS5an2Blq7MUvdN6RE+vaJW/imayiUIQz
/LlwjndXxGD7emnR9DDF9aIjEYpXiFo+d5LSO7k+a2RusaeknfQ6UeTBXXVM4UOm
qpbbxRPQf++noJQCikP36Ldyp2+Ko3gzj8k/2aPXGRg9TE1h8i9hqmij/LyMdUIk
4T5PTtTkdbbmdrOezAm429PNY+Dp0h1u1VrNz300Quzd1uJiYmjuHb8Z5Du+u/y2
Tat6Y7OgMUa+GW0ZcOKyvtMGr+FCewclx4/enuf0ZLEee7mNVbqd72/7bvMRL4Bu
PptI9041pnOUblNYqVgoyD/ZoulDJJasHtencX2b5UJnbgb9uo/2yRHv8sUMb5HV
B3JMhz20m8hw7GIQ7/lrxqSk2G4FTFQtPpdtC69pzSXPWakaRvq/GWEneDR63nPK
bOzBRWSiR5O5J3K5AgpsXBAPmaGcwtTJqCxfhGQrdP9Wyala9gw0dNi5mSYNdBTz
JVhQbRxiFb7YGvFZCx1O07JYXX8X4/4XZWZkKA+X06pRRRMPZvmqTsWywZLvj22N
Pniq48r65UscfiOIj5Mut4NogTFIvnpWivnZPXFByiA/ZxoFtDTSdGLzTqOIj+2M
28LoOzXQspzZ7+pnkqi0fdL1ovkbxFlCKOu6sj3nExRsIANQGKXyARzhte+v0rG0
oDTklW1N2Vg0DSb3uofYwA2fWf/52yZSMQj6gGMOcIrEfKyJnBGSJgoVGn2XaFZZ
UcdwuqfgqpyS/n7eHz4vQhraEXoq7KXg+JeKReUN1i+9WnG0VrZaFPN652J3N1iq
SvL6EkOdcrGMmvUHgG1nmGIkdrc1e/SHAcXB0PVBavXNh3BJKlqffaRqzAhvmw/e
4QFQ1hdEnv+VKtjsqEadClC1BtA3a/qY0yty2mmipkodnmlJ9/YCVrVfkIpd/7Mc
yEHMha78sgYzC1gsMagy/XV0XpUvM5vtTjzhQz7LSxwuenWnRBTrKsR0USFHUKIT
2O/VRLH8FNpRl0Ub1tUtMb1poz99HCDEQqhGprzEQ2PIGPAwAMULifIvEGhlSquR
n7TdhvK0XN3Vq+UVlnowF3wxeYC5wunuhzvrhJqi2mdyngMpZrJjL5wBfvqwwbOl
rW7FsgRxI2FkQFpomFQcNMfVZHTKPQI4lgsILYBdp2iLY8LtaZG1Vn1YyiCSGP5b
eDkgeXTkJf3JZGQuDc65zsDEWufpCpGYBuHZ9zyjkYJsVhKHzDujJ+mZALjIRjub
6BGi5GU8bqa1JkCoVcxp9ufa6uNN270j7YoVbrOr2ORGnoJpdF0rjtlc2JEZBafI
yPmf5MZPa9+CmDQ8WxUjdNXPY/4ZVGYKiX9aotqxXmZ9CRySmEBaF8ZlJmsrejxX
uU+0Joksw52wwBbOsOrCsWoArka/QGRvP5i746qiaH84sFJjAXPJhL918+tCSoiI
2R0AyYTGPHUKh9Fgcb1KE+e2WtWfPil3/2UOcW0bg1zwfh7+lGzpPNu5ZMz6IjEM
CBnl/QFgCdUqLhPRNsGoEhduM6PNww9KG+oBZ+5xBwAjkpKHHKWR5WFVXy1oxcfI
x4qkjXUKIelT/+74bQ0ot6qZomclZ7WCkqEigRGGNbHfLEKX5ng/dibNmzBo3pQ6
hXxdsTx1RsSNnS84TXfUl5iVen01XNoVXcHmDm0bcA6lMXGs5CpU17b1J6LCJP0M
EJnRuZPnTCuuuvPkbDKEGirrvXjSa6BH/rUtupVg1seudGn/7tRDOaYDa1xVioWJ
IV/4Sr2U/M5SXcUonsNrQHnaNUGRGyxE5gm/ZoJpprnltyIAV4OSllxg00CUNPzv
ycamKCfMS4E+qAoyqp+HAkcsO51+Cin0o6yfOw2LcxU3RUj/xYVe6Sz2OX/paEAp
4Ls1okqFxFsT7ev+UXmds2Obs8LfH/OvUnn4K6upXNptIJnSWBpcqf2NDKAfgZld
xZD+tEB7oLNrLzDw+eVSvCCgePpYmgkzGgVCPw+oNmvoKm7LhWphsFDlEhmvOgCq
RIUqwLaIHz/Z5GsiruMZv7RHw24dJceEso8GUbdErUZsX8z0NtcG0EkelxyA6OjJ
hDhduDqoijGShkfvQE+nwCRjlIWR1rDmbgwOyCdPDhXmVaDM/BO/CVW2urc3kbW4
7WgI2La++vVbQnXa1KOfRmPYrkjTIuhs05CKUmSYKrJnh/Ghe3Em6JH1hvRoAXPI
U5yv/ighq80rgM7PuMb8O5cbrDsdW40Z1gfzjcrjb6zx3B3hec0MztnTgnEFCvbz
xPBr8qJnXSozywcRBIFSviHlrXIn43L2IW3f9qSHFXeoIAZGpdc5FjpE/iOwmN/H
b4YiFlK+TjhTiPUGi9OtgNjSI5sbA2Q+/tpNdWke0W4zMDYygw0e385Ho/VoBATT
V+/LQJP5gFgFhwd0Dj1SIGG7e4O1e/SnTHiyIjsm1XyjblmjZ7IhkQLKuac7/3JK
o5wFQVzd3l3FboUpYpMeqKABWO8Ttg4fSu9kl0Ja2VcsLarO3GkVVUhZPai+uVGK
KSbJBqaSoka3LnTwoWpjolYWrCVzBFiMob+c22OXmvHlMVHuSIa2QzlR7wNru5/5
XTzRxW5ikp2rGfBa0HZMRcqhcRhUsXcYObFiJazEIOaaz878TWw3rAFPGpcOEvuU
kS424LOeyz2updbVrxRjaabIM1wtd+OY3c2hOzR6O+Y1uQO+KlaDKeAmX1hL5iOp
rAuuInjoTPTztIShWXoEAlI7fPTqLOCXJjdnCCpIgWEZoZt8Nmw5id3MMLNaywVJ
0DJTVIEQnobkSoNCfEqjeVc3a7PyFVNlmlkW1OfDJVdHU/C17pN4FS5pAsJd0cXG
dC3tUekAr6Cr8CJf4CaYegV/q2v7bJOxgzdr8zpWoD8Z/KqCm1W8Dj2PdZLx9Qrs
DyS6xmubwgpn4BZlvT5mDE6ntINJXoA3cNwTthenlXeGtvDM6jqvh+zKGaN5owOk
6BtcQTzlaruKahN/4d/C26VZXf8Fx0iHpDAOiJbWKhn7xwI18cJhcQYTnxyQ0tmc
Eg3WDGk67ZDWRv4w6FEKxJXwuWRnLwdMaSTZ0qdrd/04NExiStSEu/tk50KI08eh
G42hRE0x8aysdPJWQNuVEyIgB4kSaas2/M80ftoomJ1YB7TJFyntzxntU2rKI7Ac
lpfdbtoToQoOByVYGQVFpCp++GOyMs3/ZKUcoWEecWGJYApFs3Rhph7WKv4We1EQ
xpAAeGtKmAwTHY8ILbIX8Zc9YtJLvdTDwwDEHC6T6qjhuVJ+rjSbXdZ/qN4ow0Z3
nEhqF4w4jKcchusSCfYqyhx7X7VuOrOuhtZ2ey3I/omMbBZoYe4c6OtoDSwmRSwj
lsGHehWQHVTRfa4EdGcs05ImdZM/evdi+lKlC5PYVFLAa5mqXBtiEpnxSNBQ54l8
przEaTIgj3UF1nsSxt6Mu0TfqtdFjM3w8QirUINmyzeHrRM8pgG2p+L++JBOgrkC
lMuRDYW1ye713SUiNRTMSu3xYxCi9MdtuWj1Jzok1RgQdmW2Qy5oelMorFqa4IFv
AvrchhI+yN6F3/KfEuxjBFP4biTXDsFFlbqZMzjWtG7vWbPPCsYlW332pN/FoG74
2byg5QPn5PphNFG5MbvSK04j0ucHwVig1jJiBWOFd4YWneNziF66LfAeexlq6v+c
XjFn+b+se/NKvx8fpX9rSevfDnatQemdmaDomVO0gC7k8tgjRmkruZznGQEun9dL
Zk9PstUJ+fgoZkSzgEWV3p1BPi+hV1UoEivMDYzVdywh9iViPd5v15KMw/ymQ2AS
0OYdaJArCNLcX+H5bo3FVthhXkK216lPc5jFXT9q3x1gTbId9HItrLmHWk1RBKnX
Btp2PA67sRx5vhUC+OzaWH6PaKb3agUNPMGuFD3fgkam/QRTtUOQDn9Vglmn64lR
hy8wnuVcWBJP7VVZfuck2MaO5+QTGbVALCf0E+DWvUUmQUR6V0Zf4Vm9NUFP3/Nz
VTCAPnzVnakb747pTS0YxRqppkuIPBiJeSh1bCuUCxjpz+mFUaXXjhV7tKQrLSkq
RIWD8graDLmFyjUVciqZG3IPE/n8VQo54J14qZGRvqzQ/I3m5K3lCEyDrqZL9EfK
007v3LjbweH6FQH9W5uQAQ/uhA2gFEr+336gkScTsm3uJl05GuQWb3/T2CTKMiKH
xLlhRqRBP1sWnYq/AY1xDjnS6+1uceQTJZTTMfm9xebAsQhbfDP01aX4RViRhEj8
HSeohfHvR54SDjkJLhLwjpWSn/aoTFVg9ZhzBnvjXMNOc+lIsAgbYmADtwCgkSlb
wigUydm7P0r5uRu/QsTSAR+qkJEdi/hl3oBv+SE/XGjxIthCkcLwVpHG93K1BELy
03Z4JbFNofy4RBt73ghkVSNg23hEGJsVQc1X7vtTcWS83ffCo7n+U5JR5i3Jf+XG
IXKeRnNwEFPb+WmUy77pNE6cCfz65s/zbEd8d0PmNSWEkAxs2nBCzYYh4JgK95NB
6QtR0SnUwh5vw/2ywyNRvfP8fG0UKDqH1Z7foU96nsbSaH+AOTLgZLFxuEeBOWHT
zxKRxUaj9og+MugbR9S82qArN3mW2V9etR3qvRMjngHg4rVCMqGLCtxDTcLaM7mO
2lA4vV0q+veTEAK3rQUPkUK241gDxWV6ZEmSn7Z9OAlriRKKsrxxUidQD8+J2HxF
bmD9gSSXuLDSgRAL9CzBe55wEKac0BRg6BWNHpYHvADxa7K4VpeytsGnvPW5PkHz
XiPiTqrFJ+Naa5PHcwnTaLDYh5BszSSutbsmq2L7MDwakoTIskETg/FpW1BNzjpy
9HFZeDn3Qf0cVz2PHloO//IVdCbUTS7uUdI3HS3anMpHBDuKKUvnTH3/e3nwqunA
EZtwPO6MlDIy8SzRkVk/N6rxzk5a+W69/PpNs99DeacR/Gv9+8LNmZeywMKBIf2U
q9Z8kwBH1CDiFAP6fC9h9AzVrnlj0mXrMBE1qaUgOsBrUhS6iny4tp0akUDE4KqJ
Q038Oa16FkjcZ+KIwzIA/m9BZJDRT9wXokVwBLNHqkOiaRvg0HLJVpsaocg7+WO1
n/2Oej9O9LadXnXpUR+qGGPAVun81FkCr7WGT09Ey1NkGjUyZYg4zFsi4ExloX8O
+W0bmNYAw8YZVScJePHBdBoIWcasmzv/64LSunPU1P4vW/k2lH6avgfU1LkXldje
rsx6AJhQ02QUbWaZVH583bat9WfWPb5Ibv41Nfc+Q1iT/GHWZ9KITjLBXNkko9gV
Pa8Yxkbo1LfbUikLu+7v9vC5mVcnAv3seRatB3nAq8WZIASVbQlBqIYnQK68/4g3
moK24uFspZwDuMjgdq294nigUwPmQdGFTyETef6WNbv3SJC/1vO5/+FA093WvcFZ
BWcnhzk9OwzCk/v1ZJmd5L222PEyX77wUTBLVh2PVhqN6YA4wYbry4L35g1cPFFC
7VaabagScUY3kGwDeukp+n18IxtOlHyTQ/0mVdYrL5kK9GDV3dnZ//8YZJNO+CNY
JPnT9ivwnASuNaKdTff6TRaoTWnw7T6/ETzq3V1X9yhR8C/nDsyph2d7jfKULQf1
I6wH7KWxxgZegqfulCALF7uTsZHz2TGHrL2LCRhVCD7kL8hYRtRTp0tm0UnrsDZj
3F3g3HtKp/i4nB5CHklnn7hxXoDsXyFo+WIcZRI+Nrgn6ngmAD8hYAyYSpnvJ6PJ
MmSaz+Hz3VW6zK3niiJmGIq8Ipl5KT081qUe3hWwXIKfK2OVjM+9/uWpXxFjEyjX
Il62jFQ4gIaXvRoX3p9rkNCAB9hcmjjgtZhm2/F8GdvQD7dxBZFg6NIs8uVPxj90
HAva4AFGfIE8QeTjkycZLBlFzgqR20MefAyCrOK08uUlNLlPXpse71h5Jqwz5AOh
7sK0tk8yUK9K28SjnAzs0nBlUyrspilczSSbiZu4Vhw+nCcZEP/G6n0FFarSqajC
l9A4cjeXv76aRFmxrZ6yStl5X4WEGFQLcZ4UJZKegGAJt1irqqkbQnWKeUWJBozA
Clzbe//UcVfQpdg2CzRJ0LmIWKakwPddZsbO8bAu1f4tzf4cfwm8HEMOgdpTZAxU
0VyXeketfX3W3AQMFKrX7FpyX3pwVoFpn/UKdyiVHIkSIgUn5oNTMvf1OyUNtSix
k2PsMi/BYl7BK1+4PVGA0q++L52s/O7q1DZWUCulC6bvxKmCuludbL7jOHKYQm78
QUq8rN33Asu2Pc3WqXcc5xAgXiaCAfuMUZ9xouR7Kqw7ejvveNfwUm6dgH1pIN/9
wztwVZAp5q26BBRJBrDKyb480lYr8oU3DRZ0ziLNw4Ru9NusUPmaun3HYeaKob/b
ZtRYlrxE6ldkwMTGRNxEjrDs8/4yIg0a7P1qAR+/zkGUNyMDq2RJYnWHvfK32i67
24CPJ3LTr61riMLAAOdLqjMRlm7ZkGbh/e0qYgv1HvDjhvvBHu1pqlow6mNEI1Uk
sTYia9vvXjBMcpM5v5ADmaHYGLDWbUq0HPPM93JSFOPUWzRR5ZCjuukxywdHcoAF
037c+PoUYxhJKcf6etw3OVo1clggS7ilRSv7Rq0pd7S1jVrUC7rRQU6Bxw+M5FOa
vc9mAJhIPxmIjOPKmFphjELlMmWDfVfhT0fE5E/HmYMP/26zS00kgEsk76hpq35m
DO9Z9IktrTYx1Jhy6lAq2YLf+hyIRUOQaU+qmiCbs9T6yXVkBM9cvc3FNP27rOXs
NQmWX4vSttxNArsjJM7tjRcjv95xQt7eblj+s4YDNqQJwrUfouZCqzK+VCj5DIco
/NjE49FtomKaa4Q3J02jNkEwLBGQG2MaQh72vhdab/ALyE7eTnUKWbykeEkdf3Kg
XnPZqXcm+EktHPuBGp4Xma6QsnufFEQO4AwhJjNg4HbbAby+5RUHlvkyZDCqpiap
BSF13hHnjGFP+aeYojbhMI35Wn7M0lFYX3AEf2IcWEX4IysYKRq8d5MjmQhZhoMP
wPOUEWiSX+LWy9PY02+eC1FUSduKRt2Be3IjaGEoQ95E5q732Xhtcb9BV4cRUvdJ
J6F+wXIG69Oz5Rm0TroIldBuh8TsF18CN2pG12r9S2pD4wipl006XzBG2nhF7cot
DA9N6orp5PqCRk0JiUnRb9lWcpHwQX+gCfcGSUphxBFh80H3GvM39SpSjMm00SIN
s/6BLkV5R3FPxgrEBCwqPad3GL+2gPI+ZJe7y+K0YQs0UDxYmfVR9R1Wm9Ywokm4
94l0sCj8FD1Dt8rBwSzhuHLnd4aeequ/1Uu3eUbDRHxoyiLwRi/yC8LqGZUPsCQF
bDrjIjWguFI6ZDjEHfTrhc91HA2beeBLynygM/rXjqRs/sUMCR/MnyJi07FDg88u
hG5uySlsCqazVUbBPmhKf5dNrig2Uh2u0Zr3lTVYqIa/zQxIDIGNf4oBMCYNs9IP
ohW11GVd+G6iRDcbgxHKABamxAhR2uSdaY2p12rk9sGWrBiUyfCuFZ7aGom9/DwZ
s9zRGSs5g5nRUVv1DIp9h1KSmSymJnB3/mybIw0mPNl7eV8oo5W9ezo37BOld99X
5zFQaVCyXAzVqAt6cNuhRMWVxYvJWafc/L31//c9W3c/Q46IyrfVlDe0CRcQrBuq
sUlq/K5Pfiq/PmLY/CujqTZcb2OHSGd+I0HRWaUf+mjek72exXrJ0bKrCf1uG96/
pORsAE8I0BZ1sw/n4W+WTrZfIqsjpZhV5CIN28Vlkq2XmsvZnDIcaVPPEsy0yRwe
vIPvznoR3OfTWs67r8SM1Weo1OmbPGnNU1KNdte6WriA0rS7AX39o+04HOEcerx9
vx3xSPKzG7+y0iatwPWN3bf1idClO0tS9LVA99CkQbfRCfbj2EW6G51Tu4Dr2TzF
nUYeZ1MGfYX87xgbIPsTIIU848xO7dC8XSPnjESZCsFgfS715Blu0lRrJqIXcG1v
PsYUjeedPnbB2dyvVd2ZPpwjjX3+lcM1yPXZ70O0pW9HYGKmhUU4Bff0JdHB2i7P
A4b72OW/oXyPQpB+dgJZvmSXssCr3ry+v5ZuJ6H0wAYM0Jyog1O32XgQ6G7SSML8
Uq3Ru1nRoACBpGDcv3HiXltfLR2IWoVjjPpnvIZ7M0ZzP4Pnij2G7sppsx2Aagwj
OmhaDaW1a0WXVBHp7tOhTLQPXIb441+1L2rmpP0a671zKXw1A24YS6KJ1ICBdq71
B7AJPDCe5RMizQWLkoYNMQF0Ob2JBxwuC6+oLL7g3fKKlD3vaBuNTY/Ath88IpEj
8vThWiAvHo1f3S8yoDzaWZjS6ZAE08xgWIt14sS6kL+KpmsZcXDH+F6WUwATUnSf
v5jBcGIn7T0h7UeFpWp2QVvGpotiR/DerNHlVPTrb/jpWMqMMcgwJ+zvYw1/Ytft
PzqHS9XYDPy9ZDb7eOagUaKpe/HTiWMrtMwyanynelfgz+oGctoKGWr7SjgVH6jF
fFZ6zO4PvIp7YDPW3iEIGEYCp3YKnyajdjTRFdM8zFfA3ZcEVrcfGTRxs03EG5aw
Uv0ARPneWHNGT9tunbdEk/GxgETr9w0AJWNshCarubkpLJ0KDZMm5SRg0rYWvjID
5NFECY+JbOxvAf9QEZiF/lIIzX6MLf+WgPJTsOdUVx/iEmQKC+CAg4Ed/uVv3FRY
sV0Z5rZwgp8aCNcmD4d74XeBfPRB8MtXr1GUw0zFbC0nS6YtJ8EX+L1b3Qx7K6ZA
Wp8J7gWHfvcvzQ2CUEYlBi4wibD/HJ58M60Rxp1ZAVFzxa9JgPHzdTnkbQCkLRqt
GYuxB4RKA5JyeZOo59wrDmter8WZwY4qspoN2k1wIojsoHqsv02hAG6xI4QXizFz
svKA/kVuxGIbA+1WkM/R2Jn/uZFtY9lZiZw2wEZJuuJSz7GRJzFeTZHeX+dM615X
XNRias7+qB5umATZC2zbLLzjHSxAAoCArtnK++piku+Dysme9co9YSLTdY8AHs2D
QXI75poEpYfPo2CHq/Mxa6S+cFohwrLjUAQrZ3EhjB/2B1+OkSvUC7XooboW4nQF
BNAhEFLF1QoiFKZxaDakCV5LQEj5HwXCQuX+06y0E74bDuTmYmngDX/b06/WUTpg
rhnv6eZzWq+z/WMn4TGyb3SQRW4s3WeCDw56LjYuDKP02PHoBt71mdLJoUZ0+/r+
PKQ05whRNiBAb/XJsSUqcW4je6UMMuWXXABCz0TEf/x+0PEuEray5JaZ81zR65Mt
6lqazZoohRiQnuSKqqMys5L+Lxu949E/i69w1i8R81NCNU8PokGJ6tZEy3jNjMG3
YycEEVNr0vRg+c9zE6zJg++vzziBRhciv19CCmUQtDQE+1ngyFOI49E+iJ3tbMM0
c+PqaUIlfPdAJonbSIUMf+HaUsKInw9tycT2IQYA5aOl1cKpdZws5kMIdehXHMTI
DwLagwj+CJ3yhqTnqCZVZtavWNYfYFsgK9UxyXFikJ7fg87erbr/4rDUPPJtNSdh
GTediGCZF1oL+Rp8VcaznUfCnGrVABuFfmzu9HmIlkIO+6gwiEUcUYCFpcNZ2cdF
bsjRnF5hJZdYRoBKSeB9JSCVil3kux3BfLAO1Mj/CPX5VszAqFF8BgBWRGUDGaYG
4f5tLHyKtH/PyMDuQn3a3S3XupdFELf9mOB1nLGjKyW/M//e0S8C9VIaI0GAJkGP
bcuuqHdWD9IrnYIHAclI5DOdlhQh/MCwYaX8Rx4dRh0u2oqHXfMq/HEIRSa/xmH3
B5BqD3RAgfrIYqYQBvAg1dzkPpUEx2eQbjvzCl2yll3UD5SMCgg3zKH7U0eH+ow/
YQjQaW42P6IBRfRF5/d5AnudLBbWDg4TLiFJxoz+oBEILfphw/sN/JOcmxNStiin
ERDrh0Z9wKqFUsOpYrHe1dbkXrbHZ5HNpxv4U1nKBpUVKAnmbLgwJJRe7QQThP6H
dnK8s90dRfzsW94RJ8xyIs6JF6pusykm+Kvkp4OdW3q6g47BANqDsCUsEWSllE+A
ixJQMxWu+0fPCK43otSJnjGDcbN9NSgzdZNiCPLK29HBvfOlhKvkDu96g3Fcwovl
sb007mj7KQ4qkFUIKrG/EOcHrkO9kNKQVEm/FjwCCMhMwCxgJKgljDZrZ3aWboSE
r4gFgyHiqL7CKIxqTsjTTYc7OuVgEPjoN85jlUuhftVNN4ktV9FuG3A8aiIZXStd
JR8tkGfM/0kzBE17H0h2zalLESfoCq+C9mfTbiY2DThCazM/KK03mKU0oePqmOy+
VcmBhc0zkKPy0kMCooO4mpCvuDWTqGyHyJ0F2gjkjB29QNLVf2zB1AsH8Rzu1yIf
6da0TVg9WWNNowo1EA73Mx3eV/KqtCTyeHCnlrDEkv5O9m2S0C0aqYabu0PrK6dC
G4ovK0pDO2I6h8ztmPHwaigJnqJDa90OowdYl5xcR37SeqCjP/AkxNkol5fNg0yP
i290LzvI2dTYQF58mRarEFnjIdWl/24QN2N5w/virTAghfzd5/ryN1PRXa/EDIKt
vfTKZGCk4vJy4qsWJWgWroQFr57i/wIxVQGV8fYXOt1CXfY4EH+o1COqN+dV2FBj
cAiwPug/8vQYOxaqcfT8OWcrMnuE9n4k3lx2+FZxyn1G9cyeWs/sUJM2s/MmqQSz
6GofDcYm05syXrH1vStDz81a57yKLZRVBtht7sKqWj+jpkofkCjM+JXDHkb+EA5y
jBNatqGgks732NbqomyfgYeW/u1BDXNpPkNV936Vk7XRMBp0iMqDPHB3gTupICdy
M6JFqKF1CZ7QPzyGse3SJAWBXicizBekcSkGtyKJgXVRxIPHUfCDlVaimZYcPFLg
IePHEzBxwr1ozZ74yedocG/O3zT3MwXAusgO36RjWV3UbhZ6lC+xnZf0pWpFyhJu
PPrykJSQWmgmmgpUYrR/DMjwTAhY9i91wANLVBkuLSbDeBp4pByAutOiepK8e0Yt
NQIP6mNsBs0I5ozTJ1+mS/RtmFGBAxBJqpilH3Vtj34+tzdACSfIftvcn32MujCz
8BHrEEYRTb/SpInHNEJtDdV+ici3+4om3izy4dySdkQsw+z7lPJoAGP2BeW+a1ou
a3mI76XGsPjImHVHFCKg+XSuSv4tMQl2ghqsbNKqIaEVP5BRwcTnRXkgeaAkuwBm
LNL9hkf9RLqWJ46zO7eMyegsma6MO1vmIKSzvt4fNBFPbcnwTm5w4W5iV+/JTbNv
rHtxUSRbUcKltGdi9VcenCY9BHq+ByT26g0bVtVrt53NdNqzhPqP+XVV+2ddv3Hx
XXVFLmzJNsjKSHzVfrH+1OHf1kyOYcdadbYSSNN0kXqEBJUwzU67soFgGibeh6Vk
4Hc4WWxR5k/+3HNZXXb2CrXeyQWmsu07JOm8yUexujT70XFyPe/Mau9aa/J/fwUm
sPKigh1lEuvLbA9Ku2LlyQoNHA5U3xUnDL75RZHilN1dLbtoe6jZLm8Fzl4rGVTw
9PSThQdf/FIHojC80QPSVmMCuVdj1RCOlzuw/HzW57BVoH2u5QAqUHlMscv9KwzV
lzGVnC4zik3yB5gWEprIxmPZZiYV1xhwrZuKoQdXH0qgkFnCGUNg9p8i8EdSJdy1
xAJEN9+juLbj4JXNs2D+nGdbSBMIZdTm+uvwBAGLppGNntvSPdsadQ1AwWxI5Thz
6e95t/bVO9zUEJzsJggooC7wjIpL8AY4nDCV5GTY5OCrs3RN8u9gd4Ajox+lN6SN
HqmjLETWZt3F9UGFBGtFTxA3h1dhxAxSj3/Tvsi1pdOPo+o7ZWb5jHOddFJBqkJ6
S964fVug0Z1J3DiwRmAU0AhSRMzLRiKIWWsKquQGC7l7lm2/7jGMkgm7MqwrVOol
oFdiNavjaymkEdWyI/pnyHET7YruQNQzQZLplSDl8AL3xbGEOCCcS2yDX5HVr5Gj
jo2/tji9QrAkmdTxHaBTKXdKgAFJCz1GhU8IVRz2Tyq3gnkVxGlEyS6LuiGtQInc
Wm3+pnD6xFTu3Sec0C1IjYcPz0QH/kilZ90PFhVOli0XmHcYEFMhc1u1TZcYrdva
AWR7+5OyUSSfoF5zhaiNf8FPQvOvjlcdQcE6jsap0ML9y667ixkP/P7NE3hSKlDF
rOlBckeBg6SWdIp1T7sasMv8gES2UDS+S2qOuNddszUdIWz6eWa5EfddgP66+YRr
k+Zkh3Yu4lY4g544rtMKwtPpgu/2TQRad1iMhKCjuaSH2hdRT1uNu81nE2lKBArY
YxKtbKmHRt7TRgZKkcbrK1uTx1csI0hEnlhMpjSqcmqsQTCjCNnmDy+ZByVvItLe
OETWTm6XybBZqZJQM3Ahw3YjbEZXS57JM7B/6ulU41jxtEtrEiVaPas06yJy3q61
76msR2eIUcYg+wbxWZ0z8ynMb2vGvGVogvmO30HOWNyfRBCVleZHzp5kiFn19i5Z
TORDxKdJehe6v2uqVrMcXZaLhVJyyuwUvovuswbp6rpfKMOPzbfBwmV6g9vYd25F
dKZ69w+Nhncjbic0gHXMtc1RYGlfw0i8LXLcAxR7HZb1WBGbhOuPLkuN1ddW1nDH
Fqn2buRb6bTekIoRI8jkUuI0huPyB/lAQi8nV1ALfWvftjPqdV4/nKLcg3+qOivM
UsRh/WmrFz2lM8mK16urtpoxXbu8T376K4h2GDGwlEm1BHwK//QTtKrgKzMnS1FL
skhdXd7zW1+st7TDKoKxE6CX0MatgZ2OfHhRzsy90w+uWiuPv/BlV98N2+koOmZ9
NeTc1t/sZPaNDGzXkyBZaZyYgqhlAXl/AlLoU706HUVTx7vkRBXOpcZ+Gg6BQbU5
CcXeQ6065IXVH4q10fg3F91nshrHT9iu5HXYWu5ui2W79V1LwZ5gti3dC9mWnPyA
90pblDl1mAfCnypEck4SXe6oEqBnxFTreBm8jQJtqnJ63PosC1brZw7eOztzFnrd
A8TPSQHh1zxctrC3KXPVIRA5Y214vE0fKdxrWNBNoONLlxHJwImkQAK4fazbxkkP
FPfakTTIjVdMJ57leNaAgLxiMUirlpXTH8W7mwlY6HVsxZDGcdyfKz+Oio85YtQx
/8N47QRcolJWvtPfNNM65wSY7DvY+6K+i4ltpIPA7CaJqAGZxSvSEoTdQrIV5KO+
HwcucDU5deDDjh0zVjaKbH49iCgLo9dy8YnbMKvnFpWMXrbidoDExBotptZu11UH
97hBzUzdK4vs6Uucf9BULvGQtrfELXri09v3nZTX+NiPnxWiqe1dV/3tKvqYTHPq
ALRGSgj/OKUWc8aRaOQXzi5rsnoAw1KgxJWraAZ2//6mRg5x5CulhXmLC46trsPy
pyYVToPxG1AY8DChvLnxT6WBaeEdW26hXtEbTDtaNsVVZa7G9oCXXF5RlXVf2kFa
qroT1oYZr4hWFTJm0BmYLlYO8bHOphzF2cF52xZdxEHsiYDouLM1GvrRXTJby40W
FL4xmDMpF9H39c7aYt8uaQS2aV38/SX5LpXau2hdgiUmSk3bYDVG5X0RhuR+/CCb
pp+9JWdEV8/jXWBc3/oY9pGUKFeCUVAn9z05OGol1p1xksqwmNyDJqDMwb0k39GZ
lVT9T27IkqLVgi+Bm+7nMGQMx9VrqmzxvnLJ8vii468KtRVNuriFz9mzBi3sJxa9
ofN08wFINtu8u3G5+Y2FSS+3OpLlAhUADsjbOgmNX/soa9ZlLROZKCOuH8PJVLmY
ZDnLLoxPH7JhY3SH6ixu6QlrxFZ+RvyiJxGf3PuFME/o/5VAk94Nu+pj8pI8VLrF
K65U6FVOor07IrZ0JHAVhSEH+3Kboz+YTjGfHt0DH5mDtROnTNIKKcxmsfAih901
NE6Vw0VQ4ws9LX9gsPTFCZRCxoF1Z6eolzqf0AmjrhGJP9eq/sVsCxii18/vTk0z
5u70KomSwCRPiXld81rcr44PyljVUGHiScMzor2sEb+SUCmmVzESHiqVkR3Bfrio
iuu5a1NVeuUj3M71PFvnjYhjNvYRvF1v0zZIl+HyB5wZrbQqpRCJMh349mGE5EjO
q9+xStBugn8TLDWnqCT2d7dF+alBKVXYqScKGoipRKYUI5pv1BzzecXxZo/+v9xM
bXziw38z9tzm2UZtYRq6zluFu36ZpZtx/ZV4X1wYSd/NryWdmZdD2lbs7rdUjcN4
tNRsw2M28J9+Q+P/zVC48S6+LYm2nV7xD/jLCc37GcJ0jVWb9apHBP2GyHNb2lw4
FAzVZRNpLeE8RAafHaWiGBQm+1XIPb5dO8Zhk1XzoHXZre/7EYjvSZ+U1hGJuGO9
7YcD53Sos7HN20xOZ9kkP8r+gTjZb9F0BbyDgk+FVGIRQFRio7kXOd112lAqODo/
RK1Xg862BxxeXIAVhOD7ReJbnJk1Q5pgxsCuM0U7mHN2iCZNBKP5WA1QdT3k9fyw
jtsb96WtBYKx+ew4JGwhVrYww2Gr9STLq7WbhoB7gUCtxZQm24mR2FXGTJ7QzqvY
+8SQJsRPMfWwqp3+3QQSrYYUDUNKQs+BiE0P9SsJkLLfuVrEgC4Mkj0kLUbXg+4V
iRMdhlwU0yO/w8luXTQr2jk9mR50BfKNyIENR2NeKEH+hV9LfyLWrFAF7FA2Asp+
caNBU1PBJhxhUt8+5uzyqMNjlh9o6S0217HEJU6m0v8iI8e39EvoFWt1vR1xe3BX
LE+I5xQIK61Hav/5DdJZVxm30bCeb5oE8ZPBcX/DJro2Nu29nvhZGQ8X2rkBTDSi
WQReR7LMGsbpYmNhnkJXWXIt8r6iuzdI0pEqylVm4K7hzCYUhq8EWbc3/i9b7Nac
Fj83TjNjh1ovJFGc4q+bP+XX7PJmooPTIYRMm1qBfgk8R66sNHQZSmmApmo4qE1p
Uf9hsWrH+LIken7SBqFsSed36BII462XqpAUp/XaMkoVwaJPvFjjKGFISZZDE+1R
xtDNqAI0hnQcNQt33sVCPhMwsqYvoaA1b0wUBUyhg6JnUEUIXktJ5voJfxnAcgT6
TfzlB1ajoXpP37IRzwx9IzQXaYx7SiKujtRsXpxumldYcCGm3SOZfL11gbjN/s/l
3SHkZfgHBB5n11tq49cZEYMfStKB6i63b8MumtyoysSm/JDxiA/2rSl7kt3txllm
JlsjmqEJk9HjykQFcj2ibdlV8CyyWwWxYomPNJXZXhavU8YDFghamt3RHfGNR6Lf
ESNT7hIAStj9ibfv31MotcUem5bseEiQA07F4BEwX4N92UALV298aLgnfjb6/s2Q
Sn7z4hWl3P1Vv8zjKHL0jOy6IxI2YNfeCKvn3Clgp24d545549OcCazTJT1ETIko
3o1efg1S1N6bO9eYzNNQ16OWTsacsqUsnEtgojOXrlbdhZDt/GgFv+jzaZHlrizI
4iFr6IsWsWCQEdY1RXT1q5npY7EC7jvu5LmWrQxkfUas95Asy9IDbARwofr3TPAg
G6lvBlZa0lSyql/iBILfNEs02kEQtJcN4zyiuTsPuPto8Vwip86lLsxfHAXzBW6s
K7kKyR5IKsO8xUrmt3lXEy09+e3SJkkLqYaR56ntXE9Hqu4QSxwtpEWYbfRIj1Zd
zUxBGPr9zimumxiisLyGgQC/6owefGmLta2LNFKhZERlaaV1q0LZ5sPahErWsDZX
pqLvnHKPBWc0KAqupLV5nnOKaijlUcBnRfSUgEiTvnHaDnYeC3w/oZ+5prs6YN/W
MncMxlO8sB3qoSGuHwGFCUMOjZuXoMi1bYoxsXIyd6kgk5VWbCCZy+XsOphQ4mA6
TcxrnnIXy4J7Y1Ad1fkHfcorih1lBaN9CQWPuo5yUqzMK6Qboa4B2aupDR7K0384
7yjCMguw/aW2Rd1SXpoMzFoQEhLyLiXqq7QKvahxTso2ItUFYK3d93+g35EileQM
TtiiRyl8adDl9hb5fmYSAcUF+HX6+7VweI3k2JIGB2n6UlzIvSWZ4s0KkxszBTPn
LU9HO3EkYak3tn3JFbjjy4kJ/T6U+bPho2FoaAMC2XEjIn60Q0cSyUf1AWrb/7UA
xDm8GK6NZRLotWCCTnoUCmCayWYhsrsWuUMpaoiqDukVGbZkgOJSx9Qhgy25BHeu
dm/jGvlcOcdiuQ35PJpA/mgbGo/L2vCWesPHZe2t9EsibJeMeqVD71PCBdcAXnC6
q76QYtKYofVdrrlk03V1YjBHZIZzl418/xSd/gUK/GTu39nILMan8oV0q+4r1HoY
HXts4eRlkdPj5e9+dYjmlU1MTtyWYdIihYodBTEXWiROLpCXkDM5s4YH3ET5PSIp
zPVlaM4IDfDek3F6bPsi0K1JyqxdzR+0SdsU22EE6KBNDp73tBIidPPW0t/pO2/D
ANJfMWBuxV1J1vMfnt+fBmUhkSjBvfT4WVbk4MHKyDB6bJjDIF3D/sMXaMSwyEDE
b6GC6coVP/5YQCBQQuQnpENUj5V7kK9ctBJCZxuesQhV4onVzvLPi6ivU3WOR3uC
JweJ08FKaTViUoqsujgzpYmGOzKrQJk/R/ogOsF/FtfLIQc20nDJWU0jqf6CnVnw
mD3FqAlxqc64G75oyco7Ns8LGCWe4+RjLwlQN4m0MRpMaa6lFhAeW+jgBE0Mj6GQ
jiS/BL/O2lrJTYEX/6f/+4h46MYDlnXvVjyQKiSgWh5fXXBAaP75bVlDm04l8nUL
HRXxZmF4opEp7b1u8pZKAj+iezOMlY/wcVlRpysrFaCxjRpK3d7JIvj0M6Y/kyp2
tEM9MIF6LFQL4cTN08+jsOu0KMoj24OEllrbxpwVD6hcbnIUsrkPUTFxRxhk7U/Z
zoZVCubZN+yfG6WiKiiGzS0rU7iEw90bZrk6AsjwFoXBLViZl7QQvpuW4dwNRkjh
nHtcJaRURVUUHEhLLGRW6Mbavl1zVLNkjQtYx9l4jSpeB7vhKKKmBo1lts9HRpL1
dlgR04OG8lNZ4StK2+9XBcIaOQ8t8ydOlrW0nZAX96f69YlICbw53OMGDwJNCAUL
/709GgGk1mOuB5vr+xCkr5ID58SrgO9B8XoA4yh5cG4k6LJL64bbs2hB+d+bMlaL
BI3pYEZgzj/Nt7+l85m/dghzntZr9XuKlSDQWr7Zv8MLBo/K5C8h74f0k8WL4Yso
8I1rYI+xQq/uqS1jkAm/ekwbWKjJJqaQnEt/MTwpBp3BubqW/XU/Ywk4hZIxnSQb
/TbdNMuspBvweLhbyypVl0ErOKT9xN0699pKX+JSeyzivSz8j/GiSHYqcTrPx21I
fkteoPSfhxjVLMEzWwgtou5fxi+ijB7JNKqzmFN4PZlDGUP78AM/z4jeQwUO6a6c
L4BZ0N9TkCAsgC25yb25k0VS/bbdQiFXfH+IgZSVDcTtu/Pr8IbU4dMcBt6rC3cN
7oW5ZCHwMrEK5F5+B4Z7SezvPxzCa74e5Y3i3yi8IQqagXsaOmnLosUazMtQZOMJ
SmKQEJNdRRuywqfb7DxKQQBq6HMYWXsfgC58g4mdSNF1sx+wCEW8xP5zttlGLZ01
fRWjL+Fvw8tP3ENDsm0rP/UzlmW1RktVtl9g6EjrYQtFpMNh+fj7SAdab5Bw/G7Z
gDKLC3evev7I74o3flm1uHNjXStJHIneTkI4/fCLzjeuCQ5YANC6NxqZ0IsEk8Cl
8ANGLO5cRiNYYbib3J3mrNmeZ7jBExdxwTTbGzl67mUX4dKUgsW8kwK21cAw9qDT
FH6IwTHJwE2RPll0cdeTzxtFoyqfl6a4xIuzDgJfKw32zKuw4h2Tn74Woi1XLcEI
ezsQTGkKzCNM8IncpRxXfgUFKqGafUefiS+lIbx4Tgrj9GhlDMXAUjyx5D4du+DS
vATHLvEk/pH0lT/X7zxYCEiW8rtaT9juveQd3k2OTaoQfduhpByUhgw9b3GQCwWN
vVW8s3ijztpfSehYSr3ZNuZlcErennMtfTE4Lj7i4VZV76+SKH7lM4UxdBV+Kdpf
i28QerLzPBJI8UEnask+hVxwvMf2pzKov8yEBisIbifCCkNbZ/e7fAbZ9PQZ5VMU
eO/7xbaoL4gJFKBkSvp18Dc/7si6C4XtDH+LTRtimwFcgEeALTdl+w9VKgF+l6ZP
UYPdoOfl0XBKHKpJzZmNB0FAQoYLhA2YUPQ/8yCzNbwJQMYp+KQs9I4egJYXJPBE
zxOq0ptMjD19eTpzkVfLeACMzlaQcUKlQnegB6cRMtVgVUPkc0iLJjy6kVJgiKyH
EtoQoLnfMNhKnhIM+5hqh8dUiCyokENzLn9PiJszBcEtBI7akKOxkNiMy1PvkAQ6
hDR3LPNYmiBq/juny5lXnIt9ymDDWGURBS+QiVMEePO8191qFIRtyXyyF/0AP8PJ
yf/xl67J0awqXqwEjnUIHWKHwO9zCZAndTPHSQjYeLd8fp5K+wL6p9DXYY/3QKyE
AfIcVixrsGeFX9bxWks+jc83DHqldeRVzCsGCC3WDPhLlYeLL/5Le655PR1nKqJX
c984i4uuMWPvi7CwdKTsW4LCRBKlG3Q7ltmboza9NG/5qBx+2gFQqJ62wBXDPk2m
Rnjjq67mFAZcMzk0l6N7wDf1+OVthTj4iEPiEzc39SdoTTZFINLwqnkrF9W28fjh
fZorgzFUZxuGovIry1g3QBLBgMRIebh7neBYGIYc40YKk0JB+7SsWocRHesmUG3a
9irQljXBDxy5Vtcsbba0SCCX3lLnM+ckRu9PWt5/r3b5pBoc9oXPpA8DppZ536LC
DcqW8JqU7qt04lVOqSY/fdUZX2wuGpgwpaXMcvd2c47Yqh9+jvf0zrHE5u4Om0ZI
n2wVTpQFVB/tG5gsYMDaRCXs3nPKDe4xrUDtyp8zFdM2KImqif+wtIoaO2kOlhnF
c/U1C9mCFcRcvy3XeMvlTOLKPyqmc0QzW5ePKDZbRX6pNZu5iykmdm85H1gq/HRV
mcraSmKLFIdDYlkkQaYYJ47GkTutNsawilfPGYbf/gRAQ3dyONUQp2TMBZF86HMi
+zpc1hWNJlYRowSQAnXU+7GhpWJZTfUZwfK0Vx3zLWVByywo/bq9hcXECOQXK7oP
VFbK1D30HFMMx9cOtdq/Ub/SZWL4aNAKa+szbA1TXhfkg4xp1+i1s/zebJP8DkgH
KPEnULNxdCfYYT9rA5jFs38dhAcsnv0buRlNB6TdeYxL6biaoMJixSS1HnPw0kwZ
Z94EANA3e0Ih/T23X31nLz6hoLNXJ5QdAKW4YWNt+yzT4Lnx7+eVHW1ZvETfioQ2
6ibhezBZRDQaIgilhs+iKwX9Smr8wrwKqaw6jem25EshXkRAk2k3bk/qMeXUELMb
9oBOdza72Czzk/z0R91luAqDNxdJV47vnnrWoKZDhUmbV3ulvzsKbNJ8/itF9aeO
8agKAT0UQiqAwjy3L3qhgSbeigg5GtF4dQbRGqzaCPRR8uLbPor1rqVeEDUg31ux
hWKNiQrpSTNwC26FsA+5+JIvQonMWMUsJJ8XVbSp5E+PoRlo09Bfa7G7MKvjYSrx
xgx1dzIJ+gPyFPFsrvztumhPs8nabBpFqCcskmxPzbH2IHzNwYkw5JbqbwVdPU/T
3YDfx+pN2fSWQYPnmr3aXod3LzqSHYKr2WU3dpocvsKAZGzLOUZOLTrGYrIQERik
mczX34k1JMamDiDnNCUyzrlg3mUjyEAIXC+GGFar+1lnVk/CQZ/TyaRQKMZe4hnO
AJ8y2Jjhz9kz/oD7+ab2ls1KYFpP4ln1379CU6d2b3cCiZm289t7NoXwAbKydTJu
/+NoalHbDtHSHDOFz1iDPhIouTeSc4inUPaGZxAM964nB7eFWh1YBG/DEOTdeFwP
IdaLO8XP+qmYpV5OJbMUwMG3OeYOy/FzpXSTT3LsFJjXjZ/Fp12dgq656V9ichdW
eg6+q9g0uCbEs84aCdH5TQeF0iFytjHWwpFVwCStIs9htmZB9MglLiVqDyGTt7N9
w2adsH5MzaLWpBmgY0baqpPcHyGeARlBowy7jGAJhUwqHxi9N2FagangsRc1O/oI
lNr1UoY8pKEw21m38MYXiRpO5PgdQvKbkYXgtU6irvKONK+i3N3rRxlfv9Wnofvb
HDgjcoXWY6RG1Y/Q9oAU01tm6M9tHBh/RKVMiUe2CU3LmkwNEkh0zd8X5pTXwIiE
JYRczNjDKmUF5fgjgO9X19u6vhxTipoavbyjp4tKI8zA/y7ngq8bGcqsk0wuIDkQ
Pa1FikOSH2IhP2aDnPJW6XCmi1GzFoILC3UT1+CMLZvXqqn/1Imxw0OPbYv5TS/3
ArAKM4omQqlfwqgwLGiWZcdrdCQFcCoPMWGuTZ7wXnkxJcuk5b1lDrR1BrthmSEh
us2Z6xOq7zXYA0wYsNAAOdogVYEAvOAFiwHmWsAPf/GXY4hhEh+1rTsFbFtv/JdU
7cmxslpx2nlUmgASQFZyVLmVL47ggHWYk6G4r7auoZoWda5FE2EmN+JdRr6Hait+
mxw18wz6Hae0d63K01S2COsFKEA6cuWUjIlUCZ1AVCNhEgg8U77MwKm4uEfb5iXv
edHgIB+d1lpaoZFs8Bs58JsCAukOQ+M+9Qdi4sC/kSwrmaLEgwf6PoylGAAkzzrQ
ibma0k4jQCo9/UCsvrwYcOixRPaex7lcF450Zi+JnlWU34HSHzBdHDSdsBoiwcTB
P5oxoiyOIfTGl7G2D+qG9pC8vT7/jy+eGkSO/U5+n2m9+esQeVp4Y3ZVUDICi6rH
6Y8dEYVyvvZv7LhAzB+2Xj2P0EaE/je2uJZ0Lc6etDZhJq1MBLG7YF93XMxlfs0e
YAcqRP8WvCJUsnxRySKFeRqbUVKPktPYQ0UBGpE52jMRG/fxeKPr6OcvNavs9u/X
Hm55Fk8UbE2QxAn2gPAdWHBdqSyWhcD/Up3Lw6HTPkeUmzk+T09eX+xRmC8gfgpC
kMEnQkOIJVqwRiGEgFyyhpmWmDQEC0XQDyq2dxCbYudNau0Y2RQ/Kfcng0kkKZD/
3H8L0CNyvcq12NbRCNj2KNc/KDnw6qGGBAOF1eUWS+oZjXA5aC2d+mdqf55JkqX3
tE+glyKSrx7M4pb4e6DF9RxROlynqjQBB9WPrFVqlz8awH5TwiU1D6lJqtoullS8
Ko+wxv6kg5cAm8GRe4gxDdFnPfg7eUNFxKKfrdNXzJrMWhxdrngmNaXvIpF3QsnM
yz7sCtAWxGGLA7/Xb69PQP4sDEtn9RjYmGGkOCv8QwmRgCxV1N3rLHiDPr5zWqsj
ZdrhSvuT04v3Oh/+rf9fK9ElvlGQskGa/nBys/1H8j0OwG86bnO8qTPitsYYCMxy
xpmF/4SHgRgiN6h7XtnkKgK/aAZA67gKFCA6aHkGV4eE0ACXqENnU4OhODNFqXNd
o4zNtiAUaPczXSmmK3adE3ySXwu86hFSbpWMZS9Ry95254SJvEbHe/sYacv6Bqm5
+qtofJ6S6SC7IwRUANQLV2CJ/LNjahH/vXzih2hr0kxyH6Y7YkNFpH1gqmvVmYPx
Pxd0i1bQgDuwcC7wYn//84uDMgSnAB9TEZJZPRCuBCsMM2mQ69ijbZwIsExTzhKo
4JKFmfboa5yN4zPBKDON0s3spKIvXBVB6GjEgH3rNYR09m7vpuRwYw1NU7O5l/IC
Gzo2pVDF2isANsb4ik5FK0RRH29aIk/c/V9LHYbgSqsQQ9Cvr7QaKs51XCQKB5Zh
vkHx9TX8/N5ZONmPFSau+klWUu+JH5z1QmkcZsI9gHve8vRAgKPJbnGQLrx/Szz7
LBvYMPMHo7e1MlAYUEgt3OphJ59C/LLtBbIoy2BEcIyz8hf+wgNfqdRwnjMPk/Mh
wyV58Po6AC9DxLNl5LUREYuG386IT8uqLs7PX5CoYZ5MJdK011CJqjp/ZMoNdzic
SsqwTmfkNGL2gQ59KLjezVGCcmui60y4Vqtht6U2DODe6plfUKTwT8eWyvIEo+MA
d7kN4Jw+eQhPVdXNV9hchh0ELCu6JMSRXYZ9qZwFO6Nzul5yU6j+C9l8dBOTIHTF
DPOfwf4lE4lbVMoEfiabuHqV9YOFUdWBjUPLaX6R7HamHTS6VNYkg5RiHnW6kFsV
08A+piErq7E/ksHn1nnj51GTEJ7X/IGwLhWDMqrY8bAN3f7Gv9q8gBb3b2Htdi8K
iBAmi+BQ+XJ4d1gwHD3DiXNEBxkru1AHAa0QijmurXbMdiVWsO0VHssrP1F1jdeu
Tf8gev+kPjACubS177W2FoIv5FLyo4K+IxI+FaY4QLHFR6Xe3sg0xNrafY1V6VdI
Sy2loS8Fygr/D7gbdEU6gNnhIMStH1mnQ+oF1Avx/KNG8MrEVZbSy1o4Zvu7o+HA
aI01GGtigT1nSnVY1CFBckzt+Addmxzo0YafiKwGnvMoX2+0NZDbzsyWIhDYTA1v
luKZz1+XOvkjWOyrVW1i1WKQkzrSsrlSMZjfeZuM+2ARQGRwwyfaXihbLVWlqOfU
zT0jttkkozbsrQU+RwQTecMMqG3mIHCoiqJcV+E6Z1kSOeKuwTQnjFD4eQyT88Ff
QXPaBaOZmHHH5JLtJsEdsekGR8WBxe8lkupD2YKFjRgIwUCURQM5NT5HLRAW9Qq2
ZTLl0l6C8X2dgi9sX9auWqX9IJD2Fhck6QWludaxnmux/pY3C1hEat4OEhoGn9Hd
NdBKEFeS85BYM47Kmei0Lpk7R0sOkXaUTsEdVdQ89WmnOqXWhftD75Iad5RBQnjh
+nCNATvrf2ZI24+IksAWjmvyjq3KKnmrfyFZoWpmeuMbEKs1Pbx4hrZjPzMj0pSv
irNniexJKNF2qKWi8LDJHhKjh/ibHnS4M0FNCu1pb1UTJnsyENe4/qGjJQP0+RmF
A0dZoG865h7eNXwKHEmBjU8abfivYyB2MxBtff6F3wHZWuTm1iGausExYL/exh/v
rjcU6Qk1xhZ8G09AvVQSGHtY5j5FZ6vUy89J2GD4vb8Cx9Vfe0M4m16vwoRhZnMi
P+Jx59TcnIhffVSxEAdW5HQ8Lg1EXibEROgsH8nw+yp9YAa8pm034aELqGNHq6MJ
Dft1YzF74GUKa6VPi2C6CWhbPCArsywbyoJuyBwoWpl67qsNhhVv160NWehLeQYg
BEbVnqTKuzPA3ZbZr8GTj8rhgIeT2Zhd7C1WpuqtafP3+X5LDMOPHJ2uZ68jNt4q
q5YjVL4frafSt6jiNRyz2I8fZwMokkmTaq983xWmcCWQjqtia/2z/kTfeJ9Zl2IX
kHToNiU5oxOHEK68xCEPzOcwLpAJf9I8i+o3gAejWwxPQNnpXXu1CoXD8aPG9nq0
dlccV0hFBORE6dTVojjsMQMpDu49llH2VHUqrVxbK8z23w6oLhgNtL+++LmmWskG
bC8KjkbmqUhHiRqPje+wlODh6l8uN32N289ZHO1OMXTM4DSFiiQO66ZGfljoLYMS
Lug8qDgTp1knYf3LQE1QaIps350ehOp8/HNbYRcUlNFj/+GBAB3xa7N3zdbBdoMG
MtkbbH9CY3tBM80IzO7Qu1/otGrk0+L5fBVo2OfcvykGOcs18WHJZTJzrDvXz+5E
CTQqXeJNLv8lCOKqYW6/s8x2W5n8rnOUnAXgyLTpCLORBXK3xfc8IfSenpockkpb
BoujBSBZ6n3B7s4ZWxaD6aTuPZ8JBptT09MDZG4PgeagYxA7vH1LdLrKX34EMD1B
QWVZrgvtXJgHSHZ2xGYQ4XSB1WpRgA2X/T+BJp2ziGXJ9mL5l+xBp9dQ7g8QMwof
keN2Fo9rdb1wXggT7RbCv4AwrkN51unaA6ntBCBmebRCE+CraTRpzAURcPBbnzGh
jxuuaEqcB5rFkrN5NxJUDF3/52UORiDEIG0W0XyU2v3xsX/HkDKHYh8PJYqv0HpF
xJBK0OtA5F1pQHPILsxer/HSmiTQ7tQyN+QwzYLS/TkgDrx+flDOJC+LX86eSUK8
5jd9ZNM/upep4kyNeXMIriCjNjqE88MNIvr6r7yDFSjKtyoEWmY2dzvSptCWrmGK
V652o52bt4CUPONnW6cILfIVmF1PB0r+TCDMJ0qq1EffsER95bwfeCkgHQo72xKa
Q581BXJ8bYrraVVckBTT6rPSiGX+NZvN6Hgul79qMAjLHTMng2wNBH1vCjDqXYUe
+Ept+0q5pYcMRRG9w3VGZQu8utEYjFoN0HH5YFjBR7DUQqAw5eCtKqbRKKYfqoDJ
Hq+N1QWG0ZNfd8UO4xUP/omVk8V+L1e/Pd8PYFV/gwfpse6nWMnJf8VYrJfQGB62
SjvgTduOG2Kv/xFbljBH3UzH2m83W3Fwaq1Lf1GbJiF0jolr9Sjt9Sxibvosb+zY
1giVCtMkpL4ub1Phxv8b75K45oAdzBYNWQIss0DNcDozBD75mipoBUjZg8IwdZPq
G1xkivS/FV2yEkOXxpJyZ3FwntVurKiBtY8JBXTgn2CiCEnv+3vAVnZhn0lM/ivS
EhuYa0oq9QgkLuKc7DQi4YFm6o0JBZT2yYXGl1chfIFnx+BRiLsP1dzpui7c5BXh
tK7tJvuS3Jl5imBOU1oX5nafDCDLCWt84yX8SP1w06vYhU+iudR3ZaL8NPYYnA9z
yHZrDeuIG3YQAuwKZDat2yw6275p5MV2kASzkR34JGNdqRFPZHC6Nt7XvOEpdcuv
wxQD+26M21DNA1PXddeUuhZESCOST73A69fsNTvIcPJERE2nebI4loG+RkI3AC/H
EaEqDkmS9Of7ylA2TRohNp9AoRB1xQOwfVE7fSalujjB8e/iWrrjyyRjUMnpP9Rz
1BMbjHg3vAZVUq1y/zERu0zukYAjZJbtmpDCwSSFg3jXqis6H7LWojI4ebsKZ31u
OwkWj8X3Zp8qcfx72i5rIOd8bplWJ0iFwkIgKuQwa19IIRd1SOwmArndHZavECOO
ay6mV9jXZt9cL97gVBsEscmkkfy9K2QreoZLpFgxnUlMiWY3ajvmS1yGyaFlCqb8
Exfeur2uJJOACuPQu7epHTImYGgRE4AvtfUcRhe9H28AmsjAJ9J3Ktwr9hXW+on8
8ZMgFTdVrk/X1/aTAg59wvK3adaWaUfk7jzZbsUAydMIGbaF2bdPJsegD26whtmK
6q8LQE4yc4ejY/rcB950bUxBmz/W08zDshCpmrR+OdNvsW8J2T1TTDfUWmbYoR2T
UN4y3jvuo74m+5Xy/029OxV88+iC/PDl985eqAxNkmNXUtp3Rf+nPwWcDXZXgBn0
FvUMpCbk+avGlKLF5/AkgkCKYYB9DFq+v1OoEzQAwWIEhjWvw/i29gL9N2CKxgLD
r603+fQUxbb9X3cV9g/kAoXRQUToYmOs7ZUu3cLVkDUuuuMKiqlFA9hLx+WLEdQi
uagrUMRgq2lNE+KWQh6Z2qrnMKEoQVu5qQ9Tn7y18Ec78RkdLWtmNhfy+xGqGsoX
9IG0Ltp99LwKVBv8tqzFTlFub20WiUvRx/oQwL+UjsdCLXwmbvDyegwActk1q4pB
DFoFZtce84bzxoAxqUidPDHwncq1nXBwXTqHEpaVB0oUoSq95SJ3Z1q0mfTATgRY
ZBnKN1Q8WP5Vy4zoBpQjM+pCGaMgkuCOJv/nya5bW0H9LF45EkGygJ545w6fTr/b
1mybXwNIb5aj7lbKdPc41ib+c8CnfFI3No3jyO8VeB3YT1S6CTeKzbUdZ748yXx0
7QW3I+HYhv+iAsFVlVw3P+HcDNDef4WUr3CcqdZXiHBnDMaPcj3nDwgnDVgnPyaA
LtsNoHfpdm9WqYypkOFhgTDIi/s6t7vXnzL4pJvrSrx2775zjFZEzuYx6YeiIldz
e4M5x8K5zo0G75AZuGS6O0w0O0ydunusEw2tpRGu5WEgyC0K8GraAZlKskWbBIhb
dB1fSRx/5lDFY52GnLF8/A4uQFiRwgcEvdZjOFQVBkZ26RCEeXRPd/GDD5I+DIGS
tDedq3rHz2vhll/nlCG2byAzsTvbD0PnOHr61cW2BhXm5JsOTlVEmRfXBqw+gin/
6kM/nTqFqRKOjEZVlOUmPmQ6BumgUjVpf7KqsctAhlJF6C4TOmW9UIva+8uhMm3a
qrAyHdL/ZHzYI6je9QmtLBIa0xe4lXLiv/LIWxkUxH5sTvo/MrF1v2WUXFaXmdFh
I+0MXngrggzta5TmMdrfr0NL0pKZU84vbW0sukS20w65UMG/Gf+vqnO+F3PdG5B/
UCCmurGRCOSbLDQl/Gj+/SuH+KWuHQ1tOB+L0WZvRkOuybq2CuAeiRcSOZVTOnXn
di3/lwogJrdiiBtt6dt6IOHHAYc9EFbRleboEQCmwdvYKl/EW3n/skG4tsN0Pph2
dcXQQByCu/prsmtHumFvAOwEBMq7fLEBSJfc55bCkjnK4a6vtKPwBSNF++qVAah2
zZxNaZ/+JVJowChn6zgNVDc7e8ov7h4x02PP7IZvfk0IUyPYfZofx626TN0E718U
JNoyY5PmYdsJoeEioyYth0uYzsKOCTTLw44DZiaNgZPd0CKvBHFSEFpj5F8RFcq0
/AWid2PkKwjW347lIXyJ1Zfl7z4+0YvT/Dzw5Eetqi9uFoXzvpgP8v4Sn+lmo/n2
/OsUMKGS4YblS1Z504mpWzNoZYjLF59hZps1W3ISdMYd508gMM8B7oI/9nmwB1kZ
rtaHg1RdLsuGkShllIy20d5WNxP/s9DZmvQHv33B9NCwKHhoVf0NnuNhUKCbPZdM
E4k0wiRhEh2KtcM2gAd9cPR4yE+w0KXa+59TzsU7PbvIh4kFCCtHNI1u0KLpC1vc
iOYyLCJE2z81gNuSceruDYG63aFBtpqfAk3f5nk9vSjLUvYVMHbi0MTdft8nkS+r
eJ0WtR4oOiWH6NZLMnA0A3gcYLI8JGKYw7iTX875D3LCZXJR6ThNFbmiU3rTZ/l9
tL1mmoGifU02R7PHzd6yILVNMH5i7SDlDAuMyVW0fJx1AY1I/wP9kqI4heM8F0yG
VJxMIMilwfgaPzkRe5HIo+9YH3CwCKuV7atGGhcx0nngq4RYZW4U3mS3SS9j5dja
Nz+AoG8fysCqsTRm5fBfRv8U/5j10ZvN1yq+aHkcl4f3pX+yO6eQPLUEsoibsEOi
CXWufK02YW9zxS9Gir7XU3I/oCm1553pantbuc29CN8XNlEgdz2uRxNQNyAHjeJD
QYsb+RLOVv4EgulD48pYf5IApDpdIAhwbrOEb+jXwxKxudgrA2xh3CyiJtHwPk4F
kR4EEHxdcpp/1rHulpeUc1QTiPa3vGV+ddYCxVM5uPTL6DSQ2hj5JY+cx7Q2H9SB
y4gZ2ueU3Ny/QrIbPP/LMHlQ4lJnfdmiVpe1iWMOVUkb/1ZI9ovKujwyHFsqDOrQ
6B4kJRjRLSaUSQeLf79ycG3Ikz3vIP/HpV9Epf1KNeDgNF4I5G4vJva2xfZZRjtR
m1y3sR0iM2Rya0Z9hYtAzy6qZQre1pwbK34SzlKkOB/1VRUyo0mfua2Kep6JU2WO
VHBWDv7/yfQankC7fTvTFyVjsROuk61w3ChOUidHArzjJNYSA3HMbkzw9P8U8D6V
xN9oa7Amj6hMyryoZ1WGrKK/7vcfZD0IARM1rXAsulzGKs0meUvQr4XL4UTO7xCE
mfXvN+qJs4U8rBHla3nbt9bKASUU8dBwrcoKrU7a/kdyIzLrcZK8xpNPCuYIWEJM
VPRNPV1jdIQkEZnEolsTLwnHxmNa79GQNuiwQ6PyYGbkgfyb+RQ/ULukLrARABDG
3EhKC7uDOUfG01kup0auhvmrcecxbtYjsRVJa+CbRjifmfsLasUP/4X9YBebvCf4
FpHCa3ts8WS2H7Q3HWYO8/94Y1QQkz87imquY7oZP/IPPWyuv3zyB5Wlif8dYntb
ZKkAaZqdClUHYngKlheUGnHE/cRaiXo8XIb6t33IFxHrd6MsSJyXKpcvbJ7up5fZ
YUbzVit+qQpDKjwffEEdiazN3Tm6AzvSdjHLGvijDgkX748UlPjizzW800TVQF9i
o2+D7ezT1ndSUjZ12LBpyIrqijSVnZIuQgB6Btba/MbbEae45In4GbMKOJqq2vGX
dacdHxoaZkVQE2obA4hHAbnWjcbrV5fzYo6/Lt7h21CDCZyeoyCZT0QXlj+slp7Y
TZ298f3b7FtbhEiEsuFK9RGVjy/l0q/wv0L2fMT/ty6rJj7WulaB6eukTcT3UU3o
41JL2YtgLpzVWq1fn8hYpa5sQ8P3YswzHdyy+jYhQKyra3R7R2f6WRI7YnUfvZBs
ocgQ88ltF0jGbXflu4DJg4QhfIojrJH8+J17PwGVpnNhtU8W9rDGotEoHXBQgie9
gzeW4FU/buxbMpt//wjUFjIeSJYoyDt0KRMZX/U2dXrlx/4VKARsWYhmwVuUTW+h
fHK8fj1oIzRH7px++wKZ2Ld2XXKhwnk13bTQGS6TTiqLorZEo6apNJ54j57s+1gl
eEECajqnk/Io7SyBO612duZsfajEz5JtinCbjV9Pcs7+XR/YEuR/2ftTNlwWc02g
d63jUIkNhWXE48ncIq5wieJA2d/3G5jO+InORiMiTzn9njjvRdVWZ6rxmT8fYaYr
aKX4ebCpRi6J58QFg52J3MStlaLEOn18tBp3DC1TnpCghvbegOxdjLRhwLqQ+GTG
OhgFcjyFg1nZUXYm6imaDXUxtu0dSuzw20Ykh0JkXWBwAXNRhQpvH/y9dBREUcle
+PNIcGsL2DCSZu49BnvqX6eXoHV5SWNoB7SDLTI8/gMMuN3R2q3VCY/HiD3ncpfs
wQhLzn0PYy8ZgZ9V/xC5HR9hjJe/9qOIzMzDFhyh8bLTV9xPwq0bJQInrhvwKlSb
8LYhYa7WldfEgIoU/MNn9ilGsbpZeRDBueQWNlC9jyN+/dnZcJjR7sjd8y6WsH6M
HIfFo3dKnp/zBQl4b1MQswp6JTKDVhDFIFX4ZnHiflDJRAHkJPIDP0WfwINb+tTi
5embl3y6ePSd7ofxpaUd82IoNjhVeIspaaDUK8nGoadxighoVvJlkFKVH/IBOOtm
pauc85WEjNTBnDSr/iK90UiwE/DJ1r/pfpLv+BM45qziAXRqwV5qDKFDf0vhTI2q
DnQ3Z2A4egYgjubpF4cRDk030587PsBLuX778d0/Iypp1OkqhfHUukJjKzWi9Ue2
OeIwY7FMNg3GX7Or4GP3APAdDbWSoab1E/oULK2lLpL/3OUez0ZHk73QugKFXW/W
ccast9kkbzlPbA9f5LiaqPhLbto86EnfQaEBff4qXGiNbV2uNmptni3pmOm8fCA3
xPuEzDJvEdUKBARvkcIvtUguNVW/i2IWBj3Hon/amSzArqOScxHrg5zwCrRrX5Py
3FVJzaKIyavxeGWRQXkuT6Ipq6zbrCaG2F/abL94LrOAHDFvBGX//d4C5rL1kHWT
KFUPeuDWjKPcX+U4QMtcIxgxGg2QOsKVCeUM9ZwWTtp824RD4tv1G9ZBqSpRQixr
CtOuFRCNwnhKmADg4r0VATozk8PcGzMCRV221/Wa5XGr1IkOXgXcdM9Ojdc/wXmb
ETYMTDkzgH3T/wBxnmTnKi7FKwV2tF9yishUIXa3LJBIZklTmcdDYlkorDjfO3Dx
2kW4WWq/1j9E7XUzxZggCSOUTs3tsq39fXHZN1dzldOTToFZbLKhmlnifJFEBVEc
icUeO/DRRtgVQolWjssQ3CvTgJjghGNM7Ts0Wwinw15kZdjCZsRn1eCTNRq26QPo
y77RZRHH6t+1a/YS5rPgPD9KBo52n0yWVvbRDEpi2whQsbXo6/ClRtvpbA1+OPga
TvmyJRQF0/rZxLcPwdgVaHCGMkdjyFlVq7PNKFWpclVreVQs1UlOpwPJxnyteluI
xOVixxppmCZTS9dVYxyZzU+9F1qyWtyTnDaBs/rP9A6KG8ZhW0rLlX86Jw9jr/A4
KW54Pp2qCM6Z5AVGxeZnEZdMjKMP//NPafc5fqYnhuIqnGZL1KX2r3G2jKiWQVBK
Mni7XHn1Ztlp6Qv+eeDtiJjAEKjPoGGrPlH5gwlYBZd28vnuEg7kQskfodn8VmF0
2UYTiBuPfxFOdAr2PKItI0Vd2kbVZUuV092klRkiJYF1Nv6s4bYXVQ3Sd6ozd6Jm
q0mBxF3FIPZ//BPPVikNLUV/EtEBEwoJZ45LkOOh2C0mAkgaZ+x91R56BICAcQeK
lP2P4im4WUrVGr5BvduX7OU9YyXDeiUtoakESeS8XQUHCTJ84MJThCCaMUDAfOQn
5zITaZ2e6BdVSv7K2rleT3cwEpVEu+1jZzBpNBUXc9/6p7FFdE4sfGsUV6NAt2rQ
Sotxs9G4YeM560EUWtoWtY2jwokIdqR5NlL3h12ezbfJA2kWh81D7/M1Di65aRkB
LkFt9yDJyYFf/pSoMVUJGfwOs03MRjRNUjt6T3s+nTslF7EhKJhzh3KcVb8xY3hV
JDYSshgxuhrKJUOas+UTk1C/C4R4FA/+dqd33R9y0xolovFojNPwTYJvg+LZct+Q
N7msShcjhkmHfjpxyHk/dtMcMMbEKNaCxh3dV8jPX1i+pTH45rJIDe200RBWphK8
KJFr0HvWlNhdBMkg/nI8oi5TrrwcdCkSu6StZZUdZjCz3QfuD3N/NY/KFuYkQISX
RO3YTREN2yv9SosPiAsnPsOW63uGY1+6A8RiebKyPmBJrcT+N6Kxv7I6NUSXR7pn
M4N4RA9mFfxJvcIMxp45hFNF12TyfyyC4NqxPMhu5idAMyE2/9QRDQ2xPJpAQ20u
E4zkXHZkLPc2iMUmW0+h4iD12r7R6jy9/mI7YLDQ3bUACyZtJDe/pNKK7ClTb9rw
PzoRV5EpUbCldm5sYK3KpbOWzhfb3jNzuwo1JVpbKhYpQUHo+BHO0ZDsB6a6t+Vp
Z1f/vwOOMx7WMZ+KlmsDscao6v7CSQMJdcHg6PEZkWClcpXCf4K79E5xr9Z/wvMR
CKgDU7JLd3H4ejW8LJs+zLnwAG7kvdPRAIwijUv8d/+Z9PLo4jCv2MLSGfhCS9DN
2OPGeeWKHQ374ETm505cv6pM682L6NsCIMOu+Bwd7YyvCXvIZoeddXbXh06f0Y8T
q9X8CLUyEmtwrQIHLnPmWsbb+5//Yk3iwRvaUEElMBBiu1K2Dds4Yz1FNx802wCs
ZsBnAcbR8IQYYwaRjOdv5iqcMpgiDavE3KnzBje/qb3WTuUv9Xc+/ZTsprzltMB7
/ee2H6hXZIeHNiW5/tlmCudicTqKYQfNYgYIJpEd1OXgdVMkzSOcmEXGH7iO56m9
bu26e0subKWvoqPOpOvyqg6wCub8BelhDlu3jMIqsGoPIKL+FYhrhsqamCONj2uy
6wRRg0/9LOJwe3+P0yfBB4k9JhvgRgFRcLrNkYAPRf34FjRIlFH7cNwDah3gh0lW
3Z0YQUWzNHS9TzO+GB8yYiPPfplhRtSAj8U+f3ky4QbiMz2GCkYtMo7TRoGQNC6l
xJCL/5RPA/Bf4+hgbWFQaNPZWfgInQZbVp2QX05cpfzhoggYxpVC9L8bTlndXwb0
Ee/94pjUThIuE51SthAMiZL1+MNaTKusBFtssrPyPoYwCsKXv8fRxo4Kgt4FVQZn
8Z/YouDnEFgOIErGyw2aXjfIu2VfgsR6xJTcroxTy1FGqwzGsRtGWNzAm+EQcCOy
ipsyu6WsVNg3n9BfRLN+3zdUtLtNRx+sg4/pvXaXfOdHBNT2XiABB0CoPPrtOiik
HkAiM4i8JbM+fP2O+kTuP2t3Rh7lQAde8D6ncv5N3LEb/E+Nd8qQFEWdwj9mACFA
4EQRItWuURq8mOg2iU0OjmhZ/obCAOWgcp/nZ6uMvJzEXJifrNtpsTSjkIv3aS9t
0xLKsF3Udy1OaHCEN5wG5fgjml115VKmCfpjjggwDugpQ3Rn9shN0LKRJbmhP4Rz
C1Cie1FgYGKE2ohML+dqFfSOkny2aOyZ5idPlh4obJHHKW1erDUtL3fxB+hgrCrt
22ZPeqoCeUdzQ1olXgD0T+2F2CcnQLLLptkfGfz2a7Cfk8zMa2a809zeebaeryc6
X4mwoQAhdnuvFp8eYmKzwN4qJAq0ulxWhVoito8oy1QR6E+CUpC+dhYAOwrmfaSW
XrynyLVcab9cuVfcOyY1KgdZVWxdotZtJ9Od77t1F4fXplJp8BCk8DkePgry1/XR
T9H9Grf6SB4MBhMN6kND5ZNDwqIFyxov45ns2yxInZmfQNETK6apCNVMvFXz04jV
z0xZNqEwRpX7Jm7ITWk+xTciHsbg2XkCDQuoHw/n8EMJlEoVThLAyVy6aDQDrfTg
miLwnSHcIbJOcCAniPkVuF4XBh70dywJ2aZaUtan1t5qGv5JucXhHReTCsgH1UiZ
TWEiBpvRIdc2ZF4wBYhf2E/FctmmEQOCa9or1ekS0vStQjVMkevjSFxvnLdCpjDH
bXkpZQLQJ8EFi18b1guBK+XEVSNGORk5BSQqAzW9NglTVYzbSci1rRw8TiPEKPUW
0mqwOeTZ6OgVl4WFUrT1WPfSjPkHnYZSn5onQ9TJIZp9NK6LsSajv9rKsj2530Wa
zKYEhwxX5D5Bft0YuKL3vEJWv0Cmp7xKnJFYvraJB7xCapO9IRNTZ2Js7n3MGp/D
+WM2k2v1OMuvy7FABIoK0jRq6m5O9kZ9E6+VdL2lL32Z4z6/SSAxrzPpINbdU5t3
+vqg9sU+Hc7mKrYokV08pNJRu1V8abtvFiocpZFDZJ4S4RCO/5O72kkXo+6wQU9z
vQSe3XCX8u2V/xL6fLRmbBT5ivYh6UJeVSrzCUyxpm81sUvDT8VvRa0ef2xnYIwN
hRDrUzSC3A+p8sHy55SgifGrdcgFg5OZ0sGPjdiPQ0rzBHH49GIKeBuJFM/2kP/6
SMbgde5eRfJhc1MDCnTS+a2PXAzAeFJ1KqYiMPoElqj7QyG6Ae8XhM88TJZ97+Ik
kF0QUAPbLeoTxSbDBXw2ICBK4JTFq0qmNLXCTiJZLFuwBeEdTfw1ii2tz+oTJtYI
6B5374IpVwo3vSVAS8v5rpD/NBIambKcXjGFip+4iqvl0n2gl/oZ5G0GpRRxpJoX
cTX4QVqHyStwNC03FXmwCmOJI7AChemcwt7k8muBoDkTWgW8BjzVOMhYG4AwI2ii
pZcY6f5lDNAwgFnujkCvi6iUj3WzDgnpIiNYbUM8521Bc6SScTgV6PM2snq7Ej98
f6Y9znCcXvQpX7TCD8Ts6YQp81K940g0F86nDb8+KkQuEscc2dTLEteZyxy5pM+X
/8cccLdFJp22UEgnLlar+klhunHWEamB41edfLbumXkaaUavYE9tocWjk6FU1Go4
WVqRwcxyCqisyb9O7di/Hp3iMUyA+wQQ3jWfwgFfXNKVy9ru8U+aKVgwukV4PkXM
zZI4B+4WW74BoP5hxbwC83Aev1ulbh/1NDpu59GgG9iMNpRR5pvZ/Gv2QovHQ7xN
AvBaAr+ye2R7qi9+Q6f1hX08f6mbiy3VPHAuv+AQn0OE9lgCT3Igx0orPRGdsxSW
X6WSlTIZ3cj6rn+qpw3DfiA1BJB/r5QW0+mhGV00612VB5SFhxV/J1ojriMcmmqJ
r7f2himhjNjepgee23sk9FZ41S4ywTjvH6B+zbhfJ/1iHdyzU15yWOxirJAJEmiO
lKAe0eW5DiFvbMuAFs1KQQ53295xgoG5Nw/EW0S2YPXVcwgYytRi/8HocfHz8EEZ
QBcxM4aG7twq6b6RTdz0CQft0mOBEdimQdp7HJUta0F2fwugYaoklwb7La7s/Ywy
mQ0y7uasHE8LUtbwJv8sVX4yd4i0CcCtYibrQDP0VNQ3GvgWyrjlsSC21S07hHm2
d0fUChysFi5/L5192OqSChCV+SPT0FLVDfbIZYNvSYdYiqZBw3E30K1taZSVZuFv
8JN4yyoUOozd/Arp+MuQIYyRnkA+xIRlo1BEIMgFNkhxg9FlGFj/JL7gCX4zjfKc
hNE0Lfaq+jr/ULCuJ5Te9JR+gUw8eIGkpBHbywt7rJFrQZwQl1hh2rm+7T9jBwXA
LsHmDfBNfYnTRU0CSM8vKJTkT4MWByd4c2/DGEF/LcR1gUefYcD/BoLFo06wnDpN
3Ww8/0GfMlrAhnNQfJ9MkswnCDf0WbUzu+oOrPntYYMMwYZI/TO3c/ENQbLxEWc1
QB8wVwlNMKxby6W8QSrmKvODlpzgE5vtEdBO5wWI+vLjD48TZztupKMBzIfxwk1i
AhAa6MZu3QbeDohl/QpBzyGZ0sTnsavdFGxh1FH5tjC3rvxX91dWRJ8kQBzRAbMV
EGiNk38AkbTqtXkf++213aBxUzou4QbXeNKjxOS4uaZVdY/JbIpZfkSNqLJXao0u
CUk+FlVBn2bEtZ2CMzUCssE78Y118o+rzzjGAwvPVPmoNf2f7XgQWDcSxYoywOBa
grnt1zfBaOzZTKvuqtAKxtsZSGmMHZWB2dtIYDrCUc+NPbZ52WPIcywms62IP68r
C2fnZEJUpWUuWWeIkbKjPpF2ujESFUDOwmPBdZHq+k7kTeuoAS7Nr1bLozHvB+JP
ofvqr4In46KPzLpeHbaqe7KPYuWuxg/sFiJpcyNgBJaWe/OZf9Poet7+WmmOxaix
dWbBTKpU0akxT2ZD/v4P0XIzWB/2r1r54DI6kc9JRRAXPIwT3kCAGWJTjLDrG7aJ
nr0f19qs+7BWKF+DqWFG4xGrLyz3/EQVTTZ37Akrs7Of+hweGwaxXVui6/JAQGfP
xEkHJ81u1vFdtkZa/AwTszpd5hcFte7kc/gAF+Ma6YOR3pIqgOSyu8HapmsmVKcA
TqfjU+N1T8fdAgCx0Q2k5nAwWlJpiCvevy2NF+lUQMEQz6+M6ZiBRon8uJJkNpil
y/Mp5C28vtVsyh1JYOXI4KmFlZu5KOEi9CcsTEPR82z0iP5ls3GStNCQB6wbl2FO
kIwR0CoVYfpcykfds7SKYnd3EJAQFyBoVLYvb0+hMDE8J8bpQ3cU6fxrsw9S50Cx
0DQDehT1GJIbwnGKgWQQ2WQllGm4q91DBqjQwPhtyB/erhu00PHB/1+oUxABgp72
RxkZShXmfMVVupt+zB6vkdNyIA/Bi/znKSF16AXNVEMjJZsH/lsnnnpVTxKp8W9y
iibUl87ffQPs/xiW5/IQwe36SO2CGTTtKYKgfGkc8pTo709oBhl7NHjDRwVTh4CF
1kQkVh+h4lYyqpCuznqDggEWsD4wfS33vBtNHVUIAE0iJxMNbCaNWXxoOiOpVffE
IYe1Q/H/yGYVKKkYJM5YJTnzuDn52kpP1ciQJH5j2IWnfxP12TyhvLUg1clW2u7q
HROmLBDKIXvXbxO+YwL3pvq5W4fDQh9DZmmWFi5SzGvcqIfZLUORloKMvnebEJXM
CuQZ+yQN11VpmN5bgURKSSvIoJOA/idcTgxq0CQw1to8Ve/2A09KEA7+0NgAp9++
wnYp6sAODe0hh1yqoYaXyTFvb7ZII3CBUb/ZOCMyQkm7MIvZLnbQxMg7Vzmxsf0d
P8YQfzxDMehhdh/6sIeK1a90ivSCjxmcIHM9WaDg0iT6HziEyOdF/XK5WGXpdxIO
fwMeltxtyti3w8xX1V4EpsA+a319TKzU6d9f0k/8tyPH2DHTMMbyxggx9aVmdQzy
roggHvZVoE4LRbFWZkcluycTEHD8u+amyOQngHK+wCAdRagedoRcp71LHzqhBWnj
+1ejmlH8I/jOXlK3KbLZvjW315ybnsp+5OtIdYW8wBtEp/DA1lTquDDzAyXxfWrl
ruPVsg7dBOiTHA4Q507YNz2Q8UTIN+5WzTx0SDlrqiIJOHQcsStAPiKtK3hHSouW
+UnBprtf7+ibpE4fDRLcjJkL7dE6yDOJmwdKhek7HwRtVsx03oTlAPZ+F9iH8Vur
Z84oZz5euSk8m891hFo3MSDvRP2xugCywJgYfj2/LQUbDYVBdqtMVvfRXsh+S2Pj
P8vCffIk3wtqHfSh7NTBfniqSel52wXD/C3gdYuvMASbTre5DQvVFev0J3KDh+Bj
QPUbogg+nYw20HAi/IKpNwap/L5vm5Nn2BsoFTa7N/UOSQfwlbg8Un46fiUBgF6q
sZ6bXHo6R3txj3imri7JI/grnFu6ty2PTzgNlsE6jOECAdGohkBTkVAtrZ6w9qq9
JH4AzLYOeU8c/I7AZHHBGCknpD5fviey+fkakUPeNxS63haRHMJmjXxMHWg1HHRD
S1q6uegGjILYB8cG9VVY4s6MCjyI2AYnOUyQoJjInm/Jj/pLaFapCZksDnN2H8u6
cnJ+zmVCBKef2NGeMgwZ4wH5LPPcxqo3xIVxsnbwK6p1SJirB14KsinGZ8rofV4t
YTim9d1Lezb8llv4WbET6HuDifrArIm10xTfKVVtV8qeX1SSrwlLD6/68THwAGbX
N8YH45tGrVDsZsSis75iauyQAl7bInyf/INzyFyRvg3J/G66lcfrEulXSkMG4SN8
7bvsBaDBnGmiElwJVkIi12CVA2u/ZUS2/CJqZJNoqcFLgc/byCI1nZOYcsq6HvyS
nv/WCKoMZ/1tHwrg9XSG0onAOT+imbXBNPFXLG59Ko/2R/wlDoYIHeUXb/65wY+I
wdwFQkJxv1KtNG9yQuyIuKEOPs5YiHbJMr3bGygpPlfRv2jJrWdagBThe2wxzrk7
ziYWEd3dgJTzAs2dAjh8/fAAZxeCLVOO/sWmpdYnBsKp+4KPK0uTD4W9OQH6+0Tb
kXff1gL0dfHNwrk9zZnZjWdnCKA+jrP21nGWmJeR9OcBnuqygalLzhjCYgzw7TQF
ceV/vo1Ol3UsPHAJK9RkfjCFioajFMWxoX/k3knqSNCGR1tDgCYYKGZ7eALSPzet
AHMHOpPWBD3HUsJ2pGsay9vtRz5sl8YBCKb18hgm0aBWUE/9jTqWyKfo3T74a5dA
HLgFD+sS4NsSgsBiH/r3/02jGMXbOb8nFE4lk6Ww12Hd38QLrN0J/X77VIUkbHIq
e2Sk76IimoomFTUfNDc9rRXnDEfyPh/neAfh8jVp47SxqOfwKG0PA83o7B8XBlmm
6CfEPT4Kporq31cDB/YbZ60txQNsskopIGfbfbqDnXyg5ZbLtq2Xf22enN5Zuv71
XCbKcRd/JqtaQRAT5eyWVXJDNJmW72Q7XpC+7Ej4CEBnpQEim1LZFwZGTe1SRFRB
oaiRD+0nObD6uVL4EHVpdU3zDYmHtTz/POC+PDxeKARBBalXPgcjoIcgwdanKfnD
yB9vKz0C1HaI25yD/c5cs8gt4pL89X0ZG9oz9t6H8hvZrEVNIPSPTllSSTsG/6dI
Cj7OaIgTX5xr6P9/LWK3078lPXIVFA+zaoS7nmjh4K+ywiM/eKb2wfPMcrM8L8jI
c+5tZjyw+3LwW69W74mXG0a/0fJZfSJ9o8FPqoy+27P8WjPfe3vIvKFkdnvi1nCi
9HdD+zfbPBXHonMEQ9gIk5ZJKXHfpxOpDydtq31X9LiIznsdkOkk63E6ENhTbxWW
i5/wy4feNZBMC9cU0bfHYQ5d65sGWoIqLJaw+9XB4vOonkjm2nkm+6au9FUsyTfY
CwuFF8GdoT7tqInj/XOQqArv82HVSNJyZWzDDPoo0qRj5IikezVTIiUJEBOBhhSH
+q7QN4wipph84o2/S6G8GzzaYIVszdL0+E6BJxI2vNi5Lw8zfruQELrN5qEBdUN3
t5zgWTrgJyeBBS5ygETe/HmUBHnSm25uhbWKL2QwPj/8tmzMNmOBw8VdXSzg+uYA
0fWTBAQVlAi9MqNETELW5jn0vNYTpP4/pGM2/eaPKe8HVnAdt38INSnKbZlP6mtC
MDNUIfTz73sRoVB/ipBlo0HNuYb8P7AbkBxsVTIGY1lnTzcuhaApi8+1MHLHPfsK
T2nQtXY7UrYsN7YTIpV4hP9EPmQ3luOnmHCHbLATgCR4LRXkztpb9Rq+/VHLxlZb
jSQWy7k7r9jtp1CIWPm60mUeopiEYyocpcM5U0NUYa9HodsG59qBg0jG+DnIUg88
w+jeeCSDIEMirNEgO0qs9ZHRXd5fLt5uhj+PUUbgW6v2lVzal3kBYCkzhse3Z2tr
5YD2f7QkYXeLVvdgDtX/FnZj7bzUvsboNGRFwak61hNWIHBdsoNQrOyI4wjJKl76
3LaA69EZdrvlgJKflaWI+MNxzKzkF67dl3KxmbtKqXSyGMgwC5UEbaeA6COuv59K
0Hly0pta9nczWnuVo871Fo7DqGqMztVEQYSeIjn0PmHu3dGAGlAf3zidEGrtG0Bd
fthQb6dEB0w/X5H/fP2vtrQNs76U0OJIA6mV4eOWSYcSqkRaRZTKDRu/2KWSDu+j
r8PgfA0+mlSzxAe7EO/6FGEejRWjLcNqMe3fJOAPZVUYrVwCEjdZJo9Tx3tYUtvv
UR3n+4lLTLTW6MaBNB+zNTHRVgpNDCfyG/uVq7Jk1tn+PS2gee0Mh/ILf7Vva/+N
fYF3kWKY+3+2zm6+3dM2zAkUPJoN3YZLVeo9oulegqkgoxBiAeQvTI7kmWpW13l2
7mMyUFG2u7t/tFQqv14QIh2dHFICPxsl/Q2PJNNnhYMAW41a0Ox79aDeRDXmjEbg
xFiCH6lEI4/2KNrSbNFiVwqYQYW3iLV8Q8LXXfv2m9nFkgXpKzC8j+8rK2oeCtq+
LaaY29Zlvn0jrk/L9HrFnpa5ngkQ42o431sPiwXL3ZUmG0y1Y9oW2f32/VBq8BX4
xOHzrDs/lqFoAj6NKDI5yyZLfQhcPc5p0O8NuAigB99ggZJtvByXBIBmgUrndQU9
pCpXNFiL+zLJ6Ve+92AYDs2PfrqGqNbtXwkspN7Y4SXoP2KwnXFj0ljOWRFQQgZK
SVta0UjimqHBQbfem/20efANyADuG/LrPNsMjQZ4/1CwQG1RRqCLVwdh5McfO3po
ts1RGR/GNIVNnUvZwO05x4Md+UgoCPa7nB0OrIgwN3fppf6mM43TrxMwENcJuhqk
sH/RWrgaMYwJrH0DQQvhMPCOUBfnw1CeESQ4SSnIGm28dQzt0NpT5UhUdHDCM/g3
HlQ5bYGF3CJurG5LOA7eodQ2ah3PN9HvKVQY/81ykkPEc2tMCD0ilvO00zJeEdPi
HLWuFjYEuuOxJffAbUQswLA7ZxFifAmNTHLO6T1H5JCHZILrL+NBErJ6L74rvGFw
vWiel7gieopDCIDTwPBsCLssfK53rC+5vs4krXqvQSWhldynDCZoS5j5bFiVwqUc
1vyhZWLNvAjVZrsAINlhYfnUf2wS/inNYRjHMCX3WndkJiyC90vD/W0I9UKgWbt4
8K0WeMkQt5ZIBgdX+udy23VN2H1AtWihzO76EbLIeKIztSCaf1lu1H3+8lSB/U71
PhRzWWY6DpESxWlIjReLxKj3JGr0U5Ei2b77Kv+j5mSPTFeAUj4+L8vI8g2bN+Q8
JVmupSQjqUC7augLOzHA+QC8JaqM6m54QcS9bgBCWWItJnd4LOaziZFSvwclg/Wf
MRydfZRunLHwCinawBJcn/Gb3BkvoFRFh1yGhAaZUmSIuoWnVzOv42BqJ6Ur2Gl5
p8NMBQwvMDDOmzYg8wmFYyZkplqgaKq56imIGAHkzQDxcETJDSIoGAM3wJOSYCOb
Uj0Y2MPD4SLtryOdKBOEeSzkrhpOxGjVMlIq/RIfDtT6NkxNMJXh44m/NQOiRdMH
5/ggE8U2+zCFPrTp3CBItzpkFxN3s6LHCXE0SYWPl1JwB/54dE68751AgN9baWfa
8gTAGm9OpKtppQ4eWhDo6Oz/RTUYcRywC0M7Yr7bIAcs0Jb4RfdSqbInl5GiYIuz
SZv0khh2mrO7+dbSYAI1d/4L9kXnFUBV8c6aYls0QNCqMUMDikanN2SCMKr+bWLG
yVKhBsLBFG+g5iAiv0zE9zqI45Sn0SPPhJD8lEiWRSLA6WBZQO4CszcjZFLcXW8/
IQOpsQjbGFJnegBhTkB77WLVKdiRGVzu14+6nLyMmd6AJhD/lcnsuNGrfSgu7eed
Hy9t+V14dsvhyMj+TYBaa4tRHPwutPwEOfdnIAkHZCLmE8VVP+A7Bxfxm1hK4Qld
4WhleYDHKTXzms7N8Jhg8pRBl0ot+tuWd3059sS9KDA43MzYaBprJY7eH4Lr6GOL
zXDExQ0/N4UOG7Qtiee3PBGwhTEW9y87i+R/4gtrUhHV9CqDLbnXR0VrXXi08zlC
s8l4u45b3iwFuhKzlXUY7B1bafk3Vm8+bhfoCv4l3+D7AoUGUmjpYGb/cGSA8/Df
JrUFqtuMv98dV2gcJwHXOhNH4jdzyxcFid9RgTt5O6OB2LM/qXUQ6JqiuLeyXyay
BdMpcTRYgtgPvM1SMd0UBi3PefJpjNIQ9Gsdk4Qfs0INuQVe5EBHd9VVW9WCEjKl
YUGZ3qu6TyXbnWv/sjGnJA8dy7HYDrbVWaVZAt65U05SjI2xz0ZbjSe/E3F6XG3p
iYBqAkpQbmTjhRDubAuQVSCaCTdO54scU3xcS4dXq+2wHQfr/D1LIZihZJxUaZCa
dG8GCbP/9aridBN8MQ+NtNdRg+FU2WX7EbZy1HFOJU+5lzxern8gRzndVYi7+2JY
MA5QWmd7tMw3nZI2FieztF3/tswVYSIR/ySiL1kbRV8/MmnEjW9i9cDuPhQqecIg
WJn9MUSTx9Z8py0YlRXAuUcp3AHdsQ5j0scc8pyZH4nXq7q6qxj2UqOSqh+8LULw
Gep/g0KBF1EGY8plqc2FdMqzYB9TWioY8ZszfuvpjXV79fgHrZe8VfYITgJxsrtQ
5YjLOaq2VnERBkPhTdj7josdCg1W7cx7mzYPzR6F3YMpvNBp0jrFqqN0jZ/vGG5C
x4fXsCgqF0soKoNcEmzyMMDQwJiirA7zPOXzjW2QOVW7gfy1BJ9xSWMO5b8eyYuZ
Cnb+VzRdK3CjaLOtuZ+poKXBZeveoJL4B15qlmVHGEuQ89lU8MXWjw/MPBWbmOb4
59f+m6MoXoeWv8XjpattJnxduFsr0cQO2apoVUWVkyzTjV8ctVf3/ORin3Ox5rT4
UfCJNklFzMZ3uPTyuTnfVFraKQIz2XnyNJhx2FYTzgOMKDRMjOYIl5ZadJrXio7O
tzcODnZj7gn2XF4y0QI//QKSVZtU11dpn5x0yWjOfs9C9SEws2ruj0IGagjDD3yT
ffC0QGcKjhYWeVXcz7GnNIwD1HchlAbwPqrZilA2AmNJ2SA190FUl1wC7RBKIoj4
0Bkghm2UegTjxS+HDX3orGrbMg/xI+XLBObtIw/a8yTS5nWVd9Snsh4E0gaJ025H
nLVDNkfa0P1T67mKKVO/bfAXK3F2oG1HU3cigi7xB+/9anA5APnkUQWYqiddxoex
DEYAIxZ3c87Vlm+uY23040YVymDtbqAdhxgBEWV0KcXn/GLqq7FsgBQ2OyF0cAvt
dE70UDwGhXCKmQLVlp/6/9l2N1MV/ih1kBRQXfqjlvxzmRMNGolX4XyNqht2BkaK
IBARBCRQGwnHJSwFwbALqh+X4zFt/yPqlAgnPKIiqx9GV4JpRzKs2pXUAMtSxHjQ
aB+lurgYRM+shzdPPrnKbLu8sTx/MrnLIX6YroUheqGUREQhebyEL+hCoEye+OU8
Jn8NLajeUbcW9RT+BT7G6SBPDXohhpEnR+vGEJEC3e47ehIPf106lvpVu61/lWRq
7vgIb5Wukn9uXAmsrxBRKndMZ3Ndj4XlaP4einlJFzoNn8Hk62xUMDUbSNo7FNzF
4cLv816ziP6DR961zBhhmz9KY2jnl1XFSpErEJUFEms53338MYjijvwcp++Zgu1Y
Rk4Cl/7avAHn7vpTAyw4wLknXcbZCI1L/pVPRfN9Mg3MNgAuC97oOtSSFWCbSsXy
zzMYSchPQRGonS6Zc82xzAWOoWZJ9A6YKeHijZz0TQHl/rIcq0e4OODUGrsbKycM
ZO3YJNb9FzzDCeeHozHmICNETwrN0dc4PfDb8HejxiDTCceGZI2MkNk/w0TGmES6
0EGE03nZNgXJxaX4aw/7IP25q6P71MkJWtGXl73Ukw1McGuj+N8DQenRnZD0G9lm
jjf1DDr1ei83sikuPc4n3X+1NpdQvKGrURTIpDpIv7T4m2F3flvKdpjtY0Hxt76O
BYF7TMPnEVPyj1KRgsRiw6C8QeFcbjejn6/3DWTWrGFp1i2YuHvf6v5cPsnb088X
xQ54izua6SappXZiZMdyPLzl/+sMU3zw/CqlfwDKdiIgsUG2j4Si6qk2/AzJd9j5
toEn4X1kd9nMI93gC/AlY1AqKKjnNJq788BelIoQteGs7GTnsu79vme825eEVMDL
O9T7YacnKG6wHfGjpUr/moD49X8MuuDdFCzRVJi28w/b6ZBsV2Ho4ebQ0KLU4+uD
JLp7NDyejUMr0LcO0iW0VtEuFteRiborviiiS1r9sxv8xTwJzJRsano4EyhXDQMy
YZ9guf/9CJL7U1/SpgT2QRriWIRrQuvLjQfxrV3px7D/jPxTaFhpV1e3FZcroikG
PdoXTt/uZ9KxVqPQwWXuFzAbZLEuNG8djXuMtZKD7fmFRaF/RdNvJNApMW+8ybYJ
gVH353uKZmfJUOOtl3zB6Hl9N9v0JopP1wiZHH14NMIYwE5GpEdLw4LOOIoL8BW+
GI/t6cIKT2sAdq9ew3UsnKEwE900NhhCA+yuIejESV2abeMEYQ6FAfus54UkO+l2
eNnfgHUkGLGZwrvt0z9R+lt/2WRftks67qrYDuj2QncxLVjrSNI8Pj4iNOMd5Ixd
1IIm+7wrUamgwBoIwIiijkWkZo7F1s7cuWzo+sMza21EAwdox/t6AFnp34M1rjfG
muueN1o7PbMHH0QZbuwSd9eI0QXoeOXVMF+fcFjLTqBhWeG11Vfit9CXwjYLqceN
GwJsdMpZAecCSrQraME7wixFTRwNRRwzBtCEg8MhQL2pOB45wtPSAx88iVAl1MFG
295H15pC/zu/XxDr2xuAxVGQ984WMAqbL68qsUiu/C1ZrX9FAfBDePGr9Ft5mxjO
TvwagPx8b3wDjniDKz4gRQM6uEcmJZlfNJb2vkMi4RRqbbOZdfEaQB/5/RCf0d+x
6+YyvnNWR79ryR+ft4JwO134cx2LUbPonhDL1tI7x+LmB3KxuT7YkhkGUpBX4Aku
kADPSNUQ7BMOiMLw9CBllJTFocrUkyrRhN1jQyMqBTSiHki9KLBiLok57drTx9va
0jbBE118Hk1tKgVMNWqnYrHuntiTOx8TX4nqAK7HjtrmeczNdcuV6guEG5biLdrY
FvOatHoundths96aaRiRgyKaheHhG7a4lJ6pkj0SFl4gILkaa5desk1LuLGCjCQg
enCICDU1Nggvvh7W+CxTDfoaJ4h4zObn2lrftDZUqpULfhykxVzarHS35mm1wL9Z
3HgY9Wm4BSj/oR5fFDI5SY8ISIKsug0X6MDPdrlw543dX7fUQFLXLS8w3WTYjdVx
Y3uqtexkejQzq55s2Gzw7uYjbH7kbwnfm42RK000jPiaGnrDVBXjqFKl35smUNjx
4UBwPnJigCTJfR+6qvf9MXhxcxau5QbON4xGXHoW+2vEUqrVJnbH//UnhPc/bQm1
ufjaajBOqQSvjen92lIzFel0pKjh1dr5yxn+ywTHMFpno822s5gu/DkibpGZITS7
0CRZvPHXPJj+Rkq9T3cstlojhVjYWdI/WEZZt16qP+KPuAvgre2N7b+iPnltIWD8
cLkZm0V2eSK6AuNG9MCMrvKrjn+l3svej0/Qe/BPebQlfyr/7zd2nfk78xcXVgvb
LNlOt1gsC03kYbr9QVmtUowW6p8fxHd+8PBLPRJFN5jPJB/2twHInmqRq0AEAduV
cyUjeD3YkUopWDiBh4//+9rBfZdGyyJZDZQCzUiLTD4nrWCeEgwN0Im0Fn7UPI3s
TKFsXrduNBDzMqj48A6KH5QCicqqeybH+VQilWhVYmzZdQn4QRDUOdtpjH0LB2uv
OOFkEpMLP5EQsKIF1WzS7bEuk6nk5Hf2GlXNBZZRg2k3iq0RvDTzf4DAAyzsSRgn
YRd+wrdv1UTsRqtZMTdqgWhnQot4m7XBstFkuOGAPFC+bOsJmke6eSZNAhDq/7RS
7B7w+9dm6NnCArlm0B0JDZvdKT8eNi4Lgakh7+s9KlMm86pAwl3uPFQQ2rp774Q0
LZ/Bzga1mO5qswliySdbj4Y0lwiL2+EVMA9i5OkA+F/Wc+g7Q6tdmJrmNDiwVbpj
NF+nySIol1rq2eyhREV6Kfs4k2tGu4Q75LI6JYO6oIeht1lPTYskYaO6mnsr5QZc
gI1fJBFYn9GKcGr2b3y/wIce7jergpuIL2q7TPtAwRXFfXGyeJW09WeenYj5ozuF
ZHHtUzhfzUTaNRrst4/y1jdsyiuGZFaL6ojyN3OukZi50Na1iVJYlYBdwpYWTmz4
BUFFzYdre2uuvia2b82tNFep84xZyuf3Anooof5VJSOj1pZPKH13ETKpNq2TleDJ
oDDxpwSKZuUekelpKXdZOkVqaVWfw0JIyjUo6GnujGMLzA1vishwn2ELMPxPxVz8
pQxAWLgEBp133vOeo2roDU21sYNPKto+pbFNw/iFH4yJfH3jWRPhoeEMjBFCGAF2
+DlzFTgBizUpqel6hufobKCjn7qhG48BLPiP58j3sF6zidEYZ2JfoAi8/qciL6/p
u4xbD4vJF3Pj0TGEVn9VEpQCYDUPua9cGPYt9/Z+npHmtZTgcL8qkrgbBlfvSDiW
81Uk5vMc/9xps9bPl8Myr/wan72CUfzITK1dKcGE7VGOlFsbp9s3W0x/eGHcetzj
xnle70PbQV38d3XVv6kvBDBA4oSHJ0GThAdn2zKpXMuJOFuLmyu5s9qOJoznLwxh
6Gd6m2uCrPty/V4KM1ayIAw1TJV57YXQiaGpj9S0gjQBRnjFGAfZVWaiI5stuagt
Up8exi5aC8BM0gda5rEtSjbFkiMeAa4GZoZcrGwlGvxtWY38b6iHd6TA5VdQQMca
JdVUWCVum723eFqnkChKuSUg+H+LvK36Mst71yAq4hOilN70Q5s+q9PPNex2J8sf
KlNoZ3vatBsUIPuKlfTr7xYHfWBfqjGovAfYLsUSMNAb6phPfnpu4708jc+ybSQv
1wjBAkdUlsmwniuXCyVAEw/aq+jjwMqyZrkTR5bUyiYk3I/t5G6XMT4yCW8Wcv7Y
JBNixeb0toTExHubQpaQPJ45Af9GsVGia3f0eqaTMnATvkCFovk+gSwPIXtfcJC7
dv86/USp+rg9NcZT3b94u6EtiDMWJ1sDbJCCDEV2vhI4ov+2LtSUHTsJJ5CdDsQz
p30QXfd2hKr3N8f6gPSYML9J5tUrlj+QjukcWU4dzsEnyPavYlVWlHkPgKfR0lGB
n2GJ1c4J2zBtQ4eYRSJhNu3rxxBKdsHbGN9Y6Ai8ztq4ITggW2IyDwuSJ7Da/dRz
TnKXC+/JRpNoQ12I+ltTD4ELPH5+qZeGQV1tSiY/9O2aEL+yXbcIzn0EUvFSiQpU
D+br7V7XTMxaWMGZ660pbjLGjA60N+wVQswHFcMAejOys1TI/BgcwaLjewQlFYZ7
DJqS/0SU6ZAfIHzFnJAw6pyqCMZmbKtwr7jqZs9y6WyUY6ekWPhtA/tyAGnDlPsM
G5RIdCerpe6pW/kxDnQ8pTHKzumbinHsYL6ysxXwM+icZNqY9ZMa3gXDVfzORnrP
lEpyRYefP5HFkWeSq5UdJuScxNffXffr+KWXE3iMi6pOHHLowGVrU9jOx2LoCe7q
6DRxC348UTS3Nz67GueQb93FQcuJLPUxEPT6QRYF2d/Pna9g2NLrPsbcozSpRGrU
suPKT3VM/GRZdKKTm96sIrvt5y05ikxiFpbAOBjCqok6GvxaVuCRoLl6+ErzV/N2
g5eYFIZxAEeMZa/DMq3eJETiRZnt9xg3voVhxhEvKymhPTdLFdc6Sm+Ll2yY2YpL
MUcFU10ZdYVMnrnSyL6ELnWNR3Gi3/SNcO54B7vY7MycIy5nzEcy5J4R5a06mgWa
mni+JJFIMI6LGzt+iULPVM/A2Cz/aSEzJatu3ifHeHD7E0SUyyrC23TGkowQ3X3h
wjOH9LpIuyBrLnJ5sNOkdVV/HsHzhlkczhtRog7HJZe+6952G++T7pN7Sm+5SHXm
Lvde2yCXRe4Pq5BP8x0h57tNlXKctTod9O7t1oHW6ewRVrRFAu5KpOcXSlHqdo5g
0+lfiGsY03zpflTe92+sT3vvW/9MXt3D6KWAvJoLe6tZOrH57fq+ue3QWXDAKn+S
ceLelzNMwSnixkPh3rpUrTwA9khsZPguK/a4PiZpSf/6/8KhoWk1SSKBcVunYibM
E02/+eKuy3tp5u85DUVzgY6/s9I97MkoW/cuJSGUqshoBJYouV1xlBnhSV6LZgVr
dUU8keOsNTnTyZsj4muStCLMpumj5bpT5slWyiOkly1NR7eaSF3BQ8/ZV+8CH8el
KRTmrYMI2Perh7JPcRkIhwU18PuZBSs1XcIdk55i4XHmvpSJ7DfdItdznn2gkRyM
qbhWTFkgfAx9ap2XJY3HjYbbkSslT94VUHjkU4I6crdhsL1oNTjieLOsu7A/3v6m
vNfizL+/c8Vy1QvP1+hPrY1mbyeD3ipxfNMv43QLEvfdXR8HtXQHuhU1+IylxYe+
HUKNdzQCsgB9/4FZD8lT/X+odD5o4Gq2S/fU2wPtUcDeVjqCI/OqdslgVNtUFQO+
42+T71Z7Vp+dM/vUQJR7o+1MLWJOe3esX7pEcQ2rRD1ACT+SYnU8Xn6gyjRC1vLA
Msh2gawdExRXENl1dAtSHrYo24MwXfjQhSTjModiaFwcbNOAL6juMBeHTXYyPFze
Blx0uAs5aNhl3WPSm4uxt5ksne8W8N1q8Q3nJ0og2xDM7fBAkB4LCdl+ZXtDUu7g
CzLdIupWgQtJsRyHxA+Pk8ElC9dI4BgMnWKlAVCPQ/hCOgwLEg8Ez2pvOFRst9SB
T6QfjOuldRvKpLRB6ifWzMeDV4GJJT4E04+dG3WMZ/+ua5tFnvXgDrRiXww/v2og
ToyhuSOOgRtHQ0PXUsPCs64hwTkyJgcgs6TSeJ/4nK5AkJ5mZrCUe43s+YSp86EV
XjXRYExIoPCHf0ajL2MCKWZOnbO8suzOQqHCmwxa5kz1eaCHKyClpTVNRxlCPDrV
ba0c4x6/hu5YTMxtTTth9FGHpFBfja/nguaaOh1WkAGB5Fy5mTfNpH4gZkn2Xb05
sShtWJ7fFNWuRXlYQ61Ew/Gjt/FYCBonD6KF170ONfr64LSlmkGz+ILuAq/uLu6e
l/sBeoxmqmCHuLeWW0LyRnneflZThV/ChgIpfRhI+Q82v51k1W/am1c/DVKyY/MY
WdKNqPJaPLP8wU0qCuRMEBdjPy0EsgpZLHHoMibEW6YOYuzsvjY8+ZSqtBketxyH
JWvhyHpjhuM/muUPU724Bf0YraEQUd3STqsWmoIE2MgaZkEV0PaHbciCF0XlBM5u
3JWbRB6wg5BdRW+DXqh0HIPqT8bRzDfV2o01tDo3SK2+9fUIL6IHoL0QVoVSgx6s
or+rRXFsQQciS9qIfiW0OtVERl9LRwbB49Er0A3f9t9jOVXmiEE676mjirLlwUN3
Jd582KlsPF9ZfvlTD4maxDBsBH2QrDVDCT0qod/M/AKUJ+r1PceT7LFlA9laYD4v
nw4I16HcHO/K44DA33lNPWKK7+n/lFgwXWaDtXY2pA0YlKk7fn4Lu/xW5Zu7M5cE
LrEPa+ABdLDG0t3eqMgiAm0bAnXiUMdeJEzThfmkM+9Sl1VBlo3yMpuiHfiXVSuU
6vn8YQHNGgX1WG+6IDBvh/R0hJJYYLySjMOiDO55shXtdvfFUplwh/Jl+ZG21Ymr
Yzc0HfS5k/M6bkH8hwJ19j2jIavyFSIj/mCaZycvBKoJEThI7BCvE3He9AQrCWh4
Fz9kj7yxwPqC+WAINafobvpzYzs70KBOI3RQUoTa9pivSHNIUVsN/Woq0EEz7O/w
NL4GlfWhXiJ4Er3ooOqH7e55YF8z1OLg9Z+UEynwZJy9EEmAqAiHLOdpHjSiJsKU
4oau/M5EMiobWzT5hNxUXXKYbg9DzgSH9alqceCrTPs20t8UuMGCpN08asn+Cs1M
YJbXWkGr8c0sq7ZkfhvyuJu5xPWrAuA4jPps1nMXTwHxo/1R01tnXvSG187eFbqF
PC76bpflrC9cTDvJZEUNiPXObT4fTf7MYqrpp15zjFlcHwbGPoHVahcl6Fnrnvks
RZRAi4zhu7CYx+1zgJxhnbi72sbFaj9jNXVfZIprO4rmv3+AfpUPeDadz1K3AGKw
2bVubpvFIzeQBHCSxlK3ytAqc//GnkI2bcWM6pHYtfZ/lIXVgxiE8MWTRbSbzzOU
9smjSnM2uCFZ6XseRU7MXS9lrdlHXXdL68xjEpk2X3m1KX5PkIf5fDO18f42B/Yl
E4ohPL9614NvP8Hb1I9vRWW6U1ta3Z/WPW3F88PbHVH/WNvoORf4Ui2LEH0Wz8+i
90JRqaLWFG57MPBKh5KESVk6xqCKs1Nnj4zWyAIfvF6UbBZ6nka5o60ftCcjd8Yo
7MeOvlb3Tl3DQlFZiNv6YGmDlXl+W0e345+WTjaczZOQnrZTZ9PRgzQZVPCxoYHg
Kmt9phMyd7XHBOCMJ+aQi8yLXwWmcSl23szkyI1t4qIrUx8rUR/MleGAIGvogfOZ
ZIJDqjgT05hgs1vpPVZabgFHGDrFBYBO1zgLhLBMs37mdQYzXS3CtIBxdU+Hg5XR
tsSXmy6TgqXVAxJ356fRKmfAjV2gP3E0+QE2IY4sNGbg0qKgb2YAhcIEHyoMnXgF
ChrvWMFj0LpVYM39dzAxhyQNucOBzS105zb7CIw0wZnXN3Rbmrv+yARbej9eMZtQ
ziEQv77UxaNVX8UdvaiDuyAaj+eVttrMTK2G79lPESzsnlojeah89IzHQykGJZwk
iSQbnwvZ0Wmgn9uZ+1AfjOmBVchqaQPGVSU3r6sVth82wH5e6B+jbXO5CjjxrJzH
PmWU/YX9fp6l3BOc+cGXKugykVeQSIkck6tD62zt+jFrsnzBavuOAQlI9yLgfRe7
xIaqQ2jWUypTxO2hhkK7wYptdW10FdqchAkGlUJqevHnDW4fMZRPdsNtEFLeg3lQ
H3SS6ehcC35hdw3032ZbSctsPrwew8K3pqrY8zZW6iKmxtzVtVeqTmHazcbvbM67
2IP70W6YfYCXeSbMLIXKUEBkoW69b1TcYr+LNHlDgMmQIlCLW6+7ACF7pRtz+AlN
l8vPFtPkMUJXoWnVaWOKTkJZyv84ureOFfeHSFYJvd+r0hhgLGNOfzjB3/5X0kB6
Vkm7Vb8P1b6F4CB71SV/RrA3tJxeXUrB3udHKP2TXTUoXAEEEZrTa6vRseeIriLl
arEUMNIv55/cHNT2PVfLf43IOIZHQKAsF6auTUF3BIrE5/sT32Rxof0PXpKQ1L0l
PS+NVsTFJ0ZeD1Qy+d0//4sFd6LXd2ldJhatTO1ckrpSqOPC38ebfycdve+Us9Pb
T4WU12KRpBa0eYxYgD73rAIH8zl7/SAhjdQLs/hMrbcibrbybl4JQyxihN4sS2TT
FkP52iVECRu5GjJAuUkl4N6BkMWkrYDm79yZ43mGEDT2FUabtBmy0dDSRUIwh1vQ
MNNxowtZBSpgLHxYsNz0bFF303hLEzwQJv2pW9NYDT65ucf4rbVMTaEgK6AAcV/y
f40p3cr4bJoHwRwUPE91/0hycI5krb0/NigqGJU0MHKJ3V39GoJF56V/oiEWSJ64
ukoQl3ffQMAt+32qiaeqt1ggvAtybWg3qkfys/quBO6PxWFU4EAs4p4qLJZceX/f
qR0/ydW85MHOZuBwWFiwLm9+ABxxs1RMVrI6acQxS2iian8lrZt+8GD+cWeVzaph
8DweCrrMlECFgimx0IBw1HDLmabk2s846zuxQeUTMBIlv/JL1iSNMnOs19+F/Oc7
iaAixE9Qi6IxwRkOV1zBW5NdcivcHieOV8ocCiovRD+KqrS0vWonS5SWbNfzoWyH
vIdP5WB1x1iujKlncPQ0Upn81wbV+KWjXvm0R4K7iKX8OBjPcCthpX8Y2WeLdTAP
oQho8iLyodtUJmAhPZkPW8mLPHi0/iMwUOSAVKLNyN//1TOLKi5XTw5mFV0MsSba
f3UrBTXLfNUZQbSGOah199Q2D/lTWQW/KWk4d3Eh37LMsjXOlZ5AALvy74EW0enr
024rYT43I4nQCRpRPndGmwRwVE32N87Qb8vWBYMf9X/9R+psSYLiTUq7hrMBmgnb
mQJ+eFox1GdT+MQ2ZdUIsMEavQGLC07HJzbdl3xSo7syQ8NJKWH3NMkpA9peuVQd
62YhTLL9tGLJWWPlRMrb00yerULVfb9gTQbOyAjY4131fNk/KGB5ie8LGfn0C+iL
vjw81MdICBxYKKA2gDm4XZOwpkJ2tsV/MJhetG3V49EwhUPxStOkXiBbyNC8bva9
8kfi0dR5v4a4tQcsBdXCRDhhRXgKFbcdvj1HCT4Llh4xQ0rW9YaSua5W3d7Ci07b
IVuOgz99+duCQ9x9JJfPb8Cba/Br5sLxIhqZcQN2n2W5zodSU6vcHFIWfZLxLPKx
s7KjONVVk6CcduGB4VhmxekIcK+fhfXZwCmX0XxfsFIhxmjPIu9A/cEzxEkqkbx1
TbSVbw5Zttr8MOtd38E6X47UIutOG0qJGW76WbtCMZQpoud4P9DzuzAnJFYxrzPy
V+Jx5pUuxkjqwNMk3p9CC8msij2wZT7gBRix9cu9PYm5AWSm895CoP8UP3BWEwwM
Zoe7L3wgWZrGM2hh5FtjnYaopVRqbb7F9FWsru9i7qaYEhMKZRCqaZciYQtcnEh7
QD+qXeijrTdKxZMkdUlvmuyrlnpcVek9R2fACrxbljeLXgz8F/hyoQ5gNxbUjAst
+EkNcMMneo57vvkk8o6JBqv76bITWLFCnWJTozuMYB2r6xpF6pFrdqvYzKXg6Ysj
jMB+7Khd8BbjOk55A8ovdF+yUCMyOImT6x8HaKMkL/lnrLctjLCQE0FS4CndgcDw
LAMzkjnBOmT2+PSl4nlz6eNIMg5ATu3Twm+IwxUXUDjPjzUWbr/TbxuwFOL3qIGz
6ZOOkl7Ct8JuJx0WzPTokcIYI6WXDY1HIV5Vk5AJPbkVOWTYPWkwrv1O2p+KNhHt
TblVSOpyuEhGPTJgXo7hOJObb66HSCy4cZMwry8CuHMEJltizfeSO0CZZmv6knkd
jg3suKUsbevqOIA8MJYuu5xVTjWwfCn6brvwseF2RJ+CiczGQ7p7iUc/7rXyh25B
rjhtHgoGy02HvSZQDHu32zC3Qm6oN9n2DE9PebW8Wlpgb28+AIlbGPVhCHrMzgDS
C7IDu5snpGMFe+xhaE+igSfe1HT12V86SCmNJrGZNl7ZLFvMVQ7SoQTV1l8vAzPM
q00UBtULPKZQzuf/XUmGG+X5AArrknkg39PJZUJcL5H45XDC4xjF4hrpsdRekoOB
scRWW2KQQjBdXmBIFai+EJS2JImwXms2sZVpcw3qy6s0U9ITVCIRlxTqFa5SXLqL
1Jg8WRInM4K/9ngD62ZwzyDhPqRR91EUj8sod1t/OR9mO3NLkyavQ/vYEeWm3wwx
z5DwDrLFB8CKUj3JWrYW+n1JJlzDLkD9soxg7fs383T5oqYXy03X/GJ0h7OB8bQI
bpwmpnBE9he1whPEEv6Bg4sx7CTpEZ/w6UMhOfTITd0cipUj+8kwiHynA42/LJRf
NrzmTboVOj1SX896C5d2ahIiKiOZoY8yr4tLMBWukFmELGLlGjqdA+4r8FKCchnK
sUaoPIYPWBP8bAb8M0XIrP+jBU0wLkIU3Wzkb5vPuJ9on1Igeww0UHxTieTwqa4L
4h7np8Jovaoc6Se7ZnySYnWfzV58YzZToopY6lRYGEpvWfS1hG5IwsxgPnjy5bOw
d/s1PhJ9wa8qYv+QIs1M+vDbAW+eHRlaLbJrYXV6Ipy01C2Kl6QgpuXmnVDGDFgn
HXfQCJoFlPZNvJ+KAuWoEI+ysudKNn+Z6fYrka1BsPQ+a29s52/k9d6KEcN3Uiua
qm1fk85MgLO9CZ+Rd1VUwTWUVMIaDam51CPSm855CO2veeTa4KOc5wkvdn5sDnQV
BhqBPPP+K+CG65UNvO/q6R8tmYJNXJrkMzyKbUPfPRlxCCOUWz/e080KO9/deU3J
MCi1bST/NKOQ+kwGilL4J4vHKupy5nX5V9w9AZgOr2w47dic94EZgs4fzIrVjYcx
bSf7DnUfa6rKFH+W/ZkBBmXQ3DDtaayrHPANGYvco2FJdmFJZyf9rpaqnBPFD9yL
Qr5DcmzPL7kD7NgAV0RQVFr6T0pdhCH7oVB93iwm+D2PK7lyS/gdaBWkr+5ma8J9
NjmoRWWL+ZXlClSkRJHw+EXKhfj+ssKq5w17OtN9sXlFh4R84Lu3anqR4zRbe9R+
DpNCrTvEziBIOu3dOyOGfE+HFdySNv0GyBOf0/oqmAQBI1vJqZyNdw+GAGH5ZUJ3
IfhPjQ50E+eZleATSiFTiUXxo6BaXvNLIPcASwEyhvGbCNUX6/z6jER2TQdH52as
0py9MKF3A7Hlw2Zzsl2ujaNsiNwxG/4bwGaFyFdIWhvI6/Z5KLfi3ic/e71p0jxW
r1oHLWpPkQoDgkAm4WPeZoRxOhCRBLEy4rCUPZxSTahbSFTMVXyqkM84zHDjw9VH
03M1C6EFx8FuQoOCBMxk1CJeUT3lmFvty5zbsFjldPyepShvQNkKXDaNSWhAgsvF
rf4k4r2SeIfXoCfJPaeXgO7EFYClvnbUuab3CH9CQIkUbyBnpCVVZFFmsZRpu18+
M4YmshwpPo8HV1/FyKN1s9wBmIjwnSu+EHs47qcQJs+bHWySIhnu7pJ02SFluZUS
Soxj1gtE99lQoyjgrT5O4qSrOst0OfjA+HHgC+2h2XKQVWJ+Sebnl5P1l7r1drfR
P53wd4LCNPuGBHa4tnDZA8dDacioPAsvSZz2z5ZCdfLN5WV8L8owu/mTqHB/91vd
YVywuqOr+bxgqtGZ+mMsWLBMBtgX6V1jdNVHftRAcxWUMfSm9CONMtVeSZyF2hkc
p2spYYBYrRfvEwLHu/nohu/8lD3iSzvwVFwi4Fg4Lr9OikpiOvnkC/Ec1kOsQCGi
LUw6HGoeZQL2hJSpNu62OsHQUPuKcrp5vLa/pBcPD8tBHzuehP67AKuBknK/wzyl
etBcEGM1ikxXP1P4WJU5V7U/r9vAxAuXXRCmWvGd4dL4GTvq/iEx/gvzUeTQS6VU
EIIOo+C83NUgYq9xjSrA2yPyuBeKCiv2//0Yz2N2yu/ecLm/ONHlcJZd+/bK/eDb
b4EipA1PIYIuu0QTDGhjXLsAUR7HQKBDXJQiPNNMAw/lmrYz2SMbD/dimGhWWC4E
+JXPZxZYLAsoDRHrv27OixMsVDs5a/i1FWgVia0Q2UdjOvyanBMMmFfnV3svCtAb
fZpHrh5Nc3CamJ1ir48mmU1hzI2GiintDb0Z6ko+viNXCNT2EHbRQw5VJEG5dMPl
NPpQcwEKF9aVyfk56d44CG3wvqUu9r90+zlRVkvEMUY6FuyPszUZXVznmauih/0i
mD7HRcBmCmPwgirefQ8sQO0O0uHM2BaJwGZl5hYvW3GLRW0qa4KRg0ie4HhJvIim
HVnUoV1G2U1dhBRmBLSNFdjUrXZYz1iPim6tYJw545b/ulKI6urjIdEkKydiH5DH
K1AsvgjGDuQfgapR2u82xl9zRWI+37jh+N41UdwTysou5ujsuZiSadufxpiI/fen
h5vu0opzNQLE/xcByNHksJSn/2tpYa+aP9emJv3KwipX9qHVL/vPQVEWrBULYyTh
xSfBkJCqmL0sG8PGElLDPRy8rVLC73P/H0WWHEhzh34InBABj1MC759MmuYYcvhW
Kv9NuEVm4qgEzOxVZu6Hmn7RCi7j+dAHbas7A14QFgPL2lckQtqVsQ9Od3pMR6wG
OXb1eoyW1AxjNhYLCE63fqw7NiEehqrhXkb6aFDUQh879LGnyoOEoxq8FQztsIc/
7MdYeo/mwXB/A5jyeUvNbWwM9JxGLkhq4YMg9PsyhLLTmaFZicllBnahpUzlbl6u
8L0Xlcxka6xUkQ3cqWxW8NqZdhc2TKJoSlByj4Kc+yLjuSL0sD6vKa9VplmVOVwf
xDcXxKmvMFSt4pBc6SDQf2m6cwjeaBMycpEMySw/GI0LMzTQDn8sKq0Ssi6ySkYQ
0JuRhzikJvbw7s6hLjoTgGlrc9X5cdxUPuhDtRSqHSyHh56I+FU9rLRyrHY2Fa8S
HyTkcgwF4JHSZ7Ip2ROfH7Cyomhnj46RwRjvbQA7J00zXoj2PU4WmuzpCuMNOSX7
fwDnLbym4RUFdEThkm8jIsXZH1sXpc8xzKtDR+V4ZZ5KYiGTkDvIz4ZPqp5WCooc
OI4bCZs1xZcFWhdiQqKpC1EOUFr0Q0R+Wwr/FWz8oftwe8KBFIQK+ssYCfeGqW2I
j+DOhTgI2Wsa3WUhrNGQtBXsIIhL7zssHTc8Absthh2Bo2Hs0rbIg0fSKqccmlst
Es1Geu7ufSIk43S6W7PxUeAAnFIT8f1n6MHFdFYoZ+9cGGN1C/DO8gWIfDfrlkhW
Au7kCtTHdoK3SRQN095hw7qbSAX1aaz6AbQ1Ab59148k+nU3to0oAkJLncA7ViVj
uepetHRH1pCdP2DP3YnBy0SKtGTaVmBR9IWnjSQ/iSYt2Qi95kIkHeP6+gO+WPz+
dHacE6fGBYMEZbe9ikFb0e+MokfE04mmtamFspt4jw1AVMgqzzp04nshYXN+RXR0
ACP9OaLXfDhRcrLeYyFXLWrjhW3puLEWdyekCPG5oQGHwOOVSqZLFtUJI8sreuf9
X/mjIcIdGGbZ1cQKWeCF+4Z7TrXMCfuE+0YZyax8D7bRTPgluev+bA3SUwxdlmM3
kKNH9ae2dwhbJzJZmPwNrGjnwQtsLDs2mkCYxZshowKhz/3JeNgNA5MoE729Jd6G
4Xq7qxjSqENLuyVMu/2geAzOrQCoohyQNN9Y+huPxObty0snG0MHrptH9RRcutW8
BYCwdhm5e4PBHE/atPCGbp1e6DZQkbKWZQu0pQJqYhC5baiY8MPZCVxwIMH7RqXN
VRwPMV9srhHhgOVddHF9zc1vA0pRPa2wxiXsKQHOQGrNnHFwNZf884AU74BW27M6
rtDl2wxbmANEsaVc2ThyHA2r/HeW7b1V3r5mAhDP3pMY56mlXhiktCwEXecUB54x
WukgIDh5dBH99eXcYHTIMh4j133QlQX4qPp8b25n82rDts1yzzFyfFMVqgSCdXTv
KXFmP+8vuk6wG8c286ECP2MEpe0D/GBcQKGJMQTVaj7qwsHSA8YDsuN6KF9RUndK
R1r7dZzuCixiZiT9Pjyg6qXFYqRiCtg02wvzGtmUG2TcXrUxOFPfYvcBzZIKQLfo
j73BISNUJoJvp8eYU08zZcOUjIRYrT5TlJUIe3iI5zeSVisGabdL/gwHpnYzYrGt
qZztYDa0kuyjtdtvJU4/BrPxCF8iXeToEiNVuNGNEfJBpV/pRlZ6Uppz4BfVev4P
rOoZKSGW+2G8ePLkXcYqW53u/B88WRedJjmfXCKvG13aPce3sPHdUqLPfKBYB652
rdaFf40cYc5FLRLOdycVjrK8xQVw2WbhspIMW/BU82bPQMU//YZYAPLnT3iD/gL6
TsAM8x2Ldbj3bRIJIdNh3thIY8tf/hRScsvpzxuuAHhlFeVvCyXUEXoiuY9QXFBU
rBph/+HvQS5FkqyaXKTusoXdt9en8Ib00i+1XWKahycKsIgz4Zv1lUJO8AWE7Ofb
5U6XaqCBkj50HNZZf1K932x/uek9hRsMqHXd221/by1rM47bnyC3v7lEbhwbLvav
/nXSP5/Qq3weHnXngp5UAwb9IRNV9nVjhWhX//KUBXRRxYZ+yY9wQp3/o93duITn
yAJhBGYp8m2vTUSmVK0azkZzTe8xtUFeqpjJYznlNcAAiSeAwcTd18CCJE3nupMq
DflHcFS49Q1RMpdJyk+8X7HnjcbjPX4/Gy1JUgT9HM+GYF79tUMFprjcTvmwuMsV
ZnRnB6K1IEsCVGq6wwWOX95KOoU2deHzdtZuOsfiX0isTq21GaTRgmFF4Wql67Ne
6hR2rtjcwHBT/R8sZKBNmCvuFzeHmFMxcMS6Yz0a+D7q/76rHwOS1mvYGVd4Dbg1
MwLfG/Wg+9/VUNEfmHaRVWeAZxNcKotDkooF1G54QcxcCwXPwRIHvwdEdJGDi1pk
kJpnfB2/HRiy/dD+CuuUvzZMxMYgZaUvu7wvD5zCipSbUIzyEMF78dwS5qTYB1TO
Zjlx4vxD2rCsOaP07A2k9tNK9wp9TngsigdSgzocdA7A+xjkZrniL3+0pIwpKEVh
WJjyKAscVqEM7PhpW4aviTEPqjjvlhQr2xiVHAKHy3Z3VPQfYx2WQ+AGPJynbzfv
ZFOWP4C4F62b14VNQL+lCAPS4H05+xC76jApWqT8yU4SKbh9JQ4fwgKN8PRkta1f
vLTL0ZcM6qcNcoKNi6vT0WQkKpOU0kNAMdzYa0z4sVyQIbccE4szqL0o4OEmIyRP
Y592RGLUy/GLlupt2YBkDsC0k43mWR688ZbGIbb6OWqgloT18QtzBKvbwA12+37i
PwObC+9SWB/7EsNRq8Yoo5yGRyHkDW47YMS9zAao+BlInsOCYJoi9lA2eEXY4Mm9
HaUT/K7Qlq2pJuWXLpqk5BwySy4GH2cVTslST0OuhMZmBQG7A4EWuyKrn8O5D/bt
Cq9y5ynyaoB90gkh4T00ZO39jSpISdsTb+pqvgKKIleluku+b4F1j5GcXvSaPUfv
GG8Y5JuCtlQZp6SPX6WUllFvZiDt8VCygQAEDdotko+ZLkppPzynehutwaLWWKx7
N10FBGno7/PWQQtPmjgSnzXL423o0C0PKLrvgv5g4isz/MwFbKq3rFFM080B4Ce3
bbRZry6QhmVku73MWjabmLeCd6AY7PIq++2tBaYMpbsxo2+A2Y5Za1njnjESSSTy
XIOQMQVIBW8LtiQm9EA3ZYgrsL+jc5JmC2SRTKKjXkwiL8HCRHxsGJ1y+d9vC92A
iL8Fy1gSP80jGt2gRyQyxNP5PA6q5+QkuGQ0DVDE40/xG1GaXfWbzAdITrVlvHn9
O140jsIGVEEuWdsFPHgijFNUeDGPvhqxZMw6xFFsIzUdVrTVUF2Fs59/gjJNSqiu
RhKjne73HX9bsmMjD2y5F8Z+zLksZtP3jNkNDRFQe/qpkc/TlsuMIPAgWdvpAy3K
q4gpwygEwud/Stc/8MKXgtwKT4/OKJOKrkTEGItWqrHwLHtLpcujr+Zj4sZeF6pj
0fYPI+Gv6Pn/v/xJz7m2qnLz8CgHKtu82Y6n1wB+J8+ugxvsCNkKAOM75PTKBXSY
sEio4fzOfb6orAvj+JOMD8E6iToRRqr3whCAsh3OBqsTjCZA9WVQ3kbWVPYVItUO
gUlbKew2utBY6MCfIPuSicAAs+rtgNgf/f277wlLGRQ+a8qmblAOE8s8jnOl98SJ
B3y+dClAJ4Gkkpxn64rU+KX03Gd8+i912e/eOQ/OEkId061/zDjul+u1zVzdaaxZ
K5dzv3VRrxknKZw9xR2Xj0UIpiSKjWFlYSnccVewLZoLdzRS8klRIr2XIC55ggkf
/iWJtrHfsqzz7LYDpEHCtjlOfFYqBg1xONaYaNPFP+HW/TB7G4XtutHdm6g1f0LF
y2XUsB0nYgvmyYNlYVML15vXMQ7gZx3A5uIIUjm/gOUjChlJHPyGJVNAmTbec9E9
PWeBAKt8nAB3tvMNh+8HjKveqEgu5mEPD4AKkAyd7JAe0za/1hN49LHlyVsrmdB/
GtcbXY74xjo8xkBCx28EafjMKavIW7af/v336exVj0oGPqQAzo5YCVD93jNNha1T
nNNVocVuMHJObMXGG0X62e2/yS2bkPV0oYetcTvwJgBfYjvcH2SYFJ4QqA5Yosgd
RNszomW70jll+w0GKOMvLHwfTuphMhpyTM9TPT3BFgu5mMB7Sd26eBE2lxaDqgNn
V/B2VKuaDuykpX87B/18cOn0rl/lv3UUvzz1R2oyL+I/yFirA6KrCvnIOdKMiEmc
Q4Ge4+1hSg9msfF4RoGLEw19nsU6SMQg4rYNwZ5DT/4hf56iaiTrN+Bei468HoJV
eBNSFwUhkwubIhlUkxNNzOea74CWfJan38gfTduJiaIPoZNRtKS7X/ti8UaxN32c
Xv0fIBtXxCLBXHmKJC1bF4DTcJP+2BhP+rUuIvz8HfHub8C3KjmZgewR2T3dZ46q
3PGFAdxLD0eBRnSojhUWfzHyr64QjXxmjzf8P/WRlI0YyF5wnL4BBOY5crZYoVGP
gA0WPUvfiJ/BHZxARUFnOj2Gn7kKM+YZt8a8H/URSsa5iytOFt2PJblCAHPdR3j5
ojAt2ecd9FJKfCWKy6O46XsTYEfHVyUYC+TFi5zI2uw677/gE21Oxb3WPysh4KJ5
tU7sevZvFUpPO0GNyTRx3DjRzU7qamrEKNeOyNn30aE4DsodhLepoH4wDanNwNbY
AW1kQyhFwTxHQAK+p4vBIUnUL1DHMojvaaVjTPKG6SLU9jf40/Zsmzqm8+lNMYw0
bxUZVVx74I9/Yznx3HwLtEd6/6Y7v5S97s3q7zqa7swqdjz+BXhS1eOD1ty4hKE/
5lbv2y/XO4b10T22WCwJf1l2dKmJV1q4HfqzGympkPAVKJcvePeiVPPEUPCrEe2Q
QQtXU0NXWjxDonHpB3WuS6kOahNRySBOX/LqjvJv/61sjJw/IfErRIau3bjA1/F2
w938YOoxzdIlCjRJ45Owt5Y7Fbvxkg5E8A7YvdiRJ5PKEDsfwLZ5R3s7oBEzwY0A
t4N44pCI5Y+wPNZ0RBm7dMs57XK9Zs9Dhq9yJNEgjr+NUWmiXg4FVTwz+c7QVbnd
NgWuiXQf5WQefBb8bpZNw5Xm7E3hlbQyfScCPk939zxkQxMmEjokCFj2OtKIvHq2
LxGSCl1PxgUttTVngOC8G4gwnc/hhAJoKHySlRiKEpyZvy2XM5YzK9AXlPkWgHeA
tnGFLgBhY1QbCBTZomfnpXmV0IRnobtIcA/6zVOKGq+c+85wsukN3ZIaEfWdSr40
CZl54Xk7HuQO6RUEydoWoojI44ddRBhy5/gs0Ws4CeFlw7oPrnxcUfqGv5AOI//m
6DYAks2WL5l5Ja5kepSHs4QoP6L4dg3STmGTi1VvHZsc2yt/MyCLNrlRzvoraaFL
rHaKOwvq+/2FDN6TEj7QwBpUyTPwlBRKKB2Mt+QksNwErdZobPxcuMjV5ac2ZW3O
OwtDhQJN1GqKhT2d28bv3IcfFRPsB/Kj9jVeQ7wbvyce/qXbtFTDiLcQkJwTLNGg
QJKPh4/iDdOPCdlxaDpw3m3Xx3CqgVNryHR2X2visMj8jbKOx7RexI5rticksv63
ZImMcSHqv/m6xkcPY5A9nbN4/ylt8GudXnAEeWIS4U14BT4flYrZVUtuk1rJuFr0
49gqjhDVvQoB9mAh1PjVxcCv1IHS0SNrcjWoijnhfVxyVTlsLiuzVPr2fZkmP8Hu
y/A33549teNjvGJs7Qiv6XFEj4I5wlkqu6UDEW4iuqAdu1GFu1tLg5XNCoqHdRTU
zwC1huLyueiyKNHitXbv2lGn6Vj1xzwqR/8+PnQ2B7/C31JzFdwZC5/VAbDFEPRB
nOrT63RdJvSNBW9U1Ig9Ij/NTDNzkRHhCYlwCkwojZG1I3B/jBBjtS+ugwcQQ1/N
TSS8sRRlBbpYB1hamzEGIqKwC92OzHdG5wdUgfGTC7svh1LqHNJbKRbkTpss7y2E
5ac7TtlueqO5T9x+vmLJgeg7UGCSHMginR0T52L0tQhvzQQhUyPsz43lU3F9xsVR
k8fWVDuPcIR1sGqAd77Uq3jYqRTYPksBAfLp9+eAtBb31ATGx3s03O4nnvChrafu
YAM/fxGK5EwxTfQbQSNt3ar7vlgcknisxgBDbKzXh88o2mMxn0lPhxjEYydqHJ+P
z/K2Z5SghNJXXUXdKDioXTxsKTbSsA/IqwhCJJKAVPVs4mfr5uP+tM+oJLdJwZkX
A233e9+wBY7CyF9wZr9/v+6pWQupaIvxJl6iV4FWEEEV4KPGeBRXM5pnuT6rGG2t
I8MRswN+BmRfsGguWeOUsZGZ0bHqwaroRYBM6nOk2gpA2Tn4e6rlmHhn4/MKcBnR
qEaxDnRFSM1gshkysljC173YTuyk+WEfFPMOvRi28UGWLCrETtmbgn+dg58i8V/1
5pwg6p4aH7a7LXDSMYpPPTUEiI7BYLfrW3AZtt4w4nG2GlEOKdpAzokfpf6Blz9v
o9LX2sKRs46Q1xyYupeGcx7Yie2kQjRtBfSZSklV94+3ZgdcrgrgnG51b09pMtYK
aMJIv9GHNlDcfJfi6fFEAUZEYbROpSqsU9Vw2rdx54JUH8np9B3BuqYXDNcNHmZ7
MZAj2FFVbM3Nv+AU2N7RldyLsVloGHibLE0CaDhHuGeqFGn8yPOfJNH1od8zvIyl
8RHDzNyroK8OGzq8Rx8ZZSsIheQnr+MB1vk25vH/UW5eAnPM0fKFyW72Hy3ah+v+
TV+CbvmIC+Efwr4R8XutZvJ17sNGKo8qTaTIQk47ul7f4Jy0hzXE5H9gqy0enggz
YU/njkrO3L2hoYI6NYW38I274X7ggU/j3sKPiEJjQp9y5bWH3vFzIYWjNP/A1vwb
IwgA5OzifXgz1YdIzwo5igY7URVs//P0ko7mxPonDZ/+LW7YBXqYv25JOlz9ifIC
3mY6y5/DpZ3SaK2WC6OLVVz0mS0nfssa+tivcVuoLWYxzjwGCqtK0lQ4u1qvclDk
RIceGWy7KiMXhVZCqDQxMIA9zx9r/DAVcx2hi7wsXisibNaXB3zrKhVKdQ3FFJC7
0XYRifi7+3zbIrKo+4fV+C23F9n5YbTvuK3HWbsiC5WyGfA5v2u66cOTxpCfhzG0
IH84m/S6xysTMp0Ej3UpX2lalDDhIENN033tyU5YxbQj76p7hLmlaGxnUQjwax/B
nNQKfU8NrWfUNOFM7b5eB3vV+9VYdU7DPjanbpVbu+KE3wYmBOiycgjprDhKBIfY
QV1cgDPUpMoysC0b4FmRXto9u+e6CUtJKySGB/papASgN8IKDF+LKxxx8lxJ8fhq
VzhlRIj/ur1WeJgH14dxaKuvSlTgY2T1CKLwtjRqbJi78agcGpP4byN2S1nA82Gh
imH7Hwgk9DZyJMlSME+IUXskjkVkhXVm9ktKfg8pnVdsgyreopNvvHVSuUmQGozW
KqaoGgrv02cQjYVKiOHypC+JeWuUwz6WUg9aPHX+Q7xc5pUplYntv0ytElaJH19r
EdqZzZy0yx6MOTq58jyANTG/evbxOhZygkxNh0lmhiGucIs2++RnmEcuUlVSmw0W
fPc+EDSGO4fC0blmq8LN8TZenQ3jCjKDI/rxLgfp0bGIAQYIxe/f+lCpb4ECXmRL
6NNVvxFWIqszGcVDZcmGsCyc0IftHqsg9FcidUqVQfNqn6ebZb9F0d4l2namGbYr
uwU3xWIvc94SQ3MSSoQ1rXqFIsHZozpaqlatca+WhaGuBrySZpEsPlCVVNnnGVnQ
tgcKwvzO6zQhs8Xee1NWTAQ71wrgRQ7g2IJ1noWjgzou33QDwino6fJZta0nYzrw
vkhIlFTp9ulx8n1Ym5TT/8ytCHYuzxF9Zty87JCDzOj04MzJ5ZeJoVpMVDhu03Ze
wDpgz+Hdu/2TkQIud3vHyAj1VmkeZVYBab7BU/G+XSXNzwuMPQdyE3ytzNyFelhd
ofu7QXQUfUIZ8J0JmEzp5s0LShRE9XDQvKHL5kMIGDdmpp+WN1sNvFViLysjFXw1
5dXOCDUuBrtUcqIuy37ynfG2k0UmLL06/T/ibvcy3B3LbBkLpM0KI+oQRiVYrVfH
6FH1sk0gJA/b6e5qOTCaeXjBZiapEBrlDQ+9f2+SDsAdEvHzMUmEqGU8GZwFL1MU
ZMGhuj41ZxLdCT3s0vGrdXhfwaX2RuhNpCiiJfeRkDEGuZ14DBr6100yHOj8E5Uk
3KnGVN3lhU4+9y87+Mz6kq2pzl7H/ICT/k7MCl1ON9p3oKmkhNuQ5JUDO52y+2xC
RfiCiA+5xYTtQ6jtDeKEeh2aahOJvHUCiBbtYSIIH2bzwtBKvcKUAXK5BT9o8DZu
B/g/QMR039KuCkvwLQ6I9dpyxmy1XyifX6zV/BXkN176uROL6G99/1qtun+fojzl
7sK126UU0aRHdqNKduANe+gX03IIvDsvHJp8B5jxuHK+tj9z+zVwGEJ5ctCAPRLY
MBUCsaNRl/A5m9r29k5Be+MzzWijwPOeftRKivJbl0k82dN7i9F2zoNFH+h9VbHI
F8DlMezfERKc9KXUqlp49cOc2MKD9kNORp9Br+gCKMDRwkAhanjXGCRx+CAJ2rTL
rEjgmSNxD6Pj4Wr7815raqqbICNec8aes4h2k9lQItCmXv6OgZPgOOZsj1njYt1V
S1dU74g/nJGPtPP3CeoFNXP5wlTNG0PM8l1Ch785mUntFfB1S59nPJAMRjuysg8y
Osakp1S4TGTCKEzEeEtnXe0t51RVVXeXnSPl4F/GpFN9ltdZ6//mmsx2KDIZcpAR
Unh5G27guhlLT4efUnPOPV9shsc8OQ4h12cNH1eedWT96/GuhOG+G5IbGfsBKUYR
SdEoKKpRHlDtVZ1HRlM8MmqhykEwACw3QM7D2ve4pJceyOX5m1kfrAQtVwXwHC4I
Om+Et1K7amFSP1h93g5mQQiRSDKilCx5zLED2QKR8VS8VSVFyAgZlxO1vXOldHXD
8Ncvc3vNF/1J2kYVD0hG0l/itEFPBG3WBL11/orSQ+qdudOBDZUrZKtMxDaUwyfH
zZ5TOaNX/isBWWC3j2+REpiFyF06BzShkSWMZKBCjRtov1wLGDvw4ZyEdI8+dSkv
2UL+8Fqo4csee9V/I4KewibqChkW0NfCKEmeEsn4mc/svGDj1Zu3LeCydncT3Ad3
67afRq2C0HOFNmf154HEvCgHJYsodoW30hpSLtJknNSkuH/jsXXop0nypj+eEOhN
YwndUUhtC5TV+DXJZgO26ugwe1txRcua4LqOCUsevziwWEiRVHpC8hKIFDL6k22P
9uFPikcaXFXLtt8PaP0Ou09OfInoSZYEyruoqnkPn+jKvTIT5YKQ6SB2OdkcmjnA
aZC1PI5h84cOlpPu76bNfuwO2BmfO+OD5rx2DmW3ahbUC6HwonDFmQ1YQWe1z7IQ
jI35cFRVFPtgHZl/pF9qZu+WMZarBcbiyogS0N8lFF0i1RNnWsy+0t10xwRvS549
kVpxkLVzd7klGw0967ZlGwvUmL4UQcnznyWJLx72+14lMxzxbKaUwY52q6+58QN2
sESGKWJPVdoWidcICoqFzdprDFz+6DRfwUYyVMfQW3ZYavYX2XpyKkEk4w319IFK
5qlDdr6gTMElAg//wl3TJMGNvRHOjrCUyv9SRFmLWOmoVNS8u5dR1f81WG5gX9dn
GfK9iBpp5TAYE5cWxvN35lrlo5ISu7oAtd0frqraI+0Ry18Sls38BmrUS7qrXKjQ
bkZrpykXzaHVjHdBrAZcEW5KSTXuXMzfVrfdvO7bJzGeVGzgjIBnFB2yGb2o/C1A
97JMISSbFlqzXttIPNVSuDlQ1JGEdocPhWNzB1kKo0LXK6Pt8Sfwvjk1c7FCzrkp
uPUycocxSmf/FosBEjvVmivsWhcbJRYQ5B4yjf2dy9p2VxKFF88yEdyGSDVvgUhJ
tdFaLikoaVaYsGk4zTmGQ3E01B7KH++VL+g7JbKwHwDM8NTJ7+ldzhzBB0JaTaRr
IbRM2jCryXn7vlU2CsVRIl7+tzJA6MmoMBJbu+x8U0z3zyJUDLAsJSbF+S8YTVCx
6SRNENdYD2295bswKr2tdNO/fW3OxszZV+CyLSSSTkEEdLai/I9xNyWFfsIEngf/
w13mWlI0YCG+AH8TizT9AC+x5fUqX8NLTNVki6+HfRWmDW9C2YTbpFUmgHSgCP5l
j77GQZ6y5SJD0BajZrEFnluENr7GwpN599gcFUahlEL3n6zdVXF8TIHcfSINBZ3S
rFdlGqzkuloSevjQVMQnuDgcR/InJK/t55i+BUYcBEH0lZ3b0GKwd4WxZkGfGLog
uLn0Q+KIihovphnMSZCxoflLBAjs/pjEmp4PLVOjUOTdGfknYzNwKw29QUh/EKjb
9FPLqwxB9v7cplomwj4RPToHxgATNSSqcMrxrrv3zYCRY7qNnrlyq42G5qYjRcea
wxqNOBHk+e+5I3/14byeLYeSpUv/N0YLOQFcZppCf/788xiDlADRJl2uJsIGxhwa
KZU4kDagbDikWiF85D/5Wzqy1fKS406y+KvxTm0gslpzRXNYuMZl9nWXPe4MtNiC
YqtPpsCRtns2iyjfRWvvJ1j+BeUHkoWZ8LMzKA4lZyR+ZrcdlUEaebsTz59MRSin
1MMZk0IMHSIMouP67X627p0j8cndBZAOUXC9YzgQJkJ3n6cjSmMN/woIPbsPkvtJ
QqZycEf/vutZa2n9wru3STqExaVnMIL0Vmt+uwaH3BrqDtShPJXq/pMN/rQCPOwX
gR3khjSk1IqOcD6nhh0xCGUwTavrRpXmq4Og20XHHbAAJoAi50+5PXzL00pubAnP
rT9x1WTnmD/627ogkV2UxTx7LgH1M7VyKs8D7lnYTBa3BOMgnTqvRQstgtIZ82ax
+ofpu7JZZWnBy5SNW+sGXIFbjBuTdXS29+pEuN4MkO6iCvQZDMATxaai4dV0FWhC
9G4bq2fOs21ac9JjIJH6INMqTgjYi/l5ysb5bblR+JldhqtW+A6x8c/1wBqCw3TU
2z6KzJawV+TkrdM7lu10FY7yJlXVg9WapIEeLMzRYM3mK9ZVTGh/HLGuNfbBhLzh
qXcrgv0wRbVP77AgldSHXjsXhc2WvMvnDOFHvHme/SuiOqsbiIOpR1fBISW4RrCj
Yz4KQuGw1uPWvQJKAlcAe4ELlScMNLFLpDBixyzLVeOVaeE6XmMlgWL77ijdg1pr
iqPZpgj/zO9bcFf6TCUoBKK2VHIWZC6eXWKUzh5tTb6cJbKBibPJ5ZH1JI79oGwl
pet2oEbW3c4cBhfqxFeinlAdDFSjYRwKl0oCCyIV4rZdU5TiciAucwZWBCyeGEvy
BoeLT62C6o/w9LnVrP0DPOei7Eyw9Bnv+8Q8MZ4Hap/4ioNXWg9U7DS0yL3qP3Ck
0jWPvOVbzRnNNW8z3X0ZEm/6HWnxfHBqxpYWJ3bM6leC0alH+hugNRBwHHKEWa1H
aaT3XcNmO8IsiJtZFfei2J3YIHw4OnzfG5dUEkvAwhp0Y1w7IkNWeWy67vfkvdc9
yFOYK9qE/+UfeR4FpQ4Jy9VtGAn1HjyuWpTTD7w5tUxllCFgRk5I3fpzsGGcMliH
ELal561UrQqDDX031PG+GSa/EtsdRODOM9kGDSFAn83JZAdTzc3y7SU7zxViQSSZ
/QBZdtv2c6V115SgRscBnHaPGrhy5aIrhS+/B+OVQlRpzDmtW8kQGwXyxaN3AtnE
hxuw36XtmIxQ10owtpI3sdpF2RE+rviofCEAZpPSJ5OU6pYP+NC4fdWLbJ2/+3aH
MX3a+vs32+9A/+5EuA8cNfq3KWEi9lIHqd1uzeAGU1ES62gqNQR3tUmX5o+346W8
yPZTvAk4rMh2y1Ip0U3IkJQvsV2DSI494cfG9M2BmJET8CwUcesaxj5hCMlFzX/L
sgmr33o1tc6C2o5sUil49r0KVEZciFt0F76OhHMXzDIAPS1sOHwwycSwXcnxPK37
IYL/cBJwrkOdfBWe0CUOcbEXf/mBzsKvSFVYDZ4Agad5qAYa7UsCi0hOC+Z7OPmT
j3AqA5LXODnO77rqqyoD6+jN15+EQ8ekjOHM653ASFVCQKAAuk/379un3o/GjJOx
wGb7flEK3ICOxdZ7bNH+BoUHv/u1n6q8W7O/tJuu+y9oU+TD1f4pJdXpPPPps/i/
I+LEwEDU+oJoeyC2Dj09x45CrbBNo3E9MDXb1iVEUHjfT2xijYd7jzkkCV8cMZvI
kEsR1wvV3dXysQMj1bmRrCOUJDCk7ATlAaCeqNhPDefQncPuKR5a5tCXrE0YbYkN
YZaTz0H+PFgJ69BjyCmR9P3KGXF/je0OQQKES37JD893zWF8gRdXRm0vLxmZYeYC
UYre1NBJmXVhIi5ZD8KcJ/tqERqRhX1DJdL2lvn3bjAlv9Y9TM2q/31EfHfpFG15
ue5t4hmUW2S1tHb5Z4tVUOWxM8xE+CVrg8j2HdybDIY8U8F3SbGnIuNWguAK9Wvt
dHzLN9f6y/KjTlktZtMljoFRmZhYyBzN2d8jSf+Yi72j6R16i8iqs1qBmVvU8zyU
pI52e4qPrhjEzTwFiFhl5nBM8cmaWwtBiaeCJGUnp+VYxK17neIlpp8l/aW1BWrM
X/A5DX4+ImWNet/7gnbF36oOKJGqAqRyW8cwI1GVNaQJEPRxwISXZfOYSeJq293K
PbSyNWyElHKmqfLRZvFcoI+cS+aOFDUVP9rDhV67zgGA98aUxclY4iSD3Rjki+UP
xEvrYoAp2lXC9nIdc3Fc8ZdKEiNQDCiZw0/JxuMIPpIM4mPT+slia5FrWpmwFwPt
gWhiPx1szZy7MCHrKj5IrOlIGBSiV9WMHwVemGSAszx1jMt4DUvXkKl6B8616OGA
o1Hek9gWYKR9TPhVHulxgAIt0OL7e/YFFoKUv6LvqjIFT2Re7BoeBJbs93WH6ZAa
jFaa+FnKrNa1Fq4b8MYPk/4GfuyKllgW1wWJ4b1JRTj1aQvPPY64f/rlr2qu5I/Z
7uz85+mZDMzAa24tAjK2YG8Xn5alo04AJoQHO8ZnoPZPDUKuC3q0hITYsnQ/hX8o
j+rbxfZ4Gnm+D2SyfMZtrabXlJxhACHtb90jAZcIzSMqUl3AOfOOPXZj0w/p6lV6
CUf4MCQ8ni7ljFq6xuAz0u8sppGmLUuXS3hhLFGLd3kNvWOkzy8fwNn22qzn/rtv
xgER3bB3x9nY8a5E3uIpoyKPmKMvbP0eBEVYMeewAwFeh4uEfgBHCL2pzBuhMWLQ
1zeb/BUl6j576Ab9krcE2ah6Jxq7PN2Go0Zl7uJmDndvkI+lY097dPIsz23oUv2u
7BeHsI+658iDXONjfGA/FBEvryjUKBDY3zUKCTdkmb/IdrgHZHS1l4nczqzw4MI3
mo21kn5fA8U5tUayr70PBl3IG+Se4rq/TTl1VNaEHvMpBN+ORPR5wdXC1NSd0B5s
QvHAwtal2c+s3Q5rj97emX26CdFCYPZUUrhGkFVW3P02Ebb6ZN/4jupxzgmSCd+U
npKCPnY+hGB6rlw59JDyLH+7NRQZIzPs02FHv4waYIqnA64xCNXBTKUkYm/1M7w6
RuHP5a1p5vAA0mxuBghRUDSMIuDGfL6YERiwO2A77CqVNJAu914Ix6Jwax+xo+/y
IqlRfRuaynYkju/TlW4L1c2QA2vtfZ5BqgURp7I4Tsdy4PNq/r+MnX/b/0J3wseP
ltQmbnDt0pJCMaeGDSA5ridBziI6IWKMNbeqEueAKbgAVdYvEil38PCxwjETvUGJ
okCHXp1Ry33xBui1PYGK40+XA/5rSWTBcaqtk4WkOq3kGwKEUoh0lGekBpW3pWbW
Tc2zRwJge2XI1Ng4B0iILsk+oOQacxXqWJMcoD+JrQDKyVJQXChGtmzYn8vGK/fg
dQocoWc6UHgKK0//8MsPFGBV1cdSnkc+di/VTdyfUQcCuHuqQSKDHKsDhxIyPuoI
87N+kH4xrTth87S3w0woRc12JHViD9GCJ65bgfQkolVs1zZMiYej7EgIFK0SCyE8
YIbKA0uKd6LawUAop+SUEsgm9zmFlkTPiXZU/2tJ13ajog0LuSAu4mpOt1f4t33D
6QOYRQsnIsGblcobOphxRIYqFyHX8R25Wau/rqQdZm9CPD26pAmhTyc4Or7ir+CN
HwKTCOsoHJn/My46AUSr3ASvvKzdbPblT1TzpdoMm/RipeaD2W7uPosgDay7LWbO
rfXz0w7uMZludyS7fA8cUFrwlGqo6WzuW5VI0h+InM7McKVF1lcmru0RlAgrJ9zT
IuZV0RJ+pHfx8hcsjPYaT0GiN+6YEJA5YcFQA4NanR+2/E3R1c94knQBDdfgUYgM
viNN9U4f5po5KhGzPjJ+UhXIw/3Oafq5uM67O12YTG9ANUKR443e3ZM8xIHy2KZe
61lbkLGS+jc3rm7WdgRmAzVb35UlXya1pj52m8hf3L8f/qyl0Htq2rjhH5u4Fsaw
a0phHsT3o2li/rK63sY0Xs4yU3P7A7BXVi07EOlabqHZgDzN+ezWKWhEtM5VSGsE
lNXc69jawMRZ6nMMPCI75JjsGzVJ2AGAW7Gw5l81LDG4ziy2PEHoFlJY+W9yYKvU
BQGvgyB3Z42G/pmfmA6Sf0KhIl1nIlXkRGuiB/RYJkQg2iGanyP/WVM6LhP10VKf
06ONLA7+Jb/EYHmuKtYCfV+dc21YKZfwfykvqjhPsDGu/Xybaco/5lK4esVlSFC0
INmACe62Qk7HjFuv8vEhCNzfVxZFN7xl9hn9WJlPSC98s+d9uxM2nQ25MNg31zHJ
x9NN0jQTUQqN4tw2+uAfH8XTeL/Kgo+J5s9dWqCFV5y6IoH6lq+Im3l8DXJwaI3Q
Fqw0l/7nYUJrvICdzlDxe+m8sPvaun52ZWOY26dLzmDPaObooBMmeZTk41l34xH3
SvGlZXgsUEHWJHlrOlFB/Y354nOLaVOkQnlOuBlTMX5v0Bs3PrtyE1lL1HDJfpm3
SlM1hO8mjpiINaGaqALnqKxDJN9qXtkK3HkNjO9yIhT7ohyayiO4UAXy9KibpQ3B
2DwcI+tiTHgLzqvjBlMsNK5+hmnSxarmeCq783dlqf/SqQ1cvf60rz9K7ar7LN++
ooRHZkoEh0QT4RYYp/m09ESv/AFHMbMHloCFFMuyCmekx/S05gHshMNpjH2r2n+o
cN6ZHB/Umsw4Uor1knrlLHzpSptq1tBsUBUcbfBE7BB1QedSPRhSorgHs1ebKV/N
RQaL16BH+QdA+ChdKQfNCymlGbHIWzO2yp6D9L+m+bPJTuvmRhze5K8T3RUQv9//
+s4I3Wh4feKIIT/+NHOXeu1n7RglyoFyGw8gRCHJWUvAi5JDrwYEyG4oYFg/35Zm
v6wFI8Er4Tm9hGKYaGREE73x42ddC0OZx6fQBkmdcJkW5TwoTeBuMTuqshjE90cb
Q4o8vbBgzj5TmCfnjl0Ye0JzrjZcze4Xbkpz/YHaui9u9ijJSvxy5MwbVydQg4e+
SZGgvVgf95tjrZzKUm/Ql/qmWYHrOtXjCAV/0MSC294UqXGJ2xgDORNwStbHZcVL
GhQmBWR98HzqSaYUTmbnLGXE5y/hRvXp4a7u3XmASc/v/PrdV4D86qLuL7xbSS1e
HB8ir1nMoS+rrqzRYS3tuJsCmPaknHpNKeh/Pq+EWz4giDEc2ltgO4MzZJiU8wBY
/T++h+kelVajlnFGSvGiqShVY02TTaDi1GybDM4LGHBMC9hrQA5ztzt7Ni/lOr78
jVMWXUS9G6j2od49mPwDwitWhLdtIQFzV5CDDPtWYKYRyFyVumTfcjrF3kStlyqb
hvBuhP6otu/SskesUKEGUxgyln9r92AdUAjW4m7dxKaZ1EUB9MohCrdSegysIGjL
M89sjtckd147z/vCHBiprmRoIZzBqryteXK7tRQXY0pVjGPg4c9RX4oTnx+kpGac
bOUE95SlD7fVuEPPA+pENTdkRjR8QYhLKrrCVEQl4SdNNmcBFhcal5t9Utjg7y2s
wl3acxH/UlzkGoXY8oIhaZ1+ILqXomoeEcDFKcpY/+NKhIhLuWuBeQNTBWg0+T8A
/Z1JVpiUiW98sASqRsSo8qv+2I5QCFmjw5ZvhJ2Bv+wslBOTRoQNUV9dGo+h78/V
ZRd32ZI/x94rPijJZyItUojO8NFbG8Aol9wo6WopPLcLcHIV4ZNdphw7FPAf3Y/Y
ihHQA1XIOxgoKrdEafcQ0hun9DiKR59KQLYhMMVHrvMU6TltGrwDd0peKZKu3Ms+
wg7U3mxBURcZ0QveU8ehK2BStnGN3OUUPxSlLK9zOEoG2b+ULqzuWq2Tag/dMMWL
pKHgVGXItEq/5kz48cOrWptpg4P6DhTiqxtYszEqnMOwZnDmU4sc0Qp6ZN2O0JSI
Tu2pKvPG6JRjT8Ue9rkO2kx1dnxJPKZeCSfENBujs1PqxdiPEPYsGHor96cVoy+r
gWXtlXSkCRrqxYbC1tfnrwE9CgmpA32X54H9bvZH6obPgaOxrp4H5FFngSXy1vUx
1PJJ4LnJ14ZrYqIMMHhVOCUSWSHgrHt3iT/WLbuzAPLV/CMFBBowIadT6z3CSeSO
spII7uIr+12h71UzE0NfSARsG9bNP6+aRPlfagUzOqv0jGzFMDUzkP02iSA9sfYI
ohMnGdIVnMhx6P32fiXgATc+7wPXmCtJPD3aQN7uah5Vhbu7Kcaaf6D0PU3UQMzr
gH4Jk51KeiJb3mP8ggpun7j334c30vFiaVbcUe4HUy4zaPNFjOXVTsbSgDOImX4Y
adIO8pTLeMro8XuY6m9ANP8wcMLsLO9evwqAwp2CTS85R0kmwaZlj/Zx4h+0sct7
bvZ6C7fd3vyb/J8w8u/Z1GDMkIm8HYTa8i793xPw32mHDjdgTUEuB6Hpu6XeOZM7
jLVMglZJP32h4RXJuSjZ9XwSfv1huoUGf9TUqynbo+gJ+KaFAjfzKOzKolhnvjBH
SX/9LRYZyM+3df5o4UcnUiHsAw12YWuA5LU1RrwEXYcXfjORZl4BK+sTdgt+OPbb
whhko8AqxLOWUCAlufwGDd09r1Pnx6gsxy+ClBgkX2C+07siu8WN0cqX1iy+moL7
wpBhTGnRq+7GgcSfDCCIY6vHO523Xao1kW8r3yzXieVP1StU9UqHEKJiIDVKd5Up
M67YrY1Lc5WhP4Yt15xWQ8nsemjyflnW0qb9jYf/tz588vyqlltbku0sD69uCKIP
6eAuCZUPOYCMNfSlGXts62NcPyjGKdJ8+9r/WSghDgGcH6iGUvDPlXtPZXQEooXh
L+FSD5z8kRciaemVwXhaBJbSs4GVu+g6/EJMowSebdRUCtSoKNFzbMdZe7XBU6hA
UNNaxTtYNv3WVPL9ijJw9wuFRRrrjdP98G3fZ6TkKbnxvJvxWyLl1lvJngb3Siup
xRmTBcYvKLLmJJgQUApT1BC03vTgdoZ0ifI73W6reADWF9UD/3vHPeRDXOTadpYq
8DBd860mnr4cBzMAXwQQN2kcqPXhU4wPs2Wc/LOPionrwAy2Zy3YLNGKoXLYMkDp
b2SfPThKCHE28x3UWaS9NrPGfCZGScmoEViEjd6nCYSUtgfnucN4R1KlwwZefNFF
uHL3/7Vp1CGblb+BTQg7nz7epVYPAwjtwOxLdps+g/wB9vYTotaiYLxOYQSaGrdO
8PZIKE25HVy6hkBSCvWIIWoucYS1M9uln19Y65sVYFGrrhgGpqivFqXj+qCU1sCM
uAbcMSWuY/6GdG90eUIcBFPAZV/NntaSuFQU1p861xS5M49FqhAk9ZqDwLTD4PF4
xsqw6fLA/GAojDJlzSswHFQ/c5m+YZnzF7brNm4rqC9u1uV7OZ2hvRAU+UgFfqq7
oJdTrD8GzSIkACYiDnRUE9Xq4UnJWb6h/3cqiPgySa1WsXwC7H0bhGd4dnzICaJS
qiynb4gouSTHb54BjleWe+vn4U7OKKoTaTbrUW/XAAG179/UhhYhsDcbrW19Yiu4
OHvcFZMCcRCzTIutHOhWExCA5MdtuJAcgReTnUxFZf/jlcS/yGT61g7X+jhsjAlG
06ilD+J1dIWQp+NZUuppSlbuXE0IMuHU3R3wX7hN9SQ8j5KM9ZgoIt71sRLmy3Xq
zYkwPybc3tZALXBh9D0WG2atJQ+4kDfzjcaRO7fRza/XrEtpYn6FyGH/Mgvqa9jf
gdexZ39TqyevzAf8Xe/4CNFyI++IifYGzdxZBAUh9FRn/A5pA3qVQfP468563zm4
JRYA6ZbvLatyLjfhbMdegeSeANgEK2Ocd4mQPSHBVf3GdzahUvFCxI/rJiKBFoE3
T5H2ku+mmYhyfS9iqpxzTgvsT7yAoNI8PHJO6XOwoDOu1tHX61nMEVOdYlDzYzkj
eQ1dkj7bubofR9cmn2TOnZ0siHL6OXJUyazWyX37V7u9PbYwjjrgpeP+GEaEBZ96
xWT8WUpa9GVjO0nKzGrVqDQP0RvxY4qRq+GzWJHl4wPjUKfiYflu1sHk2iXxBr2D
8mSfwvhB09CfJkWu9ZxodnC3hlMdZoxvD766VQAPsrkqBFRoTsuCtopJASKCIUdw
XuwGnOjlo4lXsGfMA02PTlFbeZnK3N6f2av6nmL22J5AnHnyscgbQPIZpHl8zrNB
MsUeb61jW7yCMrLu/UNew8TF0svELlzPsm7jHE3lmNldbbwLukigGn+q1KpM3Tlz
8xiLIDQzwi9MOWBX+hPFUTSbDPDaidOk0cojMm52mRUE0oj25AQYJ0V7Pe5gGsCV
UuwipyXqM9eJUgSSyHqa0Ueam+P18GzDMLng8Aicac/WyNbJ/cMopPHRTmDYeMmO
+vVPSOoGpiqx5/MZFnjRLG/Sk+KaS1J9daofVsYo3Hav8ajvbqcWvAlM1MpK6Hb0
4DaJqbJCfHkXXCcc5rkXyYoJdRMrJlxnHAGmDD99fAeFiVR2eR3efQD8Y8E4WJXy
84HeMT3zP2ypHlxeKgktHlUymzO+PWc6y2aGnSu+xcJrp/+mDYse3Hu0iVZdzEZI
ebeWNW1CpctscUgjXUaDPaj3dDoqAQM2KkPpCMG/dvruHiI9NmKY52RfBeTf54ye
JHSanI+F/w/F7DZ3s6MkcdsUFB9tDdBoptPF0FbMMYJYoi5AZ9lsTbacsPBqJ/3f
hzq1aAibrw26tOtWoIAmGUhNkvQBGTjkA6XmxyWYZbKuIEakoqrSaaVXm66/lnyg
isnyiFzptsE6e5svJYwe3mlLcgfTOFOfQVjMoslndadjGiKcsliXJPfx+8CYL5vQ
BEtxLffEnAaGi6sJNcpJt9WqVSzkPnzphSnI7veZvtykca58nylkXpe1qV0Zu5KW
9iMf2kywXJUYzJ1QV+RhMkKm2yyBnLCUbIsznNiXvDsCkdaLhotaeiHp7djHc4ND
cBTxtFou0W/UeX2x7Dru4VU9koXSxuCm1XrB6btBxvzjHlzCZVEpxsF0zLBXoBHZ
/N/BajYXQzfbDpMgwHyD46Hg+bO9nWN3BeHOW4UlVjbJAuJdgNjVDMSAwGeqG6Ws
LpMSL6E3v8D5o+DD1DG+EYUT/X+aKnIQ8O1tWhVgs5Zt8qF6kMVVnDrNMDiHk0/t
y4TIm7Od26VYDNzQznnNp7HHZq5nLLcjocoBi6sda1OHjnZtSyN5DG74vnVu/0s5
+zZYOYwlf5qJ07n5eCrLwFdVeor+dogrzNcfDmcKllULfxHv1f8N3pHlXtIkTFN2
jz+LNQ3qFC+vuU9P2GjrQGmuFI6foI6bhLJ6l1RSRAyPtcnj+TIjATx1c0z0Rxap
xnW2dc1g8nwmcrOMSGQOBsmWlsTWaF5JujkR963WN4zGgw0+eu9J9hKxgEoCfey3
U7e1d3dkTcVIEsZKATkIiPzJLc242/Ddxj+c/xLqFP310GMF0bFy6uMK5W3wLg59
92TYUvX9RWFUC57c8nmPcXNiobjx0YBPuC2VZ0STGlAoZxdsN+raywQvInYDOuf2
8FVKPdxcSMkoHMcGuoOj6tJyW9E1pKV2lXSyPH9c9LoZ4e9TfOzVOelA4Fly41O+
rZVbLLSgD7v98uu25uuFDe72jD29fU9ghqT/C1zFRG1tI+tYqANIlCEQEUoQrXAP
5cX6KLfMqbUWWG6SYOts0cBOyrVaeUZhrbey5kMw6O3qDoXWz6kLEbc3zjOYHA2K
ok1Nz564rDzUjl1bkDAvYYyu0hT+rxfeDXag+5RGsrAxdU7WnbHNFCiGCcb5qShQ
2Qu5NrVfk1h/eOTtmYwugs+XuTHmudr4yarEFhSJPztWzGmdFJyTh4KDg6JPys0m
NAyrkpy0NjPVkm6503LO0zfh8eOwmWn5rWcXZ6UnWbdNpJCK+1PEau0F5HcQgwti
r0tg9rJkJXw8VGEiri8jxykfP+rua0sGpZ+hFg1yfAdFe8subd8LFyK9rSwnmN+T
Yqm4FT4K8IS+3ok+oOVwA0+saypzlb7W56SMHN4C897+GF6Q5AJjpJcQATa6OEh1
Q2LdRap7NL+Nxv4goC55MDMFnUH39USmNha/ZdD/lsaXOVgx0RdWu7ifd3CxRZF7
Snv52a155R5Izi5tjAocRbQoQCNmIQAbLClQi+p/cG29fOzMBMQF9NUO13T82Hv3
QRmxlAr1bMh6HHvrK3McgfP5tWPPPwQBGrVXZcWG0QE4rQBiFmpXubRAY28eer6t
bKnAjTnwYicp7x+VSb+B91Adf2ItaymJ+8aC66czGypcXTPhfsfLiSF6RoPb1wdm
qJwUs3iMqrVjNhw+3VTLbPZVRgzrjt9UO6eied30Iq3guK2YWAVLzGluWBwBZQUV
1NOSQu7xck+GzofsfhEVSSNmTW0fQBHvQMrkffDL+Z6QrQmfAfOZLsPTMLg1BrYD
A5CUM7NajURYomUGNyxyRCgfbA9WTc1gSlBhVqAMGJJ00FCSSJUtGfC+HJLQXfm5
rkcA4RR2ln9rvofq4+4HdAkuC0HkUhxUlJdvsLz5HHqob7ZP6JKKCzMCG+Ei8JHi
qk3Be134TMBUugvvD7wXIBvPBugVYnjrEj6O48FtJiNw3/NvWMAcuihV/+x0jH4q
gYrDZbdbx2FBh1aZGq+8y3iYiyE8lwC6BpXxPUxKABIkPiPe+c/17v0S9K9hYuC8
TtfY89NRUcqGN587006jeFR3y1ci/zHqRorc44BZSTbx6vDAOIlgPC08JwNJi5hz
Gs/bcLmywNi4eLJt7k7mEGMB6CrYddbf3Ldh7Gkfgx4MiIh50bevogbg/QIEL6MI
J5IvbXICf+LKJlMgsJYHQ1ntKbUKv7jVbmva5GDnYZKSMZxoE5wY6wmfZshOEbcz
AjTVqoI9iwPIHBqmfendZJzS4XMHj++B0qPNT2V+6m1MuPrcyHrPQuUKuf9+k6Uj
xPZoUaKgYkMHEgaBe1abdoj+m9ZuufbC24jwa9rHJkn/l/zdjBmXKH9LGF3ATzf7
yoKsSn3J7NFrRIuwjOecAq19mkietE4fjh2hhAsETZmj/zQ5mYhH93Sxtic7pmhX
rK+Asd7DPWot0powxF9G+Nnzjsk6+8QteNh/wU3955S9IARXEdiJ83wGqnDON4Xf
fvZVEvqiV/SteoOj8ezu8PGwYJp3Vly1mkiUoN8BYw/byTjDigTWFITKxFXZOh0h
ubkWmc17VHkRq/UZE0lICJ373fFW93MC3GkpucEVO8vDPfz2rq4R76e+buNhshev
doRzDg0+J0alI2ZSZd2YGVyWB6/rzKRyX3pwTBkv10h5MTQn4E7Hj1pQpTv3fzwI
Q9ufWmAOvNvREBrd1t8fAqCpoAt5lNmG6ALNAliREtGcjhmEuoFhJdYbsytnXBK0
zKWu4nQaebU81NoK6FSb9mkyduJYxyZzzrcQjEkyy7uLKAG2FL6/5lgwXNvCGRRt
jbKuHlKNpab+R9jAV2Ewj+bi4a+pxcYzTv31f+mhfvYDi/RDmngYyr5S8aUbItsC
YaMpZeZyhxhKolm+oVsnF6QBAFYK/LXjZPhxerjF1RqjZJGjciO23YBh4k7aTUIh
uaV7i8IF1a/1J140zATpKXbZIa+bCmMp12kAIf07KMn/qQD5Wb6M6WdW3w6hq7O0
TmGlKhGQsI6J2uQJWpBPoecPHNbAO2I5uCsnsJw9vYs1DAQwDbW5q4idNPpdzpjx
f5ZHuHIiNOhoAWvkYoR5oWpnAgX4Ughi62X4yuwG1MtfeyJUyImsh81T9iXsX9OA
qxsHcf73o3PRga0mQnCzoJLiXQIpH3zlJo/sXpki3nGpKskGu773mDjyiKsK0fUN
zpOaPTBGF4xt3wR0Gznr3xpy4oy/YOnqH53jvVyfLEbEmqXcgZtSTQYd29//GPHa
WoByVDLim59H/rOpK3qdCzp+CUtVj4jmqRh3mZhlTZ/6wnVr4YT+sb3YLOwnz0R6
ttNv+1CPmciH9/xQJ1lyvCuT08g2xd51C//aEoVDutTf7+W91iGmSoRz1GNGl3D9
fGxqOWW3vRJSVO8eTaww6BNLBpYzOYwX5a82gd/p+DMLTjWlaFbO3lzKTAmWc13v
ryhnxPvtYSUNioSxOsrxkPeZEKR5dzQzXHvikXQq59s/QGqmdsPmefYZNQELf6hp
j6XowU6Nr5M2W4pi7a2lve811+q/dpRQVn9WZdm2ramyqQCyTSHbLq+QIChjWqPF
60oY5t0jDu9al31FN953OUgANAaO70DpDq1vEukIbwaVpaaH3uFl+gZnG1BzjL/R
xWDR3naXNIJ+n0ltwdiG2cYOuEOrDltPk7OrdHNV4o9873+AK4oLyieCMsmtOokx
GKZZU6ZyPLjN8a9NoUdWz85An8TYISG6dDlVtie9m/vatb/7zTmGmuB1z1DA1MCN
hG2hggq5UXIY1Tim2wGY9I56sX+1xLXEP4hUYKLd/iXiRsFCzAHHAoCQuEuOQv9k
TA+x8To7Xod6jDrQtJDbx48soPMgBwcwFMnBrK+DKklgTli0T5TqWY6hSFWUaU3p
eEcvCcmdJQTidKLPq/+gm4LXWU8BTKKfRA1dPg9lM55lrg52Ap6R4mM9PHIRF5XB
lzgKjF1Bk8Uo4F9A749zLGnvkChuVpC5kUlUmm2Hl3/MRYoBMi5QZVTPDcaozK/A
5upY0uU7i6jkKnfCLRP/2+/2mAIQqdc84vxE+yztmCHSbFI+6iOyBpATTsirm/B+
48INb5YNv/iKLI3TUY+pyb1g07lF81rnCbjot2Ap4A8OXs6SRsYAETX1yvGLwVSf
f7zYDCZ88aA04SLtsNWuVV+vucHxFoa8yOAeypX+eptv1DBeUO4e3A+BcDd2BiwI
IngPwh0XYGcujlxJM0c6HCUcFs0RObqPip+Kvhvcji2jvoX9k4cm2xcvXOJNHTMh
yu7QW03WQgKG+eJXGAGl42ksriBvIGboOchycECR8OjlGoEb922bc6iClEvKutJa
UgGIPzGErZCNhLnjmAdu61JakVsB/bYPPuRcXOJydyYQJl95+1/AUfG2mY/+dS7i
T8SKNtbP4nCCSe1IYH+xW1fsh0yCztSg114BUfIQCqE8rDhn4AZftDz4yiZZLXlw
nt3Hm7GNB2bYO1T59zAusYwCUQdPrklyLIigB804zeEm+C5Pk4v+jaU2Z69S6jhP
bG0XF8XH14oLP8D0xyqDzyO1XwlxcEFcwU++LwkYDr7ZfiP7jYjHCypl7zUs/Td+
k554suOm9Vr7ozOCMHaD7Jr521M78SAbuo4Tfd80ThWuQhjkOQ2MLjUeNJStsarn
rJUHgvdf34882EAXzdon/Ha4sWeY1QDI+E4WCQcipibyQyGyQiI+OWD38wSygYCk
5I1Gmhjv8VuLBiV8AeIeYpoaPEbhWhgBsdLMDHqCwspL0Np0AqXFMpQmSLAt0s+Q
semUkjKsVGt7/SKxMloZDD5yNhxCm17zrLQogKaOeseo/imFKSS1pqBUr2FeXLfG
/tVCSCB90l68TssZaag2LbQ+WR62pJsN0JBvW0YTemkOZaaVXNSIX2cMywhWmIek
MIc/3K9CE2woNNG50T1sKHGGY2gPiSOldKDRdieMVUBY6BSZNE0RNjhrm59LOsat
Dt+e5Sir5FcV2Eti0BmO5/PjvwsRWkC0Qh0HhbNGM9uEOOfeY/JS+EiLO5uukoLM
+U7TEOjXWaCccmMAT30T1Kv1ugvjzA9Skgr++h0RjPwdBts3rXtewxatbN+fdNOl
gsd/W3ut8pi11A/3km+C5HufLGFTScuub15+gAnfAovlVEsga3fCfSjl5TE2iJDY
S2jeUlpO3EuchjMfJ1JJfvPzUGx3np6ibxMm0ravuJiE/Th4FfVIK4IsNrkJplKp
L9UUaFLXfS+ZkNs83LiLGfEpghRCdn1GTz+LN39ntaqVGFz4eOGKwwMI3qom/WVW
m47rOnBOegoKOcAIvclrPdF4XP0b9h58QYYUr1ceYHi8Jly3+ShDXk5cN6vOBFLD
+xqyEiwyCWGOuK1ShVp6m3KQw0JFxqw3NXGY03/Uh6mVlMPu6nLmKk4AmjZd3Olu
8tB0dw9xuVkQ2nAhi/kTg7VH8qAE4V70Lq3HBHBPfd6u/WYOgRt4siY4uBVuY4ua
y5+rG+PBUZJ8kRXQz1j+DGU7eX5PB3l3/tSn9OkzLa2kB9Rq9kxWrs4vxkp0i6JM
k/+OCoJwxZWh5NiJvonblKy4h2JGWFEVxkh59NlLOYmaVGeJQ/9uDStDVVS5/Iug
nxnM7ka1/8MARHR8eOxN6tniUijBaFaCZfgbsBPHZKyXV9lFAwEqHkbXqCKFIGex
jq4ajkEXPcRQXM0BkDHi41VGgoLGC+2ZNRf9DyxX8Cm5iu+VtUhFEFSBvvZsYCBm
38iD5NDbtI/C9WeihFPZYK+3x4Y6xU+f1YG72Ypym7mfyvT09IgQmYUBYym0IE2A
FRt6H4QeIZAXWGnT9Wb6qIg0xGz5kgzG2irYuX2a4qRfF1qBNC+3TSjfO38AmcCK
YPseIM2HmfKrMA/UHR3HzlJe2+WNmYd569vXihs1eoHYI+PxPM59bhBL07eCitHz
JMQqjScAkl23/gyOAXu+MMtBrepMiey8MXBWeu+CMFfLJKH47ypouw5y7UnsQNBA
bAnboN3+4pdp9lQVAQDgd4evejNaNfkRqjgvAcDkNItThqwttX/Q2DXgI43w2MdW
Uoi0OG2gRGUHsUfKGIVYEYwZLbadnHkHqhxTAfsFguC7s9SyPkc5nAA29S1CW+m9
Qek8ozvPuWPvVYe3fmwYElTj89QfkztrUfIFRL9+oUfa6hexT36qfap+pSBR31OZ
a/UHTKTvycXwsh/eLHp78DmGUQIxV5z3SY86ypTNnguEri5xkDJaKNtNYbUE9wHM
HSzu9Css3BI8PH7SGMrqCBRw0+ozmMgWiIEnT7Tq95NsBT9yTGoJHX+f3tuMRtXt
3PBYOvi3yXqUsyhzafRxVW8LxtVu8a2G/vVWKecwnTF4PlxH6F1HOzHgrK0HGEl8
6unFdS+QQptiYMAkplxnfWnvFtmNhfuTVZJ68h7CTygiD8FEZ7W9xzuxBll+URFx
2NDGwrNLwf9793FP2bFMJ2SD1LbcxIm9v91GMK9rwR1EPnVkEbp/I0Sp+IWgat/n
9kiDqsNCUD/i+miXLxeABgb5UQdALt5whiiHWi0sYK3hZN25On+tPcynkOMV6yxO
qvaglRaqWVhNwvhKNJOQynkkL4aYsx6ziEGPbr2cazlafv1ECkyA7iBT96eMK9p4
LlexolvSasME0xISJQgetguP1XxhTrOUuf6le3cTwOc23McjqY7xLIjQ3Bz7VEpd
Lv0XzwjJ1H5RHMhZVLdYNqFerxbCtgrJRkMig3hLDI4hfEa99zvnHDrr+zcAWoa1
ee/HJWWH/TE2DAS/m2aJc2HwgudnGR36AkcKeUSDM2qsYW6wRWWslswUWF6HX/nm
r4B/mnXQ7RBVYzB0D/KeRkxvOaI2X3GYwBCLcaZB4msw1kUhxN9vrb4p4ULKca0e
RE1f/ox80xm1nbIWIbLFdTLYQRVPoZoAa+E+eSf1Cij4IccJCd3HemGfGmRLmz9/
zDcxAwdWFOrwjq2CTmE5GvNGfiWU8QLji51VJDoSavckjGuF+qC3cXdtN54Lwcng
jpn6KHFAZyFA/+oyG4rE2UEHtQNB2qQla0gEQZBrYD5Zgj6C617FMzWmr23wxP1r
fUmjYRtlLw6KP2ixwR/ur4TQKV1xEYPTWElzv9m2wnsIvRvC2K8dEkRl1S2XLwSw
nH1SPoaxymTehgiHedDbjyzaLJjSBxfQ9w8tUjGxGss+etqyzcmWw9mN/YXCZ8gd
zKI8ut11LZ/f+Ih2RQl2tdR+xSmbG4RHhJR6mMGBMDYhcvLNJEk0/5+RduVJAgiR
z1RF/x0X3DBkO3lObVVPlYV+zseXgGelAVVxP2pST2k19YkMyoyFif8DlhHTyRVe
wS0ellNMk6il4ZufmIOmRJtLhGnSXfytSxNzmGO5Jl7DI0F5GH3S3eUG+ocG6OgM
ia0KUdfqAlVTkCzbwLS1kbYdPWk2JTtkR2InrXIw80IE2v09TyU675mXStRxZs5f
ddOBEauPaVBKJnEU4jr+HC+tgO6jsWpr4iWko/p5OuSwlznzuRJkP76rFbugfeHY
Mure4M21PE4XAi/24WqOsKMai1STXdjlj+u1NCoMQhdNjfJxIQZ9ElGaOJTnZiL1
aVYy01hx8Tmnwtv+L8EXMCLbZY40i/2OqFndWeiz74DS67deDSyxmbZ8FTM/P8bf
fmepoBIVTPPdCuDQlpgjw6VPvimkOYu/rLE1gi2APcCLhxQbR88vZWAoVindmvRP
JjwvcQKWSiL7pniW+11sM7UK6/lioOrV4NPVqsBUXaWe70NKwsNjKzpvw8kUL2AK
FPLPMCQ6LL8bOEsOPqfcPN8KSfuW4ZqYcA4tmPvKLfVqxV6JWCGSiHI3JPTfbaf7
DgCMY1Rs8P/woZXBX4lk87eYZVG19rung7pRLANUtY3HX1X+1J1bhuNQgr9f9lx0
CbjFtejC7ujJSI5pRZvrKybTQI8KW7zEBriU4l9G6hkBQ9yeB5G9/YbbrIOA2UA4
vsCQqsbAq8EHPJHoE2PmEFUw/RL6Ce2VlrGFCzgHpRPtjecf2PVHA9rolcdD6pU3
6pCWWv/otF+r9s7h7FjAR/d5vdd2Lzcp9LgEwbuXRFCOsFrGkNmtYbBPil/FGvWg
kcY0+pHH/MDCw3Kl3FSPq4kzyf6J2d+YQevQ2t/lB65MMtW/wBLV1tkB3gNuwL7g
6TFyGjVRtjJ5dU6ubCYGH1zMhoPbILv6K5U5C+LQSmKJvsR46Cs6yp7MKtjE18rS
FrxWRq9NZMiI3OWIeyzib0owqf7v47kSiLHh2uPvob3yweQnyYLXt0DM7hhqni6Y
uGQtwALqiBAReWM2eNfbqtoseDcffdm+zv5jMM/b6l7xE+dOTKZUfYCTesvqI057
kmQFxQIADvIhlKzD6krzUyxokf27DyLv16ZA5eBi5Uff3y2ns0xFWYr6VlRP6hAD
nbh1ijAbf13fsItWCWOpaW7De52o+7qu9fO4Xsx27hpC6/+P5N5qZ26wXNwNkenB
FJjxOaPl+CpdjQnuutiK9vn51DBY9xCJhw9hqSnLS1OJEIL28LpBpIcOfH0UlqNm
rSYrQgfILrVQcbx76481sC+RNjXPHP0tUy7aqtyBFmfkh8qGxTmsGKhvxvfUti97
iM8ITm7c2hxEvp2JncB8IGvUZaYDu5Ud36YTM6ev0qijVhcYEqoF0nTQk42vLlvX
u8S33ldJg2EvDzU/rSovPjI/n2/DD7mGNAsThzWLbPj0Iq2s/gOTOOjAdb9DgQ1m
+aNSxVyoGNN9olmHHV0U5YR/Xy11jN3JiiNd+UlpmF86QM2ScX5X99vy6IONyEqr
jsygu++s7macphzjrCJ793dD2xwcME9d7BnNBGU7V3PieXMIAzLiCdpQHxd77LIi
hzrq3ex0pmSAnTnzkayujzvhqnxNZeMs7CSlt99RaPyzfRd3I42uowDdYantlgAL
tbmLkHBicVWhQrlAKRwSQxRRMLBpfHBJSO7ePpGR7owagP+zV9m6ydJmMZ/vv6X0
dZ7XCVUAg2eetbPqpYzT3LT2QeIvz6a74W+k2OPEaT4xpjQiZ5oM/rDO763J5EgM
flMx5WxzmwUwMz/Gdm5f1C5ZNoYmAxwKtgxmdFqEXP9UQEWkMJA9YnQISBWwoiHS
pPycf1MLsJw7qIO7RQnAJdGe+uH0qPtzuwcLJim+qoHUVBIi+XDtucqdVN9UxbgN
H+GmPXNBcIbgL9VrDQN4MbIVYHdBL6kTDFhI6f0pTZF2+gYTIt0cmJHRKy2f3b5L
JfEEgvplJnZtkM03SoLCFBbenUhE/8M+HpRXsvza8MIDv2sf948gTKRN46MWOPDK
K6XZ+j9DLs45XQ0Wz7eMi4FQp675uzehBZlGhOTUS90VJZolb13LI1n9n02WjE5F
09F2CJ9zPMNR9U0PpVAF9x8Fa/9XPGTwXfz7XEOAXAomy5aJ1tB4VdpccfcX46T5
wnmeAVWGaKzjtfcgO1XxK5/UalOwZCLBORyIJQPZmHp3QdVcXMldORT8LCQhvMLm
VvkW4VCPHKE8oSqUnMn3otfc/PJI2t1ed9GhgUcI9q3NO/zoBwHaDnl/s8jf8gFh
IfpVu7TadPOafETwgEiM8FI6247vSgNSGa5MwRF4bKfwbRDPYhb4BjO1aK9EAd1c
rPPqKuwBvbFqpRYadyxWqNA7VuFKUg1gNCu/rfiJVJUp6REhVL9w/ytNSWj09HzO
/3nQ09C7S0x91ec6a5/N2d7Q1aynkcxqMADFi5tGxdQhZs4rYG8+tOf9zOHZPuXe
sXK01c06l75JcmLVIMFeNstJPateoK+EOGvNjvh3HjTpQUep1RMcN361EHaZCmgc
4aDRw9V45+8XxkQs9retu6K3EG4hyJApyJAjnd93JvB4xmVPXdhG6UYE7wA4vbLr
77qnATSH+g2kiMh9bpHLlxVqgMPCuKDHt4SxubRdNEOqKsNk+kmWnTzLt52Yeikm
y0760VYHK3W3igusma8/WbX54v43K+oG7Uu8srWSU70rovyIRaWtuRF8vXUotD0r
ga1qkeCmfbls97Ky4kBWvWNfki0UhChMk3iTYHLPOJH2Rx3SFK27kZ4LkbEB2l48
uIcz3fkfSr927y104OTdeCSRwdyFuJAEdlbQFqIONMGHc4tYIR+tYK0Dxw2NaN2b
uX1YVwAOQdjb4AlMdpqH2IaX8tahQMrSRaESXZGOvUlLcs0ZcY/RsYVhbjs7sUsP
SfigMn4xXZLD1kg55MEFYZHES5M3A9YNy+98ocio7pkjoL7xMQ8bS/EbdD+IMQiV
Zii6jjtT/1Ad/pFWIrJfUNpUnH7PIHINQVp7RJlNaXSJ9kiGNj1+0i1MwB8QaYap
1yBpJv7nXkTXiFljl20lPCdxQVfIZ4NZTOOxYv6CqUSz3aDBIubV4+a44J2M0UEV
gpKUYs+ODDm7SyXqvv3DBmEPtUPqZNFl5jh095ganGlr+UwiQXK7CVR49lMrybE7
thb2DfBITr9LI7bXFW/WOeIO7pNh0M6OgecwEfHWTJVyUjVAkqD3U2s+h3lM+2t+
dzz7OVxuZ3W7anjzJuVSi442rpXH/DrrqvfE9NPMkqwOVS1TOre/T/M0MEf9ocPZ
bq4B/WuBKy7r1lKf2iD5Gtn2jQP1uWDG99vUwyIcN+KV0Y4ZOOnCD8zymOWuRxx3
cResf6gNJJkhuKHshzPuFRqRasRFO+SH1Y4mX3ohPU23Yu+7X0/q64JD/XidFD1O
o/56JkncT+bL2xh/VzOh6etH3oJ2ob3kNxDApMBnH5FKlAjppM4E02qsms7hJynj
mWjEijN40fbXNLfMcdRI2xUUNYnx3kdakSzImhsEsnM5ye9Z67t9GEufYVoo/fDq
alcIpqKnKtOWiS7cRykjDM5yrmSONDdWsReAAH9xw2IGp8VqCYSShDavd5BDLgKp
4RnVeE2zEjxhYNjKBGfCQ6NNfIuiNDBflg4yc4V6yFWQo86wGJZ6dC4LdXFmT5Hw
UfHXctodQRX2edd5X+lmWqcWUaFPmGsIDvSkMnZ8iwzOJSOW2PUlGZOcvkD6CZhT
g6/8rQAvNDSAljeAdDH8HspcCXAQ/nB/7GMlzM7yCB1tu3uvuSglaJDkrOKDGQL7
OfZnH9DxWan1PJL5SD2Fir6asJBkPefuulSSma6OcGGHX2Db4HLkfC6XaZCDHmEa
hJi7wwePSv6BRfc4YH58RXu+iZ0SG69Va2y8NismdZrOOXtPA/sM1nTbO5GdCuCD
vEwnsMe5dzTZiNKEDPaN5okQuem1h21TAdfRYxxTZ1I4U/4izIvg6wi6KUW17bD9
OWufAoAjg8bSmmViuz3ptbmut4i/SfPNCLt7KuTd60GHcNzh5pwjTyqBuqxTEFE9
LTnR8WjDoHBI+Gx7CYzZO565IUcuVHVwcgCgtG2uGKhjqyWoFBVRRxuu69ppTtcb
QG0m/M/IM8lPWPlA2UzUr88oDLl4bpcpZc+YRJwfSDsz4YG3A4N6CEfZ8+MNtfGH
QjFwQKSR2fKhlQlIMG3UstpbldthIj+V9LaAOfYSGxCOsh9pfOpSpguk3eaefZbY
h1QvDr9mG2B8c/e6YniiQmC7l+4AX5PF9S0C6JW5zdcvnUG9RUZLmRcmLItFiL05
GsHV08wf/fS9X3hLU6DH5mZj16ybXBj5aB9NPmJbCoEIydErkYvLeFtn5sj9YGys
C4N+PsyoVLFYcFtEO0fPCckWSdrG3RIGoIOVYjutb9YCjIi3DG3e/mFYhmflSjSX
NdFmwNpStFaRz1NhByRtpt40XD47Y3a1RpsxqNHNHcAPN+xhWVFGEg7B6ud8Q1i1
5RtPOBSDPcsb2Z/OaKiLp8uHwF1qryfOKE0gDV2a2bJc+3NqMqnjjQaY1PlFbZ5C
i5oZNVnJ1JRAs0ce0OOULH9aqUrxe8wgr/hTywP6fQGC8DEEe11skLin2pkewT1D
A/5DlVpkehAvkRE0NJ12NFx5cp2Kc7OevVask0G+TUUFgyA+/77whTfa4nAeeLPH
V6Y700S9s3VVN0xMRBHyv+9Ye7qFGjaD3T9f8Rg+t6I/rBuF0CXpYIwV6lc1VWfb
CdFXUFnIs0pFfENv1VX75CP9CR/kb2OZJeE/cAOG4o9weJ1syYa7mvSHl9c2tAgq
rxv1DP8amIJVeFIPImC3OpeUjVKIUxaMDdy+xlFZteN/WAK9DyAmufJg6mw0pxF5
/YkkNT/Bk1Zpxwgo8+Q4Zg2fsdZxv9SpwFgwYKxluEnLch0x4zm+vskQGXfCjBrB
402xfLjWLTpza0/P/kZOH/cAdwmT2S/L8aSTxX+Kpa9rSpzT43eAbo5ltIjWQPWJ
1505kJN1lZiYi7WBhZwmWZsOmPStl8klNqz6VUR/Xv+OgqulGyQHVd0AZthu+Jjp
8+qtjvdNNpCCoATzPDg3iK9Iqs5N4yacdvXuvstawBKEITUEIlbU7XMmBEZCgN1I
tQ1YMsVl/vXmUJTwn5Ft0svS+cRcZ5IH2R1iGkpvVpZZyFj1PaSIUKpP9sxBT6i6
D1kWtpYFbUULtN4D/GhiYmWCY2fEU+deHK4f/MuxYDxkKcd+om5VCEFw5RQnXcf7
kQw6wTMgyjFpEMbFcBtSt2c0XplhMIJBotFmNOIUVe5hc2l178kGuEZDYgY/TWaJ
r7/Hygtrf/vOU0VwpG0wN1Mx7ulesbb3Ze8M6AcK1uJf2hDps6t1Fbh9nRm1xKf0
DqUYYB61gJ2AAXrpPnugO+2zYoKqdVX+u5+KzlKxExaamX8hu2dll1SU6kxPlNXc
F5fD508AskiQ8+H0KtI0IhZMia8ayDvWavA6nnqABZocB6EEbzEKtQ+pcNEE3Lk5
9PtD0AJqiXmC1eQK0WTiaOEPJYUWJbhvne/BzLT3/PVJYk1I/pmM5rzx8lTNcLnw
dsLCRVHPoCy3jHqpa4sYZnRyT+yAf9C4ZWQTqCrTo6FQWjzbUiq234a8AaZ5i3m4
/CrmR/S5APa339vw4ruF58i2ZDr6vvuv4xoxeoYNP0H40u9jifsBAAANKwH+wKqK
HtCxVdVn2MwL6tjcb7qzkSIFiHCcFK0QT2ZsbxHyrwijHjZak5saUBIqtiqcmgY5
A9Zf/qOkMsujiAe3+BFGhVZ7VPmvP86YgxyWKsM5Xy4ZgBmKeFgwhKxhOc9vSHNH
5xbMliKsYbUYmS1LbEcyNfhi+lGgKrtW9ant6YrFZ8Amm+ujPi1eSCo5uvNEq+OC
i5YEPeplNRzdx3VxjAYXJyDIAygFjkLTo23n65N7fodc4ssTlNrhuGbC2kRjGBLE
MjtUC6jAwNd45MTUlTRU2UZXOXCVPoAm3f4M0gTgKa5kGRtBjLnbl4LeKCuP34ia
0ktmHfK7bW24T8QCuB7Mp8YPQWIiS01EgkvMQ8gOGQjgFfo87FPD1vlV4c299CNr
3OEUsuoTudj1ZW0HD+GL9sYu18OnhWHNDtJ9T41b3x9n+FGyz6thWDFKvodJ1XWT
WppV0UskQDgVZCE3VDW5f+pb42QQitQU2VmoJRfFeCNbZMNtj117lTuq7TnWeJpy
f691ridozKgCq0XerZKBmDUJWNpEZDyZCgCpXBI0a6l3mnij94koPacnDwoVjzkW
T7wkCFo/mfESPBjzJXtZLmoKuwC3eoctthzkhvaPx4AJuH4Pzto+nbvFf+NHZRgq
YrDa8OFPFOJ00Vo3WmEs040iyQtP1o7pnrrFXefLzKHujzVgFt+0JYXRv6Eb1rB2
MWxz1GVfSaTL6/Wt8PTy+RpLQ4dlsf1X8cgQAD0DMzJjoLm9cR7Xp/U/j8+L17pG
NJQzGGdpS7XW7iCIMue3qOa0SW6yCkt9uB0Gz5T5bHIGTE4AnNOD/kA9PT2/7GK0
F7JZlKI2MFrVFqWyuOJafacApZxhpISLK8rE7DHwpcEIUn6ZjM1lp457q7vzZntm
qOuyM9Un+twSq4sjYragiZ2wzMPmiCWgtVsQ7GYIX7pw/l/Kqupr17qVjN/6foJC
ouOQ3QmJzqLV7lYWpRd4BaakG489KqV1k6DJp11siPDBdf7nNvux7RO5ErpDoa4b
xjxzlqSj+WQF/UTAZZxm9mFN7DA1OQBAHMpWBeOSquvjDiq3Obcmc4jo+g1oWwPa
HuF1zZa8xcYS2CDTfvMnVGBEhvlXslcitl5Lpj7bl57u0XATHz2AK7jhvWWUJnTY
WIXtVvhEVADcQQ9KKojQEhGM4qSKgsOyFv5vAJYUkCboSbgFphRmrvGyO+NsH3ff
AbBbEntUJ4rxPTZoKQDG/Bm17h7TU8h3y2lkaVmJYF/r/rA/DDhHLSrklLUeK4KA
muf+QBTC0qGpeSq7aUIL6Y7dD29p09NQPp5oEe1ssv8akmxQVkbgHrjPdTipEb6B
ERqL48WryTMB3h5+yvcaueGZcbdspciIaV05NiZ5nAqz35b7qdITOBRFaVKBXPQb
8VWYv5Xj0Djc8UjdBzzbDBXTGc3yVR9xw23WR9rlLAH+GjNtfIxEns9c6oZx32uF
UCr1QCZT34xItBMa4bsoL54R6rMLAl0+JVl+x9TiShJRJJhgZoHko4lCw5Mtporp
quWSjOmO1HEOp6A6DfWk6n9UtNqz0siOc7d3ZK6+1FW0iJ3RPnjpglufCciOvNiw
bP+3yH67AQglXeqw6Kadl5XEzkRbLPFzFo11MLDUsXQLNVqYCkuobzwN+SMKalEv
k/b94vAXJyVQshsA7FfLQaCA8M4ZIvaKGrCJk8AWSYuW9ckdNHZUMA2wMMGFreMA
usZPXI5Mlx9T1vOnpicXASUk8NP6MvlEMni347oV1z75jOVyKrhViUgt4/x6PTNF
QoSuJyl177bzou/1riV2lj4aU2QUIBxww0lq7NOjGnoPaTZYuBRX2yIjxPgEnLet
K9zrN1g0P72DRymFaeuz5oFoe2JtGAYt3DJBoDxXbzW5b1g5hA2G4fhXMLnsjnxE
bNxP4529bcJu1FXhdCPEdVw8suLgkaR3STYMjfDyjYSsQmbsWIUJZsQsR55R9HH2
YFPmDA0WOgjrMkAv7JoUhb1n0DkNiaWuR4xYPvYoQHPO0FLucLLJSBjK0elIn6h2
+d4rO3kKP2nUB7RYvENLx1G/zaPxhsH4TD11Z8nVvpvvliX+O/DWPYIAbxeEzeLa
mhTmnYtqjbpAGdVgmAqP1QLhuqzSlp5zL8nnWx+85RiamU7z1sSrVkgj1qGc4DpL
OvH305KnrZy7heHaPFRxXJwXW/j5ZiFPzOIyBFEfRdwJzSjdrjoBazPWGA7t6USs
lNd5LenRSI+DLaIYojjawvzP9qET9+mThAS0KYYi7syqmOpye7I+Hkc+AsHoAzyL
ycdOfJOGFUzMLBBf2CjatNr1bGqJuDUSBuJuAL5Se5ba3eQF6fq4SZbvx4e0vNRo
YA9FWWPSMJxs12iLRIoEnoMc0mcHIuEQhe+ES2tunM/zDEQ+8bcD2jGuyjCLA7v3
8ATDEBSuQ2reBHCHYjlpxCKPrnSscx0G02DiIcG8SsLNQVSV1HESzmWu5rNl/+oA
4ADmaFxw2EAUHr6CFZRNnHzOVPPlHn7rcpNhq5zg6YldhZsh9gl0hOnOMwphtksO
RMzPdqJzWYkI7EcmKxqAMWi0DpLrftBPfTBbF3Al9wUnQHSRAXKuY0ryKkGIwVfU
z1zSuDzTR6/o5fGQFtguzXPXGalMB5wp7E5cs/NoM5h1xtZFmeveYWbzBh9L2Fq/
zdDUYNiIjUABs21hv/X975Pu8IlOj/wg6j4n2jNI5SfDagpQFgNKcON2YdZNuKS3
+vcUIfWZMO5Aa2bdRgRClKs+IU63SD9qSUIeybGxWseotRlXp2woh63wdVaS4CnH
Omh0PHykt4m/NqQ0sd+QRRuhwMJRKQ1mb0O2JsrKeaBWyjPwowhYOxwUrC+gK2/k
NTvKBfK+ZLdZZzwYzVDRepR8TD0BZG1lIzfegjx/Gyclk3P6V4caR4RPNhrdGRyC
7JSOHIeD2/qJ8492OdKd9x1BtNtd2TRFzn08ptEc8RKvBmCvdWMs0wE+NnrHqgfZ
pfTePr/xTmvYZPvwGL+yNP9bx7A/iV8GhePEyL8hFOZjRHKPYT0ZpqPkPLc7hoO8
xdMLdRaN1CHMTh9/Kni3WzAmpc9I5XjqaIoBdfUcQzoZQrahh2Mn6L7du1igiOlq
eaKyrNFuNxQiBL1xjujLS6JBJLueVWcltLY9WTjM7F2UHury0mJemC/BfJTb+8aI
yymG7aFiA1ER8Gwsupgu5jmF10A7b+etD5nnpx5Ql/Ma3AnzLo1HtbRA5QqdnZO5
WjeqiK7GhFBcVkrWAk//yGtLeGhDvapCW0m9Qwc/KxWlmTt5cHARYo797gmu3bWs
8qg6x/QZ59wZqeCCs/OUM6GlK+6OfTMYkaDtnbzRDTsVoV3FlHLsqgqQJOK+TVHU
QocBmNJkUc3ZoCWaHPl5aO0yDp4SeU4JVc/+VvijZVV35Cmile0Kte8xMeL0SNej
fPvVyDgENSVGdEv95ALv6Bl3phmzsqeYxhKlrGuLbhaMUifuF+WMVGLMeMqVv0QA
vjnE2lXBgSNy60i86OsOzSQM0rq9FcdSLsR3TgKBC+NwWpcvDz6OzN04PPuDLWHG
iBXYRxforxbcbYXI0xx9d7Ga949X1NElZywIoY7TU7VwakAn8hhucg+QXBTCLJSW
Z0a9jw5yyY/3AZrxIe8MyRCPQIeiWbhnZ4htli07fZPf9CayoTfjT2kPiEXM3fX3
QUW7WWA8OcagJh4k/HyxFtjGr1Qx5Sl4673MuyJGsPzDI8Mr+wqAwJOf8Dje6uBc
COB7tqvalCPExvKKDh5IJEWVnIeXf/kjvjh9+bvSPz4+qmacdzGG8jvzZKrPVggL
lhwFDa8SY0DxcuQndWqn9DNVsotPNPIm3D14YFC0dhj76OciGbkMtZhztKXl6MzN
PvsTnAPV6tH+baFgsd6zSxfOjmC4RFad9YwxEtaOgL8rXlZWKZ03nUOHWBApLtUh
04MG5TcCSdcqu7Y1HTRjs6bEhlOjiixOYFrMLYEOsuBSustQ04+My3rvjIISCmRn
qIJWUkmQKgFv2SPl+X7cBYfMDFo5pk/0zucuEv63sNtX5uBTS41VsSnbPga6Khms
2OxLFSVmoy0Vrut0JXGUnRSfDowi+B2o4K0OYE6u1zNs6Ug9G+o9WDLO8U3WbFX3
oltjgZuMWXLzCc/d628JkknFZBRkpWK6LE7J/pfgiO+YWCqOzs3Mq3A/FFLksCOZ
Ky/GoYpTyLGAPSvuvCYKOl0uLO38vvfksha1H5MhfJmM6eHUaVrAOOoQq93PRQUI
3QOe8/rqLQwZJDpGRvtLkSMa4QjAiLO1tKtGqbkCtEW5tjI9h40S17jlo6v2wmxG
rjW4FD1Q0SfS6AgypZLtkl5WK1fvzhR+1644lgiudA2ergeYa8YEnp4omzr2XEQs
R4Z/Mta+F6pRN/b5N0/RWdfslMjYBIrGnsUDqRBlTJXUMIs7DglzYSB3rM4zgj6V
wA5cTK4q8Q+Qu2M6kQ8Vt5h8mLHoDIOc5AXjJxmMENKl4G6SxfGBcY4CJF9B/2Zk
1N/+CriV1TMRjdGrU7XQsq9bafIhWIzLw6TYrPfIlG+J1EqC3H8bDIbZH8Tlb23P
UWak3AC0HbMlg0lNFPMXh6yaUYfKSkLgK7MxZUS38m63UR2ectMbs8J8hsnBC3R/
s+wrcatyOiFwVcysZgO1jov2sK6bwsndmdhM/ZotAKhhvcOeOBogtR3jAYsV0i3L
Mmq4zeWZhp7ZkVbSFZL6cVu+IquQy2ON9ia76wGXetg71CCCfkiCb1Uax1jHAchV
hfvr+opan8UyfdYIWmq+gf/CsGjgD/LsIaV/Hfd9am6fXDRVcQhVHropUQWiO1Ch
iooq53RPXWMf/2nijNv0jqkhIMO/NuVRnPf3gOgGgVyIHnJ90v5opdRfRtT7aIWH
rLWt2clP7swOHjDnrA8yLn1zyh1KCMFz+NnvIy99OQFG2imfylivSm5p02MEUmAk
6S+1sL2N1ocZ3WpYdIqDAuxL3ZtEF9hfxjeNX61btgc3Kx0zHdeZYnvZuYDFg0Lv
AfvGMzUapWqBFQdwZySRiziWogV9PrWGmUP2IxQtWHkd548ApX1zaCkt/YOfhTYc
6dBF+QWYHcAHFW7ADxV3mIMBh+GDmjspbF/JZ8keRW5VxISDCYFklTj3U3j7FtGY
qQN/rzLtwBnK6e6EWqL7bZFgsNdYE1NiFEKUOqIk6+GH+GFvX6PY9RhyNNbBJB+N
V4WOwNb8Av78AwVrV1i55mGKPIFg0n04xsoqvi8bIe5an5ggo+8y7dfo5FcT2Cif
zNMdadG03gQUzQtSD2dTwhqMlM9a+SzxMX7XIbdhlo+LTzrO34WFMFlpWeUrXLMt
KibXszT2saLQZ/lhciElNOQtN5P/+XlVdRjH5fSi2+n2zi5c3lGRj5S90+KKRS21
5BZ2TrhgpXK8GFVO2IvBYOk/CrFwbCEMyB8h+bWXmjiMHn9YSye6DeN/NYIfWWvM
YaGXTkpogcd7fHsir6vCMtNjXG6/LMxAKGr5h9iyUSWGGQBS9urMyHY9nhdMaidg
F2uTErwtkV1fcHGG16ns9gfJsJz1r1EgP2c0/OsZL2YS4WL5FDgrBuA06X47PVEg
VOcgxYJx+5qr5KOuSWDZCkLM+2g8oFZx2rGC32egX6aJ2rKfCqt5M0kNauNo/R8c
yDwX2bEHOv0HxkCcRCJAy7TqGUfMO4a+/PiTxcvWUFJMdE5DF3suUpc+2bVpYKST
0kIXcRaSoqaseFkIks3cDoeWvu0uWLPAhgmHOZPxgcvLxoRZ/ausHrYts9SxYf2i
m/UDWwtuPGW5yMiQourUO8QNWSjF27CCypCdRxkvWrbitTiLLs6g0rDSLOHD2u7Y
3UaSRizJZ42iXp3TE//xKIUpP5YxWpIO7XxfQqX4CgXwRVEgXKkV7GzFv+/3PSAi
/y48I/ubcf1W+oacJINURatC+uNj6Z1Zx1HZI5UQtndynHUpukK9nDXdfcCjfxVW
TkTxs943RflehPi6qHXkwrbQff8LqWjHpjQcm2yOaj2HMeRN6t/Zp3Sb9JKXL9X4
EmmiewnB2IP7wzqHYotRiInRy7oikIEKqs4AnQxeqTMgpj++mjig1MZkefqUkwAf
lrvS6PO6dWrUtQolaWDRr8GNuXlWktR8X5F4j715NemGLqinn3LiVb5A4nmYb1zQ
jV0v5OkpGExBETBeR0k6S+nIWf9dit4rATAnZKT04aXmTCYzhYsR7ygq6jpwBHDz
hNMJ1RqMB9i2nzCH/UzcNx+dlJqfC53rs4VtcIJOHB4bFfcH8YHGvD4XulQhytLk
1AuHZY7JMexqCVUAV9Ml6XkhuGjdPtMCoyikOfDh8YLm+nAlSHnkePC84Kfgihwc
HIxNmALaXU0yuN1R7u7XAdkNZ50WET0P9gvprvvnk+OLeZ40W7r9EB2hP6gopKm3
j8dEd/ltLmTVS2UMO3dGRQhjmiOpYktaLz+mPlXAfwymmQmLt9JR11IwmJW06c+i
TSeUTtRRahMrUrgjFiMYc6yB0CaVJ3oBynfVaJB8mm34jN0Vs2gsRuwXqhN3WL9D
Jqn2TnYSSvBcpqrfbivd0PsnmDUOYCA9mPYOjuTnqzTUTA7S7+em+y+83WIQp5CU
Akp+wNzvrKa8t5B0TGxF5D+oTiEnE9eKGicTaTjh+3403Z23qq5g+ZNwFCtzolGE
nV8zBgz3aQ3idqpz/sdgC7dt0sJMm1kNsGDZj4qcwoc/pBf4ivxT8eO0t714lLy1
FUVefasKuaGivLLcITpJmnptVZTMHYRphpBD1kAlndNrHSuICc6Z2Jz8K1lrukvP
0lwpBxtCUuSCiqx+CtjMyd8K0iGVw1SWhcBklfee5On6c3j4IFAiDEOlwFQAeICZ
Qw3kx68r2c2c5NDU3wPjvsP3B8Ic9FqKucNXB36pkMHIoRe/OoiPqZ/5bF1M96UG
22m+wUPvyKCOQXb6hucVQ46AV0piAkBjVLmMjq0xICuXvaRh5SqzzefaIGv/JW3q
z0S/YSIrtlA7zdwJI6JockOWzwehoeJWKhKK9auW/xTwsCAhPIUH7oar3Lygpb94
Bu2r+asTE112TbXhqziKEXbsCKGtqxPAOFOrsE4i3KV3mZFYYHdFR7YZ5fGY6cMb
oWpNi42shRG/caYUKyBFYJ4WF5ROj2iSWCWraWq77x75pXCPhk6zEzGJEmXDykHW
5RDd8Kp/E8WyETVd9ZAlIeuAAJxLSzUwxOx95e+csa/Hd0pwgJRs21pETTtyLp5f
nOSMD0QgQkTYiDg884q4ImSgRBHd1X2jJU7UWMQiWyndmV27DrJPU3ybrorUJm+n
xDCBIjYkPVKnnNvO+UwOk90Cu15TVBLYCubuFtevWXEKUysUvdQal98hsmEJ9mW0
NnStGOXaUECXm7Z0jpZsGgCeZUmlf38LlJatWgSblA1y7k2bevqkeE5x7ki3BCPc
eGDrespPBR3tl09HB21VvkFNlv1TnLIdY0TEGzZPJdR+/DI+mRlfGxNvA+Y7nSJ5
McH1zua3RKjlqTkg3GWZFaGmiD20rl+yrWb6bjTJEfYIKuEpZxDDm+UElWOElwFj
iHZHtFLvPdHdzrfHu7GADvbXSUEEDhN9QRuVVt/mVFKOOoQEE1gdXgn1vbak6ueM
COQZnpEF79q1UsJUo2fe4xHqDAjHU+xHeQzbxY4iah+ouXYC0qQRbHkO9UQcSHFU
UIeIvdMBRSjChhC7scQH7M9RT18XmecVorSVQ2ERq1cDkEvjF+8GN4BgNq19I3lx
GZdLz4K+YgSE1Piy+ZvQAvu0iZRs8mEJfi0SDADs/DGIzWw7hQIJ9ww7PH2XzGFN
Iskbc5eEFHhzJoCGXaAdKG9uwycVnuKbZtvGCeqK4aINbyLtf7XS+YuVV2BBePXu
x0VpPOLlIQYRAKBR7BDc0SXER7gS4Q/3mGSxJPNfoV1aUxsYlAlZq5KtHDragrqs
skRurQCRX9GIl7JjqOzD8JsC7RAsOBmMpd+HB0UsDZudeD4J1mX3AyLElST9jaG1
GdulwvD+7z9wAtvQSVvlTORe1HtBOnl6S455dxQatMOO7cC7Ph2mGSHK5WOIXy5T
vqN/bW34mdKsFf4E+5DuKpt0jh2pQcN9ZnOvSxwxX1qFY1y/xvmmadbkV2QpX87p
oVhrFA6AE/7Wyi0ATuYsxb5W1vpPb9F8kR8C2v54Jjcu9tS1yAwc5SH/8R+K1Our
XEhc7j7fshN18c27LeBe1wq2ZDyuaCRxFtrm/tetX+vXcYlw7+cWsy4wcXOsiJmJ
MYTHKfnVHVTCnseTI4i26KteyF/GVzvdjuTPF8XaRPcrvm0QH7EIfw7YsL9ZRnxg
cyoOLW+192Yr5MzrthoHiIjn0p7gCwyJsKIqRuYa3QJBezsSnpvr8mQlRX4d5QHE
Eo/w2qmmGVzgsGBEF6UoaJSTmvR1FmTeIPY8J+DEUm1qYj5tUU5SO8z1yskack4b
eZHr156suyBaESSWcvNFyG2ral2+05BjNvgF+HMba6Eu1jLcqLpsjOzQtDx3Uc40
AeEXi8jmHPy1HPHnActusWqjxdg+hif8Qef0KYsgoPpVK9zm0lTvrJnAqFKjBMVZ
08RiaLiHhEc1Hb13RMbvlo+DwyILB+YdACI4XosD51J18Y1nY8yYFCgiysOYN7It
lmdefLd2HkreL1B2r1anOm8AfOOLxi3suCdJn6uAJOYya6eCLHfNIEL25K9kE52Q
Ei2CdvB9tgzcmZLbQ8SwEQSB0trTn+IBzItK2Apkten7BQKen2O3wMGL6/G8TlfC
VhRQxCcc14bD75rh7Cm+oYaB/HoWQfUFmCD1/vX/5lkMpFp1EX4ni3CuFaMYyRZW
vLgGa/XP35gBwaZOPokyvOsul6lH4UYAnmZaFVgs6IcGB3Opqzem01Yf8YCZKhD4
/KRZaJvP0BxposUCzqitRaVtbKjpaMzscxC3fcJbwNni8+U6Dr3KQ8LzrlHF/WJS
IJ4K9QPNlagNGy3R9G2D2NVSi1h2dibuulUVLsZDPPx2iQKKAQYGsuIv98qQz/Rc
52StDJtP1L/NU+U8VyYdVpyh/iBpZcjEELv3KL8tbHsZl4Pjt33r75M3s+OVlBvg
FbvGB74Xww0l6+fiMx4CTKarUDY9XTFFTVMyEFawbxKyujOcRiZxPXWyxiiTDZ02
3W0AuUbXBrY60CYQGOAIE99WQ1AVtHukLn5Kgl94m10tTk6PdYynOwMSEB1ma0Yr
Lt/Yw73YkNFz5OvQ8IFzEttUAyPBua477VosveLI+p276M1uujw/+7QFnv6rgUsN
flrwrDeXOLJFR/7daGWtbMV4JNelBOWFLY3UmCOZptvBH2mIIIhfJ90pg7o6kqyI
18BXWlp46UwWpAMmm0IEc16SZg7lqlgvJEM4pN568xB7f2dKbDjKUweufONREQK0
jwf3tIYGoMLcwpcOgMWPOX6S/aCg/5ckVQ4kh1GQgyAjrIkN2k+HPipUbDt+LgPV
xLRBBFmmK4m9Xmfkxmrty8IhtN3NeqpNoyGflYpiVJ6ejT50kUu5mHjwzvuXRoOz
bMvmSmzondGXGfp9ap0YmRtu+0BXIc+o+jf57wh+vtltOcpvBAxwJS1W6wMJ9MYY
/oBf5G36Vpd2ZcepczGD+F0i+yXPXzuDTHYJY1I9YEXBG/iC8pK1nl+5K8CKzkPZ
v1ynd92eXsq2NgXxN168v3mhfuTieXSIlA3u2jSIWzCY6uAtjRiQTO8tYDCvno3u
3QV+U6jeQbHHaYKTK+9dGreu7ybUKk8m17aIn2v9wPigT6dUKLkkB6rBGuNglUhQ
gI95cjVVxBJvFNhlkqNUNFvc3hlhceBdD3YXESXF3PKjxwTG3pgcDWzfRIBq87rx
GaQAxADWajHGwr6WkzDyOVDBaXjrwUDRiluri2vAWZJMjPC+sZ0x5GufsFTl/5ZE
1Yas4i6zZbR9sdAQpyidvovMZTxXH+/tKDIpYWNA5pR2eDUsdsiobADojxU7A1Mt
PFkliAufBsUvt/KuGykppVRQph4wCDBMs/pbSnWZkpl0lku5PzdJ0sNLQ7FiHGmF
ij5roP2UA4tFSv8mGRZyZZeFK5CUbocOMiQ0YTcWFFd3aRvVc/2xo3T/6cwNMFew
rtJS3DznU8pp9FJrmUd0bU0zFbUlYYShuMe1P5FxcacAqssohMzITX6+aCLG1AYF
nrf1e7snqRIt2/BAGHhQD7IG+EDj2/HqCV62IlEUjhyzkRnutlwL1861VBQ+m2CA
N/90wYRR5TB40Ylha2KplEBJzNhXsBologQH2Nl2//9HrVn2u7TanSOWTbmZp0tz
XBFL2LLhadwmxisAlYCaV3/7FxhAo6lArMJw6bhvEXZOTfp7iOquq4pGVYJc5cvI
sTg/IzmciO/wM7yJwBTGvFLRvR/di4is57eDM8RPQERz1I7XdcGcwm1gYZgt2MLx
sjYluBDS77IANswjleNOwSxAGj2j9pVt0OriMQ0lSg4/RzH7rtQgblw70TPTUmB1
EmBAwUTG4PtegcZVAgGZRrNLH6gWLldGpitXL4UufEsQ+/eAiuZbZM2NjOJEFa5u
8wVUXdqfVpD0TV911smx6B3bZkso0xQz4QETS6rc4qIeRjY88YvFR4Ip5ff2Qorg
Q9WhZv4wuekP28fZ8bbvPtv/rI013HphrmCaNYceX4Q8kvQs3qQs4QtpxBJLTHcl
O/ZtMtYuvus6VSq0O0vyyVrjiRvOski34yDhdcBwzoMSztcI3u4/kIU4V/HzCA0j
iQ0s6jatIAKfsmDdLW3Ao9p1Bji9+3H/lOG62T21nstwu0k729y9cSdaxDdh6tJK
rn2SehGKJPfSwquaB26Y131I8gpT7wXbwISZCIpcePWtuHGj1dkfuUQmhq6fv1Yf
tvicK88YsEoUDcUVA5RNkF9jxOtKwQ608uKg2r+h+onbTCLO8JZrvLtgw6egTNCC
xKxkrLoFT6lPUy3/uaEIVdsV9FAtPF42yL/DlpZLIcFcxAg8q4efKBLv+Ig3U638
YevhlV1C9juD4MSwgYh8XQ35fTvHz+aD/bjDVo3F8jkr5NvX3yHtWzubStZo3oql
m3Ys2ck5Jm1mGBR7tn2tNsgeJRv+FFEixiBdkiEAmidLSK2PU4GULex/p90mij5f
63FEqfRM0f3ir0gHdTgzJtUfSRzz11yWDJ+mjTuwf2O6P4/qdCVWvnt+V2I79yGZ
h/HmG+RTB3PUMnD9tPLT6/TO2XTkB52QuskV7/lWW7sTzfAgTgtC1kenHinJlW+H
oi64pjDKvumvaodetlUKkzl3z0u1Y6kJvervEbuRHSxoZ19dFQVKFgc7MqYTRkM0
8h3dNv7QIEdCycMSVbeoRMqxp1cunMRghkya539aZ1/OuRpfALGeiNtQAMYsWrsy
AM3UOwCOMIUWucetgUz5NQeDPjtIwkzJuOA2bCrPW9IB9Try6KxrNjO5KaNDaiKv
vewD71rfsaRFnJ2MLqy/wq0Id7tVM8lcdcGNVOqWs/2mV35akdTq/9ToYRWJcZpm
rUVmf6qFLzd7gcNs9yE0Izbbq+zTqPnAYI1r48qZOQy8JZCqa10rOLgUvPLOQjjq
Wv86qoOKGhLPVaLOil8eqEkzXkpllW8gCSs1/aA3D6GfQ5hZHIYa+PwxJc++FiIJ
ICq/GhQRa21A5mj8Y8uyG7s0+5kjbjaF376FwLHeGDxpsGuVehUdb1SQecLIVP2P
YMqz5uU8xk7Ll9F7KhsehDbwTco1wLAyWoOF2c6VVorqiQA/xrtb06emGO1tluBz
FkXHIQdLVkC5k9OtEmYcoM/BEAQNWmNDMWeo6B0aRUBfrPBIzBQc/tdEEfJ9vc+J
mmBXO9ysWQAT3E9bvxhdV+S87TxaFU5hQsxz68ejtPNL6W3pmjJ/VTIGPOugq7P3
t+ztIf/9tciq58A7NkHyYSYCz9KEgrZH6NVb/fGh9uubZXwcxM9Bpv0FLMmQV1Nq
2y6Uk4se0mIwNkLLKY9uzNHBsjfS0ZloQZmkEO/ncDnkISjZmLo/tsqmE8ttDSJL
do5oQ1Tavxv2bfjDv6ofNsRkngXvGF4glPD+4HkXlb7YhMawPB83kCce8lCz7r/m
c52VWWw+Vs9YMn/GCt49ZGS+HJ1+A7oikWN4Oo2V05tZpF/0S1GDdzGn+NxyX+zi
QBgxWZx4UnraozodbVL47P3s2CFkuxgWnlwBDHyKTUuMPdzFzNzXGz3Pek/vQK5n
QoOzuEno+0kVH/aucvjW5PGuOpumVwoYuK83gWu/FgUV7vzk2NyLLmyC3m+QKtq9
RYi0yum3OG8F2VQcGWA9/G7/fmMvhhs2gwkpT0zOodqirfns6A+AH6+kLRv+cGHg
fFmNO7ApxXA7VTMhost7+uhrD0tUtK44WKrfjuo+B3qmJSAFqQ/wppUV9K45J1HE
mHg56ZzDewr6+YHrf44nkFGg3CWsAKJ2skiI6dJExQr36EKbN+3ZoeMWg4+YmCzx
zmnLi3WqQHVqTsyfmObQNhaRlCpLp2K861jd17OmgQT/q7DErAEZQW1B5BqX3BiF
STVnhkhuBEJqIoyLhCULmHfz6o2tS63KpnWjQf4nx7ksFGJHP9flLwq2732tNCk9
xHwhmD/WVQ0ZaE5+4jRvhxn5fcI4rDTxmv30Tnemq+7/skGO18GOw9f1ZWzXZCPk
ae3Tu7hgKV7E2rOdK2b0dFqRfba4BUs3JK0gtdF6hqBFuxJn5ZXSTsRG2l2/j1fu
Chq3jFkWYUWD/EoRyFwvyk8aEHWT/tE/Arg3+Ab3WTkP5/qt+pLowsirTUa0lZVv
V73EzL8YM3c13AfrO4Pm9aAxD2t31QrYQ1UXE2PRtCZk3HzHMT54tDAYK1PPn4YW
uaimbmhTa8R1Zkq2Xrwf1w++MQfPCozWWydqto3ONePLFKGqwjvoNQrl1jCmGr0g
R6wo7LpWOycMu5KcBRH2soVdQ63ftrV0xQzRnZHTYDPsZUIIQxbTVqxkg1W0uo/s
ijdcchIz23vpj9o4Mckks19enZGgHZPHU+ip0WpTTLRRU11DwOH6m1vPgpHg5KWi
Td9Hm1vzPSJZ9gPqTvfWy5dQqZyl78+Fh+324x2HhFuRV+nRLZKVM0QFReRTliLG
OIuzDNqnivGWq6nWt3pRF5bT1ZrxH6H1R01G09HVJMXMXvBO01uAcr0bWab/RTmC
SsqQFX4b9XZGoq9OG3mQh9+OtSM958or1CqxmXqqoy+GkRlg+E8vJhARkLvyqw18
K6Z0S8WdudrXbXFOd374/RHF+TlzpPW/Hadg8yA/QvSr9JQ4B6HlDXwQsKNRopQQ
eX1jY5aTU2HL7UxAd/ineA5K/GMG4MbPgkkZRpbQfQNBS3PLSB3Qhejx2bWOTfDU
PulrWzhDDIPKVCOBI6DcfPtWQbkwHgFXFGmVaF6WLkvauij5ao3PC22atZZU3ffq
Imkd8U9NnM1qo8HOFEXHeZzDikPD84tHrnkFbrYrqyNClDo2VJKzlUEPhyCN+1Ef
lt1Qj7oQBFoePffffbkQaZdeapWYp4vNQJma2+DQuwbpTOvUtsySAKnPqWrjCVOX
dyRy43l42kuBFmznFMt2vJSnM2cGHtwuuzMbOpfQJ/VJDUtbPDUV0xPKm+ZKMzRW
7bxgEloF1nvRY04C9GJoWfZPMBrSTeqYv2hvMKGvICiK3gbV1hf+Q2j3rsCACEb/
6MoJFd0/CyynjW2CGoU+jpCfCDIuXqZBfgAzBK56gd/uXU0Tw+JjkamZ79kSgDrH
F+vSfKUqOYMEZeSVcg9qTI+vzsPuAPAG7ZiLZSab7xpJc1KgAKW3ta3fOVpIStLL
CHSUQq90OdRQanAZ/SNFE8B6B4zB2+OOQKsSoPzRrarLAfb8TVYXhT8hBG6fCfir
Yi18ew1BJ7v46NHsDpyLB4ORinypRSZ9m0twIt8XPogjLnFh860/X7C1UONwdr1h
BHPVpbTsN6WVoZ/YqTp8MEN8DokGdv4r+aM1zl2c2hHQQi9RZmEJoqv5B+jA1ofp
fo0BA9qs3INOZ3y9g/z2kE0m+PNi1nyx6N7X2Ej1PiEpj4Jd7e6YW+9kxRmenWGk
vU5Xl6ARRk+wSwokCccrYmb6iT6ubxoJkdEjsLb8UnsQwBf9GQAvaA3l4+qqYowF
RoC7SQ9wtxlWd53K570t8KF2TciNzZ1jdSpLBd/HlzzqdkQhtOapezxKwcYpTAb6
SVGkLTwEQArZ/5fJI9Tknr1m/iGy4BrtEk+e5XvAd991HUjgzF3cmJSxm5TWwi0w
GMoZqewfKycIihOGF1oMzxQXKryAZ0ffvhmSUlXTOrrYDs4GAxfpSRq1LwAVLZA9
cu2riimkGxEdfNM2CixKF3+Wwea0/gQHOuZYweQFM07nHOBv5lfyuNfe5II6kUz1
UfFX3aSXm6CmEvwPkUNLHvEPUOu89tTJzUEEHV4chRODRgBDr678gi/79whl/UWv
ej6hNeudCcVVVf6ehbXhfQe5uiqoRJKyONLCSsFANPZsAcfzttNQ50Ml8EIlbI/s
I4nd7ILlQzTM+fs26om26Rsgv1JvBCX9EjMZ/ZP0F8hZ2SlHG2Dtwn/wO4wNERyB
EZw8DTWXshfzQw71EGCw+iYRZux2hiZ7tsNtouN6nG25LSa8//7a4mzcVwWEJjiJ
0gebUOS8DYmJ5Zl/w9sMLoARAsXkWxqw16+i3qbNRWtOmvWtwpeXbG2Lg9WjqfwW
SQnd9h6jO2CIc5qERC1ZGa4+/6TFFnKWKiYVQdqHt+zJMXgHlsuPJtWp7CQWR+eN
FO3RQeA1bgUy7Z2qYAdD+9qMOG0cjPaiE7SzPDpoh3aSUah+rEIq6LK106BsLPr+
tAjuMuNZjW569T6CnMJHH8PpyPnwUuC5u4baul0Vtt9Cp5NPmsTH6XFb95y1R/zT
gfDeB4x2Td5q/NNjVOKx8uJx1yM66rLh8sY+K4biwNKCwHrsN8W2rIhHsp3qTNxW
KqlTXD4iCzxi/xINoRheCkUK1mEt7q1GLsCL5zyRtpJA6W/dgEAV8+cwi9AdAYWP
NFMcjc7fKJc7FGMNrMDs/Rc/1z9hFh+eGEb0EFhc+k/I8OWRsQveYdTAwqOaJHSB
Fy1ChJGpmzB6HErb2hEqE0FNgVk5z/2qkdFXiQe6Sp8pxXwJDBBYf9gU21Yq9QjM
JFeXG7AdYntfyze2hPODSwKTPDwXzI7Gclmpziot9NKxt+kbUXGyUUpojTyOE52p
Pf6kqeFo8m3yUg48qJVNoJDmUqiKKvL8v+9Z6iS2x5k9VVkSysOA4Ly8+uIyUcWQ
3liargmxQhmYoOweD9VBK0O0uZRaLaati5shggh3LADbOaJXxhkzQtWBYF7o8PRW
VuNq/JmIgUKJVvvCaz+UtDCKM99EfnHuK0IqKZ+BHnJrXl4JzT2EYifA2nmtxXZm
Bdf+kqCYh50tyWzwc1YaE4mQ2tYeOF1j0kRk6S2BH6nisk+mN5xUNiPpPa78+dMN
it4NdiZ0ecuJ0f2XvpLEijiXSwDEJsiq50QE0ckD/jtH1pkp5pi8aeAXcjReCSJc
z3/Z6VCRgq953piWgpUct7w2PKrTuVO4NM0oA3fsD6zGJ87Ll4QC5Z4FZgGO5hSs
rCCtxcN0z8fixprBsvTuBkbCpwLQYxyZdnnnZtCuGlHn8PthcoEI30GvY4iplcvK
BgKE1ItSlHM+Jthw7YOjWQ2T4VjP43BEzSCMR+8kQ8J0aKDkH955hF4yjRZz1RgV
o/ptrR4KmlmN6ZBuuQG0RbwhFe9YX+NE96rW8wpGhdWrA5vrLcBD6efO4wkHE8I7
t9h5Nq8Fk7Mq0p/OzjTHeZXwVECfS/mpGC6e4YeF6OXhi98o6qC0rwwMQV0TTrCF
Zng3PLn1Ovv9WYIVi+kNnzKG8y2DQtOsD6Aj+LP+GnUODezMVGCPVVVchj5RCrs6
ZJF6fIgOFh3CQMPw5sL5lH5R0trGnEwzRfTqUomJn0M8krPd2CWaIH/0shl1KGrb
aou0uTgFOChrju6/1/HjBCi9wSmfx01n2nAyre8j1wyzkE6vAXyiGzjv/pb0AM+/
DKeJH7ZXqsttm6bTrqkFTU+Lzh6iUKDSe1K6bSp7sn6PPixhaF8nRrzc8YNrLCNo
9zZrGkWVpUCZIgWfOVFcfM2rjcF1COcBOM+knDu/smX4vPAhcP6jh07ELUr5+RpW
kE4zN/ZEit3pqHrjMQCcruI2WzyAlhLLfGUXE/Ok0FIYR9dcsm6et8EfZbsLn2uZ
RGHK3JcjpdNCMgE9Yc88F8TM5ANrMwu9iOkiXAN14127ZxOLMvp9TEUuyQOOGMGW
ZqGHCnsfjgrEuHj+ttKoPJQPW9KFkOM2G/D6JG3Rys3wfwQzM9B5l7xOmf7mn8rk
7tZH3AtGI4Ia34AG2y6Xs13AJxGTixLwZRjoAmyPAdXMDBPLZsrS/x28otBkAGEX
+o1QyNHd0eoSHM2FN87BUwvMCwTCwEMrVdLHEGvzUDoJnOKXVW8WPkVsm5z2jZV1
Lj9s8xrV4Y8XrV1CJceV1ByN8oXjcoSglByqdVvLQEtGNG6oWmWITfIXGMNq7Z3F
hzlAzIKTFaPoBxmINy7nWuOmxBE3UDEvwPTgjY0uzrALkBU1bkKkQoe4uwDbhfNA
UON53f8zXiFDMe8yT9Ec1f+/J5jBQsTZMLBTGyUQP+rKBvjUEK6bRF04CFj/lWzh
1ZcSNBE7a1G7U5533FiyTNv6hJXdMzwOMn9rlLYAyevIbdtj93eCdsgZSdOUOmMm
IiauiDbvJUcp5/drtXNTZbxn6Il6ZJl8cNCRgbKpUDE60kp8MjL0zvM2wIW7SiDY
z9ob3WM7ghWwGxhyhYDD1+5MEyJET1HnNHrgFTHhpO0c6VWrahKto1ZsxjVX+ANP
8IatguuawAGPJszkp04T83zrBmgTI2JPndkXP/ZUoP9EmHBSvRFFUGWZQDC/mi1o
Tmjtfd1YcQvkM9vO9FnfDbMQaC/3bEvyg5FpNJhNSKoQQ00KL+9EBro0YqUYZajc
g/hzxd4Ltzgh296ZKN5wsczSvJlNnbURR8nDqV65L3mytRI6mWAb9YLSSzvg7TkJ
MYVdQjrIdQpmrrIHoWb4hTDnq6RXjVX89R+EyZvvejixnJTcNYaxW8/QQFo/e35M
/492G2nfOiSanb308r3c4wZbYCMcDGx3DgYBlFw4goMfy/Asfbao6aUQZUNLYQfL
rykFXJ2x9nzUTkpwM3zBHs+hdHZsocCsm0uCcc0EPYmRMtLxBSeCq4KnDwxOT4vf
vR8QrAvFdt//75bSa/8AnCSWVggGu7CdfuJCAcI346j4xS54yOnhbHpe1TWW/oFn
75hPbHp1OWZFF7Z/svXNo1vdid2hfN7cfoBuhWcRvS2OIKXtXZItKE+CDORIvNJe
z9bYDHa6hIW497kTsfO3Mqs6dLblgmZwFT8zNsy4VGidB6sEI+HSZEMpVZruyzVZ
Y7XnMRxUiqVcKtb1SGwF9os0lh02M5gz7oVtQLBra/hDMX6xsUuV1RBNtn1Mcmfl
lY27wK/4lMDbPq5v/Bi/4CTgcfAaBpivIsNcqIu49t2PfQ70p5LlaqQEKDrA35yE
S5Pq3oXtpIJHr3klB9z2jJHV5cFstkydngW4ET2RE9O5W1gd8QulQdzWQJf8GPU5
JqIstQ7snRiuRJeAObvp4PEaGaAt1EBte2EHYTUJIRXC6+jPJWUw4Ayy86Q0J8he
2twzwQUAmnRCsEX2eMiacA3MRTb7/oGoKfZ4H993km+Kir7YjX8JSoqLmV6rDP+9
J9jsfp7jJg3gReoBAy7NIriYzJrFP84cRFCRmsrutTQjDIxrYiA/UBKEThwTn0kr
4ufAptzv/A5pAH6gv0N5PFhR2Fc3KEW/812w806fIp/+ZPApXUrVltFybU86yx7u
Bb4HePMNY9qzas0kzKbwJphvHnmAoOaZ3GmmoDCE6wJp79N2U4emHwtMOdJSDahW
r9m8Jrylp9Eyq7wghY2YJcR8tWAWW9gHMFmc/akrT65AZdRgdJ/WFWT2n6MIOuti
+Hsxm83ehGq7SV0PpELVWQX/mJecrfa+2NMIdSa8O0YfYrxWPdQYsThGjD9q6BW0
h9tjn5oi4n2fBFzWoyVYaLfiSEV7qqZmFf2dX+9VaLpoOJvekHQgQxizFCfx4k5g
9R997eFkKgNJSLsOYbOTZ9i3CYeOsC2lH205d+7phhVjSPdpPpIpW5TV8XSIjFpI
ERkEJUdm1zCPoONFJekSm2e2s70vwKtFBI5IIZ0rBVmN6DTfFvkzZDVP4EXyO1VK
A8B+wGZP82ExvtFUM+Q59xDCulNgvWj4jKbmgKP+4eXT4c3rEPL6iJJ6jaxb5JfF
uvGnfQrHUlPBBZQKl/dsRuULmA/5t7VBhDe3hPIqlsQo/ToKK5u/7yZAmVWCa3J/
meU2xFR0Bg1+oD65lWvvxEAkfJFwgIBIfoF3bZhvMNV/ylZ1vs2801jSEqbO1SYr
6TU1MkC4gamkDZJu9K9iGKkBLx8/zEufak73n59o3KOxTqnYdsyqMzelkjbKStxZ
jcKfK7vzdT90Fmn2gCmqldKfAgFYDzQGmoD6D15j6rOaU7O/2LISNsbTr13/KvXm
IcfSdWT4tTCHoaBZXScSZiLLyEq0/OgOGjLH8GiqaYpERi+T4MCgzv+uu6QWIlno
LITNYHKST8y6sYMNEkr9r/eAgSMrDv1GFVM6erUrjMpd2Qg7DBfeGjtgwI+0vCBk
TdEB1iDqnEfRrqD+IQzDGINcOZbXo+1GAMRLERdB3ExqnJHh0a5xhD3d/0f+twnG
hSEDzB0+9Yl2aTVSlpToEjE2m8TfUbpeNlWeIhDJNfOhKrAqGfzbmdgNDTBXCUMz
arxMh5GK2PLI1l8OSKAW0sGZal0QdxReavthgLCvdlJFO2lrXer+BzH1EcFmxM3S
2BW0JEjzSqveTsOqc1ICB0sHwqhxTdjy20xXH7njoa/LnRsHBZYw/UQeYfgeiiQ7
sVmUVdMLjTvbdFBSgljmmDLS2loO9NgCd/Fxhz261C/7IbgK/mfY3XAihLWWMB5B
rmHAOaDqoN5DNdNTyIWkhffqkXJOj6W+Q76jVHudJwzsoLFhauUmz9xeDiXvfymw
Q/yCbO0v5Lirys7Dm+YhXxNu4qMHMvf5CcO8UBj6Ds3cXcTwRbgtXbCnCMaQ3YYT
cY52N47xEwyaYH/KGFMwcTlcdkdM3Hli2yqvMaJdD1aWpZ5Mx34byvGTly55RCz+
12n4b6h1e7LmRPEG35f0VraY0rv+ZO2TxNTqZa81XrbtFdPFlHISVZERlfdhD8yE
Naa/2Q4QN5l+iafV6/F/W0sXfmybSSjmnkf+JYQQXTme86+YhEA9/H+qqbKkWxal
/cEe87hp+9f6iJimoTDCBjns0uSGfz4ONjowMjectBAz1QnUFvkdkfRQqdlc9qb2
zDKW8zR0eu1O26TvNt4uzNWHuZf7hpPrvDRbgt04YHJvAzRxbRP+sFWLv2XvMsgz
4Z0uPjHZFk3RkkZxwxv35ESxOgG1KJv43cC9g3OhYzilEAmpK4RKmnuN5r1jwEUE
MVBu82SNi5qjYAVDzXGaCdXLNklapNqQYoJbxfLCNMlB+ipxBotesbGAKdyqvxRG
ncNPteZlNPXytmH7ahfcUyORe644l7HUhZcdYWv8lVl9QuSCDzk3JAjhgmllvl90
hvDH8TymQgArf0BlK+QFGU6+XHqqg1PaUPBnI0k48giiqCfpzOJM8CoimlJWNeag
CvGk4ndMb4RzyE+2EvMwxp3FyMYSShzQO9VgzapeGJHlIbnmnzgC8cwTuj74GQ2Y
4cpuU3c3G73bHQAoI5vhOYUWKRf27D/IENAbftYHNcEs/QiJo5yfW2TPotGcX8pX
Hn/VYbrSNksgvcdLLPdFpqBQM34IpdOUco6u/hqhx/uD7sLI5305SQs6Asa1w63L
kXtuLdVYNXmwDwwXq4DEnrFa+5/a+n+xBC5TnWkyQW+3M40vnpmZ5fizsXGyF6xI
hTqG7oNoWgmbB8qZLAf3aKAa1hqGKUvqQZIKCRlXutEuqzTjFDpfRIQJdhx5+qFT
ZGu7CY4uCinLqPXYse7IAU5W+s7kLLu5nZ+O5kWBpLLSxnbcM/BiqmY0BqVS3tvr
o8ljDGm0XIKOWQOg0EwZfgZwrA+Z18rDXiHg7ZI8s8K6A5Lp2TQcNll+1TfniqjA
2FxfQ7FkVz53WcYZz/ig0jmfG2IZtHrez5ieRgF9CCLbWD0Nv+BF1nJR3s3TMbNa
qhcAd0/SFjfXgXMzQVVWbpwBIX30tZTPGKljxGv3wZIeI2dY3H1+k8CqqJe6UZF2
19BYPUpFUj4SLKGO1vlpGXR9FWBtOZiZMz9H/dk2jYOyirvEnWLNJUQe1ZAVbA9u
LwXBUEF4Zaie4mLSsqZEnlt0Dzs/UV1HpOW3n07Yv1oNg7YKtohrpjb2sCJJKBKI
R4iTiQ4SWNSJq1YaYcB4nljOEo9WrJc0HooDOoigzG2kxVet1xEgXIYwkTcaSw0Y
kXA5TlyM67COVlsrSRgq7369X2Higg2mR2MwIQzCCDxEC5gPuXqLHQ1OrOd6NXXA
wuawds+AIyMkagAjti2IeF3IEgMaQWqET+x9NMoH9kC7gG3BSTc31/cCVhQKjt82
vtFQs2Ju5cLfh4ZdmftI58ljhED4P+GQNiI/sqby0re1gBNyw5FJKQ92Qbwgt8Au
dgFG39Vjj64tCGx73mPCLpFCWj/RSD2DZgJ6SstbGX1uPkL36bbR7vrVXpYXYLwR
rYTaoH8nTAxuAiFUMD1sOuT8uw9f9PirgNFIwE2OhDDgnZOqaF++UfSFo63rb273
j/xuPcp380xtCGIYC04DGoIgyYo3fbNhKdSwx4zZRo35AAjegKboCuNe2F05OFwj
8O2NqAUBRJK+WKe7ypblYxyMH+KimW3H8SiNiylkHg6tXu9Op9UMUKaQm88MeqjY
ha1IxYJl22x/2NzdOQ74XZhU1n2dOxvCA4DvshXsj++kap8+RF2ZJd1iPclz/Wue
PSgVntEjCFJDb1ANpHWdcjoh+YUKza5IUD2AZ4jEIZFpgPlK7T17nE7ct9wADE+X
vIRyOZQpeM5ekKB8c6aMRq7LgykEBA9NNLreAR7sOVQPxcg+Dk6dFhyWUnSaNA+b
659VFQv8hwRVv5IiWmfGMfS73MtOOqMjJz6CZmawdcaQW6aZL0pWtj6DnhbHLM1e
2k8wBTnIi24lrLT1AiGS3sZyIpqHOSz1DTK9UaUfA4PFEZqhHLt4lLDj6hnsB9kI
kypMRayv/QWQ0W4fTrk4o0Waq6ZTVOcz9UEK3Q8SoNUwJFi8cPHRSw+2GihV9DTO
Yw5aW0TsJVPpwlKwD2yJEf2vnXZAwDAGC8YzcIloGRXFBk4FE1daf/ivqVLtry35
tnXkTas7aIpDk5+E9ki7ZEfduQDMQ5z8KsNLV+2e/meqSyXwZhwulRbuisMAClTk
EIzQylJjzF2hSPBQE93J1sknwLQhM8INLX/+uoKY15ePq4l8RiZ35yhTG5+fa15l
kl+ILIaMdgEas9xzb6vvLbD2iQHXL3I6N1+Ga2p64snlrJ3K3E5kkjGDXI0Or+S8
sKW9x4D5NFIynKPdKYLZ2vsuHrJaehKql2XzZgULaKxgYycavlTIe6sOYdzIeB9Z
os7rZfpq2DNHesehfdALID5HVx3KP1ozieSiJ4IFYW4ns8nnMKTyI8Zdan4j6O3s
APCKceVHpTn6yBaeM+5ZnCZOOGqVJsb3Sak6txJjcC4q3DnOLBTFZ16QDd4fHru+
mqQ2AM35PC4aXkaHG9oE4iEdndfPeVXT3RPz+P4QL6RvZTV+qS6FCq93qHFyW33C
SFYj7HU3IFdMU7YeKph4iiWaQaAq1sOIU4JwcaCk6aN6aNxCSdOxgSn8at6B6pid
YwZRpYEdPch+B0u9MbRbOcWh6rudOov4itq3hpssvZ7zAApXdH030skgsMXkj7jM
pIz9gXeTZ3sQ4X4mMNBU+7YuxVFPpVsn+fRYiJnsVXhbmcJUJ4CuwcKwxPoqrsXI
fqDJvpj5tPvG/97vDg/lrsqRWtgZGJeUXmeq5NFJvD24YTIyCBJ6gy0cxwIjd/Bw
mcGkXeQKwi/MM6yUplm8d7AeqwjYKcqEQaEW623gfdcdNNZgDcJR57LM1g8g5Z6O
7lqa0tCzRq5Hguw2NLw2Ud12Gd/5AF2i/RbtdRty8gSJUzEcFgUGgkMl4BklOC5Q
pnlfrSE4ImbtESstC6/qrnnNb7xN/jfrCKMCu1QUkKKhTtKiaDJR4Px+6wFOcVyJ
qojm45WrWAN6KdAXJvg1YMZnr1/nolQ9uZ/9dSBFcIgC9WA8Is2GElaUmqh7QeDD
BThSesAauzgtubE1DBFpUkNtqkKsLoYmoUSa/IgbE8WmUSOrJYaNY56EkikXSJwT
fM7BzVEJzwI0vhGta6CI5D8oACKs8ypdm/7QfeqatYjl3KWtqdXwapha8yqbQV61
gFv9ImhyI1XGTZM+TiQbyhQceDkFQ2PQUUeebNON2tEYZIGhRfsxSMn2TTiEm7MB
0l+n6hMeeUaCGD0qeRRCALn3G/4Dh/h1eMgFQV39JT0MRJrsZnmspht0YY5WLFNh
6CxomYrY1gCvvzzrsnyCogKKL7ne05PhXQi+31cw1mrcdzDtHaHMEBnYm5+qlHrp
ccc6IHo3A9h7RMBOhYzAXFU7V6SPhbp72j4Jd7WOTcuYsWOAdxSdfycY3q6ORJqd
FA8tO7qDztps2IPCxoqy16p5lJ7hhcKvmWPbx1NB5oOYfAqr2bVlWL+HwF8k+mZ7
Obxx8V/helB49kpNPPH8okJQy06655SfmC5w9yKT8IRocgUVp88OupDDShzoP8UC
DWpb/xWyX/CsvEh8s45oPRm+8dF6f1gccXM6BVhRZGudzTT8HECIn8yOPb/Fk+Hy
3ozvbHhsed/uEyWajUfHaZSy6XhJKdmkwV7m4E5F5tGr9X1pA43GUVuk8uHl3pYk
iT/HFNjKTriO56pGio6NElrXeKJLmvEE6vcMS+vGNGiLVaD5nsjj3qsxIIoCLPHj
jcp+IS9U4inNL0taA2ZxtoT7u5mXCJ3hkB9PkniJKhIQfTgyJvqauoQWbI39R2jw
hcwYoHlZUnhqLPfLnl9RwU7+gB0NGwlqBI0KTuvhYmu6xVa1An7xCziXIKULL6Xh
bYBZUdU1JYtnWv8V2LzS7khUh07yESi7CR4FKBg1NXbmZ1r6ZkJ9Rv/KvBi7Oh3a
OYBG6bB2VRTsERdhEADA0tStdlcMVS5nE3okgU1NzsRltJM79vJ8Q1ImmNmuFuOw
hFVjJ80gj+dbimXzTTmp170vWVmZT3GH80jNkbSJKSurub5ukDDcRSIK5Ax6qHRx
31A58TslVzFywFL+9epNSaoZ1piBMa8ICijr3HteB7W9o6QBys96BafjDe/LrHA9
dLoOYVTYmLPyU9U/sX+mXNcpTyG2DvOhf3vLHC6GrTWW+chWKuCBNUejtDU3txEd
+AE2WlhX9g1TpfzgsRo3J1HW7s8Gpp7m0fVqxQMGVAonvII5FSHSQQtI+vqzkxzq
luWiMreQFEZ3Y9Ktms8L20E3V/xl2skvO4x8Tfe5pp2U+NN/SkIip6gXvR4S/GhE
x9dcftrhnrLRWoh0pJqjRvgc2A4KwZCNW5xj+N86kC/B8g7OFdN+badNDgTajpps
n+XRMvBLy1msPLeZnydpVfXHkm7Xc/ugpOQ4FFAEKwgV9FwLlA28phrp1gwyNVMe
XbVuW7NtCxfwS65AdnI4wvLGqqmIx0j29C74GNrU9FAg4NxjMSWUpvYdWrNwj3vc
ggtT8MlWxr6NyVVwDamD48dRImU3j1fgpvy25J+iCdvPmm6fr+DbwbDz8y8Gk6lS
l+XCPV8J24ibXK7nWyNJNpbSm0oMl9Y3Q+xcotpffj5rBiO/YjhvPRdPHoyON8SI
CWp5NWrR5y7xrvwqAGCIpfFZxTgaS18l7BrNZdjBVkudeOQm6NtJaFRqS2GDBf2k
aioEDs+Y8+dAMDuAndh2Cy/sDt7mJ82ZGvufgkrJedEQL0PZKQSpWZNuL/YdrOnf
PcvCHVeJTtvfLV//F1mU/Z3eX2/Yd9I+PzcymEmmn+s5r5ckfLXoaz3BK6+Xcbzm
WRHZE4O0JesGj8tBu0vQ/ho4qcJ0BDTFK0uGg2iS2aqKpIS33h2cFACCMVMKhMaI
3jP3eqaBGme/LpkLtlWVGi7jddAh1JtruqAXmzBCOpRQ3JAOqITQKCzPeSHCDXyB
NWalm+9dHG0JZgY/CNQN0MCIBVZ6x9uFuFL0mFlrMPIWztAS8kTGaDaBXYC5IdGB
oHux+QfBxCvEFM5bC8esqrax8slj81piyEB94rRMj99lgXtznR9M0SBzV2n27Dkn
7RxzuxagAAi7H+E09pcz5s4NVrl+fN3364II89z83VqQT6EAHXem5wVYMP7UD6rx
NECjCas5ASWa30g7HqG5cMCYGAiqoZGd6zzBkgJutfs96IW+rUT8R0+eNKUSZnA9
h1tme8YfpviAQUzVvABDvj/XeP5M5MKR4GIro67UIxgcHAdJJ9dLU3teYfcGbBOe
D0FB8K+9Ef6O/NLbJtP/+o0XGN9MeUZtYThx5saYl9Io215wJRglzhAFbNsOfHX9
rVWj6mrCJhi3qK0Ilq6teL7itvB05g3Ed12Vf/oHIjC6jf7DcCXlgwKZ283QZiDo
oct/tCpxqCquZoxg60shldjLMWiyj/JjQ0yy+do3cvdDpCiBJr+P351TmkXxdRmL
PnesZnRAfGbH+R8utqxMG/I8d+gZrgW901KLt8BpeH2rHyaMbQOIMCIDJCsroJwH
h8gjeG0vQdOcnfvl1ptD/9gfyBLJcRfdBd4QQ2EyYynakH+Zfhe9T2HS0bd5wgxl
JFWcCUPZq1Q16GFOyd9Ernr1PvHYKGiRV27Ey3iB+LDHjID7UQJfwvotmaXciscu
SVOeTQ13JW5+Fyt3TpsM0kY+ck+s63bCBm7yDrH/flAPrKPqScq0W2/8+Jqjkgqj
tpj2U0m9muHvtb8z/XUeL250r9x8944V4CfKCvqJC5BhwjXgwtNGrsYzPImMBrbG
23mbkInLbD/Hrb4Aa4ww6ZO+hp8vtweSXxpeL38BR7/aankzQLpweqDjdJHo0AVN
57b4hToFzY6nQOBz7ZxXGHVZYp0gIm6p7bdv8ynGCtzYTWPS55xZCfKrvGB6aiNj
TZSkVxI8vxOo/cBnIF4zeB1Swe6t05n762Seof/su5iP2zUr8e7J/SWe8N5uaShM
3/msos0pbUg4NNhRV9KnF7OsesrGcvwg5BUmech957RLAIkkbYAVae5ysHGDOMwo
slcZQCrSJIHf/qk33FEP1xuhqkjk38yxBdUw6C6gkGyfZrIqP7UDHWnj6JbfOuSK
49LMtGrkbNE4/IP34AIukBDqDI/Rk6xmif0F90venUZNcJ5r6jf/WmI7G9yaZPbu
47ZM9VSWfxvCLj6h2h8+pNciCpDxHLCVsNpWi7XNi7ZoIo8tHdpNuDd98MfoPonh
AkegaQ2IqsKdnokhCD61wKa1n+wnrnVRAKarTBBKXAK77oO13KhbbNQkXQPQQ9Ss
9BYDq9JKnWjGqwqb+MV/8faGVhq61AG3KEEjuwKtxKdjq3aIboANo1VZfXNLLP37
Y2boA5WkoQ1RFGZB/9XSgYXACGQDBpglwfsUYzBH8GXHvhIG1504H0dXfkIo14Wa
poIl2LViqp8mUh3oynOh1IoM+8KquiX107VKl92WMJhOdJmHSQC7veMCeoPl1yi+
1xDYCXTbOSMbIe6MDxRoeZZkC5JzPzyV9oe7NMjLvbadEWcM1iXmiEAGdHnf5wYN
lr5z+hfwdU3yxX7LZQK4O0sRlB8i7DfOhrSe9fDSHdLjzxQ2zQzngGDmwBlPZItV
Y/39NJrsgA6OG0PRMf4+ltLZUKxXMIyUsOuiNRLtQNlSxukcv/rK7RrG6q/vkBLH
X/gIXOuyp5pDObQy7huufQyXOvolD7AsQIjzIK+86pGdKtF1DNlEWrzGewL8W5Z1
zJIBKkt9PbZLn8CTU7BDW2UXGH4qT7POtFnoDUVV/QV6BOOusWkqOFIHmkYvLJ48
/40gvhHOeq+5G+TIKS7sq2erpC6cClqk2Qy5Y3eZEEUBz9jejCCRsEbcyYv7ixGW
8N+BfdQzH0Fwzm2cVQwkkHbVXh1ie+F31l4yjmvkn/pV2wNGRyqX7f10lssn47Ja
kiHW2kZYpCH46C3Dpxs5cZyQbz2L8U6yD4Vj0NhmerAdQcd16/gs0HFSKkwE8A3g
3r0fAaG7Mi/yA31YNWPgaX/4NT6zZOlp3CNb06KB+mbB4XcYlwd6JHyLa+lCWGhT
DEZAAWRyFV0gz9uJMEyt3ps2gzbWomnDq6J8zILdeI9nJzebATA+DRF923FeRykr
LzvGDIknLMGciZAtMh2QgGwbyAf87Ulu4q1WoBH5UIN4Ef8TPZU1KFxA0XcF7k+O
qxV/Pqr8fJ5eM44CXCHx3yN1WWN5gF2Sh575+wT2Tfr+H8Kgud1n+f6GMlKRq8f+
JY2+167UhUwHxaRDD9UR10eZppelr+2F7+4GR5OiMRAy3W0sQDjfJ/oy+cUynBrn
nJJex0yvtdRGiKj08eFqgoj99QTyKY7mOJWldPioTtpy8usjamR+6EASTnD8vXW2
G1FvXBtsvTDiNd2yC++6u8SCeKqkuIdDAM/4DUZFcIM/5B0pOe/sxkgbTVrC4jHB
4UJ1sW6xCOcYQm8e6mNPtYC8tqSuFQOO2tydLRZTYty2aw6fxLpAKS+zm04Y8VYO
/8amsxPeW+vKCyioL2KQylKNNeiDtsezhWBoiLXyYCe7IF5PDikwsBO9eEheCfz8
A5dEIeXWlgAxJZrQcu8FiSyrpisE3MzAFEz7o2j1vHnayuTs75deIyUDrfZFrtsw
RmBvg9VdijEhuHe3ZRQ6wk4Yp/g/xw9TeovUl/2zUtt5/D0jf9Jqc7CL8raQKjJj
pfJG0uyHFne2FtsQ9xoAR3deO2oumpWx5Hbcp/NVpODITL6vuZAqqTMusil3wnaz
JXcp4IFQT0CHhQ9+bnM8J3xzF5TyvnWkLdvlA2JRqziPhx97l9+zfz3GHxDuIKhh
Q+bijgG824MO4C1L485/eBpeq234nQDwsmwvx08MvBr829B20QvJa6NumLRf/sM5
DUkSxhqIF1+cMv+wvoanFMkaCPr+DL/T69f1jpNLsZKLm+bRh+abfML5h4h6dx2s
49+cv0hWGXu/mh/7zXGkrkzC8mi5ZdqUZIco6E1T55k349SWqVliuIffMFvG2xsj
kzj+kdBXhMrvRC3JpItWMkXgHWlMGs4Wnp7BwajF3htX8Fi7CG49BO/ekn1bGvG8
Yxyhv0EUHaRH+zvoktiDDk1eS1r5f3klflB1SUoIq8VPJqPGqBlGOFk7xoUazLsP
LaJtUg/sZhDheAVXMTXvaYEyUSP9CoM8UpgsZUucHggdpFgtMqNFS7OIJWx92hKk
j6cIU/S8jK75VhVJkoa1uUrovISZFn1DveIXvWb6Aaud1GeDt0DjdUElFx8+sO6q
T4u0/O0DEznu3YGbajpsE7i9L/ZdD44lHNrqtTbOqxcXiEe7hdmq5QyAC9nWtIIo
Cp9KVDNNIzuaYLkWiKhjERsuY5ZjDVwUt0Ry0ji/Mow589w4MR1TU8MpCd66DAtS
XGy92jrtyWsPAbTwHbZDGtV3DFGXEdjHEr6cLLZZ66DrtCaJ01UR/FFnd/+Cvgej
pWlH8XZi915eJ+V3wgRpm3sXAXOoSv0OMIw9D8qiYR7PAgIh0bTFRDgVAe8uK83j
PfcudGz1UomdRzF6M48PdyrHHyVE0gkqJeOqHFpl4HOUtjqbdrW/rPgotEMtNvKP
oWT++tBSlSsm5odnWCRgxppahhESM45+KPLYJUM4qZzYGBr1cd7c8t1hNV2zhTRc
oJ62Xz98g+3q3OGl0df3O0yAuBUo1w9ilfUBirFoEBflKmp/YM9+DRgp9E3Rr0ze
KQZQr8NJWiF1xJ7sXqrysCt9PUUf/zJ6lhtHD6gt23+S6TawHFuizSjaGyMbK0Ce
vZJPRTG1JsmIoZ5+7/W4ZZkb5TJrXgctwJ3S/ZGzwLwO0lRHbDIlUNcStOFNwzhH
Le1YVELFdLdxylLSv6pN6kwXALYtkRDeUa0I40UUzH9YI9mKjSh4/jrq3792JDtg
Rbt2XfVZ80BU6SvU5tdsxHceQKJjryRvvGPVR9jTxYmNwdUqjkmOt4NF1xkwixEp
cCcm30+wDJNunAOzO25M96Mn0588m9YFecBhYWvLqTSf6iMCv5c2dU92fqHCWJaR
JbTXozHGVuSvXI2jYSjUJ9CYVPPCtnT6KS3WlnKDGPin2aGCyxxuaTmMABn52RPr
fT5LMt8YAc6rbDmdXFhhfwVdt9sBzzmUXE23G+UEgU9OuREK5RC2QYwmp+9Aeorn
eTfb35dHttoR4KjPraZnyS5PGRUDd2wlurWjAcloquUsC6vTcXPizYpjZacVWv48
cuhZREQqZdncDc8fwXvoY7SQzs/1Jk94ufQ9T7KJeLh4jZ1KTWJgLhk6C97J8dTu
xOExOaSrUFWfeu+i6n0QSSdWFh82z5zhIJen1oVd5A7khkBrZdltXi9B/6sNUMkg
wxfumg+By9lE8a86aPTa/RjT8bVoZkm1xE1nfKBxF04/84Ea3M3CF1OJTn3jO0Bj
cwX9DxPaECPQBEAKvESuF9UBzDf7nWrkpqDG4Wer+GBPDqS9/Pt0ITp9jbjXK2AS
2vE74ctdhVj+DNUfzZjtkltbrKJP1jvHvpaUbycBQoaioJ+Gb/LFbNAmPfke3dy/
tYc2VkTNB+hEUiCawijW/nhWdXja2upZFMGh3f9D8qJWE8vEnIktqaxRMfKjjx5l
T3AcLNsFcYlHAKWRuxSSqtiOfbEKA739almVKUg6g6cUurPjOyK0Q7J97YtFMUTr
/F24UeOT3Zab8x/DhOa2BYLz4fMWHNq5Us+fhbqkFtOIpsEb8GkiHs8Gc5kJHMl/
vV33XpMZO4gHTZhs8yaFzrVetMsLpVEwqXjK78L9tS+p9GPFRBZEhppIRfkvxXoy
kJEQVkJgT4aPw16nUikDK/BJx9Qstje2EgcXblienEkiYeImXonKgqtAW4gKajIQ
XtAiDYqq8zGnZMDqbOMToGf4DMSOq2Nk7+RorbHr8bajlbOzGgvxsvEcw8xJM40W
YRx8BClrLWYEFfzPt+C7Fw6l32/goGhjzn8sO5WOjQFXh2HsRLRui8NCtJ0/5Lp1
vMgAbOBEtr9F0xTNENEko7jaavs5TSExmWPciFzDWd2dGijU5m2+FXPKf/dK6Hwz
exfE+x/nMadLUT2EqwYFM5dnc/Ox385kMTC6FX/K5ANXlgy7OAoNaVDJJkcYBiLv
Y0q0IiUjuhJ+OPSoz48F/ZvXScSaH/nBzYCi0XDK4sbCRmuflFOL64WFEN3lKIiD
UQmxmmKAj07xJILY8p7a9PO19sw84y5opAw1bV7AewZmbWCryUVr126ULdkFl3ZS
hj+YkvDIVzV7RrKr3snpmqeUefBkiSiY6m/eUatYsZJIZ/DtDAzAR4LnX0Faq+EN
cewY7Xh0A+danSeKnuLwRIqZXz2FHMAXaRMu4SYpeAdWpMKgZKUNeCNy5DCDtT5L
j8dQjPylqkmLFfXmkz3zUbHLu14dtLuM6TTXwTaqHS8QtWsfG5TygoJJLxhZFGIv
CSC2hxOkJS/xU5Kye57891pFooBwh61G4nlM2Z0cxeI4SwKPJ66PpuvjHJlWgIiv
AMv8/bqKWenlFF3uJ2VuHsqR9Y4giVKCkoqLSL33CqU4ZSwxCXtxThY5xDIMGPuc
UnVHUHBDPvfXeLvvLeAlU+HvuRI/ZSrmKkXdjVdV+Do9myaff6benpH6kuNty47y
uE50VtDs/QXycOFweH1hRivz9ZMiVNZa/O/55eeTafIv88NO6sciumBkLQTHz06b
jixw+nmJ+FKz6LkesKBnbjCFPN5wbC9aVf9oOUdGF9a9WyU1hhdPbx9NZgCFQoNA
9hkFnWJM0ge0KcTdvFV9QlgrYBKX+CcM6d4gc+ACKQoVcDL411aHyvTK9I7Chhl9
1D6oSo78NIcQpgA/rcsiCYE9j6baqRfqgFBXYJPeCe/LjlM2lHAzOWTpIbAH7g2D
DF5NmzfjRHkR3JwUBjr9Zhtq+dcKKNLlCLFeHLtR270zCSoGppU9KiH5tfWz1dz6
CRAHvopRMFp06n/1wD0YxzV5FsQikprcbKNBKNoyT615LguCT6QCHU5idlCourbC
8u6ESXlIWqHwB9q0h2rXUEniH0GTWnBSKgQhtUdOYfWOVlorrmCZIdwsVHeXwKTo
owTuIrNqAc7dC6jR9GiwiXZPtIET7AUbv2lPmz7m8gqs2Zoxu9K/x0fn9BswnK5Q
c6/Afpvg4CrQUkQjF031N4qVGyGJiiopb/wW0OzLVVOSBzEB9AjIlJ6DVPRb1m7G
EHkJKbIswhrQvhAJR6s7geOn5JDY4JSNTBUWLBDYNuRTGTHyKdFncS6zejw7vDxH
IdE8/iu0xD1wGFbA2FaK5aAypU8Zw6lU9IYM0b0D8x2rYrmmMyfZrLJRi6kIKfiu
h30Poeeq3JC0ZQqsnwH1oDc87o6VoUxa7z4OB0rP4hiPChyEh4H+DnaVJEoWF8lJ
oA0RJ4Nyb8L6bj5OPTaeXyLD6/KL/lI/LiDDvEskWk0ZKd2Q9FqdcguNvMlBa+BG
rYNKHfgFIRJ7tiLjNcuqxfTr5BX+9fMWcKx4jj1nCUsb3q2buj4xqyLVhwxdDUOC
weqTTEBw6ceFfkqLmcPNIOhn1JhAA10fm7AgO9THDLqE7t4jDr7kXvNfC4iH3Yz3
sBG93yFBuGrqOHt+O2VAGARBtx+uRJuESe6AU1oFcdKsF+O0Pt3nwuzl0rXuKSmR
RG/wwk4A+i6UrhWSMV9HWwHpvyBjp4sCMARGTAgSMy9fBye80fIcOkhQr4mYb9bb
e5ZmrbpTrmKbT+Hlu7jlkqKy7CQnTJYDvBpp7gzuZNGq96nsHfGVm0jh/hFSRL34
pjOMTVIJw8ZYoaHG6djSod8YmyuA7kmnI12TRHHnroV/HeQW+6SHnUZDgDymfFOr
U3D+k2W+ZX4k9GWdV7WhVcrxwgpMwpKUbrYShL45VQfs6DUzM7zR45eaFqtN5xGj
hGXrjHgG+LSczloQU6i/Plsm8Q8roLISzPDKxjjSFh2UZUj6es/T4o5eGGec8Fe/
F7CFDDUr1Ia1F5/e2iwIJKxE3Gp3kQZ4E4MdfQdMUVRjmAkq74rRvfJ5tXSOgBOA
Uz3mbo6Owp63qTxQXY0ItSL1OvZdyqKmwhyJPVajAbRDrxpL6Fz8Ngwo+NlnRfqB
FOBdwsCjkAtOFLh4wTvO2KXPEz+D2aLWNXNhjv7dQbj5USmhmBmW/GWE4QRcWMik
GUkZ2vNlg6kpnQZ8AMFol8Q5vjSVbsUR2ZfZjVS+gYQNrrtVOczKTB+e6WXivria
8d8a6RPOYDNDDWkKaaFPLFC+hxOWo56yrEbaHTl5bTYsUTeXOuQeS0AB14eahtB5
fB3jx15kwNYsk6FLSj4EFaOYEwSQVTUDTJhePYUuUDTgsPRymP4pIOrtzEuMN6/O
zkOh3rdJjHrWkAR9tPlLCjFsldi8IpOUaJDXgcmiaDHpzBOUHWtQjlFEk5zzNyKu
xS0+GtUj8c6F7cf1uDiM+MnesT3LpzgbsIyME+yn81ort8zby79CSGrmHSnsqvwo
dX+z2ut5baocaFptmUNmcAgyVKhbNx7OGFY42YG/XKSykyvknPO2bfbBA/XtaVTK
dqZglp3qvSa2aqAtWzILoHePy9TXKHRdsujIeEqFZzA1ruY7lXFiLvdUM3rvpnIP
kF+OEj8e+UZYw3Z0UCbUeHCSJrjq//K+lXqy2bvuTjJiFfBplAtlootGFK8xsKBS
7T+1QIieBdCu2W8HqNbiwtyxkslQc7hH6ipP5ivNKNfzyEsVSiV9FzkOrK6gn/c+
ZJugw7M+JS71TKC09Lp+vwL06Tyg4sNp2XkjZRf0escCwFT3mlXMNkNjMhc1PuGE
NgAH4VSTMvzB5pRpX2aJarjSKoiSz5YcM+KvxFkl26Y25Q0JhHxAurAN6l4wKGTm
eqPdcKpBakg/a3dG9rmgxRfKwxVimEJJ3EfRAFH65mY5zdLWe8h+J5Cs91vLj1L8
CxNVSa54zfud/r3Jjui3c50vBLhsjlRFGN0lPPFM8r9E67ck/Sz0hRK8w9d0IWl0
kIg9T52kwPxJkThgOnGzwVNRymtgotPvksdYKsSfpxOorzvO8PkiPe2VeVIyIbM1
HCFVaKc3qU2ugbrKREtWGSmknZq+6gZtxg8UoA8qRhEv8QM5fIt3GlWst8IXlRP9
jILUsKwWWI8AAMRXvbpikq/u7Gr8eF5q2H5Q50U6BOxZjbNu9fPmi7Y4/lMtPHA2
pA1RgMnQoH0vrbvIntDKpy0pleOQCh/Z3eJ2vxu6JElHKhD4ft7TrN912smMPO1t
g2EZM7PLGpQDn5DcTcZa4GklGtUkqAvlXRJgCVsmoxKIE9Hd0r8iXzlzZfnjwrdb
wzf7TXlBwWG9jfP8y3ueiHD06k+2vKAVd+IRRrP/8iSJhGJTG0hbM0FG182yuzpq
LRy3dg5H1vuyh+twJ56+zQPdh4H83LZdheApa3NQOT2RiqcnuODdAcqfOsjcQCc4
OtrYTkoBVr17TtWHxPeiTtUgLRBxfGyEse6gVYX8O2mllfVavKnptiTe4XIFNOQX
WWMs9QGQPMAu68z1WAXdekdc4MZi+Pw4NtETMmfBooGa69qL6Ud62Ntw2dkPGQwz
RSL5PcIbpgZJv7O23rbXfB0M1LnQk8VQ8bI09LkJWqjUisCor9e4TIH/z+uR2Vnb
cwAFdOfOHPh4Hz2lZpwslCBSqHZgevqXRSaFJfbQTL9EbccZlWX3eyLl/AvNgGiq
fwSZXPivcAkCQLEADnO9/XdA8vM53MCkLUaGP2JXCT50UJn/ztzLnH5pGM+LKBW9
aoejj44JpGuv1ygPH6rq4eGQHcrPu9U0zNKk/QSyflV887Gmbo1WaVF1m3NUTQGL
QfS74+zuTGCcnmYdEGqsXAmK49v/GxoTVCdDwp9NYyw+jo9h4gHxYW5JAsv/So86
LliSQxpvk1yr08Vmnr5nWR+hb8R88/zlk2M9r3joWz/WwWxj4PbfP3/05pbuWWgf
8egPZuLRfZ9YZq5JjXZMv0p9SfjdDPXWPHHSwshsNaNM0fb2/wS09j1uzdVc4DZc
VlUUFK+ch+h7Iv9Ao8accZXLxcBcsWKOr2KbI6yZ/DNajFhxNuMb76oNJ2PhWDTs
K8VJmSQIXELHk/xCmA+l0VChVaAM2DyObeN+OD9UqLO2/7P6uG+VOJiK2pjnXAF9
F1VQ+gfHzqjZh+dnD9vKhy2i4TaiST5Wm6Pbay+kezROBheRm8xdXEUOHaxBPFYn
jxFAg1GjJJTgawGdWFeq+lDMcvoiLj3ANibhXFU1yVhpC3Qi2aB3MWkB9pwerqaB
RkJziEhcn9n8PYJ8uJZ4BoWNSRlCvXib0zZrhE7igOYYUiCou3HYt6EPdaVrAZXn
ooKMAyZx45XBN887G7F/dLurtO9IBjc34UdvEopzwp4cEj4M6zFc9j2vA5mj+K6F
Kf10jSsp8tRaveXsmdC2YBliaooCWPHHGe72y3GX+ferOGc8O9hBqoQREa0hnL0E
X2sNAprJHU8QVI9ct7dVyg7j0hJriYGCtC2sFNmGP9vRyUFwgMwjIhJReGy/0bGv
oDTBacdLHn0Tim6QVwOvURcYMS9DVEHFHDgWMbbBNFl/MDp3g5WiJIw8CSsEDSfS
9hrj0EerzuWRHeYxRD5M83gxPnhOMT4mfJfI6NQAVUgr/PHA+H84RYKouFkeKBKE
r0kCtg1VqsU8N6fG2a5HQlxP2t6hAGuij8kLjYJrRMDCjxBMkrqX1VcjvvRQCm2a
VkKfDpwCJjgZeevcgVyvGarFrgUCMHdzGu3coMaUS9i3zLxvfT7q+le+x/gFyllW
zS55CHGz9p5pLxquUTnnCjV5ZEp4AAQiVkfX9dHG13CqzSl1CJB5KtfIxpWNCW67
jVMphAgSmWNoWFzjMziOS1lYxR/0/BGuKy3E6KGbT+lIrkC7iKjJrjB/x01iuX5q
nwM8m08ipP2L5hl2t4VqIxwFGz83JaOvMBQmnN93oTI0fnIMumOax7MsLUHjYPzK
ivexh3j2lRqJhwJC/lmv5zgfDNcScg7SJyb8NtIBOQKAl8D4m/Uq74MXC9dASJv+
31gZp6rUk91mxTtJado8qBcG5ecGfjIQVbwmF5ZB00H7rWWf8WQpsQ3/D5MoiL4M
CzIgnepAQF4Bc3Pw9VNpZnfDLGZ3gxYLmJwZahrxDwC1LDol+qKpksifiw9F5e5a
Y1V3Prsapoh7DlU4Zn8Bc2UzbSyT8gfzyw6PCAC1ARHDMVQHa/uDEyGsv2HKm7H8
uFWNT/SAqi64Y3tgYDf54ygO2uSmCG1D8Cyb2AugieF/rUgZNI0jnHNOEiqSRvJF
RDmRphtHMaDNdbLnhuT1NqUoJeTjIWzZATr/2e/8xdIKNrNjtEdML7sae91qRP3D
kHOKeRDsjB99k7LjYn0M4SfP6SzuH57cTzcWWryxfwCoIvL+lQxo4w+80CEIC+O8
eQzdxUKYfrIW2prcopKUBsyZair34OES+hElh2FaNZknOlg1WMhwVvdFaj+ldxxt
hCLKAFrOPH24Vh0U9LTp3jqUfhk6re5G3z+8w6l5NUkEL83/e8SwtqEK0VL9Ddz7
pS/lvq1AJpFG/VFy2WOZn+p9zPfLq1mlOdfUpT7eQODJwOc8T9gpSLTyjcQIK+0G
hApuciAhy4obM6UQ1HPv96+W73UgJ6yvbZU6k3U1r0ZgY62O/zLaPv3AUq/Lpuj5
7gGNVaVWGPCsvQc2XW6JvPJd6bxIzG8GYNBfdiSbk5vjxYU4FTFKo13cwBkEmFlY
0WsgRIBn1SSpWCIUit6NnhsMRrHirDWH2n9fZ32owpmY6SlH1JP4aVgc7K9jYHgw
LgKThbt5PQJ6mAVOLZK96tHN+ILK5OuQb0e/8XJs1yvL7PEzwYFGC/nktaWfTQg3
FPamDCHwFB6+dj52Zen7tGC59y1yC0AGh9sLR9V26T4oGHVnA8tfErWQ02QLqYYL
ZXYfunJHz1kJn7BLvOf5CMwVdjya/r42Y+wmLp8SICJBW7BYb1Z0QxctVQosZwpF
VJ7aah4/41W72SpsLuM7Hh3tbAexhdWpfDNKMhMJ/HCpRpyJBrbjr2gCBL/qCWtO
uBC3WXNBd4t8EQAtpbOWU6F33qZo8UycPS8/PxPNZyH1XZePwk0UuA4NnSVi9tAE
Y8ug0HXoEzQh3/OvpLSNksWMu3f+SHt3xC3nK74DP/jtw8US9t683FMJeXqm+CZ0
basJ7giVDq7TIBfKMiv7F3OgjRwMJZIsLPF/O42hqLw1Lm4A7aZI/9PbRGJSdxFw
OLQJ5x3I7gE3oDogD90wxnU6+pYZRbmQ4SxeIgFgewS+m0pJ5hN4PS4005sN7YiQ
XNIPAtt/0Rkglwx6EIHc+JZb0rzlIEFJFCloV4O2euyXejlX1A4UZfrQLLZHUc+I
ZV6UhScPKNu+VkqvF/PRODRxKomnQKN6mlYBWdFbOZ/R6qby6hB1X+XggmpUV2yb
XgUISX6m5bw57RcPRLc+TLfAs0TLVpWMm7PaNwkEqHurFu6DT7caf1lcxK2KyNuV
UZ4n5pB0rmh2ziPQuMXc45bGPxKkmHIKb8YvNwaJ0CoF0PRv1gK+3MmC66dR1aQi
5TNnzHWfc3YR0AvLhiusNi3KSklPIjk+GjhG1s0z4/PBioJ3PhOa+MRarnBMOydh
isjNOQTdCueAnA7aeBexty6qN7jiHtNRg3ropreZxTYnyRgFVh0pJve6WhkeaqZI
Ugh8N4LSe/0hPHEUjWyslqZi3XoCvdKqCO4U6o5jLUYzYB9xpShBl1Dwrcikqch8
jkooFpYQfUhCM4Y6OwJX6+ZZFi2AF43pGE72yN3cbe0w99nv+y2vCNPh9fSlzIKe
b+DdHJra+9z+D5TwabMFdlRulmj4pG7AOegMPQBuizr2qqTPgnABB506bL75M3UH
sj9MVTc3MLcF9Dk/jt3gY5SK2K8Y21qcZAEVxA397kDWTmLFhMkzdyXOWxlnYf2W
6yEhnPId9mDDjNJov9WMkkAsOtN4C9cHgh8+/wCUyKI2aqrvo4H1ZuEINuubFjv6
MpsiWzvVU/FnDTOp/9uzRzt34+/IBLUUcxmi3gHrhtJ1y84ZJ5H0ZJw4msWNqlEJ
kUtZbtrLzy00/kxeHsDytQxNmcmgJEVfSmBLL8r7L46hQC2I3HZYZW/yV5jcifzy
wBBOLEsXXJ33s04wc3PO8oV9/SiR4WeFyxLjA/HI33VncqUOpcOY4C9kFkrTI2dV
QDqCi3lyst6DgnDAvsBPNn0mTIxlK5kjBkl9Xm6kZiBs4/Z8ppp8cFPav42sztbg
lxZQ/9aVJkkeWCLN6ByOGZ55g+DC17/5w0Q8jgDrUxn5WL3tG56GlmgtpjE0TM4J
tp1Du1EOsTd4BYdqjgav3jEmoeNJ7rfMOv3izVUnXjUYpWbuTkrqTc1oyyEvL9te
1SGH3ZpdU9PnAHZIhP7ElsMNqGy1PbK/nOfQylcC60J0rcYe0JRuXgWiZLBX+V9M
SIdYp1CfxhumWS5kHuN3ExHmH1wl2CMMmi6lRVKe3V6aQpR7/Y6RwjLI21KvE8fx
VxHMlhUBg6PBk4xJgwDELimB6SW6aVBi19FhAV8amo1IFxWCiT2V4A7yDJoSO7u2
EK6u0x66pWY6rkkq41ojU7ffYPQsjXlJSRiADWYSdzs5c2XlRUbDMcLZ5CiZVykl
l6XEvida1UGHqRF2X+RkFIi1zbKBZLKQPfsbL5ATajXRpg1OCp43zay8SAzeeQ4f
lC0wtnmOnerAgiGVnOVddnLXilqzyE79WI9MBQ9eVbOJjjQLPqbgcVHiS79UwGDa
/zptFPfnXlfAnnpLfzLVqm8K9plBfROcuCa3hv0GCYONCAT7f3l/YE5XFMtBEp5q
c8cCmdf3KYBDFlxAwtyxDuz+kXVGHG3u7JCqNBVdR6U7DKsmDnY3aWgf9/X7THe6
h4FqER6c/EkqEhSjBflerOWmi3BM05i9VMetruP1B8m3v2KlabAp8kxsTbALK3Z5
j/XST/X6sEPALXh5vLA5ZY+YJuAE7KqX9G/ImNFjqOwijPWpet8Eh1PfVFF1WHBM
qYOAQgQu2a0hvmh+L+TZRmkFAsj6wtzZHqzvNbq/qpkLynJ23GGwQs3rVoOl/0Hv
zd0YEMalH0P3QtM4KHq0M+CWTmN9kJWVOpjBpKvtNnflEccU9RC0PNRQVTnqbq9B
a1MPM0vINbDG24/0TFiAKr7mLK3apSbLTvaDabBmv9k48/FOYUBFpGAXNNr8GqXb
JG6XufytX2TiA5wo5M0KCqJ6AU6SKPyIDW0J25hWgyTBzSCQ3c/tYXeeoGcVdxVQ
fnRgp4FJGbj4NPAOIKQTMzRuBTy+xGuivniVkGkl8izbLWvE5pl7z1qMImjUByY3
rOE+GjRprPd1c3DXPPdi65vPHHlFqVY4uKqZgZD19xM/Y7V67+JsXZ6vjZW50dyu
VbDjrctgasck+fkARBz9bhsa1ehrVTBaVsVPHX8tYk6LQQeAR8PSjr1tPw1jJTbt
jgpthnR1MaHcIsF3ka0v4SdXt8w4kBkl/xOr9k8Ub93XLnnFPYO8gxzE3eZFQDRx
IpkJ4XZwyrfDa+vVPEwnTq/KYFmWW5EReqVCpCsrUrpl0LNwPbKyFt9hGYMlS4ed
SQUbN4tUafIqNx9tZ9DsobBmxPXwGvUqXZ0N4BtkhC0+EtTPeMtDEXw9xYweU6IU
fAyD/Y71X892zVLAIkKBtU2AHz0NL5Wb9l5YU/FeLR3547hl6zBQPXiBXyEhU7aR
mydyZkjwdiBRZa5TgkySTKFdaWYSbt/yPYI3h7mTv3m1+PvbfUfV7pqEuF1972aQ
sgKgr5ZTCEnLyr8bvJtRG7c7XxvQAIO4G7eVDECTMPNtqeHBbK4JI1hrk5Uoy/Ih
FCfNN7XnxPgir0i7Ze4RAP2qnOjP17eWcYU7Nw8kW90tWv828cZ2qWk0cNWqj99L
wPNJDqchHSP+MDlftWEzdAqrFkZ7WPfSPMU4hKeM+9yGCM86wjIESL72Dx4TiMb1
ivoIi2T2xv/5XyXlEh6sQtDTrZjULXug8b3vafzo5YvSTiVLbnGMAMRU0FJ5y+Ot
KXzus2C/olS3ti7qhhp/mbECDvaKBC15GGpOqOSoRAb9/SR0ayFS9J6tVfQmu5sK
ita0sxDKmSWlQ4DzZAwxQH+f1o6oSNO4oxTsVQX1t6sDqIhlH3UEBWLnvPUc3XRv
4kW8nWwLNkHIXdwp+zeZHjCyb2QWHSV1cdWIvk9WTlcHe3WMwbHDTG04YV5Dq8L6
CisZlfBmFlVzVjlOJCpLxLb69gga7Ri0j6ErGnNiNWcO4zWlKk7X0c9Hne5Iojnz
hjIxywJUvdVJnJsFOnPvSE95Yh3ykZukPdpF6VHq606IIQPGiJMtA0QZsnxngiHg
t66yMDUlpJme3Q21B8R5fylqf4+1hol8FeLo9n2es9Q1sRQVzjv/H6FPm05cyLGX
tJzHKkDbwQYdn+FsOs8hNvcZbJ/myx+wsvrLWFE90ip6ShfkasZplXbEwsP0xzA+
zpzaX14+Bu694tcaN4xXuVGjEC1EOYzErMforGTus3L5PyE3fX2mIP2CmhN84rdj
/H0L8vlPKiCp3u2dHeI5maNXb47YEqqWzIV86mrZP/vxZK6Yy9C8kS+YMeK8BZVm
H/6QgqjXkYtP87G216Q6LIVY5dcmwgpk6FEJIrj55z/vuUqS4yyvgCQiU66qYHny
nbs2Dsl+hNPDY0jNE6iPL9twyP81IQc5hEeY9hzCceNezyz1KsH3vrElILWu+Ns4
axydZ/6oVXfHyrDwfY3n3UGXr6b+zDCWbwaFVdSfFo+q/4e22MX5aokZ1+a6YhSm
OZdkmBgPoeIip0Gm3AQMUGkxQFvEKhI5yxUqUd+L7Mq6Rn6vdhLm1FTz5XTjg8Ns
7aC2OJsjVXQASAkhtMB+9u8spv8gpkQrmbkx6EeiRrbQAulEb8ftJs6+Wu1c3f3S
r9/MEOafboBF3ft4x9rj6DR9X82ZSrsNQPbZSYZIuMMK/5PaSs1ePI2k7kk/MPA7
nrWeiEDmdyXuqAk5r2bJKSnEc/LlethzUxqxmG4ay/SkV34zkDgcqQkAwHvsBM4h
LOw+L6cBer8cCr/Sxek6pg+Kxt4DAJ502J3IK/ILUms5FGogFA5h45mTTqCw+5jN
pYIs1dUJlvA3/8mhw8Hke176gNvhl+RSLhji0vCwbLf/Gos2RpnotIoNlAh5KcCs
BvSfMPtNOReTbxqWx0cGpkau0aiB3KvT23fAhFPiVUdJ/fSGh71GCI2JxmytvxJz
Gvqx8LBLPI22hqWHsKZXYQPOOr+jBVuLXiZhDwuQsyp2Oeg60zbFveSGm+NEoMhA
HiNcODNPtCC40mcm8pmb9V+zwMRPGoRxw2bhhHiHumhpNEHmGYNAEo8yxe5foZTG
hyuRO59BLHzPMPWCJ+gkySjdiy2XUBlJnekRkQP2jaf+hIRnUjGKOZ2dlDkGCCxP
KUxtXUMDeptU+6R6K/iI6HvOGY6Tk6vCI+OPDejs8YcAp6vrsK35vrrDQDIwuGtx
AD9+2+e/wfywcCAWVi3Ke/8Hcd6Hd0/qDa52HS83LIzWzZPQ2zMvbrxJTAKcn8q3
6FZR4A15JRisI+Lhx19Q7LhUYeft1oh709hkVFwwHRqjUG9BVuyaOMKIFXMnDWp2
2Tdr6o9HdAYob8rbmwUS2bkBn3tjj0/jN01djWfslANGFvjYEYbc3YjNo/i+s2NY
gybFzuMHSn/d16bQL2B/548BHh5zEKUUqv6QSoZq67cUmaPjnwBvi30FL3FvNVNQ
HYnk2kdFORM+A6AmlbBYEnti0BGC5azs4XC1rLdqjs7IfWxpi9dITPQza/kBgC+U
cfAzJ1bdzs3x6TWEeCGKAf2Wnbu7X/FLfnSBGp2WxYopjU89v/2hPXbGFWy3sDQH
clWz+BCwGzIr28Fx45Vw1rV14l6XwKH/4xxWRVR1KQdNRxWPsjLYSkZ4vC+oWSKN
U6S3JVB71wsJMSHUWzl7rWG6bT66K/yrBdyKVhT8rFxukXLq5y1JhCSsEQj50pnJ
+Wd2OkgEVHFjXEUk02BaN6U1bjQV3U89euHq6rwzn1nfjA6SqvhvKk+HqS5qNeGF
9IyOyO9ZXGQwjwekMPxJ10uaO5pnNnRA7EGzP8hNEr2njKkQJufZI7uVuYqO5pMv
L8B7YilpAywhPm5pCHqPHBjxuLrI75mIbLVj1cfSmys3s0hvZAQ1llldqim8GFLW
9n2zIuJM7MaDRvDvuNYxQRFT4xNH7g9TlJKkmr/9fNoZnB6Gk/H8Kv4j15zkqzTy
0sacByib4mhBk+8d0j18/U1Bfm4CMmLnkkpsLDE9KKbMXMAz0KSKT/jouTBJDB4S
sPkSw5pc0UnreHJfve2d5uMrVwBDgfmxge723wmYldTW4Z0l2T++nnuobTkcoteA
l0zQgKfj5XhBfaKd0l05PyD1lIfba2QSh79V0TjTOzAVCWEsuuPm/cAYAMfy9xSC
KHjSjDAQoVAGZc61w6V4f6qav6SSoJScQOxXiGEUheCvfo5xcLTLzEGpR8E43GR7
0f+XElZtVB9PRw/bAtutkTYFhyxYSowvOOycjtMQNycSnT5/4Rop58FXdupCq9Ls
fG17hhPFhzcL26LgjMkpc42E6nhOBgPqQhMo8EQImEtSNu80tk+jZSEipkGI4srO
4fnwW/TmjCBvqFzOf5DTbNhftSAtKutru9giDi+DvQgO/CAKRnHlxfSiUlBe4/Ui
/qgeD5tDmroFWq7mMVCxwg6AF1JA9adAPOFE2gp5hnymNToSa9oJEfRA81ig9T+G
sY6o7dkOhgDE/EaIPr376CsL+JXIWglZF5/gcg+qUrgGQgd+XuO1wBfcEe9G4hCC
/r7bNCfUC3ojEvMhr2aKJ0m2hm9Jlr2od5CgU+qH7aSY/9GAbv8VxGlbhH588/Wo
o2jmPBGC4Xmef9E76xq+OXwWzWj2ZfYW39Gb0bTUwmuXRYvoCGDju/fCrx4dzNjX
5x94l0M1pelJYZLLjYvaG+/mngdE20fbWYaLxTSvhPu4SqkYJh5SQTZxND8Wn/2W
fwUFmlhWkD8ikc3L8dOnb8JOsZI5Dhi9/dhUMdRTyey1mX6q2Y4MU6DHtXa5bCyO
euteKH7qSZtsdXOAz2t8PIM2Ud2Pqh2IbMfxW6vXgeOop8OAesNpSWr2C4fVdidY
Xl8snkrJt8Efk+hDz/sZHcQwfR4qVUUvZJgghKChQ14q2T9ButiIgvOGo3NhiwDT
Kf0zHcsl6pK1c4dugEKtkD1+9obvlQwm1TnKqpKrOB7MAb5p/2Ye3WoL2/RqVVVh
RatuPke8sglWWVjULfbvib6EnTQHubUNTpKn7bu8p5okU1nmbXxmRaFGiuofTAbJ
+2XPTUAi4K/gCBT2GdxCiydzl71ce+q5O35dDKs0qr1HQyHXYEf2NWYRJfTNMwpN
stwbf2YKgDOta8iBGKP/iLPB8fZbcGvB5xh6+Wwi+5qX3t/LSv61DVLC1WdBGU3L
hf+lv/8tJ9xS/Qefq5vRV5rRcCE8N0dt6SY5qtXA2pJdDEIsl+P20OTjKPLTiD1b
KQDABdJCeiv1SBNR5bbPyjbtg+xL89Lm5BBjpgukZLr+SjIRzD84aTffQH717sJ2
LJ7UyC4/llEHzH2G0QXSVCtjhZqwC/jkCeI6NY18cJfiMc6JkFxRYBoeIabdsKLQ
u6gg6w6QslNdGObBUMXmASqGPmKi0SxxSpqhjaQ10QuCxIJzzeHwPYnKmpNebVMS
U1SrMF7YYcxvK2juOJ07TNnNsD6+BDTPdao+3wZtAlF5laDNMSFE5sfTbcoQ2cR7
6MCJyAxEyAQBVJ0OvJ9iCBSqNeYkEBwKEP+Tj5iNcHqbBmdhJ9BxAZs0OqM9X6og
Rq+P9F+W+tobaIqfBO0eOtlR6StebRyQ8PNla+Vpt0GH/Vdh0OJy6FBeW6K56Fw5
p6C5ybO3ZmV/hcav5X3xQe/xgWaRnJcfdVAXlj0d5p5CjO+sSBUUURVCa54A2ug6
LkI5SvGG9MXCCeHBsRdVM66DsTWlkQYNF2q1iMn9S2bJZrQDlyCTq1Y6Rm0aG2/s
zAnIb6s8AB7DgULXtdB5g4+I9BaW1y47SMy8tyUkEzmNrJ4tzd+cg0D++488WYHm
yPcHSAg9GjdDyuK36Kwur8Xg2vU6K3FuaywEltgHYYx4iXuitWMxpUpzMlOa/o8J
J6UYdoSFLWgrhYfwmAWlk9gaOLiEqQfJirHVKWhytcjuQ6qLS710XwZ/NkCFy5/L
Ua0HJ89NUYx25K7u0uk/zlkG5TIhNNETu2j1THR3B7L6kXwLm8sYEfIqIPq7aAcx
I53LlRDBTh88YQ1SKPq8D7GjDabcyYxPUTIW1Chc94GPcoTsDUU18IrLajGg1BkP
g98TjzlXohqQDccxXVj6x8pCcnHwNuY1GznFz4vFCKZSx0lSWms97WGWQJqbjJbM
3YVWpzcMS0VQAngB32haVXOzFqlmwyToWBk21o0c96WCSCnBUnvOQAnKfeUEj/M5
cCye2FJ2D1a0SiuJCeislBtc58TcbxEU8jemNcIrXaYuGV67ZkPheMWIXr7ngKuu
MhNnHh8bJnMWwzj/CELKFuD1yogXzAsa7wqUa74MRrT3AIfzEfT9yRpTPo2vCLj3
pQg/IJ0HKaTQQwUUmo2eWDv27mdlcybvqux1nVghHInbCmp7qvbDGKhmgZe8xhfP
UCkI3zTejLhxgCjVR8IFpCK5tOY7rHZN1huR5Slw9kap3kJkbxHr2EdgfJ1bqIz2
Y9rtlrJ0MGd4UfvMNx9uEyhGDI17X7xDhBU53KurHow/VyACH4ZOtTW2R5dourv8
3ESy4jdCNoJjsGGBVXYW4ly6XbO9iMeROmiiVPyWEe6vaIeE6zCDNSrSzD/JaqhQ
mZ3E6zMYYkMEG3IjxO1EVhswYmQwVyCFzpr1i1z7VMLwexhnRXuvBsI0wt4hhuuJ
HFlVTvHtVztVEZSB6nIuyhqzZh8WGxLd4GTMgZssop4lHR6wJxxHV7U0WGY9xeGs
5ljordmjyAFMrnDQ75QmpUqDP5waFPxXWvAYx2Y4CE89OA5Ghx1/2fCpUDYbEUUC
d+UabRizUqM7AQ3BQg21R+vRn9VzabCVrOdWBCCNKLj2JxxSwaOtsyFvkGkYwC5N
3ohZKE9iHPCCnHgkpJlYHfeY+bU1y39gyHUI5sHga8uIrd3c0AzfGT3BfIi4Z7T7
wBl+4fHcC6/8niG5o2TvmYVomZGpHlTqeDaWbv0ElCkUiikO35tgkEDVATsyrWjW
4YIYqrjwA4MAYOcfmJM2KqdInN9wjjBipWwoQjIozjmpVukwCHY8FSGaChD9ORMW
OZMsAw9pqex9a1QCtN2gIIWgbXyFFet5P29A+iTfI8gYWIQguMGwQaDKWl+D6Lvy
lobLeEKKPsrtEZn2fgLUHZZphFsxTbyxkOisHOQVpAICzc1cuWC3idKQmeyrhEWV
OqivIYMBrNk5aExpEhDQotvrDpD21KIpnPTwDtFOgrN5TlErWLnZ93YdiLVcJSa6
hU1b5wyhNsIJRwVCWwPHOvxTdFd7eEEdNaHSfZ2ar+CmBFB/yoEYnPjy6RMp5ogh
nHVLAmH3ixnlIGjn0IVz3JmFE8MFqWXpIQ3FzVJzN0NmWQzmraPlBjDYzh1fgDkO
RPuey0nYPJcgrz5pXMYouDTBIb8ROfI6nU47vDHVlgnVnc8Ha/CI+Mu6Ik/u9S4G
ln9/GZM57AXU/3d1+Wiv6GYSqsij/a8i3mSOjttJBhd5KohjssMksTpEeT182BMq
IUAKuiDuu8+PzIpNvglQO2C6/8w7vHIg7QiHWjt5ITJFU5pJrwl23d4uSBDyX2em
+VmlzEkL/+VbJyX48l+CxsAtLv/S4yYyPEonH0h9wyX3Oe4KyMziOdDMomWw960l
ghZSSlLJe+oOv3QWGW1GI2PUDLGHsa8EaJzd0ADUaVxQpf2LYoXy359m5Cg2iNbb
fZRR90GH1D68Lp+aHclARMdtD9cziLf4Ovbt+8B3SLlJ+qsGRKBOL86AVv1MVHax
iHnfZtjbATVdu/SkuvysG70OcPwy+Pqx8Ig7k0zjyYgMFoKtWkY65xX+8aStnRBm
QNSSsV7naTHO8aJUPCGY3x9xZQEc51OnsgU9uVIsLmmD7io2SYLDh/gB2xbzfbAQ
Byr3NtXl+1eKTNEhD67IpM67/qRRzkdgIfmv8CCkGVwJaYEV0JDinn9o1OkTmPww
lnlnyDW3599V25rBfvPn8nkIi7W7nwBqpKxwt1rq9oqaG3TvP0p/mlWvtipLHGdE
26nrmth2YkGbsK+IV2wAoF1T0Ex4CnLytOXifnTW6l51goUS/m0/uYTtJa3lJUiM
unkj1K0TXt/gGEesaifqxVwgels1wUp7FIzJjjPqwIApSq14NfTgVUu9UHg3xUVV
igJk3fObBmm43sVYNFYd0vuhDGH46TdKjHLP7Ilpwd0JdTxTylTGXKNs4tnZd+md
12gbZPAq34JfFIEXfs4UhJ52e2ZEIEogK0vElWwCyYGcMK7UVt/w40H5jnP/LHI6
o8PePwTNxbY2vER1MYSnUkTfsRfxaAZEUI7HgwhlGvhNIkClXu7Wccgu/ioR9Gxw
BarpW0C1bRTBt9ilHk3IPPu2gv4TXdBAJoaVsJ0e6ZoWYTrSsFKX98LqJ3w1tlRz
Zidimc3YzNoZRluoW9nzVQnU6UcIzJ4HPY5nEajlKmmH6NGubwO+Jk0TYXOqlakL
ktFxIMlgg2f5hrRweWWif4ebZXAhnDhBT0JqLtTt1ZfI5bYAj+/DrXofoG8KQIli
Ug5QeJPiVxjtj8O1yqTr7t8q2MonYqktkCn/LdirRHTdSQjX4zVVEXLAqnA5wPQw
jZP5mIcuqliKBzbXOrP0RKMMNf2Sp32LPoMGjJD1spQD2tIhbSzxZdaKJJ5s7iiw
nvKS+VS5mMQ1TpOV11Innegmyfay/atYR9UAT5Wol4UgrMi0Eb6Hr8xoVbkq/F9h
RtuxYYQ/2xPbL+Eq0IAnrnlQV5PH3rmP/F0CpPvmDYiwRb9lmNftW8C68xwWlICU
CCvvkIsj9cpoIi9LzlTnRrlatu2vD3bsk+mFP0rlnaBofGVUbjUfC9yrVhXslvnZ
Kv2zqcOYttn6XDlZyZh1ueBKrdO16P0xO6/MCQ3xgs2TVRRmKRxnN8YhNGoj7446
7u8h5iwyT1iDArY/1yCxEnyy552EEk9LZ9UoB3EdQqnfoIyzvT/VORVYlXZxLT6C
xZlE4y0jCCijy62hpqsb0H2NJq4R5/9RQg73ltnM56b+Hi/guotYzxFQQXrX03U+
GzOR+pZRn0fbKLRePzyYEyNb9xfwwuMplfmM+1dxnc16GlKJBZYx0gZfztcZF828
bn/AOzh7MxxIkgadisqdP3L9Ek/ofjjBTZ0aPgGQ8e5eGrn1JvVJU48jIre754l8
eyXqcY1rB/blYyuDfFM+2og5VwMHOA5atpqI1249Cir7xF/50eicsdJBFWthgO4c
jNConz3TqPkpP+DS0SqX/SYxFRxAj176KsdiHQnCvSLVSluSK0MdZcm7DMAff81s
yeV4Oys9M+QsjZd1w1EtlCRrdWuth4ab5P0JpD9i+voaleYhFOYRVSqQBhaI5RSf
xmp3ywTj3eyHtRwO3x4uVbaG6M7r71o5GbjyUDT6uF7/ISVypt2C62MJm0ooZujA
z1G6NFrpT3y70BJ+O7F6riFBwfky7z/j/MwMrqFZlpUjhj4dQ/wKnkj2F2FVeJtq
tro+0HtMvmUfKgp5XufQwedlxaWxDvWxwdhAbd5/JgXELvSSJ4me/nBlrIqCu5LA
b11GYoRk0v3c3Zd9dMSKiDmMN+TYR1gPPgJZJcB/evG4j9AB98feTmqTQV5eLjs0
KPw0tShm1EW/9yAveV0FBKSgRZupeFj4pLFoGecnQnbByNMm8Q+C7v3tQG4eQITC
Blib5QiPT/HFRJhYXbG6r5Z4Dd862bPMQFHHNRe97BfQBUYLhgaTztRgX6wwERQk
W1qf+8BS7pmI29YEE6cRNZ0INYh9Fv16vUprmePgVnxS8C/4L83RYfzPkc58qsJv
esTh4MPZBmbMcsPrPVwi/k156L/3R+cEhR2VI6xVbFUbKIEc2g0z+2LEKlfWY8RS
O7lsxVgdV+VBHOmTiNY5/PLLqtGKklR6WDS3PFXKT8DQ3fF/FsMRL7tIjRLft+dr
XWHstNklsTdN9fHuaP3dG1lUPdmiVBbgs6EniS77IXD7VrbAbEoPPNjsL1SyoCcp
ujk50fQt29QNE9N/f+79NxrrPYO6u2+rFIqyqKQyBgXFy/fadaRp/D7wORmOnaON
kEZhrdE8dG4fphcs07ASvERgJLqHTaNghDyRfrpWC44sUMcks+CYcG8ztuCdHoZQ
JMjtsRqDpNab4CwchJ3cnznBRAR/+SZC23kCxI1lwD9xbsV54/A/avXLwCejtmhe
RdjCOBf+OHLCTKA+/Md0YPoQDodR5jwE3ztObbuLd4Rcc1dyrYu9CJ3WtNDS7hn5
rbW08YtzQd3TIxaryN1MJz/wRyN8k8wRd43f/O07Wjq8p+vz7SLCKx3HCcqKxH+h
Bv49qR+BTaqxOefa84IBkr1ppLjriCGwfGSYJh7PNfdBIISLQHji8Q+2K9pFtSGW
vecB7R4gPrjM388MOneLkXA5R+GBTBmOpFnpjv9+H0h5OMww5OYCQ/IvP+uOqbAk
tDjuKrD4BBXF1yvnu7PVK6+XGMRmVmwp8fulfnQiRtkfnjuW5nN1XoEtiEgL+leG
F9t1vjcDFnrh52HjBpnW7avnJs968TypriJliUjYT3Nm7phXLmOv31iXgXN/YcSq
rzLz4GJPkEkJYZYIiRX5wO2FCLs9NkXk1Lox/mN80QYWJDp88+DncMhbAkLoNvF9
l43cobWNWQ7Cwexk+gdSwoKzOQduBPfckODjap82qhjMyDBLJOESzdyyXmWtvK+Y
ySMXQ2NbtCKcwNP7f46FN35r+Wur/iH0dcs6aYiJfDRtvPP806dcdNbBJBFK8GLc
xLm6R97YkyNtqr0CSXU2uZf8p2QxxhCBqAa4KzxjlwQfT2tV8PeTPQovZnMqBUyD
1F5c0qduFBPGwTWnz0Zriw2rtn8TjDqDJgdI0mrPbh9+71m59e/jM7c8FhxicziU
sATJAtUgFHeDv2PppOjYVZHeMthgfszbqaHJ5ZJUy4RckBI8M+YiS04Or9c/iYE4
WRDfT3snilziU/ezTVTCuFMYiqC3E+KcVApSgkJOqtG34jvn2N7LEIfKuetaMBy0
QV1FgJ+geGnP6uV4ShJQFdSwu4mQWw8URVMN63pD7XDIcLOgcErNkEL02Z7SRq+3
VO3ErGjSNyFduSf+VUy7eP+T7DMbI9Aun6kTXfJBO1S8ZqRFo4QPLhDGnYcZVz8c
cuZHUScMq0R5Eko+xh3ZeC+MXFksLzDNUM27YzmYj6mZ+D+ju/u3eaOyYplIQqjx
ML/AyCidoKPOEIFb+A6/jYX2H4ZKkSK04J3MeBNmlqvk4hGSyK4PTn1vLRxYUyg7
XCxlF7xoEpybM1Hc1DrCs8fsOqhiemycFaPFggorLXwQDxCLXvYaFgyZlaUYyTba
SZy7tymakcPHnIc+4fzCeykPq+BZ8X/Ele9LIe7PUISme+kfE6j00cJrZYxuH4cy
xUrV23JK5aqjU/5DWewibdZH9RH1Z3tqBfOMoyXYmsgVCJlaf+mQWp//Y1TARgn/
3swxX4zvOEDzIESr0YgJBbpsh2uavcOPEt4GRjr/mDV3qscunuF5IFgWKQuHF7eq
FYZxCZpdbBxnFYUXwQALKHi13qsBc7XxH6cTLL3ZNhqPpfmUkD09WaKb8Y307xLa
hbdC/WQFCuAANGZ+eNVfI0/iGIJmgS8qO2MYuPoQWpICWBzUFu6aeYjUiArtCqhP
GU/nrwUUiF/HLj0yTLd3bk8rt9GbFfmU4XtFUf3hr4mkGyc6NTQLf5F0uP5yJOCm
eNPwVUy61Rw7fwHmWSn7lz0i/T8nh80wt92jS6KegSR0TIZnDKyoSTFWCu3LOfhV
bEgVDSzJDh72hBlep/2fr2+fXlkAxP7UKofNC1a7gHGW/uxGpFRKPq7A/D9rh5+/
IF+NiRmGzU5VqytNJtW5ZV/7KI0yNFAIMdvk9jX9QkgduM4JVKRjD4Mbw0aNeMcw
/58I9Itk1tpFmzQ5PyrSoo5Xs1tnk62/zSOa5iBvnf8XOWqX2rc/8gIVdBu0z14O
9gGjdZPWzrVNgk2agRusVgDpB4LQySmkgT0rJRw3VX5KM2zBcZFLJhj7I0I9L4SV
9oDNeuWgkn0zEi2OSTXca7hbjAwy1GU4Ftv7tpLmz8hCgpzbKsZY/+uPQuYkU+4e
wvTeQZT9KaFhLD+sTlb8jIhly7UhUxsCetEMHSF3xlyXAmqPGXGATNO8N97z8vWT
4hCfytvHELI4xOi6bIBaqkQcZtZXzM8FId1B50uvBmiK9CiD1A5Uwn0S5ZDzUhFH
ewLQKscGpTLvI6XBEG0X/473+GcpxDV3fTOlMl3Pj38QumsyJW60xO0ld+Yrb8ZD
pOxMOVWMmJpegsqs5YMMx4PNepA9tcJNeeLhiFSyCuJuPFmA6MGpOLGgnIPi7+z8
rajC/McoJ3hsy1IwE7LhLB/IkiOj3H95jCBSQdh87DZWZ2MOOMJ19AMIZzgOHGQd
nB4xt/UzbaZ/rhfVuOYVVhfib/ceLcA9I7b7VSzVgIWP7gE9kvYv33IG3zYgZHvu
klWWRswEi+sqsKya28DuI3aVw+cjpCGA18UTNzUMGG6DAjljZHAoEvAti6PtmEjd
zjqWimHmNTlG5O6re/3/NuzQUGhaAjDD5lBihliit5Pn1OLQzTA+aFJVdNETWUAf
mjoX15k5C/pz3QCWxzqp/cgi8xAmUXijFqEBdLZRHHbgVaO+nNo66VcPBkGpIGjy
H8cfjVBoROCZEx9XqWRCIz20w9Cll4OaPHLKHn/2UngQEUpHlDS/mDz+8ZmTKR6X
GYVdvZSf8GnYjF2falIpKo5qpCeY5zzdoQGf90U53MYGert+Gol8KmJEQJI9XBVH
yeSw4/IN2mHFudORNAFZGxvfd+R/W0rUBmSlxxvO6JHmueHpEPlt8QKUWIhJZRZz
cqTKTDBoqlMat/M9i8INQhkK8+zu84lEVHHTHHb8kAJzsCd2pJXJzOOso5Zj5V6Q
Kfv4XXQMfZT6mJM15pgFz23was7RgSz2o9nomPRPM0N/uCnG/ccOxnBXg8BFyyLi
jBm5H/+RUQMC8PdexOXrmy29eTLVxSrkwXyGSi6XB/tmmKqQBTPlJ32eRWFWGddb
42VwChfSahRmmwG3h7L31ACSJOJAoQDrkxRN5kwNDDRTX6IoAyRPoXz3ZkEC1bRC
IfRXC2oLTibF+BQysXW3gsRiaH7QAvaeEzvaCFxi828iafe0VgjdPtsrRjRRv+/W
+TqRmxQTiIkRFOoeUDpWeVxHYGxmNqtFJSZKAsImAMV/xnvLCQfJ9DugKTKyMrxG
0Xf4gv2o0qXz8v/jjsLAXSis/RxrrRR4aDpgEucSowNtlFgMu4YGLwiGiyWwDYuW
yDhJnvBHFr9Uwmzt4jukndok4jE/FRZgs3jRfqadH7e5xAQisbB4ib7wtkZGzsFi
jaAzgre8zcyjzXzISf8F9lqLvn8QJEz+09FTlR/NElSFprRmetq0hlCvTKUUKt7G
i+GRaH9Gu03Zlta/racj4ijHPYoOHJLTMyfj8YGEEqimKJhWvHOWhcy1+FRcbbqW
sy2xsjq88ZZTe+JTvHYaxNSpUCSptuu3cNdjydjssnuI9z8Of39IqOcNC2GY0f42
xVaYL0FVZRXcGXk04FY6/2YMIJVh9Rf9dGf99kS66lYChL/FkWwF02Dyfo0uukPM
URJulf9JjHszQMUIVosI/bFMLK4hlWu1Vbt98+Oerf6HK9IResv5LkXbV5z/TMHQ
jkGchJsOSSQNqbrjqw7C6nY9goe5krxzOjjvCPC2JgLy98FEg7/FzB55JZlWD4Bs
ZMPwW8rr0yRgeh108k2li2ogsMvT7VSNDxlhVZUqG8W66uv6Rh09ToIWfFgsOWrz
az0rGxC5JJFFzM9qGVSeHf+fBh87BGGwhMipRx0aN7Z7JXdYll4S/XoIDfbKOBJ1
NCMZztIl456pZFiV/hhibDvb59wxrlV5zb9UeO6wJPtW4391wPtPPuwQRLjzBTGt
iDnw8SMj/j7gq2NEOVPe/pgnWc/Rxt0FNbgVbqcioTUAXM/V70mqx3qNxTuUWs2o
YmXve2keJ3Dp2mASF73I/URe53uYcSraX3SsvE6mJZpxT4h8oO2Ck2KcK+wi5Xh+
YckH3y/pLJZJe45r6Qj7NxTFJtgWP02UmfUve3qXZrsHWUAAxGX1Y06zcApDFhmR
Qc0MNZlm3c46m5RxE75BEWHcv4v6Q+x9nROvhfnmAHesKRn4KRISbfZZZoVBCYSl
VeypZB2t3NmH8AaVIT7R0VmIEujVDUV9/rnoxHiItql8rFERvTlOIsz00yVLljHF
Xi4nM2bDtnQg4R+13B5BNwjWGyL+HFsuO80sgfLqqk5WSEpYAPGRtvjIiZYPouwz
UwLzzgqqQWtc/zBCMh9E3bDy3HCGe/M5e8VVyZPV96NZyqQrk+Xq4SJCrbsFVHqx
sY/kMAGCRgZWKFlmZDsy7LBvxt4uAN5E10R1A9YB8H65lOmNGVJ5OyALH9gZaysJ
Bj8IhqHHZ91WPZ0jpuhTxAO+TdxZAq+vaBydh3NA8HK59oe34aeC8b56fMETEaDy
1jw+Df9gtrDrmLIjDmdkOV21PQgeobI+PFo/vosVMLVCfiBpiDtPa9QNRQfzU227
Z8/fUwSFT5sp6gDG0gQfDT/dvMmX52cjpOBgKVJQ5AJJ4rkWZkwoyxlZA++iicaX
UVBDn7nY9srhljMOpSrPOHfOxocnyQjoHzbC7JBeSHluw6wLtmcgKz0H/vbmqu/Y
E1cFZqVxt7d5q+RJK1e+iew8h6C9UHXpqcBVSsvZVs7M9InM4uIcGLzkejYXLqvj
wXgh5nrFGA2qm3zfBicfxgI4/v++cdLPslH/DgZ8TQLaGEeqG53KaK6y6StQNAGd
6KKaZccmebowpuo3zGN8Bx5ebnrCuE3ZMffvkZnqf//AuiQcDLRdzjRp5a423P3k
bCwLxL13uot3KocE1XGIuo22upt9ypSFIbOS21/eytt5Y6y7zf6Vh5Tgv9SGVO0g
vA+6y5mVdmV1KuD/wQbazbKw0U3Spb8BpB7N+hHs4F+HD7kFSpEBvYr+mxArh7vC
mshZ+GSvdgP7ZQMZWxz2YLQjiotfNY7ohQq5n+LAuyAM95LQrrax7LlKjcKbyxXI
Bb1fwo+m7/Vo31eyqHklpQ77QpJ7SLQ8CnwS08fdHhBnz0lX7VdPubFuCjthA22r
fuSVOGtMFLq8rnXwco7ZTjOwDeQYVfTp+UkwqzvanN0Sn6X3Ikramwd0c9xFEYAR
5wgCLBX9yg+9+Vv8XMo90ZVAwB2RrRpPM8pbaDK7Yp9RnOyYyap181VpYUsqJjMQ
vbxxKa9BF1v/kW+NSYonfBTA2X2Fo0MV178zclzy8ogo4+ExTgHYgol0Q2NslNXP
tyR1Gg2E1e+BiH/YkNtr2pCjTCZaJ9y1mS8AfIwNUFX5GapUS9c4+fnT8xVdMnEr
uXneMmr5s5HQRJCoBZnoMo+3ORAS7eBrb3bOurXy8OkRJfvDmsqejRojYrLiKV7n
8yJ7yUOwBYOzlxhN7zbWTqIjrfjZtDlhn2ysyrIYSaWdj6W9S6wchXxCw5dNArFm
Y7B6pGrGwLalqeNo4YywI4PlgmdDJMjHyBXV3CrRT0tTs8HU3MKC1uMuUSnusVVH
LZvP8PHfzr9Ip4+Zg5s2Jl80hzQWqYWceYVO0+s7MG3ZhmndaNYtBk0RHt0PNRP+
KVTEG6IGSePUkl5N+fSTMDnsHziJ0RTe78EQfJSH+VQXtgJ3epPkOY+4GVxhkYRU
Citt7Ne2mOMwAYNTWNComFGq0tsrsWhA7HweQZ0OleloQInVlXJQSMz/KtwwZWPY
tTrWgIZ86TGNs+KZcum25d1owgFqjWgqMl++2HMPwLTMUNKrQmiMdd2FRQyeEW/8
Z8SQbDwmzmTwF2jDBAEVbpbqjylAgGJrrAioY1kxXIfEQR4POQwP1/yEF5fwmTsN
mA1fEdx2iY8az43EELp1wFidJj/gaQG26jtBls1RNXB5Pe5uE+bsFuAW7hXnaq+H
M9xFhvtUYFWj0dLkO5pLNnhfU1t8iI80OPuivMNgz7ErUgRntPqRptqCghTaGbA/
VmoMFYTthwJ19RzEyEkqrAh9kdMhoVyAHthKoZ2mDB6JKmJO04umXRln5X5yBbqM
wdS7wfI5mdxO5JByOtyhyt5H9dgTTrCWx+aV7GUY9W0FhRhbjEiwKX9lT5TlbsNt
P0CpQJ0hJHc4pHhTfy/0PePWLoBDnrtQGtrPxYNQSbG/0+oxqxqxZnYcYJFU6Q4B
3oXRoueLjvJnzzffxmU4cOjYPl++gbdFVcNQtpbil9m0xCGEm0KQ3zC8j9WKpm9n
Y8L1abC+IZXBPemHBoJHLFfIUdA9RYPJfLpSJI8HoFHV9PE1XY2eFwb0gCDv1iS5
eattryAzMb2WYHRvyLHW+1EMqkY7h+2M97cU5SRZwW0SeNxHCcBkgD6IJYqIOEdU
JF0JQbFqUEB9AeAfVEVrKTXKSqTd6IQ00jjo8orWhyAhgwmfmfUDcmQAwSj0Su1C
OVHoj/UtnSG3vHCxsI4Agjc49utU8tb6bw0Bn1TJ8t6Z3imWpY3eFT9S9eUV1qTc
LNes8FmnM0KnHA5EW/xlc2Eo0fcOMk2bsD/e64QY+EQNpm76oF+sacvGXJGQHaUN
60ooN7UVgmL2PyazaghMCcygopYcXuKp2qnimosyxb4I2PGW2IROZR1mQBwlGoFn
JZtd8PWXx8qu9Uijv62TWJwvbs31PMvtXILcYuOuESvtvL+3TRB4nYE9eNhI5dMH
a0obdvwRqE6sOg3Fnhq05jYO2KxfGnFfnkpsygZ9fGonuKO9YkSR28xKhdVvpbau
x3c0dXoRgB6JsExo/KPDuBO8nDhkLu687anGvMGHe/HkTo9B1u9lTSHRSToGc55l
QqOe5Wz3lqzS2x2gVyPkFys7nKmi5+ysR9oyb37yEacElFsYIQ4K5oHDBDSsKV+R
zrrVyLMNxDn3Rn0L9NRXCTYTPayeHyCtqwROyXri0azdIPFxjugFrKgeE8OFNsVC
iJuJqgIx7WgzYOZqoDyQSi33KOt+4JECxMJR4km+XFVw3sI297TJkTMuW0dWD3Wf
A4oEuNRrAhYPMEcdSBG99up5bR+rMk15HJIABHCpq+NmBl6xKHpJekUutY6kSY0q
9IAPM6OdFCe0h7krRMiHxK8L65xzZ4pnOZ0/4G3qYN16h0lDrSyURX8RUS+s3f+5
fJij4UaXHL3VE17yKSkR+XAMRAM26mfESF9WXzn6eWWWpYgoEmR3rlVQ5Bi5eAK2
idc3HjVpryRrwCsVioyUXWbg2HPZRaPIAbpuFuoYr+d7nw2MB0HTBp4zoJYjdaK7
7IYSFkcdMGfrmUoPWZSdKswVlhZf6iHZDDVMKiTAEgymexWFSXpFcNXvbOyznOTQ
G98eEw0H7VfyZ7HZbLY+nJjAML2gisWDAJY8Xnt4dIXucx1J/liH3NwojfOOlfjL
N8Qb3aqNmCkuSDQchRYQczTACCG8a7IkBwu6eTyZ7hrsg6suo2yHZ090DHGpBdE9
iBw9zWUWHdNR9Hrpov2ukDEY3pe2tKyu9LqOKL0ZUmTXX6cvkc4r26ixGUgqxhUl
9M1d9e5A4RYvqeKozUkazPmzES2sO+WAoaFM4fWsYxQvsgJS4QqPpCpofOmqf/T/
LXGB1MZlH/C+uGOinpkukd3MJgARCO6PT5nkpF25xH6jMchhButiffLwdoCWAseH
zALP0jvlzjHmSrAQLAtLQftDem3DPjWHOHhlK2iKRDeJJfidBdx7TTUiz9mF5p0V
QZF1oK6ZKl9PpRZABnkXQ7dmEko+4gzwKQUmJlRYIODwoinGjIGpXGrWpj3/56Ma
FJAc7p66rU0cwp9b26Y1L94VTdibIPzGudx2C+pi7vBhYyrHJrQk9cdVFAj+8bL9
9/recv41U4bqj9IW+SY6cNmd/vNim5BLGNnjxO02RNker0YYi74HGnLmvh0h0rTO
cOVW20BfElCLLplmsBqIgBdLlTbRX/Qyc8v98fmT1b/9Vxk4yJjqaRaRMs/sisl5
MY/2lGO1//B+a5suFjdsh7bZJvh5z0FA+uDfjn/MpG2HL/jKw+bcEtW2J5iDs4v+
N82Ddi+B2ZfWWHLneTqe9hgLaqYIeGLs2uHs5RQi8rcznnHDi+e+NGUOnlLjSmHd
CS5Wn0RpcCK+mej7qpivs2UHCB22DM3UajGFDSSbkEETqXTkLNGG3QQhbLfeNsZ8
Y7iEDS0zRc7WaVpo9FJElrqNa3sOSshtAyCgNv1t0f0DLSg60kRCwceuKbmo3dLc
CEcGMVz/bjuotMSjWBbx20T3s/b377fJyb/x7X6lLHbnt9ydUBSUm7iMAtqpuV3r
00qh3x8PRe+YXjZ9go5fijrTpgv2v4TxPJNLuYU6Db2iwdGv6Pa/A3IBxeEYKVu7
2f0+tTbf/eToryYh0Ek1yo+gwBHSqkncTO0beCFcFY6r1HDeLCkvbuDwl6iGh+W3
M+hFpnZhEpG1kW9yhCyriIE7pSUax6LZs8M0kUGS4WB0Mw9ePcWt9M0V1YFv07gR
rdtzvpGJj+tAiKIZocOn3qo/d6FR3IvvEjvRqgU1D4EndZa5bXnAZviibRqneh9o
yJQrozG9AOzrZCqCg3Aup0+pLydq4f8Nue6PJBPuMLT/ff6Q85rfPoghKOMwlZPF
P0jFIw6Qr7jQdEyNoNW2DS2LmEHPIkusUqOiDukfA3s/4hFfHqBa1vItGm0PRHlC
f6ixXBRjqmy6VZ2Q6owh+f6q4T3KQqsxpUPaDNboZfrGZ5uIW/xx0iusHXS04mnl
WWAdTwyv9Lq1MJcgow47Ne5zeoufPcVrJi0rdGGF6Md40+ucv+BVCArlRNcOjwn9
AE837xo1GFAepRcWf3XGMYg0hccVRSsU6mkVi6r6R9NVNF23HgyNjPTEgG9ovhX5
chkI0RyrMO99tB2HjFCepRYX61reztxpk3Om+b0o11SyPf3H4OBaN/Spj1bq+YDE
WWP7syGD3QXV8IcSyAG6NGKzrURCpuuRnVNRU2UKH6bkEPPGxUm14NbiFifSDMAo
7aLFmg8s3QuXiktc8Y+tLF5srro8lccDDcIufj3KE5eKYl7F4e8drVhbX5h4JRF2
DDuLdeatTIjCXeejmDJc+/BwzULx8L8ZRKkv5/1PWvi4w9+dWckNzmIUMPnaIBEq
zAuU4zVAmjo+hj+dtwDyZRzi3f3LzEtaH8LBGu3sLC1qJarCn4UB/yfXxNhYEe/M
TwNH/z9cE0Tl4cINWOiWROd0VzvKusUOfAp/XrZaXP13T+HmUDiqcKEydmyKBphb
QKlocwOPXb85Cxvn3F2KYfG3mSkShe+sYxVuSpDm9e/IucKnd/RehaoyHqkAX1zk
oSRda7eB7eBbWLA8e1pNVW0RBcThMBugoSMm8QOxLmpw4UCgq/b3MfjZ9rDWoB5K
fhGe8Ch6gAnhatRNHbslxdOe3eQ3ate4gDx35NKPYJwopQev2rGqLN8ptjkepxIN
IVOrml9o/WaJry5bN75v38+CupzVg9jcpZpjX8hQqRN0Y7VS1nJ98T1QVdLjVLN5
SjTZjk7zjQCW+11wo1xz34I9+C4F8t2W97UU6SBSrpNzlRUzssEJICnvt5HPstZV
s6fkHSYNz79lSRT9MpQzQndn3hBiXMIfo8R0692PYm6yQeYcPArlE6k7MaCAHWis
+7H0DzWDoOluKWuQL2VLyfmrLj1lXQaISxNtrTPFFckDRFGWr4SEBw9wTaPaAbI1
7Ms5aI0mQ7c1OouocqxTNz6UZOoeXy3pKKVmHsO0vG4OLTWlief3joVQJlnSvwE8
PnLgUVRLug0J9ib+cZVjG0xd5dfgDmCYwNLG2v2pjgR0tXuolLqCixoCpv2GFAbF
ch3JNJXB3M6t7KtTLotD6F0Jnp/0qCXs+EVw9dSxw3YW/2dNsmE6rX7nNdkCtheR
gES/rAJvQaLwOAyslvLIELwyEIKXcOqcnFAbkhMwvn9aE+x7JCwG7vVhOHfoPRkL
8Wwoa9zHPGUBlPe6xVm1bhLW9I8DMnU62aNKBZsLnRMa06cPgy3mDHkaaRKpwQVg
dgkdVagrNlLapmKODTVii4CRFhH5IB4fkNifmCaJBJIhvhancuoYgQcJIL7UzAxX
6J4proSiELjK/9KZaDqyzGnV5+Ck1Raz6PTqk8ZF79AtsYCRFf1frOAs7UtcBXGs
VXEp6ysECcP5W4Sc3+n6ofjqgAcbNMBRUNJvKHoFWgfhTvH75paQI6g/OKPXmQcx
NC049UAXr1sBSWI3cjAQfbVO0waEwAyDmozcgDt9imzaAGexy1GAlk0YcKtwyvS+
7PzlFaoUo9FoBbAdelAU+8GiWUmKOpkE5rT9hH4cbKlG1DZry0pScgM6HW5L9lRW
cVkE8HL1fz+DASdLMGsOXNI3OO9gSplc749luz8EeiMlJ1/axLASXUvlPP/OkYqQ
DRMlCwECB3IfV583SHyCEcIRqKFQbgouBLPeMNfcfRDAHPnca2y/flgdxPtBgRSd
lX7Sf6tHl4Hz/m6yYMqb8LjokpJYW4BQi5C3AR3yaicECNA6T9Cexx//Wy8Otvof
PgZUtWMZrmzYCTupMNjukNo79MiXngSR95SbQhxQ2C0D883kh3ZJaTk0q7/WnWo9
hSdaWn6FlGG2mGKvAmQRQ/qur8pCKK/sOv8I7PfuT6kHy3l/sW94Xrb/ICqr0Diw
yqYW6C5Ca7GvA8eDVxPvA9LHDyyh7hMEgBsziko5ybWquLXa0mIVaa7OV3m8FgAD
dIDFPebBrjzX4J4ibhFgLxOODYkoZ0FuaLLtyR4mUW3ieunWXG2JeI7yusS+Y1fR
RC6qE8w4T0qiQ3InpzjwUkDNyM3nUCkEOBvKN+h0v7pGizLbOGgeKig0ZNzGdxTb
yW+NoNrkvA4lpcEHOAEahEarq70iFMtuLzo2Ycy6J7dqf+FSfvQSUoY6EUosyxD3
r6CqZH60y/kxnP7YnTYHylVBQQvcfvn0GC9pn48mPrYXWhLz9enPa1Ds5oo4Z6pw
CezlpmvvNq9M2OKGEQGYf9y9A702Qopq3jww55DbmOP1a1qcogBwAB+whup31+Wn
XZ6XSopPr/XQUFuEQ+7XBhg7Ex8q+CReUiuUxpmCOmq2U7LbB726Zvo9hC20rBFz
JsAzIdqyOzvbWyWVLHTVm/yEwq/lJJMUXugdX5Lle08eBz/OB7QujiCusnrb97ct
3/8uCkF2w6yXD+PtIQPALY/4DkzVxSg+C7tGF1uyakQHq/7fQO5xN7b+HL9pG42G
21e7j/8qv0DJKP92vWtDWBfzMdKqvAY0f1mS9gP/USh+KRO4In/RWOE3AI2dwpJ0
CLtRS99nPQz36ckoXXmHIYtGa6KrZId0nLVcmBePz56qtc4CW6y2+S8CDHlgM8R0
8r4GSl52PrPPX3Dhx0OQPwTDyMwaI4GPV20OImC+dNnQzKLVQVvXO0Q44taxKQut
OwNBDYqVNEVZKMkgc5yRjMJX588qAWNAc5mBXBc4Jj/HwJdmixhScsduX/y2AwXj
Wo/8wCz5k3/BN10zth8KRfPKrK5DX4RREErFT44ph+RCb7dI6XQyQJ2wqR56SIs5
ZPqGLf6yy6gpW9zMshVlKGchZwN4MP1lvv7Wph9Byp9wnCKAZ16LBpZVa152XT4p
FYgI/+9OZRumxvvArS57TC0i7Mgr8/ZHw69e8M/vUBYgpIm18qP9v+IAVdOBem+A
Y9KYjD0EQUTmhwOPigrAWXMgvGjsoM4EUQQFDMRREAGuGLmQpE7werKZB+ok8GBN
nOc5Z+MFQ8nFpYBH4I6zCun3SvbjvLC3vc8eoPWGKNm4MDaE0cRhKTqSffqB8lK8
Wp2P1+2DAxjWCIo5eqvguRL78eaHAVdwAlhRVAYkJG0qJBiCIjBbKDI8gRbD3vFZ
XxVSHdZdUlV5TxRclfLGQ1VEC/uh2eCJF2AZwE6MwbwHBfFN/Cd8wDTjFbiTNWYc
H/zcIOWCvKWomRoAd4kLVwk0in21sIYvfOXHlxJQOny9pBZivPURRCh7oQp4cgjM
qspizV0QqTVosc16JEJMPx0G+YoOjHjzlEC8MCSlV3nMXU6VEdu3NyyxsW7QfgwQ
3fLXq6wogq/oR3QEqiiysD3RtWkYz67MxKOhvkQtQbX2u2yoBcxdb0R90HrCsmTP
eNLn1Eioj3rjWAcsmbZqgZTZAO3tya3VnrWyDfMP4pl05z2d1JYh6cRl/jW2Nz5P
X4DhS9w412B+0ygDV4A7q1uZtm1obwDhxz5u8D5pWVVk2SiCB+JFP6tu7ERTuVFU
MuHGXxFXsfPAKdHDJF2QJSmDQM5HV3+CKE2DdLwcVQ8PTyZNnuRpGkfnGvxwshx8
Vi/tMrWvj+OCQ+LZ8gGlPPKKTCQgfNaOrLDZrTtnwiDqV7GPeIzWLJFVcVCFFg9m
GU0VVlZoN+SYcz2YRxchGZhhup4IMMO+BSAScqAm73NJkfUbWujc3Scb+4mBEtoJ
uuc5h4yb6VD1i761nff1Oo1Yn2iR6xJ+Fj+auMeyDuTE5fpjkaKIFxjyoh5lN+xK
/yyxWJhoxel0z+UuEfcMIm8I27cQil1Unzy5gMCX3t4C2yTiMOinkXz5rUwuepZz
+5XIaC5tgXVtdZmuYyBaKVO2205umsdxVnCj8pnVyli2F5bCq8bjNEIbsEoDd/uo
M02cZQrVWS6WaG5uqyasvcdi1nY7G/BYWbL2lExJ9qFZcTLSe3JBSmSse9VKSFEc
WQqW5kax38bRc3Wi5Jx25u3X5b822q7IPhVO8EfPLTcMi9xQtKO+mhCcgmWuG9nx
Gw3Qts2CulX7YnUT/1b+gzdky0Qzr6txpP5no7ZNXxhnxOtW6VNWopKU7gJ020b+
pJx9+TB8CuZG6RT7YOJzgHas3T8L1S6HQb4NVOj6Cgyj3pNUw/FqxzJczC5g7Ydt
RL9YR7+NpFkFP+xjZYIJI3T1LhPoH1B65b0QF1NyuFx0jJRJxWZy8gA5SiVR0OSd
lXpBciFl6izjvtlqUdRi4XTScZVoW6uqaBtZ0ZRKfgnPHoskzESfmf4RwkCt1w3i
3Pt6eLrNXfLivTF6hOOcdErSSrrdLFqVCzHKg64FMfcI4/Ffzu4yJfyESnqnfSf1
PPaqhrwgLfZezER9y86XB7l/ssVJGoAm1Rc55GMelwrZBcdZ4UN7ptUSKcmb58pT
g1bZu3ZqNBbol4+uh5l7e5XhYFMy9Q7vcaZtnPFd2KyillxKBFjgZVihNmn0dQY8
qsyOu0nkflr2TlLqqq4201Y1gGOcXNXGdAGz175LtQ/QUTlU98asB9eTITaUkxDy
AcMcnSkmN63FoL9RF9lcsnJa+2BRVz+5edcKp1igdYEH94Z1qMyMCfjM7l76Vdb8
Tvi4WaIpT3QS0aq0PA6YHcyWsZHWL7Gq5tiDd0j1SsSjsJ0lsAjXjWcpHRc2WX1R
OAo8v17ovEAg475kp9Ui3udhznZRWa2YIf4NhXBv9bjzby0TlMeAlYJH5+lfDpUP
dYtLOh1/VqDKCGdSUKJWvB3/cRs2XY0iyBE7UOMtWaYkDFbBV1qxJe1W1EPmsCd4
XIW6emv6ONpbq3lOmiXwUXTwR8MlvnXrU14NZaXStke3ytOmV43aKzl+9LyoMOYO
C8UVn9sCfYfT+0jU7nG/lcmzWAm8dwocyk0ojYiYSieVx/R0rsz+CczPD7rSjp2N
h39EmZwGjUaiAHoQ3odcpUm4GiM8cg9eKtQUG0dm+kw+jsF63QGlGElKUNV6UUry
bllRuI5TP8WuWUfTvyISXQZGndONzKJocnTe3b4k0nz5cNVOULB8cdiyZdRHyDrZ
BPTUZMq+GL3bApePN1jYAHqTIUxMDWbcC4/AMvyMGhNbFW1Qxu/6F1un0XXkJZoV
DqIF07tQER3pqESnqnB80zUZu3Obx90q23UYAx0vd5yn57Y19IknIvirlIHlSI2H
+dZf+43hKz2dI07SG/d1uNfV9cxayk+C5gHtwV4DlKXeAT2zFbqnwZnfKSBIMw4R
PsKh7xrhdpPR8TLUj7MEd21XOt6v3C3+VubLZlGbvrJLljuNj+W71M+Ojfgsxco0
6BBmKiuKG6BtmIEjwT4LU1VYN4vm7WY0e0Lbp65srB3r0qI77qgowWPRCWFHh0E8
aft1aXGl++C4wIyJV1mbi3LFfl53+QGqOJAWb8rA879cKfsNpLNN9dH0gSraaY/A
WwIyVFdoWcFNgSMOdcuQ1ruVq8VaA+SRzBDRRLH3edaJwhvSqErsGZU5JHXWumWR
PnWKo5Hm5WHxcvw3aNGu7ueTLX/TiQ3wV9GeuM0AX9SeRKr8jD5I37zPlnZtz0uy
0tju7Ux/bCkkdjrK7nwyC3kGj3hzsrU1PrlzSnb5i7QT0NmKve/XGIBSS/2CHGVC
jHrbic37I03O0j3hGgIK2Euijq/sp0DplEIDydg3mX5dPiWNR6pEYrvckBGJ47iV
0Ii/dtIIdu6mfMUKUWD0kV6gBnq1CZmMLbkpWY5qAEDnBK3BZ9zSAqlFnJ5zL9WF
A87D8fhHRM3wTxdUmubl+5+zdRBMfGY1t5rP9pvS2XV8ggGR2MFRNPhp1nz9ER3e
RgvYGs4vpLjsUIr+Jge3Jvs2rIa+s0+z8V+bdsWrcXtVGHy/19awNMpebPONwP4c
RB4KhsR2g373TGsZM3x3i8fezWfXUjUocm9KH7FTqYxY07TkyIkQQjqmaEE74tPX
bU5GplYaCDPYu1Axq9Q3MGUPRticKBFfALmVBtGlua0bYvPYZoIOJzAfgz/Vgf0E
3ASY2ISnU0wDvXHfFKNhoyocLjYu/rj7Ljtea6E1fqRuGvgaHKorHUMEJshh+kTX
2ZaCYvIhwEimPj3tVZIXfjnp2O86w6IddRPTh5ANsjelqrRF4bvstI2Y9owO9ZpC
BPFqagOZiDpWz+UQEsbDNRsR1/2KB0ZVzVkbYN6oIpoeMwYZ1j8tZ23Fjitzicv4
aDCeodbgpvCbbg9EHEOlcbh58+0qzQbuELIXeWM+6+4hi2C+hrGNbYbQXT8F9ohk
gml39jM3qxzMvjWhGSVfsidLXNEe2G05BIAXJWMleVuEkg4bA9dJTSINmd84ontO
PUnY33V/NS0PhGFuhO7jYy8pEIhWuNy6C30xV9PgGE8vN2/Iddk2QhxJgcHWSQFI
y4hoCfOUNpR8QWi2MBKR2ztONBXCjOcRyiK4cYJGTMIfr+1tNsAaW4qoGhtW/Beu
z6/ptG/YBeWYaIl3cENfFhZYtoSDxFy28sb8/iqCGV/QOIaGBSTg/CxHn3xNkibG
uvUMIb2q0TTNdkfwp6c8uw105POJvYEeinrmlhPZirnqYK6iyi7VlsvWZTBgNmfq
TlscbP1gHmK2jryliprbawtDVHnKpk3mf6H3HFYDq3CxAMF/q6hTfxjXGaZtkxja
ODK7kiE9s1xmjsmku9Uxjjcvq7xAxA2bXTyNU9Iqw7YP4sS42g7301mCFNmmgY+E
adoYgE0NgoqdREYGgbLUpQNJgCL9y3BbaLOy7JQKb8ZiZcsxKmOB90I3hdgnU8rO
mYvXe/q64VM3WBP9ORmKZTR8K1wgDf3NHkTXlNvC2YGc9op0SeHtSAYSxML4LhLT
Ix4qk37l8V/yoaDZeL6SnVGb78pZnusXFpVlAtG+/lvLiGpaj51gLssflAUqdMgV
umwPbRgFHwdefclXC9X376+WiicakDKWfDrF8wodlPYxA/v9txDAUTs2cGtduEJL
1UlqfsQNqWc+XFoGWJTyk9XBrvoHtkq9KIJUBg1HTxZPbn5jQrfYDUcUE9IKpbOQ
PRbL0YZXaf4jWunU3nCOFePj1J42xbisFCg0F4Mgsm4XolzB36hD+jB+mWjoasCN
9xUjEzQTlv8WGm4mWAHjzcXdA1VTrnZOgCwjc5S3aGBNJRf/0jxfOKZHkokw418D
o+Zq/0YFkn+mxKrhbQ+hZHGY9LDmvCVplecBW2VAy2BQZoQ1H15D7qOd1a408YlP
VZVUFPnFuzKDuRMdWCaqKRky3CbJl9cP4JHtxFwq3CLLSMIPYHDSQ9Gz94LbjxYF
fuPQEgxjEjNZyte9R5Q6Z93yR8zfW9yyMv8+G1Nb9CK6leGnyUTkWKgUpI/RuCfE
GSGPa0jOw8LjVub48aozxy2ZUuS9wjIbF54Znxx6tpTPaiS896vDrdqt362rjjDX
DTFXNV6VxyYW5vTDzlp9VMfdEY2M0qEtAStE8ZyKIRVNzhl80AuOD3cTpPaZ+OtF
Y3aLmMzVot2wKkhy0DcOdakLusbMaqwKKvIjBYpjNgT8620JXKftyEVXJqFdLHqE
fU+PmJ/iBC1jZ+OGyRHV9jfSTjGAgn/moXcGNiO1AvCLiIgS2wnPLqg12mrtIbR0
c7aq3BCL4UNEtSr4FFNWiFIR1WmozdHTBTE/vm8+6ORucyAiJmMI8YE4/OOkytOr
MmNS+lnk+SelFn5RzRxYBl2cSLQAJKoZM0F1auDbSAXtbNoCnaeKq42RbhdnPMda
T9HdFjhhIc0RP5tnriN8+59B0harPpxi+bShc46oyzBRTnI8qmxRTrIdlUE31Xyk
FRFOLrg3damu/EL2PpsIvb/5ejDQQjZ8ZRa5TRjQKreo7o5xrZjkzFDK1b0Fl130
ItP1Gl3iA+JJZdpitWTJEs1xCER6ZZKjlMspQvPBISVB+/q/zxrsUifn2kc+C4eW
Qw6dgqPX8oYhJXtOkt8MaA+0dz9OHACECZjyPl3LOfr7wZZTgNU1jQI/tYpuWmw7
1T5FdfHi8skmk2NJeDiqxoN/SdMsFA21UDHgXy20hmbV5DKsFrXEPGxmtdzXIPNU
qCaA7J9ZZcR0rtB9nkZh00VAl8L6/Mw+GeVPoPcyB1/8BuBqsC7G47Nrxe5B74NB
e3nQdfkbENi/yVN0/Muw7HdUnFs5umGIyp3XAex7uURy+3vWkLn2wbvsqUrK1LYt
Np6+3jB6ICoPHf0QMSwt9U+3bK2pEdJryMoat0PhMEoCGNZnV2Jm1DU+9o7GRgYH
/Eti/9RxTIMTnwFZI+3y1Tu9JNqq6iukIL+dNqb9qRnmsM+laN6thpfA7R1Hjd9m
sWL/1Nbr46EjX9Qz8+WZp2Ke0arB1qDuyhnLRZmj7Ojwc89zdDIXUA18w9dsaYy/
YNDn/OPpJp2QFyKTt5UXO4UoX8I1wgpv8KWaI8sVncah5d0sM0dz+X9m9Vc0TkSc
uUhERfcmkb6t2AnEJK/KAlDbYNuLalOlzPsnfm28XRez01GJFBe1ypNA1XukABEx
LobhZ10U7SrwQ6+mdlvsexStddKo+e3nDP9srS9FcYqzuS/x2K5mMwLAKnsk/fdp
/jEjiaayk1zH79EZ+FLxD6lxsykga+0iXQ+kn5HbOrfyS2rjTHlL1p9eYIqi8QNx
CgHS3cUbk8Azeu0N+2aIb5enJ6s/Y9VzjPf0Gen72pUEVL4++mnfGxajZ7XMm/Vd
UhjPN6T4Egwjjtdb3Xtu6sMrPLoTPIAYt+ud05zxFr1mNc98A3zFQLTWu50EOzto
dudbMLV76JyUxcwwOpQ1g0bHjP4+raGDQ8N0ZfQWVQB9TkAIU+/pYpZNQiLoDMWj
Xvy/1swjdPbS+31oeTMzk2Cn6CIO+1HqWGA5+Ot3MtNVelfa0EQJdZ05JMqvGSB7
la9cI+NPUT9rHev9p6qwbFPQZxDTPFULq/iHuayirNIvSls8EB8cNm/INQb9Jlkf
agmIuCzb33aGIIhxLEQ4NtFh6cpp6zl8D5Ar2NbZs7CsTCk0gobzwD9D+ml7QmlG
XC4ud4OCiTNwHQ8AkDAC207UOLlwzInqOjDG7+Ihjq8llKm3v4qSfPBEDUc9/7wz
+YQnkd4PGJt3pEwiC09A01v85LQKg+55ao6yGz5qnH9zwNJyk97kw+v4/2uT20XJ
q7jcfwYrIRTBtU40qWvF7BjMyICuN21t7ha23d0gXAvZMXtnEIV8kQfEuSs47ID4
H249YBx6g7bjQX75khhBPOGqhSyPlBX9JMsgc0pkOM8BorBB6I9ay/UcQp3xD10c
AaGGJy4jRFen5b7Kq182N617Qw+uFChNrKZ41xgGZ+Z+MLeHrSdzRmYT6LW1ExjG
knbdWBQYWEQwzxsr1q6p3fF3pf0ealsAD1wmmhDAJHI1qnzD2RXnb7uhMU6fCa8p
YtkzDqkBR0juj26gfm5DChC1zcR/fBKaCbVjHJPEydGIVGaY0DIfIQjAhpNYI0QX
Ecaqk4prj8CMX8XY98D76ebVXvqfa/ggDYYmCXCr2V9kwV+7XGsFTZFioIhzya0M
f6OqfGI9kSivtK9Neim7YVGtxFuFPc2TKb3LefxgZsDav+HQhII5Gw3PVgzk1Xad
mPkmugH9sNf0Gp3PxeGy33TG4q0ct6VqInyISjfoL7NKcL7GtvZazcuFHwfKn5z4
w6pZr4ap8ocDI0rh97KTqGjIGwedzM6DhJtIlWjec+nj456hD1Tn/9Pu5NqFO1Kl
IarBxKqIHwkSf4bFDX3lhvdNfIC5O+yaChndPUw63AcnDcksOj/wPQ6uFpdVUzeU
DyQ68n9HUlo7rPa1pJQ2JwgvIqAKXRnHaJK60t/xGVsnAtyD4AVmINcHRTJuMRsq
YatUY/cng5j5L+PZlKdvnsKpJdUhSX0GTCREZOEEhpVnVlM9RLaXa3hp+rQK7kYH
lY1wpfal3nt+nkQrQ64Hk82uWOGWPT1yzlOTaxpF1095eZOAObWW2D2Q7XLsGLRL
v+B6ys9l4TYc6BKBMD5VonbMGHXgolFA05CJOLQ1AHFmMtF36+FtU15zyykwT2rI
kj9fiCd3F0u2SG+Bl0K5NUHhoIZGTWoo7ZAypaurnwhPK5qa5gVA9j4mKqktiHFP
4g7p0r8uE46pj9uc0rrmC3d8sg5YQM2A1m6XbTu1uSYXZsNnUMLwdNr9xJSthfrI
PGBakKZqOEcX+LLeav73SLoGIARzeqtjsjCJKWr+3M16QJxDhP+MpGX6rxJlkgzj
1JGxgSjllqloTnAcjaI6iWSXLIaekfzU45ivjCriz+NG8QHinnYLdW+u6v/+oajb
82+Tm259sBX7LDXrYcLRrNoFBkjHWAC7HdDExRlFI7VI4djXnyUQrmcl42OK40Cg
CX/Bbrne6JzqZsnDkGLKb6czYhJwRLg8qIiT28/kcfz9V5R7UdVGu/z11npCzjl1
mKTuUSHLa4YKQBGPMQwWAkeBAMn9WjcZ9AE38IJsKVjbYGppHhhil9tu+hQXCoSe
Rp/oPS94/YpmAO8ACPFLT1OUGGputu44gaFnm/51xzmt6Rw3xAiCh7qn2TSw8x6o
2ys2WFCaG3h1+5nqbCAfaO3S03B6OK7KsgqBcePNQhQY/GvTZUhpgQ8U133Rf+ta
4S9hjY+MYWHWp7hnt3c112YKDBxpzy66BA9I6rDxXtgdqKgwXBnSJF9bm7mCUPh+
6kAcpyOlWsa4QuJK72TO/a+1fjhxULhc04kPmuk8ZDPWEC09fS4joiLnrCtDQ/Ip
viYwp64+KbwFxGoyN2Gt7WCFI6HIM/v39m311Wki4mI2YLAn42oWNMNk1asdiZVd
0VRP8cYoDD1o2MArBKtOIacqVSbnTuz/jpYU2+7PisaRAqb8EL0IARd1YHiEisxV
dn3mZRO8aDmh8iLX9qHbkMJjDNIVUP0fxAJYkZKaLhj3hnJyv1IgC/H1zMUoPMRV
YRZYbkrQNWFPC41SuliPRMe1q9mq4x2GTq2uUjZt1mlXsIe6yYXFC1VENxv7L56T
EGqLBEsbHTAqXJM14Ktwa2bH77LXRPCZR/Lb7XCr/B09dGY/yXekr7hb2ZCQ6+MV
LB2aC7lNaUZ8SzlddHj1OlRfqOZ0PRr5acf41C5d4AjvFoZG+EGcWau3n/n6jeF3
wQdjdTy3JKASIsYqmo65237AWkWnoqxByqNRLXEkSocuFprzLY6bwgvGewSjHHGF
sN5jD/UKpCXNRalgXhePDSA/28sdbI+A2w+t9M9laPk/k5kTk2WoipXyljGhcc6p
4T6I67nMPjRocf/Xj2czfq8Ea9yRwWhpPsdB4I6rg3kABLAibe0ZBoyhPltUi7/8
YRSeKiPMiiDwoC7t7mt30XY/DVpCEsdhWUSGZEbgDNeK2MelY9gWQUaIGhjyueH7
BLn8lJixmHXpsKHzAYS2LRf3SRwetXte/kQnUA8frcDm5NTOmqy5v9O6/WwI8+ZC
KxkMannlAOTJwdoW/8RxZGrBsRwJwNtd1296KrknlA8S0IS2HbiiSw7LIyQTQam8
7vulL+9PZm52sim3SkgOE0+Pn2HcSpHvJQFsA6JyPb5Wg56zjAw8hFf1JdEhzRPq
FbR8GWPLhLRG1do4Qr2tkRdGscFHBntUH3P1jo8dycMv7/eOpOAqxAvejZmGf5+2
X1JpIgcaBGKZlrURNgeqBeXrbw/9xbbPxTi2LwsyweBHahnNdTmZ7gAI4H3bdDgL
a39O3FlSJr4LgOkRPsMiMXgVJya6lwzodB1p75hOAX1URo34NnqH6uvysEO9NOAL
6RS0ogcF4wGlWd90CLhaSkMGRQEhwem/w21ifo4bhszKcs6F/GKXSFUoJPgAGKfw
5xTQBmCIVFSgdOVmtyyhbSskrBgw5Y8GsvLAqtpm8twMqtu6Aul0lHudeIfifvOx
VjqVWSUSjOXdj8iERLyx/VtWAvkBnaH9z2EZZTk2lgiMo/gs1VnL4nl6HoxmbrnR
LpbVgbafGLH6crUVDfq8knn/5CH+TFEusk3pekTNnoSS8LGEUPKzuUv+yERD0+p4
GZV7ooH4warabAzHk9Sks2+obWfNEUsPD3/cmgocI6jHwVDlYJuNmgcsN7kCRWQu
QpJtlvxwuA8GUvcSx84+H4y/C1PRmcNfE8VLEZBNr065Y+pcg4vLUk/NXcWyvYJl
CE8NASfOCKAxyqbn5PouCfVhLpBaC4CZEEkVsFvWykH0mI+IEptvqsSyuXV/s6Bs
2dRuyWV1Toimj3pVKY77uTgk/FGOobH3HP9pjR+9WT/MdWOsULRWRbEAs5XuuloS
ZWhAiaCxQdGnRVDdZ+ZSpnRnxQuQJXjiI9XLhjSYKrVIXZPodNZKgDIgLSv8uvTu
r645ccgZnpgQIuATZZTuYVdWsLhSO6Jupl7AcboHw3t2aOqkSW/zsoQDM+y23Y3j
WQHtwDYIh8M3YRTLT+d1pDuZiTmwvq22sOCvFIjh06lgzpQtiTneJ8V0eWUYceSe
ZjcxDonX9/eUWrb3wnkBeVb8Fb0dO804os6KON26ivf/jLw7crOooxaUKnhAnr6Q
QRIwRp4nMFGV1FgheS2X+bbb7ltkii0Mqp0G4/iIayN4kQmGiCwR+KmmgIRbuKNJ
LKTIUdnctpfUJPBgzZCerbOhG+vdChvafgW81nhKN6tY7BqMf0TiCtjcRIXuIUyR
T9v/ZUfG+aI+0MHm0J4CctDCqZQ0HW0Oj/rrhzmTWcFj5f5kxafKwkV5IKUb1cB8
QgPjaIXdA0QJCxMv20HABvL2dIeOIhU9DYR3eY4hX3WpcgjZPITtlcPAvWRzVBa8
u9fNbyHoGCbKHAfWf6es9DaH5nOHOHvP5ALtx+VbRkuHOCmDEAIoLKMUdUH4ZzjT
1MFBQyNavaqSjR0ERc4BstZ/VzVCE3lvhlGeUQUle0XJmX2+sVfJnI+0D1lBEyKS
InxpZNUcIdaljuqS5IvPKNUUeYib2mEWlYV0+6Ur7pX2dBoBxRUigZt3EWqeFNMD
T2BAz5oGCv2vyWigoyYOqHFTc6MAQC3Syz15wgpm3xjxgeXd26w89oI8jApN4pju
NhFG+mBUHyt7FPlgvLDb4gpnkug2AhSfoxPBENhOgGaofLE2POql3Tp6zzJVJPoy
H95l+A0wC5/pPBJeAvVMfEm+yh0AXHxxc1XzXJfSnC7mIpNjdlJ74BRgFqhLbcoa
EBG4Z28ShEBwN67j4+rHB8YqeTTiCREYFpQcDEd2KupTjU20Cx92MriW1wu3NLv0
WNSoB1WEPsMWR1wRAGQg8Oy/+t+rY3khc67rwNp52Sb7klZ248UDEy0/1hsiY4A8
gz2xU2P2AIyrTDYW06AxnhUyI4PM6akMKf2MTr3Qd1sj9dMsGzX6oDKB+0UPOGsv
AnKVqshLw0GgLF/bqwwRaDFqM8ZjFjkp1fOJ9HHFuzh/mq/jb06UkLsTIRA19Aql
oCcs4r56dAKJR1KsUJE+CQehpyf5gdGYjtuhFdpY8ZBJyJZeuvTvx3TRZR1gUbqM
bt9QqvrgJMb2zp1y7i35k6ylz3sXow4PGlIxwMr6lCvKwBJ0YVIH8DeoWDuSp0/s
sSavxst/vHfFqLGn9WQMGGT1buBqgVjzeGxaISpySkR5JQOVXcBRCxo78QqDHmnP
wK0wwj9bx+fLHFccJGm+2Vkb4Hq6kNctpKD4c+CyA3ch930NC41mkyhb3AkvUOeV
yva86UMzVSkpm1F+vWvKqK0xjNcQqtc3InKRJw5sCQcOhiHYes/u49dyI5ya0IvK
h1ePUjLY8QMRat3dYFNMuw4CB+4BxXBCY0OdcNT+xPQHOVSszQW3sWyOKSRIHHlm
ANW128/3gsz2sewWvWhjwGs41BYEY5sq2k8+nf32V/Dzq8s32N36LEqaiIDoedVI
ucFjcXug31OxLgMmafT170+nEMKYNwV26FWy2/tm6nNCSsEnwkiBA0R8XOQkn9Hk
iHNYxiI8fBbdYAUbPvUflss3UrtRIlBbwDmR0CpXQKnUTfmEuMMPwh8RkV+Ln954
vfRlR6sQt9/h8wwdM3Q7Zxd4KeuUyORqkhQGpt6izRGKsnSBkjpsdUqbvT+x5xUV
iprGYOWiHLd3B/EjIZEYPyTkvuNuGXuToiGzcORZtqEnxj+OuiEJ8myYetaRX5FB
iwt9hDU01O+u//VAWYAXcFHZn3iGsawahwRKqJvecCp2lyPzQa4+lOruqJTbiBYz
xEUi48zpNCPAKN38ueNLVxpxTnWsHJ4i4Gh94WVnyRXGOzeUTLtGtCO5ELXKTe45
3nIlHirTr9q/Dw91Ob5XZxcozt96Hov6KAwMpEnnIraBaUqm9rwwwxoMxoKTpDJq
xe28Wvmr4KF/NP3KPgOp3X8dc2TuY6b4PigarUKCP01jXGyvD8nknMtja3bJjgyu
aXzUWq6v4eD8fISRp+dePIvt51CpPwBrT+gcus09Fd3rGUyv99WXU/04xcimqwog
8jwjSCJH3T9Lt10h5zTLTQHThfA4366ygJbxW9bwxGIugLDyF+ekfH5G5x6yK2zr
FNWaE7mlzBBuY/dQZlror/m+GX2+sxa0FfSZ2cAN9oGPvaWyuaXymcydqHliM9mb
bG96gYvRqCPy9H8N1ndDfaK4fkqV43EhHy52LKtVDbInn5KCmZm6yewnfBs/Za1u
omssn+7xSRXSyCezaEQSRRnZ67m5dWtSf6QqZD43JHaMwxj85bMzCc8MQp/ydBLP
XkfobqB6DZQgLJqLce5msu+2ecIUVme1+7l6vHbVeYUPaB4QkPrUwKxizQRJRPnm
vA0s693gLyWYshCubIyVu3K6s8kLzvnvzfNJJTGnAwgOzZn0b3N6VAFoVlRbec9S
N3NfoyuNzM+c50OKIsDuMmZa3oEsuLgthhK1mfdAIljQTeKXtO7Ycw1INpHvxg3q
VgiiE6JTiIEW1wCNu5Tw7AvedNt93BXSwAH8iskefMxf/yIdZa7vc8i/s0pImm2m
wSSVoqvzhLm4/MBn+f3/Wa9/0J5dvnpgk8yHf7a+XxBWJezJZoXLSeXkGNXMshDg
8AC8dEKD3lJZz1hHiyumju085cMJKDyIBKvNWjNz7k8iyHPiIwN3wWPfQ2nA86+2
8koIYKqpgU9A46p+PUs89fj44vvgRqa2o3O8Ga/woQzRcvCX7LDCQUx247uUovgd
TKNlVB+zCZV5COrTjsElQccXrTM+zCl25EBZTGfDUnFNXTPeUgQ7/b4GwcDZBBsY
U7VAX6FamocSKiIt7HFPdVhIQlkwf27JkCn/UFQiyTBdYL7AFNRqPiKT9UKWoSm/
mmM5mf2yS6/BTC6CmtPbhaRImCL2AjbbST1O0a5/ssZhrfbgDxbSaQx7Qcmb6LFc
yMMyXFpSKN323TbR4eVkAHA4h8JT4M3bdPvbo99x2WJNAxVyPRT8ZKXeTXbb8NoC
M1RXuFxvYGWZUOQ/V97Z30cgInfddzKgnreFxhWdbUckgVBnFd8Ni4pG2LiEo8qT
dSINHUrSaHPMkxX3p5ycmS5+pmrc/dEdQAVJzp68Lowhx8SozLA2O/S4yKTMv2Bc
OKG+p4O0+pgxtnwggSdb9EQmVwsNNE6SUiUVN/RwWVceoecZ6C0OHw+MVod44Cg7
J3Y5kLOYgnh7EbxkIU77a8rb+hmVpuokP50xinEToBbdB3PWQAJD302tLiyNMjuF
8AO55ijPCgP0W/t0scj94vfgrd0vEcU85fzUBbWyBhnL1RMQX7pZl93bUvTs53i/
nL6h5Ni+/8Ljw6BWBEgluvdhDbMvkMKFEWPeCmpNJMrJQxFhRtmTS2Fb/LnsNVqU
uM8YyD5loVny6ZxUDK2QEXLQ0O/cpnwLhgWGbEtB3q2B7j/tMqbj/TGLrKydFIBA
U9WyWXktqlyPnbyPHi+ZriEhw9WrrYULiLA/zHeZcCOLoatk4ZcfZ4EMz3azc2f9
9M/J+CAWGBtb+Jwvy+/QavHJDSYdq9bVrqa23iqpELsl8uJkohQ88K4jdxz2Nohx
8yR7ssGR0IUhMwTHYV+uLdQ260x0tXljCAPfyAW5LGMXT6aeGtZfweKTO2LSCqL1
De1GIMsWFdPp5mgiPBK89EQEekxPtdp2PnKlfPWbDuEHTuDHLekT6ZYC4XFw0PMh
R3lnDZIMMykuA/dk9PKxYxJnquoxvw9YFK67PdI+RwfK2n3AvVVsb708zim6nyn5
m3eZhT+aEIwXknqSmW8gCo5B4n8Nq5X/E319EqaqBIH2SIZz94z1CPh5nJptIU6V
oEnn2eZxRIkJe5EhPUSWVKQuRZV6L4IQzTe3An4kZP16/wZwn3ij+K69Wa1izrEV
r3XN1586ddsSW+P/8utUydyq0MSyv+uFq9fAsn3PeGrzO2M52iGGii2zk8OeMITF
r/h5Lz1U/WzhjpEqp0j+z9LJF+6yMV7GdKJqOCCIekUs+4rwdaZlQM38qmmeOSuv
tqYDOqOP+nGloEydFRXq1lDqVWCArxdBTFZnoCtO4hy/mFVV6zpd+lpqU+oVeAMc
8ro4moOwCkFESGbtf2YgigAYuFoHUOuZ5lgWx3xSz9A9HfKPmvdhf5y5JR3PjuR0
0zJw52bqQBWRSQyA/XJoMKaTUsJwwicX2kQHlTkl0EHVgVYbQcD4GrQp9oRiru5i
n+6/KJhvc6/k+7VlEFijXmI7Md9d7WrjEs33a+l31Uhj3psnhjFuwDCJRuvQxlc4
XXOP2EXbItX8pTtHcOZ6qVH5ZyFY72wLAq15/yYwZKVavoPWfY+0uO668GLcCAtK
5hf+I5OlaLMUAQlNJ6JBh4MKzjA+WerLiWPAZxEOPLZtz1jwHw9fOh7j4jVaiJij
s1XqTwrwXe90QnRTLzmMo3rGH35KMoo23ZKz9ctcTRHRSNO43yG/x1OvQSk2Fj8Q
qm8Dk20i1O4tQHUc+nVMpE0NL4jhtKv2nFLQ+Hc4iCqsYqMARLWmnaA+VfRdzsUE
437dZ706gCAOOLJvzu4NJvV8gwmmB1mtz9Q9SxI0v0bELYJ/37tC9qrtaF2jFn5c
hqyTA4T2bjE8b/k4gJ8zVk7BuuypB6QNsIpa9zQb2c+GtRe2NKzrAHG/1Ez5tTg1
afu8EYPvfNXWKiSzl+EPuCbXPPsks/3KvEzETRKoiFSbv2qmTRuj3x3iDyITBttM
2qtkR5NTsbZm/6P4jP+3m6BAVofevPqRUxrSkxYqVq0n80iUkwoacfz6kFOv8MJF
mW3p2Jz/bZI9xIjsUsoPQpkmomKBxQPEAyctJeV8KbeCOqA5LQK4C8RgNzLK2RHo
J0OvmrT1mH2Y2OXTVTxqOz28GlcdrbZBeSvfKfov3PECm5TffpvhCSkC6YEaOllO
vJqeDlIXryTCTjK7Wa80TY6v+wIz2QkbxVTcIByAFG876VKnSj46u1LMaztxDzhP
QHFbQ3zP33Yj+8A9SoUukbA8tsB+l1iEZXG8wQmHF4x0OIPDWA7jyAHr8hkUruYL
SzeR6xgEe6JOdAtdRfFuvIR0hQNQVfI2NmuPm9hItTLw9vChf0yoyJcfWbT9wngD
KsJIyxFYhjiBvyrIFmi1XZehpBHgv3rF05u2Qx6LS8dmtwP57p+Ly5NM01HDS/Zq
hKQdrlu9/wmthqYmZD4/+414VY3OGrw/OfQD9oBz9siiPJlDq4yp8NxCuOrRkUNg
E+EBafc56UvYPldIJg7wLcqHeJguNCRCGT03c2S91MmTLTi/7eA+SJaNrsCGKlT7
TRSb7K8m4tu+e6uhnKmgpcKZ1iESBEJcaVvw4aN9N1gpR0UK5LFhmYhV015CN+Pm
L1LfpaNqSeH9wkiL/tz4WfYXZ3gCi2ld/d7/XcuTobh0T210R7e5T2ijYLD/8hcY
Wczr+0oEWSesAWZEvoBBKdHF8ghiel7RDfoLR5ZOg8Lh3mxbXuVFSdYWpq9wgtSD
Eaxu/nXRttVnsYKmg5DuEcq2RVDZnkPf8ys2AjStk06qY/nVmNO2Th9CqZwit7KT
l6gOBMa8bJkkqJO3g3S6yo038rfkaicZUkOvrkKMlvOF1qFTx+1ZS27Rhgix04Tp
GwrNk92eF5/4LPiH7UWpmNyhohFQefJteslOAoD3Qu1NJ6mC7bmBDKsjn9QA4Otb
mkAI6ByEQ368N2+n/bwZizGAsRRohNVznQBRhB9Mti9f7P7WajX7F8d4GQBKTKya
YL9TIdFqpAxAeMC7vB5gscTHkco4bm3yBnXWLs59k7lDZQZxrIpnmOrH5DFzyJ7S
6KuCwM8l82qwQTGZ4Wx0XR3GoEvCyk0Iqf4zslEKpAsvhe9UXYezvXbypV5AbMer
pCHeyw327xhJedkCphkdHroR+JL/n8+sf76SSklpCPnQ5p5VxYl1qVUKa0r7d2EO
ysct81xX+cMDH/14aY+IhzJ5Zlgfj1HSwxXgj/ExnnC0xO3o1EmbZOmGwzsvlQVf
YHCIaMKnbsRI8N1MDDfpba/AOl965MM8XGKZhM5OZGyu5UUknoVAjJazq6JRM/bE
eDGHWyw356c4iPra+liPGb9nTDwUPsWsWZBhHdgF8kFMcPtaoPZVrCRYgstEVP04
4POXOmDsxa98MohcK84bPDNLh0nLX3qfTEnsL3H70H08gU29w5wviY2MfvSKMqEf
VPGGn5dvH1U1NksaFfyr0N7eIy9ydiI/U7PsKryvy4+JkeDhLGgMIRUbMGkHERDo
yXrkbhxRAOYX7OwTH7MfIRkiNiJCnT+fCVCidoseUcgzewI5ByuNjCEIsv+O5Mh+
m5/QbWKXSKDpyFoPodLCjg663R6fT+KkeBTGxubQMadouUz9L7DIuxr3BuAB7AmC
82hzlVuFN9VC5vfLwsSnwk46GX0w9tUxcuTMda12Pt9ZB/tru3DleK3KRYIJjXqt
YlVlyuNI6MGU906ihBlXnGOGc/OhrVVpn362WjD5+gCQB4/vdUBZHR+ufVAsWMp0
M6ejuicp0YfSlZ7CcK3QM8WMz4yYNgl+DaMPxrMrsyMQ+HARJrdBAV1C5OCmIDUB
2e6oZMbQ/WcQNfYIFSRigIRPtfnhpSaV/W8lNHuNzlHYQhu+Dek95NPkm5PG/cif
lA/fQtJXIT+x/hs3pUlUcpN6vtLd8dWgH1HJaHEAvARThhQxiCAYLqh15RL5q6RB
2dUjMAP6Bcq1gNjq70SDp3yVpNOGNBBE/ho9+wv9m8kPD2tPUZrVNLsCsaf4Ho0G
dUiUy15mJjAtfTel0vBAxBKgwVg0HQIleOtTEpTPfjL64augToQ6Qctg8bL1p1Sn
TE2cHY5JS9Cfh2tG+eq9pRVlldEz6nKhNmuGtTpjtnVMeTm/cmSgizXSFFkxAZtL
aRUCHhbxQ0n2bup9qFVWruVQZX6ukjQEZ9oYy3XsUGUtYfOUaDATGc/quWXZywRa
ZCWzlQXcBhm1AF6Wfp3UVpCEKF6VPRWtqzXhfYA+2Mwcr2etotee2kIG0z2XFaa1
iq4D8aj/ziUdPTl+fZS4CdGrdaIKtHQ/x6CSgSb18r/0hnWUCtUCKjJmvvjZnjDQ
CwlmQCdXM4vOI1RVAhkcUbuVa4KEaaYWnwbC9ewA/PMkdomAKZ2Q1uhNwDdwkhAc
s7cM3dxMxQo/mh4QntL9PFOrlw4FwNUHVbLexlGNAmK56pdAJxbTCbeE/oB2rXQu
DrSo72+xkH19rs9Q6FF+QSG60CUELiMwfZL0GD3nh2WC5umQGX3YYhmYHwR+C9xZ
7o7CYTDFHw9UYvtbHaV7leJl3exr6NxxwpFVkvfxj95B9upIThv6Mj78JUKBjYg4
ULPMKpnRgIsFmlNgf1xmXswQ63cGxpwI+YB8JTTnfP62d5W27RFYT66e52lpyazS
qwvOsJ7jrfGlKU3NSIpGb9l8gZ/e3bhMpLRMyH5QcFNXU0kT4XsIGGqrgrBdS3Z5
ZPQDWq8cJSs86pZT/McCi1JM1+FBrKnK5xylgzZLk8WW1bJcTH0AY9fzivZ7enri
O2nZAqYJ09n0AV2LcBgsBateU5jP2JMQjSYFCdqurhoKvx1lhszxhIFKpYDyMXdn
/sQsihQQRY0keRC3UfidfCzn7QwgSVTemPacVgrJx/CMsRlAfPNRA4piosc1dRZq
P2DhBtUWP3g/nw9UCjEIPrWGysJjZWV0Ze5XEBHv8jBA8mKwaevfSzl/wCI8xZxf
KP8seOaMTObi12HTBxhJuSgoVddDTKXLRtIQveesGl+0Sz7Yvc7AFWeNhjzGy66p
kHgGTkoII0xvsd0p9F4U0FM4tiOB9Lxd/h45kjb+6i5UkBwfk+H+Qn9RSnLfGG1z
bOS6O1iNETqsl9u7gIFZrsmefzZGVZ8h1z1KHfm7vhYypKZ4HascBmjmbaiYCyrX
xT55foawyAG8dEZd/haFOrKv9UFm3vqOFT4L+YmpjcEPHTo+8GTSsqNFmcBMeI0T
dW/4wwuYMAUIZ2vFBBx5vBYa9Xxw165a0pH91xnujnjK5C1BD/hckXGR76VJoZfd
M1oYlxR7WVD7ygHHqPmvW/L9jHhQde6xK9U/UEnUB4u/Qc2w80piB0TGqWheaEQk
v8VWmXOd4ahhfxebxfGvUfiP3JnhES+pphX2YeHZniFWpQw6PIWZIVXaCkAvKqq/
ZAmkmkXxAlp6u7Jjc7oVgQrRFyCXU7/r86F7VOCFUwOSQykyAB7o9JRiA/famc+W
MWEhkf3ceuBO+I6kEkFUV6VYUInKa1vLW4C9ktnHognlVScKphxvi/+oRNzsv1In
msVAHe8JqAqpSH9jcWtHfO+i89f4Vu327026R8OREfHujwxa1Vg+/VoEktZgq4JZ
c6YWfZ5pn4PHsNFXxVUeBcDgCm8nId3FA+h9WC5CJkNQd6nCdX9eyJ363F6GPIBE
Cn+/YW8xAvoW8dn+13gpKYaO3nP2YPNyoo43VJPC933aD1biYKQAswe5Kc2gHHi/
3nNzIMcIPJaG/9qhflZBxBXNh5MMQ6G4koqM7UA2X0WfsM0pyo0O58kUoRnFnKWD
SYdHhpbYpOScEzFU5l6Oxi9V6xFsOMFrBAEchAMcUtSxrchogCY6tb1Cn7qA7Wut
XAjxzxVg+ycrau6fncnSk53aP3f3c5PyuzCFgPyPWLMQKQiu65X83R8of1sJjBww
ro6yDpXsUSxtByL4tRJQlESXAua4FViEq9Y3eDwlNkrQcdPDmReRleviGuWvUhl0
klzQ6RuprrSM06I0NR2MOgExYRQz0RzfeYBXjMr46JqXqCQ5x8Cs6IjZLcLVZhUb
AGjBnhF0UvTXgSYDaY+Z4IFgHmRccQepoXbnIpih9Ewk3KoFaE0S0nCXx7GQsc2X
+nzNwiVF9Vq8bnYEg/vkS+p+kVqfQja3QoJKTiN1akJHIyf2NBKlJxjHLr/irpIC
yerqK0aCwKKEVhX8STMTlNOJa4Rn+ILzske5/w9ySroPw/y7BczZlo0Jy/l2JmcD
5NrM0K/jYHcD+KnklTag2rPrnS4r5Oalb7S3q+dYlhsfxKH09OT2wrInD/Rrajg1
qu2MF6s6Efij34nfQOKvut7UnxGqOCrW1uCP7CiGHEdijZkOsHk1Yw4jh+8oDcqp
EPhAITNBhM09ylMKz/Oonx3M1380aHYFhQdJFSjlR+ShYmlzb9qQeZgsoiGDILyh
qjgfpASz2I06s4q4SDc8ianA+jR8D40SnIQd96xR7Fx8ec3MbsFawXkgvAtbbhXn
MA5ouvwoyPttTScjwDHp+qEpe03c9BB03IEaXtMOXpZ1l7cl4U+qiEuufX/N2zCF
IkpDXkQnCeXslVg+iKLEwoy6wJ2F0veSTxo5MjV28xj9gDFuFBCJRxDPLVTHJwkS
+En4oMeRvixkgnP9+56z5MvX50Fl5pxvO1bJqmEY3j7FvzdtBRPs49wnouqjHP+a
v4L7LCRL6WzD7P/BxbF/Bf/FeAIgFUGbaLervt1sRtJvGD+vgHjRI56PMxrjf0IN
BWBQ9i2iEYiJOA8gdiR/zvl1SibVTIEt6DpzX8bMOisYQPNBwHoNxR4m4JJY6An7
uA3VYRkMrKvbNriVfWn8fTKL2rzCAULY6V/i5MPi9l/ED9NRdkz8E6SecxEoGhx/
EsScSyQNYMUVrrP+92MYTrGWQAq0ptrI8LarKb+X1Ry/RY2J3qmNafMCBqzLhfAi
M6G2Ztx1fAyYmxG6+Jvx3U79B2CW6Fi13jzqKHl6Yh4zycIpw1h2Lrv/HM9PpoJT
aldEqJPe9AMTg8sTLuEPObCoiYGtWNsocBBib70QVMpIwrY6gFQ6+wuJheV0BLze
WhaqzsacOpa0nWRYF15WmtTvp7LsrPAM4tdlRPAhrLXr/MT6CJojSKcK0z2OGxK2
xozZpawpNJ2r8xi8Ltj65HlgHngRP1odybjB0xyzW+23Am/+5x1flUNwogPcA01x
nbNeO3mUfzO9U06X+EHrI3KIP6YSNYGRNupv6gErJrZ9OSEMpYXEnOpliyL03Wqc
+Au4po0bQs9J5AXga7jnJ55QbE9PZS7JS3mb2Jk8Bi2Im9vIRE0xpZIXZfcl/q7v
vKREt0JOEWgeCS/BLV37tsnNKmFbpS1/bjbU7defyL8owEPrYbaT/SNUy3ZtpnlP
veHTAbqyer17JNn6HMzyd0yZA9zcHGU3Pn2AtxQ3G3aCqds5fF9lSfmn6lpLXERw
mjs11xeIo1Jk+1eOoH8H/NWzQn7EmNO+mFN1AkdvpOFyaA6ccXavLTptTBmHZU+Q
iyodLXRRUpgEYLHU1K9QUpzb3cXY6P0shnH+xoEaUyP7Qx+Q0arIBCubgsXV8dxu
w7ySYGh2yHipepjwFbV0svRBZoCtuRH+3PM4S3tPqj4bNrrilSSK/LSiOx2ZP3gW
deQ/dD7+WSg9IAhwhilxfYsp9PvX1Byrh1RRRHnr3lhRrV7fuh8aje/F6u6X+wbk
4OK3ZAEZ5mAK+lXuie/UQZ3pnIG48G/wIX2i0X/4EFyMzqhMnAAm/a9dR9cTGp15
RlLvcPdaWBlkNxi7s7TK+CfWqShhQ9Jm3QVRetualn9C7fOnXA5QjhsPO5vWdpBr
GnU1GIf80e4F2f0tDV4fGeiZ5mzvNbHH6+awmMYmHuEwv1+A6l9mB8GjhXW1AcpN
a/XidsuYjYRAiEvPV45qxerZMW3a3BCJT3mDFiBs4eValvQtVkx6/w8ITLG4mcc6
WkD9KDvc8FZsW6dWmCWUgOoR2qBbbq/jnqs42mzzP+Bpr1cFheLro2kIbx+iZYNq
OTWiM0T6GFyL4nfDAPM7IiF4TGiDKNWIdKnHP81+Aty1cNEXV14J9yiKt31qXz6+
ypbgeI/U6ssiN6+y1YEc314fe2NKvtD1GiFambmz4rBP+a3s1/ToggfPrE4z5QWm
wlbFEhhCGHfkTSYdUQ/dUBprqFmhFLG/v5FGolwgLpBJTTnpvUJKIFW96eL31msK
BcsOUXjQs6xhNfKCr0tOhCUOY2udYz9INpcG0kUHYhXgSXeS+cSg2rth8vOS4xto
D5VEXaQvEW5J2WWMEMLoCav/Ki+jowGeZfm9gzWR/BcVcHBNFYs1yWKlj1vh7Agt
5hN+/IQHOQpKtaDQdhRewKid051Lr5Gu16k4eIKlKsanTTBoDmS1zlCDOH2/faCh
9MJUXwbRTsGg/2LHXa25O/Q4TSq6f1DeVM0YMAQbzGTfYeoQ5mIDGfZnXnJ8Pm4Z
Ghpqwxyh0qUbOGNO4SBCpCgmTnSI9qaab/8zgCbWzXYoWbLXU96uAhy6p5xBOZAF
Tt9SNv8IXG27NIvF10oM8EWvzUlhinK/ua4sE6oDRRj17ejB87/9gx6SHQvy9//9
M/TmK9GGbZET2HgIOuNjyFZvlG+TODx5IoHSr74/pdD8/v3ufLTEa7jG5DMgcD5S
m4QCu1xnW0/ATP5dRHDH7bUG4SjkkMZTThUO1+2/i6xYCW02rk02R+44L4c0SQ67
h6aMYSOhzxL4r2LrPh+0JlCAY0tQ2rjuKjnN6It1OskniLSNPw429vz5PM1id5ft
Qj3A91nCwpkWHFIMQrgsoehsCNEXnVR5x1l1GLaWbfxZp4jZgabna7hgYJMYvls9
mRvv3QeIW3PmfRmlCk8/HqXBq0Phu4kQJz5+bGjTK2Bkkd616RAbAwD3x0m8su6K
NfD6Noxvj/AVGgNEeDqYn2cVvPM0LZcX5wUnT3DqX47+9yiOIAWhX5cL8d4TMqya
Y9a6XHtSOFd4cFmWOGwsewh+/rH/Hh+1YZWFhOtQlso4LaUghAYeGuHobJibgHbX
41DplsjZjlweOKwVrNedrS9XM1kiE7zdyXMZ9qx7RZAY36PhWdokMUcUXT+CEtDc
fSGFvFKs7kc63yzY6oBSxgWGDipsNIbE6EXdu4MEQaH0TFI+nQYxFKMfAhmS0JCh
hz/uytx9qwbdeAZBLEWWQvnCS8CYPjQyWtC0KWtBUKd4zB9uf2IOy2d1wSvxDcoQ
zOeQP9svJgGf5LlsS7Mt8XEg+F2+Cdjw6aDedptfJfQuIENKIWRGPbBY3V+xunld
Ercg2piwHdPstvEICWP/F1XE7f7rvudR+5s+8zmuWgOdE6Cj645P6SZjLytPO5Tl
jvvAzYDRWBnlUhu6V046hNqGjsrxBBVnM7oew1QKtQ8+nz0oW1L8wDl0fg1b1YAW
aG5noRl22DI2k6nri/VJiPLSL6DDGid1vGHHDWgNAdo+GK0+oiI60taeONlc6eyD
j3PdkXqTHQowRIZZ920VEqv+fRdZQVNRQ6bj7/eeRL9IYVmMliXsSJjrwZ0ihoiY
CO9yj0MugY1HrebCKDgNP4QGU2vIDJk0v7nag05HcdMTaJonhmi6+qg3erXtzNmA
kSZj9C36/IlSuk/5JJg4xmElTtytIfZbAApmgMixeQtazVIaLiUx+C1iuSfN65+k
pMYk+aSqIZcJRQ+5jf/gSvDarq01gFaK8l3QxHKdf8sLgXHaJzRgfo+2Wfw34Vxz
L+zrcVg3th8yQVsUMRnK1BOafp2mxgnWR7ypl3ssC5/CvoL4z0HYy5tekF9Ry6Ba
Ai7SV4BkxnwOg3KGfvGrsLSgzC7YP1QTiHoga5VG4ynjvoeBkU42mEi5Mb5ePwz0
PKVv2HDKr6KA9RTUhWQ1E0UjsD75puR/3d2wVRahhhV2w1G66Yef9RT/Lg8GwyrH
hIOs8r8v61i/LfC8dgOG6tqymqd8Ubgp4BnCZCKRkvnPKWXd/AHk30utyUX6OTaX
rVcdXrdgHQm4WaY4IR1niGnp6LbRebAcbXQ9083ucWFJyCwotVPbo1di9Am2Fn49
yGCb/i0JJjHofdCjKODsz5/SberBBPAQ/swOWecjSyFa89Bi7rpVH0AE+mui5gyE
amGCL5BP3NWHvcT+F+SxLzlFwn8gBZXRuiLoNk2IzIVgJv+EXnQT7MurPE7oWEIT
EaPi46hOW6c6RZO3UZaHuXRatHNTrtPjbp/GKJDKOqUdPLSe7zWMlL9Gar+A5KyA
0pqTaCEHigFGOB5j2GOiApkOITIWVIAN66ZY1ZqKTo2veKcsO6LzT7CQX1kz1laZ
TpVUBfUePF66ZSKvXuseI0FI+dZnyL5VRWB21upgWu7xBgaZqZl2ZauCWoI+J4j2
o2QA+5nD387AVMyIkxUXdR1B8mZmWnrzpIYyvETxaIJrq5txraMfnn9xd0NT7DHB
NJsahbITm8I9w45hTGh4yMOKqDOqMaGBocyqdADatCeP4GoD2kv0BtDdc4rYFOLA
5eGoGkMkpZa0u2xaDOFyuO2t6TU8R+7e1zRHL3vQRj0bPde/NmeZMrb1sbTl04Bv
W6OMC2H1p0e57FJy1dEs0tVF3eOuT81st5XIRgvi4etg0+Cer4oHcl4aGy6VxPil
/kjOXIQGmkAnSUkSi/Ih2Q/YHYy4EAXpReZ/8PIVju53mBrhNvqZGx9G1XQ10V82
lIy9H8StmOdMK02kPmR41yWmPe6hiNtNmz7Ib98UTsVRMYMsGAtEHMwsI7NcVw3J
79WtRZ0J/z17aG1IC+1bzhzbZh8qphx0P1PGX2ezMIitsXHqKyY9DgBekXfPld/a
mlcGGw9HJiX3r2teJuRSMJX7Dp9NCg5xhABrlwdRwC7xUidsgcXJPN7psplVQxo9
FtW0woqZWnU/p2p4+XtQAVDm05G9gODc6tEYg0iQYKQ1+Sbn9+DMrHVRWPmM2/fN
4zsxZk4fmI8Crmfr0MqtUgTiaRYhRu7ZzTGbIg9NuPiQ3IHPzkh5lYaBh49cxOGW
8NKWcX9j2hf5jUi1fb1cbhDu0h61dqGJ19fTyGHdKbQwdwFF1OsJTMCaqBYIxnN4
QrGcTLDkl/D+kmHVbo6UX3S9bfe5GwqOs26yT0mlRs6IINkO4eXlmPbKDPB1NQFM
BT/DC7lqnHv69DJFRF8Qrn5h8f/YrM6r297WZNATH/jFXe0Aq7xKpJErz0kiHtrA
7WUvOFeC3XK+K6nsy/fA1qBR8hVCyJ3QqoeA6ZtXwK8tfUPy+cOOKv/s1n2RDATz
TJfdSsY5w1xASdR9wizlbom0ncKLC2doWvU1UW4JSXWnQYiJgE2vPqM7l2onKVyx
lSx0ulJb9ztjKNcSv2fuRYWOGZMsmiHqL6HBvx6NySijVrzAo+FGDdBpWuDSIgF3
cTvvwTovqJl+jjqDUW4kub+hzj1aJPtRZxgAYpoCJjECYJ5IikBtZir3yy66EHcU
50DYNwcBkzBteW2ZkOA5jxw4ZrnP3Go9g0c0RbT8PC3twxaz6SjmcIWU/EtoaqWm
hEWeD/HZIdNUJhtyy5fr2Zo/HD7DcNbgpheUo8vqBWAz1DsekVpoHkyXCZY4/GKT
z0JHKpSuUid5qnjqZty619WdJvVQN/2xbSPyjVMbS/YWytxshlsr3VGz8lGvLK4o
opBEnoiV/6BBhvXQuHDpmuM1Wr470J4CjPOhfs4MOxk39ON0ihWU07l92GZUccfZ
26RL5w5Xclum1uQ3ihgQ6NBkBIsDGWiIgnYDgBZD3tIo50yYKVJSzdxoi0pFSjH6
qSLkCHMkHqebzIVO4D/Fh/taHXOhCHgDaL9jXqJJHUOW+Ws+CfhRfP83szx322S0
Rf08rqW4ijNFY9+JeQybM1Qma3HwjCQgG2wNk4Qi4ehsU9kehS8PWBkvLKS2v5OF
nmo8ITIoMnb2gF18LR/HUfA6Vmn79WQ0zQZpRPpcJdfiD1UB0hdK1gpSQWgYdqdg
U1REFvXkMVipqw5URcZjNXcFQgOcsk8pbSgd9aFLEYyZQlOlEsy6RZCw9K/9t5up
fXB591obqL4A6d4GCLdqaRYwME3Js2g2zhrvsVrrpyYIcRWrD/jSmjB9M6X3tdNs
ylEMb3KeuTJGDz41Np5/XDkjieet/2cjn+VqcM9k2qehJrJIpcGfRV6N6DX8O2bB
quX2WJdgDZMamMiI7zkhSnFBRNgJ+XpaWq3dAtiRHw+Q7Kw6gA38k5m6ouizbzfm
NP9lE372GVyo87+V8jAb4zioJIjdqiYioCorEkIZjvCKaRKVn5TzKdVjlvxi+sPM
Am68gJ4wW7j+NB4QsG7jv3/RygX4ZZ7Kv6Dq6Xp2Y16fbxMKEf4Aosi/OO2hFrCB
oGwssoGCbg+LhdRwjL68Lv13KLxlQVGAporky+K5bqhhgSKX8Nwh1/K81Yb3HJBH
rbwjlDEoqYcqtrhuxqKQw4K0UdRHDIXOXvYh+4etyxN3VwTFHjoBItipVQrzGNyQ
ETnqqcAikewV5JKjNzjwgKKg3aKbnfYkBhhbeqkCyaPv+MWcOTWddiEc2b26ALF/
NY9daXL95LdZsj1G2mGCfRQ2SSeWvlW0tr/2XS5WLGkvQFa1crJfvWJGIXXTkWd0
VEW3thfYTSM+RUYqkPWyXLbeDo+6wGoyqPcJRbEpKPf8Z5FXtXTVScmuA9dk0Zyj
GKQhzyyN7z6gpjMmaiJlj7gKL59ChYUmU51qrJKDhXUPQZLpO37qWxTaYy8diXA5
Qgkys/EQnOtpllWTZHoTtYOwPxlSteJ9Opvoy/M0SoMSGsQH7mMrP6w1th5jGlBW
zAgEeD42Xif0xeU12S/vODPO3/sRccnzqKA6N++x4fynZ03rUjs0uoSrsLSK2uH3
qDEr+Ld7Ca8nWpch2x8UjFc0H1Tx3LSbV22F6vN1NXn4hBN1EBIxvbdVPu/Ng4Zj
r0VNP+1HCu1brWb0mCMrSLdrgz9sdJZ8gf1zAua5XDstbmQWANaSBiGwL+Sl1rif
3WK9w5BKWzhRGA/ZnQm27sJ96u9mE+PTYBgqWa5lKr1Ba7d5vGnStvWZcXI66MWA
V53FHKAElyLaUosxAFJBFGPpqG4YdaBpSSSrzIKS+bPCUOVKuEM4fJSBwg3u9ssn
m4RYLicvpDJEfkiKao78WhTwtqDXNmW4CoEO5D2VDD+WoMRdlkMGNZgbXDGYxqfY
p3y7EKQFfqzkTOA/9/P3LiWNsaMuLrfofNQYDPaHzrn+KUKgyENnKhTXCTWt/c4g
hnwoUXjMfHcYN/vMm1XYKBGofgjO+kJgpXrGjA18g3UUogZUIj7hbv5BYf6DCRuq
DELtDhyItRDAWMbCN0QVmt4k7can1Ih/DkIRcFHnEFDn0ClSyhYEg4xUDVc2C3E2
o0SBwPl0zI08EV3OsxRweVZYOr7G+x5nUiTLkl0b3djy6nLOZmog7f3osdeJ8bSa
R42MB7CtpREX7iNAeRNKQZdp2LuHmcLL8MXwjBzyb4yq6JDs1GA7GYwE6Y9Cv9Q+
8JiujS1ITqKcHWI9pfv7VDF0MVDq8F988GmgwGfU2jfOs+sxQ9hBxd8U+ZbJSl91
vm2qYz2QtWFns4q8zxwxhSGGKuZEub1h6r8RkDshwf3rvUKOaeUMmfWYfkJhc+ZL
hHmRspYovv234a/JIaKE6EOKQNKw1DJjnVxZf6t39R3AfMKe+l/8yEsYzNux/c6R
x4oprwTgvpA9Szz8zSu9g6+MoNVREYHM4q4czlXAn5Dm6LytEPJgsYic6P4l7jNK
R8bGvDYJKgy7a5IZKypN86UW57HfTKdHdrewInOg5PRlKW0VdkjgpJiCbWPr0nml
tSKHlqPK/XPnzMPoter14NzZAgK57PgGXgnr7U+4/tn6FjcNps8r/Q1Ni7Pea4Ix
sBZEX3vs11l62/NOOv5GIveWfQevY9vXfdSJ2BrKPwsFXqwL40t5uk4zRIGdBAM1
ZH4eKH+anyH9Pnv5DazbIxMAINrVzfvQ+J3h4YgYm1zO8ndc6kb7/djeKcyH2JrG
7k9v2T21cPxtFwLjITW7ATj3rTYFW+GT7fzbL3lPoEL/2PpL4ePHq9ldhbKCx3u3
ltMYI1Z8XnU4TQtJB1FyMNVUcyp7PB/WvmlocBMipew7ngpNTbe6XyvOsUATQfgM
A5LAK9kvl/3CNRKU6CJReEuEaQsmy1PuSKN6NuJbN9iW9I5OZy76J1lRTqnlEpyl
IA5cJQBKb7yLq1ShZv5OiIgI7uoxu2R5Uqmxgkz/KRFm0poDoGgb1MEC0lkL4uTo
nnrgO9iZk9bBEfvGJKT/wfZTasoN4o/91ADkPkx2cLBftjvfbjRSC2cbp+1JgQ5F
BfjJwvc+ob7Rqc5BQiVai8XMfnCR1M+h0uvLiz6Xe8UCbbhfhFm+9Twl34MD8THK
NREtBCkGTfGNiHElSnyDm+do4Pbrt8kD1D6QsEy5Cpi9foVqYEGXPf9rGfVO4jEs
RDIe7U8Zh/VkomiMzuBnvQYvy1qWFOLNAo40soWh2KIGYnR/lTyRdEfab98CC1BJ
Slz3fUt6p/FqADqNaDwhjBX3DEuyxuj1G85V5/m9zyUbrjEKlI7fHZpNKNzoqk/r
dI1icBPOnGtHfzAc6lc2+Fi5z1KkcZrNwoWj1ELjOe4J6wjyUib+80CgZ/QyDxyg
27hyyLRgj8KgxtB/zE6SK/Psfae/h98RjMSwGV5nXb64f8I/CcQ/Wg/RSOfwBAcv
bqs1ZjVPPYaWqQGkh9s7CALyThXtNo/zBlBDzAHVdsCB9sAAKEMq4hCetd6FyGiB
peVjGNpPt+Es2yYQKxj3Md8LQYqxwKUfFgjORG2ZFuspXpdgjZaK8I8Ut+JadUXh
MHJ9HtFqxu0Ey6Xk1oPtTNZwagcmGo1d7G3qe6jkTE4OXxFa2BLEXeGWdA83DHaA
LcjHewCr4o+3k70LiSgFP8o2ro6dUY6LqzWAWKAQ428WQxXatvLaFwa160BsflJw
nG8AI2CJVRfJjr2CPAJQ5VZ2zSegfLOY6kHgctd9eN3RZy+3nV8uatiU+4sFbKHT
mydKcFf1gUba8piRQmr12pS5sodGCh1MX7OaF0QT7j67Camc8/YCrCbWmqjL7NVC
tWizqOvY89xxlcf1CClog9SZrtVIqTghvd93VEK6SbO9A4oTWiSoJeJHzgNUczlZ
snFyfPIOrXB1f+67qB4F6BpWrZ9wKd02wOpPAhAft7gsdwOhG/lI1alPxFQzkQnK
XscDZmmVxoT707KXpxJxTWYqYYQYJpS4d6E9x5TB3TFNvPnKmT9igqHb7beiBaMH
jVP3n7RsaArKRx8IF4OXZtmW3gRvd4XPTSN4q3nN57OYiVTW1UcCdKCUGRxYyZ+X
y2MWJQla41g6O1Xnox8Q952tVGjMlbxBEYKyJ+g110u8F9pqQ4/QQmCs4O8bvIXI
Q5iTg69EP/C1MOa3262NHG6eBSCfTyC78JVUF+KfKgJP6r6txnhFVgFXtBX9nZJp
lZV2lyMym5mwpv9Oof8ICfcmLmDybht7bxZGfVmXwQww3Dt7+hhnED0bi4TNpZJM
MUHnOz/T8qr/vUXp4gQ9OQLW3eY08167OYOPN0ByDfRMbFo5Jy0URG95COAxLmbN
8gbwLsY8f8JdAke1/5rk2TYvrAXBvf3UyAKQqO+I0uwrYIPIFUTEhtCYlUK/t2rw
FBnUyxcGfP9Xt45T4gcLZUxsrENGVymik8Ij+ABs8XZxjLwxA72v5YssEA7J1vrA
A2WYW5AHGtPoQb7W7moain+ScQT4u6bclU9ZMZ1YQBM9BJxoarE31hu7zeIosVgL
j2BV1PKfDBEZC6ai3ST1MzxJj2jtzwgOoAadudl70CqeJjNJ3WwwuWjohycwmhcv
f5qpT+9L/j7vJibxnPWkKsuXHaMfOGM5nSNknkopmT2eQJbqJY5cZ4JZOUjlvkYi
nJSqCGpccf190gaNo5lM1AORn1dRj0Q93v2QeL0rMXUHpa7p+xz6GFbbm6J5wzac
fy24gzV/8d9I9dFnogBPTWnAEEJCEd5inPvbK06T3G2f+lm1kJuvwjOswqfLZ8jO
7ApgGU0JUQWfhbrnHsAO0nEEuiHTH7DwRERb7hE9XENd6DhfJ1lsJTEW0vydIUIl
Veuu8jzO6AXnx3yPcLW6senL4zCTI+zGjSPP7PZlK2Wmz8h7+bPllryRppnBkV6j
M/BmPlIwLP143a8A+iFVGgSxIYkpa9HCTaR0F1fGeLSBzYdAiJMj5EVt8mTDbqki
hor1RfO/DVGdXtmgJsrjFUy3jTIWnUmGojfo6NTrJrIHwQKxZCwbJ/8j32zuKhD2
nQ7M97CUN8N9OngEiSLXkVO1P+8njj/FXMKdO3hPyOCeQrCtSTAYAdKc6yuAOtqA
B7aNyPapfs38sbvWCQ44t7IMceYPdf0GJ/IrsMHOdWAdPn/ekDnu1ay7QZhMe9oo
pLaU3nZvHBX3EO2hVQruKxOxgZkIBP6FbHF7z3RH2kRkBCxCob5IZ755gJfC2SdR
Xg+1QCNIHx2iRBL4Csrmbc8qpMesVyJPBYJ0rj6jgfvBgDa515/4IrDp/lnEzgh1
Dj7AmXx9rV1MmRWBpg6eIB/KwVdxvevP9oqY8hEZSNWFfieoGhCrDdiMJuoYidKH
RFXnX/DwE32/tWj7NAMrQe80lXt1fF7UEtA13osUbs7nwdKdA9mnwjDjDe2aqwSE
xmtToGdPoqbFQ0lohry5VlB2F+VvcErYGULSIRbQrcSKjKVA+qYWWhAJSzAWdvv6
XltOxdQ6V3qBZxMj7WnKw+4lVi0vV0sTLrhlRlO4PzRCRAK13XRl1yz4x/wqbztS
xV0g2/BxZQ55wVvI/VLBE6iBstGNXUn6Jq0vhmfhcAymgatgz4kyuquxdzh+VFuU
8u6CZa2EmacYPzn2LuFfr9FkoYFm2x2HKLpBe/xFqCCln6Ie2tv593w/TkZcVRoi
4S6OCThjosFTQGK3NO8+UB5SUHm2Eo8bkg+Y2o5+NS6EuJtUvVRSaKs/8j8RW2iY
7sAZwm7lDwVzvrxGhhue3V/9SUQN6Bhw361QoTkg7n5qekk5AJPVyZpEuC46+JVP
ZnABlRpOrTRHAY4lgFEEOnDJG+AmnGVM53BrXWaoU4NQr25ieF9Vzxs28riayU1o
BEoLlD9whdRfbTWH6nZHyyRlJz8YCOr6bRmuizkSReoZl0C5ZmLLLlkuaWeozASC
bJ771n12mQIuUUGCEXHLp7AanipDvy1gU1RKtOeZ4OGKollivMnLpYkSrW3kCfUr
4AAbkoVcNJRdovcncC0NhoPXdXm9bFHofqjvSLqRiwAikv57bJKbD3nI18wdrajc
6bMKv4sVixiqkXcRWS+zgoGJupChqug05sUaXKusvBaNgX9/4aMKcwsfx0EqIXuQ
0i0QBNRZHB8GabGRaFFEz++RKx0+nfuq5m+xXhU+lcY/00AsjaEO+WI+f4P3zH9Y
l2BdQfbhsROmdVN5MNJEgtS+tRScaF5Ib9WRmYEXsf6F4V3073Ovaw1DGyFQc+oG
9Q7+sxHW7OEzyy7pRW4bpny2t9Q9WPZdYx86utS5RVY3OvXocdslRGgd0sySp2RT
ygv39Pcvlrv/72VlQc0PzS5GCZlBT3bnjN6ifvZYnmH5DbE8kp21XH4kxSTmAeTb
qeshnSgRZ14d7mGFSLnnhqHi1RjtLKJ4WG4RZJDUDdsQUKUm1renoCjyQdCl7SsQ
mrAzsYxVQRxLAWNA4suAk3rA69Vqg5idbQxep35BIcuIszSc5WUWNSXYl1kpG2+r
QUFs4+FKL8eInwb0cHvZda8dxGkglbN59YpkzvcthT8EDjfWEVkwtik7lkenKSPB
DkhnlZLuPx2qH7c62Wvot2tOr5TcAdYJLNeyr1LiYD+6nfc4nOzmWVNX2MVexGBd
yTktzsqk9kWaatTXlpbEjeM0FPGDMUksvK7CYt4w6OHMbFSMqdkBmUocFEl/8Puh
xA0WmXlc0oLs7aIOarCRNZoyEQdYepiOdKmwUBOsQDoK8oWFV7661kn91VXvqevd
PrDl/j+nhhj2ncd0IJpwkcvWJf8KfogEj086M1O0AeWwOkOjWdfPVph6n2M1tf8S
Tu8eu15qsMg6lG76Ue4fBDpSGjuu8lgFdnoQhVXAujaVtX9PTuFrHue8YD3NaDzN
KN9aIbwR6hymAsGatjVnlEWMbPvew6HdSP5JG1Y91kWwHmGMUibKKyAfWaRC+VKK
LsZKh+uF1vhwkERtgtES61COu3zp0l1CazwnDDfIvzq73tp3W/w3UUeFj9Y1GG5b
FLwej56HK8wRlp+90DWmbVtwyBoaAOiL/ArCnT2Z3mG3slRAOxhszkTrkQMs+hm5
e8HscU8R+7j8goiGmE8cOFZGA1/FNiRXeGEkOoE1a6igAxU8xYjSGovwvHo2EE/G
h4/CCEXBc5hXN60j+uGKTGGoTtxPLDNgl+8emTE4treN6ulbaBrqhUvbYo48gqcG
gpv9S9JWgATsIdcei4V7beOu7QDcwaqWTLqhizgXMSe2bizIgEwvQER5Y/s45RAv
gSd1Gm8S3ywan5ei2wU+Kp4pgzIvwhCOhE5Q5J5qdbuYLzG4iabPsAzjxIGqdfls
bkVN+pb3nYpNT7UPr0IeJ/p23rBik7ZbRogjfw6q1cnWFNEOnqJlH6phzsR0AvyS
t2eO9WPQYYIKF6wLPKLgLUOWr42HmsHkTgEPqkQHyWmKGnO6Vclf2foguuX7zMCy
EQH5pd6qMzPuTzVGuyYEtvw8kz2J2sMiOQSdftLrjKvuMe99HPvqYH5aXsgQiLkl
G5HsLswuJ28Qz11NKq+5ip0gNoyFizZJrMizq+InzK+Wt9plJG4UCerUO9f5zzKr
mPsOxC4kG1oV1KqfMSDb04AcoxmOiPeWHcXyTSFxpkIZmQHRyNvCC2of0nG6j1X6
5BkTgbS5t82wwQVqOsEvbNEkZ3/BhWTGtTiVP5nFNwmoT8TnUc2y4zghHlwpdfOk
oaPR1zodVxApk5k5KLOdIyhX3EWrdK0c7JerMBc3offhIyce1QsMe4td6I4+2FQn
mOOo7LiMNoAJkKvZR3Un5G4mCgQoGIXeJan6sv0pTkDjX8ym+oN0YKsORN+II4EV
fuF1w5CTQllgC4C+aHyL7WFId4s2czchkUuonfk7I+AyCpHtTkNQSiL1TRKW16Zx
2wUgot9ux8ly/9Wf6hyCN81hh779/aE5ltMYNRw6o90aOVuUh6G7yJiyCOTOQPYM
3hbYBnZkiYeIMnDGM/wQ2We79fMVedhVSQuhP1NeMP1Nb0P9e1Jx++faGeb5HXA7
+q2xpjfjL11Oim3iQRIBjyRhtoFX9mjM98l16k3E/O16lmfm7cLbKte2q2Hgfa4K
QrMHPH4XVdM70icfk7TnmGIDoLTleDQNkctvqFvJR36TAzcNBSkOnm1c9LGHojpb
F3NAFeTKU2Rv/h+/Nf0eFX7y/CXif+RmRLd3n25MS8eOTDs6Pkt0JT/LKZKHHIMi
C6lyCFOptvLARZp1JCrZOpzZ5xuCs49Bb0xTtCknZs9fwzfjczQGQfTBsg/GHZfY
RY+kBDWHL78W7ku69/ZM0d1k2WxR/PDyhTt6bbCwQ6qdCku/RaExERAvC4KxUIMX
5PmvBc8k+b4SYrH252UKE0BMoroyIsT6pHKDAShMExd9GkfRSMQwnmmPYGD5Ka/2
WOamSwNn0+wsvvvRQAmhOOWQuqaADeguyKoYY6V4V2qsREGRFNo9kIb6v36Gm8ah
HzXRxZYOHKQxB9s5EPsQI7zYFJ/d0upZ1nJNp3f4JPNj6Imeb+L1p7TcKeaEhqS1
a/48+1U01glzp/KHBVXslRxdXRNY8nZsbO5DO9ZgOeB5RomWbjWwzrP015TsAkd5
WGUowix7ORy3ySU42U0xJMa3JD16m1XEzr4EQKU97BQ3fRCryVbF3qPAhVDR2y/7
lBSGnEhqOf6pIEqvgfGT//Gtml4J/tqLOkPEwZcH2A8C2eFAq1pbyMr7lSPlBCXb
B4RpCJm7qoU4tj1xof0Ri3CFbPhVxU0u4kbPYPTI6Gi6fJ+ybXq4BCgMgo/ZNpJC
OK7Dfl0fzLnpuv8P4tfIUk2ifLAU6oq72d0DqZWme/Imv1xu37mlUq6eKGgKYazc
cYDhUM7BCx8yEbTDp1gzQI4g6Aq2jY3C2nzp8hM6I6fG1lx3+BWvZfs+4FdiBqab
fm5e1cSiFlCeupzfdgZ31asRil/RJZpIjD+k7X4xLRFz+6EwMgfB/fD5PfJJ5UuW
6LVpSGGHfMzXUctxWOhveWWYL+WE8QdK6ve2Zb3hR+n5b0wxsu9+/hzDzrD6FLLy
Jwq856PCRFRl3l8T+P/AKcRn14/db31rhInxswWHCtWSQZg/FTmRcrNYQ1l3vKGy
PPAqo8XPMQBxdqZac3wwoDl8705TDIPU20gg9cVjiI0/SW7od57acFtCOkhjgoFd
PLNBhTocqSjZwNlxF4k16I6NNvAGQdrjSPohk5lFEoRY9oTydHUi9rCiR3qLdeNj
oSUF2y0g7z65JvlRgxypausCLd21fXOrgja7uLJH6PWsCMquOTqbJ5B3TpduOi54
34XpKh3YaTK0Uab0omv62ol4ZvBZPR+0FmK9jBLcjUGJgLJ8BqgAvW37+hcZrQJw
czPrhB+5zoU8Cq7Pf+8DfmdBbQBm/t3eDRgNAtznn/j//mlE60be3PZHIPIIqEBd
EkIktDutbjYjVAluFQVIQLis7GABdEILwdBJ6EjE2pxBTPhsQNrBRhK7u4g4XZbk
w+yt7NW+8yRDYpMeDYTvQ6mlhHJ0bf7zEzaHfgWQfthlV20jWmpL+KMzMrn9pKK8
sZOdQolAo73H5oPa7Rp5QaOavp+Rkda4StuVdFJEg0sOTE+/PmunfRs91i5/ICpr
YM4+kcsKAIdF07TxUkXIz+MZoRRERuXoGJbgJBU1JkA9+7lMDOSnyckzYwsP7bfs
PGzVXi7Zciniem/FpvCMUq2edB/qmMSqLP4H8gPCQYr78XaHkqfzzN1Qs/FfKp7j
y6uX7zW5X0cb3Io4gaynWIuoOPRaBOQIy/bJFuxNptQQDWfV0ksb4OFRS6OTPeQ/
bPPFoKQtWJWDtJlF3RBSJvYi8VGXMeRRygwOW+50N8OeM3WUrhrq8Xf8wCixOai2
uxh0GQDSvIOdVf3HjAL+7yx82fpIoetAkXjP3Fjncs/fxivMhTNoALo91XvdgsjJ
e52Khi7AzkaKZVCsTcoX0IeqMSQSJFnKfmRpXYz1sm5wabqRQNaOAdPGCodh4zI1
ej2eejSvZJVB7einlIkwnm+YdqmUCPi0TYamdNxS4+GdWkUh35TsOBYJuuN90KRM
Wvj/uudNbq3JaPwFDI2ivnLoWvJIRCJ9od1Re0tdp6aVzHJY55GZgT/66jXH4m/m
glb8lpNbZV0Uvhx7oVFV+iOiuA6oQ4TC8b59VLJtxQKzrwalz5VyEHAb6FQ56qoO
zPUCNR+r2qY4AtYqrDo0Q4LRAJNSh18nGT0wZxnviWYzX4WR+64MCpadZzms8vuF
41F1UttWgitjRTk+9+Q98Fq7L4/40/mkp8Rg2IqsXBdFkHb7ORXAicisOC3oP9Uk
zqXihajzIXT3f2tU4UT3FjUcfYB/9Ph2F3OgryIDNlLNgRcSBQht5bOJhURtczyl
AvkdjJsNXa3ytPHktm5Mb+j6jLpMn3164j7hA3V1+Sdgkp08ks1PzR+rBfU6en//
aU6I5SAk4vGcEVexuMdUD83R4YB+3jMTF6WvQk9N8yQvS97/l+aSHq+TCleExemW
9K7C36IKtMxJ4KKkVHaTg6dHg8fHIjJ9lWlHmPUTPasc2pzNie0AdDSb6pmQKd0J
zBj+IA6pmwii8x72xj1xDDsKPYJ6GCjTbItltJw1ilktZypwumOe1DWJ/fXRqypz
GoEQpEroueDyD8scD8Dg5aF5BG0OOxN9QcangfQCEMJqTzSK3+L9VXDR8pvtqGAb
ZFD+mjviLBHHKmjXL9InsV7ty80RFm8xROzMclvRrm1PznDfjotJNMpBLjJmRb1l
ltk4llbpfhh2LvrfhbU7nJBXlYIH+04hFXgwZQxe8kfR6N/li+jfDv+yCDWBDh5C
crdQTrV/3hg58bOoydtv5QH+/H9Rnje7/EcPe0jjKs3eU3f0ZTWQn3ceB2FJ97m5
iiTZr7XBxiW67K96CanKnv73saz+Q+iGiW7Vvr7Hpg9RS/9FBomMspWWY1opwdmk
NfM/pvXXwm0SJZkxUDWzeKBio9Abpljegm+yJzdZlTPMhQ2sn+Ub5QiAD/cIDb3G
gQo6SBv90or794I2O9keKjEylGOAvy2/aaGVn0RRPLAuyVfdg8++ARawdF9YddMk
HddcOD7WJPn5M2Gvyeh0C/Qu6RHxAG1Gy3qGRrCVnaEzp0ld56X5EmYGBR/W8Wn1
jwMNZqLN7mnV1DU+DGhj7qOfKJJyPEM0O7UBBO0nnWqbS2aegZCP/g9FsuvwiK2p
VJ61upqHPgooY6Ti0PhmizGFsS7gNqkH1E1IsJ64QC/fIJItgWTn2cnlH7dU+Cem
xdqLYyPvEOD0ALBNXn0JSSL+u2N9oLstR+CMUbHZgk/UxfSqFKfZEeWPX/htpHPN
tz/oy6n/dLKWE9aB2YxkIE/YFkwVD7jjqAXaY4FMhVl0ECyrn3GgIAgqgcXcxt7S
mlk5KWc2k/QW5SxOD+Hfi/FBl7gyUB93ui9yl+F7guQszPBqrifNydc9g5fy51iP
d+IuCIil4UfXXhUUYtUjGFHej/Vp36gjl4mSCO2JCf0tKvMKsuMOEPzeo8cP4kjS
f6l/wcFTJTpbgcd4g8DL7BRFOtbdT14+wuLr3LdjxKLK+E8rHCP9bCCSdyNz1PYq
TexOpgV8g69tT0aTo/+pWU1gkGXIJSOaDLH0flUnXxheGwgqxJR7c/xKbK/avCPJ
mfQLZbgtnzHCv+m1Mvg697l4/vjdFSYpupc6DtDaT8BAat2eff1Ht2ZobAk4LMLl
GV7/608v7816GnvVQtusCmq1SDZLdL6H5YnQ/FVEynpI6CPif7rzRhKd3wXsvnew
B1/R40lgoeG6IVvR7xEUxU8LSSOnx/hnUkJfa6OJbzzY525uwp8aRHqsFCdYIjuJ
9QArwSmQOST2P1U6BqWBz8JI7zEjj89YTDSWu2f3m8BMqnsbfsj6uVhbk29cRBpZ
vehuywFZ0QgWRyFbHZxWyw0SGuNHTHoQgUbHQMrekpVyQK6dDbCYD4AtogLb+m+R
dec+BRU36LbnknoJbQcb5aGbx6WKYPhV/raH6VYM8H4u1CoDnJFLk9lfk/x92R77
2UyWVF9mJxKW1LTB4chejnnGHBTKGs9nN+52p4MJtO9tjMWmFnlnCxpywRiK3CMM
2WlKM41cyhCtWDH8IRn8tBouAO7YQAJcNFP5N6I3iumwqAi7d3kXaijtKxqXR9BA
aK9z2z/V5sqA+17YtDlgnh4+xj/hkjYuMSIhPNfuo6SIgd/ezyK+ptKdKPM+/FiT
LrjShqlbEsz+yR2j1+dS7uCliwuUNDO/LIi6PoQa1bJbhAFkE9R6xciG5uGqX3S/
t0UmDWLYEjhkN5+9vBsIRpZQV2PfBl6504xF/f+1cJ+xR9IcE9uCtYct0FaHeGyq
2LMrGQ8CnqK/+KyxN+63KnvYU6cSiGLDPXuQ5yEVU0QN17MxjKBh0zjD871uYxfz
EALJUtJwbbZ4qGnUB2P+LGg5Hj5l1BqXczsFUmPzV37D5P0QZbbTon7CeV0UAVFr
aKBUzbQ6kcTbe7EU11YGTCHPUlpUg/EF3h9xbDKvaUeikQdlh4Pjc5Rl4LSkdASf
G5Pk6OoXgd2yX0uL2jKt/UnoCN26s4M8ELItUpnwF+ESRHUaEds4XxdK8PBTPVbf
+0y5NKpftOTSIfFBrzzloL9ez3Q351xh9G5vWuyCBSZEC1ZxPqXDp4m4EfwbCbqb
kLnUq5TLEmlM4tYiq2tyuGZ/741nJV1eJNEWvw5zGH7ic8XhZEdlu+Q6Pivo9Q4Y
gZJiEUdCjAGLXz+vjhgTA/l7wmk1nAqTgtI1pERdAaJuwXWYH0XZxqkq/B+U33Xf
uHhQckYX68exqErGXc0Ljs+P6IUTVfwcjtxzmXvao7WKOjpUljsNP0oWQf3ycyka
yGgWIJ1At3qxDgt3ve6BILaEmrOvqTmRpJtJ8Mz9AvXSHuWuSZrbrdGft4N+uj2T
RQDzmpxE1SYkPTglauGpWsjW5YNMMcC6P5UhVoxF8/cajca9DZTApmdOYcXeGLao
qkx760l0H9B15xvPZpnBYcBVH1cxbkpuBaYPEmgag4d/R0iOJgUPcOK2CWMtM3yY
UvB8cq2n1IIk3jlskxlOVxv5uu0hRogZxPGlOj0VP7wGO0yjc2V4yh+sCfRhBn/N
u62/h7WjyO+/fwFO2bKH9GCxKD4h8H+TlaIgUOlkoc/za0y+Bd2ol2YmezqMM0SB
mnQO/O6VgwIsoxJ1VU6sdPFYIrLTxZqdnfNlG9tXjNg4PNqI4VCJJTs2+FlVDZx5
xKSxOIhJT3+l6gi7XOk2rcNz5xM6+uMVH5jgQhFOoIdxtb8+Jy8TnUcoTOAr52I0
U5AUmue94cb6CkqCYQ8EkXIR9g0y+IXb8FBPz1ckvohlhFTtCsuAPUsnFEatZ75I
MijPnnTivEiVvD45CUc/r/PMWy4SmSiTisMLG98N2DmoE9jzVVf5tqUsEyAT3SNE
qpDoMXwg+bFmNYAY/+zkm/P0rocrt+Gf5Sudfgi7msrZORTHPhJuJlzuJ8PMyNol
tBuGCgwkluEb6oKxeGs7LL2qS9BPE5DdZpnyd0aP5/JA80uRIvSjk9NLED45RF8M
N8bdL1zRV1Rj7G0Op4AS8v/Zgg2AabZUcmN4MiygPrDtwBosY0lrQ4/9C19L/dU5
+6W9XAdHBGJsHvvm2aJCUp8g2m6f1lBOZaFg19k/Ii5ygr9pYftedAfc0nvyw2GF
ZbGP3+/L8pgMnl4/bzPFTCwhG4MFoAIvSDEzTA5As9EAUQ5SGQIxXbkEqwT5qUfB
ZVUQdll4HBLAyOlG5dje3FJOr4dyZwFPO2pnxw8hAxbBTBqHYFncspS3vqIft4Bi
8gijXo6dSfAJuOZ98LMLj4q5q8Z2quhfDeHFjGBPnzsbrHhkPt3mp3IUkdV7EBrb
BRNL7+ID+YLprZWK5y5EbLGRZ6BTtUmCxed18GNympW8w88Hp3yBz16xgmO8oFJP
H26jPEl1Axj6Hpf0REmCtb06w52YVTVlbx0mP7NE01sQWE1kcar9WLm4daacZqvg
DEij9krQfzj0FU3rxkV43Pl7Vh6uLKkJ2ZDbNsVAZyHTueSdPxjyxAG+QKMLbWad
tiTSJHaGaVC7WKu2TGJNotk/zGJuQGXWEstE8kX1qlQbZbd7Vvt9KtyKRtpyftZo
ggi0MULvaP7XlcKbE+T1Gv3SeOIOGN86Cd5B7FXRyAmkNQmlsq25bL9QAG/xS0YO
xYwvNqNcONTOLylh+ZzzV32Y3mDsnKUlV57XcOwA+YA/lqQmUzejmnbTj2e4dGOZ
E24yD3L7lp4OOsH1zlO18NBC5DC2ElBwP22NwVjhQ1YtLjg3MoWW+GctHcfcsLJf
3ITwOryJTRc6tv1/cIpl2+r2kQQAOBAHxNgu+auoWvJxyEU/+RGAZhdHo7u7WwSK
0/6e8BI7Dtg2he+tZeoVV61Sphd5TlpSER4RSLtNzRYRHhqnpRIIgCh/XNeqiiMC
vPzwvufvas2UCMFk0A3ZbVMhSTAR0t1Tq8htyTPt94dwcXYX1WfMaiMy16rMi6XH
/ADviw2DhWvfaZCmtOvSuYTpjMDzu9KR/Wf3q48XQwPgZKSOaYYT/bzECasoseoM
UUKdfgsL8KeYt9d7TorSXcgW4YkHYzPT1Ds3WSNenJONaFa6nkT6qilTWVpO1565
e6GmErQ/KhbCdKUkqJPdQ9qc8U1jVMeDrDcwXlDJY9BHN2Zga5VQA+G0iKKc6gXi
z/9YIkq95x4pwvRJDvgr/bFr0TZBEPoiu1mjR2sSmUmIGQCfYWeXevKWsf99pHd2
7hVcEFhtbTGAu/Yg45ybHoJwdcqHHJxBZ7F+CfmdStxFNO+shuDHe6skbxBKjgzk
i1L2ox3cxLS7cGJnNlsUcEzu38ij21BPcnkIQSANK1e2mwW1zJzPSgL2SRQVp6D5
LQovKWAEGpQyEesJx9QQvakx011OUvbjpF2+UqkDIrrjxsYLcHi52jhrvw5Vbfl5
suKd1XPnEZucLxsYwXU0EcrlgATyazBqhS5oiqNxP1VrBRfNdBknKgBnWtLpRIoh
8JFDFtex9zvtXgMCsCDmSEQlzVDW22n16eQiaqyuXVNC7fAAYS6gSIxFTGKE1Oge
TQf3WkBIBfNWn91MqnHuifU8DiRC+YbHuZxuSP8ZggLEN/nga6NQahcuofR2Xs+h
7ByHad5yxlEV85i295iSREWmztQO4EtftXZq2YDUfLQAFKXuyEjOKtGLsd0nn4Hx
raODOZgiXBFhdjTKpMwDTrc/grPSpsUEMI3rYQ29L0ExT3XIflv12vjvKFsBCSqK
6wL6K/+c9d7wxXcRmuksd3Zx8M+wxkt5UcVnPkwvb6b9OUxFZsG+RgwIuOTZazYD
PDkvsS4pLDIYtHD90V3FLo29vIT4u72MHm0QAOnDl/A2AbsQ1+9HdgyvPcXe6TIR
0MA/To9+Q8ZVgtwqtY/xmYpT8Js4qMEWzAu2mXfxbgjJLJWmcYLOBIBwzpMho+Ip
8NNRj9M1tjgcWXkjBfRVAkx4p+zP/ibWV+rWvfps7CdfKBHrbEHJpQ76JwdTe5qJ
7G2kyrFUAa11ovnmRiAaHYJ044bmYKAXIjc8Aw30+yKEELjqmn07WZSJPGn6xTcj
l+8OmuniekpN+j9DzXtfNUkfffqZm2yy6Dwg2AqeFQ+HR0sv3VGOfnO++PW11Hn/
i0hnBaMbqyPvFuPur0PFQLqxMt5/FALrXGjd2/rC+iu4cu3lJM6i3P66yYuRABuk
dBFaU7kZB5NLv925rusekoyPR48D7dfz52F5HpbMPITXBoDryLNEAtykwYfMuVWa
HurBFBFv1Eb7G4PP1gJJ9p5kvVEfNnF3PMtEMoOipKmXYxsGLFWaKrgZQtP95iPg
BHKNMLRGViO1dqGu6QSJ82QGCpMWJVbJUpG7XTHxI70s/nxZ5s1bcQz6siTYvb9W
tvJYiApPqkvq+hFdYkcmBAMHMUrFfAfyz+crhm2KHZTvEi4tDbEQmrgOJDtoef0i
DUjBdcz6ezxPKCYFhw+dBdGwfPUoxSLnDqg41d9pv7IpzuaJpeaK1epkBXdkG3SX
wzoIlFuD2KD0tBPS7Px+f2zvSubSdl8F3W0mEn9A0I0/xE0pxZvhCBhLK9URW1yi
tIsNKTQyqUN0bt09ru1NNrMQ2tSHNRzOa/fH6ugaBq9Sj+wdN7+CbqYjzp3S2Cdi
5cA4Jk/oMoOc9+D9qOeva00TvKTO99oSWZVTpASW1HLrIdVNsYQ2yoUd2fL6JTuH
lOzW6FYsjd6rj/42q+CG5bqoG5n3P3VclM+dJwBQtc4JN+rAhgATIwOnNGrkOhla
KUCI4oHKyFMZKN4pJ3pgjEUniTgbzNKg/KUAhvn+cA3y9LShcgbiwFi0FnmqeS0E
2Me/CZZ/Z+SjocAok+j+mxATuUOl/A+s6oH+IT1iBTVjOtFPVwGzAVW6ysqq5dsl
XX/0OnJ2nruQYZhYnTuEZtS+eC7I9/KBmPEf9gjCHcHkaMZSmj5n/+ZDfl7zntcs
yQ4IAvHqTpivdEiuO5/0k4icoGvZw8oYeCS24s7+6nyE33XrVDqtoLERwkV9roBq
5SdIDA5cTUZEqsy/ve5rSLTCt9+AKI/X1N1puwEbG2UeeeuemuCmIQtH1hVxyMsT
EzP03ns7n7eujpid3hysj8VU/lZgP1dIR4Yo2/9k1GzR08gsixUOes9KNLrtNw0j
9bnHk35B1uvXr8Tx6ydA7v+ni3/Gwo4ZWnMsu+4birXc5OnHcZ8XYqx96aO4l1eZ
DN/DT8wJ8TXTuvVwspTN+uRStCMq0Rtgl2wZYTomfy8C/gkInNIohwaels8HDe+F
a904eGvP/K/YaNAA82jFbCkbv967rhnY+KSaIwqaTjKFoBzYu/K3zitlXO6DROn6
Y419PfG8kJkZQQDEQLa6JAUe7uLt2M6gXPYNXPw+2qNDSauajG2LYN1jgu6RFGMq
lHHUXkApBLDNxp0z+RA/LP1PDQOlkkDPP78VBjbYuj7WYGrAbtyBG6nPHLrJPTcG
9l2kz1vNVgjE8regHN02KcSrPbJLjZ2LjdsmavpzSPDeLaRugACltWWMSo+YWBBB
WhmrUoRdmm38ikjIaSBDwUfDEgZQQ/ZOGMaOMVF/LL7EyAzjVQBmQYQxxq0Ml1ik
90DIuSI5Ux8v7PFO6kDzhzNYWpe//R+Z3XCFqEj3STjA8EaakCpSlHvxyUBAfnT2
GrRDJ0xyTdij/RMhVmBNhXYhqYZcqUbDz2ptnb0vPOsZXHWTNVkLftj696JAG8vM
59c99s21diLfYVHQmwPde6NAWEEg32f1jl+kIfpOlMLode+Ttf/N1SsTfaOy7Zt+
CHrN+eLdPs2DhIr3KFuutkqk76sjq+h2RKXkAC58uzjON74CMrk0R4uy7JtSPG88
xoZrl7hbPA29e01rTkBvbzWCULOzQxA3QePBkgeeUKax06y96vFlk5qjYZM9PdR6
wrdJGB82seWMZ7SDCehlSpoGL9l4jKWbIaxb7Qkwz175DkZ9C52u9DNafG/FimWz
joB7yVVTBrfoZ6A03gmHhpNVPE8MIDVLQA1s2kXh5sv4bRjG+noXJDHyaaHP4xRI
IzaZP+PKHfJK8rClIFzDph1A7rCHAUv2RXumXQSa5Ui67S4zl3Oq4Jtqgrz29Ng2
ufHMykpWd16pl5lVOuRmoiWpu0N6xR3LhEUznA8VgJwJRqB8yp+LYX8rJQhOo29m
CdyUDc+Q3YJu3+qR/oZ7931GAwxjU64j8cTvH0JRo0pdsQ6i22uP04a5l2O227iE
7Y/gkuFuPTII9YEgxGLn33Dsv/0x5ZnuDtfehZrRkMA2RirLRDPgHs8XIF9jLCFH
xXpkStSs3d2oufLRSvCcwgtZhCON27L8c+XfAmcMUm0+L6I+xAN8sgVU5mmA2kV7
+YIrYwYt0rRUVGqLPUGl0g9NJjKYTkfqEMhbTAtVt3kG7PMrw7ijoyut9gBcF7o3
rVG/PzjzGKRmcadsAZBslere3+dEX0FjyBa9MgB3pwjY1EgDK9zYqM9OShUtstJK
9P+wlpYOt7icdLKsYaGp8xCUNQBLDELA19DWbr3MpCsuSzX+zmwgpnZrfSPb/CMV
mHnK897o/ufuGjwjs44GYhV3aJjciCeI3mwF0U3cwBz2YyZxdnrfzE0ZG1fKszIa
M1V9DgE0qtPbjlikKUSYeoms7k6ClpoxcW4s6tubXEqLjvesXrrP+rI7iynj1hN7
h6/CSXJFA/+ePSC9RFxa4q6+DBa4ReBWzkoYPrzHVwOt4gT/DPYjCn1DYznkPe42
+ITNsFgcx51LJ17nQp2mzpO4Y36fUutmuDV+fieY/08XSwYZT1smnwYp1rHOky3d
iE3Ids/1L8Zt9ujasbHNxdAXEMRU40ItfjQGuEA6BdegWyPjQbPUUVQG4zQkReRm
2cYr09mfnys5FnI63yxjAth/ukHZhUPcvCVgMA/397Kj+cRgE043DSmlHNoxYfsJ
grHsREugcdlK3IlSvkQvMmanmfs7a5kv+jAl3edWdj7mnYWkxUPYC9plNtJJuygX
djvwmjqIWhFPkMe6LWbVcHqMvkBRhN44GWsoqDgykS1LTJyn9Ou+cgMLluXRdjgf
9xPy/5ZixTWmMw+5gWm9PDVmoqo53AawOxhfUGUUDJzkKp4GWvk19Q0mJqRzNWqw
bdDisywKjw5HewoO3NLJ7J7YXHpvhQQtLIJz5cH5g90UMu7032KadI139/ogZv4l
LdGOGphkbFXfL4pS348RweLgIX9bH64BG9C5kqyKGjmmv7IFeZRPhUdpgpGrKk5O
cTVmkyk7tyiJYXGZPoPdy3olJZJ5Z22pcDWTN2BB/tzB7S77GHTCMDnCVGc++hXJ
dfirEACdCBSlvmsLcucMDKGZAzr2QdPDzWHckIcP8BTJSVgzzB22nkhbvq7iQCHx
kTPq5PZULWBk4I9io9+Wo00x73AijRq8h37isa/eBaeubZYfUWKS/vhVOJeW50mY
5TMeNN7/heDI2ij69gUWiIIefoLWwno1JsxcXTl3AK61jiQ0CyKFbESIs33+DCX8
A4XTTeARdjXePuQDUqLQvDpNUJWlFQIGIsYBIGhKKKzljmH3JmZRXWPR+lCYLqCQ
N5oikVGTmiirZXGbRqZC50/rf8LmOqSqWFyOSHJpMedRlofKWJWCiao5QD0D2eFJ
65yJqcGVgBsd/dup1gug9yqhkEuIv8QZCXwrnMqz7z+kkyG2xsDoGce/Yn1kNMcq
rKdJTBp754qidBMxjVv/RDgUDXRrkr0SZDTLeQG7sQl/r1GXbZnXed2ehuNw457/
ut6s7q6uGuhoqLjKWvPXSjSQQCVKTp1PGbDMlxODWhULWBNG27wQYgKb6QC89V4Q
KkmGviCjwbqBfzmHQNQx6g7HW0Y42RY77d5vItcmHUBAPO0RASrkCYt7Do6X7mIm
Ti2H2LrYf7QicNg/VX6GeHUjePd1hFU8QwJnlaU7Xw20jhlf7wwklm9SQZNj3I0T
wWnseI31Qh4J0knMMN4xAQ6lRDa6tysOLADDpFYHmLqi/0eKcSzbQDQv+xqFG1W7
w0cuojBYzwX3RQGSFrbbdx9i49pcbe2CEA3mQJFzLLKCjqLaoXGGsAYFjsUwbmj2
+rf3p+XCHU8Ei1K8enDwTo7qDttnt1Q/sF4+XeVBlKZYte5vAFvRr5fre873sE0U
hzXtlA9C7GQ3PdD6wun5fXEM/8JRsNVAJ1wamlsdrYJEcPxKYvYGMuDKtTo1qk8Z
OHGIr2rYpi5b1yecNs1F5aOjmhkPsoxvUalWHa2A5LVfHzYy0kDNyFexjRBWI7ed
bXDwFms+SYx5bDqHpZQeHUI1iDNSNzIQMlpxE+6l9zIP576zRdVaT8gIGWSkm0AJ
JJ2opGn3n4LrCcoBnPBNqeKB5DV1/dxf40dmiArv9u7fIjxritOjpqXKObZgLY6m
9ipy/2hfbncI6yu0I7Av0qqr0M/OdiYBJiblqfiUNphvC6T+4/tumbBd1oGaxaW7
Yf+8FfRaBp5v3n7zAyCRr5wIDhmi3QwrVc5ImMcelRP84SUYt8xt1gh1ORBnKG55
pV8GWy0Xv9MODwBbK1vY29svmbBEZmVGCU4XXIjpNf6FN8rBumgNcpbWdotCwGpl
o5u3+B/i8J8HEkAzBYwzJUd1gPd4AcBrUbeYkEo1wSlG1aCxf0Cy3+YGunYAF5zC
88Sew42KHMeAWSWbpFuUhuBGL3XPv2m6rhCMVA/iSQcYsM7VsCT7D8wS4gbQpVv3
btFr8ye7DuOVxmafzZzgahyOuCiZr/Cttzmri4y2RwN/Pfd2ifex+xnj19jaGmU9
Z7cnvMdIpGolP9zlEt7fcxciaoCaDfohJqRoG1QHNiaANMuJMeOL7UiAsbKj8kcw
ZptrvKSy9RYva2jNnJdVK5CxhNI7/rMWTz9zlMrEpeF30hYnDKgDz6kRL7/oBzHa
0WECgiOgtoWq7wt3ZohJL4AXCJbiD4C+KihqytTasD+hvtbpap/BO0ifDB2mZeHP
3CtwABCqkpDA5OMvnK/DuMbAZmNIq8bAsih08dCgkyxnv2w8vokXIRJqi/TD+vNn
9MUVlThYs8SMyqlJWBK9HXOedfyJeFBAJJKS3RA7s9Lms0Ba0ehIQu5VahiiDcXi
yq76OEX4L26NslkawddEQfjlQCOeVJJXe+pyRpxmn35OWglOeW2e6VtiyM8INlEL
0SpYw3F3JoKpVbAOOEwLD+VTNNENOF1Kpeu7Yt8C3Q45CGpOjXKmc2bTQzUQ7bxe
FtdaF69F8qc9+MkUHvJ892JQCvhIcwXg8Txx4W7GYfG2bU03zk1h0bazh69phrNo
1rSSuYK/LYhpgciUtDNMvN7xdfMYT4yTDlDOLZhwkzXzsvp2jqGR4uivqgBmXewI
NghvNxXDnZwFGN8YAbv3hu4n15qF4MGRWw5w0ZLW3+nLml3uGDzR7ThL48iAVGbU
nOrDdg7JvXfwz2jHkomlPE775wmUZad5M+97j6hjnxwq6+eFaj5kSZKHBFlAG5Vy
V7x7AgAB/hfigoExRlQoJcO6zQMo6G9fAczSEx139JqGOSB3t24LhRs4JBOe6UXa
8u+jEMpujeMHx2wQibIKVZ4hNgDV5bcIe2DyJgRP83SDHDNcmuck7p+Jy9Kx3hBQ
mjw22UaqOYGIz4/ecW4/6g4kOGHzcXVPGe6dWv1jevUKP22h3eOLKJiyq2ps5QZV
pWDluFKfl3MrDV0XnkW2j0ddUlnVcfkTzSKbBqp9ab2BW7Xo67g7E/1Om+kt/EEV
gFbx23gbM4+ijcU7tDEksYkk0FIuvSsmWnx787qXHa+/k/9G+iDZzEIt1LcFuPxh
JwMAVLTz4DwLVNHYiSI3bpNfxi9P+0zN8dKpxVLTMQ4DhWzoKfqIijRlf1PVTJWv
Rpn+ul656fbug7imHky3GRyhg4qT2I0SvGmHG5f/sxgf8QBKz8l1P1ykFkcE24x5
1kjM+qmouRDi+ZZkmQBRs8IM++uZKV/8Peuq9mrBmqMnypVr6+ATL2RuoOVi7ukI
Ry+QWB58LEdPJ11uE6IQmMB6y27UXnyzBzR9h0TTQPJ4fvQEpdDsUDi5KIMwwyw3
bIoEfdTmXSyAfjZgR4th98qutB/hpVzP9PDNvYs++tXqxAK0iBVXSPsu1yUybpc6
lyoo1eUx9pdhiExFhyB8toRYnd6pZcFZY0UQ8o4hLYlsR6DLiLRkgsErHEghf+/E
c6mbLvitM4F1uiLx9xQK491NIp5eT3vw7RATIyJ/hC/v8kY2R9P0eieV3K0cpZxB
4mQjskKJCAXbWCWXCWDs6Mf26ThwwAzeOiDndI+3HUlLnoTcS/oyogvnGnaIR96i
BaOz008JhlFphyYX6NkBBQObSjF0J9MxBepjP/3JyozABthk9PFSPeh9Ng3oEXuJ
bBHDeoe+dr8N7rO4KMFbsV4DMrmBYNFH97augw8UpyFi+9emh3IxhZxOmn8NLWmG
g+Mj0dyYb46UAHms5A7DRB1YKLR2S4O8XNhXSlTH07U+y6tA7kmR7nrc3FY4yU2u
MW/ZklxymO5MosZQoBFqEeINgvnVcuAIXJwirZBK3ri7ElFE5qKEc/JB/UJcjs/j
EZGOzmVVVW5yPb3W2aMT47ucSw5fWhEj4fe1hzlxmdHUeEZdIxn74vuU0D+I7gVN
7CCiyQlZxgKsJ70S6IVwtWXAtL3ZDrd7DQge8NNx5xrD/eURejuMDzFJCixEW927
3gBxHMIQDftVudvt80W8ZL7CInUChyXDx6OlQxL5jFtNh0DHMNstuHmH7VXwcIu0
rQH7JZiwNEXgx4v+HA859xTz+lslGP4s0H8whKm3Q3uLiWOBtoOEzYy4Xn6/eLrK
3phni67I0YNFbLg/81FUAptrk+CBezaUWL+jAVTGBh8oL1IrZtKoih1DkzNeoF/1
K1ucNRk5GlItra0h+Oy/jW5mVNgThIaPChcPVHl0VnVxiaFPq2VQdIpyLd0llEc0
Y9857tNi7ZoogSKY9rexi9UlzCCAr5d/Pjk+rs7eJdGLwjsWrDmDoO9mo7RjLZdX
yI97ZTmkvDvxhi5jz4H33fRGCRQmLQs0zMLPAmZuT3/Ml1UJgt6D6e+CUsyFUG5g
ZpO/eEJ54gB5BDiH/A7yt+Km+kGHKoIxKVMrpmdVEgH9IgBec3nY6Dh7GWcgmSdS
8qAQVWsh7YsRxla8dO0xmaQK9vfmnjSak4FUSq71WZOkOTsqKQYHNK11K0Pkym7O
T21au4AiOVt6kMXOohocehO6jqTF49uqvVpcP7UgYONr2z3a+OupRDj4X2AMFJHn
5gDwaChCoS7NAEwWcUVzGdxaeuJxl/WV+zpeFSXI6d9K0vSKce4ntQcU/pX6RFFK
sguuMc4QC8h6GmQEA+arAIGyi1BFw4BOMFQQw1GP2QwUSP8gnm8uj50cbsJhosRS
RlRo7cwV0sYZkQiAoCwRFaqoJllJYZ3D7LbWuCL+dPmsgZWxuSMMJy/f8CDBlb4u
uyFjRfv18SIX2fS4E78JqoMZpBoGbv99H8uYM1/C/ABKe5UpTps+LDwpDA02KlUW
6rvYQCB8qsFreNythazy+eFnBEUMTWe9Y80MFmbIb0HpElPTDxANIWmyYj+EGujU
qoM7OlaIKJ6YZ3h1SFHCVSBtyg5gl6SajHHYK/g368f0wqKoxAxgIxmraL3g/sqf
jmBbbIIq8Wpm3p2v2t81te9U/wYwFy1K1vrH7sPlRqbpz4Dd0aTiSRtEtilikKj4
vhNu8D2zEDVutMF30A7pAW+rC+kVs/pyYuhPib1Nt7cIYnxcOFCJraxldWyF9F02
XJJ5HONZJLvH8GKamqMCbsVXcgTjbTay2mB4Yhb1aqKQU9UuCNfJyD+fivx76q9O
wp+/CSrqX32bMB3Ay4LHX3Lms1EeWzPqjBt7ZXHhUySwMdD3bTfQAcXLjWsN7zsi
QQGRg/cG36z0mm3EWJj+4APPS/dEt1J/wotCN7pMP+geA6/4iJvTanrDSrwSuDc2
ZeplPFtuMjmGcKQd3dutg22z0ZBbPMLhc2yaxISjOauWo98eEo+Cea3FnJLKH2xA
xdELicEPFcj5lT0I0JwfEh44QEUA3ErgrtjFyuBaJDu9Inbz6Xa5d76rkL+hd4Tl
V5wLlRdPlTlu8k9r7jpfzE8Ymch7ZPTKuxUrSGTi9CqR3IFnzKvUyL+OwLF/hQEG
waROrDWUvQUvBGhDQi+CDYE5kstUrOeLsI00yMuNLbQr7nhRpbE377iGRgicFEIT
pfpl1hmtXgSOTDMr1x9a50QjxDTyFMn1NTzGihpWHlBAvgJH3QOOOU4hYaAb57eE
QwRvYRbuq1596x0NMCPODhu8X/QQ+QzvVH/s2JOshElCbOffU5JnrYvskCujAYQp
KuKdPQLAT584GEUY/QTA9eXQ9ubY8RgeC2Vv5OW+jSE+twY6+fs9MexTWoSt9aXp
X5QWrO616SfJUdoGBYf8BNSST43G/wujJY8aPqAez6mT3kVaQYIMnpn/AqRv77ou
wzBx72KmZKUP1qyBMBrzQ8TyZma/QrkBxbPAr2XLjvc+5a/oh6pGOnwtwy0mRDQJ
WvuQs5yBpzNtwE8EnF4z3ba2r8QjIqOeeu6AyZbffANmDy/QvdDT1751xj1J68UN
lwe/VMPF3DPzs+yB0cIQXnXvMwx7HmAqUDw/ioiPjY1Jv1KX4+pWCspuomUVRCLX
RR/0s0PdGUPZyJM1704MJ159j9jnw+g0vSTMqhyboMTUVhlhbPc8XNXrrzm6+kkT
ZxbeSzYrPjCMLefl5Eb8S2ph1FS+/bcuV3FpKkFDFlVKCKjsSW9pKrokYzbp9pO2
N2PKc24UkZqhH0nUHtJcsA46IXL9n+AjR9jUsMS0CKr+uUXM6vfDhgec8WV5bVrS
DENN8hgxHneOUkW5D3wXvTTNFl+6J7jbvLovmL/oNpv23tuvqVaosQ89t+XQiRY5
7pcB5dEeU4C9V+ucIiBgzdXfYP88YZ1ZJpvTnhPPJnlh4tUnP9aWXL1uCyyOzCun
q1j0g/xd8FM/VaxEr64Ilbpse+Txkh7/z8KGSW5B1Tj7IIj2CTCMyIo+HFmqO5vv
ECnst+ylDJY/KjPrQb1VKo3S7jxfTaboafNvQQjIbpA7xSUBcdCw5d7qLVV8uKCG
xVEuQukoJ6owHMB93I2c78CWORVjZCJujrrf3YB5HwihHvZGl/FPVvds2LMVqhi6
M/6L4kJyrq2GiTz7om1MEAu5VeunGu8RtTnm9/Yq4zRi797T1uf/rMl0KwWFd5NL
mBLqoW3KksGAFhwn9/xxVaBLUid0hKrXj0/LFP6XSiv/uuzi9ARoWbPoAVYdzMvo
sV3f4+6I2Wr/fxVVJ8dyqqs6IFyHNjw9wD+X6D7VrS//DqMwW5qK73+bLTbbK+Vp
NFZdP9CfxB+jRNroH+Iw7AzkRVOAKh6D7cgBBH0Ay62mfwO/q1oNiXAFWORklxD3
ANFctZzIqGqoCL+hup/qs3jbnc/FmKEyuBcun94+AMr7qNJD7BDHJG1EIJnwyEnT
g0OXdoMCE3sZoa9UvAYLK8sobub0t234tnxp9i4TjmP8ARWGm0wIIV72ndiOCSkG
MgIxAdZHdIpFL1MY07q4DuFkbnmcCi5RcPXlw3A2vLQxe2NErFglPyhYyR7aywym
cFSEtNVvR6hSgm8Zzou6+hG6pC4ohr37NXArmO9JNakqaHTpAPIog3/+Of1J8EkB
+VSPRomFMcwncu6w3rVYF0+29f8udmda0rmZCXryaFlUM1CEpHzkkQCz8ffpE1/Q
ALsWb+ft943EfvpMQKVRJj3O2/mpCGbAbPv4cFY1/QPwr22xGyIVJlEbae5OwCMb
kelm10s5f9lqyE4GukjAXtcAJgXQQLLcFc/Ww2DIYKMnA0Yk9PPmLiXtO1Zwak55
aRUdvHMdw3YRtAdw6fsWTIEmTZ2bpyhrnwu2eAd3A/35O0tAkghC2nfjN47CeMil
xMjL9L8FypPX4dLKGawH2DwAt+wZYHr7Jsjp9HHa45iPaTYDnUMGjkr/EyOAyTxu
r2eY2gsSfvGz00h2Q0MVsmUcFQNeNY8OwjvGu8aP0f7R/dKEgwY6s3n1/ECy4CVy
vtW6kPsaAkCbcDniQd0fiBOV61iMGsCPU/mPI4NAYe7vjG2HxLsLmOapv8R3Jtfo
xleRZ2hWonQnX/ICkNd5fl17Cz14Q0Oz7Qaa3Y0LU4/gvLlBbHcI9EbdirZb5vRm
pQMqGmJrQJt8H8gZVPr0ZJHTDrW23QdcHiDV9N9s9a9wmFDWatruZWIVf8oIG52o
SiOvR+z08KIlIUOav9/Wy7xPKTP0yhHcl2OCvkcaE5o9aQNtxh7WOhliVxwoYMcD
mO2LvIMnCDvIT/dGE+9S97JlOxcJgib8AZ8SclRHDHXchNo5ZUH7HHYruIR9h+AS
tbkh8HgtUO/E4nI1kYms8rC+mGDF4Hi0BbZVBsOjTf0mN8tayELsHVFg/WVxRnTf
GK+ox4Qh0MBupHjaZsX+QaEsqKLCIyYBFms8SxQQ8Wf4RgkgSokibWflrejE910H
r7uX6xoM6s+pVaWhe7y9qvwOBDXWVFicY3GUvA9n3G6US1HFl4W+xsO+0pvkhOXx
kExFwwi1FxqIFB4iughx/dcjjfuZrs2oV4fECgQRv828Zu7qnV2dQ1XjBPhoNYne
vHgnaUeOSA1x13zF2D1HQpWiKpryG0FIRGastFMN172TDmkVX+5ACsA973xzw1kp
JBjpu1kzmtk0qvVQyJiMQxrzniyCNU/upWvTKvBJp/UqYwZ+konhlmjAK7b4zv7g
HIPTdXr1CVELBNTV8HyhA/cw913mSspuI7kIOSa+vQIYk8NNtMNnN8EZzdcy9P9z
ZJ49oP9cpJpYmPbOd2Wr96QZMG2a2bGzM+zztjCWSmb+cMVOOYFDGsbaD5do5JNa
ICEkVeFfKvxnG03VbgTwSnDm/VzCOT+2VzfWX720F+jOh/TBK8M6kuNEV+pF3z4x
RMDr4RRB75JYeqcNpzxubJQX0LcD5DCu+v0fKEhfNOURPSQmNgQDgyhFYp8vMLvR
xfJWdYJIelhfx1Q9sNi0ARe0zwQzyyMX8ySEmY6GWKySOcJPGOH0mL45nXugpBlJ
cpLErL8ISYhzwi97dfAg6QwJPlAQqpiwMyIdBR7IC6UQchpdX8yccbiStCOwiofQ
Fl14a0UM5XxUgow/RRYVG2CfAoW/yFEL+5yY45nw+nl9R6RP99/EoctNTcMiayYg
t6sBr9b4puJqfybUZZ/Nj6jvYOv1RfjZuZIbKabQPYt26UBNjVcv28doksRvmj6j
9zaj8ntwZ0zGrDYrXZ7/L4LW+Ozao7hqT6cLickfrlRfUJYPs2xoTC4tYgCsOUD6
ERbTsTrerkXPVkXOcOxKS14WbWyIsWPtVMUR5qxfvcl2/RBNCgWkPvqm5sTp+9o4
oTFNhckkA9/VM1kgj+hQ1JKY8+99Tnldij8+OlGyxpRXgYE2FUGeQR2+jzx9b/ip
FGPUvYHuueU12jlTS5LOMq+CXT+Xa+YBhF7p3TrcLrKPmuaHRPqHoR6ZPmlPTaQJ
sf+CkTLPt3QGVxG+5hIQQFQDti0V8FzHXSdiqpop1UM4I+q/n+/9uA4Sa0saPQ7B
NvhoGnpuJ8Vmi2JXdNNyu4CAjkbAqEoVSCnuQMCBpGxckcTRJlMKWsqeQfx6rgZK
dGe67CpmDLrOl3N6W9nZnO9rkBDsjJ8eqYZsp4V4dyc/W4F+I5VnRfmJ+P0cexsU
GOS/AohCEegDdK3kNYSzxSAp6tVI7y2kZn57jcGEsECDPFyHNccBLrYt2a+7yYWl
7ZH/pzz8ti3NIMAG6R4X/bHc7As+9/ogQDO5CkEORNT15jnztXD5YWBMbGf6A9OF
4x8MSE2904GgdxCXnK+pw0MCEFv5DRZQD9nMlT8/2qkkbYyWrvy5XsOTF5RU8gll
mJw7iRy2wqh6S/WRLwOkz/BMGqp1c+5M3SNGqinU2kvBYAzVkjBVbNmTvpd5odLg
H7sTgHVpSScgOdNAjovQqzFB24ofMvss1sKoVXIPsS0VqNifNtG6GzjTrT13m79f
DaqHPM7+WYgjT0yhzubJa+cklJaV8wcE7/Ee6AVwOyUJlW7vULfXTy402ROsOVV+
fEN+Le3/hWf39sHDDab1hw5+8yZPlGLoWrE7PBRolRy427Xt35gYvevwgP6jQGuA
Mz1KkkZhLquI2UujMy48QUMYxnkCuULoNXiw3k+vqYNpsNcsKVMGNnHI6lwZIBCD
MdjK9wO58htf4p4lqJrjVBrWWtDMbfGX1qxwDrA9LfZ4oKIjrMzJCQ3Mn8Evu4NJ
F8ajgJEViN9WjwWSa3JAlPxl/ij+srPg2ZcUNGRnWbbNpDh4038MxEah+SXN7Fyb
YI76rqMFSuZex95L2InlpJjyrpcOyeKpl+RJkdH+ZJSuOFz5MHxwcRdn9m2m2yqp
30w0SRefKe1wXezX+0bXTcm86cIqYhy2kQIEnhDGLhLhgTBIl0lKZQZjsszXhga0
OkavZMw1gc4/3Df1Angv/Cy6FCJV2UHzzn17jNQtAEwLlwNrJ3BRvrCeq7Sp0u0W
LUJuy8l6NYoPHKDwbpfKxYHCRxqwrizv+47m5swVlXgBNky7Kcpswlv4dCHINO8F
S7HxfoSyzjhtWoarhSgVwm1PGbBeDun5Vj7O++zRa8paK1Dn+MGWetPyU+B4Q5aQ
TKEfeptVDlHzgpVGLo/3im6UafHDr/NSu7tyN4f1+Phuf/6E+v5d+aL2CGydXABj
YWnUkQbvi0TDulWwsKA3Sj+2HODezLOPH0UVgVk07jF/osFPQj+UQiNUW68zkZVw
C6kQ+QYt7AX6x4/4i8H6BR1/TWH8z6equu56xT2Kj3ErZE8Zc5bTgZvCiV/ouy+1
bPhZI5gsn2ze8X827HN7oJpkA88aGLMHfJjiaccfRAQ4M/D3zl3LdFcaCMcZ5w5Y
Z8fgzaZx58To6vCVMoFWDCYSf1uFdPev3A1EbeCGVAf/JQzmyouaGJv1i1OOpG88
7xY7CI+5xmDPvlB3o7hunHJqYHoLMftJFv8/vKCgWER5ZeWJ8/1QywaHYcVJRqSk
rDMgIlcMIF07JCmYSK/3/6//pJ/y9gZKjEH9DnOnxXBCwv9407G3zd6Sa2gTG//O
pcdB4ZzOqcIpnGsvRTN51CIvTogG911Gb8wHJbZh31HtCgX+z6/qXF9N70b+sbLk
Biv3LH7hUg9ZrTDs4Ic5OdLfFX9Ntbq5Qv9baHeI6bHdwA+U/jnvCZBsWnFh75VK
J+jr2mvaz35JfbVV4A4H0jzGi7JKMIGLds/yLoAR4J5l8f9/RLvhYm4xtW610/hQ
oVJdHpBs0psfFzIl/G2J9yisGINCbkW4WTM92KgHqErnvXI8hfubQwBqzj9J7AUv
N4VwWaWJQoFKb8cZue1FvFcXzd4wFB3hiYiu3nUM12di3MWs8h7E10Lm7mzMUZ50
Mv/o0xJsjbx9BcxObesvuyO7YSxtEcBSGDMd7IsBYJrtsaQ3u2lsFq0We7aVdeKc
huWwLgv4x0WBKu1lqODTJoMaWXAoPKS7HrzrQjjfwVnhf/4tLbnyNrCuORb3INgc
O/jguwL59FEdkljaPLxUVLGo44shL9c1wXJabACGj4cOyezBbQ45cpm1qpOoieGx
6nFIE7FprvszeA9fcuMvXro349fyc7qy6lbLpo4b8f9czrtZZ2zgGTo1hCvi52x4
xt/TIJ0VLPUXkl+viplp2kLwhHmU1rGfXFpzrcppm3tWxJVWohiexnrU2joJCz3i
E5dkwuU6tcNY7hWaPQW2KmcdZ0+BMCIl+HdsIQDrGAfiqJhq6gUIwPkaFPtmrUZd
3ZZk/Zl+qd5WAcQAEJidlisV5MhOBoR/czOD4ErdU8hyURWWd3u9HYzME+P2nrj0
D83BWmKuVp4PsNgBWXQc0Mq5GBcqXGTdvZC0X1zHGS2qOXdlrag32whr61EEJEOC
OAAHtJuxsmKPYhnPB5FpqUw5zgh3/wHDJBFjt2pqOMvPnMJAq6VUNDHdB/huKoOa
E80/6nrkPI8uPOBAIgUxM54s8Opta22kGLvJq/7r1ntf1AQAt+5YOTo4jxsZSJbM
neBXZNicekD9t6MFhVyiKUH04eylEB58J+axdCo1nol6e2gstajNh/tpNZBImMir
bIBneA/g9tmW3nCf1/Q6AdKjZfKI9y/dVjXiscisDzoD8343cvmCTKV37JA7fCio
qOuJgMgXDJQWM9BFw9eT8OAd7199t1HSAph4b0SvxAX4QPar54GNjPMmN4eHkBgA
7o/bZE84Xtu1hAYLu5hqyc+NPGu/hBr9W8tUPwWn+zUS89kZ97ERLP74fAdQNnXN
SQLvvXrZoVBp8/O1mT6tOYcdasGmqcu8wFIk+U3EtCnIokx2LT+OtbKdoGrd2Yj8
+4eok8+vXVbQOZUJtnT4zyr7048HawfNroKcB8P1ff+K1ILyI9si7/96uFCAEN7E
KpbKqAKS0eDztIljSlzIJDsLW/Ul+tYjo8GTW2R/RH5m/6vosip5mYIBYIdlrTpk
7kuJ1bM4J6bx2HRcd3DDS8hFiRq/LMd/F1jot10HRJ5UMCdW7sDk7AzAGhiGOIg2
Aaw8Yz401M3fKqKu77+MapNPxsuQ1VdTFvO6O8F+ZXkoumWpNl1j2mKd8BE2iLdR
ZT5tpmSg8TaZNqjZXhWeskJ86QQSLblNzPXYlPBoVtMK8+xsk0rjuIlLcET/tI4j
0I8i8fupnjUICFZ3XVQbQ0PjRMqnODKLE7uMtg9e2km8lNNCrqBb3P6IrZvyJeNc
V1pAuycxEC5LiQyNe0xVIie5BSRQq/DrqHqMbdoP+h2+RXLIlUBoJXkebvFkmSEy
2jlvbuHCOrZv+A6aa57nu+M+pBv3/HPxVjXST+3yRynqByTtL2UMhK/PmRh58txW
jywF+zYVgnYBB3/QYmMgDhtLS6ujC/eSO+8kk+XKE5afGuctFHLYQ6OPuNHwmkMm
5EzMHE0anmyip8MZxqYXhVpv6XZI+P/3Iw8jdtIWnr2jABTaBIh1w9IhhK3yh0F+
wJ5TQks+efIiFG3u2/zo6cy5W2x5V6DI/iwwK8gXi+crPpoZ/p4fdF2x55XDgdPY
LD8uMHoZa/eCAaGJHHpTBPETuzwQb5iqZVGJTE+T5PGQmMD06GV4aXX16T5Nv5yG
DjGa0vb1+/j32qhbhT22BsIr308KG5EJgTl94mXUoLU17+KLt0nzI2iNH02s64z2
v6wbQMNFBuCb5/m4NonKvxexRRt1afbDUwVmDI9CMHfVKg6VYiv5XefW2hURONcE
5+pwJlZytgUgUC4GC2/3O0fh356ouA51MsaxcLkk4VXjFeV7OFIYNQ1K5OTLILXQ
8ghokcee/2w/YGr9LYPymmBYqW9ldY0oGcYolhTgKHmHdb1zvfUFRJU1EMIskRz/
38DAO4hkmMgkaF+u9ttF0rKovfwCGBLglzxjbbE1X19uMidr3OgdhwktwhEf7ifp
kG5vF8vtvAkF8dUKyDUikP1SYz1DamUSqZc4vTBDXsLypBXEllnrumUvFYJuXahk
Vn45m5JgzuuBjmDB75N1zhljMkcZRBoVZT8JHmSy4ysIuB68xqdLWuwf1lGKmiKe
IYtkRflybi81Q8IB+QcbIuxEOj5sHXESHlTf+TJi34dK/pfYa48rfj/MTCv9VeUT
q8BHD9AVQeh0zkuJzvSBUJgRMl1I6WqWp49tSaMLmI1GgZS1R2opTE0thKP1FmXh
3ApWNdCj3SP0U4xjFqyGA/y6dxbip8q/qu6Qp3DXrY5iSvbX0JmKbQtJOi7XiGD2
gC5YSV28upHDFe+CMI2tIO8PxTkQiiRLD0fKLlOpC0egrru0lbYJn6z56M8nnc/C
aCxrkVImV3bvOBi2F+s3lkbl1Q+q29dqVblwP0YdoVUKGQlbsn/GdwoJUIQZW7sj
bFsGiwu1HDp6wGH6buNx7fKYJyqiLOHgYkIUxN/ZVXB1kq/A/1g6hICThkl2aMb5
9/wC5kCIH0jJjxR7/d5EZO1kPs8wVxlafyHx5hwI5iLtyjxf8fNBzUZO3JI7LLU0
ptMP7cVhvhtrCJQmtJiVWWjB4eVzy/qEsWKLuzNr9yyif+XuusMe5S5fGs/dRuAp
KnpI/iHuzyFKMhvzwMuOTEtwKUMnS0rp4jxE0dcKI0QJIJd+/3qyXU6p6kaX6DTo
fBpIW7tHrXB3aj3gM6XX/O5zRj6IfEJseAYBtkuNmjAZdWlEpYKfEbW/QF1uj2eP
Hg1VR9PBXmw/VTz0QApEK4Hz15Ypp2z9QJMSuwasIfPmqXeJnXjWi3CqjuRbcyer
t21WxjF3AdysAVbb5MdKb0q4y57LumpbjIdzaDr601+b4yQDcp6ZTNptKEG6xYjW
ZY592O3q4W3uw2hsFeL+pM98CRw/9k0KS3BH2G6++vB7wEoS2LxdVJId/IDQulvu
w+zT+BywqUEIDd81Cb4J04B+/GW5Rka8druhXaDeAqc+n7vYD/VcEm0GOYBI9DGb
hNCwMhFyqojIrwBn519ISXZ+U6VzXaOfou7TlFq+Afs/PTMT3JnpXPrPe1UGIP+K
ErhYnd3lGrsY0y41iKAExiqMcozaQP3IO6+wXUX+q5WJQvAGmRR8TuszmOCccjpz
vVEUumLW+zJ5sz0ZPOSNTrpZvP4Nhg87q5pwi/pNPhKElO2wRZFF4XfeHmlhyB7Q
bXKfdo+MeCeuBQt7WWLVhl4u2AOyV8WZ0Br2AWzHUGFsJ0hkP70/i3YxB0/n9CVp
gneQnuNQfhgDCw71VxkkCAsYl9OcqJjJNNDiuXGjwTq49sJLcc5DQqmEizjgJOpp
EALhw7c3c+DlBz/KDDgh2+03xVTUyDqBqaXhVh3emX5pXfR5xmYjhFtQz4e+EEf6
xHsiHwdmI9QILrHmQHf2FC6SbnpGBY4hiMYbsbokw1nHvWK/dv1BP9AiEOohpYWc
BKTSEH/UQ1+fPD0AEMmgcUzkaK/Bldlc9ifd9Rwql193M7RUZT2a0Ie0s3hGXkaQ
BYday1RaeybLXH0obqzeTMiek38skea3CE96U5xz8qIx0Ks791E+Pz3XqIe+4i42
ELptU6ZwmDzf5Kig4KgEmq9R4B5EHWG+pPIulLVrUJg4rH9RblFvrlMCG8zBa18P
Ss5qNXyeHzdYWIn4HENlBfnQnoyJp3cZV2BPA/MScQsBM8AjBgl4El6gPZ+1KlBa
ZKIHbCcy/TbFxCwH3Shm0r4HpB122dLqjF/8WFPVrr90hkjSCOINVV6opg/ciZ4x
EebOs1e0WjJNAmAPW2DB0VzPHVMJOSORva/AbL/vuxME1Le/8fYBm+s51dHFBhfI
5KJ9ZnxLlppoIsm97W+kowc1rXjMblJs4Z5Enn0RSDjQ4r7WK+j6ruA7ZRl2HqGt
lWBM+Suz+2IC5QCw9OIJ/or+QUKHKn5W1Zp/t+3WaHb7V6/KrEQdT34Hq9f55eaS
wAQ+bBlU45XWebmjbMU3ORa3Ah643X/qnbWPWkkJOz3SeBAYDDRHRf2Dj6iQju6a
DBgCxXuHJ1N9l6Iio6tw079YA4mOWcrdLF/YbkX4Aq7MOb/mc+dRxebxPRmkuwMk
Em8hrOCLQYWECbaMXxGDb5a2Sjc+c9x+Cx9j2EmLurtdj9zRht7HE2jw/RaOmIDj
Qd8COXq3Ya7NzbA0xF8u2osta5ZoxbfUE5CoY1QxQhYlAjhTlLIFvhMsRLuY2JA0
mX3E2AifGC+R8ecMemnTg+UMzNSsDqzsSvqxoOclEGt5QYosmnG/enmewrKcGaRZ
HH0uvtBFIj7eU+t9sg8QCpWg+R7KMnkcwyT5pDJzOiZaattkCOiirm+NsB+AW3vG
tuSBVcIg9T6H0WLa/w0w2Xx71FbfW1XeywGgEk3zaDtW+OuNDZqnXpkUA1+MZXvT
T9v+Qx1LkpYOdXSxZAE8MvrA1UVQ9cWo8wevQeV/BwJDy6DeKLJzGByLFA0ZaMAq
NMHWsbwDwckei732aSwTcL3tqJ9iLwS37CYJORBxt0m5gQAES5wpIgdN/o3YefmZ
lmQOfHBAj2xC4WAHBgxgn5RDCDVAs/UtdlVFeprDl5JaA9WKhVRtPw0GNAwWAATl
QeKyT+HJ7bDfHdiQsUATgTHOn04l/haWKKIshzgdapO/8gTqNCR35Qy+upAAOraJ
878o60EXufJNibo3Gf+W4Ndh/zp7LWw0GIiUqyqAwdVxUpOU3J3W4YZDEm8IScFa
vuaBfDtvdOgxzAb8pnQlLgF1HltRPR8JVjtXYeEEz/ua8mzar9+pUGuvGjc05V4P
SMsbDXgA2pRNDEYcENjNKy7rcXjR17fUY4figo0GwTiRY9XnLeDNoVEuot5LftcM
mXn4BK8HiIkUTUA/Qcv3vXfIDUu7h46Eu3jRldMZUDIyC/G6yzImQyKz3yxrrmKN
V3ItXS0okHwT7YujzDZ85Poghu5vdx/YMtBy9zzYURFYgQcwNAfGzGErvn3zGO9P
y0nFXa26um0yoiQSvpt6IWyWeh+6iI/Gwg1VcZn+VPZy7USIKpM/zUBfEFFXvIVj
EEdAGRNeYy164I+OcydPZA+GeTaje74x+SKXKGUotg9oX3jbNU7o1PT93dEhOTDw
B6KqqmSnrcNviztEQfKoyqb8I54Pwls8z0CxrxYN0ydc4dEXJQjX2PNw/IDbC7HC
zgc8I+9bZLLQvJqN0e/uHVPL5KzAkukA9yGSgbOZJM9kB6fH1QcoDeYbrCXwpVsI
l5iPoBHnjovd8XFIendukaPeFjBtJBArhqpY7dr70++9ORNW2d2B5Ae3BmxXWB9J
O47IT3HxDiEcjAVrXwNJVEZROd0bDtals90X5/zK1v1ids7IFuXkfNVGc5XEXMMK
aZHdPrunRlL1mJw0jVieTnmQU+cCW6SaRUdK17jKiYEX45jD8z36dQZ9Y0utjYAo
j7DqToT0JBjWp7R15fZU+HxEN2W+/ebLYl9Kfrh9lCUtZ/67umQMHGfcdTn8aKGi
FR1WSeZo0BYFWvpm8lFHQv18+rUly8VFmS4K0lX2sQwOvsV1qjv/ld3RrjXC6GZt
Bwt0xsTpxJEmJ8Fh6EsSkDqDUeoqzhKmTqYWNlz9Qt+P4/EyxxuEoykDTH+J4MBn
t94rtQ5qXR3JYWE+FiQWLVyLZEj8SB7v0kB1CutwjJMnuRw6pHWjPbDd1kkFGB0A
rF1mf4TTvwMLDgKL4Kx+5NEYjnhoAipeHszaxNitYlSQ1kQ5tsG2mW+DOfIaubeP
fdHh+5qrjrPOaiLoQy6bU6VJyrmWQEIa5AYcvw/hyyjMgde9oFahXJrMFlz9sfey
jtlxDe61jkoojMLK+XHURhd1puFVPEL+vBjR5yqg6fM50KZeRVMuh4aKVbEohlyj
6F5D9BR+BGfqmlw5semR5B6xx5rloUx4EEKwzqYUlxflVLsw+COBSUQlbhIRdMP5
5HWn7sevTFBsKIUCBsIy4D/U/QiISpVAoIQ7qu7Gc5OQ+cvk+dmHVyEKQDDfWcbR
izVTH9c9oXC2cW1EBT747dek4VEY2gcLpLF0XuJ5cBWSRr7JZoUv+BjWYSFSROMp
IvWV3MZ0qrN8uvZHHniu+1r+ioykuW4aBdpRlU78fBERi/P0JnhvtM8pH4+d1sD/
N3fc3o8XjS1SpZvPLtwfWnMHSXBpTILS9L3NpLkCmE655a6y6cLn/DBV3ZMFjQJM
p4GE/M/weO72kTEPQtEwNJhmOr8Iv0KXADeRbfsxPqE1JrVrN0aw9wLGIdFTaVHj
3LB2Ei8BWaqCguUDBzFwl/44gGShmLCkPyFw9T/X0Mzw8mHsuCfqosDadQDhy7y1
TCp8BYij+qfArOjZlmtZV1OH7FO7hwOWGe1nmxhouJSbHSldOhOComtSMghrMJoo
0pzROWEgiNFCxvzlDZh2iqW/LLQFUbuwnJa57y/GzDTbiX9WQZjSXy5VzqKLrcGW
qoRaIzMXMAMGVzxT8WAixoFMPyGYwKT3eHRu9i9j4zilvJcEBqPKYdlIyF6czaxA
AjjV/w73D8ScNZ2t9dTbrR/2e5DiigNKsmO2ZKt2kSnkWVE1wJj/6urF6nMTs4gZ
DRlZJw6C9EiAaOHe985Yj3Xn0WTzGeSfpLySN5ehJPRPz7WXieFrtMuW/wpdhEIq
T/fO/QoBP5gShPojyZqZElgWPSYKPKGJFNTUHQzX5Tp5iU9EtO3OmufyrHz1A/cY
BNDUFSX4xXuZ1l1cReuZYr+/L3T+Wk2ngq8+f0Mmhhp04VkDCnJgNpBdTNoB3s0P
z54TgRP8Hy/mOAXPA45Sb0wPbnqpxHpNfSXDubyKEJgs4DAhyYpkBpXWX+BG4W5o
nyUNP2DzxMkhijpm2CEUiHejQ7y26q7p3aU0/c6NtWb5jNNHNus394Aj8QxvRuA0
ik/ZL+zU0ARamThnTAMvkM9/HtozoWgfErNLrjJ2vgDVedO/RtRCeEEogi2yBZgZ
e0VFTxCOW0kaitsc01NVB4hANVdVCt/oZEZLoexldMiMOXyl1qqt2jT1eG6lwOoC
b3eG1Xbux3jpQWhpnlLBkaysv3qAf7iBokNWGmxoasaXvhRvJl1PuOLtOKzhAaYL
A9gX8ehBKOK3wBoACyjGWXEyjxxHLloYlgWd7DNTBpxTHGG/4+bu2uRjk2TWHRhu
mNOO5rfl35079u13kAqaqUFEgYF+jnWj2wixxSJcZGs1aW7U25Xo8EguB0vEXd6F
Y07ZX/PuQXHJgd5Zkvx6lnqjPJV2RdTuZuxcsRNyIiQuvdWj0gaD8UCQ3HUXw9It
3TOTGxJhHD91K+i0pa/6yjj1YfLaBr01TJYPBPZG46aR57lsjve0Vdp66a+PUdhP
9xGiod7vIDDxgqcIqBXp9huNAvh5MMVY6CMi4/ZyyJ/sa6FIlzzgZyp2P3Hva4nn
nkaHQrmDEMYijrQllVDE/hx7zpK8RwSw3vqtv6WuuVmnQtucEp0kbnC51Xca9DPi
o3xRHSga7Geli+twtBue0V4C45cjZasKYQ5iyCacIs4qz96OXBbjZ0UAiNpvT9Go
k8s81MPX9KDEPKWyWNrA6CarOJq3yzRbnQJpWBP3AjUzGrzGplV0ueJgAuRgSNk1
DIzEi1VK1h4P9skLU+oC6oZWyR0d2P4DouLf9rUWIQwXOyj27puuh3DFzD3XFA/8
Hn6mTf37Z9z0HnFS5ZxIQY8+WDvhTft3a+U5kZkfY6EoCq9EIiu4t5mSYEI98YWy
TKc0RTjigZj0OovOufEENNzxf/WCBX31pTJ2e0I1nR47RqA+JkdMnn2dkIGUckLf
ANZzNbBS8wD9iynxaC4oULj616OGoDNinFRl41szu9pV3MzrhmqsAMI1zPyClo7C
lV3Ykyx4C15DkE6hEcJaavazyeUAPPfmlDQl2T1Y85wTV9eFwwCLNpaK0Og3UseT
iWp+ViAjqKZM9I/O2T4rzAJG98d0ySDN4rE/2ef8/g2waje1dT0E0gQd7qPbfOgO
g6yRn/1goBBA3Q+5VNUuOZmrYwUnmyuvZQlyowcxYE4dBw5Us1pLUNu0/MCrSkjx
WzMZHegXhQrqjzTvhjc1mMONXqxVl/tpz+WJCfjxvLm5tWn5LM2oG3Gk6hpAd7hZ
ftSQ9IUBDnW1machmIo8rWgrEcH7rsYK+lZz8Z7mGUv2tkUZoUdXimHqfz924jSu
RIkdyaXBjTb81BswlgjauXv6RBC1myeTLo29SelFWVf7Y1T634TgWFW9czacRGZB
vnGWJ9QY9y1vN5BvHPSYBP8xCdthulQPhSYRFBf445QFwDTkFKMPocL05dHjjE7C
o751u5CHYr+Lhg1P0pVXt8MVAJZlsvKamGidBm5h1gFKPI0lPhfmYCJkeHN3aY0w
E/cGObQWt0m+/mnBJqINUV+xwCEeqmjNyEYZDMwXT3hb+tAzM2xjZIUDBmFcobDi
ZvH3bgRqC864ULsY74YNDD2H+Cb0y2rDrIqpfVrktvghjN9PcimvPzGqLxKojGVy
frQOw5kDxhbx7K85ul/qRPgI6mxtblxbNZISbbE35U+i1pZGbxzARGgoz1dtrHkJ
sQA7RrEg2kVnwrDSYsurtC9RTAmv7EoQUhRrw9pJyaTf65fu/Gp78W0N9bVnmTOq
mqlddPfQ1kJgIvqE3Lk9W/rBNCBAhZlou0UCT2TJw1hUTtlsCmipG0V+WVj/F2FH
ds6+HqN8eaqEK0fNlpxji6v1752ngp4QwfDnVa7iIES6L/lUu9fyCu1tx06hViCx
fV+NGB3WNOPFO/04LygOqoX5DGjeB3d7m7udaFBBFJJBxfWOPHJQ5SlLM9dwujMa
ANCXuPYk++o+EIaN3iB1kM9a0QjC8bnMGuLElFJr97W/OU0yETEuOzHYf+NVs1Pl
IwjPK/HKnnIvwyhaZCgQAoFui0uXJ1idVmEmgqqjFyJXov+Nx/k7PfiM/H1u+L/n
Tm3bItpl0YNm8Z4Vy5dJ1Gyvq4OsxbEzwF1aZEBAdorq4lGFiTQuz/lVpjIuM6UV
7A3gDBxmfYSk3ZReM3h2gVuyEIfxK1YSBqkAVLJy8PHJrmecrikpCTbA9KdkdDfg
coOFLvAJutbzbfWZXTBO8f/x7H5Cb1+Geeis1IzD6W6RFFIo4SMSpcSpWwCr038I
TaHZBEKJFt8erhpVpRi0yUvcEzN3SB5nv9/yc0KqR90gkt61I/Ja0zof6wI1s/1O
nkd9064sjLKiinAuTUcTB4WnQrNv9zJx6WM1RitX97isG01gZpL0JamlZzYhd9Vn
x4Osr1XnNqKIRfO7Sbru8s9naGD8lizbqjPsDw+dLIynlOgoYKQ//qju/lou0iCT
ygVPqtwZIuq/63TGgXyx189uWQoucKrz4nvp4H58L6QBtNpFxbmw0sMPzYIz4fT4
N4Vcz5xsWuBqsjmqQP/u3YaGVhPZoAJdO3p9PjMLp++4N8i7b3vqvTEDh91JNkcV
vDhsVvHqAC/SUw+MAd0/lunOLUPLKFqGtFGsE8LCLQs/6kytzXgjHO6h23dIQRCe
R9liL+fHvX843INBUlCpH/9hsdF8Y8EmO2kLf5OxZ93bbBt4hwQ8FuHvDe2CDyay
728U6+Jx6UVFIB1LKuOiqJj4gl0HCY+jemoexceez2jHp+YTR8/lNlQRFEGdFEmC
3XvjboBUSTeJjGYungSOIt37FO+KFd9VqMP8DyqGVQy31scESIN1LfggEH7sb090
Ef+qbzVWGpRE5vNxVzbmMokY/pTDheQJvJMyNzlWx0Qg5zvAEhh2Mzfsem2nTnbS
0o+LAbhIpCBBTSN88j6tT/zYCxTv8gSJd/86DDVPLyOSMTbrf/ADA3ixwdMGbf7q
Mm/0LLXoTVgvU7HaWjZYLbrjbmAKqDcH8pEU4tWrdQWw/CpdQWblpX8k6JeIbIEH
yntgRZoRZe30Dt30moGBvx+qaM0LM8EQS/R/xk0Ey+VnvcIk8fiZOyVF0G6JIfo7
PV9x0KKefd9cyjerdklnsrTWxgjpTkri8PHehSiLgoi5iquBtLRcyiba+Q7A+H81
qp4h7JPp77CgwYu3yovho+gZE2sOGzPl+0CmxqIWpraIyJQflAq2p3kXtWFoxChJ
3YURmzcblsUxE3wgtchoUgdEjrdrP4JTDen21pmzUyVfYHF0Gja3mbRDV9qLCK4K
0zdmayncJ/Jq15XE3VdltBknVrai9J9XTRoyOFJKGyIQl7FDg/Y4hMuF8X1bAmfX
cJFxQMGfIjKEFS9wJ6JcHjJCBzes/HXbvwPaXImgKNT4DgQ1M0WIrD1x7PXj9o+Z
U7gfRSybCJ4gno/ToKgCQ04avy2Rsao6oOuej7+amnRLxyDQLog5PpxnUVa/2Q/I
sZJvoD6NvIfMTBihfUSH0gc3rzhLIUzzyAtJc151Ca3Cvfa2zBhaukyxFyfry495
+SHwkXQa0aGdmo56xm80qE68Osw1dXj3FeyKNzD/0yqKHECsGREEQZ0BjHhRD4t0
EACn9uLd2sT/A4dAEzOZhioXrzZTVqh3NYulTk5SFqaCwQPTvhDls4EzdCni1ExS
rGwv6m//PuhlBCD4ZKD6ErZR4HpV98sk7MxLwHsfCOoepj5O+9V0jcDT5HAIttE7
MSkEDAOlfRmSy+KEq5r8KOsBIvSJHXbySaO/C6m7ZIgyBIPZ9V0ukRuGobxwuwq6
oXuoil3Hs9HR6VQP5rjBXVEkcZYupwRXiJz5yeFT4pXO7UZdXXyOzwg2mhg4ZlhQ
ax2uPB0P4mn7uv3bIEmzfR4JP9MaSxp1CIrS4o4zHyqxc/djQzo3zKaEDTTs5mp0
zFl5H0CMOIZ5c/mVU0SJ03zBZRnc1iWBYHPNKA+QXv1CWkK/J378BHWoBGGU2fHh
Mu73bnYnmdc8hjSNLsIRS4UCYF/XK1/DpLCxpqM+Bm7N8aZoY2vDipsw/Yl4mhHa
Z1s5yL0YIdIkk2p2VTqba68YWpcIF0Lfqyy6NzzjE3xl3k54lLDj1qUl1Qa70rpH
ttlQQpN6PxNC5p/UGScEaByUlv4w0G2gzN8vBZY4tXq6HGrWdsUJjlsu2zvNNJ65
TRBIgr9xLU9iVc5Sm8cZSotZoYTu/mn/qluC+eRN7ht8uM+6hyOo7Jde8+Y8l65m
xcAvau5jUEIUsiCBiRFNlG6NlCF68AsuSXQuwJIRWkko0x3Ju/GIKUpD2hRaoSBr
4cWfH0j2xspmiYwcq264I8YsQLA2skrhspOckOJgvmX8zksAF8K08lMk6UddIvKn
O4WFUDc4i3k0nS93vxyGh6b7M/Ej6q8Eq8etfo6A5kJSnD0Li8aPifUkKuBjaVq7
Fttdd+AfDTV3gZfti5RIKQJBCE0wwcbmippDZO9+YEOyNpAm89YzzWS49opkgwfD
5m76OhYOC3W920kBsNxgJRL0gN/UQZoO8EloYOyI4ywavD170ATd3qoSUVa+IAOV
nnQzN1uVzeDGUToLAlwdBSX3LY2oFQF7d4GCmieJbx8hJsA4Y6yWZFVT/su/ttV0
cSajd4ksEnC8VkDsa+ggnSa5rDO+xrxRMs9hSqR9NhjhvQT7XUzMJ67igv3UCE6w
22hrzyms2I4bwhoVFV6r0FEV1JhOx+HyU7PgqKY9xxineOJRLVVZDKVSnVNUm9l5
7+yyD0ioT507K0RJl/geULETlI8Cf7lOm5UeH/qtTHfDpax4JAhXNVcuJWyWLDL+
ZunvOq5iXIdv8ermjq1csatoQp35dQEhQ/A83k7Cs6jpsl++PqrXEia0rnjV7Iah
w8G/x4dBMjDkOpAl6gl4CqxnSYt2RBfacYUYKdekcAgG9bV36Kcq7p2D3lYYFfeI
WkAQSd0sofO8Gf1OH4QK11whc7byQQ5x8QvK2fQ1icEkbxzO8OeZrSs8z5oZVhTm
/f+SVI1cJY+M4vImeGjSU0VkRsXfDfeJtTHrX4DJUNMWK+CxN+gt6kKdHmqidyzM
Z/yODGaqejvvu0LLOMdJnxG3mPRJ2AmHiAmFDe7zEGq6U1kq6vmATDJ4QBArATKh
qdZA7fAm6Oay20BUB5IwXx9BbbTt/Gojoeg+5j2OaX3BLB/sJyc/J1wEjac1QYT/
hQ0cUv76DfZ2YMse1sunW1G7NhgtmI392lRqW4j3CmwjNIGmwao5Po2DATm8sRtQ
CdZS6CSQqQJVd11Pe2d4poeAfcQBx+B/QMQxZCgmbPnLXz9maoRNOhsqfCimIvdi
2DBkXic6svBeofkJWqWkDouDBUYvYjW1Odz8W+oZPO4kCpmx8/zGEG3TrNJY7XTY
pc5jwiWPLAfaueJMDt80EjxvRQXGiTOWxdF8t6C0KDi64ZoJTfT89CowyjQO8V8M
QAT+7h2zdded7PGmg2ZCMNazgzpSxRhViOBLxADUBQzhdLXVD6y5DgPv2E/vw7ho
EVhNu/LdhQTFimDLXeJtxcUtJSgjZUikR7dUG+r91NB8j1hUzVCLDF1nnlp4OXTb
Bqo3+hu9sh0z7xgw0EsBCGfUoh9KNKMfasLjrb1rwf7X9LUFDNfbegQQmYmjLYmk
5Oeo2iQ8/wZ0a8U01v+FtkxPYY6RTV6xPknEKeZn+Chd9Sb4JxVw6uBKvU+a8Zds
bTyFMA1qOnGQDKamAh0UD/iIMTymHSdY+a455gt6GCCJAbzXnvovslWSeDFWgrum
BV7mvqXDINEiJCmxAoPt5AUftdo9L8uNKr1KWBXrLhjEj5eq2X07FkDjPQEOMY/H
e+rsXy23X2VvbIL0+NRqwt5Qv893553gc2wlPYZERx+3f4t2piWymQlqkfRz4L7B
8JsHqNj9q5U8cCm6TbPfz0WaV6hJLOtmsQSyahpsVNdJRP72fUZ+XVPwhRIgg66A
vp1UirTXmOyx/T6WPvqNrrUzh3CxI+4/TUiRghkjKzX25Hf8OU/Y22BqadlylYso
wbXM48Aqa2tk58AXP69+rxH6uSXTAzD4rJibqce/fYbA/+QEC9n6hP/rKiHTaNnJ
GI/PBODsS3AMuYWaUyeiKI+JLr6ZA8Bwu3/z+C4GKKBN4PxV+/mu7207F1v8qz7/
CQfG0AfMLvGsGBe9mcrgO98ZCaMWapu666QeMxW5Y57SLhZFvWD/Koo730y4sD/o
32/e+fbegX3AyQXyapEyv5VLqC1LRZaEY4ARFALoBXg7AoBZ/mntF1W7B9ahCko7
P9/pzLAEvOLR83eYzHQhVaC9qOtnLHgHVSzgppIsuOovgc+qxHRisn9IoVyPrOpZ
J++ymbrMWMGJUERRlrYa4nGlSjkneK7nvZmfMfHqMii8wY0ipuk5I06ArHSrjaDf
Ph1ry/XoY3juo7eqPrA86pqtUZcKe4sEy7bF+3LlgNg4n2cYYyq4pCSrVzTOjYut
3bLOvbX46BeXXSVraDdwgTXpvH7B8iuTpd3QyOjg10r/d04avN4ZF8C00VAxR5SQ
proKayfXJfnX5zhEMXhpL52A8Kuraq7ynsxofvcxMIeUr5HhEzOATexEZaSZYkyx
jZK4yl8ENMTo3FJZFh3uXIG6Dj8vk04E3IeYg5L0BaN3jmM2jWx0m77lF96E/mlJ
r2NIbHt/qWDNBK1BrgSX9j7OCxYyFw3MjveCiFarR9FF57AEGoWi/B/MSnWj8JIr
R3pHno/w3aciHyxPt+rA/smpGZNcFc/quxwdxcnqCVIyPgE6iryI/mQPvHhclbos
SZvq4wWGJeZFnV+K9k8tjC1qBB29hseQChiQ0MStc9wL4we5YtfNsBD99W7K8siD
Z2bFfxsBR+ZdDi4isD0oADGBH/JT1ew8fH2++tObZZleOfuREqpWlOdP4WbOwJk2
qbjwq8J25aLH1QGKRWXVt8gQLBzRuCIMK6H7bGTtgozaf1F4BPSgFN3s5wvYknmC
K8APkVN3MAt46Snwczio+slLEPnJyDAtVYVNeX7eQh5skSVTYvRFowHlNwldbIe7
wIgf8CbFBHR6G9WUSFOObw3Lh02gPa1hlz/p8mONtM1MvshnpLbvCDtEFrV9AKrH
+uslx5vIu3AU1mjVOB2H7i8z2/yL0k1e3/ybBdfUOmaQmvWwYSat3P84ZlpW8me0
ev6kHn9g7S+abYnwt38m0B8Yw4IpCxgLaEVOK+3kAOsjeii/qM0BpixpPwmLzf/u
KXk9WwNg0GZq0ljqdp7HHhjDrbi43SDxOHZdJjXEZD2poXddPsPdoOgb7zpwZDZx
8DcEpxlpRLWmI9sxIw2N0MbzGKywDQUtiqSY8TV3wl2ohCzeLuLcTU+x+ef9R3I9
FYyfS4AP9HJCedq5q3VXmN3WaWyzGjH7RUNU/gUbcFcioHT1ROGSdjL1+4Z2kUIZ
9LG/W4iyt2De5mSzONZG5yqE5KWG8t3n07IfOVTpiaztn9oZ6N6ZTreysrlFKD24
07MYQlP9g4eVNeebKlvghZHFs6u02M0fqN/IpO2xT9m0dwpPNkPacd+oXRiLuqkk
IBGRv33q89tQWokGk1nsrOQPNTvVc5g0j0DiyoNMLsQDvwMdXXhpUZk0/JWu1cHi
OOXAu43OqsOO+S4SUdc3ZlaHIN2qus4lOY8/oubzI7UbgS6cyPXoyzl+vIjc4SxS
eGUoQrjyxWq6FCHvf1VTFZVyOQGZBo84F1yS33IPNyq3MY/iazRY+ypGzyxR695T
dYno3tDDVCqyAIOtErj2rw9qT+BvlYnTpz8i7MbMoX5DStHFHtKSn9s29JNY2fPe
2NjSpZAQfGo7DKaEmtLNH5GlKJOyQ/gW8vhOUAVRMtn/4a7ByMam9chZV4chK2QM
MaJW6Hkx0mLcpXV+h8HQIb/evJQMXU5lxJb3ENZabwiq7l4YVKwiwB66ZWEF3f8P
qAG0jbuISrJ+0uFU4v5AqKWS3EQ2njW6kH9dRsdL/uP7IMwWRjK/qNYaEX1JUT3Z
vGGYhw2P7qGjU+i0qylYNyyv3tOi3f8KuYXN/1aPqVzQs4PeDY0+5M1DENFxOfEA
0WKYyqoR2r5L0sdN+Nnpi3yd0SB0NEWwHu3fWZoQ7Gj/4C9HiECHjjQoNxPkk0yV
uUGUd/Txq9m9bmJ2tY9Ka2XDCfQWZcVBe6pl9GalILneTAcVf35oiD7gcE3FuEUu
fk+qXULjNZCOfOTSb3alMhcJ45Jj8t+YUokejVld2OwyGLabI7AeC+Py5uBvbL6h
U5OrOGHW03Hj3cHSbI3RfAdf17q0ZDaL8CHkG/ZqPI/QA0dfVY+uihzgb+OX0nqx
5o+1htsdr5WlsfsznOgvWTwzIZyxmZy+JRcoEYag/LDGnYPO6EETaorFUeXoVZPt
ieAT5eDqK8X4D6e6Cm7LB5K6s8NOnx0h/59shuCkaIiSTLqSTtzd9lWmEW3HY5pO
Jd+Fy7Q9tTiajLn6GDZxIknwMndxMi2n3A5g4U9nuxubF38a81BCYqFa7XtpYZBF
jA1iVPCoEHFrEmqA2nT/uU8HPKYdBtm4cm0gdFpc4ey0AHvhEcnzica67fspkoxE
BUDu+yyN7DGbmwRHLVeyL+5PoVGvMeCHp/diXDK2Z9KHhNlh+3brLgWrJtARo8r0
GbmJY8DWRSaSpR4YYYqdUqhKKLitUmE+CsFRuIEwQ9ut1jBddcYv9HvEysZsngbz
VHWupNwC2u+4FWGby4qNMV1ES6Ti/QzI2Ib6MhuEI9cK+eoXYZoVsapGrlJ1NG5j
ij4dJngoVZ2xYJy5/qxOshhHWahqSS5bE5Ed+6MS8LHLmdpLnWu8m9RI5u2IEnkx
UTxq8ATudmD/FxfntVuSkM9ITPcBVUmkGA5tETfp4NiNMoO6/V4T40+QLY7JtJs/
w+pOxESzzstCZ9fpvuU4tFi91Q8naGPkAuQbImV7FtrR1gvyyT5goPoy1EDUK+nt
WDdK5YXvATWbjbJK25bkmeAAObuCcNh3NqwZL+G3Hm/qXMXKUTOMNOq86bibRmj7
U6zXkCtddqLcFeLDsKUAQ3Lf4206BSnRM7Ut1FjPOh/aV4G1s2hyxTWrWiNnq+44
H0R+GD4CEgI/YRxTOh9bfWDunzu/POjumDt0f9bLNxPBZNY4soMg3gRKr+hUw4Eb
Tir58EtlZ+UGDqFjfX84EerG8r/ed/OaRwcuQbaNCkeRGn7cBpxLgYKOoUtmaagf
4VcpTpSnnQfrXp9L7mzIaulxqhG6Xc6pYak831C4/Ddyi14Gq8/2cKSUCPSz2VyG
s49xVmIvIVMzNW6e/6kruK6S/lMT8B50xNF2za2GrIeyFHLdY3UYsG69ypIuRvwI
Egc49iKJGjmp8tSefiXmysYSSP0+atn1NbFssE1W9Xw82RPwYW2h3jpbZa1dACw7
ANl9b5FOcsDYzSJqde7Gu8BBZmhid8ZkXiKEhQi+c/k5IJ/j/NQbbsJGXfkBrnbR
t7+yUa+tzNpROIYMaWbCrtKwLw2vkbSJlY7dFPPLPDt1pOke6ktVSjJGDg1TglA7
AmZRZ5/4pWMRrHiYwx6/Nc2TwqC8aT9L+sB9JDhrDORUoWX9WOJzdOGmQkQGizeI
jMfz4qbQSzOzunelt3FcuKrOO0SwRmm2qdC9ERpfQQGe5JRFlq1lEuTSFs6wx2/z
awGdGXtKcHFP6HlKRa3xb6h9xQ3fp02pZUS96v9DDeiJpkeET/7JBeLlo7/PeY2O
cfQfKdttWKzNaz+dKi70cILLl4llf6LDYYLuJv8KkAYp93Vlz4V+lWFjH/8JB3eE
IwWV70ppYwQD6r5dQ9xM9bNRGE2e85bLinaH92PYf6n1beltFor6nieNrDXsQ9RI
e0Tz5fY4wNzyRWebfuuLk3OJnvqdw3XzeBW2rytczRT23veXzV/S5q/w9Wxcwo10
HNegAVqV9kps1xrd8gOlLOD9NJBvnwKuNS87KqWc0UbOgf7G925w5rO6cpf2hvfc
GCuOH1Ko28+WlglqBgMwxt6A8JZb4FRM5UtAz+bzk/fdedgDQ+LZ8LgwqBMwhImQ
bfNKB6/eZADQ9zdr8qYentU3XUeVy/xCOAWUSG4ksXgOa26MjnUtVCJ8N9czGli2
283LGNXUPadMc33SoBhkxB8LaPdbVdhcWrqYncQyJcHRkewp6ESDN8vVD//bgj7r
O8IWAS4e/081Z9kRFCbftgAJg9ivyuVz5K3ulaRuZ6YLTkm/48NGKFeflOqe96ci
I4kxGMiFWzSuwowlP1V3NyaqsDlYhZDtladtyDtv9qeYR7OfewM6siuNR8DXDDbe
V5kOYgavpM+j89Hcbslf/l7bJhL8ySx1HEE7xhX5KYFb0GdMy/tA/098i7FqUvMn
NUa0mbelEEPadTys93KpAtuoj4mg0oc8tiQ26H/dIUKOhQ+KeaUMdjKrFH29UJvM
iOt461fo2/Y2JaOCcw54+QYIhdSJacVQ50ZMUuaULKqxVlPtaHANfFcVulHuLJDs
sUWC/PDPlg87N3zC2WA6vGDNg548JvjdbFTWG9frrdQeFuGToEMkgYqJDshFwumf
PmYbfpfJb0e/0oKY1mNenl3aQqLvbWI0b46rEL0kD8WEc78YoT59Nd98inPaiuL1
RgMomkRNFAjhdYixY+ZPIMqHZKmWJo7I5GWlF41LI2physfH25wRwg+1NOP3DTok
jMo2OUG/18MDH+UA9tKy3bC8W4wU8JHZsMBk4WV1tQomZwJSoExPfL5XTleovhgi
hiQFjUdFRFArn3HUanXCicqBKL7b3v0B3/i1XzlRtsZf6rr7WSXiie4YV/4GxVvz
V/GR3AJjN0xi25G3IjHDqTf94Q0cD5SgBIY0P78u8/EgAvtaxAVd6jhNnJyDZ6++
uBt3BM6Th5thcnZdn9bMCrioV70QUXnnoTetHwZD0vR3ujYeM8BhRapQ3H48ZuVR
FgSGdH856m44GrhrTowSfILXTX3TMVCB29jl14g8rhpkZ0UW/iEoly5k8kerf0jO
BpGW5TROGHwriN/O7d0XWsq5u7xqUA/Ov2hSWlww3LXg4sfb6jWHVwTlK5EjL2Ch
ZDW4BzT5fh/g6E5OmWuZ6Lxe2HGwcBojo/t20dJSeVga1+Wd7axOMtVouvx77QSe
i6WRbMYa5FHOK2FPPyNe1OXqFM3BO0nLfYadAKI/q/xxD8TWVLoAEM5sSHE1hWl/
keGy5RI18nrXMsjQ0z1nWiatwOsl0fcBdBJGQBAbkj2bTXiirY35O+0DzenVX3HN
EIaO5H4B55OxvWM0tGtr7G4iQcE5wJYZrWu+k7dx5hfLyPaqr1ExPYTfPl+ZavLl
CJ8BbqbkHDOUp66xFdQCSKvBumH01XjMf55R5wiTC2wbmS7lsG1ZkyyyKfOMjDMc
RRgxovSrrGG8WuEaOSb+53sRJ3fe8bgXuU+RTSW41345G+e5umTkmvQHdLB82qnl
Ay/X8k9whj/vsgC2im+jNT2uRddhuljUWQb4dP/dJUZoajYTkFIZBJDBVuqKRsRJ
E6GgPG9x3B9BDQr56aW4a+sCp+cdcW8oUkcegaYFGsPoZY2VOoMoSbanRIxZX4bL
IJJ1OGklM9gfCFZKi0UPPxeGGAaIY3eNPzO97J++RTY/e99T7JbHzOOqxcP/Po4P
7aNuikL4MJqByMRLlVndUMpjkzOOtGDQBfWD+aCOO8MhjiKjY0JqcSjsCE8Tei4J
h7jDAIoHZ7rqU3WUOij/QENh0dHHxsKM/83xjHmlKJIpfA32zTH53Il6F3zG7DVa
kDZKTlQQTBkZwv+FKzYmqcx9nwudNj0jRgptYo5cZQElIG/pQQ7oMOXt6pob1hwb
HvCMAtNRG8XORMZDf7lPznAHZBe78Dbvexh0saM5RAZbTgtHEuPH5B9HaHscWcKD
jGlMMj+HkUhQw1QirHlPHZKcyPTEa3sK58vh7xUNZeViuWGvhA+hD++Npj2z7KT+
/OeaR+BxUi+Fmlsbgo3OL9eilBU18ZmTIaxl5XBwGdQqFy4hTMNY9icnvifYbN5n
Z0zsEjLC6jEe6DEgJkyroo3+P/ka6rHlUuvxW56v18EHWRfLlhIpe4AH6lBCY8W6
nm4rr9IIfvwUc0j/rvQBdG/vvCgVVva2OoNcH7PXnEqc41Qyy2yd0JHgoD0bWg0M
REinUIpBV87wesNrPkHUw+oYu2+5zJcrcTQ2E2/vQW/GFCY9rtr+il7D+HhpNnyT
pNthmqrfueo3/iRRGIYyBBSFq6lxAl/yyR4Z31G5yJtYJbrqdylpAwJUsvoiKQj+
1oSPA06rPz7vNh8SXFEyIg81eI65bUt8aJ4wTDgIdlYOL9dDl/Ws+3JQAU5LB67U
fP8ZhahCbGJkZV1DJfBTfEhcIAtxzIy9QWnhU/xgqM5iMeTCAEz7JYIxVbc4s880
5BytJ6HRI61vr6c+Uqm3XWO470FaJYUA88odAopqB0JWX2+mePVjTth6FQ8rd0wJ
j/3wbVu4GLT/OphIz3ZquUPzjvfTDEKqEl1CKE6VfAbgvT4sa/p4NB7FdQXmGvoi
2AX+j+tYW1MOOlNo5l5Yzb+ZKkvCMTaSJ+O5AWHciGuz5Y5N4dkqb8morrZEZSj2
Dv2aDsu8TsDk7p4r3nxtRJgthU0sdrcHREFQsKPppjq+0vAj8/1m35cyvQ4wLQ/5
7a1PnMQI1WHvfrRHrirEZZ09oLJaX0zk7RL8fJ5pkBG0IPMRSXugNyZNxx6g1hqw
uVv2lcDMtTmI0dee9G50eN7McDxWJwURaL4nQb+8rWs+rfp673jKBgG4ZXog0LfS
sE3Hra9FoZ8hjG35I8jeGP5/i6yRzf9b/Q9CLXIIsRQzV7JZlDh5RSccdMP5wYIo
fj7sYRUgG3roli/IvYlj9uwYRSFWpHx82AWzIWggX6tiTua5s4YzEPWLQrgszM7+
/isvXf1NaCSvzFEOkl7t+Juj0ljBmeAjMRVZtLW+BAOeVVxuMq+BH4/61bBx60nv
flGPmvAEpr+cfxitZEAxpG44L+Jl7u+jfmR6BNVqCqCb4Ftw+kJkMRzk5x3UXOeQ
kKLno0S/5QTQ/kqw3D1+wv9K1tIF9drafhqa0aw8myGnlYDm1mumt2pnc1vXVjHk
1aCIhW8EUAdMoVcrm3zNj7Mlw3SqrqvxFLLZ4J9aOyEFsg+dt0R2BjDZZxHagruq
QSUhBU9/bk+/Hy7wt/1fkuPTFa7WZdI17nV+im0RUvd7aLEjB/By/QWQ7z9Q8vVW
VRtZKzbNjnQO8ouVEz5GMCv0V5pAol0ECImDl3c5iCv8hSiyBj24F2xJIQzsYx2Z
LGxNcZsFBWFSuYB97JQmcqUPv8LfS2ZwuXqpQp1zUanaTyNirkEktVOyLqd8YSqd
oJ2oGH5EaUfBHxfWz9xbpILTOgrh4R+Vy4le6PVu5u2q/4BEz08pF/Fn3HMzVbW5
5qfRvZNXEgU37ffRteXbZPkYqCoS0XNvVJOOrNb7mtdFemcoNTlAXleyed7/+45q
azWijcEqSg5qq2uKPpFhREL7CsovWu/3Ko+3V0jpUCCB8m+SUxi+xyd1ZGtTgdcL
tJqEh9cm8Mr3a2D0aCLEdBZ6kZ2zQ7qIICduGZuP4kndsYn90bAWJrHbmZJfQKzA
jCkFUUdSKCFMNDHhE58R9sEUcEzJE8KobXeSvcnaA3DZy90U0AMGrZ+nVyRWpSwK
bi3+8UFb9HMS9AWAqQgR6Nxz8Wo1/cm1W0NY00qP7uPuhzGpl7YTlMxIcinBw83R
mjDC212WdygUcoIz3yTjmBdncFkWcNWRzwCGxeEYjZDCFheCkvzBpvar1po/5xhh
//wSSrOhgFARZSZI6Y8To8G0TDQfZUAOaHxUE/zNPNmpd7Cd+zae5N5F+Fmk3Yox
E3DQXPgEr2tq0IHMqGgdtaYgXdW18fZIHZdzCGt4wAL35zMNDZTf7qpl67ERF+EC
WkyCe3jl1DrhjxszAxowcGqjr0FNwikUGGu9nvbI3f+F59w/vFLbM4z5281iI4v4
P0tE7u3MIf7ENC2tN6VegbnT7XTJokLmeqXcuhwmf69z+0oYmUjIrS7/xovVjBXL
dvnX3PUyudbdwBJTfdVqaAlBUZRvq040zkKVFdaqhbBxyRb7Hry+yLKHOH3rTlrF
ksmgByyfeDCeIbT1bJbTY21ahxvi+G2iKiJ18JpTotk0YC/yJLcbgp0SKPo8ufQL
EhSc2Ii4TCEgov8eLpzqAmywl9BZxnT0zfJI64S4D0JacVQpMLWBCBGRLAy1Iy/z
rfmUqo650q5VPjjA2f8JT8QlzqYFtDQ/tlJc5ea/ie/g9LlRPeh07zPNYydNnjFY
UXO/jckm7BKVcVX1IbXKKGOND95uNSDUoOvhO+CbzP1WjV/4gytyYPIFqOU40HkD
+nK5aFoz3LL1dLxVr9Q8TtbIT2/y0nLH8+0SFNjsCkR3vWV5noGMlF7yvL4tEG4X
piEjElH7FGvW0i32KLuJmOkXzRcJ3xfLr+6HoXvs2rFACp5VE3EivomPNS1JIPHE
Ega6wgdYCrqqS/QH7Jxeg/CxdA/giQ1k0sVSVpTMJ/Kg3kVxXDSk6pbgygl8uX4A
SBeffo5q/ckZbaJlN5AIVsyH+R2+RWL8FKIQtxuX4cYkYBIaXOuDFNpZHr7x81Is
++clp5qBOsnfwstZQ0cbYuUKKcuh2EMTst/rPonMZxLowHo9GrgOrTlFCu6eHKTe
Pzf4nFhciW1k2r3JmRM1JdegfB6Bi7gVPqqCPjOCI24NBnnyaBErmgSAs9VFm8vX
M6dDAbs+frDQ2Xg/tU/7thC9HTUN3i3eLEstqXQiYR0/nD2VKxRYKbuUERgp6nim
oNcWFQ7jOS9PRWmvTeQwnanG5WS7ZlqeRTT2gqHWoqP/6eBG9ZIeyWw7PDeLz1TR
BfWHiz8JE0QnKDzgc5OoZC1s/HyweyFAsfaWuzqopbocn2WpZ2vFluReh+mbHPvH
TP8dAALkuPjcGumWyH3/l3XcHqgQ3J7bYA6xaX9YxP1SxzKutJhBZeBCQ02DsJs1
azOWTP7pvlJc++RqWbZcjPz0hiUh8/I71BBd5u21J+fkaIAJhxGVlHMAdfkQzHy9
agSCUA1+lqL23HQrJlrq8TeG9mD56t9tw6OxgTCpmmJ++Dc9gjGPsppT1Y3G4coi
JQMhhu6PsJO8zHajQ9HC+WYCwSHv/Q9g0LOomcT3t7XDCvswtZ9DTuPWwCfrhKWH
eMI2J8Q31JcHblBp9r+obB0dJ4pbJqhBZvLZ7SrdAI7K/z6GbXU4ZD5DCmxZBfRb
JwPa8n9R78sFEy+PjX7yNn5qXNtwniWONKCsTuIMd8Q2ZFcKcQqNoQDrSaOLjADc
mXahnc09ltXECVyYiYS9mU0HkoJd11Jl+xfzKyiAmAhW8TYrjFnvm/OtOpBDe8nK
JbzMz8ciiLtrTwwAynsJS/RVcrMtry/2NDYGuBjM9BxwBfQ8qC1pAbSKphUZwpXo
/g/wFNiZQb7nPaQV9aAUGnY/xg0nuwQnLxJxBMdbWi9EkauQHEGvZPH0CDr7ig9U
r0QTYCHo0qP+Ablip5t31fZTlVQZlxGwi5XqDZR92gSjuzxJHrMMBKQb6SGzZZJo
1ZIfY8RMSJiR9vRH3LnK6Qo+BhFUJKPKJD/NN/1GLvMxTe+vbIC9FU0n2nHSVLQ8
Wp6Udpzj8zhW5bKEDHJUh346HfR5FpdS0C9iXLiLrsESWCz54OwvSr1n+7wWCK2q
YfZ5+e6+UlaaLp9NUEPhtiJbV1QaoYQ6aUc4zG9kcuP98vBgWtK+AQiQ9q5Gn0p+
11Z5YIWLJaLhHqnB4W6fHowonjIjUNc/Svc1jRUNDu3bCeNUc7NvdxKiM1mjXoG4
3MRma+2qIrL7JbAodqjwZTQ23fx7zG1DZdqndXZlTW3/q4X83wAXzOJ6p3Bn6Q6d
aY65Tz8CTGTeB+Rin9Y8o7AqpE3TPtWJhFh15i47LARmHYCXAFH2oFucyLgRmCcq
vwvVy3uqlkXvvtkbUxdDoi5AWHsXpitKkrQTwSWexRwjkO7YaXrAxZm3NkO9cxtO
7G9yIkCGtpCyT/3cFhb8Yag9oUzvFHb3dP/ntF/EzabbYnA/4Q8FOPeJLnvwltjh
m/Ypu7jpa+fe5NZhMrzRxDNw0Xhb/RkfqNJSSXfYcoFBprzopmtandt5QZ5wztSa
NKEXzxKekvCRPUME4i4mAq1u1bWBkgv2q0n6WKWs3b15ZAg0IeMeIIYM0lyOs1Z6
c18FBjBvN+1Y1sLpzWvrDXfGsjiBeDsivRLYoLTX7jhDVfgTLdPrsXlKJW6EBQJI
jMZfNcIqRj2k/jt3aV0GTEjJPt+ArlMJOXHboSVqJQo6YszpO1KCAo8Tw+TlxLMV
yoga9HarMJyovn/UlOYe9k7/nY5IunYaA+mIriY+HNd7mMN3fj94saLPakAirV/O
enzimpqMyDjZLzjjm+JE7nGzXgHibocqOu4jFNpLB6lnJqJktVBXZelA2Sa6lO15
5/Gs6EI39rphktoEp/ZZ5wuW8PPLz3oiXr16qCNBKBZtQqvCDalFa+fQEdYWcODz
elD/vsSkKnRLw6VHjtCeBj0b2TQb1ATzyXepNPA6+PV4kiCG3cbz4n5cRrQiZNnE
h5kEIVFlCy+Iid7flv+ryGaQ3xGmPnyHxsgk4aAbc+ZUztv4YCiaaxHVSXvEOjLA
sGKZZQ0q/P+Dj2g4xqfhdpuK6aeO//mnllzolHD3uQE8sP+aBMBelh3DnLwxOHop
gJPiv/4lYZMU1L/ArY4AQPZ9SI70e7kHdLiphZVn1Ktef6lw45oC2ZU+mmmo1egF
yPDnASgf3xiBbYGCLBjtTBaqiw3qNMkW4b0Z499pURtcgapQKUKHGzAHwFzhvIWn
prJWgecGTr82rJsmo8g5/Vl3Y2NPjXQ0M8/wU1w9oAMKRkE/K7KQJDIy4wG2nMFC
bsed4Ops9ksji1rnWWa/rjVsmwZQcPARpNzEIJQdFeuIDZ2/4y7hG9zkMFR5wygX
CGm1sndpKHvUBDGavR4lzZ+XeBCqd4cx/lUshkHX0NsDElXb2flGRJYNy9h168ih
SaAHtQY2axEDExZti86G/r+KNpbc/9bZUcMt33vAfOBNX6zQ6cv5Yi5Ulx6iEv89
Vy8ZnLUPLcdN3653lSN6hCa3gEetcGqkCh4BTbSImd1ICu3spI29/8v7rHdOvy0H
hVGETdhEuP6D4hsg9ApDjrlzx/SL1DnbdtQ9Rx4y7HmVUNLL8WbvGZZy3KOyJQ74
u/mlQMYdHhjsan2fRzfMGfSEtoTcTlkE1+p/V12AA9hDn0PTFS02PqLtk9/TEN4C
V1nPyrMQ4BqPx6tLJo4ompezcoFhBHYBoYQJYP8pbiyMTDScoJMaGIg1+D7fORz5
9BVYcibkSz5hWuCPy4nGGCXwPku9hxby63zPNlnEj7aIM3bhQA6C09DxjL0RmgUB
2Uhtmlcu3Q814/H3rtcYv/qU11D630EULbNzv3VSOvC/wnoX/Mwo4lopEt5AK2SN
APDnQxUxb87Tr2+iuot7ESSFUMVkagGvX5LTGtzzr+PPFWuaczf1AHZhZ2UDBz0n
ZoLFz+dMdwcTCYiXOoXH94eWLT7msod0dOUNECUVC/kbFoy/L0pAjlCGhq1onecZ
2HYqfELSLdPNSRT5grMTWAlhWsehA/QMBtWkM10PiztCU44wt/CCTPVByC3eXztS
mzUtZxjdD2UIhnv3K7/pDR1niyTzVpu3qa/4E7k9sFndnqwr3klIgYCAYr5kxl/j
0WiOzoYLGmAeP4PmQIm03KxeLZEbmEpfKxcOtzRvMFBGqtdWo5UVCIB4oZ363M+5
WF3Qv57B441iasZhdkTozHADA1V06kUe6+5QV2Vx8C5vtCFH7bX4qNvLGddSFtO9
EfOQBhG16ATvNzJ+MZzjGCKe4O0k9S+mm4JhUSkktWva5DQItwFzaATFSRzDWpRs
10v36DPPvkmEga4drba/nz8UsLNedEdnJ1q31DLJudm7GsHlBHf5pIrnJZacmFrI
XvbYPp4iy/VcuLXm3QYEks8mFMOGuuyN0haS28dftbX8Evg0kZBHkV9mYeCkb0ev
qX0sL8tACcY0GfrH9lgPXm5xClHoMaqLH/WdQvILxMrmK4r9FK9c12c/dXKH71Px
yq4mCOiz1yRaPA8v57rIIbLjRScv6RCI5qanTD9h7E5LxPr7jhX8IMDqY6z3Xm35
xDsP8IrjeHjkhIFct+V98c0ftPnfk6OxxsS32drVt0FFS0KHWPeubsNVoid4Is4K
dNWg2NQf36FvQEcRPVagqz2YdJtyRtmzslTEnDaKzd/10kl826kf4jx737Hy/4Sz
yz0ZZYvZ627LhrV7YXNIbGDLO4YOn6Z+pbfLmzY9yy40F/C2bCOBOvVkzrRDA5zA
k5ARQx0hwWBjsV1loqVMAw6933iCT+p6pP7GxmfcDf/5X4HFx5TpUD4L1d1HMVNJ
+VKaQAYbGumpDAkx71IeHSDAYXNHa/2RcbyK8JTioE5LTM7iYLZlK6RP8Nwhc2+j
40VSYndsLrcP9dCWdxUgHjvKimWTdHVOid5WMNJ3w7hP6SUjfNUpHoQzp+oAQUIh
dUefevvShrIEExn/otolwbZsd31Vdhuf4DqVkEhNO/EC7VTu51ztdVeN/ePzJ+l+
fCVibzeZoXhsHzeyem3kAv/df2BgwfgNT6JWKHOlGOSousWGbEZh1bNu69pI141M
vaQ6pvdq47S4SdXrQjaLkQy3GbX0uhPDq+3fbhfIaHpajfXC1FqWPC2QV25k/Vws
/Q3R3ovP9yEbkDkqfTpA9omdn8iPI847646HzYNutU5oJ5+36BsSaCnE6VCPWtvN
GGQ6DB4agaW8R00a5QUtbUpeacuWQWCFFJYG0NQrjq2Mgp3M5r3BC27iNNZV+5NI
uNUQ+oTSNlSoyQr1tJfZcSfCGpUkp58aW7EgRGStVrkTPQf2EtAzDtUA+zZGstBW
Qj1jaP6QXTAChaR0AGOc6eGQ6WJ79jpk9YOF/R0PcY8Nmu5LO5TnkRQt8SsaYGN9
qRE6VrmVRkthcakCNQ99q1dm7EL3PUITOC4NC3BIyqKzMRL5FWUi7pWTursEI8YN
LjT3q9wjJBtgELPcNQfQZ7a8Yvxt90DmBJ5KEGuQtnpG+FySD58SEb4eBpVOacpT
5I37/uPDPFae5KFvHcPiYRq0rMXeBdnoHUza6my1f0AwRwZHUC3rBWNrdWXMF6ki
LBPZwQOZnzcO7mej88RldkOP40iv2jlRfU5pNScc/hNeJp5dlUCcTQLhefd9lejR
wSinuzAwy8x2gs33w7LJYFqnzUYSlYnAFoJvUWzYxQWJvdcJWFfqVT+XkwaNJ1is
r9B9MELuaZ1PwkZuJs5cfsfeh3iVHTg8hSbqCZmN+gc7cRySP0LdJgY3bXyQ91sg
VlTwi46PrJ8SNkMlto+fmimjZNjlSGZSqv6+5iKkXarK9WHUzt7k40qUaqsHPBZx
AgX+v9Gv4VYCOgYSm4Bi5R+arnb6QYiM/rQFnJeaLa9H1kJajyDwOb3iuSC6r7MO
L10IuOf8xyVYh+QJrGdCICbMWH0+mUH4VguopQ9vmp+e7BiSJjObhIrmJyAcrc0t
LUBRff2/YRX8XGvm+rk0wnE4g0fi7T5JU9bv8tQ2tntwbktZqYJ28ykBJhpY+G+W
EuS4W2S8JZXFZx0GDMFUz2WP8S8wjrv5LJfyZWUASGaC1F4SUzsjQT7+BFmEIfS8
tuvq6irkVzSFrm0flDVQGQQkq0KhLp0jGRKQwBToBnVfB9pcKKx0YMT0dWt6Siij
cUNnc2MVORZ1SIyGecQolLteWSoR70PlNl0/uh9uEbluitXmlz6tnVXPdUMeUQ4V
/0GYMdXqbHPfAHJPeMS9hDtmBdlQfJFe18h3ONSJs9ipUaZKxsdOjRi9hKRCv+wK
20EJRUu0h7kRmmtTd9Rg/3g0nQTc0sXdRMTEJJBypLMsj/WcipveWaUVZsbqSeIr
n4hd17nX5h01R7VPYehdxwBVVE4uZcYfoSfxc1jtJXuc0/6VHt/BYpRLgtPWT9yC
dWM/W8xgWYPSnZf4LmAdYVCxeWbd/0M0U7OSBiax0p+dmuS/221FwXgeGJfXAuZ0
HMXiUFSVS408TOF92eITi61tXzIlw7cOWiexkH22u7uhRJ6dVcI1hNmMjkpWPr/B
jOrjFv8DMrJkadEX3gUqmmWiaDQGBpI4BidhC74MY+z+1O4p7urwSTQbkv3+UK73
o+Z2nCSvJPp8FsAUe/0j8Um1loa0F7wgxIkjdzLDcvkjDBdVJzFR3XJoRMt/qrHS
uqcy1AuZC/dcWHaOW2bsgHP7KdL3tOEPb+xP4JNV90YZRpuxe1E/mJqaEuf9cvXt
8drVils5FK3jDJA7JncjymEjBXayp+mDhv5DVrzVpEA3cLgFIF3zeOp6VM7p0AX+
hncw10pl4bCs17C7CEahiGSDfP5Zz5dO3iG95LkE+mpeKlcck7RloZv6KErwNr53
8ucctdzJckkqMZ9u8NRk0aMzu7b1AGhfjS86kfjuF9+uTM/OFdzaFCC6jW8kntSf
V1PksocUvulmsK5nHoMYaKStzvBkvtxxghRQYLNkRkFFl9F0J7/AkziBXEfsgdow
sCQWbNZpLgkJgdkDuH2eNUI+Vq/cFKQ4X6utynwrjaS3iFowYFWKyd+X0xztzIbS
kC5Hoy1kMJ4q3Jpqej/bwX40iEE2Tb+f5nOTlzGoMGm35oEn2T1Ojd2XlA5c+Hys
z2iwSAww6JtAyyZk3IvUoCB7t9sJPY0KHG6UKoNu2zl3KU/6Eqg7Y7gaXHSuYwLk
+E3iw9Y0FrPFFVa+2IVDZYhnbM5FnPHHIPeeNea99JDmo1lmdUEYQs21N0V1O+40
4R7osCU3Q2iOKM8S+x3AqPKoC7haWce19cLs//DjaVS8tGtuCBmwTdOVEBSlCPFz
78k3p2OLwINjLfW4BHfwjiLy/vQlX49A3HAJetVQlEEQvm8283fftvHlDhDGUeV9
M6wZUSaKFNRifRIIu77Kd5rgdYqfr4ujn8wq4WZLiXS3mc9IvIjD4jOCBcPw/HXG
R5kimR7G93bnDBl0xpjTHImMuWv0aqYDZn9MrZWVP7+QZxJz7odPyZlvAz1Fpy0/
cjXTnGfZhhE55piLfhLJGl9uhLCHM25pxpKHD5hwRo+LVs3Aaxv/rxnLV/beLSuD
MRE3vOY6rx09yt4fEMPymYILwnxlNRSvH+EtP+SMHQebEa7/032sJxeY7g3cLMgJ
PXxSumchBuQTgdMFce3FQCr7PI7FrEdMUKPQtI0HSBZIdavrYnGbwyPqlLIpxvOi
mu6kGGY+YXMx5nwPWP4Hcl9R4VLZHaY8wF9jXbfdUUnXI3f+jJZdabgwyr0qUhAm
suYMZidvKLjJDxbCLLpeG0G7iRjBYElVceR/s7zKgn+933YUZLGhevTv8vosY/+C
rJGkhzXqCN0KbT+z5cZb2D+jvWURwVBp8u7pGzqgwN8vPbmKvKEH6GKskKr3YhRF
BmeK0uqCmPWI20C/Rl7MzS2zPgRe6EgyTyZB6/QqCyc/MpTdKwUKHsSuDNyJm1Bk
k/TPsr76NdXGzVqHlZR7U4Yvh2V9FdJAKrryabnjfBH/LzMUa+CIQHoqSmQNFGrX
oKyiLXs921HzKg1/qN4rsMy/ThQu6pXI19iVfVqIBsqOHYpIJrDBGQE1xZLHM7dy
OT9raAd+0KBLseAtrAywWsD8h17/HSnGp8DKDyRijqhOjLyBpoI4C4YmC0IkQPfd
rVwyjR3bdDeolQXt6+55lsiS6eBYksHd8YNgUVyFj4rYQWHcMbz6d7Buc9QK6eTI
SHeLZq0zDfpAatd6ukwHok4Ez65ZL3g4Y9JN8AEBoYRB3+9ZPSDVvk9yPBuw/1jz
uvNmTXu+4k20LclAd9jGnqhx7GRV+C+DYaXplh6tReP6m+MmffcgXZNNhguGmGAx
BmfXS+hn8mGNTo1RMwtsDYHj2lttvmX9YPlFbZ3aMbnAz0ZqLE9A4Qpds4Eklxdw
UMO1ZG7IfMOIQw1RipEYangqjluMzetXxl8Od0oWw3Ao3ZsrgdImbRP22/G5GPJj
3176i5GVURRTY2tE2xpHjP1ZHgtPVkngJGuXiJ+7rBkCtJBygmZURMekjf/lvw/Z
j4b2CXPM5fWADkJEI8ytKYne2oWynoqTvpGjuu1x66Lb0rXh9r1bV/Wvw0xnz1PS
5MqRT/KDR0zio01b1qjNHYWN4RICVYiHo32LUICOotiFuqnIYvV5mlTOsrykFtk2
Eq4T4/AXn3eU/Ap9V6yj8uVBj7kftGMo5UNCgeQF7aPTbwxGRzwi9pU4Cr7QoNc+
5pXUafA2csocSDC+WSBBSepKkw1+m6b2GcyKhjYaFXpz1Cf/Jf4LR2LZTrWLqsyE
BFHQWYLDRzuVIP68qjh1buJEjPMUZ/MxylkMMYZ20ToXUqozIQ8BvYc74YXcwFhQ
Iwr0pFqpu4OpQhCrib5i7K0p4BI6wynMPA+5aUHmMl9HcFIg3lci/KuS8ZRW2vlb
GMnRRaEezZUOaf6gzCnBv1aarrpt+hXvwCa9S6hYrjvJD1FtQ9RaG2n4mzn0KKq8
wlvA8EyDdafu2YqZTYNKUX8rh2u5kj24vqYZ7/EeW9XlF2mXuRM7mYd8N7QJlUie
aTvo9hrveUKAebTvyP56x5GLtipbhOc45KEOXyLPNv0Oj8vIMLDHbNokzn5ZuksB
IUjDeGLZMaheB/K28dtrbiiYWOUsKuc7HbgK3PaBQEl6gQlhudddU7RV1QwAv71J
d3pBGA3fqmjmZG6QKMQbsRCxsAJfpPnXHxPiU5hslOwKU6soA1LO2yqN2z4U52y4
9mh8YsAyMNqOrjtSj4jC9fbjewLrYQJxTTfnQ6bbVR1U5S226EJOCfm6ZQKzzzL6
72FS95pBxiLGSb6HZcigttMpZcBM8JOBs+ZtlIZxeqqjs2K0ViCNe2GRizEwkZ/0
VSy4I7+h8hyhb83H4yXKdW79G3gdpmdlqrsmj0+ng9XtUuIDjVROFc01F3sFFDcK
swgTTEi4mgqQnngDKgIZ3G6OrIKsn+ICfQ63CbyhU4ND50K0evmZXaybhBlDczFs
QT23UQwUNNuIO8DgXE6VILhPKdQ55RZlxPj6BXJAbGZaU4or+XnZqAbvsm3Au16t
7Id7aASGW3NNRcqyflVl2OmYUE+8WyVn+aLbtFrJ0MHCvrfcHiSJfpey95zlLjJj
PUHMAq9D89iTHNQk1SUIkWXUo4N/3NS/5vBVZ3foVaQA7LywJ15iHzuX/Bz0zA6E
CBEFAAAbWUVGuKxp3xnOoTkazf9VNXU8L6UFJDCQxAgLLVBvV4gujcqaBzAC9qqF
icNOv2g+/Yj8zm5rCxLCzanjHu8M8tFIhz0T22yo3wkV+5/dZq6nDwVRg38LpkQl
cHFZyaBP5f4Yc7OTqv2P7J1oE8/cDkH04LN72yGE2+kXdUD65P4wHXU+9CYK0FVs
8lF3BS6Sx9E4oZEn0T5wn1ARz/+g7OJ9BPFTbzYb6AfQ1dh8icSU0mmKSIp2RCb1
EWZWukrIW6lf2BEndL7EKj71hTQyfZPUIlksHLYfCIWygzBXJt4ZyCFXa/EcSNxW
3WEZqmYkwJGl4ZZSVnPoT9QsM/HkgOaCQjMdp8nTLDxGnjtyN/a/WJvwBLfoXzaJ
yaui3dpSud4JX0HbDGxLtAg/L5/k6Nd5qeOxqjUp/4bAKoyCh0Y6CcnXsaFZL/a2
70XebNy+MliHWa8xqpdPr+gok2VwJQ0QEw0K6cei+XyLFh/APR1Wnxb2HwKxlxMY
IoJ7W/UZpsXH2wxRCsfTYyLKTeLdRk6wgomg22jLZqZq1KcIqXsfcTfNU5n8MM33
J+8o70BOI+ZNX5N42/1ZPGH3EyYeNpichUQ+VlcyPhFJfzf026todgOotRzL4DNU
gWwoaUcTQBhs50VnrR2GXBqPZ0lhYZOmXRrArZNT0Rvvi+RSXyhqIt+pn7Ou6/Dl
XMN9pdrrpfe+8Lvb2RXvNNXSQu9YpBuV2iVoe5QtNOQvDS5isWBlSw+KnxJRko5M
jEaj9eZCZ4glLTj5EUFzbiWJhhNaZ1+VgUrG1ZxGt3mWzlU1DUaX52bRJERiX6gS
taGmxqCW+vs8iLa4JiMl/5vLtxsL6e09vh3Ws29f9hNszMicJMtQTSNBdh7t8YQC
XFBYbYH40wuuc8+b0oe6Yex2ejTMcMYILURRumEWQMNNvETGvenE2i+ds4+iJ5S6
pJlJjISvqByiOBDj4lTLJeL7DZrgrvLGe71wTVrX4rUXZHlWgRnjx3VZRb5NSKek
ZuuyTFWpcvqmMvLuwZ9ESw8XI+ENtaCuQGOtc6hXpeOCe8SfFziBLTCXLYLNW/gh
EuHwy9u9nTUXCsEUQmVgCEtPhJLhw262XP+t4e6iOPnTaNSgT5aJJnwOvjT0wv9B
vXYum22xHHURAAFRY3fQOD3w1iOx6ZuYnFuFmVK0HO26K1WtfaJKg+Az8B8wmAfy
tEv5IG4829efvvhbG0hqgavBUKIC4N6EXI6UntCSRw68Xc1WRGSuQXw2g24+T0jy
spo2soGae31tAwyWBkO5QSkwtRMavIkh7ZoVCK44QGHbOHKlbeWANgQ+Y6oU/BA/
4qleyYH4SeCa8G4GvR/2d57UvR+RM0TJpMNaejaXWzfsVSl0MXCYgZYRrG/oZgp4
IffwZ7v5VsmUieIaxuc4YmLkLDnMQKYfT38e/LscNswmZAqpZDRyEl5atX3QHBzg
BmAQoM4LjydKiNhPy/5HHU8T4jQqOW00sJc3ZE/IuFNkooUsAnibAf3NKvAfNL05
o046GVGyvIv/oZgvIKJh5VTARcQfD6mrcJxPwTxALs8BZz8NnDYSGxIVs4hx0IM3
6ckgTw/YEUDs7lVk9VoQmB9zJ3lmKijCiZKtvfpIGDe6MOXNZjiIcOufJRn6RdMQ
Uvtn9l6+uiCNKD5mH6PdjdlVud+/5giWkzwGoGr9cH5z+CCRmTY59M1HxFP07fyW
AugJBTgXYZaL0g4QAQTjrmrlhG7SZRiTbJjKhBnvEhiWe2rBv42m+bFYNw87gElI
5M9IEAIK4KilEi/e0rHkyRbBYMsP9vLRfyOQpAAfTd3F0b2rBN8m4+UvlCJtkH+d
8JopYnO7NYGA9/7AWb3YqEkyDBtbXGJWan+8Z8/rfmckKvsjXnN54AB85rc+WgI7
PY6KJhujB7SLpBAoNQsnVFOm1b/jiZcVJV3ysZ2rU082+u/tKwpDAHjjY05fwVqd
JEUBlB0wLcDJ4S2BizFR5RxxzpkvGKbRIwxakORr7T71sctYEWv3vBkf06iGKneW
gj71kb7wQxshJKDfUQU7PE6sIWWmHpXuD2y0+sdEKv5qn461TwyhAQklZZApXKIn
xKAspVUfImLtSaw3qNKk/6IbaC4fcPixwaE+ynpCHbxSkQmilttDPQFKFroCtkT9
CtiNfo1VAhHXfJAyQYlvx+fBEMxd8xhsO8lyAD3JevkUmyc9szebZ2DafbfjibpL
sEEMgKq5ZXYrflA4cC9sUv9VevgWg9ps5qubYlJ8Hui61lRUpv0hQZHNq9fewy7s
4DHqV5qAVij9eAnefWdahCM4P8YzRGmsgneuu8ksINqh8+kucFP1Frr19thKZlpv
P0eE0LlRMuvl1sIQfrQSyO5pSVBhe8AA/AdS4sxSJk2ZmANQFeq4pL7r1iTqu++s
VA13utp9gKc4Imdn/Jy2KMV/vg4dkAfDL4DJloHV9XCjLSz8bcdsmWcyPa4P9hjc
c1THJ9o9kyLPMlarVAlY4L/cW9khgJI6bQvsOjzRRt2yqxWAz0v0ZL+ttQgvygGq
9cuxdRNkuAIv41nWqg1S0LxVU21XCFnnOJ9zEahrlIpPuRzHXEFVKeN5dnK/+uMj
NK/wJ2wgR6N1gQhAydpGomSJO85tabAiEVPeTR4+gGlk28ivmhdSJ4zjQPBA/Quv
vxmiMiYP2v1M2qroTLJK6U2yqgiRRsY25WwoYszlKOWGxOQ149Tj2rjSJYn7E5pQ
zDVswMotYzUOgWD07ajGjjINEbxPEQdS93Stha9zjTC/6e0f1cnGSJXGwqu7g37G
JbYLUuYdXuXCgsOogG2+Hfr0qiBeMV8f2aKXoVCRlMkS9206Uvted+EsaatiwTWR
Lr0GQOkmaxKon1g4HiWDz7TJJwwDYLRnIM3f2zCBoc78GpLqIHc2/UkoVmFmas1X
O2d7uSJF/g34zn/mxYEFEniO0I6P3KoY1i8YC6JY70R6Niun0a+Ui25Vsxot8yG/
7rbv6I7/Bm+BAvaMGCyA/Xc+ImiqeeeFsrs2sMzWSjtEBW1cgLH/UuZZgtq4BMU5
AvfTDpssk+qQUrUIvPd9KbYlUyvqfSdvegwjLri5jvGzITcaya08EBOgkJidaG9X
bbpThSvS1coMsHWMxBRw753RC42cFy0OVuAQ1okGMZeTEXMGzPVkpKpOh59OtASa
UoLh9tgrr1csygHUPJ3/z3+SJVMOxaP2mW44yE9aW/ipCyDv5Mm+HWb6qJ62Xvm2
kk9ekpLGsjnXdjg0iPUri+jR64Ev0rCON3QBZe2QaPiknQSswftUXJ/frDdenC5O
Rme4vNPt1/Czkxp+f9JkyaWAXYjNqGU6bJCEbdyVtr36B/rClEMR8a21078JV9SO
+A/HHKw6aNmcVhiLk2zqOnDJKXrZwCd5Lm+HCdIiDT9MEG42FvvMJqnel4VRCCgP
koNUBL2hO6FHuJCp4TLNUCVVwC2Xd7+Gb2HMku/swGbRYbTySIjw1eMi1nUKsZdU
XE1IgLyjBakFUy+ES+4ODr3qf0CgT1niGbZZy6NBxY5vX3sP2YJJJld0+EkDyv1D
OtU/L9nXPK9WIONFhZu6j8CoHVSzju+jJtEca5rtaI+wnc5dk80vGzDQnep/+1R4
qUtbtECyYlwHRf+XrvfWjy+8WiCfGZ2TbPqOBqqs5a0EYivGVuRFMamGMoBtBxRb
AcO/34HnnmuGkmY1zWq/BDVBKJNRKHvRJQbh9NbLL+qqI1clcUpY+wBg0ZWiq9+U
2VtCeFXh/UerOvyEKoYSKsoa4wRmAwZE0JnWQuwO18cpItdBsjEZcyzOUMGSecr5
5rf3+ak/7tQZpitrVBJMN3kPMJmec1ANChRKlGnuV9R+7SDVPFq/Q4RGvPiG0NPH
zlUVl/il0LM9dsWN7LtRse6paDdkLZco1Iy9fshwd/ZzEdU556WZU7lpRuq/fugX
IESoIlPntc9TYtd13p58IIRSND+gzOg2O7CZd5ydpCc58ofGQqbOlcZi7iuNAkEg
dFXqHR8teVXwWz6IvPSTVb/F/Q7dIEE1bn7i5wn6MroJ++oarHVMlOuRearLNe3M
6npM+jL1l1qoHUUoe8QCnUtV/cw8mXCE3/2bWHtvJYpKPF0by/CP+6vpKHxqfcoV
pUCyQr6h1/ZIkpHXc5yu9riZ2xAVWpknZVUJ5j2ZUOqDF5L+JDlkF/0vL9sRiApX
z2oVhhSI/d8ce/vGlf6MWebdbS6pVTYQpHNfSb+GtnAoshpVtsu9HcE8Rx5tjcTX
Skw2Pt2HQ6mH7PtHy/8SLOalcn8BmeX99kvbpgQB5TrFK7GpcUUanrwiu604cZNa
BsZsOBJ7+xbauJaa9e0iFP4Fje/KnId6FN3ZazcFTB7M8oBwqSo8ir/1e3mpZcy4
60J4fcyxMcsu2pJNyujEPt7bJmwWvkKJ/HxDgmavF/+YSZr1ljw/zFcaeTMhl0OZ
izZQAx4/3RP5jSLDENYIcf92DwbdWsna3T+xgV7VS5E+DgVoGtl1IIV5iULWNtCN
AkgEYydiVekzYC2gPIGn7rnHdbvEuo6Cunv0DID34dwkFTt8yCOHtZnbmcEmrfMy
30BXkO1pPd6hVibQTFwI/CCiuF+oFLWPK7QxE1+S2SX+bABdzEHYRT2NACSBUEG/
kr0Y9Xyw7J+WOmW5hicxvYY6rfyXmzdDTmk8ApANxSLnrzmdEF7K4yzJqhg8PPJe
5Drrq5+FDYB9kkRaYKfwd4PciuUqELB/FWlfp9Id1CXpHDf7xT7qTyUkYMovm0Ow
xXhEyodnmpmcnF2IsW/Eob0r1KpxOxmiGMJ/1o+7VOdd+uDYVr5V20vJydEIu+99
/ux8iLJnPXAeD6UCZILJwf10wYfd4KFJQp9lTxYsmvA1FGCjo+eNGUu2dx+P5nnh
JyXLYplJQK78dCwng+vPgDThGI2JI13Feeugd7WF+PKFUFz3WjofxTDKfA5tMw13
T+aALSkPiO2IsMwkV17rp1gvWqSvUr6d5KQml4gOtWBn+mdc2KJwy6bl64XDTzRv
Doyo/65ggEHtVOCzmspNukL8uSItrAE8m3VE2HvahDPEsh4q96cmHXE0qTjqCI9j
o4S2tNKLBuZJngt6HEa5WhT9pn6ZCw4eK+AVMHYUXmfiF1EoTcO8/vWXbw0o543C
r58E2wL478iZralXv6TJjajhhVnRh2nKCpz8TIUCXN8mlnc7ffkOGXnspdCgsXy5
KlfIZfjZWm9OR+IfsSVTtdVK82JZZIPYDZYnU7gf6gsBxKbd2S0PIlVUzon+WtB+
jPvaXH5/KC/gmOsAUiiUISRIY7Mu1WOfr3AydeVLGonSe6yt7HuhJzbtUW55MxzU
It3w30a+IA4lDMDh0Ug3SH8CkBeoK4Z8f91xaRtlY+jnINtht1SFcn+oQZLsnPP1
foSiBRCUmJYxumrLx22FGdXHdKP7RYU1eAtbJZY1TRaX6twwsbzc2cl8YI4Yu5V8
++F62p0KZsLNdeGf6m78yxK2PJ/wNqfpw/a9venbUsPNkNngFng99BxOiTjE/pPu
dmTLjBw1ldX4b1fTz+8+YPC6Dy84vjCU+nBl42Hskoyx3H3LuBjjW5BNlbW/Y4eV
U/y/Ja/nTSvrgLSAbYZCgh9hbtjDvzdaLs0J/ZTLwtimbAIBsIEIZGXjg8gN9+Ox
YONqS3Qf0jM0YKVbDBsdnsZZBkDwkvysoKKgoAFZbvm4t77mP4BQM+RVAubdFW13
5o4uTeE2tukBofdNROIvz6XPfpu19u8LN5GzuGJ+C3DFfS6/QrY/mJ7tqeIximay
mxGFOLzfNSosPY2tusD81gxaAlpUoF+a4Av0nGZ5Yxcr+9DNEMZhFa6z5ZtPgm4y
Wi29oroEEYJIOe55SodPO3B5jdLfUSLF5mElGv7Heqhu8an3Y9YSpKm1AfBFCc/W
fJl60gc5x3mHT6JGEtILv37epQCzKP7uDsY5Jl8PdVtp6RcTCBA9TUiv1pSLGd18
nMJm3vuhcu9ijCwvvx6BxWXWsU9HI7Jw6ITrBde/Ne5x0pv7u2/P3fdizawfhgXL
OPngmBkyoJhg3paucIgYIk4UVQi0dzVBIhZwx+rmMpq+k8dzPxtdBu8n+0Kf0kgQ
FA5FyWfvQ2kHrLet/ueidjghcWPOqVeEYSPqZP2tOD/ZXTuRa1ItqVseq+8sCl//
bAW5VJX62MwluXpKe91n3nsTPYacujGyl3Nj5G6N9Ahlw4caoCkOjltekxR0BOBo
Yta8F/NnTq/tBHW0RdP/rOaxbi3UZy1gZGB/Ouo0eCe5gIBI44p6euojXfzof8Pz
LNHX64NHpPvxm40LoxqiFKp1v6tJlb1N5/0TgBoKcEY+8yPpneH6HWhqA1KxhsTS
BUpUtVcXoXpTpZdPUzUnmOJI6v/c1JLbe6F5QhBHYI/1ysm3rX15lgWwWG+/GZWS
6fLx0oGzmnietBSbZ2/W53RjJYGB3Ne28SI65QBEPHIsH5c9X/wU8dD6IJEGiKUd
PtkaKdnrrP9odDvddHTXn9GHU27MGSm8YqKoouSxV90lEfI1hmPar7Cw38NtyowD
h40ki7GWfVm7lpGDIMOh423rxPh13tBrkH6hc7Z4s2sdYlYLX40DrNTQ8tHrs5bo
zBYLHANEzOVHDY/9cJizG2ep79+Z4SburRQmv51LP12IfoC0kh5MSNYjk9caWJCv
wFUNXajEhdSsEjZXyc/45LTI7xhJnO7xXdGzenwd2f2A13MouC96N+24ZOg3wBE9
UR8epa8Ksm1yuto/QmZU4TJBZwDjgwMDMNOpRpF+t1ufqzVucG+BRRP+Jo5DCQtO
ep90Ih2Q+aFuVecxgh74EeLhxBSBO9SHSuP/pxlkt6AcnlS/ykzi+XmbRB3nsqdX
8JkUZvhecNkk5+cHGZFpiY6HDoKGCNBJ8lvPqQUsyHE+2u+iGLo2MN77XWoMVag9
CK9OHF9aLQ+WRZcd9KzynDQwrlLeNSnP22Gyn8pmkIfJudf9yamgcaJ3HqlLfI7s
htKQ352Jo7FK0Tx28OqGGg3rW4YNRMs+djqJmY/TdcUSqeLlb3xny8LELTtt25Xz
jlQIhbhBrqZpu6pkmuojp1arhLL44dB/8n13kd1qvAqUNiOElUqJOzAoxz8JBP3v
z9KkkgHKj8LhGDK7bOHCLxhucwgoZb4O5jBVPsV1pw4Jp56XvK5Fz/rltasTOET7
Nsdje8fWeaQ/AK/+WSfj9X3tNBsAMKf76AdffQ73sNlYpju/PqVE2bLQIbfPEEer
Ce8bHYbsDBLthnFVnnXqYZYQ8AOPBslLb55amjzTdbo0aWvbrbMf7RT4eWT8Ba28
wqD4kYqWAicELVgUnbbVuRpI6/9IOUBMGelEbA03dC3j/YC5+fnyuvU9lmk15zEJ
ijXwEw93uQ/or53cIJ6Hs5zlsXUhOVQ972Tm5Qn83Vo6ZNBU597wSl5qtp98tRu6
W11baadJ/lKUkb8aPTL7SJmC9qxrlHN16mstRdFaSBqVY0kM3pFaPmU8Cq260r8X
AZtAvRSHAqFgdGrzKPaBtgaVdY4vH9d/Q9JIVwc7RkF0qu0c5V20Cn10LPxyutv+
Znv6coJSI2odRSBPM/LaUo9GpWeQM/+6vzpd0P2a86+CDb3JNHWWX0NFXAnRxMMJ
7OuhpYK3ZAl56N8zH1LOfdAC6oT+qRBprig26vIrauSeLvbUWZnH1HQynHFs6jMa
8NcMsYjn94D9VEJBnAQChkXL2i3sdFY8CSWvgpwXRAprfM2aVhX6Ma8H2MUJXkNi
0US75sH5MclEAqjW1fPPraPyF+rcQg4p8EHyokIwVfAYNusaOsZ+ZfXWLmVE8p0G
O1ASevATu+/CYKSsywM9yPin9u8SrCTc8/CO3kw75Q2ad1Wenl8ZSfVWjtU135KJ
EVnePW+myDEZucRnMC2uiTglwctmqhhb2Obndv0MugUVNop96DSu4v5iSn94PGVK
eZjLC94DUUrKHzQ6PIqixrbuKMVFJmvpsv+Pz9bbk6QRgQWxFn7dDVsJ6pB8XeGY
zUdI+oxS2eMqhOHyvcEmbWJRf4X1HmIH2MHOVqKlyVuddvlS3H7kbXVOxRURYYKg
DlsaRKT0oTUZR7AJnTM/BuWH4PgXWDgi1wGuLUY0PF8ZB1H4q6tt7ffGcZ1iuiYm
zR1WGOlwphTsfVvgEUB1M6IxBnpWaZoweSdJJSIs/wceDjTd6ZAYZSH5MfShMxLO
NvE4MlV4cmhPtw2h/HfDHuDwpdxLejuVD1E5/6BlDwv+TRlHqYuqZnZyQHHAZ7F2
/R5DeZRktyywc4gFMW62ibJkzNDgevK/vq80qUwVc+mur4h6D89uXiD/fqBcDn4L
xOl6Rqt4aYqvyPxMxPSDe1wzjUJMDLQuXHYmJ5uCm+Tp84qk5LLFwqHg6C1SXg+c
w7dxxxfJGxFdGUebmkysFZwybckV4mc913upcMf5cC42P0hvnyaoetDG1YNuxoYg
TjgxqWFAW14zggwRJpouDcNN0KuplUaIncr3wiCm3F5a3Dm0qnsQzP3MWzZrnDZ0
JCmUbX2oBKa+j7kwCHF8JQHNH+A4++BPjLNc5Qqq0KNrw/YxmEJlgV2KIdMn+zN/
P9g5ertAZ4KdWOGKMhfaTBYlpOzAQ5vor/4YD36kPUSjyGcD5D+mj1AT855StnG1
uau3wBaVle7hueccwcZVWF/FU05D9dOklYz3A3IDKUvIJEmK71Nz66BgUXjqi+oa
Rex+8M1xy+FBLQMyJWFe0xdaEmk1KuCql7kFoPpsK+sxENYLi8x7cFndcPQWzYfD
oRV4hFUKkWB6vT8vFMEMtHItKkTqWcsah1/q27/Y/wJuKZpIgRvNzc3KPk9dCjoO
DZ3Rwhx2SscFKZZUeonyKV4uxBNl68NrtJElb0cmemrcIQmb5kWdIBRpxmfZHktO
+/GoD6JI7S12iB85WIRw4rxMjFhZ1XQ/1Lrag3KB7gTlWUeR5mkTlvSHrYCUShVu
ttUGgxjcXZ1ltgLM7FY7C+nJ3zQBmWw0gN2QsOo+euWuOgdWy7D6CLayRwlvBteG
xWZl8dq5tAAhHafwoCI10B0+t2BV4IH1D2ut48QEs9KH8uBMZ7YZzFwEeBJaFdcY
og1cM+hcpLPwCYsTr+1nreZnsocvBCTwCuUAUyHLoWQasYm2wplI8iDO+GVEj1KG
k2+J2jY2RjtCc5e+kCRNA0uj8OrHHeIZ3Cg2Ad4BWcpxzDHOYUIA5zR4MpgtSPjC
gtfzDWCGMtDvyPBG/uIod6MqSWMR0ZKJlAuQDol8r+B7dN+IIG7Qu19PvzViswTz
pn6oFv4dfZ393M1RBUbHSkatxgSXSwwuP+GyX/oqKzTgYRactPiAhx6x2cLmwiLY
R+pOCfUccihiF4AiT0u/0O2kK6kNymYbGhSKABXchmY3SMVFCVQZKs2+CrgGgUpG
Qz6/bvcQnSnLO0u8uLg/3Ov3TToh6MeiO6MXqOrUqg+PYzNPt9+wBrHlyNibjWSW
vTuLZh4XrREmc+3xy76iDnjifvCUi17k0IYlIYiBwspps8kctN2gxMrv1Qm+Anh0
DdLoSmc/VOcRmZOf812pLzSr5Tvz0RTgd/nQ6Sbz+EEJUquR6D/hohDow6OJqqaI
ddwlwRPnqronUb1wnDk5bEk+4lEJ3gRS7MwGXPil5xTTegYwwZLFoK+om+pbtTa8
+vqSgDsO2MrXuxdg/pnc12P79d/45uGvyhkFRUsl3R+0/fg+PzSgR6nAGdNzaz1G
CT6mZ5w3CeZgSqJPSlb8PFm7HdXpEZv382akMCsU8Xpp+dLYOULhxCc2/9IujmBb
CXIGLgPVx3bfwxXEX/0sWqu1gx0QwIcWUq26QlyclUP2lidzNtJdy+GWdrDISH2G
4Nipeq/zeV3LKgv2bXmDw51krqWAKO2+S6yL2TVOPf771AspNmyGm64QD6DoYzf+
+fUenVndJgKRxddSAHObul0MBHPEIaKzi+C1SwUMiz/Cr7q9kYqzqerjKsHxjTBT
QVQ2WX7qS2EiL/Ptihb7xY94Q8x9T4JpcFjGIQJUL0wfiexS7jtzcpZnn8LLLETE
yzCnE9CbHhr5MVMvjGucosYYIzOcWbXZvdSF5ZdvlpKRKTKPpSCAl9GZy2OcqqDI
63OohQyvxYZ1n0ul76wRUp3LRJ8KMVXIOU14ZM66eupniGR5Rq0azFqkK5Ay/uvx
5aK5dqE0yxLi0WVOLidlDbPGmxikh0puzNCDtPQRrNuGggKfjP4MMrz+piq2Mel6
F86vQ2RX7NHpbNXL0TTdtj/Ww/rpdDVP3sfIwE/4+awPSTKouDkjFdiZEWN/e+vM
TcfnT0EZsJBJIiTuByKYgdT7T9mqqeIH6L5ZWqr6XxX57cirQa/IDFzxQfx7h9Cz
HC0btYv5aO3cQDod/pwhlHdflN0SyJ5i2FtPDiT0QrQNsPadlzpsgfkYoPYwjYD+
Pcznf+bj57EQCdRuxLs88WhO6r7j9AQTYaQm+EjSaedf+joby/Lp7yfax+gaAE6Y
8KYZa9s9H9h7fKMzNeZe3gD0IUU2XSSyou4Of+e5ktxHI/u/ChzFZXNfWNXgnwrC
wRznn/LQXeJA36Dhcd/NzdWMOW6RrGiyTXVsgxAFf5uqBg5dPlvAsMCuKexdpuBC
+FmqGJI6eHGJm2pDgigiX7BA5JRDCTNionjiKK/qmQDgSD/mYky5nsx4AeaFhgwc
cBW4VKRQwx/qYUdP00R85r0mZnh9Y2XtYT6vrtO5ees2YBiM2d+9UKYawfG1Utvr
0SED2Phes6VIYX8RUPUDYty2psWznwuBD8CJJn/ogLlDMUz29/tXjK54e+ZVd3y0
ZvGx8Ll+CqH2SdH3LMqb+vzXxluPs+fiecBVAR0IUSUhrX2YdjG41cB4xRaNtao0
BI0RHbuta4696DheH9ioda95SoAdfZXQvc6B7j+xL5n/sfexELNlstvwVNYGlEb8
3AJc6byJFlDwwBx1IktMpwI2l3iPOJs+VyKox1rSy68/1cM7YWOZdOLLCsIkjKRR
Y1sppY6iAnzZJA4ycuYcSGEIyK9jvrxDEjRdrkK0NJsPv1ItTSXks2dLS8MO+PGK
NEldcNp4q0823polEYgJWSBPQbp+pokK00BpUtkzCDlThBce/3ssGahOIrSkqtvd
jhtlG3pBvnbRYip6wql7dsWH/RArdCObi06xxwAQ3eyf+Y6vi6CBjlXoVEirp5oR
iVVtR+5QyNzZ4utRuJ6e01W92HdnGIL7NtXtMGu3xyRt9NA0L8l4KXHzHVQ7Oea2
B0III6FGfFPg+8W5oMa8daRBeBarethDkx9djEzxQXSvXnUMDL9tbjikV0Cna+0d
7PON6EBC32UB7+ZKCy8SwzFqV3a3pbvh1a9iO2T1aMFrZfwMQzGr2yc8BzUXX8iF
UmQKfRW4rwqjyl46uQKazff/Axwbnk6QDKpLDH0Km/ArMPMRw72WJeeAbPuEeDys
JSUNoUAAJ6OJxcfpRIujqbbf2G82UY5jo+gISMcXqOTJ0FQcS/rFiLnFJod6stcZ
6pt7md8AzJho85874UMqVOgVkX/3t/6UWRHyJqD2mmKi2rySh7fy4GfcplrPYBOJ
D6KlqgQgCiYmDR8GJELlyPPhV0idbYRSZeP2h3ZCpFbM/gmAJmY+R+YqbBYaA/oh
bypgO0uFalg7nTjarrHxzex1ASNU3Mzm09IUQgB6nn8cEbTFXO80935v80Pt/MvF
NYj/ZBJE3P99BHur6O+OSbcJRjYaX+FcSeBhWG4YaXbW/x+1vKeAZ3H8P4RcFZUg
AfG+oAsJI+kNkbhCEtkb2AMhVd11To97Nikw9JvOaJWYIuUMhWsDfDYaHgfUqkJm
UdnqcD6VhKqbR78MjHRJDOIiTijNtXLkJsotpb45o+B5Sam890oN4SCFjHOISioq
UYx1PXnv/gInD+B6JzmeT+hS7nGCvqOlm5KOk7EkP+H2f77q73XfOwTYjYggzKcQ
kd4HY7AciHQVE1PAOT7ikUrv9MvR/+BHtDOffwOfJuNz/bQiKYzOOaAEejLQa5I/
6uC2sLFP8bfHEsJ3W6Bhc29BXShBab7Jv9I5GIeQkC2s7IyeYleOmpLcHBtRq72v
mVGH27U9e982v75BIUhmoQkbUhsWH85b2j8gKQuHkoq/MoXDt+rIPPBy6vmiGtSC
CGO8pw8caTo8pQuowltkW9zOr3iBDt/5i5TTMtELHeTJp5mik0wfoz1CK6RCFaH8
LLZ0EO28kTGBcxDF1GD2v1kvsQUa+UPrBKM9twwJJeTzDCe7SiexC/ZxtX2US1sk
BWglV2QHXacBIX8gzlq+Q57dgiEyGOawd5U0TxjIClQUL2XtfYxoky/PYo1R58vp
US4pZoi+5hsGr4Va9mkE0FMG4qZWNjzMy84Xl2Lum/Ip7OcUr5qryP7booRaBGZN
Hy4JD+wnfSj8T3tB9jefOHvZvdnTkoxVplaNGz1rRLT4ySrBeGiUUAICYDve8DQR
6egKQXcjv6Rkv14CVcqpGMSGHsis4OT5uhaux5PKpAdBnA8HaWOSmgjlfmioVLaL
tHrC66pS+QmIH71s2XSrG5s79B+0E+wtYqGqjm/qvY+7mUja2nqKquU4YwrDcZm1
fxSJPKjrQi2EN/meICkp4oxAOuyeRnFyp7qbKOUp60SNnc1kvkWzY/IyT+RnGVUi
4ToHlATauT7FSzArKgu7YcRqTQbOIeTnRfCpXuQmGBuz2sDxCnwf7SlC5JVMdI9i
AZ1h+0PGFM4M7qgB9QeIL+spddWZzla/eciaNqs6S7irdSrFagjxMRIVZFJMwM/E
GyNtzhZTd9tq1IeddiZLWvg+IMeUEAK6JV+coL/ct7Hj9b9FRqzgpAc5yb5nG8R1
FrCRejwQYuXHjFzjvjI1nxbAioF+9HNz6HoUPhhl23SimkA9pZHgcE2WkX3dWqdv
crzboIAMUAkyVrIGsWbNh6N6N4R0Id3zlPKCgcIPDsoMVa2RCxc9lAhoRpJemNIN
jX53xFmdlaz6wt8re7jva52PGFTh0RFu+6+vSQEpyv5gBwmB/QnYgeHfIkL16Td8
DRuLSD4byxPRiH+cQ+l2Kkw57+Zc85wI1Fe4uGt34BR0uUJTK6VJGtVGSVNGqMPb
3zfgUf9yNJJES8sgM3iGuf7u4AdXwrDSPsMyLcJ+qtfXl7mD9Gx12DJh5EVOZ43m
5f8hAWLmeF0h97yWXce8UWNHo9BxwUI77Ra/eYD1L5yYRuNBrmLJHXammSODZVja
61vsw/OpmM+Z4ZkfszuZdbmqz3CP5gwrsiQ6KPjaXeJEcxQpvdzb/mRBoFo2w0Sd
ZuAgB5sX+Nvmt1/2SpMNbus8K1OeKCkj2AJNpj1KVhsouvzYcTz+M0+6lFhXXYbH
3HbsVnBcoX2yiyt3Fi1quGJl/I2PbrjUqkeq7M0vZLv5aZMJx2q67IM1sLWmtC5E
NKrXzJ9Gg6sIioZgWA6X3mDJNeheM5ZKEcbRwBhs/W0Az/NyA2BA8cIy/W9Q4RWU
6ebWayEOAYgi9tIJQduUuZjsNipuNTm7bBUrndnHy/DGQ20gCvbUvO8qnrQwMlFO
cKA1zBci9I8hFdZGsWMS1KxAuWIfknXw4nl+WQa63WmfqWPHMBtCLN7jPQBdkzBI
r+CIpXQnluvFMJMP6qR6QoBn3M7L6ihjm8xt7gVIHB6I0i4cZZzH4HnL2jochazI
kY/Yqci50kvVMoEgRtYBMdh5dUTzUMNnn4/Cs3fQbByFiKCwBebxTUOEOcxU8I9F
P6IACq5m5k3EHNuKhYYtZLsReRoI2LwlaTPbUQKLCNh1CORA3OpS/h8hxz+STAzN
vxMp+w12IdEiPCwtlFC8naFQ08KcLJBjTBjQjnZjQElx4jpACWOyvmWPHeIA968n
HV/ojjYHt0Zq7exvy8etEaDuR+QVftMRAw86ArLi+JRLL+NiO+DwoQB4FD/HpTvY
gSYhNJgiT3n4+00iqXnXCIW27nPn4+PSqeUjOsE1rSCZKgY27/c1ph8rAE46/4/+
Q4/SiLSfYUgO/qwNZN+tO0nPXlatkGYOMkqci7VkFn+FpeX/1ekL3qDrzSEbNcR2
b7tbac0DvMTgDnrDNGhvA7MWJ/PDVcbsQCN/qRRrO/tGkcaVoouR30jqYhl5K5FU
e6DGpjhGRfvsGgofD+0Qow3obCo3zz9AM7IcTPK4gk14Tt9+FlAhR9UtZeWO2+np
5i4FlrZChIsLcZopFRj3PieNA1uC7H0DNhvG8Fxga99Bls6QGFg86THZcn2CpyGM
FUgG3rRXoCm4upS4D9+dkng08ujOsycv9AShRM5pUTtgCdQg+bFMAf8RefaHvL+D
AAOESvigZF6UqmN1soqWPTKBNzxbas2azUTz780/4/0ouwLQ42cPLk5fJazoMWq/
9NpHAh3H1jS9cxZoOw4GT7q5910q6iAI65b0FN/kZH4TvHnmZPveR11sOoVyGZ+3
3jAuuXs45lFOW/bJ9lsP+FOD4YEtfdvmIl6b/R3akJz9X8HrjNWtpVpqHiDJQAdO
6lSuLpAckd4hf06tbHebGvvzP8EPVwFKu20XLC3r1bBDTL+TANTLTy5A2ydkyC8u
5YUIn/E6uNOKPN72sc5DkOtPh8bGSyAJZz9PixJCR4p11jzp29/bsM7xhD+jHpk8
AgR21LTWWC+1U7q/+SXn28whDyuOrERMiWmuWSRkd/rqGCYSS57f6qeok5Lhh7K4
GHnDQfUfaN/QBhuQsz5JoquPEnWF6VwnvhLok03DDA895FBH7Kp+4d+3AdpPUftB
XH0UKEV+lWmjGN2upZWAGUXi+1X/OQr2JLDtGI7/2qWU4rSPYceUxNCPdmEq2OzZ
bi8Py4O1IoB2Lgbf3sae27bPRvzUAXJg/9126I1HoAORpq+ueY3YbwUvFknuc/WL
wbprwGMY0pWobTl939yOICB2QGhYtenhR24HeiKiPIV0D8T4wzP4c9rly8SmPlJM
1HjmAxiubb/omW8yfkXLhR7YMjfnHBuZubuM1lRvy61UuDbiMyAgIMMamsraM1ip
C/2H+qtmXi08pUkAsOgrp0q+J5Qk0cgsKvQ7+k82C2W/1SlBPqWv94S3v+ywVGV6
vc+04vD5URohrEcExDtmHOsPjJnvORiN2ci9skootbpRzAqm5dsK8/MdN0o+dom2
idV4c74yIimgo+RRTvWCYxymmrH/K6DXAduXbVQVrDGIoHE7fC5iMiwKlkf8fWp0
2VAg97dAmdpQhJ8+FBbV3twil6s0sHiVeb7Eh4JBEiVaZlWGF8EN5oWH2+FpmUJk
9mHT/YSlPO+QpbOn3eXh10sCRjnk4DVpSPD1CFUxQZEM5v+gQI2GjHZaJ4hWnpxX
fqOTInUjFBKjqpVTMqgnVo07HUU1N1AOxQ1w365NgcA5HJIk84VzK5W/PX69uTqq
66b7em/uP45wtXHucZqA/v51ejODbac4fHxxzSUvxe6lDb9rTm6yCvJTz2WM8Evt
zqrUwUo/KLkLn97YiqMUbqOAlVoQoWXknBHEYJNNN0chg8YUbXm3S07q9shEGbmU
uUiNqFP0FY9ckmVocOUZErvrVbBI3e3ie14y0Wr3KBvcXitmtYC1MBwMxqWL2cmv
/+OtMubYfaQ+0/FyX4X0Rcz72OzL53X/TM4/oG+rPPHHASatQuW1Omwj7A2RetRd
SKJ7mxeYd9DO8p+xnSvfQ7KyFix9l01iX9XIJSwvLjU+Romqh6G+JtsJtGQsXL5x
B8EEpiIDUl0JApTiJNkIMDCl/GH4oAZK/YybjEeSTmnTnMwxhy5EvASQBIYO6S9H
nghJxWLe7BFGIRsiD583pCdi1oPMGbeO3BomWPUAQz9vAzJTrJ9B6G9LwLmDTNBR
DZzgsBehjwt3wNCWyB1NNsNIJPDhUR/HXjdH4bFMCcolbv8jtsFG9zPX2YZdsgpa
lob3pW+GQrX8CS0lPKBDjMWDRDQdIh4LB8jsAqpe+ASuSpyKriiY7yb7JvqC+URd
Y4k7RYEJG76p/buvPS9ODTzfEkm9tXjJcA9m+E/6MzfWZ2KNJ60pXaa+DsEWyQm9
+Kapaf4/wsnW++2t/A7pX1SDxCcF1KuJP2j7t74r0qMa3TguVDJuwvXf6kVDKd62
o0ZOyDuHVpaWdCBLEuAfJKED0CF8h5JADGmZ+Ne5jVV0hmradv4winx1VxMVUeOU
g4CwUhfw0C50+Iy7HzriHZS/I8Nm2jaCjhOy2FI0Ugj450A+HB2m05u6xpf7DtDw
eAOE5NaMR6xRHc5QDkJSigO9l8qvhMK6l/54A0wLg1AfZmS98GUzXJ3vC5CKiX9q
9KzvgaTpFLjjgPNC4Q8LyVfV1dBT6zrK8MqNaXa94We8s3hxZOtU0qfwaYvmDiyc
DcHyX+uzKcwEUNWg2APlYQlJwGmqB/PoXmFFtuztrNOyB/iP7OaZN8ConNnw43HP
o9rrKJ4XTYRze49Ec0lrsDTT+NNseWVsWkDnHdwa8xKt32G32OCIfvCSq8KmV3Gj
Jys084hJA4zOvQclQcT+mZuCSa1EurQ/lExiaFkm4mouJMvrRkB6pHkCGng4ETNt
xcGgKFpg6KusQPrKOn4zj49Sny294MPqUWDfR9dq5fFVs8qypYq3vglmSSD1wLr3
p0hvixTxlXmnntwsxzYGzst6TcSvHUxR8mnwh+JTEu1p7kAj3N681BbKlVT+Byrx
99Ry4k5pWlTLN60ja1QzmG1Lfws6wZ4PjuULJVG7FzmodpARd8mCLPhlDJmke7Bo
Bt6tJc46vxXrCY3UzGq1FXmamz5h7/pW1Pf3zTSlTApbvFLdpckpTfs90ZCdRhQm
LPACT9qW7ihC5Re8fmHKPFXpYhZX+fh0ja7+aDvq8QQFQn6A47NmFz5cd0Vvs4pZ
e8fbIW8q79duYQzzAa7fTYOfS0LO0CTaB6MhFUIPocFDXg0E3zc9ecHVgbwrapvl
M3e9OU5tqZnPpWSb9w1j27n94AjW1fYBypehRTaSUTiOdeYtUB3yodLsbVTefeAO
CerXMvjP/3Man6K5KopTVY1fJUTlcOet5WqAsI/tq6f+gY+sE+SwhBc/Fnbo1Vve
PwHps1kh2y6vZpK2JENNGIybtBwaGOaE9Yl4FE3UyYt9btU/0GmRDiw1bXOQEwF0
cc1i+kCI3m2IffHsPOLi1lA07KrhDjKCVmixIwJ/nrfg8iOeKyHsfpCR80pf6rni
wbRsn4g7jcHPCVVRf8Gd19Qcvn2G/NKrBFxce98ReIS6AHzNPwguf47BE0mybYfW
aCGWe4aBNoMtm8CVziUDgke/6zeN6wce1huyyaQMbVl2tP6eAOO2Up6dpbDM45Qr
B3+mRskvqVjdk+JQjr8STNXT12X3ItlXcAv9pAgaRHTRwwX/vIpE725VDd+ArSBx
GO41HgaGfv72xU6tCSyqisjnUTXE8n680R/zCAzlNETjNmUtoLtLrsVmZDSrsVTp
QBhsNdS+XnJO0/+121B+zuFmE714i0FKMtl7HEBBgNHaCb6SBUba/UX4RsB4wJSz
LyHWnWaOOXuSP1/TUEBZTfH4ZB7KmwnndBnvQI0/8mVOgQ8U0f/prd3v2mm+XD6S
4yTu70jbXyuz5aWitvQJMTpTjxDsq7j6jswrZGjWfyYTQd/7cwtxKLQ6iz1iG0WB
PtO6lH+1J/PX6pRuSoHf0AiuIlZc4CJSIFC8C93umRC/OF4rud2erETBjji3mqRC
4zbliBoCcqbND2qovRDSygOUdir0lMiHvDzvqR0o8D/CVylmyJirqCQR7eh2Deio
Co01w7oMlseJpWiFvaE/o/LOjXdzKaFaGkXGfyHa6/cEJ1LS5Lhq58WKb429dSQf
4DhnBqOhkF7VCHwxZUhcB9V7WDIaYl/oVWLLJbjogny63YMcsVOG7/9Qcd768Tzv
DhlZmo5YJqSDfyLahNU+ZlG4SI00NfJUfuk7m6U/gqTjO2GS9ntPmTb/429qAEMH
rEWi6kiSYhmUs4QAK1nwX9MgAx+/JG+LXY/GHP2dLp2M5GY+TJPIPW/I2C5gFpJN
pxIsxdJ6xpqVvHSrTCm0fYv5sV6f/ODlfeSumxPpxHpy1TzuCbEvzUj4OLiv/nBj
NEIVGY3DBj9ij829xfeBLiN1t/A39eBjWvSrq8Q3FmHVrIrLDaKAnz6JchDJqLte
DJzPrev/iyav7YbRRAlZZh0Qoojsn6sMl16giFvo1sAS8rQeF4h97rT9T5d2IZgG
JtgdVSMNYijd6Kj1V6Y/t0bXXUPs1aVfrqovdJ1jELFcjhSWZnwY9Ev5II7C6Yor
6cwOU/eY1Wc83sGyu7Lj8HcSi8+IlJQpVuo8n1kqwCIu1dzVNZxpCA/5CrR/LqBt
VgTaGzw2kV7GCc0pCm09LPYvBSX6b8itb2qOw804OE7By3lu8pY+VOVtuzL0WtOB
bW6w0Kv3BSL/QYcuuja4ko60E4CrPcsZbbVZRb99SVMQdAzzd/jdCA4u2nBbZDTz
wSiT7W4DisQSaMNgExk/uBZAyNo3rpCTj92Q0qZCls6PXgXe2rUD+ZvOZ6h0BOTL
2KepcDvtDNIC+Ay2JL+gXueStztiniOVcKAWxwgknA+he7DhJuI7DeJ1qs7VARaY
C8mrQ7sBwtfPcw6xTy8iHMAQYK3BiExnclJnU9KBSzADb4NjsfM8ek77RRyesuHT
+K1FqqfK9MLQqcWFqEYKDMujdAV1NEi8Xb9bw4r/rNysEoXR5iCVPRljT/6NQFmi
DwxgV0HN0Mi1DHJl/4Q3zObyFj/sJmqisUoN0dBMKVjNCC19J+KV6RBummlqvdTb
WH7vbR3pAhUXGc6iXfrXBAYA0lBq0/llY8IwQxy7WmHJ8oJO3h/QKh3Lf1EK4HKW
J6qIH2uv/2kg64lCH636DJL1P0cbdIt1p02hi3gt6nb14SoGSdjsStaXYh0FkgjA
AZjAp6j3FpONVacYLZu4oNW79lI0SvVF5DyAeadL7tItpqDIlYQsq7TXyLrjbyb0
HaS+DOpMGjZZwC7CWT49E/2iBcj7pDSb7C3TM136wYzS1LQ3jAUseUsjJKsTXb3O
GRwziNB4daW5XpJAX5EYDQPxuf6N27hWUBuhEQvJNEumgnr8WphYLpNduSFPHrnD
T+qf5O/lYe87CA35FAY4H36c16QEERUIpZ8m6ctvNQoMncCNFVXD8yOXckQD5mMR
Zz0qVQB4LXI92nWNlPP8RHgq2uUZLbTJ6IbbfcdwgzpJCpMr2u+vtL/WPGLoXtit
RfiYrVd9dxdMUytK/nFynjRPJhFxHKjuHwxZsLSPcOUbo0VQyPSPkrZA8NSkjskQ
hR1EiVIqvR1FJBIvuAO9fodwzAWP3XZWPWZNc2EKbQf2fKWLREegurMmOYv1oRvC
GGfs+7nryfg4Hxow3TSz4VWGkcTno3HPTJkUCq0+K7lZroNUhSdZOoqSynBQRcT7
7U1/08Gw/66MkQ/zMpb6lPUBYqIYa9LLszB8fQEVM+fosC85JIxWiPVptbv5i9V4
i9kqclUx2PXX8kKSNoA9NAvSVd9L7RsZQ8raadOCfnRCIVr3PF08emh2K9E9d9L+
fhDnfrWNBXowNQDdB4WzhaOp3nKN3MTK2O56tB3TtowPIoI7CybNRWtfSZEf83Km
L5VRObAR54lrSFr8zDyEX7l9ASsUTxZ7Ux+4YJqeTREJ0H6MJxmlZ/7AqS4g0HDe
fs6ORQarXsB5dUek9IVoj4lyxTENx10Of7ePo3A+fTT1Qd7OUyaKWrvAhmYPgDli
O+U2KH8ml7jg13Yz2wvD7WJBb4D75r8xP2G3dtUbrZ4ipodl3pUfv1G+J+CWRXtG
PTWr97iwBc8oTD7yduVthnpcgmLQbqAIKeKkhcxbjJ2Qfz8guPEydVWKhe7L8SGO
UIgVdfiiHE/+Sb/t3Z2DYBH7FFwF0IYt0yf5dXqtWVr9/rbUICTtgAmYKAKGB7OK
utU274XcTluRXYvw1i6GJChl6ckbw7VXOfkKgj8O0rAwqac5JdOLiPcFPa1mjdhW
apLC2w2DVOnsLI3LAR0OYaPKqh56XElRmWESX8k5v6iSKTzFkS5HICqzvTJ8hWBh
hwNV2bQAG3mpgbuYvDoGBcMA8EgUOidSLJo7/Zv4enig5F+B2N3/3VzB5D7QBD49
Jr3wKzJzTbq5R5Z1k4yLNUYc4CxmAFIVumkKMEGofLO4lpSoEPctUksDoTPDJ2eo
ghqoUr9i2pAkguVAlCADOBtOWwVJauwYM2odcVrTMXofM2ScF9l7bFX08r2iroBy
2vxVi05s4mdgLyOq7k/tlB4LZvIu1/bL9V+vNrVeKdgDS1oJpQz9dEZaeGJlS+xt
HmklGsURDHBg+W8FUJS6Q+DPQ/DBOJZycX3vODK37kuSDSkTKb2PYQOsoaghnuAU
GPOSHpApGC+Wb+sCZSw8i6Bs2jMXHrs8YyP7gPLEHg9RfgcSLNmaOwyKrXwszqbF
KuRsewoZ9L+IY1F8QBpCtf4YiofqI2+2NuWS/tQtM5ud5jAeafA1YVzlL5NeVK9T
0/N2c4FW0f9MS3C/c5RqJTzF0HLZpOwGnK6lfcmw+nctnlZtu+GRp+eq/MmXRhuR
HjW4waR8mOwX17wnlIYgsJbg9YQfbJFejl1ivdoqpcRyYgFEK1Fe1Nbfs0gw7pXh
19ZOCcLWxf1OZ7uy7V1YGiCDhflr9n5NcbkjvHoZeFzG7cMVui/YIoqJKcvkiuP1
XfnBeXI/CSUqbGbuXYtwDyg0UmAI8OwWxjdFWD3KKjC5JkdEG40gq0x3qoY7hbMn
W2EzRe6udiORDYkumlgyqFyyI15utS06RhXmO/YZErwJ7dLA5hUA6qActLAItxen
zzORIPS/Pn+DvzMe1paQCn6jU7oZib0msmxTmG/A0rCvAPtH+DbO0snYg95+2SRE
4tMzyt81gCCRyHgmXmNQh7mzTaz+KBJ8EGsKahWijyOtcOWs9ZocdEy73PztwDLH
cL7rCGRarrgX+ro9OBWEiZMWDZ4L/RIehLIzM5Y3m0fv6uwEsl7L51W3cqkr5ySo
JyRMs8PBilH/QfrUI9Milor4v8qYZy7BCOa3P4GnBIaHXHee05c3xfiVekHfYQrK
XZxQ/pxuNZorByIJOqkSc3CwYDoE0eh/X5GoG1LzNgB/8IkJRUFTGhcUlGH9z7HO
j2M0X6X2LrYXkK+gbmqVYCElrRWCzdut2rVKhm7J74NBeOMNgbWirGO72vBqC+p9
Qh26AjVGmtNnmWtx8XLBjfUxITYoJWR4iZZtLmZ63hsSMyp9MSxeJNKWHPkpGMd0
+ZjE5tpMepxJtFu85GZNX15/BFvBmdS/kIhSPAI5wHI3qyb2OBWl1R7r2N+/h7F2
XAefZnwK3vTK0VAhVeiWZwinB5e7N2h9Mw1D4Q5QIy0h34E1bhjyB5pvnJvhi4sC
WTNDNG6XJo8JdhTb/sD23W0o+JQ9uL96/d096Oqo7rTok6wu9gNqmZ1ChTbx7+1A
3ckFySWC30sGPf9jXZwQ+UEXXjkC9Ee+VCYup2xaZf07e0WluFqk1/qkgHo9rXJ1
stAYtosJEZ/sWnlHCrjO57T5jCt9UTvVBPdykszagIEBc9rLslCokGVotN1YHv8M
+dOO2LLF51N3QmNM5wduYNmM2jJUcbJb4uObSZldEhGwTjQs8FeieK6oBboylUih
W/fcLLh5x4eEi4SsunK0Kg93gKQq6yyGbVsQJVEWVEFf2FbMSkbnTSAwnUkB1rVU
rEBNE4NnBNTIKrgWQCB3Z63UTaw6Q32OO7Nk7ZhzodE4ivcny4SZugxDmxlb7xRJ
p5dp4vEHGpPPBV2aSdMnKoQS8OKp0JNQJgM+8VmRhUKQbguk48UKqW1vtp2fXc/m
oW/yTywJ0IxoVE+PJcz9wxKSaykM6XmmmKPLdur2E+klhy/4SqJkGIVF3bdu/l8n
492+SR7JdgPaK8SqKCZmb5X9JglR4H34Q71q8YEbHE9pxkXCP/nUkUu+ZzMCjEb6
lxX1g68BbEQhs1o65ydvhBLLoXUT5sK92BIhmaE4wiN6GaS2VWOWavQI2jRcaF3j
paDB/UoydpWNvkP828/F52kiJoXh6qO4A7AiASbN4q3Jez3cjTQ4z1cWQkNrM4Oc
B0IZkc4ety1ER0ipoJA3zitlyw3EmsMI3hQRdSoNU/7PZh3rydOW52588BlyRktv
vWmwDcxqJQZKtkq2VCmvh6WUVODltz+upa2iJvBOuchsgT+znPusCUqFpqU4suqY
sA1eEMRbfaU9i+8fxnvmdt6rNSxHHqH3BXw1C5JkKn+Pq+p4TWBwc+xNspny/N2z
DZWtpNYVMkuYWi4OwklF+iTOttTdO5gILSC7TcaG9gwa8z5OgG1OySpWbUDUbJ/v
DJFBTin/EixgXxjeev/zcQGHjVx0C2ScDfK8YihDV37auLzEHMAOsEfAi6xyN+fL
qi2MxFLb3nIpESKNJ4CDcFMcp5dxiVolnTuw9wG5TCn2XLJDnQsKmzFlZz82Y/vs
e6gSJ1sINpLrnGcOlouJH1/8Fqpe8Rhmir/h+CX4Hv7r2ZI4ktpE2J4okLfc26wq
jYwq9z4xlRzNXVkGCtfs7bGWZfXTZTKmGFodftB6XFdkdJQW2cih4B/9gTnzIAFd
S4z5NFGMyTyAAUT3+7C9wUP1He1Y/R53V+hs9jJ7MKci2UIk9ua5XG0UTGfPNr1x
p7DABjMXzsrPsxt8My9UccJ/xXzAIjikmdVLEN6D2PuCdAufnpmeZ7oVNc8jQs66
kHNE51vDUzbox8Dll3MJnk0bal0bDOW2Zk3yWG8ttknB4aENgtr8BzUahaaBFcxh
fvydvkLGMwErYw8QqslZrOahXKUjQTgqoWwUtarHndJADaX90N8ReciMaO3znkK4
Gid+sxiGmWmILuzCLNDVHid5HmxcXuPnVIbOtRVGR54XCB07iax+8V2rQwAhxqjo
gn2yg830tbmu/suVLboKwTQvRCRHdG7YL0UnhuNNK5+KW/fZNcaxMZaROUPsWvLw
Xs0l2ouWbdaiuwUWtSlYU+zPCDOQoVQn3Dzx1VZRZWv+Jqi1e9QVT99umlfm57n/
dsPp4hGlGFgkdy7U/dKwgTyOaVl1+vljOLISJYvtkuTHzCqUR60M/A3TyQbfl06Z
VXkdv2LzLWo5vCtJPI6ASPk+98XeKijMcbUD2CnooU9gQNerRdyzpejiBoVzAZnl
l4JPeGmgAdDOYCd5Z+YjeUBHvovz30R6LgsEQv1PoDu9joa/0EC8ya+yunFyTsNb
XPQh/SoR1jrO1uvdIn05dgN8R4QOGpeXaLnePZUhPAPrJLGKQD8pnrNNudUWkHuA
p9aS4lnEOLLh0c4saK2EntPO4J5enjcnj9drkNlIHAiOPUQ1ktHTEEasVYlI4m/S
2F8Tz+ke8x3nHhKL0peEAvlQxVyGBCrTDyCoa8ZGxlFbAmFEPWMiaWKyBm3yGqOh
+/bE74RsXh8RNLXjlzQU+FQ+fxGGIF8t01m4jrjh74rO4pJ5HbzwIjk1KEjiLXAH
Vd/OwyEc5PlmVBPB1Cxnpkhl4nHKDCAyzHzg23A4Sq3KqLu1vORjcrc90r8zgXRi
xlPPoYEqzQ4nhCBNvbbNvO3aECKdyeOM97uBE6+4qzzrO79x/jdeMB/ollPQlvra
6fvFVg2wywnA2kfoqaREGokuk5N2WwPPYTwP0ngVXYuab/N4KjCjJNBZZK4zJnfD
OfN6BC3rBYv+AWz5t80Xi263Mg9NkV8THBzyjOTLJh579QXD7H3OlEVIPH32MpeS
Uew/qKZrsCbtd11vvD7If0mLx0YJixFfoHgNi5xwet6zQS4FpOdKgB72BpsNF5/A
qiuiqkf4lB5VzfUYtzmgCG9LRgkq7vruuhYEh5IRrq0j73cGaOOVdk6Ba1FRZQyv
UFMZLvglTZfWFzy4i9sA5Ic59sMmLtUbOGMp9LPFn42zYo79sRnagK8dA4UtXYC3
uQsjj8dXWg5efSH/uv2BOB0turFp2J1i0XPNGxumb41uaKEjl2YYg87dfcYvDLbo
BfmsNBqvgxUUNoUubCZ15z/LCtfp9XDo+Sr8cr5VTcV2dEjGXT3M6pCFZLVS2n9r
qVHO8NTN1t+3K88VvcNt+rNDK/cjQKiWB7SvJHygZd0LVwxgQ9qvALJ5PNcRPc89
IdWN40+FH0H5wuJBHIegNqWnuMnFg8ouJIbl3OJyhA3akSNwn6MtRdShlRVrXwVJ
A//x+v+zBqEKWKm+uY35YgCbEHOKS/0wsxy5X/SV89+lGxF/bgOiCa9aTuUJh+Pj
AtLWEmrxDPkN/EpqtLHKCwT9PwbjAqsiMJbfY5IJUrAuhdqhliqbiSpNoSH6L19q
BkbuNY8cc3KUyjUASQBFugBV9Oo3+ISUEDlMLLPzdCVruz/bzKJuktwbJczCXJi/
s8sxwBKRauYu/9WemPh05Ft8971My/FbiymzR4PIPE90F0xNSMfXerf5vv2xBh+M
siWxOFApjrYjou8tVLPVl814PlNzvs7bZIwcYCY7NXG/K7UOKI8klHs83DuvGJCz
l+J/QOt8a4pZ//JI0oC/MC/LSsUtSWZHmV04PDxnD1GSNlhC3Mqke+pOvT919pwJ
mDksL6Pen9pGUOB9QCcnjd8MuJuJoN1IPrv+ks79ou2xqK3x2idpHrOpEdI6N9M0
Sa2U3zKBUcNkYz+L70eL8DXIpi5EwWTZG753GxL9HxZ6pdmyB/NuZVpUlZK1o+wl
CkchM4DIsS2GI99MwdfXCDwb3Y2FiNaQutpdJSao1XfFaD0fuYmVztg/AUjgo0B2
BVQzCD3uGVf0GrDzfAGCA5sq9GRymsQ9cJqzJwXPEACXVyK38LNwOZyUTdZyAkTM
WOxdEPp8waw/Y69yHR8tp/SUeRTj7KHYCi5B/RVIYLS1ummhSPPMYPUAw4Hvhz3h
dHTScklCAEYiJf5eBYN823Q6qFcfHCEuqCWr0KOdnt4x5kLVgxcjVlS9ylEbDew6
+ecaGgLhSizHcbF+6seiN+3MZWTB4iTzWvAle1g0uJxU81SGVNEChpt0BF41BsjS
fzt0/oYcI4dsy3LmHTNsU/aGeT0svrzWNoO2cJ4YP1mHwDIcd9+KI3sLv0t2P5Xf
O/YdplFesOD+1gMUqPZqlJ3t9oB+bvzXoWF6uyf9RCEWQUBrSMqUujVI6S/WynqV
Xrdh5afiZDUTshAGd338otyoj/gAOX82xpnpjEcp/mxU2gaTbvIt4RmdEXQVS4o+
vB89SW+SkswRlLTj7nruIArMX2hoJ8yHeWDiQOM+47QtQbt5buMamjsHSpPhAc7P
xNVCJPVAIOlUrSgNOLKn5rttoAmWZUzgeNQxjy24oc4RZl1qg1XbpKw49LvRBkZp
sBKCkQc0dwOFn6sj09jyhHbwN89EWkkqaSqLjdkMdGLQJvsC1C/giF6EGKm7GgSE
nYiftvh2fUQYKdZtt37yfVdisqV2TMbu6YYH9vVMt9BUyl5IrhQOm2Q8H2dzM6YN
JR0nlClWKKoXNZ42e6kGgUOM/3Cy8xAvmYLyOzX2cl950kV393iftLOiFWDqWt1v
ho27UM2zo5GTuEPhofyqGnP7gYMSAZ7AGZMINZIphyidN3PtNE4PcW4tt/l+YA5J
hRitfJK4orvuXaS+Q3gf0Glgz3oWN7hZuw9gRElItIdxbzj1ekWwuT5RZshNEM+J
ZSZq5YQdb8E14lLWKIO6jfj8v2s2KyxoHYziWW6iwg7xawOoN6xCq2ASXdzTb3Qe
jqverVu4OAVd7Bk5GtDPWDue4Y68MYtHB9yR/VQPDBWRFLF6L7KlVP34mDSCQ3jv
1+/NCITsbIKEbpQJeqR/7YU8hlXXMrgshFiJy2dMtB7UfLtqlgSxtV/qcQYtVYGw
X4AFvlVOOelhdh2NceUcMFQFbrtE5mo/tUywLRFY/zKXABFr18tpcsRQ0epBOxg6
/wxO4bebuWpL7R66gHAfv1TeXVcTv+3omYx/9b0o2BmIJjp9dkIoR+y+HeClt/0t
NmEIB7v8PPY9kHMNbr5L5bnAHewvVcXQC+bhUDT8hLWbe/5256SvM8XgxtAYY1bL
2udtjlamEZnljDHx9bKoJtXeMMO1rznNL4n3z2ZKF1Dx65hsCPaFih8emKpEuCWa
R9049W2GiSxUjtlhKbfXddEU87W/dbw7yufsGXU4pv0Tmq1uTOGhTi60wKgQO9d5
N3e5G8nL7hBZEko7rHfcPxU6mDMdPWl59aocn+swPzk+JmRmnKTCo8X97CrAxF08
dMTMJEuRXigHOUPYOKGSX0z2KphTb3D3++eUNj7HDwa5DpWqEACJP9YQ/LLdraN3
tuNM1b0IXRJAT+5S7n2orWX2oKmU445lrLBXCm7VpV/Sv+F9og+Rp2r8fKpgxoyU
3ixo/715q9cC8EnpY2L430GW4NsFLjJOxyWXAUTUTw3yMOlPyGsCtbn6yg4T1hBa
qgOS9JLoEmZZWAuGWjyZtU4wart2sE3to2h8G6zQ7Vjy2waMCXznHcfLuKPxEJ8Y
b+wpBYEuOLX1t/IKYyFpVWzjI6tmlUgqOqdl3O93HJ8kmpaQH+4YgJ7TJ1b0L0LY
bZkONElm07ZGQTwMRFm7qIkPIjRHSThMV6yASOZt2NGORezbkthrzV8+v69GYSTJ
hI4H9zpgB4l4gpYfmvbTPPZD3clQ23oPXSz9YgKpweOGKttz/mti1P3Q/+fnavj7
/+oEniupiFFj2+Fh7WUDY/Q6woP9QPFH8GOvczLa+RRq6iFpd9ifOWSx9iblttDe
TFvW6mLQn5gLCPo9v5tmKW7CqNpLrsPnGeQWzVdFDFN9dF9eWJ25VgaP5jqWnWGq
2xsreJymPOw4RWLc3BFCAo9tflbnidz27uypekVo1VZzdr/nWni2R7MxROnFXgRu
qYk88Bhrm+1FDmN2CvoMu8xcLrhjyEoCKAm47PrfWBSaNvpIwfIyGt4yUMFsgYWM
P+8JGCI2xPYlRPgEPLb72f2vhKRn0I0FS5pvDGN/tSHzaAuUdoK3zieNZO2pcIwC
7hKaxxOmThwHmVUzlVliCJi8v4TWLCiU1reF1lYZu5gwg/jpxRLh74gKLqlViU6A
RQIu4dcQtsn7AFBt6XzptYWsVTnZ6PxY7zkpjgLRKM+ILfHs11iLLncfO+mbfjcT
HVzj8VYCMxw5buPkBNDmzOH3OoeS/v2xXcTiSb6Jmz8KvY4CyzMbBhsGNTs3ozgG
EiNxxN1B0BRY8YYcAIv33DZZH3Bm/e18LUxfG2KBsdHdJRfChhRGmQvAPOgtShS6
LTaCky8m2/QD2/e2rUwLLBRHxEFpQrLpN9en0vJaYrm5AlIu8IoKoqb4XPuGCcQt
32nJcPTyVrNXtvvgeCPz9SahvPBiCYsr7CfqKKh0sMw8P5xoLHA8ahHMj6bVCfgs
9fZpYvth415mO8mbDN6pQrrpsUq//nlf6mwNNHETuHWMcNRrvNXPCiGPasLZAhJv
LjxLcGwYsW5rT+NoUs1mV8HvXwL+13gkMZ0kMbxbDGwgMXPNzGtbDqrVuZEJp6Cu
3YeB+lro234+dPSWmTH4Ke+k5jMEqs4yI+8WilZh+NoaURL2b6rm9Siv/DWrYIv9
5tVjq0j5M2NIHMk1QK5VPe6psne8o3IihgM7tMSGFf/AXX1+/nK3XpyQVxe2guOH
/wwnEIKqVSINkVbiCU8ijthZr7s2Ktn91BYxP/kOFzSURDTlUULBgB7HEFbHPWeZ
FxazuXRFEqd1nnVpBKEBEnw7Gnb/4dX1674enS4m7QPX8dhvm4W7ab7+8lNsO4+G
5PmkV6QjM7lW/ZDqFPO+jy3RI2oIuh0R7N/Pwto+mhmYVvw4nkPLkHfKb851Fm9+
9izw1hfP4NaYkUbaF6its6nVAVpGLUSqHQgBh/rEbR5g/phh77nIDVTwNhHDvNBo
u06/ppTS6ZKctr4XnNoXsIeytaITsTYORy/jLA53Kf5Dy0tJF34dD4aRkBDdMfL4
gEgPxXoyoISh9bsFdRTsJn06PnPuEyk17MWLZQsk+RwhROySvS94Uqu4wdo0Mlne
SN/eMAE+lIZcGE0blfqG8ir1P40iTXKQU5PvKC5T7TtHyLPtbUmIY1FaINLr5TQa
9q6vwmgfLAq3CsB/pikxlK+PMSlkaRKdcDoFFRKIhQ6s9Yz3iklf4dNzZ9GVUPk3
mOyXO8epSd/57I5n24a98SuJDSCPEPGscNJG8lDUZax4Pnh19vTAx4GtBcsDDsnS
Rbr9zw7nH80iiR1nRTx/Jtg3/l+vgsItkav6Id93TfF+tVnAhQ7AxT8S+OQD0qgV
VTxobdy1jAOCxxpKiK0VUgSyTLeX1PEudV4B7mGxaDvBi7rAs4m8G/8Y86IkLUeS
Q3x3W7go8HlAMlYZE+8anwACwfD4ALe29lETD7FkaPBmnVpvP3WY4mE/ffPEwhi6
5781e3ODDQ/CRkXlW8JDAPLfvbRLGLAnVEIOMHnd42j/oW4YjGV+K84uTL+oGWLM
s6u8aQgepOq/gkLKempXpDN/ciUkZ9RZjdAGFOL6xMkXMHk0ZQh9DWPuY6uh1AHj
z//aFKiGj2ssAME4dAv6YE7hcqdYZXYgUykD8iXWTJOiWWcA/Ab+lrmEO2zlewyA
EblIUHOc9lS6UERr+00s4UF3cv8TquzpSzMxr8+xAagberWRPYIJoKFLLSR/1Q0A
38YYS2Or25KgkJyfsioa6xy4PH9koSTaaWuPF87pRGeHR/Jz5johCMavmFlM6wxF
25Mqkw8t2oLjl2DK4FMP6zUTdg66OgLx/rgwHjB/Mxnru4N9u4TJOlmRLwJF+8mE
ypgzLgu5MJVT+azcWdi8tK6MCLj6mAbwMo63HHBodCbUDVYioRRwOhMLp6OnzC/M
cJPd7kYXMZ39AEMqHg24N7EWLiPjyr7YD+TAsZmMGJRIAQ3gfs+7Q6vSrkG4JKvj
AbOC3+cyN0+rxV2bNv7exHVs90DEYcThXNYV9EpnnMZ8fST9Aplo4DIGb3nd8cYe
5/A3fSpDf+j+SHBBlCD9CkTFRDhDmjAVsj9XsXel8pQjxSz0JZjs8W2oP4wnRkgq
XMadhEa8T9gOYoLBj0y2DB1Nd/V79rjrbeF7JSSwyL3LLZSgIZMd0nInkL6Mt6I9
/jWf2TyLdrNHWa/8riS5xQYViTc98LCTXba9VT4TtLO78452JfIsBd/2FHrovqgj
MzcEPxztb4qJxH+EsB+SQeGQTMwo0JjLjmjvlKknNh76RQOUl8DJWso9XKEQhAm9
5de2/2DVkeSE0qmp7rxGHsV2guEDaImsXpPQXxyAbNVHjbu5eSPYTyDCEujSNMJ1
jMoHn4N7m14uBs0LeysZBNp0tnt5UUo3dcAnaNl9/DzMTCfsOVWi4uspg7MOHpJi
IkxMF0sWBdC0V4be0stvxE5ygUNvT0TIHR8iXBWAlsYIetLCyzH/pYI3nlfHyRS3
lpYRgKCbTWW5TskbEvnZz4IlPt5LaLHl8N4/g0j9rJJhek1YWOSqZQ+rlmr33FPc
FzKY6wpz7UYYQEmb8znHWxokUlGdLCLy2oYiXacP0SdVs1N2OQeTtljVlGgXZ21x
GxScqD0SpPzNivlrfcQ+uFLmPeJVn7418cRzBR/w33lEzgx4LV6mhhNo5EUw0dhH
4/nQEmY/u9etlDh0yHxEinnqVOSRybn2NuoME17IFbcCUMl3cJB6qchXtHIAuwui
A4DVKlL1lgGJt1FpJQDMAmfYYkPqVtDhExkT/kjXqSwfqQ14rbHvQ3VzSP9DFi9K
TvEEPSJDfqvU34QuUge8akFMbY4UmTt81Z3c0OR7TjSHyXmMm5tv/QHfoiXqvFvE
/De9j8cv6XiCz6qETc1jo0gOAKdpll4HI6AEZk8Y0RffzP+pFltJ0TTtu8PbOHCo
Nw21xjX4U0axE6lzDGfiJyobIx8SJSRb4fYffCVAi54ZfZc4lUqYdpM/aXgkqdTe
GJlf3OqcIhCqLI5PlyK978gKS1vd4HHWl22Gm72rU/s3Fq0EzRFkO81fmZ/GTwWq
4NJiS/hdMO00x2M8oNRsGSYdefmcDdVDvsiCH3S3xpkJkLF14EJy4YAIZXF9e+tX
xUQB5S8JacP1FJhObE3YY2xo6ZU55I2sFTV+fFSCLHYHuui3oVyzJtCmqoBQfCgq
r/GMlw9yakmF6ymfSulzOvHHMHAiwyefdGkcPHekeFxOdDPdmP44BKLpqNkL4+cY
rEwupTgNyTqKdER9/S2m8BV+eCqBOx7O7bf1Mb3EjDdoiVDJSET6qqFvu/k684+/
hpVpt1KdjNTLbjhWkuGxTZ7iv7a9YJz3/QBEDJORJOVHHICCxsPhd3JTj1+T9cM2
hUH1jNHEu1zB1bOIYWLB3nBHCViKhV2rLutVazxE1L0v33QWqldyyBg1K2OV2Wir
n7+GPBqozTqpBHBKeXzABGMIrcZtPvxnNqv8II7cOOpRrI+nFfDKnefATaVsx/RL
OtS8RYK/4Qg46X3P+ZuZebSN6oO9L9QvQEr54SFbtUbt7bS1Y29uCB7ZHv04cM5E
4FRXaG4P+7m3DAIjlc5WPg1DI0l1Lpur+zoGFSq0CNDcbzGjwxdxPeedhX7hJzug
jFHauzJX3QMNcN+kRODNv6duczzB5UJFkgDxhafofP71WyTFpeiLOcBi+p9VZVY9
UaQqrTUIwyUvu6HVt6TtucqnVGJCarjK/BNYmnN1qVmQNZaXPaebwcUTretal6eV
6c728uFaOQM3RWF08L+ggP2B3aztGBqlSrsF9/pSH873CMwcvO3C4USB0JQ+KCnF
4+CCJVaMQUEL+W49qLpojWVnKDGXiu/pTL/UzSprZj1JgTCrdDLRg3gGRoIQ9a2T
RzOLc4kjFrykpZRkIq5Qfwh2naFoJXeNUQNjG+e5jhKsMQLRbAeYHL+cANREVlGc
lT7JBu69w+pPf6o/SKmtpxDupQBrbfxS5TWbEcxtA6bHYFwQnBdBzEQi3flpOLsn
576PemvvhOxD7iAUC0leSiCuCLpy1kWfKg6qXdgp789xry0m02Z+9G3dQhnxn5BQ
NwuDrXnjvvXL7ir+V2ZT0XQeASl6LwIxOc0JN0S3NbqK2obErCgqT2tUX7+13t01
9/Vx2trc7+u1XRFmjElqQEFi4PpjdmUeoa8GmFQIg/dWtbsJQBpuzPPQMiqvv/FV
oqJbcQssxm676rs5CDv9DtOlO/U7i6yfsNkvLIUUxvNSAWmn+KO5WLE7Tpp21T3j
aFDjSt4x9nj8uBRGRlsajwdECUXgAMf6iR9ZF8VmgCCsgWtZaBQ92120J7GfkJpt
hmntQWI+9mpgP3QFdn/hN5qncN344fgduyIeKYNvxKtyVKsdaR8PCAZ0oFQypE74
BK0uQ/tkFeLrgdgAZvm3E/s0/HKWqSc5TA91KzFEWIdYmJRBTfMizl0Dk7Y27Rih
F/9sGo0cgE8/vdobXNWIqqUZPVbSj6GFnJW3eECxBC9MGu4LrPE1hZtVRPea59QG
TgIK3sOGu9zxVHZNqbtG9P4apT40IcDxt+P6FZtPois4CgSUv0R1ubjB/jUSmkfo
YjtRE4X4JTl9P6n7vBwCi+iZhSQav5O13uAf1MOIl0t4QzVVM/SN8eM38HIfePSm
VQGSNmBMv5klAdm/bMvBUEUMMcqDVDuAzSq3Ztkt9Gsapnmq56nzunoQJXAMnXNV
3AIwZl/KF/llgVs4dfs1RxdMj8quxE/yKl+D4udHsQ4dPROHJ8NWHPjho26Xlv2L
gVEnpCZPZJrQKr4H4ctNHqQBg6kCn5LfMJj+tGdzqp2bwTnwePz4wngcegWp8Nb0
JGvgrnHZX6tVkgkywHLYWbrDNV3cx0xb6/qdWYjCOKyd8q54RU1kInClHGVST96K
5Y8RxPwVcvbNY7CXuqNimM1OJ2Sk0YXHmJWPuVisQzfrd5TMCpI6FAT74mSsBFtR
p7gVIcyq31Nsabtd9xtGjAxsDgxhJxNCcR5CQ0ghOUNWwkR/2YqBljiyq32JDJyS
U+b0QZEzl8a0JaBKziAfoaUc5zs0jz+9oDUg+Gu0gWqr2+ubAK5FucrJU5nPU2OX
nVa1UngJw7/4pkfMggFk4IwtJu2+7R7AO1PiotTN0py/7i8oVM/TRx5r208OtqeS
H/B9OuukY4CRAKy241tIottiZD8c7he9gzRvTjbWRYG51phxh1WbMGbJfa/CKRoe
c/XJEVwcqAOwOIiYNhZk9PP3bzOkyqQGYK9YExClHYt7K9V5xpTqoGFAMYCue/kg
0ks3V9LpPRJ8h+0z3NAaUEvgsfy5ocS9jiyJEERK8PEQJMv3lSBuQI4JZ/2cUlEm
Koh9vBi75kbHRRNusA5FKaqeMb5plgGQlmBsE/da5I8M+ANhko23TdD+jlHD3TVL
JsYg/g8hd13vhyxDCGVBi60u7TIAI/uo0QzWNMfNlR6Lo3oS/poAdO2OAZw4k7kI
86r0tG8u91ua+zy8iehnj25yhJm5p039VsJDqv18IYZIrggTrNtY2bamjX0CNh24
iJajHkpmGUtd0rfeqgSMayNsMEw6EhX1yPDuchbV4OGbbxZQY+DG6WL/NhMHWYrw
1KXwHtCWqeo/cRRRx28WG1ogFn210+/paigj+6vM9TyLqNDHAm8TytBKgI/nWn8I
uLByZnJSsDWWDAHoiqkQtPnSG2EeLGYc8FkwOCv2gvCTE4OaREcUUAhc6nliSNgS
/ZEOgm9CaZ1S2cOvYql+JbaePmAWax/bvnKI6yddjSuweYutxddwWqQN8wHBr67M
sO8NbvR50u8LYEJWKvy6o3BtvpgcIVuZZorT9DONeh6QUJbMH458SVBtdURw7Rf6
Rx6A9RdQatUx2JN2dyAOAvR/HX79bx+3laksLC1pRrVqBiaVO/UurGYkpmfC0/5w
gaiRqzKQTWdBaCyYGH9V5y6pLEWUhL1sRYN1mWbZePC5YlbaD9o7nr7vQfkCZ/kX
A74wpHAtPDpbs5GASngcEZHBgSj4BNXtHf8rdhhC9fHych/0RBzqfF2GtZ/8Q8Hb
RG30rP4RBXOvUCysduDfdo2h7+uUXaQSnRhhmAFtJGNe1RP4B//NRbD08mb7q7Ey
RIsW5JojXFM8ngM8RlvMRQqyJix4xC3mKmz5RiCta+3KCZO38Yhs7NwiVwNG/L+P
pIsYTiGs2W9E85VPumCi7zBbF/33hSfbo1WEs6r2/IUlAiQ1akXC2wIKtMczcaVu
zGQz1+uqp0P96ul2PN+JgPM20v9rR1wrnrPenAZFgklbFb1mXKN57eovnI9DsV9t
CrDSPLNAgKhHR1BOFw+9xMLTLrnSOgZ+f2aghblF5JLAZ9rcTwPkYNTdDUoOPDj1
7DBwwKoKtIdA9Mood85o4CgoFUDTHK1w1TYkTAOruSoz8y/MdMdfCmOZCbiRjria
lT1sE/70lASupbmYzSIGPEk5kqk62osrUp/L7Ic6upX1H6nLMMnUCfmmL3MinYVQ
aiGAjMOtJK9Xr6hLN+J6RyqAOZFqjO6rA0rdOi6Eadf00dLoamTFTNgq5AnRUlVS
ypeCxhGXR6Dnyx26tkDUFz9O8PAYD6BLABL6JZQAhH4tLZ5BjYb6EvoeIwbOdICM
1X3bS9PvltdfGIslOXgMqaGkfJAE5X1/6er4r0Lg7+usApMM3G1cW2aevzZegTmY
KGwrOvGR9EM/y+yAME1AMFXja1gl4OplGd0vaUeCaPdljf1yKbJGK5RUAYWwirIS
64zjrFv5IXmV4yVTpvEavv2V5k2f1yC0qIEh1UDGe+zCXfkP4SWYbcZ62C5gAI9s
cNHxJ5pzR0yla4x2kwq/0Tpxn+Tt5SafgZ4mtvpx9+VdOuiC/tN1VWdMl3Hbc8fv
XXBPjpeGat/RPPdkkSYwbRdbvk0uorEul2vCsyu9l645HgoboGNRs9y4egXgQGuQ
wsqwvsOBCxMJa6MbR9L17zoqtGKQ1L/PpYLM5zVGmraqUhAefMyutJvEUvljEBgf
WYSQzAkU1kKvDdJtsA67EX8yxDDxBMBPpV3GZRaOqY4lOlQoXbotn7lvT/LJR/I1
chRLr6CVeZI2nrhenWkhbaV0aT6e88wkWF87/PuurN2d3ggJR4Xyqp5JMMhajLml
Mc9Ue6nGCl0bXMbx3V9AIITm54TXtboBgXM9T4lDsoyNjIq0MiHH2pVpfqDKsx3U
KJhgacDmmIvCQJwQyjEQevyBIOAmIBH7MiAPIz+IVaa+jFBYxVmmVdXErhhWUdaL
lzwpaIjXvggfyBTK7hJ4vKbRKZbPz8KriP/BHiKkAFKSvz1FeJrnXcr3+A4FDKJO
uS3YX8rHnevq7vvRIVrVW5VJ+VSm4GlHuIPAVq2+dsSw1NYwmcowff/gyKbUWu06
V+LDpIk5bEYBzeq0mtw3ehpEtaRXzEQJnVXsRQTr+uJshOFwE6Zo55p4JC7Wtigo
Bl5C17zHOA3BYHptNOuo7TBJZ+j5CquEHCrF7qKfdfk7Vu6kEsP/laKOfGgJ4hr8
sOlo7J3GPEewI9E/a0e0nGr3OUXEnAAq0yVA7Y6lHRUO/OOGnNiLpHE68t8cIkaT
e9Y96mw7nH1YN35KwB/Oi+Hc+3Rb82lyUNHeM+eGLxzZhryk223gvgORxwlOb9Hd
zpHB5Zg3ayJgTRLhlVDmGsH7ehr4l3hFCHUUxRMHlL18sdEqPftnbR6QZLoOT3mu
qkhFoRto0u8WsuxOuhM3PksPzXRGA/iSEWc1ucgRsF2aerHzC+QI0LSoh7QSnAwL
StDhad+KFfdU3xi/pIQI+4L+juuFlZsRFEWudXEsr2dmR/QnQ4+q/IW/wFjyiIUg
I5dNg0uen24Q4IeQV0heO9lke+vXOWsj8XutVNCuXQte8vJwja4xlazY7Yxl8M+f
xMiegQtlIs1f+w/93FZmRpFxJhggwQIfWcMWCsGvYtju3AEV3Y9X67TjgWTemOev
l9MR/s/WQDrAmXjUoEpIafSX0zWyPtVLXjGK5HJv34E7nh4ZajB42K5q/P4D/mCb
jqOsqrYN2J19o+7QcdrtjjzUhb9UJC7Ir89y07rd8ZuQUum8ItgbiDLoARI8xwEQ
RHLyREPK4nI6LGSgSvneJOxVxFY/OZBWqMqOIPzRnAGxrvILWHcASgzwwAVXBX2t
L2Vw1Y+QSlSp1iqVOjt3iL1x5nnbS476JYst2hccUOm4ziZEF0TaeI/Acy7fYc6H
c1OjePB4wXBq2KHwczKKJQUnqnLSv0dOj6fqS917kFHeQ1aX1ZSk5IHFu38gLgmu
7KkWP+5jNQCjsShPbpEVJN31IDqk23BV9QQ7/BVjtu55BNaMJmSBmTZ4sPubUBdo
AAQzR5xH7be46lfOPhDj6bEWgj6QoWv9BwMhtNqSPMTEfPOAtIO1oxh0Ukib7J/s
cAlGVgDQkaoDqyAwktS9a3lo+G9C5wm+jhWXlnnqbkKDWpF9y7rcH94fb9HrYZc4
MepVCfznM4opFLvflQfLfdxjFl0d0ZmYLfe6L70NsQi7r5x9/6kNgMUK9uHwGU9H
4l/eyo+kW5Z3djJsUDPToebtnCuavFttgPKu4FoxjJRsUKTkIco0e7pD6FYCV8ib
2Gz2r1ZsNjrZkbnxd5XQ91s9NCM3ppJxDr7gRwGSSzI+rYxnLt7X9ps6WQydGhtZ
5XmLTxzM6bPAoG3saH5TK/VMlYXbxuWKMioYPLthhGWAbHsRog1dWFkmZQ+OXNJF
6ozGoqIIdAH+UxUEchmc2JHRClLQhvEBw7nYDGzqNetRh8lpwOmcIqcJ5b00tHT7
oQ2Lw4SmrY/AFhfR+E8MPnxoWhTuh+v70DFy6LvWRTFYKt51D3EFgtyrv3qh0sCD
zcN1f/qTYwBeOaWg+2wCtDH/zupWvbuodBiMQ0BM79Xs02RzRBl7PU4nHsrsDe5a
XgII8YsTIkJ3dBC/jV7utO3GIV1gievru4nUtBWONnRtwjMOD/d8cj2oYOR4nGL7
yFmOCzsbYF4zUYw8CevDOwqSshfIu6YZgm6C00u5AjVpEA06JZJcLMemseVeXn4i
RYNb2LCNcEGmf170Yrwy2GNMV+SmR7fnJxJn5DPddSmj2a57qR+BMaBCSDWn7CKV
WKPImSE6y2EaIyoTjkiAQsgiIVVORTkIunt56gHsavrq5SWQcbr9tNxhNjhrIT2x
uWjS5BzNDZiw7QFCTMHqqxZXagI5Tc1hqXeI9qjxLxJleT68sL88ls0EPNUCf9ow
8ijCPZP2Ss9TUfy1QGqkZ2fln+YTYZ/tcWkt4g2fH4nudNzwxEuO+ypxbnMFg0Sg
RxKE/N2hXnzXG4GegjIvN+BlM+35PYlqdaJipLpTwV/EmLIc73kPUgD/bLlTBR+Y
ZAxdYBip3HLiMpoHtQvdNPxcaRRfyxsh6ZoOxLPLMxXrksboeGeRpT5X6hy4DetU
vsYEg00WU15pEIwsyg5/q+lRacNsSDB2B2rnY+T+JEVb+M0dDwgJhB3TzgUcuLt0
61YQxlAG/XrnlMjw7+Je3aSXFjG570E6Qym/mSSrvC/G+vy8JV7kNV0JLNUYKwKR
zj963aEd7kfUD6IVfJvPmgt5btgCUKa0NAMKE+0b6vPnx09oPgCF+AgE4yqNn1A6
PZ8J0a/B4F7CvkGZYKDUMcde8/GX32EAdD1oK7B+E9xDMS46JW9aOnhORKzJ0eqw
9z4M0NlqdoUHwet3IP1A0xeVoYThrNJJF7XKAFN6U1oAVEAqI/G1iFIafoY28A/E
WhcGY4BVoMKkIrsr3J7bbCCkG+DuLVUdy00pGaCELnHSStUWxLlTUoFyI/zye8Ii
0Wo/fOzkb+BkOeiDXHZWCLOhNB7FY5zWx6durXUSP1ju/XvP2PdzvRL8SRJ2t8KO
gScDaz8rIrKItxCZwXGYm8MUY6Q4EezIT6mbkRGxZkh0Us0wj8jxgntU38/XkmXT
uHD8uieYsbc8WZ/oxEzh6dK5jnLYrNdmy4BxsW9AhdQXWOUFr5FHyy6hIQYcPNA7
uyb5BZysWmeeObKFpU6iP+/wIeJuvhvOGFU1Tvj2HAhMLwB1JXAN4aUePwfSj54R
ZafePMqVC47ZnRCErplxCvPqOX0nn04dL8Gef2oOaWqwUQ0Se3SD2em9i+ZfY87G
dN7mGwGIKM9RPuB5V1XWFnT1F4gYCIQh5VW+2YFIq9klTiMNtl1qSk7FNNOJKt3P
2QBCmZ0ZH1VPx58yMK5UvKRDreaINld47xro9OMg4Ip4w+TkoHe/DPPK+kmcnWtt
qoGb9BeJnOMtzmU20Zrdw2ENLP1E6XcSzZnuGyZXVQbAZ3WTGRYzMTSgn5D1Giz+
JWwdEmuHGLEtvVBpcFy4EOD/E3fGXK1TMy+XQ+y+i3ZwxfXu7bcrWg187EnGcl4O
KUGCWXH6o4nwZkPCloqlmfBVqU/WL8HlXv8M/6rxpFn99G9zwNW2STOuWQa/q2Bt
lApgP498FvfqfS6UqtsqULEcImIlRWdhzFpli2a2qOEh0S+R0+xBSEyAwOxgi8L2
LFskOF7Zx7U+JZ5U5p53ETxXm8DYmTGAVqKbaDFd0NuMAPIpQN31150OLa62206O
iXwg1y1LgOQu8HjkSF+JSVl/4xJIGhTDIhZmWx6QhWDwslX93gtM7DiO/s4uuh1j
pVM8GpADHIDU9t/hnvhvzALmZ4IEzzQAZd5CmuLB0c0mJf3i1uyr1aAxVgV6DtCB
rj3MWLFxLGyXgeFrMFX4o44aL5ycTfLhNJq7GLZw5I6Up+OtL24EnEZrzMYok/8n
nAvObN4xYuGXIKGLxplgKIjFbNPgfGdagD3mu6jTh1utfDCR3GeMqBDoNUZGyBNT
5xZCi5R+xiCvZYtiNoS5gczqZul42yoPdIO+Sd2z0s79NiShJD6nkH561fhcVBM6
QxlEPuJ4wvp4henRsVW0SWJ6xwnSnjr7SlbHFqEx3B0cT94b4+aNdlgmw4041MyP
lCh18S8NUzdFSAFu9TZpUMggQMs6JpUK6nHoz3O4VOaN921RP8/6abMyVrumJpuU
xfo5xx4Jreuj8KPK8zwaJwHE9/WqvZFqDxDyR2gj1Rhn4Ik5CrTUa9GuZIVncbSH
fqg8I6CzBtopIp+XULmDD6+Xhfdm8sb79hu20w+i8D104YsPJQwNgk9pwBFeBNbg
x54ewL5Vxmu4iHZU+/a15Ox3ZFVds8JsPrRbL1GBhIFUSoTSJ5I22pwBDFriElVl
F/G8kO+9t781oh7QDRzguu33w0EcoZ3bSgrviih9fMKtnqra4lRhbkVFCvpgPpSH
yDX7U0hh3/OvGxHxdvZ4eejVWThDS8SBV50eJncoBidRUPKML50p2R5fB6mKMkU9
rg4EYz93wOlX9Zrh1yNrHhHDGaVlEgOYgsY54eV7wSYwgzH12tylVP2dAgk8aGg0
f4S9dBaICo/IfTrubRYymtz2HLxR6wO8vvCtJmqxMS/oN+0AIY4oFVvGpeJPsgk+
jEP6wF8pivrvaNfWFBt62zow3x983Q4jAFZs9So7G/wUl1uqRRu8jPjk12XKr5sm
bm1scOzKBQw+yE/mUL2SYel1Mqk4We72SNNGqyCAu94ol+eTu9nyuY3Aw04s1pY1
m5YmwDLVCaUM+Z6+6G2q9MYm54foNbxXtoZp9rLTkoRGFnXBY3IFTjy2Q2S+aPqf
wkyTZyXxoJwz1DvCPKCONthEmyuKwLj2K5Dc+B+u2gCSFJXn4Uoul0c7j7qZyP7T
DnFGtmId97T0fv8ED4G2V0X1M3NCxoWTfrrgsdM0SM0+SGwgEHL/t2uCoH1lNoQG
r93etpMjcaY+tbLbOqX6iyfYoGe+Hbsbth4/jZv6S4KHQcbX9s6vQdTXpkPpFBdQ
6gTkieIGXd6dSvxd8YgDsnmFegd7oOljyTrSuzOBSZyRPcWf+Af49cYhg7AgfQGb
0YL2C/UZPj7qR7kRbZ2Oyp4FFYZmRnPw8MWZ9cE/Nln0H0HNjPzC/OnNgNVqryDH
XKR6nu8L/wsrFoHeLBuNbbRoICHG2tnfaFqiWhu66IZHpagnkvsN4ZddEclLkyW2
c+dAYuqZcYY11gbT23y0QVpU0ICXlqxUfvMHlAQETGe9WLZ+WyWKT4cq13foBLOA
9/3btbS0tIYQHACPV8r5lNvygN7+0GncVQ2tOFQX0uE75bXfKA916sOBJsqTwqXB
2hCRbjRBe7L2MnJzfAOg+QOBrr49E3LlrwvEzw94XZcJDM0U7QicS27N7p/M75TZ
ZYmDYdx8kWRUVHKkgPJEQQcEYuRLrxJVHpn1CoVIfSWr8D+9yqBC7rdAB7HSEkkM
18Fu/dG/1olsX2RdYtRy4OnEuD+lROXZqwsxotcJfnTmKTBl724PJAsY6B5EHRmT
BOfq//npm9nFnem5N+JLnekgkgma9Ug+fsv7PrbZSCUUMQDNhxI20Lm8eLSkaTSp
K0ZeSOSRzGtQ+9/eNggkQNftHHVrr5h/dy5meylTIHaLhP6lqP9oBR10KnpSRKWT
iaX5BOsSBfcgqjM+wMzyFM+bkOC9JrhKO0JpDhnG48ZBqBU26tGg6+k/9Wwok2yx
LmW68COp+315fUs/xufstt/oYrHcuNCl4qOfe3nnNC8kdiZkwWLEkZPV7hFx0Tyz
q3EkB48hMBiNIu2jkxE9JgE2H64/zCRKQ7kdY4iVaKS2yo5j+Yr5yS0swwQ61OaU
cuxWw0p8GfKQ/cPJBTvVnVviG/fOVGNS7A66E0AdxxBP6OK3ihDJby8d3BEgFbxS
6j80Fh+BgCWtmhdlxgPndeWLBiEBxZapganoozvtitYbP7KBqg2GN2y0hIbeYtL8
g4ZVwH29tdki6YaZho6Y8XTn/+o7uERxAsKQafegU1ouGSn7P6Pu/9ansoNRUqa9
92WNWX0WXScINqbBeEh/9Fs7+iEWhEx1PUa9Lcw0Wew/P1nfbV4Om2tin6ljCo2e
aRdO2nVfDooJLPSV/OqTug6baMNa5Sle5uHBVcOFbqxYjCQtmVQ1OOhjCvGtRds9
qYKbCkAclVMT+lrCc400LSyzWX/Z0gwW8STgINN++16P7VreZJUJdFZ+mgw5RC3O
mF24TEh9r+sEgrtQGTc6a+51tYNk8FRZ8OxBdG8LVYa6DDU5+EvRVcd/IxvQ2fEJ
dhKVU8yMrC8qnQIDt+FVlcXMC8NMn6PpzLS6AbaGifNSkzyL31Dkza3et03SULaa
iuln02Uhm/zGKyvsueKhxdlIdgy6cnNF9PapPhceH7io4FgcOHQj3BRmUHpBZLjU
JOc+P4kVzxuepZxCPOrdJS1VoM2TobiEHTkx7zjxbBUZT/eljD06gBjCtMKePOA2
ZhI+ou1O4xgbtRdgkZridx/Pd5c4b1RIiL/IzGpoNokgL0xRqBmh5uRjt6JfLOO2
WK8fo+gzbiXRZ1xMrm2r5q3MZgt2f4+r0EdO9vfeNa1qtJpil5qrBLirU1Dd6NZQ
+Cep1NUinMeJ/ijkLSm71+84SBsetkGzDwRecsGuV8dLc9LgDkNUDb3it9OBB8QW
kd/j5zOdx9UePlmTHbHWyGw3Gwf4mrmKwx95KwQEzPwynt4xBFpi0ksOu97nUCXL
Cs9B6mqw5084/gTgN3U65dj3B9Z0vVmI8wEazeL+TMA6aZxCCMvWfqq9nWTSGFnj
8lO44bdU+Y6plnkF3HPfos8KfYQUzz/o88HJNUIfHK/p9eOg19AcXtKY+Zqmv0uW
7bDFQtL3qTsV0gC7VBXqJjolP6iPAGK47zKlcj+OA7RW+IumDvt0/Gavs3JZV74v
tASPKYjyUN63nzCJ+Xviyn4GLgZ1rMuVLintZGjZCLEn2iIT8zNK74+Ld8yQxJZ4
T75Bs/wHqZut80e7xenbmyaPvVbR1zHDB8uZz3pJbzKy8l88urY1I4tmBO1/NtuO
4anBJP/d8ODuvse+NIBLJ0cHP0s3J+V9/MqBJ2B/Y274If4OGxEWwTxjBdSGgEdY
xh0IUTCUfCBCvRCyvbWl9gfpFBR05D0IBft8ZAsWH082ulXlkIkdJMVO6OVmJDVK
6xjbqWAnnh2e/MI0eCowjPZnYb0WD8aQ16Fq7BnKKAcAxwUn8WwHQFpFXyIwEIga
YKmDNDa8XIwXeiJ6UWNsfQbPcc2/hzvlmQ/UPYEqb6GQhBPv8mu9aXgPw/uQPEwL
yRobn4kmve7IgEmFTl15X4ranB2KBN2ELCOTZCikTAoR/SDRlnwj/dTRSMO4q6JB
mQXkATKhEpohFAaQtAWYBDW+VmvvjOIycuPY+pCKu0MTdktwTTQNoS+u+ntiOGPB
XAfNi4DzbvlGkKhfukLPDNZnROtt/EsB7X0PUe8oYUcTEyCQmnVb9Ep/+1xpokl7
5Et5VHDKFcv54MmOCVi6zD2QCGPyFSVjq3u8AMZVXTrMTow7rWjpJVsU+2CKOLpx
ZjazHmDQmlHW4ynM/razUyNLeo37fX9jLlWuEHkRZnE0rDpiEVDQ/5U/3oo0CkoB
xz1DRjOewyjvmqkFFaTcvl63pluIMAXjUN2u3rb7tPOKqyO5s1tTXfX3tEmITLbX
0djoACVZUZCHCUDkX6qIJrBcOm20+OWwo6mmlGli9LJ37o2zmDp84amOV/Hp79fO
D0J4jThbr9t3kVnjjDs45YoKVEswgHNJIZwwtTMRqg+o0dJQnHtOxHAPZO8ljGDr
CKeo3DwmHT9cbNFsVqZCxIa0YULIwxhc76oUAmm2IJ/0nrilw1Xc6jH4nEVdbwWY
6RdMY+L1mYYLamsrAZr9CoKj7K017vaPuUHL6sFzZ2Nc71/wNnTPFEs1xKg0x6Oe
Hh52I1c0BNd9MPrzuQ+qO93nsDViMprGay2yicxi0OXd6QRfL+skFKjVhx5qB+uX
Xk1IM88Nw0aT48gjFkEatUM5GP5B/d6Nqzju9682ALARW1T1CZMbm3hTpRt1cZMz
suYqZVfFFWfVzHgOIdhQpK9W1Tro4Id3gYfodyFWhL6iRC8Ja0wCfs+i1LNwi/IR
nLQcr7vJf8JcEgHe3UqLQacHLnJ+1ERwq3hr0+MxQ6n8to6f/SzIMKRjXbdQUG76
0IhC8jud4WQuAUucJBX0IHMwDm2rTkDXIW1kpA9W1oE9Rq9wabNN3QbyyDUCuQD1
ELXOpL4jUjVg+mOpPAR0Frj5ichri+rWUW5z/UMR/UtREIUqQRKH3zaqrQMNwjVJ
j6ByzpWVlbl6o7Bk+1UIGCYjhpqD9EhKzGJCoQmlMA+YVaFXgZDJfiCOzjPO1Haq
gy2OyJmnT9ha3kUuwPF2brAB83MJkc1G4potyUaIlcVB6tbugfO2CGFE6PMfxNNL
jYtF6oZnzwPF0P2hpYToHmOQ5bCgwwZoG/uz3WWRfKIKngyAr32tQ6TVzG9hzxMU
/RUlG1aNouO7QaXuP57xOlbP1rwQ7lY63T4lDW1FDsbfA4aY5p+1wYKG1O+t1Ve8
JjO9s9b+drOqjg0qIsmclb7sXkZozkqAH0IoytiUjq8hIQMyKgVKssipk2RNXEth
pOZ5BdgYdOBvpUb4RV1JCLWNrgx8tKYzkBq1qGxSF2FTJ1RTW9eBHkiNTLz6klrU
TrxQ0nBC5wwqWseuW+FaIrVXfno7eOanOneA5fIoGPxkjkitN/BXsnzcAylcvTbT
/GYlxJ8fHr2ZLtRA3CFHn+Yd1kS7F2ppnFuZv+BNWPrnMYjbQEk2wtWJISUF41lF
cBe9A5vywzAMmD7FcHw/xWcbuIF578FmpEFoJ65nQIzfY0owq/f3AmCCphn73sQB
Z37Xdnt+0cy+PCogXD6qBd8+NjbeoBRQl5x6ZkeTT7t5F9Udt/UJ9ivXY8whgDbr
rUyg/8WE75tlWmcEi2TMV5PI9HKsjYKGIqvi/bosvHd24IWxHeCSFenKXl4Tpdvg
inpBti+tyuSAuRCjznSut6bziDqjGJ8A0WZmUwHM99zcTH7BGTXSAet5Zd7se8kj
8AMGeOzJLaGKrtBTu4ZS8SDgbXB6A9hERP5+i7emw47OY+lHFfpABs+emDOOTkoE
Qk48pXZYIbMVXqIenrCGl14T17NIbWyV8hq0ItwIjK5y9YokX5f36B601zVXA92D
yEzkYIYPkwpSikKGKGOFDmkIkae4CXPBAg+Fdj33Wfu9g7IOjv5j6On6xGLXWCba
YL5mbxmlX3Pka5nLWsrSVqix3DARqGoIJbeWnvsqKRqJwBDHzdbZ2kravy0AbIpq
HJRIm812P6hIUUeTGiG3vzAgGP+GqTZOiE/YGljqLWJoUxPin4koQ7lFat2R74q7
ur42iM9yN7ehoIv+P8nk07N5HlLQEd6wmUDPiGRsv40n0i+npKjrv3mw1uQO8t/A
mD26KRL3g7+93+MXEiCGuaRj8WqHlqabHcAw2vtX6/TuEEOcMbhFzuC0uxEL9Du8
HX/Va9YYhnWDXaEdpBNr80iZwJwH+/Zi7lyNldY9LQBEtQm4iU28Z1/bFOrh84DF
huIBI16Ty74lTtLAgdkzeWpNMaCAu0v6rKlLWoT9eMVmut+ZCAlJ3c29FpLj0NNw
tfrHX9Ta0FBU8/8vOjLrvKDOmjfN0tTYE54cK0JjK0G4GbUTno82hIvupCA67V6S
rGGtL29LHmp/OXkWnQpIw/bzrkEs3SE9JyqdhQN9ybQ2jEG4OQS0u4FS1dtSX0q+
fIS28jLY+UCTmlnU5MzVbXXZRjEWKJp/CeUF40CmLiJ8mCAWMW/FZvf0MKMeEZH+
v0rqFPrCl626kkfvICWdOFjWfA9gH914QstTDBIthciaj7wP7/ZxW29C2kVXbS6V
oAhuBmnufu045wWLU923vR3eyMOtV4wMQBjlEJBslFeluQK3/0cqgIidb9kdQUAk
qBNLDl2G2gk0AQvsZiTjQIIOf7nE5HfLlM+6Q1LxRbXjAD3mZiaeKwsZxymtFCGU
KC+UkqqtKuYtRIms2Y+j4vvgIpCjTm5Lk3dgu9/Xeok7zmRpzHsOU6yaeii8yaaD
LM1/nrp1FtQ4aZB9BGG6bJ6pMFcxh3N9SdTXssnXRAVdhPNJT3240wE7vz7V+goV
aU77lCw7owaGVnbcIX+d6qxIh00vXGsrmvxaEiaVH0kS8wAhGgEv2gq0RYqOw9Qf
Yg5e/fEA8UyU1g8UHi83E+iKo40SS0Op/CpkUKbUlfnvbGsX71o6vGF2c/Ki3XmU
VULI2Wn1TVwFcLAWic0Z9Xr7XPN8YVakLPM+eGADurqgB3Ov1qD1C5eGGrTHcCC1
z18VMZYCZGrn5cXtmD6eIf+H4RZIj8alG+GoLsTmIoWZgMrO5CHmYXY/cUU8Odlr
xlFLjNiCFJMBqDUhUpZhpf0I3GyAaC8ji6ntm67htBLD+ubW4PO83UFmY51KcL2d
BlAdjbq29tzTpBEwW5/0FWL7FVb7bS5xmgsnEvKt5JdzpG9eUfULwcbu8o/7in1w
q/lHkAYt+SKLKLeMji5CJ4mz1JCZcn+oXVmCrKvf7w3MHRuciIzmrHxlvvsIVfcJ
qGdU6RKQ4jp4oEm9uCR93dPa6BfSs0HvkzqBA02gqeICaytR7pH9sxZimlra0lZX
IECzD/bQOTh6+fV1hrTBVpVSw1YiGhADRlYTZnjQxg7d1B0V5fa1iZ79mTHTBntE
biERuB/OYk/JuqpqzDj1X57iCgidzyWA7D7X/2q/lS4UD1DYrSNmd0UUtcHCWq7e
roCuxHxuAnaodbAC+hzL8BEQqSq8f77rLSE3yId5DoypCzZqgR77iR478rgqHIYh
x2t89qyCf9wgxNnmxNSV6GV9y2VC/2fDuYab6dYX3TlQ1ZJaiaFklEmBjBc4Twif
1+D3NEm0WyQjLs+S7kjwCdBrqQLi340aw9YMxQ7JXgd+e6XAzicR4GdSvFag9nTK
9QGDlh5VLZEP7trpOAwNmoW7dAPEPYBx1baE3Lt+ctHrV1Te6yW+iVYdAtpMCzY5
TJT/NnQXQ89SvcVLsjwOHOGCzQiS2VSBQP5mPQ7jZM6OQjCtcJU35Ja3CU3FibCO
QyUso7dC1ujnzv7pcM8VXYPJOeh+jgkYrj49e25/mlrQrJOCDySbkqbi+0Z4Cb/M
tg03zHnlro4suvGFz4wE4e+aJFn1Qb68+HA3IYY0cCH82UMTfU60sbOI1Q46xhGC
4XSu2C+ZQ+7dMm/DoMiO6+ER/LeBvMKzGqVfo3W8fJx8EvnGkqIOTH2M9DnzWo8I
EVScARa2+1bQFH9w04CS1uhguYoyvv0g6hananeIdXD1BDqR+KD767dpmUUPNchJ
8shODhDknW8k9vG662DHhOyeLTbffjaX57Rhfzky9LdW6wpxS06ssT2fYAmjkH/B
6QqogrD5qHoNcOTdqJcLLo7YDODnqcXnEnS5HLqaxf6SkH064D98b0Ldzip+dJwx
kyPnuKofObgVt3MlZQ9vMIwbj/YbNiqhaIABGJONBKxKCNPhmePYaPntoawn50SP
waKylJLEub/xOyoHix8KyS4eAlqyUETiclR9haFUc/ml6tGscdcJ8pwoIdkl63eT
6KBAQSdeHjqF2DF0E9YRybiqrp9go+ngYHnQezhLnHIH8ASAknTbsW9nIoInMFLF
lVltE2EvwNhgP+ImusFkJf5I2vl5X4j/jvYOa9rTXZjJgdHhCd32B7Yim3TfGWDL
2F2dlVdog2wzTJwCdnvKz7EBjLxoMbUpq4jBcQojDfUBlmTTy1sY2ym7X/ZRbSSO
cl5BxJZURGlhO0W/K7ZmVVRCmTArpma9IgzeyspoPsynKFImW+xKmxCEUrEoLbM/
2JTY0817bt7o2VwwL0TVFqm4gKm3Jh2WbYowlV5WLz+btZCnDMBZIOPaUvjnQQbx
WA/uzJksSv32Ryx7pPae6h0D6/IL/1W5WuQKcFiICRRficoku4zTnMiCHXaaaVPP
T0+4d2A16w6ckG9Kv40pqeib2vWXx/VlvQy7ihmHjgQu589WX2vIi+cRF2etttma
jXxymCF+0se7I0LgWLnQLNEek0VJTTahyEyGvQuAem2UsLbMQhft91WcD6Jc4/V7
AA9AjYif3kc5OATVx33mGtoim2VAVMkpvJwyrAY7ArLzsrH3fV7RyJh+hPEFGkg1
SBWDgzlt3xyB1+DyZDAMKQuzdEc66MxcixLftpo7ZYdQNdKQD1RFE1poZDzbltpd
A2vHFoqtCGvAju5fDolJLlqxBAC6zZ9qn4KPWNr3U5f/wKqiYfTleE3rf1C3MEu+
pE4LRb0XBZZvbt9wSwHBZXTRl8/WDVH3PUiibcHPWjazBbVHkrmLkvdqHgclyIoD
4hiC5ve2DStqnBMd+Oni9NolLEWkikbciQ2wVTfeDKPTjgkdoMhVC207erXya0Gp
UGMLQgWzclANpuDUxTh4hq1h6HM5zpYcmpi9J1nH+2+9pIWQRNCM0mt8PnI0aigU
3+1W1Pu48UI27BANGtFOZ/EUpGb2QNte6TNFUTjOUNC1Cz4Da2JlLus125e3weL9
8XU4kHm7KobpfyFGh1Ep5AG24wUGxdVVJQn7m4zNE6g4XV5mhO2BHXqfiPj6nqOW
NHyGh54dnTdm8iJqknVPO+h9Yv9sGpjpG93Lm5SfgIkhGpamhDBcxAjrCoHfECL/
sPbQ8OVOOXTQqKhaYPN3FjKRYeTdbFYNH3mINyeeoU7IJQqCgoreSlswwSfNsand
UtmWx4AjSMfEaYD0gbdoBm2q82B2Lbif9NkJkEQw9o411JTKdaX3t4T3s0tWhPK5
dbZG20ZTFjeCLO/J1hDMUptI6AXvSaDYPYtJHsd/Y1BJJUzBuYd243vOpBRbSWZy
eX8NxSYQ35nd+NP7eUK5GoRBNBwv3Xne8nTqR4H8WYHbCiF0MuQE93bTcj/ku2Gs
jpL8B+45zLmk4X550DFYtmqaCKP611k/SwR1Xdky8/yDYf0hbeE1LrwqiwJGVqkX
CKLFsZt/NTDhHmmAzS99aF0BkdWCnaQq3BNM2INLeKynStoIkvgVcoyhLDH4w5+A
UDgU1GMSnr5m9vkcMiuqOF1KDS91VgTgy1KW9mAYimqelL69LBUqpcBt6iaY9fUw
vAuRNr+KwRvgxv9JYEG+yBFih6vDcIArxP7QrNtU2e+eZht0yuuHjQe3pSCY9jih
dzAzskSkaRJ3V4WqUsRFq4OckVItDm8aYDtaiCjU/rBH4fGu9r1GB83u0szSuoQw
JMVzBWt3YCJKxPw7wAUTb7o9Zk3kbmcHtbIB4tt3V3X2ngG7p3tmHTBbOFgTKFJq
EW+sQvEPeQw4dn2zcpUGh/QcfYqTs2Z6o4Wr/vSuRytWoCSIu1EivTIvBGBlXHsn
fsplib9NMaDB95dzdJ6MWzGkcqiPZ/9x6P9aHfhBTKNTnRdgLGNFFUJrxZpD0fWL
XmtzhgEhTc/zcdLoUDBxk0D4+kduHrOiTGDHqJehVX0dvFq6JVXLqaU02o/m80wh
c0eloGlhJchypPUyYXk7mQvZAZmdCAJ6zaHl5teJ1ubdyqMleg9bD3HmQ1TO0cyh
d9mFL0He/ye5SU+QAmmdZej2arI2gNtTPjEedKyw3KmowyQ+khPU6UFy/R50KFm/
/ObFH3+ZJOY+EW52cPfUqRaKVvJz3Wh1qF1O2akUapls2sCh/UXVAtcH3PxbBZ7A
QPuRjbbcvz6aYTdvl6cUbs/XjL3xwxhhRn8/p1CZLTIQMVEYCITPGmDuJBKg+6r7
Mv3nWGFk/8pgAZaq/Ic4/dvFYoVKUj+hchjCno8cM1cGNjeNeTVXL+0YnfiD+3rB
Z9MXemomcP4Vm48Dg75DXAbhr/1F7Swn8ZUVkspH6DAsezy/IyDsBNowm4ma1dSI
pSDLK0tu+U1zx3ui2sL9YUFtuwCHwf+P8sNzJqFztPFPE5igsYkeOxGfuvAf0zpN
SNoQe4Vgjvx7RSxX8zCyhD52KAe9urcpylLWzuXAFJpmujHN/hy9m/MaELHFg4Vs
+PxKwvDRde1WJZRkZYESbon3j73OvU6c5xR07LKP0AiQcdGafndi7wrAZHa6din7
rZz3J8NWr3Hdu6v58qk3+w08AeOFz/wba4uLd2x4h8LE+XVJ81yLal35oLV6ocYo
7tkt8TWRTO3MKri/7J+NlayrQToIU76ksttKgDdWnDVNEE1+AhoRuLo+zn6f0oER
ykCaKke4FofW16ZIEzsqNtRYXdOMJmARNTZNhdUWG6Z3+KHu3BVlv5q2tnwJfdFk
wMe6QHb8648Wm9kSOluwlox8Txo3i/Hnk8W/rsOEGk2Sf8mreizh308+MvvrmFkf
MHL3c5ILXpRmJKlhUP06aRMDyt2QzlC0vCUgVd8U7crX2wxtCFLcrS0lZShPRD6e
foG4zSE2iSTqGvFUyjuNCj6uUhA6Lemdj12BxTCKZ9d4NzRcLBfpQrYdXIxzBHPe
x464uz4i+vKtpi+eAerKfRJ9mBaVA+tLQ0ZTk+D4r2ARUMb8gq1U5gjGqHT9bqk4
8Yl6MoaL2ZKacbGZvKMLjf/CKt7NFGemAB4QA214F4OgsUazlyv5tbiMGBcdB00l
gzcIbPICJJEy9jbNavX2zt0pPfDPfyc7x5jnRvrir8soNKZ/j0YF7VdtpoTgCDVJ
CMBku9JFb2k54d1cs0Fo0m9FNuz07MQXBRB6i/GcwKncU2bsLSgGLJMDEfyzT8ZQ
y+jmh4DB/l1iQPh2i8hADXWPwyK/aXXae3LIjn4aptWKvQm5ClGQROb8zaRMvxi9
gQgOBlUTGRTMaXjZXjLded3Yg1wh+ljhjbhirX94FQy+oaAHDIRYclCPAULrVER7
YXrlo0ieDemJqgWaSNg/Z7a/hRmRS6WAjRDnjJgpXLQxD4WMXbNwIpxpB9prIrzc
vw12uxWSs8npjBIKXpWCoDp+7xwnvy67gcGqposV96VmrS1694ZMp1REPnj7Ya5R
lFvu+u1gfH2BKAQpcGYtIycoJC/m/EgPE5hL5eCOwdjqSVF++DaKllMX53LyKlWN
A0lBZzeEcOI61qBwDsSK+0x188N8qJrXvUGyRm8AyyZusAgRExe45M7i4SPIUq65
CJLfhbzWECXXVvYLUnzqBRwwDf2ISG724d5InoAvlG4f7Z2B6y0IFebwrQAAZUBF
Kh3nKgGPqIYk+eh6w2CpFRShy4Bg6SM9YJFN4lkUr7BLsJ/fGTQog0VCQF1WTOpX
x0/t5loSQJ5frUryhnGHq42MzYMYjNKhoUK2dH7HkhP3CYxWIgRg0bbe5t62A6IB
n/09NYxL5QGVZ286igtJyEjS4cyCEDdyMvPh+aluD214DGYjcxoNI9VKiRlhtV4u
m0GXkU+6/LhuyPkTUKqnVy8jhVXu4NVbJDyJQOZCGF/Rv4znHCToIQIlB3lSmpqm
mnM9sOxDUmFBF0xK4EBR+W2BjAeQGXdb/Cjiq0fhuTVJcLs2A1qUNAJjvneQAbkU
Zpiq0b/wuhf0XJ4f2mjhIU7XWtSE4DltlpyTPzmapjI1TSSuZPBStJ1LM8Q2skDu
KZk9qo5ITbjVBKOWRPwK/ZZh30Da6KNE4ihGVdaOnTKFrM5tAP5gyOdIoyCltofZ
PUfMJG/WpWB71wqfFRKjcm9Z5TC5fWb4eI7WaANWQTMRbeGM0pYB4sjpexutEC92
XXoFF/2MUW9fjUypjIJlb20nBMcVsWDKzOhJLdUTCr5iAowHZM+N54iC/bcPSnLI
AxxJCH4QF0I53OY1gO7co4+IhfN/o3eEORy/Ik68GmMFgHbEKIC6rGuRl+aAKhTm
h7QZ+L4zcofd8bsVv/kr2YtZ7y0vEbxTvv6++v9bO1VCJ+iaR3c1af9BvuObWSWA
giw5pN2mJOvVcHVb2Damb9baEUJwpamgK9B6MeJlDPGu1RqVS9Z5W08SWCCIbGSO
z64CCP46KAhmw+Tt3gYeKKJLCTRw1OGnD++na1kFDqurSxA9ndwp8IWFkhCkRa9p
ax9Rw7k/qCFr5VO+GhCpRw1uaxHvNi9WBWSVLCqweQFgQs3CLA4aYBCsqfMfjgcs
sjOmOoNQpUxg4lgmdR75nulIRzHTskro7u5LPSwCccTyqpwzyh5185Ck/bjPz8Lg
c67lDzMQVrOQT7qpRhianHuG1AoY06yZHZBVpgt1xHlX0mtG5/vRQqSNcLFfYJWC
MQY8tcxldcepo/prQjIg2PZwfoCEfr0rp3urOuNdPhUCsqqEvOiuKrR0+SdM5lin
L/kpax3pa+3RC4PzygijG5zhvsc74VrkwPP4NwF2dc+99M0oSk6ehcgV1OuU6pWx
nZ9qd9JC1Bjvp8rlvSlSs5sbF/riBSftB+XS4w0TLijRPV554iYLipdq++3r7zTa
HEWbzZotdxntGPuGgMulTz8br5/QgPk0H1+QQewM0R3x3DnMC+SRj6o1JRnv3XUg
OhfjeoHVDlsEWeUhdXVcvskMeGmAt1Ax1Um/TT5bJnW8Ecpz1+z3Vi+gadQ5sBou
UQtdxPn9lz6p1eu/h2ViaiZLVYjO/gBkCXFqXp4IdBBk07jamo+n5gnPHNXwjW7T
FDoHYY9xZiwrGgwSV3+Zj+Hv1Sgj02Q05fyFiNC/bEw76YNRl5Zkxs+7gCRbl9jk
o2IxQY5vpeE9wJ/S6oGue1CisGg1pDZ+axrNjnv01jJnF6+mKdtIxMAlIgBardQ2
MTFmwolL2egjtnsjYP/fHz4poEpIxaNaSd6QYBk2g1FT+GBE7LX84LPnIAB9JYSp
oBYvMVSMLbIwO0n+Kc2HQ5isExqa5YKNw/QFFaZ4R/41ON6tZLGuZ4JLf5e83bqF
02WB28PmbWerDEeGgwjjbkp9e0ZZui7xV9h3R7cblTtLmH6HNR806BwVAnl782zC
1LfJPjU3xoR8R8h1jJs5vS3bJ3KM/VQod6YkgBrXbmtlpp2TSpOT9PtgqFthbO76
xXcwZ+B9XJEcnsSXJAEVwcKOSRWwZOF/meNdsBVB/lk6aEcejE656vXvxh4E/sG3
q0ZX2YYaJq09TpqE/7DvGi8XjevoDOPylhjiiN8juZmtkNkY+1e9RdO8k3SdDuqp
XY67Y1RKrFg2jJgfWl/sj6kkoyLxJW0uTXDuFOQHbtoWztBoT1jUv46+cIorbtWv
dJnzWZV0lEWoR/7kEDzobDgd1eDm/FnnwGmgkZaDCiyON4e+A2IIVei8XA3LiFGv
obgvXr3w5xltIAjBcn9WujlKqzctjL1Clguuefi8lKyd0d/khv2THqstSvRhOW5H
M0qocqYowXMi210CBL9okMa2oBn3/43vfOg6d8UNKVITD3gWLh8cXD0g5fElVHej
RnjBG6SzRVbdZwjEjrohDBSdZGPE6ZWy7ZNrYXoDTzmAfo0JFBTaBB2KVfLlUon4
c59EIz/rstSdC8DHybcSYwau704+wUk/a9YCou1XIOCDQkzbGPxvZiDZmNbxao07
vU7Tkme8gWBD8ZA3LX85FHBNOpLnukA7fZYqTKl4vEkr/YbE52kPAsRA6gT9jKj3
tTykHVtUQrn7G2E+x3FfMEGaoH91K1/nHGzy6ze1L4zRApcOWCrLMDBEu1prM06r
MNY1WiVoNQY/01MwC3oCqz2ttYe8WCCFrMXNhBlavNSnUXXknWqEmGKX6z6ZC1Fx
mtWDc71otHsq9YhrxRG0O2Jwc3ZZ/Zc6sZYCBn73dHHnbzMXlqdFKqZDrn+IEI7w
YDYFxocu+fedE6C4LFo+rFYYm95i0Nx0pOdpIcmT8rAcQ/ZYz5I7GA+K0X48HLPy
Dvl1iJHXoLJYxZkRgKkEuJnDj8Ce5XGT+LMUlQDZxvSYhZoonzjbKwW+1YEwmTXX
q+djanCR6Ncif4iFejAMJXcHksbfKo7ESt06TTDVQYEblUp6s2U6H3LPyWhpn4dJ
X+EZsx6evSzNSnkqQMnj7WbPFN9lLg34xVaBA/lPmlXivSYvhq7lXUU9OCPLK8Mn
Y5UzywL0xYsCL/rb3SxZE+g66P8kYEVingqQ9uPDFAT58nQcRONilnEXz1IHWg2o
fL62AT2NvV2J0T34G03f7g7Ty12OcqKEnrYpoxHu8V8mkjaUL8FV/WBw6Fz5VjUW
RuHQV7yz6v7V9svuIXBdXFIQlWOWoN3U+uAYzozqA66A5bgQLACvpXkLhoQkAyUg
uRRc2LIgMpL59DGKkVEvAIrh7ABtM0gfQtrfyN3egLT2T9AXbL8jc0GgaMxrKayC
Ev5qtPtD7Q6Zuif8rkArfp8HoRHCnse9ts+mXDER/rLc9Ncu0QRRLGarXlZFpNU/
oKBuXwMKpYYrosgr3VwrNpnI5I/HefEupMbah9Dv3zcFj6M2JmWPGlfxOqmoOCev
8vhPxA4D+2h1+3SBflqyKWDd4II4ezJNVEUEYonWC6B3cuJbKv6iAoKRl4tzK8Ru
jLr10KglhI/FXu5GDAeALTsOmWC01uG61AKBQ4gi9+fPWl7Eikzb50HQ5g5j+gCz
urDg16a7On5/CjVyXpAC1/vDOmlD/BbwWz1yRaIgdvVtQnWYkZe8OeT2ZP4+rY+1
2k+TmSLCJwSE5kUjZwRWP6EYQGwXOTvAMjE2mQm+UYhl16lJZQJtTm9aQ2fCWNlR
J9N8v+BSSUiGTk6nNzRvJE8yYJVaCzwUvuDqi4+QNpE1QE62pYv6y2EUpOLJRt4c
pbTmUZR0yrZz7VcSlhrE9stS8ABwhiDkT87zmOdvMpBj1P33V9wa3ntSTvaeTzUE
wta8P7EZFHowYzHvjaVSFAzKLR7fv2x9d+HyI0jrw1e/WxUPPZd9bZNdg1aRT0lN
fiQ9p38LkDLGED0fJ9tSSukC2lW8efkcizXPOQ2i777hvPeXomH2Uc3rZvhFnWk4
9cNuQoa7ZGLBR6xy2ABkT5EtHvgHB3RAASO62/VI+yf2BA1o2KdGLWCbSwUxb1i2
XEHURgz+aUqZfFom1jZEXIhziriil1qK89BERc/c4YWO8lBvq3r6I/Daq3sUKO97
Yx23C50uVe9IbHuo9+s+Po9I2drqvd22YPxhHcm2pXKpnd9tzQTUlZ4B3+3uJFnD
jl5peiPyB4HYUlFv0gixd+y33OxVJgGA3kPsZbjqM/vNyYQONNGthlPOC1zO1cEi
XoW7mZD3eL/wZ/wUg2RntG2nfz4zpo9t2ygwIxdKzbebyFVNvH2NYeD+GCpxXvzr
feCLcozBgJvA9qv8IC/cKtiiXhmI/82N7O1jNdbGd5eTCRPHbBW0vbgCqXen/P/J
w9AGBh+kfft2FH8kn2EQLSfkNPr60sak0SprvU2286+/xJEoV2lGRbwKlxweHIfF
bQEh0NQH1ZIjGvhPaL6Odr3g5MTnLOri1cazKb55TRmL175CR6Z9ZaGlQYhhied8
ZgWIZ4FGC/YmEwSZb+rBpkLSegqe2mHv0EGg8SkAPm47eFednsg6Yk3c90k4KEjg
U+oR9vckrb0AzJL2/E7Hbm9fm6q7QHDUSwOzcq6J4Z2Dt7aIuxgPzx19Hp098nFc
07fM+HkpO+KSxDOFj3xbyGkqWdhAo6OZy7c1NOp2VskzP7q9D0OgXRGe70lYHzGw
O4uflK7DxRgX8bv4nRkyy5n5JRQtxV1t+hJHrfQy50kTynPo8lLIg/u6nAzKmFot
SDBMEE40974j1DpVnrvTR62dcU47PQ5WzFUG+xl/pP1UBLZ+MYejr9WQTWqqc9ah
tj5pJ3KCWAQGERR59it1QGMZfo0yZkTM8n97uTc6EUV7Lc5GCcExhAeDIC9LA+Ze
MpxJc+UCHvzHSxek38cFocsw3W+W5xnOrmn9nDZx56o7Pnlbw4cKUu2WAIjC3biy
0o33AYAzjYDXi1HldGFZiap6Ico6OhDx4gOEzzbo48w0jd/8ngKEyfbLxoc8pBPB
iex/Y867BThe+hJnnw7VRZd/NXdSl7vnjvASECQsJ4xW7/v1SB3CeYv9NaVB6bym
5qL7Rn2E+HlAkqb66pPTLEIXezwVnFA+PB5MQkJ66ROuFAzsqEEVyZzzX/WGHF/M
68VXmGAKIBhdyYhnctzV1pQY6es/0WDk0pqGNe2tT56z+POBZ5Ad5YpUkom6tNKx
rgDTeVO9oF7+/5mlWAjVWp8tgdjNq1xA1SgiMRc0WZ3dsCuy0K2J9yhD0lmyHJy4
PoDfzgItZQYiitks61+w3GVjIhBJLeQxH5/QvA0Rb9xm76s0za8eTsFdqeolL4h/
VbL+bBHCtFDzu1v4eOJY3EycPLRd5PFSpkWdgQI1ihr/uDB15FdrkUoyshsrHGVN
Lu+1kZ156ad30oChPshPUzfxYBUXdoEGsb4LQ16TCMkQzHE75zDmWG7K9hNLFY4L
ZAtzNQDAKSpU/G9YZh0cViTL+W68vmTzpVT4ls1JKeAF6DisEtIZ3kP8dj26tsGO
uFYnp2/hPaHeYI0HVrSv9efezEcx61JoGy8+Vx/NBKs5Xo5UReXEPned/mWILnSW
QukEVjA16G5qGvPdyyYpXxHZSHGVrgEAYLEpVzszCsNkNcNU50gd1IPrLBJFCgfw
z/gX1UPqrf4A7hggZBNDMK0prHtCml2/rkm5JLYfxC710N3O99niPHqJ7vmaWmhT
453+BoAzAcEmlHT6oaIcrIS5BVF3pbyhpNg41uIpKLhZbrNBjHB4WtiqWUQ3IgHP
IyP/07LvLHhgV6nTN6Ik3BFC/utzx7ZN1ZDocP50xUZPKQ4KxNw/uTaSCO/Tgq+l
aAa+G4UqvaCTpeiPfLgM2Sb3tRhKdQX90QSlVETwh/UWAhJjQJu5g1gFro7d7A4J
WYtqqmfPNZJ556cp1Nk1X0e4B2aiAix7zP1gAnk8ksF0x2+WWeN4i+Fq72SF/Jpw
zOO7zE3m1uod5ISrn+axmCZDT/EWZBtAOgYDXkEql+WCyBYVH3c81NopvQZKZjIW
VqzW5gdqJ0mV0C1SschN8ghx+9cJONwjqDkxPz/vxUqMiCr4QRtu9sy7XbNoPCL/
Dlop4GvWMDTi47L05m7rTn+mlPG3/XHjm2cojE1I7qALgHMBN1aJofupV49DCKae
Owz4U+SccZ/Y6MeyfN/UsJv3w4s0tRJ6Y4gU6S3z20Pp/VMOoYwhWALuVaRgr6mU
4YTJ2O8MgGTQwkgPBWQHoIDSZpxKo55aUL427mJvWfhouMRqGvrU1KqDdYgd5DsC
G2SNFsFvbp1KhluCfcYFfKK4tUIjKV4YVIdAR7/XnHjqw043elfb3ut6XX2+5Ql+
3/BVtcTWQSOtq+uCms/MKw9Kg571ClY/z1gu95LHk6aid6rVtieuN+ufCtZoJnTn
OTAQkxaj+xc/DmZAP+6pa+c7mjAodG5xXChJkrJKlkTEeMLZx3EuAQMBqgQHERqS
WucPInB6QvTMAtM0mi5y7p97P7MClvbem7qs7XncpN4Qgq6ZbsZni7CDwSYNpe+F
M0y/eUHJErl+jvSgd6RPwFh521gJq3sA99egup2pm7T8a720lE3/eNgflCpyU7F9
K1Pjghrc5vPPm61mN6SK5qpuCcjzRri/3yVSg6H/CSTeVen+qjXPVhDiW0VwMpWr
UX8iFrRqwxpN4biEfsHC4Yakv1/YxiAm1bFoYjb4dSDs3C7wT5iDKrrq7QjvdtVw
FJu3edOFSYlGsYKZA5+3hA4qOS9pEHCWSxCD9BudH8F3Yc5h5sbo/fcbALdedr0M
WlZZv7x2u509U2ILDRHlYX3UUjPtrqV0GtKhjNZ8ShReef9LnkWceQSyMX1nfwLF
WLtMpskJxJvyCaAeeTnxyQrjofy0PyW3fX9FD8BWLIGvoe4a+xoo/DxUow8fQ8jh
JUMeXv4H6UtSatIL2tMFhD7wEg4Cog/stzplpMli4fNqODzNEi0Fp/oktQOI/ZZn
EQhj8szcaUTBZeMNBPDRKapqG41E8RUHMlH0YCepUaFceAeysT64XwUAfWDEYzsi
7KxGkcLEAgtDUHEbMoPySI4wD7kZz3oSbkcLXO3szbTUwyXBmh+iPCRuULZxF60l
7Y6g5JYrFCoyunM0UQWUijQtBhCNuIdoPnbigK5sWuSbXgJBUW/GvEzN/I0RGFKw
5k/Z3ZL66tshZFY8c3dhQZQmLuRp/Ye5xcItSxNMeVBijqq381h/Gr7wBmLbf+21
PR0Xo5Ujdw/hS4QkzzBOGqm0WVGg4MXa2a3VHqYQrfqFfoIVMPBhQtsKQlV7F+ZV
PgPHxdCP9qgSE7RITSmm7hUsB52bP0/zc/66Y+JPMl+KZ8JqxXEdk59UWSIdSnuC
H01fRcnN4jdMjDwghj92YgAkkcqGpRnSTfH6fYifmuwODD2qnm5z+dkfiiVgffOm
J/N7aYMXTXzwFVXyvHE9vJya3xCPpIV9SOpEfHBp5DXoW3ysT2cPCKeIgvICQz0k
twRWU6825iGBxgKe0XWepFWsyadOJdj06sHkpHFQT41WTrxpyB7E7JItpfwhBquo
Sk5MQhiXbngRGmwWwEzmqeMww94fu5iYXpfHULFfH+h0T5Abgwcq4aK7twwUodiH
j75V8KuhcRcVWLhNL2nEHUbetpLmcEVBL7JQWBfVWUpppOnoJ3oQr1KY715HQZVg
wJTV6PCAktqRIHM0mXn+O2rw+NPzeUowRuDW32eTZX/0eZ9I+L03lvg9cQqzB/Fc
0nv9VqjsrWhG3ZisJT3P5DrKAhZysCDpmWMIiz1X2H0OfDpakS0pgKTQwJcEJLu4
6ItxxUDpZ7HOE2Q6oJGlVczmeuDTgTsRXStohG/FImd9bQ5suEQIpuAfY3qPH2Iv
m0L2f8Vw060m2waCdU/BYvZb+3c15PtJ3sZpgLUMUIzhUhMG8Tg3sdm/B7yMHAPc
XIME6AJBJaZ1yb8o9fgVK/N7hH0pfNakFACgEQ3/dHLjCfA99VISUvGLqoiBPjGT
ZOlKcEoggcAwQNKbp/1796SNoO2+OiFG20WiDo1T/JVfSmiaKonkIilhFq3w2/qo
JRjLUzGXP6zDfh0xaOPqR24/0Js+0FPKs7RbpCdeva4fk0OYq7mq7ebu5hnDTrBW
2eglFGq+svsgd5XMhiYO23FZxoXk07csJcMBYCpZL/Wi2vdppD7I1AEyOBzZii1+
zsGEwwwo37n8leNzbwYPwKjlw0szpfT0lDlGUS/oB35GTAd8lJikP0J3dbx6m/BW
BZCWaIXecZKNHblZopLbargtVD0+t49K/0TdxdSYVLSPozKEX+PkYnuww9lXgGz7
8z2nQjh57s/Nq3rHpv3hSUnNg7x/sxWmyHpiETtVrqDJUzrbfYdxpXTtR2UYuAx+
LKeeZqBdjvbuQNxOTMp54HeggzNoM3THDasUYnLe/B6jYesRNC8k3tQMkvFrzMuB
Bs+k4MJnK5+CKLDOuDAIc+Gp4WzskAlch93MDq4QPX0pWcP5M54oKAmFKxrQ5+KF
YvvA6aKOO6Qp+DkWhvOEGLG/pJSuJ4g3gME0SkfuucyUAyschK7ariS5AqE/vVCH
0eZ2qXONjvGvG3UupQ5vgSB1LpIMTPwUgpDuLLr+23mrsgK9in8JM7/eFtXk/pQ/
0huMdsPzSQdV1onL6U97sRXGGu/8fq7QJN+cM+c/+u/8xe3bl+FofdAmhN8Z+oqj
N8gNTM8twN2EiOqyht4H8S7JQiZoroOlBIvG4GGCvCl6CJO2EbRSbhhy7TFS0hKm
pn0Xv7UEeFcXcJ12rzYPSlyy3uiHbrY0ENQ1dtx7cG8TOQC2Bdbs1iN0Fz4D5ife
bVFvJQohofOWwc0VojnUfO8MGn/kHy6m45Qppga/pzv8wq3AIe0akS9Cig9VDnzZ
Tn9uA27QCBdv6OO9+GDjF9lASsFTw9un8GAzHLViR1fostdpfaA9P4oYMZRyLLFD
FUTCek8WalX0L/LpfTgZGdG4gEiyljcUd2o3uk1y5Ta9lOuOcM6Z7BdIkLZrpcYw
FPqteonuJNCi/P1VApgq5yUho1ep6SNQoEVO1FzFx1l31M2ECAw5q3xTdnytO9M/
FQ3qIXZv3RaVaHJDD9eTS/VehD6SLlXF7VhDFn3qJGyzXyKyFzNQuMoabaJeXL2z
mqwModajxl+ZW1zeITUPxJyw61bi+0/cGgHBEv0manMELknaK6r8gZVs6R9bSQUM
Y4lKCdSYs60P7FZHs+Y9IOcElKFyAb0qfDeshd3IbPTH4eiswHHLQ+6KwQlud9qN
f4uNjoO6+FsT1kjxdn1PJRI6cHavgWtzeYOLSEgVLAlMedgiRHexmJAZm29if7b/
IYcY1bdjzzlu3mjH7GjX7oRE5EVXrD4vKbuz8X+Z3GHQhY00S7+PwziQcFEPFMui
8ORunAVX9opVNpeuylfR9t69WMj77f0RpSAqpOMtEn08OSYfXUqaqkaMPf+uhWt8
IpJm7ZBnTMVv0aiYT+1U7yhOp9D1YI0EbHSn8z+TgimWw/JWUYPeoc8NuVmADD6B
y5WgYCKeMew4r8FxLnwqfSm/PlfLjDDiQ4EEfrzTxUxnGuOrJGu24POBi2GoQZ3d
6X6RDjTb8llvnOgun1qtQXfN8cS3ZnqVH2Oj6SgJkiu91aeOLflRKrmToOg3XZYl
Ar9wb8alGfDh6dnuOFBF8sIqJc9eZ0bxZ5OXkp/JGtOjFz6TxnC7/Odba0m5qVYB
TTXIMDqjkaMhocnunhxZBR9AOZKq4WLHM69jKIIK5iCv1+0lLXROK4JWn6oJFcDu
4H7EFe+T6Dvo5nf/Hl9RHp2Y+O/Zc1sCzFhh2TglJfZQw91RxNbizOl93WCFM3uH
T2mhPYAFAHXPvJDMVRw0wOik3jT33CSfbtmLjnWkOiJsvqkr7wIAw6e1oM3HFH86
mpsGeRrvjOmipXry+YdTPF+nGOEv2xwOZ7qP9HjmZ4m/Pp5JocCBOXEIQmOnJKDN
lSz6/boHXKzamz4uxOkyPEsieO7iH20n6s1jIZ51XxAz39uJhqEiK2H1cO2kzpRO
Y8enj7+yAlA8A7x2iYNGkMniz6a17dp7lq5B5YbCddmYtfgNPplmmN1gT8oSI1Xl
o2LUkWQYG++qCvA6ayDV9Tb7Z2JqGb4I99Hy8dZ6MV7Juhd9y359kNgiXxwe+E45
vH8Fnle6PvdmQbFbrgQQco7JGAzyvQ49SBlilqtqXHGdDg4YlNPpq9W+HvM5rh75
27adP5d0HLD0silnUB+dNPy9eRSFyIfwd5aT0bN3fLBJmCIyLL6rh/h1/4k2il1/
zNnWgimjyR2/D0hopxSHrpamwCuHTQM01dzHu/NivZL+gWdFA50qDNzEIOCH2Nj4
7luAlVP5xwpyX6iOvCEIH4EUERCKThg6EpomUILzkjNWCYGYZUmKfg3XDt1tzuoC
i3QQ1xnQo1f9jzmQd0VD78NaN5xnDnjJG8agoN1MJbmQeel/+i9d8iPlZ/AVGctU
gY5HHGACNs5JAJ9MjzGgSyyh0xSJTAKeLPMcgcn+p+jnvUzPbDlS6VxA+jG9ULAE
7PXBQy3t4PL9A2tZe0XT0khwwsfE3UKlLcAbupcw8rGW6FAKuyQi6IO5oM8Bk8b9
OAHdpGohNpuvoQ+yNBKlkNKbiD+qxzadV0oaor58p4A+TLqFxUVawY5JhBnBVbqc
eXFXSFTRNkfNASA51vg0o0ywU+H7wbn/tGM0yRSP9yXsTGeVV7y7umoFQX5jcgn8
PjRPWCG5pe6S+ctyICWAOeJTYX3tKO+ckhwR6bhWwHlYFyJjSS+xMbgsrUaxBxGX
YbWYVL78kx3tJIicEVgt3nXrRoXJbSKeyUFfhzI7RJ6/jUvWWNYXvdcTncNVjXxM
fPDaLu6AXMr1daxPswe5JCTtf+N1vNoyZAcGzc6suB4SfHmCUonLeRygABtZBmZQ
YuExm8OipEBPUvUC1yOuXsCnidJ2PDBY/ULYxciM6RD6P+vGxa3n+M8qmzUAiZZ2
/CmqhVvfPyVkq9u8Jl52CogeXyNpoythEtdJmFg2fT815cH1n+hXB9m6YBY/9iy6
p9SbtDd0ZUMhMX28Q066wPZUmmlJ1AjKq9OVh4L0VqLD4hBdZMfAt6KMzpV1qCdd
nJh+efTyUVS+mPMB72WFC1LmHZISwfIXPNg9p94YULadDo2YBEWY3GmsZAAiPd/P
GjP04A01bBKro47FzEXi9gRo7nvu61u4dbgu4f4SE6N6esa/3xmEWGkRXTaTMUwz
d/6bIoFwhFue9WhbZBreeEvg0U1J/kBWeeGZNlAbyn9+aFdBR3E3500Jv482hFRr
yP+m511NOAMV9WNvlgV/esSEI82aQaNeHNgrflAy6T8JZIIN5hqmesYPrPrUNW/p
3Lo29NLewUO7oGLIqEk6j1OJPgjELUrrt7zMG4mioVKm76a4wUtmerv/TLTyRQ9F
QgB0LHeJ4ulOM0Y7BnwbrG46rfHtOTuqJuEd0erftMH+zQhIKBpbAhmNDGwL3cMx
h47exMGmR9+REusITNCvgq+aPGI3qQnRCWQ8qN2Kpc3p9UY7NnShVHSad7IQZJPS
aGazHBfhehHyTfGTBvybbUToZzDdGGIFQQGykImqaAYCCDG1ugj10S5JDYn9Md8y
xPa1uav89s4jXdTodD1U/KedYq8Qsb+fQOZri1A7CduBQFj+y6XbrQeywHhBx7yC
Q8I1V1x/oL3ksx2tLzdf88vjgIMv50zG25xSJ3SjL5XdgUc2gXT9VjumehRHVukD
hjGbCQjd56/K4JgRroTNBoQgKhj7xy4BlmsKn9JvDonS9eRJgVdess1JPA7tt+O5
ONswZT+k1JQBP4DRhNF7YvhuCgkLO+rTXKuuvyLiazrjIyc7K9NDJVJkHhqyEYj4
s3qcNilBaghMfVCszyB+A1Rdk0tc9xuvI3TT+c3xCQ/mrF5ylTryxkgJ+P2sfFM3
ESKPNoC6O4n6ntMF2vfadcX4OemmMrrcnQSQzowzLAgjniO2aeLLxzIaeXP8usxh
0SX2QBQ/EgBsG6jL5PDWhZ6xbfvm54P1hdBzM6unN6BA6FV4yIVZ3TJ+GofN6HzE
DIzyO4sD0h5FHiSJYnCYmxVyIoZdSgfqRWcK1h54gFf4S/LbZ33Z3DXYXe315N3T
Quuw5gDRXixysC4QxfVw62VGGg0GaBB9ornoByxJWb/flh54daQK42z1r5yAsOJF
G4RNu3rZbautt5oS4ol5IygRaACLd/JlYldBS5321JsAvrnivhxAkrpVDmmiz/R/
CshrnQIhpQvhf/9eCICJVexAwj5lmHOil+5YTS4N6RFkNF95zGrUlKPKK3Z0ZN4k
uWnzD8bfBM3G1Ry8bNJficY3/dzqxPm4MXeAzMpyDK2qH44Hc2EUssVst6oIPcH1
NKm8jCGhkpkAmnLH8+gpxM5Gf+UPJGMnPkUBwq89azJDpqNmv5NYr3z8E8I6YjWp
oTnijb1lBi+qlNXhZeXbMzZugqNgtk+/a+0E1Z0pDfA0H4NJ6NvsLzHNVNRrXJdB
hwawZ1zcwm5JI7eR3UYkjB94QdVJ85fxsNBQvja1baSoaJQSUFzpMqsNItMfB7ml
0Fg4YFKpUpQk2dai2rg9nHk9jQlyuDAbYLkjsK2f0WhRbZWVseZ6+uGdloZXl7kn
7ZesvPqm9BuWSXdOnqJxg3n2B+QjNNA47Gk7GPsedA/oeslQyj2z5I/0hWJnNUkA
RD4alHgclRBQjnApFYEz8fl8VCGBvU46gSm9dFyHVG++KcouPXRrOBeRigWctVm1
btDZo0vdNSPaivnm2RB/cQnrPgbX14SY1RiGDovfcRzsBcEHGaCpwwaoXk1SiXoq
ia+0q7B9t4Gz2kDAzzpdSTu90RyElrP54nTHbop1dj/jXiQChsYQCPbSqJrfA3qj
q+Yyk0RriC5cVpZrUcK178c2oEaP4HRL7wvgF22o55fDWP+tbZ+2M9oAMJ3y1YM8
T12xrZ9s2mufvTcSiftitZ92v1xcxBwsQHEBcGdR1gc5IRtiyUrxMfxKWBjTRrAX
pX8VoD6HrvA5uCUKvfUV2u6bXypLM8yM/SdDUDq5rkuUcjRIeYaHPsvYlw5Ju8GF
BaAtxcELp48joS/ZBF5S0x3Gqys7cDRjGcYLCaPBbXrcHv+lIlicIwAzw8kk+DYx
cokAdxzjuaefQQXa5pZZGyVncOGehOQn2SW9qQKEio8CSRD7UnYt2u7gEslF9tLu
fp+Ratri2VFh1Qo6wcpIA/ls/lGUpuB/I2mJPFdevcSFnFfKaACfkUMFL/BnEO7p
qaoKZk5/sp5yqGEtFTVHsqj8AJYK9HKmsSo3t0OCfooAmgjVCi0pugdHFQQV3RM8
rQfMlCiqzovaabqV2DtZ6G11PSdnqb/egI1tyAp1CFfGctmE+sxqst+Db+GfUxtB
HzIeiYTRFxKO6uaRTs2vxtYymEOjqB9T2lE+KMvQ6zY4mQoF1Uf+ksbsJ935OUJL
xe8GWLCXSoXbkcsTx9q0RtyndXIPHU6NgPtlbJwBTjIm6eHusVqP/WR9P04Q9z5h
qSEGHUrg8fCw8qmd8ti7dggHskMtqo390Mh43g/GEqHjHnY8MDfEerq6O7wrak2h
+t/Qy95RC53xi/GXrebg3XISV1rGD+YxPZUEvMxt958IzWLiLUYZLQN7cGqXlZoW
zEbo83205EXyvUEx4MDHxQpie0T+MDzycAPH6/TEHLOwyjUyN2H+tHIzOjife7RU
l8gOcbWhPX3OCyYBCHaeksxl4jyUld3Sg5omqEvTfcrXhOsAJdNxkYZymfs9lSO+
XHLMrjqnyGEzf+auXVy3USUNs7gMx3hHglny91t3p7UQRvKcAvXKuhekGEM8HAPs
3Y4fZw65c1gaQOyqvlnUdocsEAUvJ8fS1EuouiSt8hbAJ3RyCC+DOS8/mOWC+JE/
JYGDSrVSLfhgQ2ZwlJm9uO38j7A3+OZPIrijbZDz43LtD0lioundG1skXa2QB7k6
LLTE2FvUTNjl3YCqxv3C8X1PGw+NdQDL4IEyT6ZF0O6ZnGR2vtkwVoV8YtmyK3vC
4i1WMjraFsxZhDXcC7gWBU6qJZyCiqm8NQZ80oSzalsvLMIO5KLsvnORTCG1z02w
MgvQdnHoyyUNNLWGhO2RTEp6r9b9G2J4V7tAoz21amOOrfaoEAXrjYIZwBLVtECt
Ad6moGlAz+9hYtrngj0o4ldLzgCGqBWFEwkXKvlOSzsSgNylDUSh3G6fW8tDYYhO
6WftMLOU1IJsqLrP3JMP0qn3yMqVfP8wccsxy0/sGLYpZ98Uqp9dAZEj2CbHglZO
useuWdJ9mmZ9fcj1ElEzSPeS+tsV3gOiuyNTdtS8F/qjR0uKyPRAlGGSRIe0TgFp
0ERHdZ8N8pPqcNAOE4HPMP1x/6AVGYoC+wgoeNf8wrzZpSMN7HvXdhrbWJbuu4QJ
43Oak1xu7cKgVl46P3umyS71TzIkSVkeTyJVlSaQyslTvdJAV2jK74U1Nlfcn6MM
xoPYOCXhD4/iJ4pmkek+OXe1PnyTPJexPkeZ3Fo9wkiLgsqSNW0xceDZc+PBinKa
UnCeDUhCAjy9uBCXGQxU3r3S5Rp9FaS3XMRo+j+0MFN911RL1jNLwojs2Mpp6qNs
4qFQYwaer4zWaq+31KfAKxXclMSfKSJW9ynHHciX4q5+7IVcEdP0bhR501c6ylR9
QB79NYGeJYhE/0hASUqpP/ykDzVNcNzJWByiXnkYJuhd9goQLHD+AWkDsC1CmwIU
LX6ui1y6RDBVuv3DCfI7jJ/lBG4mlvgL2QgcAU0xfl3Ijxzps0BRA+64wS+FifFt
TaCAnGZKJTMqFuPFyBJo8A47Kyw/tnh7Wl1r40M+2d8+B2GntgSOyyrYUkxVPldA
9IkMO7R5Pd5xq4zRXcstWyMCPhJg97Gv9cx24vGe+ruNK0paHkR9W+xeOxQKSlK4
cWN38nasSGK3whVBxYkxhuLSj1k1kLYN0VogH99lU3qjqoO4GdUpMaH2tnjgfyn2
oUEJ5i4MHwruw5rb5/mRGo2lV+ockVbutJKuoVg6S+AFiSNdfi/rl1Ge3FVPUYC4
UTpXPTomUmXXlQVEp0tsMZ8Sfu3JSzuQNO/Yu5+Qkg/wE8snzoDMI5HTPcNYS2eM
lEOfvzMGPHeozXCwDSuJr+bROxG0MAeY2MVBujZ/tqN1YN8Alj+oaKOyCCddKGv9
E055Srdav0YNPkf00wS0STslof4FjlNA1xYoG1Ooo624bmOXaNNw1xWA94MnJBqv
iJWHR9R7fE64+j4UGxuLyCoFrs0RCowKBUnMflIfmoY7dLyf8ExyDIWEDdW3XEI3
2bQ04l6ZVjWNDF/IKFoXoPeLuvFmtvt3lB39FA95G7QpeSD08mAjPm5urPgEy7we
kdGLhFq0H/ENgKRdLsIm4G6D9SLtQFGOrIASfUpsU/4crS7FQduu1Mxe++ulSMWk
56DOsZMY9AvQO/koqZN2xs7qWDYJq4aQpSx2ITcurSlKbXd4lPPQQSEHeSZ38EtU
bZfTKBJdsfBZjxbAoHLxfCmsxNPc9OcmcHGPFV9zBUQM/LPcbQvdZWTNo1bagvvR
QjSZk9L7WjTtpGvGP+eduJvA7kIe+u6t0KWhGRhHCqGFWZdRUR7w2F5WkruRiAOX
59W45cpu58j198K0zZjb8CBZzUmFHSTrwatZNSQeePuQl7wYNS52az1XAbof8Nrc
7AezclE2Os5y9ildAW8BpDaStNHjLy8/Wab3nKwrazIggt/Ooz1eBgLBKb9hXBW6
CQP5YDfXHB78l8NlZpf9o6lAt8ip7pke2F6OWJ3enktXB3n+BU0uZRxvytGn7EgE
Xe0wl6wfrUWH4Sb12AU/eIHnvWnjCdIgEyiLfARuXUzK/HMrW9EAbC/GPK22p88E
lrbE704bqO93QR5RxH3zojFt9Xg+9ewj+uT/EQEWWdPNpr1qP4yuMcIOf9SDTB5T
LZx/Dwn/RKQuFU0SZ6xyqjjJyrYMwmoEUkLzJwmV0KjyS0XmY1mJsdpc5Ai3V28E
xr1xInEoZl4w/lH1OHE3ZD7l7mo5sGFMOkiWrWaPgpFr1upiXVGNFIHCrBaVNUke
OyiWxocmD6Xgz6jiZ8i1mVospSUhquFkgNw8OKZt4bwTX0PzKGC62TElC2Hgitlp
kzVh3EEXHV61EcxLzWm9x8YMvGSR6frkCfAn8IDmFTGE7z6PVrOy2RUzhYWDFuPL
1u5ful3h5kTbNzMLoQncRBrX7CTVF+htZ3ji0J1v7w13deX+nwTjVy2oPibtORZt
9TJkj/3sCgg65JarE7ghswDj68UGgA6/YHWNjGiBgnFudKcMciV6EFwFHnbA0ya8
8vaFImQ0rj1MCTdQ7GDDIE5zuLGSd0UUxSO2OHjBg+vRzWLuDIyv2/CSjktWOcYg
DnDdga4t8Ft4LR6J1AeaoKbS6GYVS7ebfDNw5BDRa7+V2ZH6m1Fj5bjbcw8Nst51
0bC9MkZ4V6kSHy2qbATLJJesWCME5aQjiPqv8MqWa0uCU3/iY5jigOdG8wc/LzmJ
KgO8OG6w7g9ACmOf0q1uEXvFW1Bs92cYH5b5fgkXMM8MhUurzwLanXEzM1CrkiPm
WCzmDvsR1Ztmu+araz7Qir7+XtFkMZo1rNtNNUT1OZcZj/NudlUI/lGArorMBsxu
9M1nbi1TtRo/4XHmZCLwTyOwYeCi3u9N5oI6BrDvl6saxpVLpo9/OKj5rmf7RrRK
HYWZihC+dRuVi0FghCrII/jLeWbfL+SKl1h9LTN7xQc99Gw5wxWN+8/ZwBR+R7fe
1nfgBYZk6IwBbT6wqVN/WxatOYBDIsWTbmMS270xYeGQ3lGwgaa7HZBe0RFOh4ow
dsVgSaTRvFf2UB/vEJfP8DdKo4ku0wU13+kqjfVrcvpWsJZCrqGyXnkq/FsZxOdj
ZraVtmp/Q0OS7jFQyMBGg53h1o1MC+dbC9DGpJHA7Cr9BmFgOvfukQv5G3LIl0Eb
aHY/EJwNLtaQHqoaPFYpTjku6Fe8tvFboWaW2xhNaUpkcZ1zk7bPzteuW2wcOQVI
Qs+3Y7WVoAkSeo2sKwPkpEamHf4BOE/r0ddCtJK8yNgnMDJ4GyFBIi6v4r92/XO1
5lyh7pBZV5RDuY1yRixVfRigPO3LNzUJXGF2QZSNKVvi0e888ZJ00Sd9TeP2ThPS
uUjajIqzRVXkVz+qyRLiPNQugPsK46Ii6H3Hu82x1k5/IVOmhvhYWgrVU3R75xSo
PFT4PS5EvZ3xkofKbGzunSAXhAdzR1V072PoJbbVw8c+qjbwde89gUr0R8lXFkqm
8pO6Luw/4LLtC1ooOQb+0hiSnGXnqMB0DzL29l9vHj7mm/k4IzNSTNqIvIu1MuLS
MJtdcMv5HewKwg08mLAc74qoHVzVZunDotNhsZ1bbFMM24eg1YgfsU4qTi1Sc1Qr
8inX4vi8v8uZWExjjbNKWeKMpYhq9d1embD8YaF04Wqznx59nKaBqjpYXkKCQxw8
4otlfCXDMI6/ybZNtAjWO9z7iHY43kC995YyK3Fas1rXBTjczI9PSkr2sLwfeEPW
mFeop/5pTwzLkqO0KCabJ7nGWPWFA8YTbC+Xn+e4hAg2hGJjAxE9K5A2AIxrEz6i
r8Bp5tZHzQpUuIvcvuy7GOOcHvFdj7x8t0aaSM+AAu6ahtVyJUU6e0tnxf05xCZg
Gdi7UqpFJev7SocrMUmF7GcWGyzsj5ikJA/i2FvYqeXfm9qFNV38+eRpkz/9Px/c
XKDKd5ZBHFgUCfRneSVgm+/wlf1J5JLtwLil6SV10Raniy8jjVNipBUPLfH4wt8Y
rRUesettZ3RqbFd5Ycb/yhtVZ4H/N9N6zuUn035YSdfS/8Fj8mRO9wqIXUrZADkz
1H/ejdc5VAC40KlBS9Kf78I/Mau8/mQFyhGYkQGNwB/D8fWSx1crutz0foMwCszX
mxZD7u0il3RyLJwxfOk5UrlfRdzIZadFE0Svb+6nikvA5ZZIJXQ6hpphAn4DlfYN
phd46lnfogilOBFjqgAb0BFIOt6aaLfmuRoO2hyYe/RQSIUO1ibK+KBIcaOufubA
XDH27/3dsWUN+fXGDWtlZkj1mLbQj/1InXzJQ/8wlfw8+2UbBlWAF6sO6o+aljqn
aDkkEwYBF2DPSgC1kL0Jy/i3VV47oXImiXe9hObPkCdp1c8tGdhtSCN+X2JjqW1t
j+ybzEWEGhIl8R8Ym1UCMmYZ9uXxbyWkbSaUOQEWzulEuq1TiG7X6R+bduNswnhw
XK4AE61G1RzJoI1YL31iVcKL3lO950C7Kl8ODbTYtgqdKEsY9lAILCvKLTq7Unmt
fyjcXH6I8ahKA/NDWfkSbJSRR0zJwzUHRwLWbibTaOH7C7UffNn/w009PYMGiGyZ
XZm9pF1uijC51fWv5c4EmRJKfZkNCkdGJgETifrS/viXhKY7YbsT9aZuoVBXzxw0
G8/XL/WWT2xQ40Vo/v/ON7RZ4i76JZPDknveUh7HW3z7QibXBwDukBPkdNvqZZqc
hSHfLcnYFMIDiswanDg2YHb9FKqNjQ6CtOL/NI4D/9Va41DfiM82VAnSx0JidC5R
jh4kt2D9ehl8XJ/ttttnSKtBzBLMO1yU3eM2uAoU2z2kiIi2Ns7fGIPbnKrq458k
Y9BGwUGUy5xekgmznn1Rgpv7nakFtWZEng2M3xBbDiPLBL/0F+i6QMLUVuy4tSCr
aYBYujEGHJCigQMbSAtAELbm6zxGNchu1otN/1OGQ7GUCu4aJG9yIiuycqqdQnQw
fDk2NAmovs9H6+vJwj+08tB8EGTrKKGQ1mNITJJxvMHt9ocXV0HgmOtSfn8SsR22
gdCJKravnaNtxQsEn9W2BEUVmyRSByaU/Ir8xJ2kGB13qx3UVhxQc1bPd26+f03f
d2M9z43j1aL/ZZUXtqGSmccWYIEakoCqJ4vKYYT38efFbbxHLnryI35/qOpKXgrV
fkoBcdVmU79q1iECqt/qmbsJVZgL9pYFwec6pFz6pEo8hXseyh6cSP+mfiEnAzXY
MdiB9NaqFBQ6/PBhfAseIC4SlBQovij4I9HQqfeDJQ1XgMmKa8+btM5xqHYjlRie
bJtffpr+cDY5UPKrKRHI326YntRd8Zqsz/AnsZqiYQlhk8yyn8I7ZNFF2WuDOnSR
dOPTfmIyMHRM8+tolMkqiR2mzxZuJk6Rp5FQleHspApQWr1OI0cl78RitzEym3+E
bwKbu0vgnM89Ctr7R/b6TrqYicmjRupk3TElixya6xPvXnWOCwdM/jWEwRELN7Xa
B0N2NovPTR2/wOcZ19mQK3XojZlyd1ncJNTOn9zNfizcS0zOqBVciOfGxU0C1s5c
9J2FPB1FD0QTCMbZRcFMB2JZH/3rUF3jS79puz/h8PikoMX6/I5kxFVVdzZEZ+PO
GAHiYOfuh9iODjagm4LiTiRQfmgleNyA7haj+RrnrVQDWWMR61zhPjq1XR45DChX
l3BcCt57OsfBKLtBN0VNWAdBbb4bW07Mt9ckjPy59i7po0DP47Jedlvsi6gdkEDZ
0OD9mWsJIbdM539gPCwhI1CVt6N5oXxXMQrECQJZzim4Zpq08IZ7sV7RjwNVCxkD
MbO5QyWOs8OurqDzKih4JsN+HMHTandQw8x58o6uDj2Asv+C35B/jVn73r6VuJWO
Hdkiw/kpwvpN3BhNk8gx6EbmfRNmr3QrJwPheF4IG0DgChVD2TUNo9SjEDPEpuSO
Y1KyOTzEpj5TlmfoKJGzting2gHXD1pzt0QxJ1a2WDWdd4uqHZshslKRn9jTse6z
j9Gp8eKI6g94vtOOeN0PwLfaUowd66KIwTjFedH0Cgy6DlQr4pWkPzd4G/i9RiDu
6XbM3BWNUAQS0Vk/Qj/6GP6xyFgGIPHUUaEp4TSeoyHl00qHKSOmBClfvnobfuYS
Vjgqez37sOIHrB2OoR1saKqJr8HDnBc8yu2aL78cty8WUUnSFGxIiByXfzKQctgZ
waCVFQONBkEJEE5jSrR1lKvIpRhDpKMwlbvee8Qm/idp6M72yk/5bqoxmt/429vu
iqoULNsxpsXqCwvWsj0dRk/VsT+mel1tc0nLBzDd/uYGFvPgUnUKf0DnGmRXRcgg
vT5o/a1tqzVCWfwM6+qNZiZUwjMqAnYdCjp/aieQnZuinu8uH+CAMGlvZoFRtg5z
1BolMo5Veth+f8q5Dej8eedTFCuFeDnyW/JifeVFlVwNZEavA7xl2aJo/eINS3eP
wNXXlyRQQR7QFO32Vm0PXU6LYjocp4F1egMgHXJ8cyHLvQOlX5UCnuV/Q2r/4F+Q
z4b0GAQFiU4YtBg1UuVdVlR16JR+OL3zoJZFcZZHg+g78HVyplfglmORuq2HJw/C
YKzboht1YrSUJdjoupBsWvZhmia707KpEaXsfDfh4gvLyPSjsngqZni3No8koz73
gIrn0GwxSMa2Zfh4QvyT5Q9ojRFIKGNV9CNTXGeRP4UNDjsKtAQRs0aszr8nD+wN
W8Y8iIS+GpWI6i7di54GlCSwvG8aO8ngL61ZZSBzVaISdasmXEh7wT1b/5PvbGNU
gzrL34KEQBWDs1gjEiZrqOP+50NkD8tN2ZL64j/7KK0z/ESa+CjNO0JFXFRYHf/8
NbhmBJLkafblFdDZqlH3DiQ7EV/yBFtQsthT8FF2XZ8AFyuZXE0HSI1bFkqkdF3V
Td/izhRSc6Ko3/a8bsjja9zS+gETgjN7op3etgbWtm4h7HsageLac/f8HISV1k9i
WNxBhK+Ku2i26Fu2r7jkbCONXDwTUvy8Q60JIIu8U13EWnw66yuWmxzzb3itWrLz
RO/lxkPnXRJo9fwf5Y2usuoz6GFAwi8zOEwz0OpJZEEfuaUwxd1hWwN8V6Qfl7n4
IW2BjdGD83Ho1+OXNAlWfLaAcJhWhgPN5K75LR8D+PU7ZqRCWLb7GyVstvbUWK4r
eNHtTAHK/8d0p0MYJUy2yOChE5eFo8c614p2H04bkEgVfBuN+4LMy2Paqun6Pb5n
zS1Q3zQoUntKByEg+Af28eWGUlix+rJU+kyU+AUKNo4TtLW9v5/eCwFVC6Lf0kbz
Z0lyd/LI8KJ0Pc+CHSUCU9z8IKVw2G3Yzmzrg+cDJmhHQhJypg7J6tPAdAlwZ2EU
XSR8S8dyJV/WyI2xD/Pch6wdaWpY46GFf/ysPZE7jA1ZvtplcTFJTdnZVzY6cyRA
PdOvHjpJWwuECEsxnBuYxtl8GWNIk1qagKEpZlBaIm1ypQwDwi0XgmO5Ri4SBJe5
lzlB4c0HEoyibxW1ZHsgK9HskYzCpJM/3v7+t9mqPYM0/p9aBjyrOLDi2VIeZXCE
yV1arD9/LZ52rQCVc5uNANTXKV1NRS/+MAXEVnhNMldd9O2j8DyMiO7wKfb3dhOU
lqTUszJ+PNSA5z1dOhbosTObZmMCgFQaIsXTPhwDCAgsXPXsHcb9+0QuxKZXYZ+N
Tc0ajVJNSRJYbCbfCNncvovySjZV903JQURDEf7U7HRLTun03gpO04/6tkdC0KF6
VuWmjnVXwK9vKvJ8D5r7GwdMfkLHl7iSnwUjwqcCQAqjuUVvpzmcUoRAMNQjZWYk
SfDRyHIvjJETpOPL8JQ75SRbbqQM8FiRF4Z7xnNJ9IeRFOm5lzodiCNLK3JLLCrD
z/c9lsC3ZFDexCfG4aM/6eKrpbpyvTJHkeqmcopu12fF9uMeZVLpK3zByr4Iv7rk
tGGLo6K39jHZNSY6nn4TEuecyFKQDmOUnnZAvsJ8rmh2kpDDFMj5JNZD6vc2vJ/I
HlVUZYn+ngOM28WKwx/pm1kcPEb48TDDDFc6EkEo8JwULmrFWF1nvZMiusWqxK78
1PyMhKAUfdpp13125K0dqlRLtwdv0VSf0OZfSXjKqH1EtR3JAPEleY/vuijJVKMZ
qtqCJ9UR9oQ1v7xWO0ltqaK/PLI/5GTgINxCSB8xRM9v3H2CCLV8Q4t5JtCcIb6B
FUC1iMsQs334VLMoKSp55JxnAo+OCiRgrSTqTYH+GI3fP7QnuaQ8ymrr6ip1ZyMR
iW0JYXiRbrQ6A0zKaFh0mKfJgyWwDUnPJztDAC4/8uWZM2yIgTBjWmQsqOXA+Kcw
8ge3vZPIC+eyZEZBqNGdZwIoPTzWanP78rPoYsSVfnPoT949MIAlWCKbkDETu6ID
n2BomuIPCeBmpfzYsF6b65/kZ1Sreeu0KJpzlC78uKycs8OgKmj9IMYe+ZLST2Oy
hq9iKSjsUvwEAlHpVHQ5xUa/z+bMTZZajENOaO1gZAq6MUi3M8cli6W5qr8NClcz
Cq5pc+pxjtyF8Vqti72rMThjS55cOJG9MdQ9iWDg4nK+oqnQ084aPSeLv3GUD46l
gQvPuN4RAgyK4EmXkmro4Kn9EIthXRk1TNbNDYVKuo2ECN1ipAi32Y8RklUbJnXy
Ma3JZm4lU0tx16PZkEHU2hekr2obZaKpY0yjY8H6akEJep5hyr7IufyLVcqK3WpJ
rWQ1cKEl+9xj/tOJ/Pe0Z/dkwz2GGKiPi54U/3yFNLhzKc3j2DCF/TfU49blcw2e
egQU/JuP6K12dC9yfwZLhNhr9KrC4wcsw2gm1zfsS2WDKEa9noOEUjm3NtV2VlJL
9Hu4Ssj6F4chzgotwuY5nBIKAMCV/z0uaKZQsyRAubS3rR4MMzehVYS1kuaVZuO4
Z/V+cXlMVy4i+5SRypvgycDhkR7slGSEWgV95nZLXpVJvdjl+5LAwX978Dhk5Bqu
fmfD+fW7hNZuNL1re5ayzhWvGURhEpqLPN2rb76WmxOLDsZX1KvxofxDQjULhLPx
sBbymxl66DIZB7kXzMpUUA2agb/qAlYtK6dGD2gT7gmizcxbRqYUF8KRWYNkVidI
0tQmS3IRWNhZChxos/nuNN6sDdOvWs3rXFHvdbj/wMz3d/Z6Z0Hi+Fq6TMXqU6yY
WLI+bObGRiyjtgUlpGHzWDZUp1TMp+9G2jlqc1occT93q4Myp4Ar9vW5qBUmoV9C
L+xWOtnGvc0AHvmxP0hqFYiRknvwZ1wwU2q7KXVQoTfUVrR21j+LmJ90Z58fExVv
4Er4BTjQnN/O1HMecIyymXVgOeZ14bzB8H9hKEs/L3ulu1Bvmh29E4xJN+74+rdz
VC2b/MFG5tMJgsNjYXjk0H1veZJ1xlM2CGUxvgLb5NFPR/ZjlwBWaTIqTBpc4GWz
jyKcvprjwCLCB2rvMlDq5JN1cpoR7NsMgJtJ+WsjUvXhMduysy0Ce6uIbdpF63is
z7QQD2DKKrKE1wuV5u2j+iLyueL5JTz8Jiafb+i0N3Z2nSmIfZ4Bn/HA7NgSpEJD
/j9DP+lDVeNXqIYti+wlah5gxs29yqBkg1BjxiMYTHlXCf4zEkXj/0MoJK9TamXs
BbRSpALKtTtRuyJ0ymIEptNR+nM7nzfkWhO0iofkd4VB4HZm3WUtcO+BxDtHU/BA
MibPGZBlpD7UJdHvwRgcjmLwL7JeDJz8uMA5xcQexC2jEIGoHlNu4pbJxR8ujFkK
YRRnNI08rsFPezZTjYTweaHJhEp1VH2NseTwbfJalRT2gort+M0XPFNKJHhFslb2
DiZs0K80tnpjRhfHTsAXYCzZqLTXb+zBmQE2Z6ro0w4fw7fzCMGP55VvUmxxPPK7
KJp2zDW7Izwd0DiUwMCpUtcTb/Sy8aq6210pUsmQ7WOs4kiMNNJBzX5nA9CHEWtB
jhxcK4x+hk/jjZZHTVbSxIJ6iRJYr1z4klvG8NYsfGGIlRnGSsriaTrGDsbCozAm
6cfc0lHalgwVNnTBaldjUTa80LjGkWk87p0/Qzg5togH0hWy+zbJWIlYk8z6Ef6f
PbWaSDCpcMU9bZCViHiJDQYkydnhdG+JeUfHPg0X6UKrR6fEql5H31ta6lJZuKfN
72wotR6mDps5FD/P3iF7+lnIvY+SUXsPJ71u9Db6lclqa7zcqtbN11ARmzAHUOjZ
zCQHzUpgv7KzdK7rUz7cUBCAPMt3g6sLhoqfyleh4lpWZ4f0B6JjCsg6LGyt8IeS
m+trO2aXK76fUrjjllV41v8LcuajOpfzAvDXKsMS4X9c1U7t32hyUfI7YmF79IQK
ThGrTrbArWcRDnDx0WoymyUkuK15HacGLwYEtYEMw6U80t4d/QNO2/axsVBvJj0t
airRzJMowcmRs7v/xuQ2ufWTzfrhVFdM/8VEiQSYBFZDGCiZyUb/u9mWtOIzvUFt
HR+NGG2T6h7zWqBJNjLErueBconLyKUygCc2munjlv1vCWqFPF3bTKJgNK65lKS/
dqvwF4N5sFDo6Xs8oawh7mOew0KQgVnbWyfNpPc5S42ygP3BKV+WHgiJ3Ln5HW+1
vRjjeNESS1vtOa2g5QBwIJAT8PZxM1bOcJAB70QNojqcenUAPiZPyMAJ4cGl9Vpz
Ar81Jq7MK0PO74bVG26ZIvr4GguQmPeeiZYwVbzLnukw+3siEVKeYK6ah0P/cSWu
OLSWgDqp1Ay83SYFcSELkBPcXFrczd5KsMsYodguogjdjfYymKfjxB5rYefYJO09
MbE+xz6+MELfLJiMakLGfmlwcm+6d5je3rxzKogrynOSYM1Jn70ZhCUvC+TXQPZL
SI9iUZ2C7jEhIPsoitR317mgETa56iL/aWmaWXA6uB+RQQNZEb0DFhZk80qkl3C5
Saf6JYtToKnhTb7DiO4h6I35RJyIBDYVTfL0C/i9N+JXLAH6QgVk9TMg4A+npTrS
bCc8uXflmSSFPxlnGcx/bIGGEaegKd5BPJH8abY9SHEVIrWCQj1yeEjwcvu44T4G
tHi1JMZlLhA7BYGktG8mAjygOdJlo1vtpBySR9RfVfHAN+jq4AnprF4FjQsmHL/H
O43dn59jsGqgTQtWRQqZkLzPKVNIZGmwQ9Rf0d2XiLA/HQYbbVLOMwgsjrmMBhla
vy1gFdiVbDmPw5u7Ghn3tgclZ5CY5lXv7kDqw05jzH3z+AR4dzdUUoe0r5w4mXJ+
FODDLFjOLSqzyOm7sRU2GVBygt/u3MxGjwTw0Wp5W7oUz+KuIzrgvLWNaVDkUFG6
QA1sIWOKClIjEnwPRF4KmdHEUHmXmw5yO7pqT20QhIk6Hjuwd/y/2/KhQBe+uVbj
Nm5y43AF+hJB1ap1FN+bhoaRfvwZ7NpWLmYMx6raqBlQnTBA2R9pXe3Gwx78zzbP
iNnshg2bfuj7tlhZTukW6GRy1qn/zYsTIrnjDwThCKw7KjqCaFYjYnnHgfvyEixN
7DoMB5bq6TGs7ESunilo/kmYUwXR/Rj2UL8W2Jd/8zIHoTUZJS1gSL50EpNJJUwD
rIW63G8EWgonEgl6CSXhM6753gSclEIvHCgAFRy+PVVpj9+EqECo+jekiQgpQidT
YNFfI3Wxvo2u5u1sgZJadlEGDjIAOvPNnaTsepdHJs+WaWQLu+FN6BcnJktXvZSY
qF7hR6mInuv+iU7+2lA9uW3tb7+IT2cyjgyP7f6vxUEUghfIHNCswY7S7lEpTRWp
C1tt6siwvHduLdBgP6Z0qVbaTNm8WsINVzuQ3CQcKnjK7kSMLRCsCi8In6mix6ei
JAHawSzuKCSdDGkRuW56OrxOU/OPtVrisYYkwlbDBGWWpPFvW4TBSkOAHAwMoxNo
YXJQxk/J87Wstcw8cVRxlvhQMrxjVY2n8/lc9WqkfD4nuK9SZf4GdMhB0KH5Q4dN
3L++3/kqDTuGxIWM8hudINNRBjxLSY8XGrYcJ26NtG92avFQIFLjPSwB3+D5FUEx
byLckMlVaKtKtvgwxGgl6iEtq8xCRwtcuyYCuyUPQjY96kncKi5b/1z+Mh6zejpC
ZQexbYiQr1larovNfPHcX8jSgrod1zalacyWRcrGqFkncQxyvS6EDVfClxVIQ17n
BsmeJClPwaa4lP2jDN0zPXxD7LUlYNXFyrwhdwwR+j3gUUP/D1qiSltxWuHQG3Yo
jZ1e0NtAf+BcMaP8+mx3exXL8z2mml1wKPwmIVLreHHipUIdogYBwIBKfStNooTo
mLGmOLaXf2sQHr6xq3bblhpo7cjggRKnutGwpkH9AN1RBsD66XwoOWfnmkanH50z
f6NsaTz9Z4Y8ZS4vdzlnlDWxtXBKYAGCJncKB+A75alFIfr6bEvEi1CJ2+ptGaAV
Uf07ol1QUCu9H0y/0R8QGrbeF581k9J8t9RQGnUcQ8BFuJ6tDG8hDWbjXIu/qldY
tF4IbTopdpbBDHO/bpE9TRew947eIU+kZ0br3hcDCG2VLeUr/DepjC4YUQAcWd//
O9iFB5vPFjPtw66VfHoV3dA21hF4lXQQVH5pj9G3PssA7ZQ7XoTOtkexqK0GlTeu
FM1pHvp7L8Rzc5ljqFO8VcVEmRPaoZU5u2mOx2v9nStrgWFa27YBaNX+XoLeoHKv
rTMz1aVcSA4ir1AHQU7n3dlWZYTczL3phXLeOrKKYZS8wffOsAx2J0XtL0NlJc0R
84n4nlTpg11ghWiHOm8SFF1mEfkISXYjz5K9TfjobjSIs+gXtSXiqf3pZANha8jK
Z20H4QRvUvJfZ+1tmuvjTrCaYgz7YpachIScPSscH+ClboRfGazXJroCiMyDpCsu
FpsjMit2jMpls+VOk+VEPG/ijsjwGThasrvhLUQ4ywdouBfmtoPQFx2FYFsJ1RkY
QIR76K7q7lom8I1WVM4QBq8t3saY92pxOQp+t92J4HGxNq8n5WDlz7cebHKeU8T6
FOAoOIkDlA0Yk6JxTjZZGbVRUp55AFOeAV73ibSzvtj4pUZpYHDgIUHdiJF8RcS1
AugO4fv+8AKQfMWOTBJFp29S2Iv35o+xdotA9GZnkNFaf+38IsaO99n9wVHVzbO2
vBlrk4fDnl53CN+y6GLSfQbb9cbN1ayKOUHkpMpDwdp6HrdpNd+AOaZuSPvahx7m
T1hXrVPkjauZh6YN5F+UwVXaVPsn/F4h0AQRC2kUqfH9zp4/JAX5gVPMaeTpnrDa
HPE1hpvhVttdx5A8p8wtXv8PZKxFdpMkDMLw59fqm+c38Zhzhb79JF7MaBZR3JI9
BoB7GcBtEOHGPaFZXoHc+wODM0JoPlhYkeFfEqmOTP76XYPCdnHASbdukndCVV2e
MR/QU3OZQFv9CvPRgjQdrRg6lMDprSPMU7L9cq567VfB+Pas/N7CnVtd7E17EAbP
ntGHCAy3nViC/2Sdfe65uBuKb4ZYhFS07yXT698ZOAivtvF5K/VpLnke6hU4j35j
lh31rp/9NaSIT4RVYFe44wgefz6ux8JmxwE5hxwRNyYCpP8JQDAV7zvprbvTbNSm
6/I11cAhlA2ei98D1XtNBOh2BSKdhpt7Bgv2yK/qBLAQwNCEFpxSDc37NYOwLNNq
yVyr+CkM1+9ydfuxi6wcQO5n43aaV93+ZQZWzu6SFRCa0x96HjXQrxtqqnlH0iOn
XkGgphL2A5Bs4Gvcx5TJsfxm56JL5sxf54C1+csueiJWTul08fJ3xY+s+hPHTwpT
fehyX0KhI5jQuWxMOh3k/BDHHXuxSycLAMGKry/uvPEV55D5bBmaPBjSdUl0PZQv
jCgYwXcREEZ6v1nHsMuCfT9hFkx9JUa/O+xA0hYod6WCafSzV85PPGhJ76WdmE6H
l8AXypTrkFcapcboGbqOiP3jK5t0WchgWKQOSKJ+pHurpXuBr38V/gEgvgZh4JRU
IJqaQoOb/bxjyQ7yG4U9Lp0bD5mKQONkLZa9IHXzdk2P9QIWc/jnrkNAw/oBbkNX
LRTKCM2t9jMjGmUu1v/JiIBYWH+phcvgobkonxax7fMRLFL2SkigN/UacI4Upvrs
KY8B7eYF7mrI/Q+B0K1Ay2riJLgA81HygY3uBAiedHIfSa4K8SKD3xwaHlpWStsa
o3qxne1MpVHOecVrfCHlD+ilyYq8Y1du/HOn6NWT5Zo7b8GDpyQhGi58XuOIIUbi
0rFnbTmgW6lEk876zWP3hS5YvousY9xVWZLJZhVVUoZijJniq4i/JqN8sGefHLbl
Fc0pfZY6cWAhPkL9qv8DCa91pCyLHaqgx9EKtsvs3sRpesY4eZeUFuwVn6OoKaZX
tm2aQjJbs1nsePXklJjpMy6gDzTeFY9odS80rhhO15AiUlwldgbn9SdzwUf1mn06
ft3AcxWHqWzNHKLTBgxVJpp4sWYD/4Iz6LJNZIj4RS3JZ8a0GszxOaT81/SjQP4S
378Nz9KgXgQpP0uTouJ/CIGH4ds8x7GWEfJVjoeVsqag4lVKQIhp9lL9cKBq1tpq
u0YtHhYp2OO3j37q8CrplOmgGgMNseJI8USQEaUQo3oBt9WJLsS1r2rbSUmHN3fj
N4DN/C185UIEDmu6ZiA2cZoq+PQH028XRurV45c9nSFBD+15X+pQJy/GybbwN3RU
/9zztU6bHfkx8vp34t9NRQGKY4hp5xQeMugadQFUXJCHAzsDVoluk5AbV+BZsEUx
7d20g/KnGkAkpr77I/8/wyZBV4vt9hv9eJwcxXjo/VpP746bX5HqiogjQJoAV42D
5XHbt3AIFp1WPe4eZU0V0BferbgsF4e/zk3nTSHonlLyqV6mqc5v9+rDX9EUo/Wv
0H8u55EICiQ9HM7YE/Sm9RLZCLQDjOqmQhO3mlwNUQQs99MuHD/6TEOKo+okbM2K
ogODkaAzX4myUTr1q4di4tnlDy9wWnAz3vk8L0XX1GlSKNhAF38CDk+T9O17dOls
4B1T1hNqokzxibkrGBhzAtfhdtE2tK/QCQiH1jWYcKQ3BLKsBStb+J0MpG9fD7iS
E+HOtg4+FvMNS+hNm/668QoORhwDkvHHAnASpbBLprA0brIc/UietI8t2YstsdGg
DHlvwHxtS9pUwc7H/w20NO3bKIScTZsr/tKVq6jybiM47aMZYGEsil4OU0xigcWF
HHbx72DI+aQ0kh4G1rDEHfJPpV6fRy7p2c9aFag+oAysOR3BopVvz3vrg7Bb6WeA
K+ID4tPmKjgq07Ae00wsATrAqdv5LXx/LkOJNbsUtB8OL+bdfZIBytacZ3iqm/Dr
h+N1qfUFB3WecsGRibIW5qDPeSmIkPctTZSVSxKYpP42OozEnMPcDzJGorLOay/b
9CexLvWkK5RZTxjSIbeJDhrkfRUpoS47yEuDJhn4cU5DZAstIAOhsi1uejLjeL8V
e6BdbqHxtJ7VdjnecLjW1xMwaZ6Q+kM1Or4OqpVL9rcgGgYbTh2uMZr5TeSbAD+Z
90y40mqNcPjuZ3qTuebdK9RbEj/wBlhp5mTvJjucpo4RM12QkqlLzbhgywRo4tqk
0jTvvbCxenHHBxll/TzcR/ZJqNVN5ZZQMzgwyNuLxhXwqAYa3gcexHg4xKJdDX/+
ctNzf9kA3L5VUh2cZIq55uKMpX5kEGlkWd1ybdr/dSnpLzyj6EPY+QEu26POG1os
iU9913DcLNaGhHH2bbP8UFGZJxyW5JFvuRNHzzMTuKpNIumm1/uwqwh1ZRUkgvUD
+kLxTjB1DB2CQwHHFqbAdfXWEE3vLphegJV6OOhYpNyMnsSW9po1Q5KRj0wtuPbV
DXCQkAlV3Qb9XL3CTEhLACVOsgxjHI9C8y6dPC7ImbqZdYx+EyThbngDqcLgiR7i
Op2oOk7tOUjAgtcHifc+SAZRBky4Udzy5BmL3ESflj1IGeV9h8hlswi0TXwAiKli
1kpTH3x1xg8nbPWkjeEABcNJWwd72lovuy26238b5vmKrgbJXdoCIhNWY2dMXUkN
todDm3dJ9WjeZjO0mtWg13Lvs14lLeEWWY0ZHc1BJ3zaruq6IgzLmC30DbjNManZ
AP/sQzxJh7iBL9Ldz0trCwL6RlgUtlldyIxm9wkXlopH/P55+lo3rh6YsQ/3NuwO
1Mf/C0Ma9FcHiTKf82mNBYe3s67fOoi05JvXUYIfXNB09/lKYsWyLzE/rbwAUlyP
NElpKfryRsBplSF9qH+8Zc/H6vbi+HWawyPvzYNSvuppaHHRhg74Z8iYWYMKgeZD
pQmtx3A/upGSs3LqU/V5o0/T1X259DqtqTib9XNyrYICLDp8V44ucUWiGOZCLoC7
vmgeTty+Z82mvsw/FRvmjP9sFDm7A8bkB0Mbxmt97kVYi/9IGKVsVogozVSyzgNk
OaRNLUtgZVfonv9/Fwtq/67UsvrNeLygWmllPhoTJi1fmn8a4BEtremvC7ucdpnP
d+MImBCfLLFV4BkGV7aKKRwABbDbC+Z4OXkcyUdMcH8ahqsgh8iX9FOlCWu6yXqK
5hTTStAoThWyeqSPs9YAkGkQvr0Lu7hgAivsEBnHZm2urbgau/Sm0InjawnH6Dxl
PE25UYU4fm6TMPOz1nKQiCnHB9LtOhr9SptqbaxcCDyg4QQaSAf54YpQ57U5uz7s
ejeEhDir1KmWuWAqfKN3gWW2EFwfZyt0teiAOHV8+5qjrt/qbHHhGES9bZRK/V+s
HAUvUkv3v+H4mZQ5tVTb6bay8uPB/a7GMgtFOuhhKjdfZtSOSX+RRCF7XD6uzBGH
v1x8Phb97byyJa6+6XpAABrQROF5GcMcRcJwjy466JSYWbnxps1mrLET82rkAusx
tuxorb7BBv/aMayp/lrANLBC9AGLtLgPRNOIGQXfDmzdPOc06iS8/JBi0tJuMDQB
0szHSBMyCSqziq/Qh5fofjujZmS7x4l4wmFaEbH3SMpcT+MLtkgWPGxvepko/Q/v
Aa81Aynfn9POb3dLeBrUNHGOLHMeNObcRCzbZ34mmteeBeH9SrVBFidh3AsRYxJV
baa0mpUM+2LWzrHM1/HKwwbRPcfS8sUVrdSMA1IjyoSrJLKVlZGtkSCx4h/9e7ft
jU8EaUFXriEkeNBKQdrH5udE7/WOcN4Tz+bSItc0m42PqM2CWYmjNJQVsqK2fh/s
bNWDUyPduByPglmhd8Rk+GyMj8bSA5KQRiGGvbflQIt1AVzVv1ax5L7qwTsN2WsA
O9SMYD1Poz6YVm11BhnPdvwguS2N/UmoddfwPeoq9uTPMXnctCirnl8+7F27AWic
JQT31CL5I/YdxdfUYrftWajW4lwzoyASivNzwb9M+fWT6M6N4dmPH4fggYxT/GnK
2aN4fhDR8s9+JYEf02GNqkQqnUvRKMSEY//InUro+FxU2aa7/PbDR2ZC1goDYSBA
3zri4neOl47vtPIYAOUH67hliYwQRsaoSgegrcuC3RipAmc3Ebum0fL++GF3ctVL
3l8U0DnVvlgGGBkAOlbeiTxnJ+voYzGYtiO12hqkarm5Gp9foTJhadaEHlycHkJA
T9DIjielibH8mmMtrsXneDr7H9ZHlDVmw+FhJT/E50oNykioIFR3RFe3zo5dIcEn
2DCUbCZMjqAbwneW1z+eaLm2tZBqTXQGux+08DhjSY9wm7wJy5ttde8+GSxSeceu
h+qkpiZurbzF/pL5aovv5ZAkCR70B2iukaqI+SJUnLzq5Xs3WlKxLkDNC1g2voU+
rFqgyXcMEgkmDjRf+SB5DdrpLojqBL4w3f5q4iNdg/roEYD//fnFE8/DmywwXYAQ
cFUBZUJJ0IFjvUw/rOP7nPyDxahvyoDANkuausQ0v+23g2MzYIPR5OpqsDPIx4Oe
kJaKCyvVHSdrMqBOu7yciD2f0Rfpbbinf/6ToEuoFcIoMfJu7CGf3BX9cEu9Z1bg
QLjI244Fbx994jzsCP0wNMNltqra3izOJHsKuS0NVgSM939fZnogb9/zfr2+myap
AMchK/zxSnp+7YbRfaIFj8rK6SH99wTIDUY4Qz03dOwrMdgf2H8NqGixD2RU7Bw9
LSanR+LBfWBXiBeEXQpifYET4wSTV69HZmBW2VrD8Wn72XK+YeubCheYVVqff5bl
BOwOf4Jst82/Km1SRI2kShWeyeHZCD/UY3vaSMBsPPwOrtHbhSIavB47CJUk0cba
fFBqNml1jrq7OdJenhhvEX0SA38SOd4ap9Rk5vyUFVAMQ5VefA+LhORIBwKW66Yj
37agiU1YhQyO0gAZIQT7uQp48h+m7q2iQvwTWv3S6IFLD/RYJkwgXeAqxbAfgZM0
VrkMJ1+a4Pju8mbII/rL7kTdFkbuzLd3vf//uDiEqkv0j7yAgL7mofqyr3HtxHBk
nzX9sN6385HT1kvaK5QwqBVbgK0ZmBI6FdmiRya0VLWFW4dg63Jwt+G3uoONzL8g
KpwQtdC2mp0c/cQGPzbr9H7avUdHjjhivicBKV+gS6XP7QqxAKaKW/A5n0cf4KH9
CHgqUQASAP35hVdeayopFnt5xv0LJO/fh8bYjKUh3fMwjLcAQYzQkxB3pV6r4tDt
d7H6Wgn1TDl1Aqjzs1D79co9Y0b4EEiy7u7X6UfvlnTYSEnAYrLMoK+xMFtJ49AD
vnu4eqSSWD2ENUgnk5zBLuQU1kdM+l9a9K/+v1V1AbMaWvV+PquXCyF/+A7YSZK3
AM2T3FVo/M9gdKruVddhJFR+CbzBOFYfFwEq11W/2544+sR5KUyo/M9IIWEcPSD5
mmXOzshQbpiYEYuBC/zYT2a7deG/bYhaW39HeS5r4YgXg1NqXlW1gDhLJxntYNyu
Sbh/R8YzI4fFBeWwKBCwN2gbPS0/oQSoF3TjSG5NTBUtkelFK5pcZ8xx9EN55YAa
8WpxBs1mImR6Nuqr1mLQwXMOqC/ZHgoVy7uW/7OLsdIdG/t39g0Pout7zMM/bNiC
JFp2eNN8Fp7nxV+0LHn0ND87bZlPwHGVae1K74QG5UaAHCTzRN4e4Z9fg5btfV3j
N0u//FwY2P5ISEjJOQai0+AJV9PRrpN79J8c+q17ggUAUlXyzPBVxGT6fZtWCqzn
ZuwC2kITF9nENEMW1EdcDDOzYAKoqv6YpcWGGtPW+bwjexD2n/GD8s0XV8eZKIVa
7UzTecf1DrHhR890l3tPWz4eV8+p83KmBZdiW7tGFKtDhRIInGnW5nF6ttmJb02x
w0xnHwe4u01KcrR3CHnJpJEDvgeAOVP81o3hR4xqpu+8OrQ12P9wB2P3Qi6s5lxD
3wKUUg4wD10lftstp82+nllnKs3r+1UwUFtRkKQnWMSNr7HIwg0EjufeJVeOkLsf
oA/ij47+sNH6CxUAQRALKyVTMvmrx98sPl0/uKROe16+tXJweB++qJQRR79xdlDS
Er7DjbcqcQslEatTiUuBLOsXHZySW3MB9wwm3K9CP9r2xHZEChvq7Bw0Ww7uzlUP
qTlpEdiAAy5zlFnzmzc9QBKX0Dmtv/U3PPSNGrlPLPQkGjspd2RTSxGkQVcWngRP
IcI+nPBAEY5mfoedPIJOkwgCUUlNUjW/Xe1pGABU8hI878n307ORxDvzfHnuX4KX
32RWfcE0Sb+odqzkmmqCZCAAd65tOA+RROAGMbluk3wRp1QOm4jbs4f9wZ0ehuv8
JmfC3mpCHvYDfxtcB6uD5siDL5JyijrcRsWPTydet5i/mlN3YfgJcfL8r4pP4HLk
p9vyK38zTAGpLBmp4nDw+YFANvXDEk1q1ttoJZoRdHr2kwvbjdoh8SU2VP61rgao
je6sp4CqtRUQoCy1r/hz7lxLwAfeywdQuBp9LwNuze0TietH7DoK6bRh6Xm/UAe3
MzXAmdB62H2uJxKnWz0g6uuiIcoPs7MhIz7ruxSj0f+zQ/gyKB7XgLNVdsW6LLwr
E+HnrblgJGQtBoXOXPLBCgGYOeubpVLUFEzsZQRW4bgd5j+Rl2AKeJeC0PnG999Q
oP18mbYq9nEVXmHT4uX4RROukHyTE4B44qVWm6M1Slts/Z2aW0cvmFOIr4m5mUvD
z+LP/2KArq5CoTq+dRZvHIoBRtV3hM5GKdinnjxa9Xb5N5BY8PkZyAflePfr6QGU
ERxa/E8yT4+aSIYW2NayHiJ/qEBA36xKqoX8v2a5WdTpx+kXyVFJyk92QIN2Nazz
dt3XepE8MtWAKVxYgcPpen5MjFNWx8uwuUQz53EjsPZduwbFJHmtnA708iTnFcWB
swKAre0e3cE4zZ5oMk9haNF7kgL2washJdYnwcFXIwol79BIumNU0eTRxr14frQG
pIgVDzqCCSzP6OYmzMBL0FUaCUiPdcA+z8v++OPnq3umozQ5EFEK6UfKdhzF5Df8
oVTaJUt3nrIA5zSQlykFdh/DExqX4hWJyfSj/A12pEWITFzqOAfR8CfaD4Pr+DT5
ChqDgZQFYE3qwHfNxLhu/vtX7VL5knQO5Dq74SJqrdf/BSB9rPMlLOtCcQg22fW+
LAfupwx/tzHzPCHp2tWoVLdSFp+NWpYmGDmpeyuJYC7NDXnb0olSUF4qql2pNSF6
TTZSU6Lq9Ocaui6ImAUWKN4/BDtHEHzdfYE3MUATHrGE+hcMs/Ghc1jV1hTvGPHD
lOIlFdg9vUfMBw70I+eyilh0C5JtCI7RNK3aAPPRO/PZb5RaUqSaQgmgPkZcMJTc
b/k5XmRaURRl4H+81h9Z579TsZ+aLs1TF8v6jbth7uszh+zyaNiJDnrZcbC/xGgE
SMTyCN+NCjxXf9PMmsyMTLC2Q5woi/Q0eZaJLeNkpExtaJkH7nEKbPf/SdeAdbSU
CnUrjZPcWajr466NBAyG9lL1PXML8NlivOlqcVKIQ9RPiGDokAhTQoqrSZo2wdiJ
PSsZzJ4ckjmWR7aH9NC28z4rhQpf7mZIa/ZdKKy8Ae3KmyQglTja4E3EqmOV7nOo
7NA4zJtRtKCrOR9VavcSgwIYS0oK9zKzDVR94aEcwmij5Qwe2RzfChzxncMjAlcP
vFx4nKfWXtkJpVt0XBJMBrF+0USJxLS9hqtjvfUOeLTBrh5RmuU5BfjAXcg7Bujf
v4ZjWo+NbUhXIDlBkQFcoR372XdlztRCS+AwfCn64Ifo6x2oSFvL7OTCW5vvGoor
rtkwuxB4mGBcvmeUDBAamiz9AM9aHO9qei+PhyvTlcW3BK/iYcNIzdnHHWgrl5UP
Swamg+9rnCD/V5mDQDPAJtnhElEHvyXzttMFQY+ljNuOnBcCcpuWjMmyPgPOJXUy
2OhdVo/088BP5Ws+Vl/I5rdQguTwuT1qfo+gRozWF0aXe3uEciHxwnZP2MBR3CPy
b3u2P3PrSYy4upP6MyRLtA4wjgfFQ3dej2RT3loYJ3yNatrbd0wP6s393E/hqX94
+wkipWtxgJQCNHpbpFdV43Lp0Ep4UQdknIAa7uPrSRJWjtOZ+q+e7HGAG5MQv5E1
TdhLDnH12TQvz6d5YikqoA8Xc2gmXC/bZ55KAQJrCtet2W2mNPV8GOSr9eWT05vJ
SmHw81CuvoqkmdwPREd7UcBj6EKXAYf80zmA7hn2/C6FNfhicjKNi8yq9Lm5Eue0
46aicRcxnrYSqRvheptwizkqEt7+C0TIMCit846lsUNCdojRwwrbWXaEXkyqXtaH
hMQeXL7ERzNTB8UVp/arA/M6FgcqEE50X0u3GMSZZIqIeJB6kLl5Cof4ZWxcKJ4e
BmePd2dAj/gmO8yN4KQ9aBsXLLUpasW4oOY0nNiLOR0t3kaJakLV33dpwf2D0a8e
pAei1a3eKrLIrjyzvG5riOTeiMPxyVu0xnLBZ/Ig27n9Z/T3u5BtniBziquc8yiw
SPJQUDS8w85CkSTCfov75gfyhx89JSdW3HCJHJpF7jEXVzvJQw/hmCbHmrAZfllu
Jso9kH1nIkw5CHcxtPfNkCSQJRtdRpmCHD3pEV2NhXyjEPgG/PZ+soxkZuDDdpIj
wwywqD3dsxWx6EHrFosjjKg0HTsmErh3n1AcyOCrbjwGC+yolLZ16F+3AMoETCc1
IUBJfXQMTl+PRdsMhg71hoBULJSKxyqS+HB6ttojVed8o4QyxcnuWb7fPLSyPqBH
EjLBTVbz2BhXlH8joF79pxB006WQPmGr/WD3R7nomODlu/HXlXbNozGVH1gIiCWb
Px4IynjJ/q7QPdiknDPkjZ8t5uBPx/HprXXyOoQpsBM21CPCVDyoLHB0Dj14w8Qw
nrH01xzCI6mqHr56DBhHIio2/DxZGlkpCeh/LETi31ubWsREawhe5m/wOKFiPjAR
/A39O7SS59hszqwIrSNlPPc+eJzvhCEKUZ+vTBSRypg7uVmOV0UlAO5w+ynITqgV
CEfuNDExcJhUOyaDtrJp+nIGBThIkWCnCLL5vgXUJzOixWaYpRSKOIKb1s1Rcjzi
aUst24fYP4v0SZT6iiasjg2sk27RLlV1y6+JiZ9JsfsEW79U/z9l30aczHx/s0l9
zmQSPVtR/cTz3wKXxC6rcGZ8cPYG9Sahg+Hp1WhHtAzdhYydjEfwpyIQmoBHKkti
nBNoGM6y1HsiCVhMFP5x/MlvJsuJ+J03UCHNQ2jENyOyGVmnUjIe9GqVxPdlrjb6
JI7VGJGw26S472TZViUezlrNDTl+eQ+9MFB/klRNzTirvraPtdLYI2cJsA6YR7W5
jQMaEAW4NgGpYMsGEKeb6LCHE1Lyiq7UJNQXelP3GvFFhBVxU3uQCo0MqfX3o5fS
udkqgqQeMIWrD+D05r8HHOaxTtrKi3l/hEFDKOpf8ZHa9Sq0KPlEfOJMSwq9ZyLw
RH8vgJliePOlMluo7MNBIbs2Owjn8EwsAutXceWBJOuRiEvTmj2JKYbKkQUUSLDg
szjic+MBM9M5X3jkTaKmzThvlV6dSE9MdEzyojsAlmPBgOPA+rdt9XkIcFHTJTJm
STo83pXaZIS7aFmayDqah5t2COnDF62N1JSPHyaFVQ5fFJYFhH5N5NflBV4h/LGa
u1JR1qvLw9tQUt60GjgblfN0hKPuZq65kfM0MlD7AQqP5BohogVqiRG5CQLpEqOc
6mzsME6YmF4g3o9edz89eQmyknIqKLiYoqUXrgyo3koXVNHjN+bdctD9L/DMd1b0
0OihcAcoM/10v/3WUMTUE0NNSvEyrUtsE9cNK5jY3ZUyPFbrULf40pT3fQ+nQNj/
o3YeoyFrYQCusUZZCaX8TzHngD7LoKVX5OwqBhwZABxyLva42jcR+HJc/7QOeuaF
KhXCjQ5gwR6Kqnc6WcXkAc7trheo8PtnPiQhxaEuvuvnONorgqMY+0jxuclQKBQn
a2ftLOy/mpXHIsjODK2RV1hWH7wTUipQY6bWQAtWFMVdcD2cN4HWrcqwOfMuMmkj
JaEEKGGqj1/rfz/t7ZizZdUmWsRS4+YtV9dg62xhD7RObO48JdNaJ2lAZi6V9Etx
HJ4lCEc4XgoIfabCLnW2eLBgvQJjIYn0cuzBMyWlAZlnvKKxFas6MtF4s8uSB+rf
NKukKnjHq24+1uPwhnJl5hFslmleWHSJBTOj66Eq2wPwcyzheND73zwBaTJJyVfb
1zH/NSnXrBa83n2xkjkCaA55tJCJmCjYXvJuSLVfmEeewZ4X+R3RBHRFGCNXllYd
JJwdPw569lMLUNb0UkMXUG+/1vP+d3xNr1COuMIIeD4M4EoIImogay+gQLWf0Yfi
3UG2QiS7w6XAEpolnH+WPdWr/7MNK6v7Cq4qUZNKGEUt6eUU0NByznNBsx316dh9
2MAIoQ7tLp1egaGUviPZBPM8jSzt4vqv6X1v/Fsvawe0vPcW/ojWu5StlGWMnLP0
WdwjRGLNSClTkjJy/6jICccfPUiTODVFLNrbc8RkwhCe1Q09wOM42GusWa7zesOL
Nx6lS0u0Kj54uC93LFVDgvdrihCOUSNr2V2Rdl0dvLANy5dXkAM/xZdZNuJW+cfJ
K01Vr0VTq7+Wcc9bE1DMmtudJfIsREjPvV7Zw7wGjZ4U6nasjE/mnKf+zLEQNeDI
ItMaJY1e5thOGXFBW1ftHnc0LlkowiVJ428l0LOpUsw2jugLjApbzIMQR+eqNhW5
/A1XNHVUvJaPZE4WFoCQUtvIykjq9+TKr8hMvMo0TzXr5/8jxYgm+H6lZXeBR+nP
xDfR1AVKh2n4mBpFkgz+WjFThqLAdQ3tVhPG2qx1BtkqGvBsrMLF6Dzov8gYOAHh
pXEeXj+b/EudBhrwvWwikasoPNofAFX2yT/X5ua0akLh2x2VaMLiAaYtd+0KtMcN
v2m7kLkMnRuzY8s3Uc3K1zSDskMSxTSErbJ2c2hh9qf3dP9wX+Xe85TTMkJQMCjA
Dxp2BN00xavV0e/TdqisWOW5QfkFpJzLknaEDZtFZ8NEuhIc5C0s88anaUvs49FM
vy1DwBsXQwd6dPR6eedAjg3y9LFrFh57lydI1cmxDogAb3ALW54HaoM4Rb3dliU/
4O4t8u2RODGHzA2sgCU993IuL8qRE3bGFqxWer5HhNTgOzXoJ6zpCopx/WDll0m7
M1QmJ2Wmj/BRDToG0OlFNbqxo8/Jxv7gOFDgxtnFtZRbEZc0ZeeCI4pwO5eet+Nv
1+L4CVW8HcOj9AWcD8whU5+/NjL6Dw88G5OYNAD7U6AxFpY79uAYTKQPNTb05rig
XXvjLuqxucsiszBLke17JnmuQ8bRCQioqqkLS3v4RPba3gK3XLUA6DS6j/Axuj8i
eRMLVuboLrMqk4AKgOU4gxuwVyyR/ZrGXGH942ktVFRqOE8MiFYtwN8QvZJfH3Ka
dzliJQFImFvKTtikfOsoiQ+PIUY7Xy/EWGbqeR2sXbRM1gOtZg5ut6c+r501cWC2
bsocElRYb/15h8wkec8aOP1PgNuv8wQHBqj7UxK1a4PsAhlDjuTp2+k0ZW+UyRrX
vqwJjTGCTLS41zMyixMFR6EU2+usWeR2rahsY+1YtySN/YmvjbAOf6E8491EpmeA
/PDSsxGW83DjATmprmB4M4gIrdoo3+PulUig7b0x0yJveb10BhGC6MDyKeyLhNDU
xC4t9RUvwTtPhvyxw1slBYAFUy5VNVjFVbJ9POg30RPy+xsZiyUVYNlr5NHx70SA
512V7BZ3xBIL43z1pbnqdX+SqFzpOpq1swDdIUx/EsDw9PTiwWYGFO7vwUaLsmEO
PfV4bsH4BiaOYGOaqqyeO1K/U9bGxZZ+eS+qzCVDDPBetWMHkaQcWjqNXcsUsZc1
+5Q15oPGiUtvG04+O80FONOfP1lJ8YSbqFx+5nkdxS/BZOT0AbqjfsNiW+wScw9h
7ClrpBynhHwPTtOmNfbTJSown2o2wPxJRzqtaAcWxY9YQYIuEL7Nlb8ujri24y1b
Gq44dsuCjS6JikcUyiJMG8dwsvGLKYpCyt1vVJrHIGJm2E0aL6R60/62h1hlVVaR
uaoCtnV5Vr9XpxXlx7CxC/Fs629T8UGGiXahPwBxdDKe+Fd7hj/fHkrPS7nWqxxW
64mp9WTJFdH7jzjyhcX/x5GCzGORC22zBOsmJ1OiHZ7oK/xjSbQyQEsKGKvNZw5B
kpb8lHPA3IbIOI76tv6a38yqd50ZnIHCGms6zGV5AEwjDBWwb/rKwnvJJ8fIsLTf
kqDWWS32Y/2WQH1CrZCKiDqGXpNNa4leae7apL9VSMFIu+p465m5vFfwnlsmTuaq
6LnXAVPvjljqVlPA1viEVS1DJeRBUDDdaAu4Yu3Qp+rkVyjDHsGpYWSbNgUkvVzd
R1JT/jcdL1nNVC44wV4d3nx1YWgGGdNhDhL6p6VP7qDgyMmLspjHxOokI0ppVfaX
nSyWbUgn7VVLhCwRvGWKAmrhxK9kdBreNO6xykq0kWsGjwA6zvmt06zQhmzJFIKp
r5z0oVDATkjvTMEyGrv/AwKxT1E4JQ2cSoYYQT4UYqqTPGy30xhQF+83MYHSp5Ov
F6jZlgzOLae0OMGp/utsQt411toPuN9hgmWaTHxiN+JH3wM7FbgP5slcUwU9KnXr
FaySVBhpsxIV1woAow0dWWLmhyLmu7fpfql/UPvgOOST7yi6ScwDktSulSHdhLzY
ZgwQ8ADvaTxGVc9WK3mH/fnUcUVKlPUVQVn6mYV+hlN30XYUN8PUmWmxOG3t9lsd
Z+U6DsqUDG/YNC6oDWLXIHsqxvnQ8gUmvXJ1onZVCFLshjlwrrv83LhZSITdsocK
76Y93h8chh6UZsRDMRTrNd2qmZpEwuZUpCNHcYtrIRskxWb3Fp74RLnabsqtFpP0
2i2pvInGWSH+ugv4W9SlCbAYSmM6soPxc1wbdUPCaXlZEpDQNto86FKt7M7Uvi6F
MpTQAwIrQrmw8BErxOy4cPUMoLMPO7GfMkqGaB3NSY2hvSeUTcnzDm7k2o0Dufkg
itSA5Am5BNiPeRGkuRHt+cgQMDvzPu2JQEcLzdkpYTYrWD//2ABQ9as4se3OSgGe
4I2GiIzdGdr8sE3nKp3OcmyleP/+NatpuQxbmfptlSz5SMDLcpkTg+sWnsrRtjiO
cKFKjyaO1Djerl7LalffzUTV9uTnUoz5HcdH1t+agG2efLhhljZyamYvmFNoPpN6
jPjP9srEjZT/ms7KKxsigUmwC8XUBfFGkG50YDQyc4cR82ZWZ5Dl2iv16Q8m7h6i
83jFYg/j0w/H/Bt/4hP7mTDnutRwCoN83jmZpPQdwGeFUv9e8SnhAsXdSyiqZNmF
1TOufqVxbmpIdSSQ7kadrfi0/fYUk5yGAsXbmx4j7c4yySrfPKkEGKzlqwAtMmDo
7dAabUUt5kDwwUbRV4OUZzLrf9/QcfTZ+rAG4q9mmKWSB4g7hacJDE87kLta70wP
bCkhrYIYHyIBezhbGEg0H56HTFN57JuJKE/tn4sJXcTlAQzYTaFT9W3zLEUcHeoa
G4A+ddFs1BJ8LT6xJkMMuGr6TjIfN6Xc+uuUc/rFRJ1hN8GbikPbgQ47CGVMJ6Jv
6U8f5b6eejhSVWEXxNlgW67dmmzOPKX/ad8npN5wBH4Je8fQmZtI1CcSzVjbRU6C
dg3D8tZM8II+1OnZH/Ym19SH3JO190k+PdX3Fbm2BtUExNvO5+L9+ldCWCxhUe2n
OnMf5UfQFUEFHMZkiIw2EqoNG4sZIeNUSORHpT71refZuPT6D3LRpgV6LQlti5wy
O0GGxiz/nBxHAj0dLgmKhu4Rmk1xkM3hX96kjMZz9GjiKR+Lxl9U589A8+bv9BLD
EdUmMysMadlW7P5kADc9BxsaZ0WJFp4zN0N3oMr92BtL0I9KtKjTScPCr1O8toQz
ufqjcYLAvjXxew5WNPp86wXlsQrUe8wMvpO/dQtKq/+Y6Lh02HUeBPyQZ6TJrHAp
8lfqg1DCITpRUxbuJ+rAx99kTjdk4nPE99ovgiiiWnJ7LIJ/W+McEIxNXWWdg2Wy
Jq0TWN7TjqoYjjnQXxHPzs9QNV4nCWFm6lbsGlI7YUCCoQ+zYD5wuq/z9hcsoZ5o
SiTRzOUC3LfEo1OsuUncMlpsezidZ9V872BDLiw9RwQeLcqJEOYJ6a7zRfZYX+v/
ubko/YMVzO0LpRso6aSsLs1hWxFbB20bsatlyTwBN0iB+AChZJBOgpza5gQaVmai
2KCeSB0dHE0ecj0drLJPqgbLwaXa49IVLpu/zUT+m9HPFBEguTiI4xLGc0YyWGD4
8eOJ9b4vGbi1x8Cv4jHlGPKHsimpDIAxBxXrCewGELRwFmvXSIJW5fxJIg+yojAM
+czHllQGi+a/39Btsu7l2dA3794Oah6nhE5lhibPivjam3zIHm0+VbsBet7/VKmO
GWcpoUdz5z+fkMfLS+HUf3kPbI+Mb2z2fS3ofy8YeBfbtNKysZod/PTMMwxL4hP+
/M7BuOLbo/6Qir/45+Fi8c6s2mpXD4lIsRyya8Hs+fJ9uT1qnRVygfcMyx0lFDLc
pPyI/5/LvK9CYQEj36TqXcrkIfjwy79zks1ljVD5V7ohA69uHO28k+pBeBXD4u1i
yi4nujpBPGJkAU1AAx+54umOsl5Y76XD6A4Audjlx++/wfDgjDlpr1q96mPs7Spu
KRxN8awd4u5ZLNIIt4z+ZcY1tsFEXNGyyqCY30cpW4Zo7u17P30H0rWuw8ozU8kU
TztP2RUZJ/4NVN45MvfLYXw0x84Jru+antoSz64ohB3otbxwrFTX5uaDkq28s5FK
sQBYvLweJBDaZWfhdQJGjSNyxRa9kD4XOH1iHuXhxsC7S/1S7tR3Co+9DV+fP43S
DSFlkp8eDDe4XBZPRZv+62512g8dcjfI5PbImm2V4X0krF9mtLgjz/U7fOw+5o/D
zn92AhEslEJI766DqbQiNMmMxycLudfIUc8DFCHvU3H8R1zBiUdvMQPBAVBlp/LL
qn2k5fqMDxLJjU1btQEa3MdwEULnpRFwQOWQLG6y3soRUBaI9ngTfgs8fY3wzs5p
ycRGrx5nbE1g/QFwH/AKoQx1tolHpBe5NIb4bQ+HAfw1ZTBtX80Wj8/8kGvjel+H
nMixP8L32tSVH2pd39bRHWkVISwXk0Lgu41thKoalNxe4NG4bhFxtcMb8FYxeBBm
h5Y4pskLMdz5Y1usrPh1ea9buSYdJFKQCk0v+vlpEH9/1w6Tne0c99mLrGra+STT
JXjI4YgSf4GNqfWsR77oyZRWEIaXuXFtk6EiADA2EWPI70pNVlf6hEHLrDHy+nh6
spm8+HBeGbtAz7Q1KNAFC1ddcZPhluihJltWVW8BXMLZok662QPxCsKrNTZEtlb2
4Pm6JOj4KcD/gwC7id7/v0Fi0fbcqJxGe0S+SlPegnBxNExET6iqdpKu0rJexQuF
8O71iUW/UqIuGwYOK+qAWPqwr63/7knMAKzzaN2KAxRRuv0+yJxgi2o3bjYH3pk9
NZ+2zXrr244Scg2UjFbBqC1LW9A7KG2bNx3iJjOLSmbc2g6/gn7Fea6i0T2hkAqt
r2KWnPkNoO4abnlntGhSbxexDLMkZx6HDK9yQDsgm/rua7SnPvDyWXViNFAc+lTW
1jmlJ5qBgbC1x90BO/XaCD8ppiMK0Q33x4mANEwwM1IeTOwQVzTLfsUTQnC0z7rG
PwXKq/vNGBTOU0gE0G8Bi3Ieyk60Y35ts0Bk7jEtVZgcJ+6OCCCJGO1hLrJ3Txqp
EPyraqF8808O3R9fAUBGmILxWImQuvCCbpH1qQTxgT8bUMwWvWx5flhZ1yxhr1Zx
wSeaBTXPXDcwnLrJmtNPTB7xm5Hxe0ehs9m0PWxgb/SQyVRB0NIcpQMiaYYrkkZo
lqtOpHdv0dXi56hkYAtswysPDAkzsr35lIMvtzpZ8QYiVp/lEti8uD9FJJSbWGex
rVGZ5X8/TM7Cnff2hUykv9nMp2tfIQCb/HVC3v+kwUWAzXG6m7+g8qc9vyENSyt9
g+TNEHF0RXhD0QQ+EG2wyxZ1yEAxBtHW/5bgkCZ0cS75appuh3hqjYEXCg26Gz6T
dTnuXO0YlRuMY+G0PysZUmofrsvxnBDUM44+mEvqsqYWRsRaO6Kcv1qpxIDi5zad
N3QhazI/uzPJ2KOYq7QcvjZ71t67lWqtnMwuhBSmbMYGXIf70kIR9t26xTkymEKF
MUw9OZRPRbUQl3Q5MGAIzjzVA6+y4+olMRctAjSifAi2/QQdBfSp4s2AGUM2Cj6L
kU2ZX25znYLNqr40/aF6RxYAPowAGRIiLGH8DvDMEqYJINpzAX9ywNpX8MaF3z9z
+uofygwn0KuM+WZUj9hstfdN+Th4StZJlgGzbM3wY4v/iT2posalk5vW7x+3zVDU
xLKVN5gzlOhu32wHM1ie57UYhS4wgX6VrMvz0KCbb+ej3rpOyw2YX1l0stG2gsFw
bIUTOpizP09UDghbg82jzpPW4KJwe6fe/HN7Lyy2debM1kFT99jZLg5MfqVHrLmm
KN70ItqEJ7hP6zo4x+X3bjf4B0VeIaEZ3aY76B2EZwN8cVjtCecghm2uraVKhXYV
RwfRcHjNyFycEURKT/pp+WWWb2G3pVzksduQRaY4AxNIMSFzJ8ZqjEejJKGLrONn
xsViV24JZ8yahMSTMtHnz+rUATQX8wEe4y9mhmQLzR35OtkuR/nrGOMRs2PqjCEF
6tkaT+ox9yhOaIY1ICXcqOAju32N+yO3MBDLRnnYDv6dXKAvlMDL6cLfNVrCahlm
ZtbX0SkMDKR5srnsXqaDOgdkUVdayUiMPGjX+G9mblD6Cg3kOsq+oMvvA1OaOSGz
1ab5lMjrXDNDoWRXHCWuxt9CMum2kWjfaw/RW1nOd69is8faDOIvA9POeYIBRfBd
5WL8l1Ex2u2Q/3CnFJVzJhUu+KepFYC13gYiRdJHzZnRgN9lFxZsynNYhTPs8Jyc
TTN0bnqcaNuxU3kmunGuPfwQGUxi0y7nb29YjrDwzO3mYixlvLDY8b2qBgCWDIJU
nNYoBVZ3zDDK1fgnBlksScoPBeryv+MwFFIa4HEXho6b0Dym+E6TSLg4cB9w5XFU
7G9qTkLBilKHJ2q0PSpNMM6bYasjjoncamHQT0y8zVyhrjxElYjoLCw7/q/fcY9K
bQW06XCwptVL91ND8I57cGqayf9LWrb+GjBeuqinslYODbrdw0IejxO+jteDPUyh
7ly4xyvfsWRhwGLqTQHBWds8hZEgKgyOoZAqlc7HE9R7GisyllRxeZhYyGrGf03N
qPROhvyRDr90XVVaaSl0COKEWJN9RHYUuX/udFITvuUp+9IbYZcrWfYsB1RZ8VIx
tknPgFBdMInfsrMvSwjFQLFpbcU1yaDGlgO6MJFdskjSdB6UK7DC0tKslAo4eiZm
89tL+X6GDpEJBbeGilqW9xEdwkhCz4HshR1tHVBQw3cYbFibJpQsS71Yh8PxgEHI
cynR5zV12o44uJIvmsJzjLQYCWREWcItG/Yqf6eFjSK4w6HdrrQKj2gY6tvz9WT0
glfUFoTWheOPIcKuNEch9W3IYwUO+AXCAhG075kptDemMwBMCpF2yAvjckRoTgoY
8+kaDUDnTV3N29T8HX3XCkjni/U6D0Uzb1/+Ip+vmqZWXRQnhf+fvN2iiYmnw0Z/
fdkLAQQ2cV2nRr2uz2jkejoW14r20o/vcB6mGTLUWoo8nnRpVvZfhEOtrIMB2fc6
5oZ/q7XDCJM8k0swLOY5cXIRlii2Mp07Wt2ppYiiFoEGyVY+jRYfqbgd4k6y//wu
SzdwXkT7bZaPJOeI+19izBQwYiB6AE9j1SbAvdNos4s9xYf0NXjrf8rRVC0QcGX5
V+8+BdpU1rctUeNFpFfPpvI53vONk3k2I6GLMtBV8Wjrc6oX9QPrfU+uZJu60egr
/K8tmwi+ok5OoYyuA/mo6nML5dNBqtF47j293fQ35KC4FkBvwNWRXj8zz2pq9sjU
SWbJXwlY1Ji0QTBYMoymCzyP5MapqOEUFgKkLEy9OLC4X58tAfSZU664FLDctvIk
r1pOgLNsLD9BIxOOng+dZ8s4oN210lVDEYZ09Dl7fue6M074PpbRAjF15ZDZG2mG
8+/SdSnywJ4xplWI6l4tdVjHdhjBa2b/E0oRaa1SmuJCOV9rbE3YNOvShgXRmiJY
PkJeKc1+57XL5YBpBrEQOqgymchO0prTJJquWUCEfRMWbNOKBl5hOrzXqAhhGA6Z
S8vvlVP+ucMSaY6kblnlEU4qWBZdkGvMJiIS9NA1NPPD4Az/M2cW/9XpM9XqzVfP
wybjBOX6iw3n0mjHBY/k6ikKbKU4DkUlHSBOiuTrSnBgwRr3Z4ehSodRqPaGT5M7
gmehE77uyWZWltobXZDkl4JLJjt1uZnEujg2nzq8+R/n8xSoArtdRzhXq7R0LZ98
Q5OjG1zpK/QmkRbIrMAlaxOE5gnqKyphT19QzXg+bWzTLx8dLLSFVEqmgSSDifon
j5EyyV0Nh5nPudyJwOtdzxiwr0YMwftbQKwaaDebPztHEqjPLYq0JcTYezgx1jY0
+3DlHMbA/g9+41TbAAVe+Umf5RqbA2C3t1NWpUnRBN5PhnvVjjrkxCtYqi+hpUDW
k+Bh2Cqy/kLeTAneEVmQbIwMDmjdoXZ+l1uh+XaQMIY5GxQ8COPHuQVg2vReqSBk
D3lxxSy8qPcbdj80w2KqMAW5m5+8ViJWNfQCuRg5hnPSkre3C0FAvVK02zlZVcHL
DWxWvB/AYmYRgCun0iYcPZjN6Dbq/d88qGx6zmH3fkE5O9xyn3AN1vYmdtAqx0rk
yg4SsZcA3p3vq/Zon2vbBAbWz3hT3+mMJzJz7NzRPuCDWoTXFEKzfLs6J43/lApM
smlsreT8oXhwjoRlrPWW0o5ZyhCxIhA6amTwwCxFYWvJ3Gf09jtsXk1dGLI8lsSk
MccOM+VN8rh3Qm/uQz/eD61IEobjhGLFmll6JXIDpzIDcBRSVg6hyYJafs5pTbDg
Gk90RI2jdYATIooaXWHKWwKdAbsFB2PfpEerab4eY8HKDHrY39L1OhGJsWhVTIpZ
mlt+ez/H44FQ8biTdQjBfJAWHW30ApD0vY46TNUmfNbyX8zi4RN74Ud5YbIRGTZc
UswCMW1jF/lWP8Ajc85f4UgyusJj2SvM8tKAqHm3s3nKG3bYacigyU6SrLm9TscN
iV75yb55zxhZlUxfR6Tb8s4fHOfW11MgMQmsrPNlQwfsv4z8cTpqct0dSyoQ83B/
UA8OiQCncMNmn3Ay1A9KqC7GTBzwz9tk2Y6FxPRZvhINuFwi433jANhi3vrxgTk0
XhJDResqdRpn5/jTGXJNMm6oxhC9mtYFu+E2iQIE2FRkW1NCbNX2BbqbM9+2EK00
mrGOiPXl/CLCZ4yS3d7F/PUWEXVjMNV6v1o74hZSpx8SH0A/5RefTk9iRmCR5bvc
0EqGJeivVa8xuX+jYAbQ/yI+0w0LYUfpx1FREEBdKvuE672cZJSJakTDSw7DCT2b
siudikNYeSQaDCK1wqIrof1KQV1F4juNa3Cu0cpxcx1pDpAISEW3vApMhYz50y1l
N93tr4uSNmHhwYiLo84V4p5qp67RkuTZ/gQcTDXwsli1tB5uGF7K8w4W7qKtAR4o
p1sA169JykoZ+vZ021umThO+9NNY0w7/es3OEF18+r/8iM1l1or3v7N/9Mw0JWzU
AEiv1iHiBLpD1zdrTm4sQPcHy1bf5rZBcXjjTgdBOnqgN/5bDag2DHuOTMp4n0K+
DibIR6QDFMqp6U4tYhjnQEj5oDT+keJ+XrQV1SVvwdxxurbbCa5EOS+qaSfHgeF4
ZF5X6njIAlYdx033PbOinaRU1weXt7hPKFNzjQfksFW3LDRmONykydT/vQpaKPz8
tw57SWfxJE8QMaE34PAKQkHlIJrvagXO8S4Lt9jGadzeNmxwl9SqaZYjpp/U/TVw
IWVFc5XZvXaQ7qbVuXs6eSZkjDjNj2Xv1eUOLttijeA7xEhkirxIC+ZglYoZLSXj
SaFSDNekZmnbLpiKEKIysc9BjZ7UCu7Fwn/If1mLZhWUoUGroysThoXe6ix3O+Ts
4dINCmwtRLE1FTJqvs7bG8jrQpNkTD7uYB/sbVFTnkkEGwKvJrwQaHrm48dN8onL
8hRvsS2Bqv6PC5ielcOhG/RYJythQYPxwhWO0dmjRk2qeSbeUZ9Vp/VuVcM/2HAC
wJkAJ9T8fCSsIqwGYifh/KABLJnDvY5SUWVmmdEGgQV0508gLD1QCrVSBlU7MhYs
ofaewG5DybzRmKAy/daXjbyf9d1S/Oa3XJFmksMedytlZkLNiJZfHhl6UhVyc9yN
cI72vi0Y9LhFMzO6Isf7+32PBNNOkrETyhL85+YzsvDoPVzRiruxo/9zfVUMcdnr
uLG4fd1fSUcos9suYcIMP54slsp71iTMzPMcFyS7rP7/n/Uq4dTn/g8O/IN8rpPB
jSrjsjVMs99Cmiuekbl3lT/d2EBAnkR3iWlY/DFSK8R6innHX8EsaIUNtn2SY0km
JECRtRefVbwoFEUqakWW6+vn9/+hIDQYfICVOKqFj89zIOwLsMtrQYXH9CCstV2C
PEUf9CNAM7KVVbudrg0mOpVI4rBERu5MZCLtCbfqlD4FFMJYrAT9cSKA7f4tXHJD
cvR/I5RSWEEQUkGd0YSOZ/gv+Amv2MFjECwSJdK0HDRr2PntyO4d++vDWA0eW04C
HQCCyIunLPXJV1jXhFYd4jJi7rsOnXryRPTacbCpY20C63IZB+ohNnpuY3dbOnug
6ZqWZwOgz0EdZbyAMiG5ST0uqNvOYC1lA0WsjUKjVbzQ/oHpzgZjINKpxgryfGns
ZUAPOkfb0IXxU9/t5Aja81VQXIIiv81pYuTT4s+R/69F/Tk9cbaaHjDBLshadK6Y
Mt+NcqKiRJ3ByMSyR22wu1ieibsDNQraKdgqfnGXpFu6rIPkyt2vaGOXIJoM8FBV
bNNs+7fSssjZyo7bSi5DUiLujM45mX4vxMW55Rj6RKiGZtpmI+fxTp5vplMo4Wdp
6Y/VZEJUtKBo1NBr7GC7HEHxMlYuC0u0WcHseiJ9q9TPVmQBJ8z0H3s6Y8brp1p7
4JXuXnpwvO4VgZqWo5p3pAf4DP+MY6Cp9jFBjpRj9UqgYPK8OeeUyXD3T9Iq/Lyd
R8Zja9N2a+u/EJbe64QwhJY59Oo+C4mHrcz64FClap2JJ48o6LTC8Vj+fJrrirWo
cgFnD9BUXt63yuLt+HzWdljlNas690912ieL9JvTNU1P6KHSvxkI9YOihaIz+o6P
rz/taNd7pDdmgBECsx2QB3hjqSmJifFGpvr9nT9GFfF0L1uw8HGtq4NNmyuBzJH6
pPpmNncT+fqpx3tOWqTwPdiaNVaKwMqUy1bVsX8/pweHUT81aaT5Kt+7qlhDq0k1
6sM9CE/jq7xnMw1grfpj8Ysqfaw+QjbyY3h5mhomb/onbtBjskFORo1BO2GJB+3p
PLLygCxME2J4QO6yt5OVWS65bLLfFhvK91gQhZymOfl99A87/KaIF9rg7xON6250
9NLArQpGYqal9GHSMskDX8KfNUoelV3Y3zDiNMgDb2Co43AA+hmZQwBL1r+G/R97
hYA0DQ5tJBCJt5gqAGmTJdCFre72f0eS6AyxEiYPq5EFDqjImDhdU8TwQ15RRVL1
PDiQBcGdpIcp/FWDspUC/gNzxzSWU57Whm0qIRSMymPmpj7E7fzbVkU1vmfLqoRQ
JnPOMJNp59POnfwI7q+1BPHhI/9y55ZpTmNgLacuFJ/gvgxrSfwazTaF/TSMBwpx
5e4HKzHulHHbgxhg0x0jywImH+IDQXmiOFb2XPKLAdCdQ+KvVBj9GP86LVNnVC83
pHgh+VHRXl56ZliJrS6RwdNZubOg9bpqo9gO4QIgKuxQBmdJURraSuVjM7zYDrlG
KD2AwQy9kxQKvl96zLWysq2JQYiN/eXi39dSHIaJ6fmQCJc+Lr5DeVhKfpLEFd6G
AIdGugUwGOURmrGSz5ALEFzXhcBRywoGMc7B2hooalPUz2jW5jNWdXXnCtgXgSq0
MxrpXeY7hJvwshUDsp93XBRXDXy2g/DoPgMUiOxQhSRTzuV57je63sPRGeFvEFnV
dcZeLa+WJ4ZqInzkFDNb0rWgRcf2ew0STosOv+DPJaDauuK3bjonk8Qxs5ffRqlW
pEACc4HYjZXUjAdNgxfFnbnpMPkd7j2Od8NcoqvEgOEgb2p1CTBY+7f1RSmfFXbE
C7v6R/xnj6SZfWom9dX4RALRtgg/7L/ve4M33gd7jCFv8H4tUnVMN4e1QrIbEuar
fETQDwOC6Gsm5mRzpc0cIshmNcIM0kBVyud+FRFgqX6lABJaCnNej0vRSLVJ/+ws
yUqUlwdatOHsZk4YKz1Fs39v2Dlyoa+b9ihHVc3aMARnxF7LwtkaJ2FS8poR1HNn
jeyPf6258CUz1QkODLCzQGhTND5kXOEloMFL5US2UP189/FvWdJWJHjTJuLC2+B2
rWdKxsMqaY0dz86sWlYLadLnJtAJOs9zR59uPNXtnh/t7uDwFOVpXh4MF3bpOKHA
p2vMJNbxQn4QhjFIVlW6zXpYH0cLSHWEM006kEONPSW8TqfOqpAE0REVjxOYr4pB
vNRNHCpGxG1kKu9SALe7+pl0rQmUGXeZR9/gL/Ee5FOnJ+LPMIhmM944bbijwP5Y
Vs0AW24SOyUcBimUH6y0KE5PMH3OUkV5JOPgvX00QKy3UoT7K0uVru9QeUIfn2A/
5SNfczxQe9PJ0dD/clztjDVnTWW/FKZgipXCD3oRt11j6uZq2eUorjz/vVFLmShK
pKrahqu0LrU3Iz/Z/ll4QIRtHLMfCf1ddLwj1QxEVdascUicxe9G9zB/UZh8+jLc
NyxgeD5m4mufzlPQdnOWC2R1IEQG3Q7HMGFHTFMiNKlfIdtckB6BGaebbXuMLfpg
SQ3lBnv+QNoJUv02Nsb5SaWT126kSQ1uRBuodaDbnZcv4zyVT9RjYMUP7cChlZXq
9Q+EmYv7cZ3DwtES++W9KRpU9S0Q7JNhnrB6yeZ5w7K8QXbneo9Qx0u7HCrwhBo9
Oxi4SsLTuqQmZGX14fQUsrumKhYxeBw+Zt2b5YsqD8pstd6MdRE36KgMSOzwF+ww
Wl5u8/Iu6HvAYpQeY9z03LxWQvK8QYBtKb8wN6s/p7Yyx+0yA0Qt0WI2yKw2OETH
h8vUpcZq0O0jo+TpdrzzQYMoFdM91IolMrmORgxrAW5J09huizYlfTHwlM5os5QX
lKqGFPZkbH5tCWBpQoEfX6gKj2wEeJNeVHJ1gopE8cdT1UaF9jVfAwXrz3NDPnic
a1QU81WCv/5CYfp4bUaH4RpwUfnu5jFOit/feDRQiF0l9rDm9AUhTsug2g5rCRzV
PZax14g8n3Pfzo2vYJOHT5FCzOZ81vb0+/LlbwbJG6/IG7Mq2TDrKlo/3XxKfn+0
1GKmewoVq2+OtRPCrbt7AgQCfJjssqe2GGYNm66YgUdZqvCsVWaVCVbsuQ75zfxn
jGN/DDR1oK+LEmmFPAU57k2DKbA0Jd0p9wCEI3LUg70v89vAqq4fz4cWDGaRjIX6
N43WW05xfa3wK+TGhI2NPnstqYw3bOsi+6wVSWyKse9vG0K6B2Lb9nVIGVIrpji3
Iva/K0Bv2jDx7DCc1cOKnNaQisJbEWAvyaRxX5jY+ZVEhqnmvwham94YDG56rCud
BgDXWpPAtvDSBFRP9I18pX5rp+9cGgp+YWz+NgZqZcXfCaNj0M87iB49gqk/olY6
NaeIFnvdQAvGAxsZGD55SlYjn/nqj8Olcsle8iFWuPua9IRdRri+/tUNI8ci1QzL
m2Hlk+gOnYHenIT+fBZYXqv9SVaqDVcVQlJ+5b1193Rc5Kd81LN9rzTZTcNj3z1r
qbVEdlcjOZDBj2tq5YFBWMGLEkzjTxy5vn1j0GwjZDh4EvjF5B7Dc1IAoBjeNlA0
LIgPMS5FfZiPIWKHpWJDIolUwC3nhXxKRN5Bnri1UDbf5fZaoQqMz36NEEHCNSt7
X+vy/P8+QX4BkTFP84OMchioRgRHVa7sYJxnC0MJSemqJfh4C4hBBen8vVCQi7so
HJ0mwe+guMKqq/YVe3zYK7wI3bIvsE5mEtC1SARXuxMA9prt54dZg7RAJ6ibE9e1
mUkZvr3ZDyXQYlIKGtYGI18lvqXPk2Xvklnu39KXO9zOH5KD7EqyIAqNREsPct4t
9NtM8wFnnGYtv3zmbWO2wT17Xj/kY0wjgVPyc5bICXV4SKbzqz6JkNua8OR2ADp3
yJExmworgYP0A5HTI6pUJiNEh+0aIsAhunuHK8HgsMMJhoQsDD8X1JxsKz7EofV4
ggBKZJRFOwSy6x1huy+XfxXMdRWIMuukRBtwR3eVLGM4DQgZxQ/22yHuFXMYy237
trW0nKy+NL4S6+KV5HzxOwC/lpLAxBtGqDfLfiXSW5dd/YPpopV2x55yc46BGArW
2QTpLmHEuBDXfjVrrv7gjyXBWQi2TazRL8Nexl59El+zp7lnda5OLXioTJpdKPN0
KwIgkO0z47LeI+h4+3DVwfQbZBznPs8aNKmxSTbVEGllEaKsmHHNvIBgn/LZDTU3
tNISzf525dMZec4kDee05zPftJb0asOJ0xEOcNQNAn6Plb3wBPEBg2BD8GzVWfhU
xknSY4t0SvimTPGlaH2RVgiI8vDyJVz1MjFSxTI5I28tivTfGogloSCmmeYOf2FP
zaiC8gomo8LQYVJvXvKe0thDq490bhCdAYuQtwRtdnXTW4hMzYeXs99WVNCwCcA9
SIGkzg1p34IiJwtAc+jVNjc4/MfiiecTzOGUOdiNzNg1ZjNLLq3AGXU+yxS0kbGE
VXj2MbtdMw/YJLd9m03koAieKQFE2dlJ155xrQDi1BMf5v/3KDsHR31/K/WtoiUe
xmJawyAg37RhdomwQGLWQXLYglREzQYMZIl7RFvEequ3YFL2fk+rpUpLqok4Qu0o
zzCG5b3WH9B3kTD+UJTXNMMEqm6nenIfncdgkHb1dDKFEWMlWSO8gyiTA48j+9Do
Fmsmlr2CmdVC6dPcqialTNy2yzUNArQD1Bk1B1DKab8u2QzaBxw5wLeCQbcle2x9
8eGuGMLjXmFoMpAIlkRAKqNfwwbEXeFLzqg2XMgM7HVBoQJsfyWqrqYxW/TDkL6z
CoRXohKpXd+yYJv6EjG+IUn4xxI2tQJ9RRnPdqeaSf672ElgDkKK2lOhA7ezwEzp
yhPYhr+2E0bTIsVheUpe/qb0sfe/x8KFpbpokChtcRQtNkkeSJZtGgzvhiSX7NFI
loEMXp378qgU9oH7z8LUV5byERzg5hxfTucAZuHKIV4d0PaagDswfZLgpp7QgXYK
F4QdHAkjpAjg446cbpbdB5amsJYvUo2zoNK0f53cwPOHvVUq5J47MCSXPnoHVH/z
4x38d7vS2wyeUw5wewlAG+ZfXL37lISLpHne8Qxz9rjlD4jtbIlaKWhol5p1O2Ib
K22lG9eKNKnzO+im2D/06LzUFiH2nPGQRFUwJg/Sgyo89YHkHvA/tm+WndFbzy2i
h+aYn587vD5zC3IFGKoTWk5S6wyxKm50eveT9xAP9jRI06h1+ayfcjtimABBc16x
eeyiUFTvlYrNxDZsH0JSpGMhG7NHCVyYMoE6xipnidLTm5FfmzIvfeDK4Klup2NE
Na9qVqSqU9orOLS5mH3AX0cYBg0SPyyrjsla1Ty4uUR/iwB9B1SI5X1CMYqQYPBs
Ob3HzbJU0Bf/LlAP64/uUz9Crf6qufRkIbeuEsYq69EsKzh1m37/WThLWwMhOfPu
HkF/xduNJMQTCxwDxqSTp26QqaVURRlZstNcBZHvETMSyUCPHMnuJgsLnYdtFOHf
KjsxBOsXJlyeBjd49YIlVKIqhyemngaVa8lXEHtNK554Hqrkl7jQT3t/PLwKiQ3j
pVd4XkUd6KppdTioKydyKy61mMR1JPJEfhZKn7h6VTie9o1N5T4EBsNz5VhnQa2j
L3Su3PLDY7g+29VXDvWSMfq97EO/7LE74hJ+eKQ9JohkytMgTqIDvKAUr7D7w60Q
n4sKklH67H1R5FDcoOq/gOq4IJhIwG/ECOHdda8ioQoyJGCkuICfZdCmNTjRFiS/
6EJQVL/wmHvrLTlH4FCk/AlbrCN4B1ExnGFnLWu9jPKApXDkGXDMN+DWgd7l8n2u
xn8ngASsg5B8RSBfPbR2SuxkUTNKjeNm/RJagX4ErwS8lgWpxx6xPiqyjYWBDuuG
e2XCP6gKUlPTyvOe/cbFFP6EwVzeNAjyfS47H1yAynRzW08PTxiBS7q3TpH06Jg2
45MNttKSmxzRKsaDULxXMuATwlJd8P4E+UlsBlEFLPjFJKQIIh5p76Iw8Ak2BeMe
cUi3RNXnrNT9psHk2SHUhydrQv8uQGnrUNsv7Vpic8lq8HDsbpXZZqSfwmkTJrbt
2LvRlJl1rTy4ISnNoqtsU67nmmsa3NGsl5bY/09B2iAaPXEyq0q+sl6eMWAOA8qd
4ttqQ3tihUfIuNgoNCWc33qiecVI08oG3yMBaZy6nNHjnKuRxGR2I8k6wbn0F33f
sNbYpveUhfbb4WYEG56xMsCteAaw2KSZZU20TAehfhkcw53alxr9lovaEUMl/wfe
sOIZH1BvEjdNjy6ynWe8MjMInpmwgAduT74rNDIGzofDtvifMOUcGjBI98Omq/ey
CQX47/9y0Cs2m54d1KcyZmQyrJl+j1zjLverRe/ha5zJOFT2JzsvBAfI8o1YXJwc
86AOvGtb2mG6SQKgH8C2kROOeOuHnH6KyaaXHZhQT09nylZG+eSaJ0f708VS62Yg
7bWGJZRtxCIFknFjknzplU/dEgSzRosc83JP4HCfuN0ceKfhQPBeBuwNW8OTMWbJ
xiSnA5TCVOf7cKp4o2c4PdeL3li6Mq+b84hPo4Cil13dyn7QR+tGIKpwrzWrb/zJ
u7dv3Ei3pK4c0GUZyqS/i4tw+KIWRgOWnmhs63/5iy6WQ30tl26uN+0wauAkJcTn
zr2L2JCFhlQznBCfeD6mBTahUV5RRR1OABvD0Kdm7ZY6qfGOxa5G7BGc0RHJYX8/
/tPYneEgnLgIHAEREriW7mPym7qkMs0votzMzHgOvCCKkhWreVChE8Ubw3kTMjEa
2gz40H88lCx4sNHULNQQbWOF15aC+1F0JGaxxwWuen4Xrh6c9bkfaabRYBADouhD
7Ycu51vgk/+RDjYDXA8tTnG//wnHG+n8ADWd6ozE/e6vl3VXklDGTfsiT/z+dyMI
LVIHkiE9EY3yMui29U0hT4LBxDTT3atAN8mbEk6qMa58820TUGAHLjBp4DiX+NKs
YGMiH37LDbOlyo5DJ11M6R4v5WpT5nkDK8aU72WhiJL0mSAyolxhjXSGajFADgxr
cRq1AHvMmhEoavKQK11orZeoyfSw4KJboccRn8QuGaOULxXiG4HL3cDigUREqmOP
dBypTYgH0XKTquo7URgsFKXTM6oetxjIq8NwFA+Ys0B4cY1vI+Wy+SDLAXRFUFkI
beXB6dBegNLqdiQmq3PMcU/CmRC7xh48dz2eLe4ZTfJwWBEi72oIvFqyipkC0xZm
F1oKg4bHsMhNad/qT6YNtaA10ugVVtWnf7HDPCg4o02mr+IESXtINP3tU+YsJ4MA
ecmwB0hmzEHmZuZPt/VdJOpXyxTusmSD64wsUk0dvuT14gPSU/dbIjib0v4kV0jd
VXIKzLzGOwjDSbCUVFBCNvXIQ+zxAoyIrsLpi5zgd9VowBF/kUrjBpV7c6zWNH6f
pEKCdfoDvpW9k2x/Kk0BKo4jxCLg4aT/WcYZpGHDVbb+YO6j5H18HlretfYkp5/j
zHX/hJEah+aUMJGQ2kmlBhA+7uELLpDt/Y+LwAAjVe1cfBfGw0Fp78LhfbMfhjBy
bq+M93X82jzOxm50wlrNkdaWMUjpdIC1T/BEkP1AJ9TJ0/eNZCdpvsUn/E/e0kiw
wcoqhxZrqtKqf4J369xCQCz1T5f3JvVZIXhzdYoGi+1FcvG+cACdPh5305D8M+1K
kr+CZYN0j3iNVkn77vGuhOD1IOZ/dqoGMpGqhVgGYcUTCCTAGPvi5R17xo53ZAeE
HCHNh7PusDa2TaRixv3e0d1hQU07lI4/6LZA7iT4/byVmB4kh6oM35PkHsTuuXva
DYPDAQOc+ztwj/ZA38NB1f48uA3VZuOy8NeMXVOvOKJVSP9qUtydNcVOEVhd0ciI
Io91GXtjvvH35HpyVxAX2RjHNuKHzT9TXkmc+gtAKuX882tHpIIPF8F+FRZ0x/XV
D5IkFYM6aIhuEZJmBjNsmJ5HJ7FSESWZyvLNvakS8jWK1J865NJHLhvo2HL0Vb7+
TDR9QgnPwcjHrdb9ztkN4VA9GUukKqhpxCcbrTvkUOuIZrSU0qFi6mUQ4u1TpRJt
yKCUqPVGYGPHFDfH50F1wlvPo2tIfGEHQnHfSzufQyxqXWE1o8SuAgqlzTNzOhEn
Fr1ZifjdUfVh7o3E6qjPbcA1IbV7LMASZxdcjcqvMS6xTOL5ABvTyfBsppTtKuCU
w+gwuJxv6z1DhVWwInnhEmL/IEGkXPwLhsbfpLP+zSsEjgehk05t6R3sByFu+VDW
d1uoh/fVyZWw+8JIG8YcZjW6DVln3sPvqUdmYtegJt+PoMMYNLIsCsCddEzFTh1x
0q6b+4DkuyyDKB6dwSz7aaemcNgBKGhSA802qowsoiYacbec0lSjvsBR7VcuQAfC
dyy5BfrLzxhoLlrjWQvUmskwSuv9wUUkrFhlHlmyrptR0tHETv+sGpq0eXvV5gHD
WFOsoUOtATv+2RrNSEF/QFVflWo06d/tDTL4zzJeo9jUO8gJE3WwVB0YFCCzEoWI
zlwW+onXkefdc7ccC66wTgIZeJ9lgDQDDze2CoUp0rOzM4d51IyM9ThBs6AiXcuW
i/4MUQbeDJ7/TBbBWBmTQQtxCHDoOj850oZTD3EYsT4ZFUjyglBkhKSBmrB7atdq
ztlrp52ArZZqiUVng9MOTwnYFG1YNlr5Mpd22kC+raT3CRK40mB/56vkbX/4GFZk
XzgqRkl6rP/YWXTVKXdSee4F+BHuz+KEQ9lmDEANeLwZ8t9Ms+VSbArOyJgUk/m9
ZEwPEoopWYUD4EDoXtpVD3myC6ko30OQ2C+Xvi/B+y0eWac7jSXHJvpY4WykgMHf
jIaA8g5fBOeQgQUZtXPUwKX6KVmaktt0tLut/6J1LlpvXUAeYu3LzISRcaiZbf8F
qjKFgnk3lTSDGCdR24tc/8nd5bf/0FObZZieagwUJDmgF/gVNYQoo8FnUMbXNT38
dJzvqVMT5Xn6Rxlw0xkZJnKvzryBArn+/xGDr7iJIMrYcZA45ht1Mgfd8O2ncoFT
JdjKPmNynKOkZHwleGGOPgmIcan/wJmuG40aLwg891rMm9QOiqA6ZW7ecYLsrwT/
Mhq9mKj+gD1++6eAKvKs5BOlL3bhdRkNqSYnTPiUlXxnyJ423YSzy9gMbWzp9rJt
0Il/1soD07nXUIbfUWFL/H3SPzH9mOEUJSKra+ar4dak0YU7XVICuWZYLx5QM+k+
i4uWgkV0PDDFuTEOR9UDOy/6C1Z6kpvAd6HE/6mM8CkNBW/+J/V0WnSMqwd7EbXs
6KCF6BSC7gQcuP3bGF6BFwcQhNXf5qTva9a+hvV30KOM5gVF+oArYNplsr8IfYR6
886d1LRNeqSWWZXB0s0oaPTI5ahsf6lk8C+v7MDeJkikRqzu8GYcvoYkUk6V19fu
ytJ0CSRZtGFMOtzf1Yp/ENACPtreSyJqrqbHKRFo66ywLJ7WpUKiPM1w+XcqIjFh
1iETODrbDrsFno2e2JdUYMeyD+jl4saeDxU88xB6WV3nkKM2+kFVKQl4IPjL62Ef
5qIN6OqNe9wvZbTo4vv4OtGKoz6ZNchRUt81yAdIpdo/agrWVE7ctaTMqbroUP7C
y4gPXWSG6IcqJL1ymNHjd37q6ygTlsztGgpLCRwtW9kMj8IxdltwS3rB+Ggynu6G
FB8vA8nkM5MDE/4EjvU19vLNVzk49XA1Zs0wcmL11cy//hCS+PJj+E2ODVUY3rUf
Oyv3MmEFhHdB3NYhfd+181aZcNgUnWTsHORv44xEpT802WexVl991vl/V0K7HiBr
4Jyy7fJjaW3dykerss/6rjR761eGpeUWvp+2W6YfV5bKr8WpXnD7zK4vGBj1y1ot
xc54l9F1oa+7Jgss/Ip11L1apxvGYCRTuYAGesXsACL8P6uXmSC1zOVvIsveATBi
/8aawsVxQRGYvim+BgxdQNkTsWJbPqOvpVCOguCp0VsnDSTXzv6EDHrl66ZrLwJO
1Oc1RyhxvB/fR//Mh4ouopqxG9pTj+1+h2bg4cMcJVQscvP3cIo2TNul8KViyTLb
ge8sqBkYiCSzS2CsbvsiiIgy97nWpvPyitbtKu4K3TS8h+/qy4xtv7w/aWaeV1Hm
+RFXfKgT8LC2IZxxbWWkkTDZcMHNagh6xeiyuJO7W/wh8bqtqZFDG+VAnOPM3dKq
dFBO1+Weoz5lE3I4ddaVDr/x+Ms5XLpTebe9pOS0vSecQ/FdAi3WGozThHonSKoQ
k5cVCoLFNrJGXvgf1TOzRWQopX83DXvLnmHNhj1al8fdXyNlnKIEEb7BeXn9orv6
XNUKs7IbbvcVu+VeItfl7S8Sjg8LG2c5XC+DI87ssgi/dn57K6fPD8yCmETmb7Qp
EpKF/lufbn+XWJTcvoNORhlRKTQOiVsRij45Ch1hcoui5UOY3CL+bqz1vt7BDNhd
3yM4El6YylZvpJjkUPUweL9T566CGBQZN+xWaIH+B1//yOtSSyIjuG7vNJ7P4YeY
rr3BaZ3Tzksc6MbAnrZjsO8zr5JXEWChY9OLb/PwJfXAli6vqQO/Pc8umbIel/R7
qTAHykY6M6eiigHh1IpqmUcvVfpiVaUhzexBVckGWaAhn9HQL3wNpPVdbSZNgmAS
0WpSRjFYytOLLZf2oIu+/Ea1kYfNJJk+tYkpwxVo1eMxWZgfUvyxy4YF03RgrZ9s
UvkL09y7ze9A0h1CGq/WzK9ceaxQWna8sZVNjCUOZ0gTx23138rqMUw0kd3KyUs1
J2CDNOSR2a7ysS0TiYF+MlHJDhTcBaQ/5t+fhfCv4Kt2FVR6IK11L4YdyJMg2E/0
ok81rPyb9XgrsfCRktFSTGRvVQIKp5R/wTjQ1oG5EoCaqEz4qTPNxTdpxUCdYIWJ
5nO1buMUCsfIzBAfq6D40Wv8yNFwDYvTeCziw0rIDVJS59hUvnY+X+W7iCuHbUUX
rxyN7+dky6xTtZgeMWHbW7Jg62qhGNAmRnNWKaw53vAeQbB+UQt1IkgQp5UBUlIN
0ddSeUj6J3P6b6DKhuSXuXakFLDsBJlJO5xJNytHGybZfmnJvXAkaZcQDcjW2YiJ
tSJBmQNOQaGuTdEe+yK5fueAUwujI9dCzpMULFSXC7u/VR67Q5710/1/4OdNth3q
U9wKJDex7R+qwXf/zJgyrFtjhvXj0x5J/coDINvJYODqPjay9ekyOAE3Y4rm+V02
AEW5h8vCl3vGAQxRDq4Umb/h84do1Ia7Ct1pYCtF0b+QxcI/xZoipq+AQUurRMio
DDcp2mRV+I6hJ7c7nBHeuLNrtnGCI2j2Q74yqo7Td0ME5MyvfAY+sx96Yo92K2zr
L9GO1+wCMGjn0qMEo3uou2FAWJfND/NrKh3hp2LNi0UbtsQJLQU8fjHjpfRqwEUt
S2SuQy76Ijt71ZAvdcDAOWNV/c7zvejpAl+f+VzB/3DUJVatGcV35FoEZ/zsQyM4
BizvRmE8rQCDJV21Uc7uPKb0653t8dGaqH9ikTU6kbMK7W2opfwLlRg1iEa+DjIh
X2y544YTNANsPRNIiOOfwLjeLq/4mEdseWuZu+j0SLwLndBVeM2JHaB/gOYP12lA
GAROYEFPoTVdlNsjZNMcj+sLPT20Bim+HKgkXC8puYlvyDesG3DAIoNQn5uGcHqV
rE2VELNwNf1tAbSydE/+rZfhhiE18M0eFOu128jSVX0yogz//XyqCGihdZtvnnfy
art+jL5cneu+P7Sl7ubUcU7E+Jn0DEG+B1ZDfIEGaFGHZJl9za79+bVi0TvxLn3c
6LgzQ6f/R6vWLVgZjEP3gYUdCv5x5s6wxu20g+6wpo59UA8BirKQ9gDp2gSrM8rE
Ggv9K0a5P6PK6+xL8NhBJh1yb6lQTZ0e+qA5S/XXUdvm64AuhKLLiAPUZDAkaEe/
yprNvsMtTp1PxVr1g4tyLHCTgymh8hAaXKG6B5U+UjarpfFhl0lOCLclgQAz+ucd
akP4DlIfA2EFrJqP5VW1AoMM5PKkp1Qa/XtGfqMqiYxQFmjU/299YYgjQpHow2u0
5CVskO7Au5wlUFKIbB1lFHeBGliwF5440N9hvgPNKtKhvfcBu3ktwRFbhSnI69hz
jCYXd6v7dTDg8B0rLT7yw+oexk3iX7p3uGVuGp5/4q6rK4D/Py6twWSIZ2aoMYTS
zJ6iuJLsFLPrBEmO1qDFiRFOza+3mTcRVivPMCtDm0SEUbvIKBi6Jwzc8q4LaOES
wUm8VSAk7qMCG6sPKlcjL9pPyfyRBK6kkRJ20u6VdiiR1mTUH70uWpCy7cU0Wc80
HHy+O+lCv7IOpyLD6vwJwPMI5EXytkDT85MwrnQjCo30QwYlXMW4ZVu7lRrMDymv
/2er/H8ruWa28tiVhwPH/7lv58crFFVgDsjqp+0P0zGJiHVTUlm7dUUueqTahwOs
TQMBv9m8IG5VqekP/uXMbUGg1aZ9QnuK4gD2lGsOHXysb/7Q0P8J1fw4ERHXjTrv
fGsIS9xi5lgVHpQj4ROc8iWpexiNL2P/wBxW+7becB8xWZfUvDm+Eu6LyNXGQSdB
z227ftlUZDdhXPGxOC9JG+KTsMH7zRpsUHyzKioTXnqlPdK4v23CEKO/Nv3GgK8J
M9q2ZnRnqDzJWqZgKFC18Za0Axy9D2F3V/lDbvUuHTfC7p2TlMj/OCzKN23GrDrg
1Oo7/BxgdDDzUgILUgMRsDq+NJ4NSwvGVwewB6lrMMkTbYo+EVE6JqedVLA69Qgz
fjutc87x1vQ3LA1nWC5smakyqhSUUAPauPQWeSVbezF3/zlOOPkvHvUbhHNB5FTE
bxOq++LGWuytF95mW8JAC8h5tLPzuO6DQhe/Jqvr/LMb7M5voufVR3aleqNMNvsp
TsjT90SkO/ObLGynaYvyG4D/sBeTy1kGz/lRH/8CFYkuzXmNzEirfkJJvtg+ijCt
JuCMoV7YLuzI4sTyT8mNV9XKsgrE35UrqRClJxgIoRX4VoYynNSzzxnIuJhBa2qX
/e63f89oArcPx26Pw4vQP4iN+DrAeMgUPK0U3dixlviaUqm+EKBI4jCajGVVA8X8
EFiPYQnujSYq4ShQd7dVfvY9UGyoBAh7k03sFz4eRcOmDTmKgS1VJ1lbHexteiYP
MLRccngeneEtNYBcy/G3F61OxTAgQU2MEHyDwuz0LiGjc2JpoYJvzJEhUgeqqp86
sOCNh5E3hErgzsD3Giwu2dqg3vz7AodALCRWxVt1X7BYBD7LI8qrObYnPnzfP2ql
ZxWfY6GfQ5p2bvAdFj+OF6yvOniQXSmM+uWx6WPk2cX2HqKbHzpm6EKIF7J6Y7E5
onCgk9G4t+aerf381dkqdmdri7WiXwLgft90mDxAL8Uk/SzebhOymm1FFEZQTQnr
YBBnsb3wuPH2YKYMRffTySHaHwCJ55QirDQpvr91o0bkWBzT3oZSV3u/LwETDVdJ
AN7TK0nM7GB4kTfmIlLCUxnetn0txOn/ocTvAZU8/uSU7IaOLoF6lbuTqmMN8KoV
AhhVDEekOZWL2Dv1RRS+Z+JpLtj+r6WJV8Ltltdowa1H7wxEvY0D5cKs3xyZEMyx
cufE3UvLAhdY+NsKZclITD/B8m9xSobXy3l1OzMlHMXSSPpgykWplurt2l4uJwYh
4zuWkWfiOcmxg0bE7cJfne067ngUGw/1m8OUvE+NwRi9HEYY2a7OFZzZcIGFUx1z
v92QB15iNH7qVP/ik1603K9XgJc3s0SB0R94pABxx8JklCBaOSIu4z+LBjllULrA
pauDd+JLwssYnbToJaNZRVBCXw9IGUT8Z+WDp17nwlDgO/njf4W2uQ8ayzyhmyMG
v4NSOeI9Nr1uJoDLr43Gq0V3dH79UD8ZQphHFbr0yptp8u5LHQ8CZgG5qxZKwVDe
EnbXQt0WRa5selN3F7W2/ROUpxkI2sggilqy/qrGAKfUoqhTPtxDh8BxXZlss2aC
av8gui9p0TK2eOU461uVlInSvwzSMCFOPNusxgpO4CoKWGbcgfdwu19H8thgpucr
D5JTB0KhwCND+o2iByx2kg1nzmK6YXzhAatYnT4I7rtMQT81Oy5WjKEbbpO+y5b7
ErLoTTmmNez/Vn+XvyoMA4DQfwbigEThCVL0/zllRz7oL5E7JKXCS5ql9brD384V
iyNFAzAHo+K6e9Iidj92CBqsYqgqWFsBGM0vJrT1ZE5PJj6wpSWtE0jCVKylR9bT
khXL8OFAi8jwKpG2csr1hviaAD+RsmK1UtUpBIIn01kQ86U2G6/iLqSzATfLkXrf
kr8XQlRcPoGzTFvlo/qrr+GOuPqw4OzAqDFvHhz1CCyOWzKjoGn9Xq578o+Gqeg2
IEcDg3tmJQhtN6OFuj5xwFVQmNSF9fqbiAz8QPpLpstLnL2nme7oT6yt/zxBhQ2q
GLPk+jTofhgLyiWRNMEZxv7ZSYHTlhbUfkBjoLYJcMBrFb4hpgixHU7CJn5+6WdO
RCU3Y7D+g6qYXQt7HcrEj6aZDr3P2YA09/1zh+27edXLxt5j8okBZeTD1vYaAs1Q
gy4sM3NDjwRmjrpwCATlVJZLRTPr+TbcoPJhS1qcBtnAPjf1bahGwNa4pVBgdFKh
ivbB0YbA9cB1Sh/nIqZhSOdiX6WeO5ACR7xhopHNSdRS0J7zEk2MyCpPbDTN/twk
x/E9b1gVR2AiFiThdv/pEZSREZbVwekOR+0LxDntTZbtuZrxRtiPeArW2vdwynGt
uGOuUhG1esfJcTJ0lYJh1dLzzsUg7hzVrJQAcBwZAdyxqPfAXWw/JsNx2fGr7X4a
4b/RITZgcgj7kOhn2MoT4XSJmtTsV9wDyQzHlonT1+ApiYTMtjE96wiobMG1ZA34
y/Kd627RSs7PL0qDsXPMp1yWmCqwZK7UCQAElAGqB5QOM4lpkmUDGPgm1gsq4WFO
kVclAiL3L44ZvJoqWGPvkd/7Yn9Tz+qrLkx15PlAMBhOCj+Clyu86dhkTd6FSq+Q
SMmKclVU+5ghV2KLzV3NxleYFVtl7kc1pgZ1LSOhdp4J29r78mDJbljnXQpXGAp5
8rN+hU7WkItD8KrGDaljoClWnCGLGJKjthMT7gnE3gmiWmPL9ES3mCSi2QB6rJma
V3PNICTb0as4q1+tNY2Pk2iqM77DZGts8SqatuntVpdxJ+bpC8t7Oo42xwiF6ADz
OGvoESpi8jGekCilOq7Hy27LxpZWRGnSy9zm9WXF0yhnULlSy9y8Lt/zzE4YjaKR
zelPYoMjT5SSJ1HPecp8Zuj23YX3bQVD1CT2K2b75Nxm3XONZwRxxLBoad8mTFjR
A9FTAKw2qSjKeI+WkglaV0/R+EFXYTOn/rNBWHp1E//dl5ShMVdSlhiVHLZGQwXQ
09qXFMUxvcJgVUyJAD1MHT+dn08Ax8DP86STe+sq4r3US11DMe/mCOA5ZhRLHzjB
/AzLnyXsL1gEEcha5Jm/aRvL7P0vbLih/Bq2UmxoAvbPg/bYCqZnpCht3Cvh+N2K
3m2k2EFNKRillWf98n1lYSsUxpAeK8aOdEsRZcHI0iS0V9zGe0VeuUAYUqglljDG
R8bNgiwN+NYRSNbY3kLPLyLX1bxaGSn7ZS8NJyERIbAKv+4pxU3AlQgVOCjc+Ufp
1hb/BW4AqfznCEz1FtWM7nOMK276nSz2eUjPEUmUqU7Qpm5oLrOGl6zu38pYmtM5
ish/PuAta21745zaiYgjIEk4+Bg1SG4cGdimpq6yd3/sV9Ku8/8kR1TafsqFZf8a
KHhracgt4bWJNi6Xw8SkFbQ/zSNCz9BigNPn/FtO9QijbQqhf8fLY8hgxj3ZEcCT
PPl2/uBns7ir1W5+9+yKokhQPm7cy7DoTQp58HCrgzhoOM0Wlh/NO6sSMkiW3r7i
XVUjgRqgaKt+66cxOB4kwTs85dcmBnSVYE6nKHNEPqlP8pMreB1e3EhDEmsERP8G
R9rYtGqOCmmoWJ3x5O62FnE9gJa5nNkW2dAv003UtgSbXj6Qq4assDuXFCUZApZD
yhCIY7Gd29MzzuI0cb3nFCJNGhyCIm5+PzXxee+SPjOZiU/xHbREuH/1xAT+hG92
rVBXuSY3snsm/XLMG0jIbpW0qe24WPmIv4tsNQALoNBP98W99390YXim45b1ss3l
gE27KpDKbQdyxvutvG2Y6gUcWNiE5V7INkS4bt+CvSNiaVpmz9Y+4Hrz15LTs7rQ
U+LAVfmHRpYh0SYLEWNE9MruXpcoPIozzzzKEORAD1I3RFkW8zEB9BaP1T2zFaBP
J3w1DHNMnqGVdQh2tYGucEIS+c2rrtG8bVHwxZcq7uykXwq9mv2HFJ/ymSj788j8
HJW798stzlJylb3YT4ZJ+RsMeJoW7Jz6qAqiIfAsq7/6zdi+3aYlIsL4QQRldqJr
sBYbnPVLxAjwHcUWEEKDmlX+WYHvwfuNEzkXPNzMOwUJnIBgIJKqpN8rCMhRIt08
pUIBJnWKGBCo7cfDCQneNQZjzN4NY/Uc0FbxjB8qHdHlzhgxUddtvDW2fWX858Q3
qxQ+UG9PuLWNJHL5DML2XvJQje+wUMbMrMHSOw+cJyBU4ousJseBs2VpTnBs2M/l
7erbYwC5DXPO9e3qNXQ5mHuRiSs66a8UCeCu+f5xYtls0bRcmilwd/gid/tvUpNu
oMgM2WURt3jJ6XkIyK3cxiPxexrQcVXqJb0CEnChXu90HIscD7Z50+wiurkItNi+
fCKmKsZAAQEdSpOLwBmZOEKXMOJgy8rl6ZmU0g8Ispd0Hdiq80NnaU+KQ23qzfWg
zp5ZX1hnLUh28FoAzQ3mMb2WudJ3F6cwvx6QmfHy9Z5EQUET1MPiAPyIxBDmvAPg
ChhfjC8a9zheCS8Yjmqf+CSsWZswMBDQr6SGXs5t/IeFO6OGcyS63QMfVXtDfCC1
uCdRwF7y41uEwlu1EERFayvgUgYETZiQMY7+sFV2IFKzNdP+/yUs7k7pfVsXrYKo
c7u1kEfmlmMcilPp2DIos01MZJBFHsgCoE6nG4JAjojTKLfX2F5GxcLACprA8tPf
QNugQvGECpXgbdauY4oIWIinw0msRMILmeBXyKaUzIRq5eXpPw/93we3ekDaMqTX
AAZxPRVjg2c2F7Ecx/b8kp7a7Icqo/LKT1SbK8XnsELC69u9Yyfmbe62tB7Ij138
4Rl+EZ7fIm0Q/IyHHWb0NYtVfisVkv8yxzA+x7EhMPBCwHQTgymnrZGsYspVCUXm
A+mW1MTyh3RjKw25qPrNMmFWPKd3gud2ZVOTLHOu3+X5MNwrgMI9WMDgkPSPfZE2
hwTmzmCeskFb0zOPyfWu+GtcSjga6KybMXXyK+vx+sqJOBIjkSZ37+oUvjcrFY7j
YNfZnDEveimyWmpgQc7ltMKrnO3Rm/eFnRQJGOrBhAfoHEp1Kx/324lE37GfCb5/
j8h0Uvu2YACB0r0AFxH+cmnCNOfxhT3rBsKtpHlXHyJO2VF6bv/KQ96y3tulllp4
RRUxOJa6/YCXk053zcIOiP/gC+E8Q7fLCB6PKsmkjqsDKsk9CHzy31uU1AbmbzxO
MlexZFd/TZLa6SCMs9tDFn+ql7az32wr5irWPufjQl9dJva2S5of4xq06zi/0bat
JtJfAzYEy4p9BnvOtY226ViOW1Yq8afwfOP0qWl4RdYvW9YzpY1dbLuKEezhB+eq
OM+6PJu244Qk1O/PmTh0+hox5dRyo4G1eI6/yhsWbuzDmTXCUJfi/WxRN9K/kuZO
ILFaVN35zUMuR2iK3BtXVsr0PRPFyx1gcoFL7+s+uKbDAFqS59uk2H6EX1Z/dqxH
Yfwh/H8/+r3vjA+wSYSPY+UBT+fNynJEV9/774jkrDr7zPvnOs3b5jYaMnLvQFJI
mdqb6ASzfyA9N9vn7Otz8G0/4dWHCM4bqcedvdkasnOnsUN/YRXxFnZEsJ7hcjPR
co6SKMy1iO6PTS6nDW7HwC1WCcAueHKhNkknuJfv3YpYPHDbltxHsdvQDNWgR+7U
qZDWw9M7cg6+UW4HnV+zMWWXePWaep9HqSQ8Fc3PmNHaxuvTbNhzDEvDIgegM+Y6
8XIZYgy/qvpwwJwHAa/oCz2iGiECe76ci682YQsDIgHejljCdJMS8MN6PVln2yqB
8wCLrVj8x6ibKJ3WKMCiZY5jDAFuqLSSWwpT6YZz07G5F8cJSmKaGUhOovXW21VJ
hwswJM3VR19CuxNir+tpMRaOhzzpA+zbkrmOkonhV/1ACZNljaP+wVa84UT7jAoK
4lfXYWHw+6lHH7a3x+qy9UT6mhjOSX0Exw/qH9qI1hKSkf4/9ecW/CpXQ7SA3L64
eskCqCTU5OWAvc9km7ITFotMDKoBSRzrjz+fhvEmaijIO77yGfpNm80cDY2CYFqW
oAZIjT5aXxcOW6+S9g1JqHO4hFWGCRM5i4/z2A/P3YFSV4iRU/XPveQmTQo8Yl1Y
lqAxwsd2Ehm7GJNAF2Dk+c/CGKRd9++RT0YsDvh4Hv2pAsuxNcsoUkdgfz685Ovr
pYPHKwF++DhPoNtlFGnHVVdaHbGQoXWBVILx00Y8loSW9epSnFhsLND3fCuGNqoi
Oi6+9WZ8+2na9b+oKIW9AEH7ziiEXxoujEmKwrd1ofCwoZU0j9yVuu/palGeh04H
FO6H2HXKFHaPvg0qqaBG0zH3IuHJ3NWqh8Q1Y4vb68cHCoiFlw4yjh6bS3vfkM1D
IHeU5o0kEUjNdUQCWCdb/bSwNpkTA489rD+zqIJModYHSOFGXIx5lWERIHn5Tx4f
khtiX03b7BQ71m2J+ng3WLMdtSethEDrxgOsMkAEgY9KOETu+nx6J4A9Q64rJQ0T
0qQp7N/MFQUYdn+1VJS+OLS6iijzg1OXQ05rivCk5SjXMR+Oo6gHuvtUrU/PN6c5
eG+w8uGug3tX8jZtV8v+Gu7YtgCcI21z7V0zYtFM5I3BWq0ocinqXpq/FjUUjCiw
hquOMEVTUG07dPGgCkyDFmf33boxl3dlQjExXzpkePXG/YR5fRVL/4mcbGMQYlrb
+YdvT8O81JQMxAx+h/OSluRRcjiC5jL0NTKsTBUFguOI4F3bk6fkPvWTFAXkCj93
Ij+XyDl0dUcGiCqqggzm5BSuNlBz5iTDwtXdJNkjakkQc9DDaPJpU/Hn/cwhemg0
94/6p+7W0AurKsq0AgsF4vTGerAWpK78ys0S7eFoLiENyIOMs4WIU/TGNWAJs6lm
TGXlV7VO2YHD4sIati+7nA6+I1DAPUT2ywMfTJe3qw962JTlHNSdmfZ8jvC6wMtF
06RnZRctZrRfFQW0uiLYtmknEVXvI3oV7K/8tSzHlmqMho7VkuS7mVpMOriceGiD
n8zcTZz4EYvhKD/ZqAxzWKeq9K+W69Gj9MVManYdZBFIv+sya/Ex2txwuGpJ6z1u
7poXMTiu+jEqUt/BhaicvvSXVUfmfpS+csiXh90pR2fLDODV1Y3qJs7+c+dM4NRP
UpfBl97mWE1NAGj/L0j//uHtYMA3Ps/U4Hzvs2kqAgBMUywhT8trgQjresZg5k42
ql0T/M5dfKfbrNrAG4uiB9weeOYrhZxQ4VgxCgaYFqxXJTJRI2zsrBcgiMk1fIJi
Yy0Y8kzFPhyQgdbS8LctXr/jiE+DoBwRzUCv4rIBIFjFD9zzKMPONHusl1p+USDN
xpxjO3NYHoeagh6ucK/jmpjyfd5y988S6xEAmT6kz1Unx3xZyPJPi1Q3t1bk70Rg
wlpv3RpYRhO0guXvCGILu35MkZg+NcqYulKeONfOVSi5zmxnxkUb0DN0OKSyX8Wh
ydZVg409CBFNo3HhzkNYyLEKt9zHClkW0AOVf4f21YQMhlfTc9ZDp1Sxn5c6wm4P
ARMxbNuxUjF0Nc9l7D5eyZmiOH9IoryGADw8GWNzloVcmF1evp3D22yPIgZi5P32
UWiq8WwtN8so+jIJFj99q05YvYMs4O4PbuyaQBaUhN24wVULoNmW89Uw91LYC1lA
VGPtGOEffgtyHncDwzF1/zN5+nK2AwAZpb59o8CIoarw4y6poMDTIPpKpcWkZ39E
YvemEdfPYe81BK0Agb2PTh2Z0yu/ncHrIShXBy9BPll04sCogF9eqlOZrimWPQr9
nZDIJnwhvT88N8lltfQMD7ILeHGlZvYp0KA0nGlLxOMH3fYdDTeEn2wI55GBwzpP
FLWQR6JvVMtYI1l/rkggAaAhSGh643VAgVKe5gO5pLh59Lz9LBLRhG11nWFpacRH
/v8VmQNgosee42zX8RDJYSrWZHWTZv7FuU3/aqo8yRBeY+njvz4vlAXhVJiZQsyH
QvTjtJt/H95TKEk/I5Kr93ikNsqr/AVpo7ByqlxlF+Y8MXdeBodMZhcKrZqplJX8
b2pO5eAr2TjwJMt4idiQqHL9bMF1csSJO65aQRtlLIVAZVkuREnQAuSPr3+zdVI4
gILrxa6bPHasKnOWbh2ACLiLHAK49Qnj49zX/3kK65QDRtdf6yacnl9hemwrppyi
Jt7yQ/IFr3yQoFrOs+JZIGZM+JEtTp5SwKMiXtythWsZ7JPomWoQAYUzlie/9Y4c
yhV+1WqbwKKNJknpSP+1q+yDu0IYNDdGG50rXbZ1cTwvpnwMgnHtuhQv9xyrZ4Ku
yEfjzhAN3KefsMvwxkkL91ABS8QHN6YI4X+8/vePU66jwOzd4EIgIRfF2eyILUug
P0n9rw/sodKcvnCRF8Jz2c45zRr9Ph8V6koF1IOTZf4yadfIuIOhqEw6UmB/MZIL
/jDDqK7OH3QZqbtXHLgAs71jjhbGWAZw4kpGZ/30CDTjDiGqio4xJ8f36IhxLULu
BPcqdlqsjKBnAkZP3Mcjp6+jC4ICeLV1WFy9r9C1GWE/EJkUgGB9xhZPGl7daP2E
LyaosKJmUM6VgHqp80yfH0mGTaIGb47+A9n7lZ2u6yANoHD3GEa0Zgy1RDdSax8P
50xN/mKkVPXqcMA38YKhOFm+LseqWtKmSYKP+/q9mjWuDSxcjZp20Fod0nRqfBR0
O47fd/qijRwBYH1FniVLLyuObXV9EwEFWzKMtiBKgiPasqnwU3Bboj5IjHI4LXjN
Hnx7FpRmcyI+e8tKUpbzQnomcthZaMsGmim4jEe/JEEm11J6ey+P98WDDL0Ig1lx
rzlwjVaZcNq59BNtgWmpjLsPZgOOkQrl5Z5vf6QFbhQAdFx7dyEq8ZRdv65IfVRB
dXiDDDsMfjmpJiqT6cHQRHwfqdipS5JaWupeGDp7bJbldypPn8V5LEVKB7dr+K89
6ZLcxJv+28YOOEIdNCImpiBa5Oi0eCNBEgqMzg6XpBkhNcvy1UKeOpjQ630KLn5j
3InwRjkPPU6TMLH2aS/M5DfAxUf3t9jGKeI6VOc3+WgZrPRgpGv3UmziJWL3m8ju
1oVXK5B1QINZu06EN8HoM+QmP3yKnrAY7V2bOS3QWgY+4i6LZzpiPxIe9xhkYRJB
i6LK8C/ZLuubjuPDMTp7fdYi9vsvERs5preuiDwRW52zWxFwR5PIrod+YM1MuOwQ
hr/b47hls2lFpFyFArN9hSjJfejeW7qEwSMAdIZvNAGK8pV1lfoe2m0ksKl8jo95
gCZFTKH8ZLBZ/orlDFQdXRRIiNEC9v5wudaDCu4sGtcY9Z0O2Uqrvaf1bRgLoalK
8BBYuTdW6tFjz42NPvu2KJgx7nxr2q1mq1BZF7RgJr0o0QEjQhFcaUMwT/bnUWB1
SPKowe1zy+NE7CFq+9V/d9swPKYJ7tdQkxmoDGTBCrV7Q231QWSdv/lbk5dQ7Cv5
ZUbHEoWqrVtyQch9how3B2ePjx7fD824wOg25XJcddH9HrEcVVsosDgFyKMRaRYG
EdS3z+icElzIzUV3Q013LQ/udw/B1SQeyRzEe/zGxT30fNOO6rqrIl19hqQT6nl+
lCxHFxonIHqPrpq+oN9BmP+AQwfLG/oi8Iyv1DGYNlTczPeYgtja8BI12x29jUWc
LSV28M7F1k4QRx5C1uOrOB/OJ6FqrkuH4AlA+/c7hqq5DBAj2jQ0tDeuWW4pjjIV
gnkNoeXNmcmVCibyW4N6/ztsKYjHIFMnMQkTUhJ/zt+d0B7K/532Hu78ZiRA8RbH
ENJY9a0BQlUEwSM/rHD6tU8amw591zbJrEVhMjJ9IxuYCFFmW9Nz0l5q4SvOqAxM
ULb+eb7d6ofK1ISjaFyEgVBQvB59yCjqf1H6IhInoz0nVEDFQMvL8FwB/ksszKMn
NnK5Bp0p+X+GDjnEvCx+rwJ8JaMEQMyDuQ46PXn0NOUaDpPdIiqfBmbS1EqUbvr8
0kiMsSaO2VAUhLNr06p/T0Py95euBmnAKtPLyK6ZnG1uafI2mvZyQRBhTIKC+8K2
9eBZTtUxVj2zfIVvRgHVASYWd4eWOwLsZF5R4UY8f8txF9qej2xaESsIjPL8Fl7+
u8MGzb3VMMKR9Nq+vfRsHaqIelOWbIjjPoxGYtCwtQ/06/AEXIskATK2nKbXOD9A
1jUYGacmf+oRGZLrQsngCTtTEyVWRdDlsTI/EvRHoAH6lu+N8jbVvS5REDE7cE49
6an7t+ozU9ZI+gt8HpjIl4u0L6NgCQFKfm94+jh0LUxM31FwYq61bKUztl9uXlmv
KKzuEDS3G5FBGUq74X6OjnAWS7Ww+seDq9oGvGssrP8D3Ihnc0YR4h+GBWB2zVtR
ez1wIZjJzq6L16kWboCPrYh/LHgR00DfbhrODPUZC8TtIlUtUhLAAblDiDfBSPIu
tCbmHrShzYcmmt7ddCtLcYVK+b15W1VpHmQHAvFrqNwheXhOdAb7UJRWu5cf7nE6
An1OoQicVt4feB9b6HES812Hc/6jRVbVpIRQlBAPbTvyJn5+3EIFKDn1n1I3DjmI
Ev925j1RckimeOC4aZF7TOC268WSetdxo1kOjsIbAsAy+V7BhO7XQc1vD1u5Z5i7
sve4y5v5b9idxoNJjiGa4OFK4Ow9nKhgwlS4vCFYkkBK9KKN4mOd9/35eQyfN8F+
wR4OhbsZWOLd/Fg8JVtJWE45Jl4JvzUjFC8+x3Bmzo9WD7YDsEfiw3Hq/h5HHcil
Htak47+CIzxYMgYdnA8h7/WivvzivFBS/FAa5bOltQJtwLINyeJv5gN7nbkYF9UR
2/pIYAsOAZF0f6iyAjBhe65eoKIAJgIX1JlX2imo2iiGbV4mMi2hqSJGxsCjbirJ
7/38Zwd7m/V1BVCdgWUX2I46Nkd742FE6TYbSTUmvZYiJUWoqdgaJ8NiWnyrBT9r
d10lwuSaF6Z0lesAEcvHcC9FDSkRBWfmeEfDgtLQ7wgBqLUkdE3vRaXxNK35Zaxt
oCDoH5a183MQFBTJWlQXph5tPnpX7Hat3rZgituIcGeR00rn/QuRRclLiQGarOPu
NdYq33LC/efDVVdjEMV8ow0fhAPnTf1jpbnXYVkngXOGksMbUWxhjlzHUqShmHCK
6hc91pII4NY35p9EVptYFZvLZzY9Msq3MMQ3yVvwREY/WwjvK1Wcj1e9JvhyV1UO
ko1/fmLUdn7B/qs/vq9cmOGwWBwMHmbWlcPjnqjcB5YNy9ZgKYFkbeOr/zyqnwNc
/vXQAFcMmcoRx1uxbsl0ae/GgK3Rp5gPMLZDREzau8HJTXdIiFyU0O26rAEibdHg
wXQ36d6appGr4mhFxSLb4BFfEHKMgDl4LaqKfq0Vgalb/JnK4fbhYdxKAC89MQjl
fLwBNDtD7fQWeokQouyL/ceNye1D+xuBmOSwl6hsG9ohsFMYqMIgb4BwFwLxrrP3
9szNrd0nbBLC+icG8XxY8tqo4/h10aXOO+CMJ+W8uSoclCoPgJ9kQtrEmPX/iJt/
y0m36aZYEd805D/mGwLWAGsgZQa3s/P4Ik1+K/slu5M5ukZSAOPCoYg5TmwzIkgM
ZFeXjeq7ND0t/gidtchKwDOfeWuF3d/Lu8ohSDCVrn4EuvEwdfvh4tGErd/8iE8t
R841Do5K0wvWci6QhAJ9D+Vm68yDap9vVBF5emutjZwPdve/qlx/oeOPNXLhn26t
MC+QSOElduxw6VWUHm68QHsejSLbcH/DUaPwYWuKQCAY9Guxa6LTU1uMPlbSeZ9r
G19Nv9GT5tcshfXy7fv51/8zg+MnBw4G9GlCN5WrM4bkTiIcxt56DlOXTvWdBOFG
3zPsvungrY9X+w7+hxwAD9v5SN8Hp5fe8e2zHNrS7L668OkVbXpNEPqXiWBeJZQa
PglvKuPH9s07kBPLzde7o75KEo7wHKBHv5dINZ1a0A77pN1BJIsBONTzpIY9rP6F
tppncCoGZKxSdexK5+EsLgiZbV+T4g/LiucG/n5sgfrnXxipNdyeGPXihul6edFN
XUl6B19PJtFPpa7H/eglD+cc4lnoLhAmV55jQnfJUQAjlHO5kBSdLUnqJrm0xILV
iPvrQYssbW0s7b4S1vBNuJkiYFe3ErT/Cy4c1c1T+QZ5fMwt7jYRXTgOmL8g7GCj
RpElC9tlEMLIBFqhDvmkjl4A6HbrUxwUnhJqk9yHDrJ2WVRQNefRfkwC0zdJwV+g
B/StJyJTekpx39A5zaC2JYAmnpNQRL2xS1keylH2PwSclTxZo133vqSZ9IDA+3uy
vvxtRT/cyw1zGqqb8aByzc9gsGOg/V5xXRqpJnJhC69E5H3K25YBlAcTwlZeGqoI
XnGC66BNQkoGZIgQ7R8o+fmSRpTTxEl+zFmd69WXxgkqJ9EY2KazmzKIbdQsX8Bo
1aV1yI5N9i+rlHNqOCVU0jvE+5GBkliSoSxa9ath/T/xS1x8OuUbtw+WEjxSwrYX
E4Xb7FnhNv+6vHqudixzvyTmLMc5sqtyBp0bODKasByM5ImJXPFUgumHAkNZzZku
BDazfdJgIs32Iy0C/Gos4mTBm7X3ewFsgnzh8HTnViuHke9SkuSJVkG0l/QWFK/d
lrXd0uEMd24nsZxItkLv6MdB43Xud8xZRrX6J9oP05V0pvDUgrCkuPASon3iNuKq
EIyLI8yPb68SV3prUPdD5vVXFOGvVmDuoWZSWAvK7WFDrB5jVpF+qeeIInu/OX87
AxZBYkfno4njgcmf9OdTg11OfKl86vetqprOVRnx7N4ywhcjBoamF1+9cfkMSqY2
2Or0XtJ9WBRjmmqkDQKMxBDexAL5qzLGAm6pXY1v9RfBf7t4uLGHVI/8FEgMP+DM
9TiAxPTt60aKDtkv45teLRbalZzHZxYXIN8SWnHWG6s/KMtVopycjYS5C0cCutQz
UEP6iHNQUCqJTqn6tfMHY8GRH1spEnw7nOCCZuKG05UmmS8HPU0TsaREjN2VJG+F
GuHOicFTWv3Ux8EOQbyJ+d7X7SvUVCRfPfiT8bHG01ldbz6fdu8nfXZiROS5JVQn
X8AY29YTOqyQ0PKO2PTximtRbRoV0q4aIrblkl4mrDOUwnIKea5bLvCbZruXH7N1
EVMtgGxlZRJ9VNKXQ+e+47GambCar4iULmxkzvE6PriwkOrO66vgkVIID5L94xJF
pTvbWtu73Y3SEHAkHnRf6q5qJACHrWy8k3VMZw7lHbPYac2isb7RzOycMuvhn7xH
uk2Qa7S+3Hb/2iUgeL8obWCMq4xpcCHytw2EUiwbwy+vTtemZI53/Dlgaim5cvQm
8FEyWBdlDP/qlZui9x/j4BdXci1sZhpkczql3ncWD4xtaSgdmKtm2KWUHdl/3c2Z
m1ar+AS6vN95g00SucVgZgStD9EiLD6HeLVzxJS2jcGR9fUWbGpvHKKTqR+cX7t8
PB7OCd7cqfehb5UgRRXd9oNolnA9oIqfKplOKgg5QBeP3a78gaAHa2R8BWLmtxHe
6Dnjp07KllOql/aEhkyXqwiWQUv38mM7MKgvwwnuQiqxZFJUeOJFJKdXEApGsrPU
PZpt6HirQO3IRVc16Uq1j8XfTs6HQMCHnX9i58dXaqCiBL0w50ZFNl1I+lzyTDEM
wUM+uekezt8Nj1a5RH+iI+Jfg1Deso2sEXh6EvS5r5w1RjEkNrCxG1SIuv1F1enr
OitEwpgZZzXZRmd9rHStqSjCBeXYv8j4nYJ3Vkb3MmQyLg2mwRyaM1PyLCfjN4KQ
iY2xdA1L3gkduJRC5O9gVVvxpV4Y068ja30ld06tfhr1SqZAvauMXnBbuez4sErj
WCCPa1d0B71rBuiwN+BWJotb4mJfQR2rxDWTo/GQQZfuVl2JIc5Ozb+NJkI3QX/5
3pcUJCoejwTdcSRd4I6trvTfD1fFHYJld0XTtosnejHTrYOIv1RO9dPxSWn34O5v
uQX9YkQLDrtDUdAhLDXGoxdbni4ncbArQVQUo2MOAaTJPKaHEGl9ATFAm+7lNz2p
KFyDqU32w+06RAteqkgKZys3XjfS6gsbAJYnRzBUovmugFluRuYfSouzXZFMeoF9
D7Lm6risyD+l2vQ216ZHuBHevc8tfof9glUhAh9FjsGUYpF23ZXsZG1qdc6HaALN
nlOhgzj5PMXwfxp/j/28VM+tK7fiwFmXrGfntPTtA11iLdzq41zuikY5nQUtYPvO
jDifLw080cmwA5+4+3pkIoIWLv5IYpgp90Og9viaBexXq8q76PNZs+0u64jM3gj2
xYz1+0yj9khKCU9ifY649EK1/ZKyPubqdTYvqbFy+h3W+3lSRDBAwP0QrWyBnkuf
JRK36TrNWYZ5RfxLFFL9kR2Re+96u0eBQ2b9SiGefebtgzAtT4pVwlCMfWlI4rRD
giCWMTq+nI+sdjSoogDfsuAjsRDd383BMBgMpwKDbnEnaq953wCitCQSYxjWifpF
wgiBUZDqMkZuj34UZjGGEgsC9BdPo64Vmj+w/mptkReBPZqynu26XBYlTSjiigA/
Df+q1fcVS2ZqxFK01mYg5NXdkKPo5vNE/x/jIWnL+WC1v5D9ZHyWHJmtSEgl0KpC
NupdzkKUlEl/KQ7RUE9R7QCo/spRp9WqW5OaefdZ1nmsqokZuRETtx0TrM6C/Bfu
taXWna+RF1dD7/OLRWTdJKeS/LKlxPpNu6jN2T7UaXna31hbvfaBwspIUF9rlDCM
/ZCMfqxYJnoRR9sljz8HRdKjOb7mkfRNGYMVTXZisaYzgUsG3u40GP1gRtkpVF4E
1ztgxBeTro9SSA4FWvVDNWB7PbaTMLmEXANiutVPEcJNr/FEHuyMJALesxtyqxtU
3MygQoxxXmYMMLjxTpH5XzJ4l3BicLaVSgqh6sNgHXI6DdFeoMka4KyhZ4UWTUYb
xyNcMnuvDGxthpY+PfbjDeC6SRjE7de0HL8mr/gCea21LsQQ48dwNJbkW63BqSX9
GdHqe0s3y+nbwvHmmmTQbLOlSEPBDY4MZGKx/lAhQ6+L6qjc0iRQdT8/OQF7P6x+
ckIOpCi/2D/P7FmVIORU9FBPaz+EoG2VfFZNfbfl1QD4/icltSaWgm0VWq9AcZ6V
/cIcbMNFv761YLPDSjSuFFRb4fDx83aHiJcQIRSb2rqZkUgiCYFiv8yjkxKBKaB/
5dlzQwgj8rcScmsOjkN9/0tQ8egx6bov+HKnyB/F7Wx538luyramDYORMoygaDuz
QGIcKNanc/38l52dyluuLnBk5eET8V36W721RcTaFmATw855wrKy/UU+7nfh2aKA
PrCKCQ98BdCZGnHQZ4SVm3D8lJXdnyn+4LHzK/sRjlR/uPYyxW7goi72QrJ6Sfh0
TUhvjNL2m4sf1uevgTagzMySI1qpIS7M5/Y1fkB9CheA7MsGBI0nFeW6dtPhZ8Xr
N8phUjpx79Avx7dq4GOJqxp4c1R8aFsZ/RUhHaWuWMARXl2svzkvpxu408DBh37j
/WpUpN+rhGf5/r4rxn8yeJO+cvl0z3kLPgweDYbWEpJ7BiSx2/zawQUdoe3nK0Fp
usufNx04oTIBRQw5rwJNFriBc0xHLb6Xq+6yvcXfANq+9hzR7MgDtseC3mXT9eHQ
dxJbidkQdU3N+0WpLrwiTZAGfb2H9YC3vRpB0KORidv7ZXe7V/OqcxPAfnbGwjPr
uCZKOal9z3UR9clwh9gIBIEJtPXt65MTo8D01XaxPoYJcICE8HN/J/non8cmlwHh
ZggzqYQJD+EjiHut4Q9+nQRKXkZxhHJnU+6IQKpg4t7NHpQZF3e554U6bDncSxda
sBNyJk2Zs2dCN31knrqVb+t8CRZ0QAhrO5rQVCYhUAJyupqV8Vbt5rpW4TgSXi3T
rKuq0iXMNektKv1nNJ6BkJUfaP5I1GClDhEz4T3oE/3fljgQwkXzCUms67vovpVz
az7/ti3JASKT+g3hgwQNuaKFSJ+6kHzIxVbzhleuNGsuzk9GOlZk95eGZx8uJp7W
ATt9D0FIgQH0s4U4/MTHsyncY2zgfmkj6B60d7rBzpbTB2EXIR7t56n7jI1+2p1P
Ekq04HaMsGCT2jG9NJHl9wHQYVW4eh2/kPP4Eg0yu1f+QBffeP3tXJJDAx092rJE
WFKRNJcuNGyzr/B1hNCLOUhYWrXVILm0UClgtZpETOnvPr2B3ymCYl/AHA4tUioz
8vZ+G8MGaurelf+DqtJgV7UU2Hol3uRqg96MaORx2iYJBJlbrIMuLQgNf1E92WWF
7cA6O3eDVfsAdqi241wVET4GrUS51QM+xH+xeljRkF2syxNJTkmc1fRDzr6dbl6J
bchJnF4rraiWsStkTQ2xzgVytRUw6whMxUpdfeIxDsL5loc2ldqLUcNr43dmPqNE
eYeJ2CcbtndXUUL1gZMciiAXE/N90Ckp6r0GhlIeuCexoCI6TT5YIRKI3QsTLeUD
uaYuRddErrl/8H1pqngfzaaZOOI6UfoZcJIFKTzcaKDDRWzc57vfqDzJfFNBaUEK
7Rj0PQW/4Wnxy2iTmX7zs+uGE1Jws/0toUbYcle3ghg4T/9O0Toia3uuT2g3i5CE
b+M73eaYQVn7skrJNFks5dKsvasbdxMLVy/rZlHlSDpElMHekiuNAZG/0In+stx7
Rm6zX+yT2VehXhCWjGdMpoLxZ0lBPIFPOgGvksUbq9fclruHETIadGY85ktdovdn
vEKjUP/fknIBPJrPj7PM8wM5d7+jrCvTa69iPdMF12ZwBKgQtP8DTMG2NCP2nY6Y
wOmnDBOQ5IJ7Ya94UoytHsjO8RC2u2nkRbrjbQcKHmjpFQ4/iHfodCw9NYSvBUrz
iAHxSPAIhE26mO+TOlRAyon2UXebDVViiKWDUUrzLPSgcDfm0XofGHqjsR8brNUW
e81QlIwt/m7HfzY03NzJLKqNoYhu+e3Du/g9M+FryxZnZfnwUS8pQuyQ6/yE/AiT
QDgsY490zikkaXZMTpr1nOtLXYm83Em9+AMMv31WfABIOO6yjYgRC8oE5nhnnqQJ
gysAzQlOMh308ySfCI1rOqTTxLHhT/OO/H8EyhUcBepok2CaMun5codgQj3ttEvN
DI5I2DF1IvqxcgjDt1OiPN1KirG4C4/jpiSc9t8986YbVlL4I0DLStby8A0VOSdr
KF5C3Px8ZTOoVoRI0HVDlDNbRRdF27qNaB7digu/DgtrJZOyB/ETu9Nhilb7AsMR
ZhaMJgf3unCNhU15fq0TXvbJdCfFif/i6WJDGRuwQgoXUiOTWuZ6IqxUL931WIi7
4ARtqI18IWaPtgUN+XLpp9gqzELZYaYrTY3as09tbdj+KsbXuQcZmzreVmewftRi
+uRQfY+Zq3yaSLZgE6AQEDCIuO4Npj9T+rSIMts33hZYH150iSaCjgx5eglNrraq
0+ghlcDYBkFQiXndqlNIdTF4Mcd0UZCLeGzG7gkLCS33owfLGZ88tF3uPeX9XOYZ
TsDaNwRHRs/I6lIWYCT5ypAWMqlTr2NnEJvTuiFIApIQkUZWY8GvB/I5OFDU0EnJ
lm4yxPVeq/l6ozOx2OqrZIloyeBw64uCn+5gG0ZiuSGqtKbD28efLZ/K9G9dtEds
ZVWl8p4bDy+inAx7hQQBUunHwzRA+oLyICEowV/Jgrvi0QuaViKdKjhYy2dAwaFY
xzHra7dQzVU0SmFhr53R29lDwbfyNlkKALYLamv/TZo54KOiRSgXlj3nZSvAliJx
ND7KRchU0nm8Vi2wk3+JLvZFmVAHT3rtcGJeW/JdKg9VDPvxdPlvy7IvPIwMbwRi
DNNCBfZ8tLzojrjQHyuRgk8OnajK3dBKKNpz9QE3MLvLt61MxubSlWMCgVUXobqF
RkdFdqrkgmooegA6BFSm/ERuHisCYIHh21jTGKK/2cPd53fuwn74TITfGQa+N0s4
X6I73DORwcDfmHl4FYZrG2dkVP8cQHKnE/yJn8TDqCtDcQK8j7gIzn+ZWU00aLmW
NDX366WuBYF1JwN9BZHHgM2b5tMNnxCJhHFMzV36aeUTFXoNxTIrb0Czdt4wteuh
qcFUjrF20Kh3gm3X7HWIlLcgplm3hH2fUKbpfllGCXttyC9CqEb2QvCmecfQbhNj
EHZFeSrp4weRH9K9D2AC44sFgQU5LGfsEjWIVU3/u1h53aWV2OMEuZQYMW9PFm3U
aXD9KLgVC7xSjlkepNrtWAnaEk0LOY5EwDw22kcnmVSsPwLCAm0mlR48szpJbnB9
fhKGon1+EYPqFdNqFlh/X7IGisNu2w5UJOx7qbmAgbElB+jPKmthN6n8gAlRwue6
vn6OaxnjFaWA8bViwoWrJJnsFJwKXYaaZHDJcrtJ29drKC5bSVtSufx5MHGQxcLP
Xy58pzWSSEv2G+0a1BNt4QaPjQOa/z+Lc7jAK8JHnEnHHrdqeZdppf3+pdc/scJ8
liL7jrW5GUITW58kH9vu1DGO6i1im+tV1kVsN6JOLczn4uq3EICignHH9g+UOEgb
263MclNDAxGTb7ZtILnrqBGE30BI7v8xyCfbLxceEjNhyyDNqKgLicy4ETREjjfi
JG1HhztKeNJGyTVVqNB6LwHgAGU2xQI97JpX/Sf6HwqKvYmcPROPtVtBCvReHXnT
DvZh0uAOfeVfqB56Ud3cVNZcC5Omx7PyoEw3sV5zI8QaGM3nYIH6pgWb2CjInRua
XVigA/PuZHyoqp1fHLIYQtJlllSUyOeqFSazbHQu/wmxmut82FrIHNflLUjelLvV
vHkYv+uLBuddNdbYdZH4nHcD1RvXqQje15H8JXf/AYpYcVEn8u9iCHFHekmCuQGm
gMLNefYmg5n5+QkPzrOmx9fQVlVnU7p+edcm7acsxAi3QrN24LZWywVOOyhrgWrG
2lj0pwN6C6sjbLUbYamRcOLi3+2JICg2rxL/QyGuMw2OTnJ5rnswb3w36CayErNi
amqIvg0pW1w1gSNVFuZeUJDlWuZNoI/pvNVHZLZ5cLe4PgqW3CDLozm4LTlfi/fr
FHqv9cJIfCGQZ5CHtpQ3GvYCyPTt2XHAixyphLNCyIZJ/Ik/iUwf9lQ5FI3QJ4en
hzYmOUXHtB6emgmC+vtesTehWAMSGRhCl9MguZOGOhaPQkH7WXUkTwZjUW8DDPeo
CbnRQskPp25a7lvp3PX5goaQSORIAT1bKCvCvdTwGH59L8+wQismDtfY3iUOG/yn
tJSPB8s9TP528gS6I4wcM3+XPI2xDgqG1FqnVqTbpXH8wPFGEDMQcxYZtq4O+jKZ
yDjDfnqRYNXfOHiCmlexjrrdoqhN+EOrldjitvvY1PfJkDrMvXlnuEpCtY6Ceduw
uhPwv/JNDXpDOc4rZ+9EvF6i26niHQiXt5qBCyRW0AtxKxXQJiKIE44kizKO3jgu
tI6Rh3AG+d9120PgrjpSRBWthh44nPHIVft6rHhpkcetLjg6v5MKyR4PludbgbN9
u2OR4BSLpPwOp/AAYNqY5BzKHL6gTwA24vFCMZG8oJkVUzutYDpVIh3OTA5yldUZ
6UPxcR6SNhW7s2aIBbLGOWthYevV6ZHC5P4s7fZjHFgSUZTs73eofb/N5MNYdEm3
Wst6VTlLjScaGOYHYGY02sNtYi7gsyij0A9SHh/PuVOeMIJO6BZY4oE3iuAAgSWs
DSQq7t9jDLwpdptnra8327jfebPTv7xkG7f9ivFidMjX65KyYdLyn+l6Z0EdnJwK
DU/ELk96+FDpmnnEZ2D+HKIu/D31OGze3LeXzpujpqZnQxpfnKte5AieO7XsPlYY
cvZjxDR0NcdXJ3WDtVQ8JywaMCbDf+T7Wsb+9kyiDJKtxwhIZuupb0cRj4kYSmGX
vfmlTzdJyOqJ7YjRSe54dlQFsKJRT4K+x/ZM0c4K7tLsVSQanDEMGpSHWDZIDA8d
MhuqkA04gTey2QhVVzSKhrqqm+LYnEChjVz829ceovsIP9TjmBWqk2g3sChG4iVx
mxJ2/vLuMvlvNbHE+7Qew6yp+jVdw8hF9SiMBON7HyMJQZP3BS5nc6sZds81exf6
OlGE1VYNSEzJznO29u448U3k8F9ctF9FqMM2vJMlSkgYyGxAZrg2T4e9ANdTW2Dm
fH+cKw+8QLwwMi0iHWT9dpuq7eOZXFNbrCFf6YLnzyWlfP2EYgQIG4lo8BZ83IFP
DFTDjcvHzE25H6th9Ve7PsVcG+Db4658YoAGNNDRm/18i2WdJ+5AnejLuQtpwo2P
cBwaKCbW7wAWe+WhgM8h2mrQyseJpZoL8uOd1ocZr0wtbjfvr5yTRGYe7Nl4PjUR
kN6aY40Hl+EK81og+QMVPKu2knLIuHHaQIm6jlSYeyhypyzC8kjdjlSftdZK/Q6l
3JFH1pJ/lfgwH7GgB7xZoqQF7TynvSBIN2p6u8mpvHMUy4Zddx9GWROl4mYSNmLo
5poYHHOStIGLbDsBRJAii1b4AJYASW76GSISijpQ3eOQaoXHxrxU8tVJLjm3eRiW
zVDlUXvVOkOAj085e3baXkpZ5M8cl9PDvBQMUzE9BrNm1JzKXMpZRwfWQ7E4Kdnp
rL3x6GCcfmoSUZqDqyO1tKRC52DeFC7ZVIgP0AcHj999X0ALM8u1d68VQl1ttmHd
lh5qvGe4AQixEG9Zv0Se87J50gKfpUADBhCOL6GIB1VLY3f4YdREJ87BuRdm8sTU
WtaSAXXh+/PH8SQY4zMdMvFqKo23/PyYEJ2AIdMaYcLnLaRJdWse4V3nYmpbBwwy
saX+WcQjieZhqOAIeY1glNlaejWBEUoqan5PeJAl+wPaEx6kgxNWxN9SsgdiCbuz
IowPOmUzMN/Fsfg0iLHhh4G6Ce04RBpv22rnRWtd+gzlmfBjeD0GlNrFQEDU3lVh
DQURQ28N2j3DrX28LdiAgXYsE7eE47NEu2Ex6lX9NmfIz9hlkqED3KcbNRFoiUSB
F9WZeC8VnItvIoK0oKYSS5bCwxPkQvrNLv5M9Jy28OP54prG9jLhDdfhxqunag9b
ybW1r/Xh75wW2lW/QcGVHv5SxH9Zf5vluZi/z4IFcUew1fCF5nY5j0NFL5U4GgUJ
yXbZIk8CwhBrbPNQmygREps4aeOf3U6Slhe4jp6Grr2JS5o7+lBTEOH/r0gHp5NS
QIAzesOf1gMXGuwdj7lybz8kHfSYTLCdE6yczZ6sFYvT/GaxuULM5q11tPxfoiK9
TL8FJjqUZuxgTnFfiALW5bJjUoXEAr9Lmyabdhy+SGuSrTO+KIqTM7Yl0n/YvhIS
kZs8MJ4YvVeg2wLeoN+DFQILbS5zGxLxf2ZLry7ewTndAaAxwwKbCq0oP3f2E1Os
hv1PLEYd/tKISQ9OO1fHCxxbpCpdYUZ6Jh4QpoILWXAvexnwrE8wPSrrTki4Xd57
gmxbQK7BCchtCjQAKhXEDF8/iWp44HyYbP8flc4HeDI4cQZXgs6MKDX9qZ73ubPs
iPp+KIR8AvILfy7g/C2TcIGJhf/836ce2EhJ+WmAFQBEYHZ/g/9w8JtCRHycAydm
ly2BLN0Wz++fX7kj0frBaSSGxj9JlSmOi/29gJEoPq/ZzWNRq7sAlElq7HDNYeSp
hxqwOMpYBetI1AP83Kv+d87lTZpzxYOCisJwJPl6EsF/rYjlS/F/R/RT5j3iQ4Cb
j0urKPNO4jiolPY5Aqd0EMR01QnJCBUNknjgoo2CeJhsD+uLAZJ3NjCiVKcMRRU5
KBP37+DTfmGkj5LNr2+Zqty2fHTWoFEtclJE4Xajv7vHgXRJtb1VhR7UC+WCUBxB
RDgg1WaYjZwgDwJGwrRQBU5JJq1pbA2sBBBnFAg9baGh24s07coTxevBeofRWNSb
dNtkvDpCyQ98JKmYwFZzXGATwGgigcYOeMIXaR3FsOPJ/ScYdUx1rN8AoPvYuxiB
JrXf6EqVaeKjNKUFVm01miWl7hm8WvBPh5YinwYumgU/T6x+WtuBXQRG7S1rDglo
VitG2trbSnSjemEyB44eLZBFkD3RdPzQ3ceXLXwM6uxCAhXjzeQi1eM+KW6s2nH/
o4NCklDGb7+6EaNCqH2W0meEBpu0wyxRIkd1YVDIKlFRTThe7umwthiWY5tbJ5m+
aupfDOb/Rjzy07gpJc6d5LEmL3CEhpxa2W9LJ0kMaxX5UAhthfJIceKGiRKNyLmr
ezAbQQdxzFtYik01ERnz2MgEnddjmnRm4hMo6eclyWiucfWFXv0qvrSpV0ZbACOl
zNyjsnOSRLEIMPr+fwyMj4kfod1HodBajeVHK7z+YKUVP9BIH5U4WluH7aMjeU8p
jR0/nOLzAHDpCoTq2BXBoyJbgQG1NebFL3w2okjF7nkq7eazuCT+ycBy+eobb54A
a4pBhHNa9eeTyE9xP6DmlfcuQQWVQ8fR2WNVvXW+kI3i935ZR7kuC+46bWXGRAzN
nTytMsbQ0rscE6spr1m4pOASbTp7J2skW2osLAqehhY5w71G+4mK1swYXRZpSpq9
q9AleVmsYPAk2iesg8EYmJeQ+n1UEZifahbBHhOsQNKCtux9tUS1jKN9dIkXEJD7
TddCo9xygH9X3y8C1gcl+YgV/K++mw0IxsxnCtVstXF74fq7MZnLumjYvu3ZHSRf
fP9zXmgzDbgWLHhX8Ubm3x+0m908JzX9hxtlByiMLZfT0CW/yiL7/9XcKVFeI+cK
QbIL+hyDoxOlY158fN/qJvP40W9SY7HUAIrCt9ZuNmX3GNr3Yvfj0GZbgOgnKkno
KtCnWRBwnLgvmjM7ySpYe7+KkJh8efj1NFnKDDJhG3A0nmMAlTW7CUOmNvElom5f
mjAbHzWWB+bUXRoqsJyEiepIz5gmhUsuGKDmrqinGhN0qTPET7Plq5bPeDZE83EI
lOpECMEpcLNveSfS9UYC5whksOcDz11GpveNBzKrv9eiBEvflZGkC7ecr0ryqcuS
EjABZODXWxUBBXKngxJNyfe74AR4ZEapYdQnW2FsnIH00I0W7ixTt3ZgvApEW8Fm
SB6E+I4h4MkMSWay9WJbwtlTeuyFg4yClo0ebAbGx+KiGbt56tVQikDGCqgx1TAC
p7xRQ0v0dQi3YZxDr6J8kPXYsJSMqIca7likG0v3n6V6LOCrCF5p7nWoN7lOGolV
smtdXyt1akz8WKnASm+V3tLijBs9o+y6DeTZgTyg5ZaYOjjRYhigB3pkBrgcyh+a
csyMpSqXuE8A5AUNKK9orYJcSMlqybZ0OtAxSTer84J0gVbLXp+cYCAza+W+YQmU
vKIYt9r/epo39TjTFnAevAmwzNSzqw945HOQb4Eaq+q5JF3mQCN4EtvDWMcmBY+A
fBq8RcRbV/gsVXlVxvZu9+PulgEkGi8yX0448cfTsad7iN8zKR4GkS1oaT0yQcjK
5vt2mTm/H5cy8MDQjIXeSlkMvv5ELs9ZpHQ+S1LKC+Lmh1CFCV+rR8lIkftyaGgV
mH4oSjO/3oSN41p/qI1SWUbfZSGvoSGxfrpOcFal5mKrmsD7F2AcR7TlOvPkwT/Q
OviRFHjEBNCTo4Z1PH1lcXBqqt7ZcVxuFfUCa22xmgeCNyTRc+1T4reCIO2PstXB
IjkLuGEmWxlxg3mc9nZTU44KutRAS5BZhiVS8c0qryjrSTPPHYt0PPXl4mdv4y6k
qvyvpIdAPyClzrCMfIOGLFsILrMT76J+xrfjnbRmTHkuXPkjmZ7R/zDzVCeJvU39
0a+wzSGNHTJMGLCk1+wXNH8HwZunJ9USJMbO2M0MxNu0ElAeUWdyNmKGmfD73nKk
uQME2zZwvmIQgVxHXAOhb9QB88j2d8mpWw/u+fSTGFv4wwIgvIRzOuLE2KZpjZEv
GZCklz9TYAppSV9nDBX64HQ9O0me9fjihS9AvGWkIKcCCccMLodDnATwyJPrhaLy
sACRrVYimjI2cAO7JPCIr+3FSFtfs5M960Yksb0ANTgYkwE20Mn/5Z39w47iemSz
GSdQQFKgyZfZHdYk7DdM6zJoZ7r2XYj9DvRnBLQLfNk+jrWHJIwRtdRKSK1jKRbI
wRAPab3o9y4iiJLci/IJ5fLWbpy3FWusbNXFbIVMEPU5ncA4AfvQJsWHmVUgLA27
cb4pNTtYPm3oNclGqhL9WVICLtaHBgmErdE9cQe9PZcE7yDOVXMQJergGt6Lgouf
2JeRKJyOsgPJq99fp731YMqp558l9iz/HfWbIsNX5E29kE5O5ro/zGkVy6Bb3viB
fTTe24FHqHCyst3tAfnNyOML2c7wC0jfq0msCMPvyPAsLk+xpqKbkH4rWPMmvM0x
nlFmrqxIwATFzoJzsEX1qvKl/J6w9QVdqhDHZ7uwwUklviyXI8LKZme/cfWE/8vn
nnmajWg0YfKNC8yZElP2+3HBi7tlqzeDyXl4iFXeTX7PXk4LnqTOR9SUIpCSIKsn
KdzRvLOn8UeFzVR3E3KNEOxoeVz/m/IbOCweWcR/RiKXKQ9DAX+0gLwcplXg1nwY
lPiBnKYbpMunpEoV944bjh5BY3CWfEnSlXQHrfSbz3r/heQaFgE682kbnD91Gk97
WLWj98CCAarIcKAr1YnNY8xo5i4v77wguSur0d8Lg62Z8cvmMe88XYsnImFLSL/V
tLhMJ81QH/v+S/aJ2W53YPLy8oOx6nma9T9v4yQzC1UdcQsQ2VDNJ2kqwYLxSgSE
k81YVRXsggcd6ZQ6NoPZ9qHmbmKg5cMc6rjhCchO0TVdTCVjAPNYexxF6fLOksSQ
6qOYtvgOMMBfebMPfhtrzZJjLTeVPWOY77gZyroV9EYW+gNntaCq1T6MGb+uqSoW
HLcqVE39PALBAHrO4M9+L9SflU3dBL2pgu5aQHY6ulLUfzSSWLFDKuXaWphr09AY
LhPEpKNGMQqESDvDDWqTiL7qvGwbQA+LEY5kMG3gUVEWlIMYgsT0wKncODAmT+kJ
H0nJZBE1i2X3rrB9/1UC32wc4gB8RtKFbWbLKy8CfMa2eGJY9wEdnYBNhojq2Y5k
bR74MPa5K8fLfL+/YZbIdOSxVPhKu2dUAcqh7soYc+pbSenWYlu2WVIHY0XV3Qhx
4C7eYZElRXVO2+UpMS/igXnxtPUu+wMKyaXjWoTaDJPrL72gKBEBb/J/RIKg96uZ
ovhPIIQ1lEMWkz7j3GOFIWB8OoSxfnZZhgeADoiPM5Q2dctr0ge5eidbghDxCT9p
DU23gNZZjoX7B3MwHWnNszi+ZGz0KoJpu5bJUzAQcNwOdOfYxAq6k52HVjU1Hho5
zChTgXCgm+ZsuppDQUY6XkV+H0aJZQ/vqFdTWSbJPJ4X4THlJkPeMndJMN7qvqDV
BbCGbRSaRhEBBZhS2Eq3/f4OiXsggYPaQPiw0FvzIQDRNLdwqvzd/cwoazEt+ejd
2f6is9cQsGqEphdpRX2VIhtATjp3NyqpNP1KX2sR8uNrUcACUa4hb/cmr+TZ2fap
K8AII18eTCKo0pf8SAiQrmglqznfrF5kEuOffwVabzODAkdfY/zI0RFiGZ/qiB46
gKVcKrYxkCFtdK1XrxkA/iotGoq5OzDA2nyUoGXKZ33T3bi7ttDowm5eqBAlmVcg
HBQoFrX/xIRlqv2hqXebiNX4snvjVi2yqsya4AWVKJRq7Z5QjKVGm9eR78MJlBGR
ePJvUPXYLG2kXwsQK3F5DRknVDFhamEyTu3LzGPoiM++sA+tX6ifj2D+80U8mucV
9Tn9DoZx+JLFgzSXUAnYM4mPsHVJfiKYJ6w7faeh/F3cU+G4bxgQOZJ+EPnNlUAC
8WTk7KlfbngpX/DEwwfiM683OPcdqyn584PkxM6vN3YEBSUvHqszY4Wrn6Sk24u2
IcnXvp0vgEoB0V4GSgs/bZP2mnDavV1QJUQU8lVqFfAjcvF4mqPJPIz7MJE0ddp6
23tDJ77vqwyAhIElIidK4hiWRYUZZgXIE0S7h5tOqI2CEIzS6O1Oij7ItzRnK5hX
JM+H7Jbg8NNM/Q7zEDpnmWCNqWt6ZMyjCTO5z7a27XUuswod80Vnb6n5Qgdc3bLg
6GxkRE7wTxaXJ6vjtm7b6dDXyuDBaN9HIVNH+JUdDqif/8DVrUXFTr9Mi1woQBqN
VBxbmkkgswvImBdKbm1Yf+mhCIag7Q+1RKmTE1nipWEF7ObszZbfnY2mE56a4q7A
rzBLEmp/9NbjOJmNFSlC1tmq3s3jqLCVifTIrK6t1qtQF6ga3FP2WR1vIASu47Va
s0YwFsAcDQvOfnzEaCFcjyXpkSyAUFB/5qvUeOertYVW+JWu1xVOjrxzltJyNzg9
h/blANDQLiwaNWd4yQCLLgz+UN9NK7c3TtmfpSNUzKTXg3jD2vfv4IGeaPfqfzVo
MGTOsvmugaxLN1A5aS2U9L2Gl1+hga/xuZcMoPpRQFMXR6kuBAswYptZDhE0IPda
46qkuQH8XZ4K4p3xSc9H/AXOHT6+sofCKtBmhZya+DiFiDbAz6ylyem6lqlJwcqm
Yv/5HY7zRDLMXrJAFRvTzM6QINv2WmSIkwNg0dzjUcH1vtsJmQHImYK0PfhtWcCp
rcdo6KeihAOKmcahV0mCvwZd9Vd1wCselxa69Tyy4SUP3fPXEb1/d0s5s9VJqn8I
ypl8AGGraw4Tf/6dnijTyYqVcgasnigK4zH2mvkVZ7U9PN5S0axrQgaL/QT72Wxs
pexYyPlqKcg0nMIhqaZg7CMFiPeNK+6tdkNvSV6TIb1qTwfpGO+HvWzQW345fZg6
OPOcS43jiABz3cOt43/xZXT+nvg0CYsWAcr2znHMjkVOJb6gB4LRCH/FyRkqrr2S
tGOHM/WJu/4GpvBsik5Rx3EG3lxKZj4BmExBM+H2DN/YOfxxEYIzSr+RLKTczzhr
ADSWu/MVSsW7Es3XUgcN91gUx9yI1DlVuebf7Lp/yaNN7mowNM70CmcBHri8dmcf
Yn5Zya8xizvsobZ+5oaI/J+AR8BuhtSF1m9jHF0Nferi5UhrkPGjz4xHBXJgHRKh
3mAE3C63oxvUJo5kZzI36Y7ZxqvJSvL6yOyFeSvAji2ixO4cxKxu8XBt9voQu/qa
Drnd0A9ehJ9dJaeuGYivVySDeNy9U9Ssfi4IdnETcrR72q/jaVxGOtc37C/0eOKp
jGJK0wjt1EveAbaLBZnGkSiZspIazgzPnPUBjEzG0SKWu6mjNG0++r9GEeZig1oC
t0uQqFtatXSLbcf+K48ScABBqddxaWeTihO4ILpPs0VVS2W06okc8l25u0oV5zwt
9oowaG0wWI2ztgJ4RsnNZ8aW3dwFViAewPSXaTyuFGNn+pmMF+VSLg4d0Fy8Yjn1
h8lsSc5/HFe4jWPoOuDStXkgjLk5tviIfc0BtKZ3jpunMQldr/I5czQ/lPCRza6o
EtL9YlCe6dZ0ahFnov3nhELTHXqfRJGZENg4aT0IJxZYFd3apUfbJZpFYWTm2qoQ
TFdS8wG6zAfcOv9QtkavT6q6HR3u3movMvUn1w1TuLM12GMlOdKiK+xWJFC49hBs
Zgjj2+u+xivsK/P1kxVBs6pqHVV+zm3b5sUVWyqU9ifo3AUA/oBfrawSTGarqEbg
yPUjJI4nyJeS7VosX0NF6r1YNoIWDzWvkz3q1kW01FP35raP9RGETBsCIWA304kp
ylecLHg+HdCXd/pPzjxWl7VmQNo/pKd6JtCY1JcOVCVby7heatBJQwdLc41vjGQZ
XSxtHLwz0tNzgSVDLIrcTQeZH2yJaB0vsiNf1ZtQlztfEcwTa6zbOYsxv0uq/gH+
0GgwpvmEUB6SWeVDLBlRWjzc96KPlXGC/WIYoNLy2JKn3SmyGlpXZiV7rUYs7r/Y
Yyo5j/wRuZvB0g6XoWqMG8+jm/fefcJX6PtcVZEK4/RE4dgX/OyAN27DIIPFgrrb
YlvVbqB15mVe8l+39S7i6qhul5kyQoLRX4grb/pAYkUMtLicPrIo6pyLxQ73FwYC
3l0GUCKFMrAyWdmNnXuTNvF/zMITJ7Bwar2PUB2uWFvGpEwXgxa36jDKTL8CX/DL
A5AZ7ax7ySaZ/UnE4KZHStko1289u/V857ycAs4/oFqV9CtuHyqlALzp+4qKfiU6
be843/ntzTgho8tSzN6KLOU30XYNL867/qztUIQULIGSHEbOcZ6johnkDq0Iol25
4CQC76U9o/3Odsn9cDhQ37IO9DB7p9zRasEf0Y7QSVRoAjp4gYlZQltCF4EN1GO1
2JS15GxDf4idwKzW3t9dpm/zW4H28RnZHJDwO5UhV1YFid4GYyXvk2huMmQKk3gZ
lIKgwpAU533NSNkfkSsld9szdVBxs7NRbWskkm4w8gPEzbZcPgb2xcrKo1d8Ue7I
Uw7slAuemBai4whZfPKr0pMlrHmPmGaYFlpa0GnWEejW1B2YroV/exGK2nDH+yMG
sy0hJiSZhJwXy0vHV0b5wB9ekKUG/umh5gwaGleUcJWoE0NIL0e8X8wJTHa5f3BF
pJZ6hDXHoTPIuxj1LRYijmliNwLx08+sF3csqbUQKslQZ2Ab1kB7m1ygaUEebd2s
RqHsN9YLVwdPLQJAEhgqurZqzcEfeyYC9yOthwpRK/9C3EhYCTqqfkCwJiDh2Vq6
kuCMqIaH13462OXa00QTRICWK7HOpKiaPOxQ6HPMOWVIOAhgC6WxAomUzETWw1HN
nY7bjWFQtDwZqibPUT7zMbty5dNh6PyDyf/YJJTTLk2xznHQoIZBnROS6mhCVVci
4h1oIw2lT6PZsaFvmCiRidsJR5JP4Q2+aZIJt9BXPEA7KsQFzV5fmDAdgv3NjIEo
H9Aa0Jba+bEh4Q6rrmECUhD3c8ZLCoXY+zUA4n/fXDT6VCy7q4+jTVt9OIdUm0PG
FSlMoKxRWEzH7fxvyW+v2AltHMbuxGtsiR6a9WuvUJ3/CNWqj61w0fMlUiLK8eFh
cw0rCsWY8NzQNwv336fxGuezg0S0Q4aKNgkC5R6em5W3AvJ+04LgqpzivUpEeb23
+6pMFLTlXqWFTI8pDhQDoNjPHvjFa5h5rJYjU3XEgwfTIaTHS7vQCDM8dNg9XSYK
kbQpB0Q2XAcZUcsa/9/HhK+s1MUfIyqa973Yo5OzhbBMf/2iTHi1YIkZIO8Zy/dB
atfIpBJrL/Xwa+r/vjayIjOUyzrJzngmeTQY+02mz+w4hvahu6oKWExac2VGwdci
G9eT6rfxh0uJ/PltA/cSSuqr4u5xhhIcw5DWBGHuPOpQZWhvskNz/8cvjQ7Pe58K
Dy44TZW+wDpvswU+68s8C+gnOHbMlk/OEOXSccFd9X5rm+dmxhbavyW18JW6YQnq
rwaDh5ZritYZ9IE/cmriVCh/RWC3yy3XK/EnXU/aIRa6rWigR5unzOljMtAqrC1D
vqyswoMTLCdZ0pH+Et+FxVtIrw9WTMBgVkSj/o9mXQkXdAlo19Ms+de4ZLl+vnCr
/jMlr7BraTagA/FXuIgmx1g1/bNssFJDmNRTwPpprsRHqh+E10PMrsm2ak8hiDN1
3kuThuxsnuuR+R06zX9eTKuFp74HmQmVGizRH17C/GiXqSdjTCbQyhMBcK93pTJH
7rDbjXoghpPVQpm7Viry89nOwxNn00futayLsFwjAhxKZUHhwFQDkFyDfl8vfaZq
NfZFsZaF1O0Zm4+hYYcyMBQTYZuRGQjcYIm1Z6P4z+h7x2u20gr8kc7Z6TfNnaUc
VRnVFTmT+KEZ7YFSyApAYsDnk//ok0ohQCgQX/wv/DU+Wo7na1S/iYlrcBkNmkNE
xv2AX8FuIPHvxTEDAvzGiAR4MvmKrTk5GwDiaNlG7tv6ZTpv/1CrFdQP14G4Gjq1
RWmwujznyhifTGyUL4p7W/q5VQ6nNWavv+V25y7dn2GjYl0e+Ijc/NQceUtAdFDv
dCscRyWwYfkBa54P9R9OiuB48EyQ0YUHar6GhvLlIbBB2E7r/gHGUw1xj61S5Cyd
UBauc3p7RuokhwMLKq+BYy2QpnXyqrPYOxX97wNS3SM1PLrENR05JFzzYBcl6lnn
w6Bryedeyr+IbjSwzE8jrZX9yVEsjx6MfzqAzjVS9jdEleQAsDZNhm0XCt3GtWz3
6oqMDow9Qjw7V6ID8R/Et3MJh6laaydfCZ5SeZWoY2dk2XBx5e0zMTgwJl3ZsaAW
ocn6NTlO/9V7g+0AoAvY1QQxwYZ+oT1a4nCFRb2UXnk9UCg49xbbg7HfOGv9pxPH
Ont8r1TXaAniaS5AbTlIKahD+glBxE90POZ2PKogqtvRBhD2LDuPk1gJA/F71Z5w
pQ8sYejDhi1BMk8Qd23GtJNLy7G8GGfq+Vzn/vq/mRfE4JzbKmtUQBwgUe2HYpEO
jMMFwbCQbr7QvBiw1Ppn2NyJHqo2PNX0rr1o6ImqFflL/j462FGsaxfI5wf3yGrg
NhOwMlXVuvhX2vplUU8zX4HRj97x0PbdVl6HPjDUJC5siTbWZMFMMxpcTmQAJhGX
YaCjB79Gm0R3DRm1XKwd8TWqDhqnUDE/WHMn9hdhz66fw+h1M6gHk1qD27Tpd7Ff
EdFl/mnM9SCMj0418hd4igecBcbof704WW4so2pghMle3fyj4BJnLPR+HTPJ/eBb
fXd2FKbYqd2yXZgusQWCOdaQmN0eqXVmBjqq1SLkXmo1ZWS2L7D79PprfhAwVYe/
BuIQ+/MMxtkcSZzNz7ql+p2H+YMenLhjMF9iFoIB5HPeb1/LUINuoXgt2KagqHV/
xOOEQnPDsvrK3fDggNJWbR2f2iMBeb53FHjxDJDVgxcmmyJQCkJ245eV6VoCNTJd
THitZ4G5rp/BKF+nzNHba/37mpSoeQpZ8odSkt6tEnlrqfqErEarPpLqYAO7zwG1
Bo7Af25JAIzui2V6VR7/Ixm16Nd7iXQ2A+4D7E0WmkvwmqyvN3KPnYfB/DCFRHoV
cyB94ZSbeuyGyjgkL7hrkuFON9LImchOUhmn0cZ7GZzxYtMMytgjCtZS/2IxDFzz
Lk4O2YBLJY63haBAK7p3XWiNyQI3YvkVZFs1n3VZosniycdcbakMQrZZX7T7OKhl
p74ykUa7cgaDbFdDkm2ZdXlEdcCyKfH6dnLVpfsaqaZWnLqkfYCx1P4/Lv+v6QUV
BupG37L7WdTXIxhCkcWBGbHJ1Lvp4uiLBXuB8VbesYswt4ePtwQXoQDG2TH0O6ir
7Hy1uYCMlAZxwgoxN2bs2J9PMyO1C5GbxLZQwKh6qaz3bMBJO4mDwSFO/CieQylE
RByaoCQkV2Rwmt5fK3cd1hSeZeGYCz3frPZgcq/iUf59xkFOMEHsixJ9ZKmBp8TQ
iOwPmUVlBAB6+n5qAE++D4f/urpf5VFp9/UMCe4xDhnda/nIaJv6Ah3jly4Q70Db
kv4+Qs1ahSd5UNCBaWpHvf22oSx9pvsxfIK/2Hji3Kaicj0fARlFTRhGJnCGVqqP
1PGPzcORPRacYQVEj0pBEIsoANaSYnD5+zgyGidEAioam5Yt07fZBpek+jeeFQC9
YBkpcAwzYaTpHE/z9JvB5LWa8AfiqexAWUh61UzsKkTaj8upGkXV8nPb3pHwdLDk
iQ0pBNtFV4Kl+Tb0B7sO+LOWQizjQX3dWtF9WdHLdhcEPpfYDJWxTgLgvRpuVnkG
DB7ltHxt5A2v/Nn1JwFkWETHmK3QJ+7dFZDhjS92cG+rvAJ+GrMhHe5F8+kFZgI4
oox66/SzncDEQ6ODFmjD2A8oJTher1m39Fjx+Lnxm8KU+kaR8k+2bNGGsm3LTrC5
oJeWw/1EAE546AN1j4DCs5lbGg+2mgIsaLVVmWz0tOCtJj1rkbnc5RNsce0kJcLj
YK2mUgc9ZdkcKLYAeGsMrCbvrRf3EqbjdwYUnafUC8AmMZmLSGoww4bpQK3PRv/R
tMihHjl6iQJh5LPgyPv2YY93qfaW+BtdZhoAefwg6/4qi+NbQjUJtIpMLysJ1nPh
RM69/VhZKWv4ujQEnmMhBIq8LtgfLmi1SQLWjxxVGbd9yF2vAdwPLs9j4NfzKqf3
POQko61D5R7D4HTbjfMoKrZAEfPUaAw4owytfPMn5ZXz0VI5hbPyX+6cekZ2/9pn
T2sRL/Yf4TN0EB2RW2btGfGlmHlkjAQzu0yqsu/MyZEniwXYGtFSAb6y8YfVj3Uf
zzYwAUmxgkO58zKTARtzZAvNl+sDEpoiZfp61c8H6O4KfHDKt6gv9b5G+ZvlSVJ0
OGD+P8gohNrkEk7h0Eb21Zecg5/AttlLsCujiKqos0XLz1zODmbCYLq19PisUJbT
zcKDcQ/f14bO5KKqrxU750V+UY2pBYFUd2KxFV/4LYa1rr53wIArpVysfjpNylB2
RIxFtrQCh4IvSogDe9u6czeLMXvCxAnYrIpQ3XyfnoVLBHiCvfa7M56CfTHk8ymN
quK2kTBb4Pnq/r5e+29pa0QAIWOgQfXI1L37hWBgEpLftF/jCaP9WaH56+iowoam
xa+aTA/QnTMfnUhLNNqzbapSvLKUrl/S1qhc8abwQ7zmkZ2p98ZwHo1qSAJmace6
iWFcPY26Ac39UjABFcFS6HGd1sK0p2qzcQVI46wenYxT0Q2GeYO4DauSplyTyOkQ
sPveRBvc2a48q7NztUkgLeU2/KdXcJFbSMl8PK5m0uouXx85WW6Fu9QK1d71nyNw
OSYGwtrTYHKWo0Od27hbRr5mKesutXM+btKONTpGps1K8EvdnT1fYim+UeDvEarw
a6ebLmD1fsNakhDOJoljoQ6r/ztaGnEi53g955JRc/BVIl8woVPOOr8W/69jhkhb
Si8iZ3Dn6gVztL/Wz60OeWNEyj74wizPBP63u8jhOop1bfOZnjGuzW1Aa1qRxdyp
3Ai7rqxz1JAj6yedUoaUsscAJJ73fzUxmknZ8tQfROHR9WY0+1qs7UZivBIUkrGD
KPShOQdVYKO9UFrIRzUyJJdJKR81EnZkcdiOuKsq9EvUKl0O8w1GqVdmV/CYOqn8
rBXPr6TNfVSgYFAIOyDTnrcaDQF+DXiHltZ+U+TMNlgRLJUWGvZjWyiYyTKEg6RM
zQv2cy262LDnk/mR+had6h+t9hq3rsPORMQRCDtaw5agWjzr1yXlkESW1Z4uYYR1
gNisRWgPK9vMKKLNWqg+81Rd36vek8Jp2EGRWbpuyWEO55N0w3PL0LSJGortfn/n
k0rOaDKRvg2qSvpQS26o5MtF0PI39EPPKNoXgzAebF770JThnAiXHG+mAUYDomU+
HOvVjzhvdq/5eGNSSVlVJtRfutjthTUi6fYhbLUKk3wXG6F4QNUBdgs9zOonzSAv
CNkZDOdUrV/XKpclhRoZMFlMXqETRU4NupEKG+cCsvlgl2rXgh895IuaUay7nUdu
it33zVza744s25ZMl7MFLitEYqP3jkeF55xGnUMoW7v2aqA+hM0iDfAwR3k0aNdw
dURnhDK1cut7GbwI5eF+afmUADCc5IK2GMfoONA0CE/xWKMa8IacESm9qn9Fpfyp
oxUtSiEh1FWFn0WfZ/ELgegRSczXtqFPkDmLKhREOatxMrsy7gfou48N27Zv8gZe
WveKQd6tOZ+yRtdHsvT2kNcJZk/dPBlQdHJqWZ8YghDyk+HF7q50gpHd2zXUF3KN
gOtqF6TAJ3LtQ015aqmn+u4GGUSzM3GfgjvpZ3UUgPpaWfP8cgZxtDPSIcDf0a0m
2A/f572GqH90T0HAQW+Wfz/WSuMa9LZzr95MWwp/qvuTHx9wcSdYYK1CM1JgyQcB
3twzt0cK6HKVek8OGJfmt8R32op4xwvDty0PIKDiLE5H7kVrI+fdcKd/I5+C9i/g
0jgPMhDDuxqvz/DUZs2CkOFjYMgeQkCOpQsjvqZw9PPLvi/Xxmg9RzPpvOvKtM6A
zEkCr0BY1B9f+a3J9t6NWsEIcUZ93x9UeecWBBxqrSytx4T8q+X//g4qTVNUuqy3
708eiK6sjYwAvZATBbTxkBWkKEqAYb4GfUbHzGXvD0m0rUklFotYI7XpnGEKPKaS
9OouCFN1p3VpCYzRYKT4dM2EdmJz45jpvheIRgVyHOnXTlUbiBjyjrnKS2rJh6ui
XDgSE3Zrd5eAG+EXLG6NEUGPYm+WOVqtDlhLW/KyMwuQZpBzmeHWamXNK3fmv7fP
so/dAWxMUxTDPH7Mn++gDOj29LR21ZokaL6nxYpIOlJX31jS//KKl5ixQRDyCqTG
EcKaAi2HGYbJjehV9+6XKib6FslnUy1DSp7r4D8bmncon/4M+ggGFzBQjqURExnU
HHXNOCME+MrG9Xseb2OuqfyjEGpX7ZR2vmPVKrrfNN+s4Q2963i6nGcie3JW+aeT
/+JVUnnH/ushpRxmkXAFQ/hcGpgcJG1SRdyydkqOdGoHkYs04uRXMwnIYL0nNnp9
BhA35Qz2Rhv3p+dUj9vnrLkweNF+dKNqZsX1VLnfWKGuRRVSu9KHI25L9La0QHTY
v1RtffC8X1KJiH6I3k9kazBYhwCQ2DTAaIXv75u52bI+c8RgSyPZP63tLlTivogH
IpK8EfiM1BZavHEd25TMxtYvFsyrX93vW2blUpS6/dpXMZ1pq7IUKRxXBjxM0qB1
9Xz9rblk9c1d9w4I20ufkq3hle2jfRv9c/NyNTwY5NGs3329hP5MAdaZ7v+J57pc
Hp5VH1BAH9sjQhs4I4iLfDb0f7QfoAGChSYsF444zKJJa4C6MLpVOF5vMfuHpCQ5
8vzWJ6YReSXI6emvLN7fvGzx6jDNZ3GUg3GGKOvYiCkU2fmDStE5N1vZ082lV5oi
fR3jxH4gSChRAvqVv4VtYaN6hVOJb1JfloCZ7l79DKsOlFhn6s15Iml/AHKgcNxw
Xf+bTPKIHsu9tdyfJ8GeEFGnthqGZwJLL62S1IiqT2gyKdnQFBvRl6xgWicwFzw/
HuWW1nTte/YCBe3R+FGuuUYWcagUXfEMMEBLfvHcA+ZZhHPumMk6UfnBusn97xAH
SGcJTcaYqI9t7gL3TlW69GY+4OJoz35fDSfcDlT1ebK6g99T9bICYsdq3mk9aT3/
R5oWX0+2AWwp1YXGc2H/OsNyuDPQ/dGJXRv9kpMiBCKEWGcj7vEZKIOmo6WSY1cU
wJtv0KHC7/9SILUochqYYC9s2SRv9sn0fnmZHPKY93Zq8x2/Xesxynw58xjvm9XG
Gn2/lfZDOFVFhRB4O728XIlX/Q9qqGqK3kojy0cJnds4zrzqcPbOYm03Z4Rg6TYk
bgl0lCjxeNNPh12OjTyoIwqIveITYMG+Vn88dGzRu1lgbpreNML6l3u1anfWo9TR
170zmw7tJks5/6KGyizHRD2NZ/tE6U9zS472w64AQX8tmN+TqrAL1a5k7qRqti8r
biSeEln2A6LnLQG+/o8c3tCxOMdeR/vcwygzSCCH6nqhX2Jzo5P9mvUIFC2NzdT2
pRh2CSz0TDyydsEfZ0Ob/2scUgpFey66GJp2tRnVXhtYuQm2ATcdXEo5sbjr8A9p
9GjptcnPpFtd2Iz2DWSylXG58yw03QW8Zuw6AR6BdZcMa0k2FUigqajDx7IPCwbi
5cZ4CAaJF9vt5/xS4AqWsMv9DZHgFm9FbuwUPgBnd3807PrhfZtA4ZaBPWjNCDDM
RF1VQgVdFh/+XGD6ohzzp7xmTXPFjyj3EkKWm9STN6zU7reYUGM2mBFFnev7Foy4
YdYfFdv5PocNqvXXjvLxgDn5LqQ+Uom/if1d1Y1TMKRKR2A3WH6dqy5k2XWYz0T9
ppJPdZfAXHaiqdhBC9BbDYYsmMt6jFqkW3vgzqxgKpayt1lohYErkEBiWGdzgNiD
1+TB1/3RyKJmU+7h0Us8flWpCN0mBJE9gUjIIG67J/jPzgzucGaOe+3XjOoOAL4l
8ahaBYSXz5ZqhvPql5eHTwqOr5/rHL1TTbdlVwR1Zt7nRSZ6klrqC+eRBltnW4JW
2egkvsiEnBf+GoT8/45HJXu+jO1tpZN2L+i+SwRy9AICxGftlEMKkRI9X0xO9gWO
t28YoTsxQJQyAtDtwyZoV8byDOJ57zbYGWPq2cKZ0MAGb2QRkcHiDhO7mch8GzU+
Yp+C/j0INxcVx4p1whLhggqPqPgqaTUp0t9WPDCLg0dhn/JRa4kELDaoifdgjyc8
/cEOioO2OSXG1DE5N1LJdLNMI/YPYPdhyd6JHh1x2ndXRrAXzy+Wz2D4PzL83NdB
w3V9ZxjD0GMBJYtrWKiY8H7SpqkPoVOC6lBX4KctR0fKXF+b3QunQMBrXFwqnBWm
kBw3VPt1mP3un5rLyk8jCYtdE+dx/ok2uq/VxGUjPBpaeMs3zrRYNkptDWZbagFD
qR+BmDTI/yiZqIGmS2D8BGnE07q4NfRR8tTyfbN4xGUirv13j9SQGO0+MxkGCtDL
OFDB1XOgl/6v1Jg/Gt08rV4RcUUItJ1Bz+0WewN1Ae05HAkNY0nofWZfm9eNbjco
RsyOm/hqzFzTprGIbnCpjq51zsspShJk7eVwq12VxN+v/NRnKL9wZ3OZTquEg5oY
SgWNyOWhm9TTrJn2sFjFfDHqwlY1SKPThcz0vKh7DTCVdxuq8HvzcLW0Q+XghLLU
fjG6j8FKiI9pgs08BMqCAl4hBmIRnP8GqDz50U3DnLXhPziq6WMknJnic3iaN+SU
7xsweSeypgDjYkByDHLvaD1W3a6XxrqnCmnXwT3GcuL2ScTaF0iCpiTWhJ2eYUY3
vxYMHJTFuLBBNp4gnpC5+yTPZK9QWNf6aVAkvxAPbrtp/8Eilk/h2kxa1qzTbK0P
OMRyX6Po3iWv2R9t9zu14IuX99HVvav/rCiwu3xqc1JleK4i6imwL7U2nj9AOn3G
hQGaFeGsuwHJHPN3aeHMpbxVZw3IXNRtS2dETiRZRMrTSj1/j0GZuHcoRKKYuU1d
4+AM/McZLDGqV3vegzaRjlhS/zzUHmzr6zPl7YKxEs++jJ9800w4nYSWrjgONtvn
JnPWpPD4Sw1U+osSqTwxhpeqUWChEIs5IobcBA+8iC2VmgPNHDG6QGJNJDuOTs8l
lW7fIZcUdVFSZG/W2vZqLtqS21gUOJy8NY00Dn8X/PeKqok7gKLFknScdfFZs6hK
XEYgqehuV/IOonS8uqeqm/5+LZOiTpMaJiSrCrKzVHtTK5GPY7pnqBSHo9IeqeXv
lE0X/4XTZNfNkN+yOMYU2+T/MWjI5BKiUMmIkxfR89j8A8fSHFHHQ5oMjXH5Cjxa
fKVLOFFSg2qIhW/F/88ZXaJPcARBRimxLfKKqLpfxmXu2nNFibiunJ0oGZ5Ivybc
3b/hoVDhi03Yzxsp66IIZWC8WxvS7K32pyBjYpfqd0FEpnP/F1C7mndkCnhtuAhH
0O12ssk6ic8tUCaItCbcINmC7xflfES6MzCbJRsrdTKeCwkUna3jU45+QDVzj92V
b5/NZehyWWqNDI5tCYWix3bn0CxvHB+7vtXP+B6F6c3RlqPEnHbwFNDlsNtpVAf9
hxz/nWJEvNdcLvWVokCNPtrN1J8iRFv8SiFb/gudfSRtX+aukw9FMfCK4MS1Gtcv
K5r9MszmHVzooszBdGZWjCP3cgBZU1O2lhy4pcjN5cXUPfynx0Y8VmCtLkxMUvit
73yp6PielZypqHS2hudHVF39TjgGEDvGKfd5DRtj3/UExy4cXnVKKlOZpcaHgZSm
fW+EfPnLwML/wPJPGkXhd/Rd1d5zc0F5y5i6Udz22LV6hMVi09eiLsWR63e4KCzu
Ewwpr6l6AGMPnZ/AlD6jHiIFlODICrzT8OpkJ6qE6J5yr8gnNa8j9MevJSkD9doK
gUjlWv/yqrMAKIaqUkvNpQFLL4ucN0dt3/svbnJBrRIFR3TZelEeO7RhMOmI9jyw
L9apJ2Myi0la0UoplhvbuLsOKPHWkghk/i/Jn9M8e7aTYNTOsUEerFkOM4Vl3ux2
Re4MUjLNS76s0k9NsT829hJE2+VigJnUVL9/PAT0oLrTmBQ9XvEnYA302/VORFqw
I//gYN7te0elknZm2t/QmEhGh9s1vFB5Yy6QcO8cvUsFb7VGfheP3Vbg6eOCIa30
FcuFnPp5p8872v2pud7DtwEwEHsWT9CG3ts5sxfaglOgYcrIxpcdrqgYMkr56rQ6
tGP3gGW2FDk4MudAX9sKtsF7aAlcIk7XH+0jpzkPhR0mG3jg1isGZE12P9b3TNSm
sX0BDWiTFVwr0mVPnQq38A23aY5HwPGs1ghUxiANQN9JM4um8M9KFbHEZZPU+W8V
zZd4QsmohDnMUTwqEFJmDdRUNTnm6MzPWa6fQuHlXBRlZ9++lQ1IBN54mJl8Nstc
JxBB0pB/eafTvaH4Numh1c/IjjUCsrFfKCVeHus1c1XvdfYFwrbJzGMHZ5BxPRQd
RQN4xh3EbjH8OO54vnBLh4tlLQCXDV6jGTBjZDS34nM/LfaRGBepG+Y5l4QRfOCD
O4ciOQRuT+vRUS7WM6wkmVnvNbQ+P800kakMSmqU5cBExSJVT2munM98FX+AWMB9
YsdzhDXHU4ZAZ65lUe70y59P63kQxENvBtkwrfwrHhV+OQ8u+iTR90Hc0lUqzXiP
TG5xps3A/h7mIh9NjRzBliz9VvgcClgC1uzXPVXTPju0QRguMzpTVgWivclvTRQb
bUNJrmiWNr9NUqU7+5JgeDjap0J9JFrqnxffoa0gmh92mbHoDjNxFNfQw8tfnvlz
FpgD02vrFqs9xBdLD1wUR9J5WWlLaaQrv7JxHqJ5KGO1lrMWkqoJ+nw8pFajNJ46
0Io/umLC7IfrqVh6XzMS/x/QCP3MRxg6HmgGi7+PNR6GHVQDa+JINoAqsa/w2iz7
OHNCYO1y2GLsLhW7WM8CdI1Dheu6OtGqubFYeUWIl6OSDYX1SZVInuOC8G1DMcLS
FlSf/Tt3dNQovY4wcgmNxu4L/i95mEiIEemKkJ1bBYTkbYkv/cZj9r+wRdqZ8uA9
B8rNsBYz7zyM48TPetyVRT3sHEHErgdxyWQKr8wG730X13jd4WQu3tzBufAJ2omL
escMqDCJpLDo0xPzxW9acV7Dn9wH7RpXdN3XEvnuWaSx2d1MlSs+haEI/XpSiV3Q
wGk0QZFga6CZeFQnBFB60Ejyg4MflADSbIaevU2LeyeRI/SLZUcrTwW/nXC/UwA1
rkpFJiW1JrvfE75qiPAqwi52KeKifVevdQPqpUrSe/MtWu+EfePoDd9/4UPUgboW
ITfXhpC084w+QOENav3UFgXMBEY9opN6qlo4ALpz9x8y3GR3SWAETtrjW0qljkIV
HaADbId70yDhGL4uT0q0Jhk+VUk5gX7lPZ/Ee380M5FI5Wk4EJskeEns1U6NwshW
QJjYOWcsGMgs6nPuHwrdAkiNqV+BYTGNST0/Lt5Zo6bPnQZwW3PltKpUUrbmAt/+
76uuG8+wT8fi3OrU9kVxrv28yhO78DE+i4OHn6/h/nFj4kHWIgEEc5fc9uKtDrgC
M28vYEG94nElUZQblP2PTcAMSbXqSm1vcKw9i/Q298Bfk+SZlW/b4ZWOixDkzsf9
b9sQreucldDoR6ue3d4BeDaPWE2NPYxfRIyF0Guv4+Lgto4QDbVrQOY1Nk0i9Jq/
r3Fglx3C01MgwPqAtJz0EFDP9Ni7HkYmrwphFZY9xJ854JB3u3Ow69R0MhMInKuG
2ivIJTz9jmKJKXd3uu/Wvzbu88J5My6JzBApRQvMpgAut30UiBhnSK0bdQTZ+Br2
DxlgA3eYfq0VthGzoWdkTFqmuTnxHoPAxcFhPBFsoqWyH9bDs6/oXRktcR0MigBR
J3UJnEGDWxPEmMJzkZvNfPsftH1ly0tyNscBOvD/9G6rNCg38MOqZsFQcuNYtjwB
yf5bG6XwzUqh5QUSdUMKnyZdCHv0JpyU8TrjoGlbGYjvKyKL5UiPmDcp6PD51AQB
FEN2ZKPIrzv+2Crmd0glW/GSJWlGWeLSMfuP38eqQYWpiRKiNuuu+PF/RKr+v90H
WR2paMlqK696xxfK4RpqgEO/NS8k9X6h7DHKT21UykwDOezruu7EuWc/F1eHVirH
4xUIvY1grI05ntJ7yFQAaosn9CC5klVvutStwqdcYld5eLOeLknmugYZB5+7ttbc
9HN/pQit7MZQsghUHfwkEgLW1pU1/iJCzi9kLs6JcznmqeOQ1LMnPkHSrmobJBKM
gSGKR3gzCtsTfQZ4gP/aNI8FNjUOQm3vzajxF8kIC1v4OTaqo9VNsNH2JZ5Gb7hp
Ui2BZGiT7wWlszix8BRbcFeuHTihySaLxaM4OpCOI81fHEa162zqP1U0aZBHyiTQ
Ej8PGxO4pCEuFXdO8YknW3URp5AJ66ThKvXNHTSRWtxFvEb1BIeCZ1hqEC6Z6Hix
7wL0WDYy8odgRurvC56+2LKbRl7qbl0oViSMlWYI7hXSTXuyx2+P/D8D0jGP/DWT
etE5OaD2jrfJeBfS8NjfSGj6MCN+REoK04K6ngy8lO/Gx4REfRYPDx3b3DrK6CSj
6yjXpvKaC/GVRxUBiDswn7/YKYzJOgpbAIt55ytCkYdl9iZiG5Jb3+yD3AvFuNJd
UNSPWCrtMYhAZCPtau+PZiPyYA+l3ydR1s7yPpZgv5VtQ8sO5ZrsOiQFONof+cTX
kjgyjmQjeKzApMUREm/lfXutpQ0VzPOUPqx2f+Xa38oMeXhqYVQzX3ngCdzIoozv
LdbWIXpFXYltdDBcPhh2jxoISj9M2Dc6tR0b7HO4Cos4hYZEA3jg16tQp3dUSFyh
+f0iKb7Slbq+TKkQXk6JcKTAQe0huR5rNh5V4+Xj73BeTpSZbkAaFDxX5YVDv2ky
mrAs89wCvJMZj77qvh/Geb+4y1fXXhd+DEXjAZcglte2X5niIsh2UqYS//m+Dc0/
xwAKRDjpPHdw8AhlXIY2ZKBAn3UY7QYQOkgP7lwcYGZ7v89bvU5RmPvetzXFHrZn
jzKtf4NXjsNqS8tzQjM5LYiz36BX/Hppa5ebBMIBzEPqVOhvH6Qi46kwz/wvHq1d
uKsZMPWhKRSs7/B+4saMxzfhlgcavpZfy2bK0Y+NkhZo7fZa+BDn272SRWBLo2Hc
jTnI2xD89at/tcDOkCMtt30jWwgdmOjjVrFETJ7wB/3Wot61IC+43zEo18YCMmdt
V0hlt9wjIEbIEycv54jxKcaR+Nc6WvtDkCdSil/fsri4FbWAA+va52s7CZc5ILV/
IjeE5Tp5IQIngOR+GoWK5hggkc0d4A9hA5iS6HmVoFPz39xDNXXamKCdCY/0NpKK
1tTaRwv8qacO69day1YC9b4SKX49RTE4PnnNCRILLQLOeC5AZNUOkow7e6Fjq9Ai
95tlyFR4G1EcnROc0zltS3nM8UuhYI3em4N3ToPP7/jP4dJBD8TCixFAwU7IzzS9
yqkHzWBYoNtI9/aORR/5qA6D/H7WimzAJAZ8gxTAae3DkCd0g5U+meAUFI5JPm3W
imWe+eDC3hZxJOwaYeEBOJCuyudfvNDqeS9wwyh/1vK2SFTlAyfLkq0WKM2Goro8
/GJrp1NYbzonXLB1RzDTw2dAmDkWZii79lcXFZDYi9EnI3e8j7G4xmCkDm2C2Kjg
SFdlzytUvS1+zARE2ZH7BUHLDd1cleJnXxF6z4kOdmIAHnZMYrXRFa2UoCY08P01
t8lgEtJndPy+5pXXPYdB0tIh7L3fUcFqg/CQk6+KjP5jiUTnAjZtywDE9HRGm6K+
W4VGW4XOYiAyM1DEvnl9N4MlVQO+byldHmQiY99XT8MZnO/pf6+AxtYuVGtIH0oE
ACbsCl91Ej4aQvvB1WmUziaX+pEwASh1C4L/8NpaD2Wq3nSf5Q+WG0Arv3LfKrE3
rV+91f/S9t4D+UBT3xg2IQ0caRGL9O5MCY1pj/5S4AwLhsZAYcD3UrNEseR7XJ/5
86yrQZnXSfuL7OWEwLKlxfN6Jes0xryyFZlGCMrAB5jb0QXg3EPgQeoy0Cdfjlb8
4mBLQBsoiZk+0fBCHtuoC2ZeOrxYvKPvwCKiWMXKUyfDHe2jljnzFHBa7CcB3HrH
1XK2v6Xfcac3RTn0bih8wpeUtKmJCClZNzqjsFormCvLkToTGSf2feZvl1xZoHHQ
4MV9UOXugw5sZq/3vYVvWAz+m/KWnyHLxn+MLvxFn6v96a7F8zt/1Ylw8V6I3uUx
3hYvWFDQFu7SWPw5VSBKKTdnFqF1TLgHUifUOrYmX8/3ay59/N3OR7L8LTYGZ2Gl
+OJYrqV+nnd3UkDP8qxGYLp+sj6qaLh1KEAEc8pC4GmPHTq867GPf0qdQqB0Q1VK
SMRKSkOh4f39IBWtaVAPcWp26t4cxsXlDcjX0LUE6Fm62G4i60guyirL6fNL1BuX
rx5EA41oWtKOjUqyumJO3XMuR2Encu2R6w3BC0etUA4nJLNXaZXS0qm1rQmak4xg
kIsiX7FIFkRPBCcwKx3Jd4FbTaY4jW54UE0QoNbmjYjTkBNiqppamcGsdt4GZiAL
8IAhwSARdup9yADCxNjnlUG9V0885dzOpPuzyPVdbGxe7eBWJfoDNRiUN2KDGCGU
rL3BLK2SFrvqHQalhtJtOm8o0n25ugPILpdxJMkPj2IploFhC4CdZbDB0lEywhXo
D4HY0SLPslJ9agWcQWrOUJK30IGpElLwKyTlghhSNh2O+TE4l3BWwwFZzPPXw6bM
ot8RUhJfYR14voll0I1W/O6oEghNJtRUgY/HGl3ESbBSDKkNRTTmrq1Ee74I3oIj
Ti1SyXXnp2NOQN/v31qpaFvlt3lMfOM7+WfgLaUApWq8dPNCubZa60kBR3zKaqfF
4yshMUYsSswprwCzCJNAMyWOQS58Jv/yHMHNcGlCn80yIo/qwMGvl9yQ6SnaCzKg
4XGEUz4HnGyYkePhTIIvb3ZpEmsuLpzeCxMbFAiCoUuqSFjNytJYFmopVRQ0Z8D8
L71UwS+MRrEdI0BbaRGl0+VT4lY8TmeIgnsK9SVtY3qrFUE1F+KVtXKlbl6LHvA4
vLaVOMGkCGl6Gg0qHgGD727OttEZe85CNYqAi0L7vBPAASUnIEBkUw03vwEULVZB
ELbl6RBeoY8BtyEC3IJu9ilOAwRiUtNW19S7Ao5QJ6qcP6sq/9Gdu9JcEDjbH7Of
W3faj55OBdTnGdyllcTf5EpHlQhkpzeDu6hQpwYrDgW93mE8hUtj5xCqGybzYcy0
//FjaKahWfaSCplcxbNIv0SdOgbPv2HljlwqVwJrzPP51mMV97xTnLGbmDV+b/sd
ZEsyokTbQaPq6jI17btUVQBfYqQB/zQ7j0je/XjXogIUB5uALGPnP5q16bv7+oXt
gacdB5ZCEN8Bnt+l4jXsEdRoh0lQ+fKmMgndFWKSLilprBZ6vKRB8pi3H9wWGTOl
kc4wrIIhY5aA6hmX9IFCwFm6nCmH4bU3bGSYv347kI8/nu/osh9EMrFx0y1de+WM
OwU3y8WH3dyI+5+Itj8iHPgaiYfTcB/l4T5NB9zlogbGGR3xYiesuW9FAbNMbSt2
hbWT9Q0KxM5IpFYaMdFeAHVTbzL07Thtf8pXjuUTXvowYdv7Ewyl+sQfd2C2qk+C
7v1AAiLELTTKfGoQ+wpXk56WWMJME4rkgil/dYdhW39WysL38IwTvhnYg6bYX31P
SVXXT6t19A1xkSAgD7XhKEM5Ofjjcfoc/AWoV+mTdte2V721/SIBap4d5DbuanHA
01K/2paazu1Nhee/unG/UCH/pTg3qPYPh1iDZq2EhxTPRzjJSX8w8w9wy2rYAV9h
L/9z7MfnD5gvSDi8Rn1NF/GPl1GzdU2qlLoccHcyfmxyZTJn7wODNW30HGpGNa1c
TiQ8s/IUGJY5uW7r2NOqhy/PDjWOiH/OsOt0r6mqmZW4lMKTX3XKDri2zIWrTheP
v/hBMXslx4fJUjVnFHAsbPuLwl6wA7gNHDTZeFSJiaocsV+queHsUikyQXz0wnbu
UO7g2GneW/JTHr/ryf7A800fMH/Vx4gSHkqTgJi2tbWuvSb4Yo2U7nEP2BqsKZbO
PfqSzv6/yauxd6qdIxtLjagHt2SLLfWn+Ibrqh9eXNJxZDfGL7l2X2ZFX/4WDkTm
3IouGWan8hiXvrxnUQvjPTugJ6tu/zSfD9V35rSoOvGlewOEx1JNMyrLimX7dfbL
kvoMkNwp6PXMxtdayLsUBse1FwxeA/TK05x/zKRWT77PaaYozpPfmCCb19dWkbKu
MMNnbQ8sC+mcXwDBRn/GMJPnirfv8LJ1xzgS8sPONPNlXGI/jGg8A1XGg5PM/DvW
NZcHsrSF1cRtC1NzY0SOYaTzDLvb317wCpai6t2Ps/KAUhTOb8ONOWIAtzZ5NA2i
YUYQQdfmoO89cAkOVHzPmLTqlkF8YwSyXspiSu6aO7lW65t5XW9orTBSr9ZZehd/
EisFDy7cDIRP7EK2RTE/+XpCssNAWHH0RQ5qLZxDK9HwlyiEGkoRlFQCisBdUQcB
WtWo2ONq4yz/VobiJ0k68jgUbQv7KETatKbwquvnCeaPL0y1BElKlsX98i7g6UH2
H3hGVpD+3G90o7Gsn5ABRa9NtfxjBxvwrJAoNnFmoUTV/R3FS+TSQMkGPMQ/Mewb
6fKY31xS0AG+j+GecBq7bDSxv+VjwAHXcPVrUafCkc2kGnP4G2sMgthB6c3xZo2Y
nkE12sFPLRoHGkpmgTeU6SvNvYSKINleE247zVjWKH/RPP/cEn9sQCnmf/c3/qOb
YSA0saCi645x1iXhSmGxhyOOb0lvz+t34JvE5TH2Uc/u/z4ImBe7vwCABHyFE/QE
ig8R94sTVW1CQ8DXk/PSn8pe2Wt9RcYL/ZwsLvjq0+wHn6dnSWtI+ZGEE5nUzu62
kGMb/qP7gzw/5NbvvaGHbgoegA21cUw+Sf86zJHXc1nQ79ZWZXXgT3+WHJuM7Tn5
Fu/qwEgkOYxZaPEXuxMzlAe+OKaom48CiKG0E30dZYcHaGFLjFiK4dK55SYa3fdN
WOxoPoK6JyzOEFTUkH46oR5p8RQ276XvJnuuPGDRBPlD74tbhr342TSU4qx+Lvlf
lfeKkctdWS+5YTaMvyJUn4nmxJrsIlJrpZorR5xNS/j2C7nuKsBIYE3tpJXWrG4P
PSH4xgBnbFuqRunka60O5Ex8TdeDmB81YS4C569jK4vFizKjkPSfgSpxDi+cbHeG
yP89hryyJyxOHMrNqSA3gFH1eL5bc1QHz5W8B10EPJZ43jgTPsxaWQVPoOsZg4yJ
nQbhC5MbBTvmIdJcaiixLyyXBRxebRsKnGJ5eAzyMtuzOCKMGNj41HJ4/ph5q4EP
bqVpyDkL1ksqUyDB2rGZ8OgoA4rcOoK+LH+haOOlxBi/Nv7biFYxPX+k+QMEEXHs
zHnP7rZgsSwXuAG9bKjyZZhTxIYqieOZm/LassJF9z2MjLPPIcWd9T73ox70BE6v
A2z8ThGzf3syzRZkXrCznA9oBqyIxrJn5J+dGGGKZDuZ3xyPYt6H2q9QOAhFPEEf
T6wXWidplqWkr0hlCrgTPPHpISQsPOtpZNpgDOL+TTvYDIiP3g0sBRmfQZekGGmW
cDgRr42djJ1xcqCJ4GZefPLGirA0iwLZ6OT00Lf9gYVHmYkHMch/CVaus8xyoR/a
V1jZIAFdygqSJLH0k13XbPgv38K7aK1Re3v4ZiqJZgj3L+A7lnJxbMjsJbpIt9m7
2XFWOMyO2oHKoMJpjLHNOI4c0JRC67fXx+V42kI6o3xUSw4FXi2yx1ZCP3Bwfnb3
H+yv/3t3m3EvUv3FSwV1x2X8IJTMa30DwTnuCLgLac2tM8ouOCm0KEEd7bdyPKeg
L2L/aPU9HnMjSvwY44G621QHUvv+zWgtv7bXU8mqwkgf/EUow2w1Hza4k1CSC+ob
sKZhw7soIyrc75qvl7YlqvzX9dn8Dk9SSWta0UU8nhbyit06TLhJHB21sBmcHneQ
5GC8T1rxR5Q10k+aexl5Nivx9XP7q4YbmjyQ0XzrzkWOD8v5OAghxz6MEQnl5NKx
PC2qlL1BO/e/PJVZ1Q3LW2tiGANH8gew3jAdNKo34e61S0cxn8y3mAJ+atWUV7UK
IEVQAQ32B3QsXCeHOQVu969i6CbGJNnQYlwY4TgXvio6NBep0rV7F99XZU6CQmus
esEG8ReAMRnKQ8yIcIp9/ir2HFzuis1oleLEntI9L0dkEwCd2JMLhvZBM8S3IR2X
vXt3a1c2z28nqjf1pdRnepkfgOVX+LjAG2dVnurjQ+BJN1US42GRORB7cqn4QYqA
4j5+oljQcqOGk8TXCHKgq4oGXmQ8oVGsDhGlERNeosRVG/iuex1+O0E6LQ41LqVh
4GFyn+8+bdl4U6V/xanwVchHAeWL946rmLA/g0Gcp+LSsNSCYlBn9n8YxGgXbwz+
3UMRmrmav9VLw0u7fQipAZnEigDbX2UKSVkOFSnsDy5cVjpS2caO9QPBXEopmH7Z
+wyPPH5bjqeGVOlV10C6ewBEN01NjHEHMC1JzkAAJJJs3YrLJEW8nqAlGM6b66VB
eZSTHhSwXnGJ+vTKm9xenL6pVsWbied2HgqBsbmqpcfBUAb5rIyaZH2zJLQW9rjv
zB7/bAiK6+zWt7bXDG0Afzesz47Abxl1hIbZw5Kf1PWPqTP1zR1mlVxRMjCZIcIB
kTeH8kKI8l3OrsAI2G2IRdeDUNQM2v/BocNyaDYQQnw4OkX6q/8imRfLbHGtCDFv
UPNuxnkbjwsfoVghlOxexPfu/n4WP5M8jAuI50JC1yXkOrINii9sV+7QIsZqVin7
R3S/E5D6QHV29eF6+HllQLGhB7RFao7lZRRNiye7JyMqCBGlZsG5oX0LjEkMxv73
bkOI0Tstlee5M/ZM9CshvSSeCTu7xWHGPn0bjvOzrWuM0IsN/6CFTksCPv9yS+W3
5Uxk3XTxlNrW0hNWNOGtg2R5i87EPnrlBKv15b5nItJy8nPBnTnzQClNooZSPpCE
AZU5V41uFUxnEdkx0R3TJ8Xj73d5nB6CU/gjvE50pSep7w460fBp5xOvM8xbp0Qn
0EzBQ1JPP8v2LqZ9oFTol/3LRigHCZx8JZxrjUSoP2qt9AvQSLUJhSGUosQ7xIB1
09KnoVGGfIW32rrG9/RgaXKwCfVXRxyrW8urD2esgwlIZ2x1oi0ZDH2oxC8cdcWA
CQK6yonvHYy2UCrZhf5uEqPzUEX3ZJuUPa78awjFeBRZ2EzQklTo021wecACk6KZ
pz7j+boF+I8j0ElGw3i1i+RbVSS0zKWGd+MIzSEj5DBkaFN+lnC6AWtPs9KdBR8/
WjsJni6DBMTvaiVx6aMHzBfdoKIoEZZWuiUHfTRDfnHHobcRxKaZySUGC3Fj+evs
U35GBVdnsYpZgFx8autvSVKerWg82ylRLlx0mndEO5ZkATNG1TPFT7GVw6J7uMCj
nKaQrkqxf0thhEwQxzn12FK/erIMZyKDLq8TzKLask3Hh26DNXyogPYOf7Tvqj1U
J3otP1O1e+O1bf9nqD1/0SNCcWTX4q9WOXYFV8atRSgygoat06T28CaReeWcp0vS
gn7KslUmgEOon7FhFPK2g8GtZHECfkwx7r2ioiOD4afBDba+Z1q5da4Bkv4Ep79B
Uby5uh0Y8sBwimKFXY+m77RR0iiBk25c0jVNX1S8xM3nJHxyeme00YB0NdXoqrxY
a+005+y7ya8p925pPTBTUJfDRrCOxgo7whdXiPlufK1bK13Adu7eCPeVvznm1Rnx
QlZHpv9AScwh1FkllbssEkzzIPal3ww9XqUGF1NieuLN3UU4lY4DvSnV2ajpg/MQ
Vgebcy4BwdNxAoO6yxgKYilqPbI6U6ET5YTMB+nlbJkGGZYl5iECxYez0nd9+hGj
PAlavJHVOJd1TOv4s5nw7fZbwpTbvyG5FYJ0C/Zy28U9tTE7Y8w4UCCYkP/E8oCf
HFOCBeKntMP9YnzaO4uu8HCn4bLR/9g5lbAU6YAiXnJGia3Lz4lPmLV/37IoWuhT
FLZRFJG/OGi22ZFM0bq9Ryq1WT0fe8ZU+V5Q19lqip0CeHbsVpE3mc+6CSYZm/iJ
rQf51QEeXhETehKYAZVmfmH2nZ9e8UAJtWFUhLEaN78wyeux0tKuA/IS5fhXtFXE
Z8TkQKUkgevU+frgs70zjZYAu0Qc8jvXVRb05/awZ5PVp+GurPHh1vyevyYQqshL
SED9V+V3lj6RuZeUWgUq1SzME0cXaMpasSTWc57ro9/YH2OTSBi0tnmtZEjxLrTc
qlNKNlnmCpVCXnxJs3StcM9CoCvBZ8DYpMgUHUCASGd3BnMVR58FW7rMfFH2UC+n
ffyFP5o2wfbCz97ljPpqhNcnWL6LYtnc6xu4JoB1RDWFJ+76zfdPRvLhe189Gnnj
bDq77lnAL6Tv69hvn5BzYXS8ys9bhTzNtrDRq+3Zc66x2CuhglYvE3mUxStYyIJO
+I31zhdAiPPEKeVNL9NGqdnA4EAW/GbH0KdKMXNFXxf4poxwUIo4LyyPobmfkCDF
rMC6QwaUJ5OZLdBZN6vPZbce7CsnByJWXD43/G3wWBYqDpepmzzsQj3IbFgw1dOP
idX46F4Iax/EfpEKhqC/DnCn/Zc6HmFUc8xMWXmAOXXPR4WIrIIw47QByiALB7sI
jyEh3O0kDhMgUtLDdm8V+yh6wH+IbVzOO8ghWWDeprvPiUaEeytt/P27wm9lQLZW
5kBfVtujnTS7pIMjN7jLOR3ujI/F2NwzkrGuu1YoZs5CfzlrduIH8javW+O2fCJx
S7B/AmfEKM20gQTdQQkGGgL463bb9HLbjoR3t/rXmxS815de/AqV+zCtkTA7xOv9
2g5YZaHx6fCVwpoJMBCtgp5+mdddDIvGG0PcC0ueMcEWXyNZZ/hBcQKOpWJc3xut
dVsWYHrm52WVkJ7DfkP0KTB7lPYYHfvV0LQyX5/YeoQPFjU9AkvjuyFe1j6wmRyI
/WW36yjNeZT2nC+DC1X6EaBxGmIFJFUPDhal11UFsm/t8zZDT3Sv5MBXazAY8k1H
0QLWlahLNerLzIl0Sd0Lwc7MdnRLsnuHxr2IoqyT93c4g3WnVhxUc7PPY18l1eCB
YEjAPqYZejpNJejwc+IJMeKT/oGvrpH+3RSLJl7rteBVxHy9lgdRbwjVZnXnIsnF
GKXCOVRR0vNQ5cLn5dgDJllmzTUVppIdMaJz5d6IJCu7tsUoj8Oe42QMhwEbgv1o
cu7jCMXZvuh8vOVNHllLdQu9Z3yZASVH1rRFWO22fPVbP+3qvT29FUrOKU5w28cB
3zcjVfMIpqQ7YQRNmqr6b3Oc0alf9DKx8+s45my05MKwAtBu8/TPKpXWCUl7BBj4
I9ceoGyGONCtYWNuB2AnG5aOGOf9ge0RO3CXe2Ml2MZkd6TTkpuoH9UJd1bcAHCF
mgnTKoF3TELopcKxQcEPS58/G44kajQek5CFTwKuGb73c/A1mpffXicPQ5Bs/u6D
Zm7HT/YUu+7FQMnJ07KsqwaOJIgykviqZAxOMCabHxriIhcrtbSuwftq6dV8G+Js
XmeVUJx9BdmGyAFSnjIawOD2cLLEpoQKyg3NFhIsYoTEyY2oJ7UtFQOy8R2JB9K3
ehUpHiqL/pay8uaHrVZXSud6Waq892x170c7PWQOSVHa/1/u8t97awo1C4BAc2tw
1T0srBkLoTx/y4/xZGhNYDeu1SnFxLMNGUYZ3+YUOgyH/1ZZqpZBKW8fnuEBuEnr
8yewT+KUUffSdWow3sMcl0XclDd7LhAmR8ND1Ply/euUbVAMIEgJwhrHe2wJ44eD
0CFIyIlywQZUj648bwDGfN/jkKwEjI7BZp1bNfPL54ckohvGNdoiK1MJMujr2qOT
4P2jiroGPhNXrBU2md3TQqQq/CYFadV9IwBr8Ug0zjLVV4x0vsWWhWmwqYgC3fhM
VH36pAFktUoCCbbGnIXW7FWbfyBQQwtrgAGfSTL8anmQPS/BjRMDwWVd+qr76rIA
NeuDt4HClF1mX74zwX5v1hCny3yV0CKPRR1l1bNfnbt/uKIMsxPlob9B+An8iwa9
a+Vj5hIpo8tOsqW81aB69H9fzBYSALaezJfaHumsEd6iG3BhrpExOOVjx2y5r8wd
N4Bt67c5iV+fl6ng4arv3FlZJ6WAeJ+S4yKym7fDg1udkWmJXW6M2wpqNEGCa8js
5c3k4uHVWVq9E0G0xR1BpOtAeVYIllalzLBrRCG1Jr236DevuHMx7VkIasx0tihV
j523yFUwYPrU/E9AatJc29PuQkQh2hqFr2E77Qmgi8gjWhaCNj9EdXhE4yUop3YA
hV4zpW5wNxFF8QyM/47jMq125oXym1tEaqaI7cxAt1bcpvKSfXlGWXsSasVMZLnu
9Rp8PAQdx8mTmIrG9LCXAf8F2e028+6ZjIDa56mERz1jD/bi+tetCflp0R3XIkeA
+l30TpldRxVi3ldvqNe3M57ijCFV7GKPZloHEjvM4pFqIPSNgPpkpphQ1/K3AkHy
2RxNxui4L0aChgSQYe1V2GkpLPqu1KuMHvqudAXdfwyEYaJpTfHMWyt7faY46lN6
kFjv3Vk3rfw1oNwhI8c87IgDmvu+KdH8C81nrgU28Cc2/h2ZLHLjnG6gmHaU1Q4P
yLjfNn+f3XeRFwM2qCvQ7U/TQxDX5Yg8fitrH/Nxji7qeaR12OYVf/hucwVSHzXH
oLwX/teFeeCOiLnMXUAANLvlQuieZWIeszr3Z0bOph1xqGWZMpkk8VpI5Ak+oQ9u
N34YR/H/1G6ZAnO2wy2VDvPly46dCTvO4IVrZPMg1w6uz0dFIxdn3ALTqlTcciyi
E2TqqtNSYOpUY0rPCpuTJ2UI0tuMa4KmFX5iyMOo7sGwG3/vjSQorbDjHUoxWvmd
H9XB7c0tkOm5LoRxNYSV+ZsHwdQQ3I8XvAsPYb0B9erttvWGs6Q6RUJOdecmv1mV
LVQM5D1xkkG+Qq1b5SZhWN7V0RImqGkyLc5uGIvnBiwUSHiioB8VbyXG6bBIEQt0
hIM7y1iyeUBXVaplqYNkDXdIYvCPQ/YEArf6wiWk9fUlZnKMarPk0gJdRG/uJ+29
Qfxf5mxEhS6nYdQ7jVCT3KjYJxeS7m4CaE1n0Ehgj/qRGB4AJsS6+GfacSKCYKgt
86GdJ7kOAf3RL7cBhUJgh57DBDolsSkVxMQSfHQ+VLSxWWYXmzCNEPdIuGVDVk/x
fE7kdkxOF2J4PoTE/4Rr1fBqjo3reDUjKAFXcfPOHB1PB3seExVHcYx7tUjAkPNN
WuuPIfbh8sEDRbV+y+kiNutC/R9Ldza/wxDCp66Ey8+TyzGctaPslhueoTm2KcVU
Hy5tdCblzdqS0zt8pzWpVRnHLrFAltyzggXwHjyytnoCF2Hx4UyDlEnRFhhVeOpc
0YCEzGvfom0oP+dD1wYcWq8jUiqr0iaYJiP9Jqkwapj7ff0J/szjKpwlgj5YAjw6
s3bt0sS1yj1xISU0qP6EiW4FeeLcx2QKHOWkmMifA7r6IjimD6lncmJJD+Lz4SkM
CWs54jeW0fYXn9N9N23VO4udm8MELJvlfn3sQY3dkcJ3ewoqWzOB7r8xBhj5endY
cxVOz+NZ5UloxuG/ccZoY73N/DEkYLM0/NXxMniZDycF/Kg90/cqedFFANkzC5kq
WNH5N96FuQV2Owo0syb3fgKuA/I14/ytShOMLjUBxwqqR1a9VAo0hEsq3tqUYPZt
pON0igo0YcVCAKHrFus424eQo/YSzm6nBbQBfPkwJ1Z6Ze/VenTRcYlidZsjFlU5
3o7+1yRMaZJlMSgaXxDAGXQQPlhErnEf+6Nv6vmxyhiU3sbw43RSc6s9MY5L7RjF
NADLijldb9oCKtYOKH9/kKhl0Gy+9XwZdgijec3eUBm1gSKDgdesGYpFNtxGyYmL
7CQmNSvYz4pE4qBNFpF84u3ZuxO6KJwPWJtSpkKmoD/EOGCOcBjciWG1dgHYVZ66
xKa3+85X23nbREH4a6jQbCHV1G9gXeR1nHTUtxMGkWe76CW/JR3mNx0Kz69ZXdRe
DqlnA2GMPL81VSGtJX45Z5WTNokJuRMQXIsYp1ihfnlVMSGIApKZvj7/6QZVhzlc
4Q5v0I2mTkBQXjmBGschidNxS4Lm08V1T0hYS+BPymGRZUc9xppEVR60XmnHCppN
AbdRl5mXV2d2gh2OLEnZ+3pxeg/keHbT1hv1ggF3Bczmgbl8t6K7hBBt3RbYpTpG
Ul3Rjz8AdG7CDyj2rrRKbnKf3B4t49PmQC98UydmBguSjDEOXyO/oQ9VwtjLX/OQ
pIwl3iFp++2D2mwbBPEhSDhVyI2NTALrpDkLBZDDq0jR+6RJYqn9h9hEgOnrFYJc
9oLC25ENOw8dcgWKIRlQANOBB0+UK1IMvD7c4N1/jiuMZo9C93HFv5ox54o1LpMl
QyfOZSSSCZ6ePzaU63Ne2gSa840kBZqZjO/vXroCbAcfdFGp9uEEHS+HgQX6oCJN
WXyfhuoOGRJ5MW39qOF/9asl+fXo4E01b8KO0mdamyjIdAwNR4C7nyPK0KfGEvyR
MtCdNyCY9UDuoGMwW1HYsBNWSk0VESYEUQL5IPQ/bUdfSL0Trqi+ugUnDmiPrwpp
Dk1kyUmE07Ks3mcDCL3xCiM9/WFnd2yoqhOftbUWCEwyj15yNm/tFt7Xg+JyvGYy
ELPvbiLfwHxtMW3VLbywBIlFZ2H/afTFNhCACdT+pZm5Z2lZzNu0/3mFqb0exYRo
WaUIxrdDrrzpiev3eusSDNkqKOGbOoYB8wtrpNfqT+0C3QuVYK24I2ZMswx6WE+3
HeCgqgH7RNIIRQfwBOTEOWp7/MGo1vf06c8D8YdSGiNC80vOmj1pTpUdY6+zLccI
3S7EYAWbKt0QAmp9kzKurW5VAXbDmuB3AU3jiomd5BunJjqEZwFdFASUAOIgwFUj
Vj7aLqwOzVeaB9bltZOLVu32FMJHaCUeAYN1xqg63bB41wH/GzCn4QUv7ZuH9Tzc
VyM5P5Rm8NfpEjIdwlahqXeMXm6/klFK5ECGyN8rVhwsXA+eOn1HQZ3zc78MvnGI
KPsJI/SKD9U1oXNE6KCy06CX0eCt27lhsUNpWFSGQ/irkM45SpW0Eiph5mgGgnwG
EkQkIl7FCLEnvF0rMBGJetF0Dowkow//jyb4hHsUn4oe6hWgDf/IxCdC53d8Q793
/9c2D6aj7A6jj0Dpuajv9jY4wq3HGK02mWQxSyQId7EajUM9pTi7aNcxqdvsY77e
7wCduvEw0LcU9cODgXOQjo23k2IYqr3FxNNfnFIFukDVBOVd4bfoOKlHc4LsVS+L
y8DIAuVX6QRr2bMteD4j3gyHWD31gHfn6kWqHIFUak1OdYbN9+Jo6tXA7VHDztGq
6Ad5ZC7IZUQ7NU/PAvQdkADEEU6oOnJl933mWrErCk9nbbitH9R0cPL0MqdvoiuC
P5suJoG/29IrdNWctUqCM74L1IP3uCKR/fGHC/49UqH4QTjaL03h1EwzcYG/zSH/
iWSMs/76faCnxEfP8/hDZ+n4gZcKgfgkJp7rhyJHzJm9LrS/QQnH+j2mcB9A3q9+
t/xWHDQqa24gjEshyRPaCZ5qXhq5B2fEq1rrMGF+6s9RrEXlN9DWpKpEJYV/mm7n
xNeECvd2s3r2ODppvt+b17wxta5cVsfOyM+3Gxl9jKL+wAld6wbgNm5mxsEOINS6
1zolSpqhUlNJV2w7z9RNAbxVPiZbb26X47aybRQu3QMzGxhSW+c7nEXPjNDNuJh/
ltGk4xZy8a1zg3fN2O7lVFoI5pa7lEnnw00xUrQ1T813MQwyLAWca7THkFpJ1F33
5RmBDCbjumUw+2OwuRKGkL2sDXFxjTPaGvcTV6WEjNzw9VAgaJ1doKxXoK8tEKfB
7hMHOkMgA5zA95KHC+IPtfvNFnoopi6/9ya1u52XQAq7dR07WtwONPyd0kfqnq+r
5D6THM+z1+nHkaBevokUamcThkT+5K7weGVg1kIVR42CRpoMy75LqZAS5uw4ZS+1
ATta3upxNuIUX65ZWNvK6zuXXDoMWtKiuaVleJMlOsUbeYaBp17C3chWiKQI3tKd
qtq7mewZzr80ATvEHNXC+wxRoFaNGPIGrZRyYItVNzs0EgiiZoH4F6eQZXByZhSc
6G/X0rNCTLRNOGEX/Y4iDhNPNmrCTkaLbYGKUw0+I5e8YtFmihnYqz2dXh1u5mbu
O1M04IUhKP2dQnDDNKg1IXIm1tksVGeTmkpjY+UrQCtvgl2igAiXRZI8DH2UF5Dm
oNseb+XZxQynGJNAUgTF0XP8CT0CrAunIZCxVfj9a+BC4b2f7lJa0iF5U7YC8PSD
pbXNu6PHpmwdmM07RTostpFNt3VFha8/40lpIcAOwzvdpcYP1ryXLFq10EAyRGHk
Ccl4Z7U7eoL5h8Y+a6XOT15fxUXBpeeTh/RJOoKJGc8/fouUf5kAla3zOM3CzLE7
7SqG77OZZ+BaxiunQCyUxCK9CFMrwDcZ99c1ag0fy9NhCUv6SBkIACPO7dPTA08f
FI9RtrQB5FOvnti0Snh4csAsEeSP//UK59Mn/vKa1s56rp4vqS1d5hjBt5X1k8cQ
COHEsRz9ORNSLGo1jTESdCBD25+XLSRxNFWv78N+QXrhITQhjJN+XIStgU82FRH2
mJPjWA0IC7n0X3Kide5Ne6kl1X/tNkngTVnwzj7wx+h1XY9UOEqtLsDcyWFcK37Q
1tgBumBxSKZKz94D/ZwcawHEEjsxr7FO4YiklMPTOsPSkuaiu+kITIUIDvrk4HdG
vk9JWmaqqFOrewdyOl7f7r6nvrWrjYKtIh7wNj5GwF/KDdyu3c4s+tT4t3q3eXqi
43epfD8QzBySguqbLn9JfMNv7Jwd+c3grrJzOJK95cL/EMk6dVegIITOWN+cqK8g
OsCvVHPRG7IG6v5uvJ4rdLC9xA5KnVrNaMgQpc6X5Gi/OALjDWdA6nJCqi5Ad1K1
fpu4sQQbQ3PUrHqpXRm/EHqd368J6ZhLxaAVMmtAwzIle7cFfHNO4gsMkwmAFR6m
Lm/IJifDgYPIrfBG8Tf3TlDw+8hVEPbZRGqmQYc8MbbDXyGVMkTQ8Io9trVijETw
dbDmjpUfAQKvTSWMzBWQoTIDLmCfMKdk8cAg4uk4ktBCsm1JR01Lnn4oAQuQ3UHC
S2+Zt/0dYweZHD8tmFm7AV/HY/WpirAIpdgzo69i3om9MaZkMxyUeXIcaa1Wd9Mq
KCy6a+o04f8lSYlIPJs/v1/9XBfahH8SNagHV6VXGCCQbneuH6s9Ug6Io+ayw3Ui
mx5tpLq9MvbW5GSf1rr9jMRenRZL5RMqWZbqb4mVem70sjnWufY4TDYU/N6KSVx9
+ScmsegeLwzbATcx7NkjHbKE6o39A7e0K5xAQ0CkdPnR9GADjjgv0X70Plohebj9
+PMNcuS20emJ/004WBE1RXQyXMN2h7WLQCeNhQMsLf/HlJuKHAlcAvk1O8fWTw2/
WQgZcgFvtJiZ9bPja5p25Qe5qljjnKmDxhQBeNb6tqjx3pYGQERCmoHW/bBV4q8u
kOb6QJ7UCjnx0VO202Bb9t/47eTVjvcQnvSKD1US+LuXf/wthjhIbQxE7uyuT65U
yWD/qcF0h4XGTvC3abn4hjTCaYRIQQEHdam5Q1fpO4Rxj+xxvGX/lgfUYZlJeqAM
tsixltmcZ2Yx124jg7IwCbAWMDouD7c3/EDVaBdBtFQmnzE+NNGzb8rotNZwwayM
JMYJxkoKn0L6DaG5elmo/BCOKogaJ98EN6RQOnw0HIgsGlvmFuvFgF1TSd1oFYet
wNyWrhM2ue4wwNuTo+34DUUml/ARALQbLuFN2pyWpgBQbrfvKnjxjnYAtIW6iWeK
6S0M1S45siinHbADKPdPW6wq+CRlLZrGLpIMjDRzTmVtDK4Gjr7FSb1Zbn/5lJuW
7e8v1HA0J3y6qSeOA2hiZEztoeQoP8ITRZY/ZHE/EOO+SUKOsU5P7bQ6cKhuxToD
MmPuAJHJMd+w0D1DL3HE6TjZ7TuSmnfg3vraqsj5IyrTkb0ea3fnDbCClFZVVCJB
FUddClhETrtD/vGkzbWw37kTrB39AK3W5MmlvmE+2pZ0lXdlXMhd0rGCMLQCEqt7
RmZ6sG9pM12JKouB9l0WgPWO0+9e7b3MQtB3332b6ikdTf57h9StEHoTm6fHWhde
J/+RZJGvv/uK9E6lnMjN9OvDY+qK0QytNzm3DVwhYWAyOtrzPRJdkHs57MSbpt1a
9eOdPCz53UyWAFa9fQBwK3bR22k28hqYViFhMAqZ9hBphlb0hB7z9NpueoZHT1Oe
Onv5vvP9dKcqQSUxqxFQdnvC/B8Lt9rKDh8vk/69Yzu4ZqMs2JWL5IXTJFvNOny8
o4xb+ookZ8YX4lANDnPSMsWGv7osyYNcppNhn71I8KZCVaei1AJJ5Z81/YLZjEei
i2zgPSqurXmN55UsKTWCGbg7oGQjXatPCjB7qGOrcXRcbNyITP6ff9URn9vAwRgq
5ErGXn5aizS5nzk7U8peBQH08Uo5w5A7nI2c5cen2XGt12NiJFoM1VHKvTAHvaY3
ruqdX6bzQk7OET3/AL+6e86C/d06K4d3Ihjakql8hwPe1Yc9cOJnN58SSKjp0zXG
NRU6vs1I7kFzkemHEP0F22xOqM5ZxmMX7XZs6NVGMIjp1xSI5cNrqT44Oyh6R9eK
rVT9cPhBz0QXl9eTotBjOsn6Siyu+Wm4O9areRQvbsQHrrKds66at+liCYUthVTl
qn4GjgyoRT2TpHxsNUdqtqvSS5xlMWuwaq8KhY/jeXwvs9iD6kU7igkZDcWEjVF1
fgzxh2zOBZqKcIdAyqEaL9YmMabSHr4K9r+EW3iqM3ELtnBUZOEuXINj2TLV6qOy
8grm0pm3+0GIxfxjr5Z2VFfgHahONKiP/yWdlBez0G5pxx3XHKDvyLnamYIUS2AX
PDMSF0whSe9aSdyUI4AHZG/54sv5DkrYTB+RNhuKxWsqOjZgAkn8LGAdiUgeVIPa
Cq/Rgu/b1dy93W1nkqBzllo4fyogJBilRHle8fGSs4PZbUsEhIu+XS1qhgn+gJye
UuE+57YJ85G2FDt0f0D9JGkYwPT2ib3SFT3sIOyW4AvrFklLGKoxiHI/vnwEgvMV
61TSy8dgjI1SFYX4aQkIeNgpA+XVYm6G2DwEeElE3Pcdkmmr5z0vdMInBJ+P+tOX
/CEloGPwgFwU+VTCDdIWAH6GuCv+ZRiAI/OqJ+SF35r0adsQW+EeogfhtZHIRsks
CMN5gb1l0NXJUIkO++UGPlxoUeFUJQacf2Og5vshZCd/eAWa0ro+gmwd67QQqF3G
sO36k5ypnJ027sdMVs8XlXjPmYdIRaSZn2Srlo0FrydV4F4tzku5xNHBQrK9fAmR
F8EMkfU+Bo+kHpGW0KVd2oCYb1d7wCxlZdk6xZh/04/IFRPQMj3mlz9i7Z0vStfC
XDj/kn3VIhiL/YNZeANki0Emwci+GooUQTCMyv6jPPbMi5rsfCzFdJVlWAsgsMdT
Vb8aIy0QEEYJDGqv9T9UcyLFw9jJOxFFvcZuTOpJz4whekoL9eEdeEtRbNWsqaOV
K0MwlEO8/r5Olgge98UVD7nawufE/PLsHSTyKQ2iDhiOAm75r+nOFNCwS2aKaIoN
uPNP+7IY1zMvjNrXnWL2/uynVtU/uFMRCfnA+kINIKTg8vowfcCPLAhv8Rpxsnuc
CMk+tdD1bHCAdDhzw+t092Mmldx4kcQrfRecNIqkKalsX3oYw71WjVqaSEfdDS3C
1T5hV4hrAjNQrehCYp1xOEzzSK85NrPpQyqq8OJRETFiPHTh8JD2G0jVz8pAtmeH
JPR49xlNPSXWfMEZRlyl6cL7N3rA/q3MVu3gwH3GcW9G93iCIZXnHY6kXWun7rKm
C9C2sIsQRdLZoG3kMZjjFptdrvMuVUcXnP8hckdXoyBPQ1AEUqBkHJ8ugcscp1ee
HvrqvXYx1Pk14Ma5yAYmMoQY3M3ujGTVGp5wDhbdu1XCuSHL4n5wtLDzXpAaz5UH
xBnYPiN/Lfc3Hoz0a456ffKbc6+fp/DiMbN5+y7elF6OMdWWvosMcrWi6Q/25Lky
TMXEzTc1QHxQ8yYdCSC6h2Xyn9Xa+qmWXIsBiItehgW6MTdCJXjqd1RDE25scxeI
h3B/592gqyCgq8NYBbJ0J70fJ2LdKMnmYYpLj2Ks1C1/gXi5QbIeMMLN5ZcuWyl9
chNJIuO2PL+UklR8OqZAkUrFGBahH97j+gIUq2A71MkJJ/U6SVr4CITChe//K/Cj
5YIp0Y/pxy2TwgVUmj7K4IwbHWzj8ZWqkwFajuunERxKCYjPfhqvw9K//wJd8JDo
hyfsKgZ3TmtNppxZlie6p3B9bVxQH3hJ05Nx4QJ7+qWAZ65sDX8H7u1W9Akm0Xi8
1ic0SKQQIp/e4htLH+/T7qodPgU90FgP8qT3yfwEcTr/LR71EyonbkHtEDVlFLDq
HDmDYQlvztT5wbxoC0+rezLLeATgadtXNAqM/QYFWCSziwJutzO17M9xowdsckv5
dRgbFBNVzrjvMWwzTV0L18zrmT8+STyTXzo7XPRli+C2gcgOC0ONtZsUSn0JYE0D
lo9JfJ1FEEY75r0GvnDI+0YTdoKPJpj5SOhkDojxUuFjdeTd7s/nmJF/y0vbOnux
euxUoCxrPH5ZH/F+MEG8V60kj8++YQ5+Bs875O+jchchIYwFP0mEG9807JcHstTV
c4uuH3eapggWNdSnzt9SrsiQiR0YhoKp2vLFxUK1a0687/VIaFIvgSlcsKqhjRYj
RFkz3r1ai9woJi4hcm4p6fvF7rTfpqClJsbz6XMiJgCx1w/LClDwobw0/Fb0aiQb
4V4luWSkPpiuKS8dBogISqzdPYjmP6CVP6LZylfm+VSOZgz8BxjzO+7vx7DJ/yzE
zYgtnSmv9JuJR158PBlL1UW+h2QF9x8oudmKWfOryuDpZkygDD4hWqCaBi7SWqOM
+ZRua9Tpk5+7YkA7DybVVKIhTLHl9gIcgpSDxZEVIx8L4s1aeErRKMsoE3InV94A
e6qfqByPSVno90NYGFv2EiQNJzqc+9Ye1SEmwM2MyKQ3+RndlymnuRwmtYOnT3ud
ljH2cLCxtYINmSIFoe4PkZiL3Eit3pCGIyX1qi/Yz2vmBu9c7f+7JKEhVQpxOuSI
UXoNDLR+GmYFeuQKHaSV3uEww6yWRBhGUMatDlh/6PhFgtkzy3ZWJZi04RM0JTGU
dB+Extiz+ro6csYnYpykxXqqSQvJH1ISTKdgg5GuLU3Froj2LBfkE+oz8GEJVNiY
5dbvzu+ivuDGkMsJbDKMtdtyB1ErY3oJPZcYk7S/KfwigtnU8PjbOgUAoGuV9ffK
kUZJqfWimtKNzza/qFQky3iR8R30cI2AgduRFLxzvI4nBxYHDIqWPqCyARs78RLO
CyBuTTcDRy1r+KcHay6rHMTW+3676Doe2K2zAo0lDW5+HeUrJcl+qhv/CjUgE/9h
2KllbZr3QRUuwWhIT3Ja6+m3FlP+WqIjUOH4rPNTdZTxAgmITn8hFGDOt28BVkly
QSuIWnQIFB1QT+KJGTwXn3xza9ML4BYhSqeRZuDiCiehZk6YqybJbUdDuJGWTYuM
S5WZ46CeP7GwoNAyNTZIvbGMR5oGYKFbizXKymubKDA0Xu2DOuXmIj/JKb1LwW9j
g9LAAmikDbbW0QFh+pKegxh/almDdJI+EjMaki9Dj4cPLpfvNGp7QT1LTEX3wOOe
XdeFfvpCCTvTUkdI4Jk0Z0u7XVWqtXrt7bi1sMpyZnvOi2jFnLYFI9PDAf97U2TU
uTO2iXbvvO9MW4ZQm9PFaMS/P/uFE+467kUMzTKhsmO7q1zxDoQjNis4bVGh+QWr
JUHW7bOqZqigFEp7raehKHQCqNC7fIq216T7bbM8AeUE1JOEUy1KqA+Www2bf5Ny
RTnlSqaupMskkQ9ySspH6hehwS8erMOm6gsnaam/zMfs2KGyfAqpNK7wQo3b4bsi
Xi5kQ8esboByI9hI5whnY7bNFScTNPIBV8xXKZl9J38BaJwooHVO9r6BM91Qk8qm
iRtZpTCDYHa9EAD1alolUH/uWsQzJwC4ZGUBAzOW0SazTlAuzz15mN0L1mVytXI+
CdQAKHmuFDRfUx08LATTw0OeRnIAGDq0yovfztdrKWjOa1IKeDxn/RAStSx98toS
vHQh8/Pn1U+IXIbA5K6dTsHXtQEWFYmMtvaVK8U11X3KmbsSjbBwDP2/1mQxYZlS
G4+3rHIE4qDlOh8w29jBrzdrqz89WWm3colcFg/TiMaA11/Low+tSgVpVeXd9lSX
0r4cr2hyqOkHP36wpx9AYNxZPRAT0VMaBgaZptUJajrgp00JFsVEEA07wA388ugS
bKghK45vMA4GrvLWpBDkar36giD186Os5jCxdM7OqKW70F5/J8QrPxV1Iy/MJNit
cZXnras47UlTQ7wbkPCZaL3V8gDCmQPT1nWqQY/+MlPjchyn5z4QGs0KXtoKv8yp
Sw64EhtcEohsqNEVjEAuKJXY7Y8mrABMM/kbBN++ECinCqFpDsZoE/PaRn2ku3+Z
8DsEvD/bhh33/jJA9c8xW06hoXX+kVuLFkqdUeEm7D61VFXFeLTIHSAJrBMloVKj
mS+SnPbOxz2+h30pgK8Dk/KQSasF+zNb6oOFeDnXz/wiKPSxzIbxLCw+b5rs2giF
1vf7Xi3iXUvHhwHPc0wh8BjoAoU23jwdyLHxmV1gmE2rNWYbjYscCJWDdBiezmFj
Ed52E4Rsio6W+4aEkkDwsYo/3loIp/GsEPw/ny0uSE5QjzfRxNspT2OAJyaxnLey
ggoRd4mTMP3nYXryCZ7FVxhBoXyo/YqW5op6bdl08YABy5xg1SdF1Y7nStGZym9t
Vzg86QZOzQ072yY/1XSCmkpFgb7ztAtDmLtDFoaG5vTz1ChJj61gKKk43ZqqUXKs
Hragz2nQvZ+bEWblzbUeImM0dTRBBv6GBYJOsfo7dJ07thsACLZBe5BwGCjXPLGT
GsgYI84ZrAw7K8Fhz9cCuLkaOPjgHzC9ZUBLp6OEUJ2LSykBTAE99cQVm1SA53RB
WzmcntkNhAlHllXgU1f3oNM8illGcP3Ax375PASQxNJJMJ9BPAbF510q9Qop8YDD
0R/8txALT6+XEv2ffxCKzTJ6moFjMGlPAIoSKzdm8RRX1EltIsP2HO+QBeOX+/xD
3yWK87ODT27wqrlnIjhNfJ5h3zl2bxcvtQo0sFNYg2bp9oOgSv7CEH9Kb0VyI+LS
zN24mV7jWyPDLmzQTHtKld1/DvM+K6Tu5diiuhQu3IWcrvAg5rrdTBC4+0hcggyj
5pHmnP/LGrjz9DzcCPIKaWTSKJzWTH/yyrR91cxWbs4UAQZeg73e986ILsuHswoT
xK2AfBYz4iz67L1Ju+UVvw50bHVffwfLiIoJ97pxgKjXL3DOpD6PO3mmsaFuG/8q
15lAy7huykc6KZgVjqY8FiU7ydM+z8RWFvtgQhW529SnU0CULB4ZBjFRzWYoUUyy
jNFwgFSweEvbXQUyyHCs0RFkTRXWHBCfVSCRx79LXGzlnB1/XuzjCNfZJbsJg2Xm
Px9ya0W4n7eeib03H41FxU9W8gAgSuVmJKUBJFEbXCohiMO9F4VmVoHZNepg2B1b
0w+G6fzpmmEcHIsi2aTjrRojSpwFhxGcUYElIVXgALDT/1OoNNLM/AFWgoUiGgd7
aJO7tXY9RerR3n8Ia7j7MOZGSEBMtQ3FNWo3L1DcPGH2ZKjieda+ifTyvAGnVmgN
wTX+AQZsnC8zJJDt1yyZ9/FHCxqL91kj2It6sVQkkNJajNE2d3GUz4DOMp/2pfwc
wCW5Iu5Yi++xKDiTg8soLjOvKcIVsKsIB8a61I5t2rYkiJdbNr4cLaj8l7ZMb4vO
Hm4ITC9hinFapkKiu9TGJq2NJX+LR4kKqsWr36SBzLSo6mXaGs4QJFzB4GnMXAec
06AbvQCzhfRimAhoE7IkJkrfwv9ZLuekvQ0HKo+x67HdiIk3nySi8gzoS2wkRNx1
S9LxkgTLVUTzNPre00RJdG7LqcqAQ6VZGS9KDaltRqLnVLWIMWrfvame+Do5IxIY
nFIefx++YewxXu01NLwEoTF/95CetiM90zKmmr33d7Nva0RZDQdy2bm4QJU6dpA5
Df0n1ZObO7DRg8THm3m6GZ+tFbNzD0AM26YwCYVYu1V9BiHkkT+/pxnL16GlyNdn
9FGf96wwCNl0bC+oZsNijOZL1bgVYb+cjagrkscuYaOf4sVn1Ssy815Yq6PGoTWa
xdVlyFuSvMQejlodzFfy8QsI+ebTdajhVvLc04ADbOKTBvMG4sySs+CrtyXI+z3G
xROtAbwfseRv/QRJp24lqDw3GLDKa/5qK12Rdexd7WGyaBLZmijf701v1DDoYtuU
P0eAf9XIsWHR783+ufDayCzHoyVQasy5Zpzv/5EKV0SxdFSjUkOzjgi93fE6r6G9
6kca2mzezxmCBS/zquzmJaPda4E8PD+Ta0gYxLlQdYZ2nm179+Z+hF4ORTFx/V8K
9COXVsLkF/wqAf8GZqmQ1U1DJ6OzK9yyekSVEmgVF59LULKAyJdZ7L2o0OEMJN5r
9PipviYmbSgyVUFPT4UI4WfPkzNOipjwxtkl10I6tXFrZTtWyoWPzvFkZzHvKFEB
fxdLbpAy2QBYwthpfHN/o4VwM3s3YKxxoHWoL2pvIbowuXKnuHvwlilHuBfntVe1
e4HjG6tFoOxPhmDo/XXqwE3t8qnMHeNDMeWiPDZcSWdf3eyUMj7Rq5vT7pzO3PAw
xRDSJx/pPi+XjlRG0aXigAVrpC8ezoa1omJaAzkuXKepBWZYwsalfPcRZYEAbJQy
seGKHiUsb5iWmWtaz5nmSxVVUwXwzI7DeFTVjllgVwaMpY+ymnITHkvg91CS2mNN
JCB4C3mE94izCUyBCE1QvhmCN24biymDun/al5432TUec505KUsVi6ZE2D1PRTp2
OTreSrbicckp/Eq9eGItiQRckv3K7kQ/MH0xHG39eghRncpECrMuGmZHAMmZC6Zt
rYE0FAiUYShPL6jMSqigihNijMDiZZqZZPIIlw3gza6xkhZxSrMaxKpzfgmJg00K
8V6ypKTNrxjVY6R/ulWA97cLuqF40yuX5SuKvzP4Iex1GqflKZYWgjVUN/Y2VP22
G4CEjkGfo4dqedRcQqJcRIUVVEIJwhI3K1wiLxFqpIJcGMgJZVJcVbUbMIRKwIrg
HCdBTTNMsVndbDZGi8zWK5HCSxFL9VUzZMqtm4Q9ENCjGGmsSxguOivHez9UwnE/
CXMRRRtH6J3NHE9dtJyoz88xA5crFirbLnEEMCXC+mTgXGoV94lCNzrTTb1sIwPg
xJo//1Uk68D2o0/Qnq9i5JBisns9S/PPKdwdNBsyTBTvPdPxU3QdMk7gVFndj+7b
ZWlNggcAMEGRCN8JuoedRhTzlk/jG1tc79xLTc7/MO92bjQBIL6+r+i4sjcBMEUS
XyycU7HTpKNAs5489HpI06V09fVdW2lwq+rVnJlJpYt6XjNmpsp5Vod8528P8IFV
akbme7X1DCHE7VYJPW6AKYglSZSHzCWRF9ghMUyTWzEZDIo5UdjEq5uT+smkErmE
ONxdN0UuOyydByUIm2q8rrwzBMFBJ9xFMGNnbMby9bAcNWx22EI4aF/our/XHM3Z
Gr7azIguGzZpo0nExFQgEb/K/V6ah7q2BclNXsMuEHmMI/44zUboJu2471277ObP
/CveiHawipYK8TF6HYGMWgoq0XRYvt2d79Kywbw6+6MMWH8FK8EpOqZETd41Rlsn
oKDdJ/HEKATPGbKnNpGtglzgkg8KWLh7L6zaddwPEHOTcd7JaqnhTRuXExLSpAP0
nyPzifA+UWeaqKQ1nCw+A4fwT4KEQwHYRTjHOodjScRx3OpKmkaW799FLv9igv94
ePNKiHKXgStIXrDddFzMrLTuy1854XcLtL0AUDW+uabQs7npbvI5BLs+nNs4NEor
zNLiibHHnzN97rO9z2kfqx7ErgwjocO6TByi5DlEZ/5yFCwxBcJ8IhzCIX6K9+sV
5djoeDfOJtWDZRmHnRpB7TsDB6WkcazWT2O8sqRB41etH7VYS8EgjhnqV2zJamJF
dtpvkEACggBcdSjI2CfQKnWnJ9UAR3EF1z5yoTLhtcdAiC7WsmVYSPZTjVJsTavH
NkLcwJhrn9MuUz95oDY+/HrjvTcGyQ6itY8L+k7n2IEvz+g1qsKYmJ5ngNAC01Ji
nCnZg+h0In9Tv/hWAxTUA4vDMhBMPOqn6NwbvfYcOX/I+gq+cA3rfvtDZVa8Mp7o
K/mIJrlziT1fq2QmThcx/3mY8L5Yxt2rhCyA3rhwWPem6J4Am3stwBVOusYaJYZw
z/nJbdBX+NuBVvRLoQhhS/5wt1hAivM8Ya8YXTqQc4zSx4cJ/oIpw+NFaeUNqybs
4J6iU/CTXEqRpY7uaiFcmBNNKPmWvvs0N4pxkTGst/SRG7RihEq1m0t9uMEk6kNa
KNjfqSELuKogtqsvPzvWvhNAw0LKN1OFLQHH3LbKq7pyMYUJ6uLl8XbYI7W0v3qv
r+AZdPzxuyhTtm4l/HwBDQMjPC5n6V9nMZ8ZHBRIp9dE8peXD2TJpK05yeoFwT/9
6QXGK84uSGnxcOzXbQd2JSFtZX4ln3rldJF1/syPoOZKCxUZI6NeLu2mc2kPP2QF
Ep/7Vm9xPTxfsJRR3BfhkJ4gHFQEALXocfVMR3Urt1skKxw29jgKOvzT7Nd3AYdM
Usm6IJEIpj42ePxOxUlnifAsk80/HKEEQ9TzfswaazgrxzS8gF0R5/kgdPBoipyW
RqMDvVSbk/l38PNO0VKkjOT9WF6l1RVETjPNZUq/7J+pFmS44C0EhOek/RZTxluB
Zb3kevnxP7eKQeIuWzyspFxhovMzOINiChOXNcYx3JxYJqm6xKPMZZhk+hHEZUGV
rMDRYFy65ymSBLPJZK3fsy7GISETqjjpipTwaSsXJpxETVI+IQ/g7A+cF63cdtGO
fFZ6qUSuJLaZwenv04y0bCvG41ysBKAWRrONPe5kE+AlhIchP1NBTee7KUni3VQ6
6RHD/tacpGwVgLTS1A8cvBjEwbGPycrfZ+DRjjyCin+HvjC6yODlxUhw38a260Ab
s+0mBbLx0CqVnAJNDB787lm1hM/YHLB1UN9YGdVsPjDrlzePTxYrywf1yrLIoJqH
h26Rm3kaKj6Rf3wdPfavIZD9OG/rB254In26VCiijrniwNq60gmic9hLQFKqK532
fymGcDt2alrQBkH/Mr/xjl6xU1Oz2MlxB8U5lQS+lPjkeMlaCBM+jXA2C4EjyA8f
b923Rr3Xw1uCRwaZSHXH/lcWJNfV7/FfSaVn5guvdS9TgZ25IF6cA9AKKovDP6X+
EP/qjkPiXFJXe8oa5pud9pvUdEQ2GpDwJicQbPEcIzBVJ8ngEwIDbIGxTZ4grFL+
kC9UdSmUtYsMlukSVFpRC1L4uXYtKOGnbxC4DFqmtmvpEK4qwfjNQiKrn+7CkMnS
d4Pz01ErMtB+EUOj8DToocze3T519xN8mL3NTyZddl9KTqyxcgU9q7LnCHttajE7
rTLuWk1JLMZ7vO7gVHQbbfG6yeYl10jgBfSgADUzAueJK3q/0e5LkKRLm6IoKZJs
b5FzVUVcrGtYTtKwR+T0q2dbTJtegjLuhhl6o8JTFzwjmgQb3wzw33HgkQrd0VT3
7SGDD1sBcOuoC8Dd2z76g0yBNBddiHns8aD9iqOoYCTErR6+EVVV2M0VpO4soXc1
CrHJ4NM4oxnvhgR9eNryBgYBnvCnLQU88oUja0c7wa/VglTt1gAqxVgOoJdFW5bi
9FaiF6Z8AcSnLJoWc4OjNpSKHdkuVS09iA1zRpY0dAglOEyTfb/wMlQIacgUxo1f
OiT4GQkED3EmrLPEsgUL7Ja/bBw7mJDMASMTIW0arcwHU8La2kaH2znvm5VdcFWY
mCoKZeiwbBABYFSOY0NU91Hr0BIw6c6mZ1tRJ2zRPbzxK7p1bkY3Sl16bd6FBxe7
7PhD1Dz5JweMq8ZSBmtvP9UZVMhNYrp5S0PXizASKji/t8CtbGbHbHMX3tyvpmyk
ZfOrZtez8UIuGIQEhHlr+84tU8IWoM6M6276KyTKYsbfzHdO4njRft3SdVRbbQv4
yJts9S79BlVtm6rjqvPiQcFO4mUTDBLwxHveFm0S4PjQ09PSlPHm3ea7xvi5gquA
9+hkB1cnb0k7IidFZTGeSg2PTwGWDCfmbZKqj3KBIF6mZJxiBjbeDqddThSG4K15
ZDm0XCrXNFYS/SapQ++Ewqm2jWCSSQvXuL6suA7pvNCZYJkY56b+vMjosZp/vC/e
QQKrwUxQFxp4jnYexvgb1UXl2DmoSHR28aKvqcZYey/5PDE3v6nj8r4T72fz5P8u
66FCa5FdyUzarMC+9/6ta6VNgOiZO/hdllyF/fhTL9mEQvVZHhmfCuMnR0Uc5v6x
j0ru8RB4VrcKHlJziBmFbuHci0c+dOs0T2goAkuFwsIr1+WUlATGA3XV7qyTrRDr
TGn0JN9lXSenaqcjPeZ1xSMrkHtw+u/1DvjXAoFeFAoiBW5fQpljLy7YkKlbHndJ
9uM73TmDPrnY+pQJ7JUJJMvoM6djLd1faYRtmcEn0aOY1246I2Rft5hbmf02tVWa
3VMPRIgkSrOF8uZVdC9G49dpsV4kaVGmsnDRkL6aTsYLUn/2orOIKKS/FHdh6aRf
hFLNdn2xx20F+1+OR2xOKKms2/p1pXVsQRoSuS1jDQJP2gn8PK2v/uIkP3iLe1o8
pCd4rUBMs3HZq/Ug4HYl+cnZ/dJqGMCIXEP3kaXpLtlDOc6QuZAoF5GC62gqkv25
1zEVHPxwYW8z5FYs8LzxcmRMDYZKt9M/rQrMuug9BvP5J1dICbPoAJeD11225GLC
Tx+2wlVtMEznZ8Oc63PLoIG0sBY1U4711U9NkU9CnB8J0oRBYPJdyquItQbmvx+0
XiaSaDIrjGIFZhRB6um+cpEUSEfqkeiY3ZKW1OQG5r4LIIU/z3lZtvUb6UpgOnD1
mTSOhm0PKLFPR2n2pzonGjIrG9jqcsEZCz3mA07vUZHlJq5z+ioJbCERJd36R0Y2
dcfGl2fjTBy9dIXSp0uv+CiwutSeDF2jlfbihomAWfAtj458gNjZWEmNKuLyHHy9
/QdZqkiByI5Gm047gFC1+fsUDDPNcmovR6k5T86GOemIqY1Pa39gH+BiBewf31Xc
823MQQJG0YtKJ+dS2y6wnQMe0amZkVstQjlAkQE9z0vzEmHwJ5Q2puN2DQ95/jw0
6pgi1ujcmQf4N+u96U/lY0ICGX6zjo9cdfaEHwdCSvq5CMOG0MsnI8bhYUqeBXQR
Vp0TeY7HwWe+K//dqb5tiEEjb4mWDG+WBAebl+o9W+KtNwu4FTUgWmZ/c5mWfB1o
LW+UAkFzFtpqCKK8mBGGYOIB9v214VwY3f+/dp4zo3aO7MpD3yU4I4VB5buh/yB/
/QeZKVNan6vvfIbP/ZO8Ff07tI3IuL3NnVMPLpwB+QKN2MxJxPkzvYqvzVwh9T0H
ybjJGujA3bt9CYQ7qxCulnpqRvezIGIBUPSkZ8kskXWQKFfob9+e0YlgynKrpfh4
okhRkHkyzmVMtLmJUbKdt/rDscY9pa7D1hdQB1lKSAK1q50q6B0IzN7ziLwjwvCQ
3gBRL71qkwNWhHb4p8O811PJzOOyn5gt+orD0W60qkNV1fyurdyONB9Op0Pxcb6S
fvE8FCoFkNIR09vrMuUuYqDFUiTU8aWY8hs2PUAFGsC7l8f3Wz+4sdeldGkrYhrI
VWpaInaVZN7ovruk4scVy9bvj1DOjb98jHrst+qL8ReGvTcP5npKvK4wGR5G9Hs7
mhJ0YYObwCH49+6BdVnJtDKoZ/rM5AgtJEc+pcTABOYL/cYe7hlBuOm7Eo9KY2n+
f/Rw0aQAMpAeSimGz4KHUAThlfc7gLsp4KFyJESlXOHwpVmLISpjnMmifC06mx4T
BI8wZDu8rLdV2iot3ofyTl2hiE6p3OcdjDLK06aITz6arKwp74SQhp7kNTEyLuoo
8mwsEVkbX9HRbLkfh2YSaRPInd8kxrnkxeJbG3a/bx74+LlzItHdt1c8NhhnU6mG
yvBN0OTXCbc9rGg0yK6s7iW0ozds4s4sLxtGxJq4G29I3rt8GSKK34weyISbZWaj
Br2ZztKSeAaIy3zxs46lEk79ktg5Ky64mllmQN1VjKyjF1+phQ24App4lPXjBLsH
hC51t/H3acvQudhH0VawFCkhaPu2v94QkqQaaEeF5hmDXe09UUvqdre+9YZa/6ZJ
GPKxgF4+0Xsmc2QFHpkgypbkVH8C2abzH9EsBOdAarRM4gVXz2FS+q0USKydnaAj
yRytH6Jj/Jp3dvxQoKjXiSGszqxBK8vEzvt3DS36pAMpszAV7XG24aASItftbZY7
uf2FdDwuPZC0lnhNNc9zhyX76/fdyS9afYz0czuA5crwZELOxge09hcHRDPg7Awg
WKrW8GqZoK3prHLZqENcQjov4bh+yIQwBDWl86MJepkhgqyTuIqLJkji1ab0FdJZ
ayWzN4mZnSFLZLF8kR8LQpj5CQiM94ZKjo7krjanWixqBnvO0RxwLlycdKae1MqU
0X0D/EuwI09r2cRbMdXC7ZM1EGSIlCORYqvYDGheFrGrp6PTABVFuylQnPMszpoE
YOrGpBKlFhJjClk5ojS2UZ8on0Yb+j08RG04tRBYbi/0iguKIQzZfrwICUtVs2+D
zuZXOEM9Xc4i6CUPEG0WLn3mby31ZSg/YmwhtkshRShkLvPfZv7PV18gglx7M9ec
guhG65GqRSJ3QWCe9zGtOPHHAhOrjmg2mtDPMh8aiVp84JwkaHx3UW8ccbgMuBV2
pbpth9AvMxX7RvhUPmlM47k7o6kkx/jz9swIHaxb2dVEMd0gpYen5VFFiOiy7LMu
toUbZC6SnIQaM26oYuKphkzB8ixsxkt4+2HW6IZ8JEptt6wKeA+h5IbApbdu0KJx
P3M1UwVv7aocMWtktA34DL+puRkch3QML8e2aFbAjGOI8Jum1CnvvScdPPJ7cT84
IroCrK4M2yrI22xW2UZR+1hlCtTjb28SodBNHmdsCh+ZK0t+m8tHzSCfZyg253G/
AlanAjrWDibvcszRl9KLIAj7O5lZBgfUK5UvFolQhaZgaG4hd5MXAsTrzlCV5liW
+rcp01P+dXKoIJF8RP/T6/5ehSQfLvI2I9VqFNw8MfsCtgSwteAvdVnaI5jYI8NR
s4XTdBCzf1ZEYs6OlaZ5DaJfFid2zSVtxSj8gjVNxmGhrUPRvGXt4huGHmpC5ZiJ
foPsuCn2PZ0BBcJdxhNccMGim5rceuQu1OQhAAr1SZIzzIn3TpC/Wk2ecNh/IOVb
ga7nSGAXlROn8Pcn9k9EguJnJphr9351W9afi2Ze81TXNQxCBGeJ0DLt0v5QFm0Q
4SbCHI8HT+FH/KuTYgyjK1iH+umALgb8COkMKc0+wldwfCm5pYnA4Ruf7628Eq72
jX9Dw3flaXdnCKKu86ynZy9UKl6dxL5HGTcL0Wx8F5doiBSefQzdgCV7albJGFLZ
TG96biPAgpQcIaVPPkD3hx9NCaEXCTfnnlI8kZQOAduIrQ4E8U4kAf65Krh1abjr
WMYmRemh2LRlRW6hPS102zjjWbOMmzq+dgjRay83PWFiXevB/WPOqrvvMRXtbrrR
64TUOmD2gDXKMvqANuoLBTEmqfNkta1LfHoopmCGSSV7XxJjtS+n3/Q4tiIsIb3g
d3olUW53KeA7VZguHrEdIpO8RUZkqJEnFe0MKS/r1y76rrlqilegWuy9YTztrE5z
V73Mvj4mfuI/eQ21mJxYHuYdfns4AEdAI3WKJPyN/pXkQklbuY7qZoa31zutgXVM
p+IRTMZKbMeUJez4y7UTOK3DeVe0R32B8pXfM9DaHWv1/CyZT8JQSgnHYiny56ck
bg8TXv475uB+Gi+QHlkVIjRJ1jfnXduN743hteQxOgm7u3mB3Grp2zVjvXXmuLfb
OnB5FfQka+P/4nAJWY4invJVtO1Zi2tc57cLAYs3GlDWo3jIvKUq3fbGFCjpFS/7
YZG6+bhoGmvJIAUgkPxS7XuYmEp5UrBxVi4cuMXYTjn9c8HgSRfmhVAt38whnXQE
oHQF4HxLHcvgQZXusJ4BAUzegA+2wW5CECqDZ2qGM2IT8UNfEVDxdfxmiM81oHiO
vrmZL2V6sov/SUadSNYWnxAGubKNQgSLmnFFJkNWI7F8MGehXkyejHKWzuZme2tw
JDdG0jjirhQRo6cyHWomwUsQKW0RM3NrohyeDVw3l5p203ksP3E7DMHi87PMGB1m
cnT2gyq0zf4QeSlVZaPYQ9AP74hXmstww9mOCJrXmcuXfZ8jRwsJnoX9AHkPBh8X
eqGvmlezi3sfKA9QB8zMjhC83Iu6qNz3uWpAQr8qBG4G6YzgseKMcLKDYC4pQLjb
RimG7wF0kssx6gPBW4q8jgHBGgwnWK0gCWtAjGuXRxW5Kriz566rmS2jQdwu1StQ
KSWvT0tk+mhGFvSpsnTRmhTFmA9EFQw7nLQLfv2ZyULBADh+NhH9aFsYkPcUxsfm
dFyvS3bxorSyq3IF7GrNtNU8PA8byPRa/e6tS8lMGnQAwoaPEo7t2ERjfjEJnkbR
hqakvzfcaVjHw3G8Y3j4CEp+R69n/2s2XAFtmfokrqZlBWmQe15T3djy/b0q1DjQ
DQHf1E0hRlL3mVNvTtTpmW90HFuHCegaIZLy7G15y9vI33idvbA6XXsRawAkegTx
ZogdaH+6ivbwefVKWR3809Snp2n8/YZnQaYnx2EfF/if4NkSo47grucsQC7TIQgu
Z8CykFS8Dz8M+VDorD/C4/OfJQDHcJFjWRHz0+e8KZI4QXASyCz5B1xKwggsA5nr
FD+YF9GXCk6Rky+d3XSLF7D21p+/C5NK+J57L2LZXTiXmSkEOvZZyTMb4u0HzC7e
1SbSjPQ0FEZ1Lq4MQW3FI2MPnRIf2t2Re/LmvGZRJ2ehZhIwbdD+PiJf+yMf6tko
dnKxh65nL7VC8JnlPzDwGua2ao3pMUyu9md2rb4WytlpT814kdsOrgtLvdIsw0xv
PapfcvRV8/MwkykH1N80qUMNU5yrkg9TCQ8awM1avCwHwnzJxbbf/JQ6d5Y18UuO
OH0mLf6TP1qiJGS1iFyYGqvoTfk9RdBlZzIGEa+M2xs4tC88Y0o8jMtd4gMUby9G
0cyv0gDJ7lJxU/MIpW9g5lYoFyo4vfdk0W0cA98KOdHdFOgWc0wKQPjqU7n4PWiG
Az+ACWovWNO+N4X7SAlDHYkjyZm2DrbZEfWQ/xEspGDgMBosxradVTumMylcztOU
7/zfvJqwu2KBf+egfrbLY9s/rbRoR7g1U0ht3LFYHV1sjVTIew7FzoMEhloIAu7E
OfitdzcYUKVAMAbNSJeI0gc9Ay7dsbm2mvmt+CrhYegi4L4GgragAOhOeB1NE8F2
qqGbFz7lZfS7462cOYBOUjrxk+MUBz35hwMF87vZzp42rCOiur4yI+Xh8byglooA
+xxNmPbcv0BbFbCk3WCqTNUwqBf0bI5H4Kf3X8IqocbJc90IwaXPgJZaz8XNTp8s
W60Grsq/EAxz0FXsHHAwIWaQnjTiipLzgr3QN9UGaHazahEGAL94i1IKqpcOAXvm
4kAkZJV2G3doHck/ONY5rR3N2g8HDJ08li1Y8AjT9ksfhdGvnHdxoNw6PF/YQPLP
HfRiCVi2/T1zoKtotZoJxHd71BG6w0sCVUo52A32XYpNOdRFieAz8L7KZxJH+IW8
VXBRzGARPDF7X20BKEYEGr6i4sxD6VSJe9tbDxtU49QnmtfquTOQYAPvGI6L71kl
YWQYyZmtVU44eqsaMIvLD0u+UgbipguaqUebmjk0lrbQ+MbUD75XOocFdgm7ghTf
606D7J3YukSYa+bUujcS7XMNQ/K+MXAnMAkDqARrdh3BObbp9BrlzAzaXVUXetwK
htVwZHbOUHrxg1oiw9BTKVfeAjHXA150IMO7VMMzXYTRvSGwpounxxzqteUml9uo
nnBFZF7Q9JYw7qyeNajSG941j2lcERWi80p4ccw7m0b8EvpUyBNXv0ENuN3GKVYk
CblKVgTcu/I/IxqPScRzMHt9VQomCvtJTBndxWIHZHUnhSI7UottKPio1pyurZ0K
lOzpMAV1ee8uTGreHH5xUK+ZJw4Mu47UPlhCn/UPZzjCFQzKuMKbdj/kH2N1z7yS
YCBpIdfvs7pzLuhmMCd9/HZsyO5JW9g4MG/Vl6+9qLX3oZO4U0QXgpG0BHySPe1z
UIviQSqCCCXUViekFqNLIupuSthlX0diTztObt4/aASOAZ6jUK48yqo0c54sHeoL
w4FppjWMwK/fccfHGHRHRzfq2Z9WR6xX4yeg8/WPD8zvfqarQDNKJHjbTrpl/7k5
wrTJ7s+ECF1gf3CZiLl7BZDNQ9oQBhic5B5gq5Jhh/bE2FnzS0OSZzokbGSJrA3E
RejFVMkaE+gkP06/11MUscTI8v5/NRhiQN7uWmWqqc5G0hZyjQlTR2UkuWIb4g5c
VIgxWTa45L5Mg0YrsvcAwhAmJIAen9y7R3xFqh+7ptOgZ+rzIeBBHUopW3KfpfNI
yLOjp/mGyMh8s+Zmyo3uUfcXmOtrVPda+xrE+3HQ8D95vIEdmrIJ8gf4X5Jj8irE
4N+18ygvMzUbQDhdpzicty+M5xw3rjI9aBU7wWfDL7sp867XtNkvbmTLVRgzzJvN
3L35SNFDa3dnZ9W8qQKFVqyrneM3ISjZCUUEapURcOsFn5o4fnjQzrMP8U6kgaO0
g5Z4ugBJRMHS2UTb+2g6xO/jsVqRoLosTuk0wIs0FjgLM7CZV87OzaVeMl92dgkm
b+SZn+yVT1mtNlM58I2CiUnr20IhTFUyNPJE9r2Sc9boM3qNRsEhcQ2sh4p8cWIC
C6v7/yY3yAZ2Ja/WoLQ1EpYRRop+ItNcfNHVe2pvfSI6+cBqN8KkDhEXOqxJOnEn
G3EiPckRZK5k7Pr7O61TijHsQ970ckuZXrt5qHeA02GZ2kv3z75C4g+jyVdCr/Ek
xn/mVv2hMzHjcT7N3xDSraJK2HpPiBz3wyKVAY5B+50hFAH4f8woy0GAMsuuIzV9
bKUwJ2cXHagjJZg2gyTX7h31AeQgQkE8HjSHcWralJr+ciniIzvV9mwItPUi8K6h
BRKceakZ8hRbkdqS/PMV+Sl57KIPAyWYkHmOKBNUcdD+TX4+izCNK0+omUPnNDpf
N1myyYFRHbuL0e0GxTU8FA8UOQk9xxWBFA3IOQOQzENVWz+yBNtxQYY/O7KbeNCE
vJNY0+vGFevPinItSgs48TiJGvCtso+du3mk40FdIk1XH1pPPp1kuR5XnmCYmW5F
gYO5FBJ8gNFYG49d1CrKI5kbz7LAsjakqHs/AGI2wcd1RDUr/g56iDr6GOUxjb3n
WIFD5p9e7g7wlJ5XvgdSAw4vA7Dl9m1YOSyMlqI4zUbEA6iBhmhmmSyf2wO2O7qv
aoEiyIa8SqACL5oW+hgADmIYDdqASoYSl7j1k95bv63RHzf+VNrkqU48euvhz0nh
Z9jybc8fgwU/Oo7OZyyJSj6C+OrWdFzZxyXJDt3Jp8Xf1YdZ0OnAXBFblOzoA15s
xLmnumrSrovO5Sp1eK8CGjldJ9W5c5tBinUCRf1xDGsYzmbzqcHPVbAwi60jd3uh
I+giNwkv0q2oPn7L4o43w9a1IGbqG3hR54VohbtcHgnunqzf4ZIuwxNnlPIfXAby
+3ZKRg36I5n1PggImm2y9lAC9SAbs7rOYGx7gqczbgiUijFcCDGsQMjTZYZ8xZ3s
f4tHknsamfGpqAOUHL5Lf3n+YMf0pb7NVrPJfnEgw6Z8iFTwvYubscBm85lJRgjX
pCDpyHmD7VGwuTMh6NaAmZa7tBv5Nk1xwpmDYQRO5Ar9KMKZmaVE+pldRExEOstp
zEaFdzYCj01/tCJLpq6X6Jo+g+ZcWxoZKHOj63/lM2EGTQqbKDgXA8RwsPlqUGMP
64WN1FLcgZv8/b/Pkb6+t9GMNacNvg+fsQqtf1Nl1SyDljJxO3yIa+/XAm568QqK
qpGei6Ki39jGxa5Jn5aRyM5HrZayQQAvxIv0I4UzgFEHE9RTtPi5FZZKSRQij98A
Mt1cq+QFloDcqjO5R2HvHBFcZeLYwbmhEGssFXHfOVxgn2VzaJ4IZVw8HjsUKg65
tkdfiC3jLpWFOakk7leHk/+kIMSWKPjls9XvedsSSd3qzimzNLlcI3dTeJMDBInW
0JZo6FeRzc3qzFJ7JSTu7dy8Ij95wWzgzDQqwfcCI02QSli/pGhmebdIHR+aCVOk
rQMoC7dbA1yotgJbA6oOZx0tJWakuZxEg+viAY6TZ9jTbmOWCMNSh1y3gtAcaRlD
fDaBkw3cAUMl6/tDJEBIG+Q42F9f90PHwy2Xvfx2hTbSaxuFX11KyIcyVb89QxXF
9uHzv75cv7tsx7/D1YbPp0OdcRWWuNdp64H7Sc04GfnAnZSvAVZRsqZMEM1Wa0Sx
LIv0T+CMqD7uTIItwlgYszojBghQMIE876g7kGbiFqci9r9c4Mm844tgTyQLlVVv
AOnGSDEDTPZ0Q/qjsiR7RUO2/O3S+b6+zJYsCH7hzHB+P6kAyC7kIPTSXXRprgnP
5DijCIgsxs8iZAyz1Jw8Gy9yKCLR1Drb8DknlGvThOw1auTNsORJu15eyfoywId2
kkJ+2gikqKkaL+zS9FKQUt66RfsxtGIMwZxerXjtUbzZB/KEvx81OnUQTkr5Q9PN
a9tooG879IJhNeJbu1uvBsv2bKnTfq3xHSTqlSzuiRuhr2nA+zi9v6Jm/M7GdLD7
Z2JmWnnB9/5WNyAS6+n2pLdp1XOkM6zA016kDFU9CQXuzs3TCTulGj1qvHaVAJrv
hTA/7IDVH3crSgQaoDqstGamkwAuF/JBHmKjiO68BujMjJEybdCUbbKZnAJjqvhD
JA/fl6aodwUgrn+2yGxhmY7x7c6gKEvKt3dHOHVygsKw5/TTz6fRRxLf8IwkZyUa
iqi8AtYIyY+/K8QB2/N0ihxc7x1HWjXUwg+SSK0DURX/tGWV4pK17giH2z5UhQS2
XdORJEJSaMTXn86ZHU5D4wmVMSJBgCyOuxZPoIjd7KvPCi2UO7ccsJQplrBgo7KC
9MQTQp6x39KVnlUtzkZ7LRnYN3vJFcSiZW3sQFdMM8Jfy5y6Y07trnFHXoMHC+wm
tuAw9ZagmljsnFkTrYbC14VgtN/m/gObW0xn/v01NM8OGQ5BHjZMj574o+vMYnl3
ILEmkY4B2C9DFNfIsWBKw0Pd8BpK4//73b5tXMY6/c0le+T3AjrDO6GujFP4nSkq
yD6bYe1lDOajE3XZUJVv6g2+ChzNn5VjoQAe3iDrUtiiBpLlTB/GsvDi0SMUZ9XB
B6Qt8KD0ZqqZ2qJ9WGvuGRLJLwwyhi66eCgyNIL/PhlPvs8Z+kcKPrWLG7XyMXp3
Ej+Nq1L/e04GBMloQjrgra3xBrdYeJF050ausRE2onb3WOXooKKzfbZhDZMIybdS
Z9FNJvJrPVhja+CBL1EnGtib+Ffn4dIxREmnFRI27A6vjQGA2bVzqrtUrwiE5w7s
EU1qLWl0xRwwvPb7E3Xjd6RJfEE5/KQr+1lmZg+U6SHmzMthPqCNkNuE/SnUGa+U
QxC09OA6GZXiatsUWpVe6rpU1zun9rpLtjSNK/VRuwBcZBPEGMmxsP9m0pzIACeX
3qoHaxDUw4nO4mxxl8Rc9QLKZOBrJRn2WtjLQogoGAqASCLID7XUAgCOnsqJ/pDZ
6WoKSw4It6vjkytncard1fhLBAN9KIUuiTTWalptmcB7T1NARWs30CReZFtrRZpy
H8taPMPHte+cicaBAHIkgVBB3gDUAoTACTPJMJEctfKwgN7FLr41BcEaVdOS+Bq6
bsIKx6FqnymQsCU5YHzA3t+E3CunIykTOQHAcbO0TRDDyP1jQUM3LkDaJQ9aU9ZX
p8w0il2WhJ3brj5nHnM06zEN5g1xBb/h6q9et2tbBCSzsu7wHwf67KEgL14NkYWf
wEP4mCmFwgPwCsj3bIUT96pY5bKq8QuxJtmLTw6wkEjuzN+r4UsDrD85NHO4ngM0
tPq29oVKOH+7V5y9/NT6jtmprSA8y4ozICAs6hur7RAjT0qCBUQX60QZPdREfxcz
etLVYJSHg5zECoMDuu9yLqsg4hnfp1WWJ/vAfVwwf0dfigVS2KN9RyXcBNh90j4O
2NE83qgeE2vsAwOtWFppcAnzL4+xNVISEcY7jLCPj1GQNdT/A1IuZVMKqjRvh3qt
Sl96aG7ec9WrNYotFx1rBj7ETh2rpL0dGYvtocgEB/7NTBYfp8zqfiU5NuKxJpw2
zSQg98XU6OSE/1i9cvD/RiDIWVZhx2ixBXKl1TnJhlNuPXdnfuJX2lUFoQC+gZNO
rTLZbP9HZUmuFI9rWQgFX2+CmLzSDHT/0cjj78a89eoi9ViSChJ5TbQ27H49jnGG
2UobXzcHkMiUvrKP8WlTuGRa0U+CIWDd76N4GwIKr1ITPWHrnyRGDm2Ej1bf9zIR
KQ7QccV4ALQ7frfgqBi5HEjHDKWAGnWy62EpqbxZ8FoN9J+sKHZXVVXExjlQJP5h
m1SrqsSXVFonFOdOqAwHKbF8kbrnY4tRH43tbwdYCdOcpjgffIuC+hSR+oHjP7lw
KlfdLVw27tm9K89vnk+lDi0kTyAqPNDnRjaWJHCkuCA1TqZMMbsnlDYS20DskLzD
p/QNAsunI8K2Rg4EgJjvBNt9tXbWusPahi+ZvFebuM057G9poHyXopTUMmDvh5Ex
teZGjEHF2Ry1tXJc4zUdR0SumCDAU5fPahDMvLClzjkjBfwr1EwmIT6xM4XEUPtt
f4TvjEvh/0oSMmCxNBZsNWzdvV2zG//SxatWlWpSSf4gO7xlraUFjmyTJJPWvbjj
nHqHyrEP5xgLsjSsyttHjdrjijoKGpXhr1glei2vYqFuzzCalQa3BHAzuh8ZK9bz
ziSARlMKJGR8tzNZNc4tOH2wez/fj3Qb8S7uNu+sxBYTSfEME/gss0HQn2GY+HeF
XeGT7W4utEw5jIk8SXk+FA5riqp0eCD+tIICu11WJou1Hsp77fBbUkzIlcioi6DM
UpoKrZzCsL5Ccavq2Pmp4mJ4nqF1zpU76f5k5ISGvTNJf0V/pahjrjes4KtH970+
1wzF7H4AZhoCpAWbyHbUvlukHlembVAlepJs/sTbBgw7+bVdFx1qALguhAnLA6ay
1zxMOg/RV6FyZorifg0qUdZF9I4qlFHnZDX6XQ6iuMaHVgwE74oiemvj5CymVGfS
lgdfm6T/kyV5Q/ypI4FFTSfYEw68VnuvJtmm1xh2EkVuwvaVzUEPpgH5HXOjYV/d
RTpn7y3AX44nRUIOOgSBCHoPsVGrwx4vn0wocKaZ3L2S1Y9elQLzdatANSnqK3so
XkeQTuOXzGq7r5yST/W1d14qTUJoabKJ+E83PqsXdHAf8m5z5/H3GdXHfvErflDT
hpWruJrR5V/oP+m4S7K4jEbWWevm9M4AjPc9lyqImO9CAxFRp5p5j/bEudEX8O+0
bXb7PUBdemT9/65gkEZOhUJY4rnJXMGxwXauYl/MdhiPLdXmvuFH5PBqMjowKP/C
ZEoTALi1l+ATSDSNZXTsD/PofuvYO96eTQ2W24FC7Ul6HXpcDQ6FDcnXlbIplfX5
E92VJ8eBWFxIUK7JT6VuSKi0PW0qDw0icXhtntyPqOPYw6PnJNoXdqzb9chyAaEu
tIoPcdD0k0URP9R7hDdD05SLR0LSK4vKHeu2DhUjpbpsy/1+QAJeRe0RcMVkZkvw
NlIB1dkStVMlws2G19Dj9+e0qj3IWhMIFo/u0QIPQxdGhqpz5TRVtc/OdQrhWx5q
w1GCxX7bdLpVkKVc1qlUtAxJrFcabBRU641+09HK0i0bJFsLT7RT2ce1mFi44ZP6
NTfwS1aqVknOEHcuiSVjEHIMHdATy762p+17FMESGe915qWzY69xR4LjX2jUAtUT
QGFK3lI9W1ilgJEMXok6biIU4Fq4mQzI9HZhZ360y2NxctmB4VUixgLGAaJiiQd/
5UiHS55H3jNqa4e0WCgqGaq3AO2CjJQwjqfHkr8PmDtLxr3IIlP6GQVXN4UlTEo4
ttVp8cIMrKMHdOtQCbki5wXy5HokcfGswyoD/fXiTxEJwrkXEpeAjI+daE3L+PPT
dW4mvv2tfOA5b1cwXl/77VauUq4jT+U7RhmRnzvfEn2lIEG+r5MIsOuLmu1rqYXQ
d5lg1Z1rFArjru0tALbrj8C2UT1OzOeGdly7OOwhI7kMM8aoLcyV/Op+X3amGCsP
MQH6XIjiJsYZi1SGsdzpiKD0bJ/dnUkt5IGFI9GssWqUM/oo4iDgNp3fiCd3QcKI
n1TdIgnOVSHYuJLxqpOGBZCrnc8Q6T8rjKgeEMDJYIjK/7Q0qwcESfGPsZ6lj2Vk
gD+OMIbKdaiDV3gDFZe+V0M7krYHChSNI6XzEx7swZCDVvFQWTjRNVwu5XflCU/a
yaPyAOJ7YoJ27gWbUd2gI0xV09R9YC1xf45kIBFnKExFcRqanrrsyLk4BhOXW+C6
EFvTw7TyQ6wwEqepRmN+jMpYMvZdF3rOZhMNcYZjR8BzFPhUvrGeqzxeXvHDQfXz
Pvg/pxWQGJpo+53c3t3LcVnKFoMNWodO/pUMOf6Xga8cbADn78sZjBKgSCwCT37I
Xye9gajz5XaYEMn4t94TbR+o8mKydRLVZjuHowzlXzBaynemeP6uwTKzIviLa6h0
pFFqxN3NZLVYmt5n0JPdBJyrEQhMiVIHa9/B8LTnMGh6bp1AqB0twc+mWjrGBDgr
x/iowvgE3f5juBRwtl6M6g/CuG2YgGUCWZDAwtnlb2x6D0KmGNKBDZb+1dSWtmSw
A/QKzl/7rGxx+/gMk4+NhEIys32BxH1qlwMBOYXolXAnTfDthOwaAcg8YGJCdxGL
vh4lkG1QBD8bFD5y9jbq2t37rbaYTMpxe3g2fcFIm+KDGAFMcpVYIZ9sN1DkKxGl
XVzma6fGVtBDTuUPDF3vtZCb4hnmBz5wSkKi33eLiV42x/kdVfwBq2lS9e/MWE8J
LlG7MzS7oMLGjOdlv0pWUyiPMW/BD/1anamqAHroX1kV1F14GGgMOd6emDqQmtI3
PNOC5bZ80LHfxJ+SubDDIV29cNpTVw0/IWmQ/PXhqK6snqV0tpP98iJLCavhtFFY
v4sWpFckS9rJaafZmdu/gzdamoUrgWI+nX5hqaqIkvfJF9oZWlaT914gMAF+HmuZ
GycSK2Uamesizz9Hv7ODGfaaLnyWXRxiB+WwCWdN8kGsajqgEEJwWkehtUxJzJkF
+Vypijo5y6oA33phFSWuTR1xvS1Zl1oul93AlmuXDhNXc+2X0iFSQpEhJqZ6WMHV
t57Otf9R9Lw2I+6irzvMizw1RM7/GbbnANGT/9RIYyuZ+zprEqbKfrZMPlrFoZDh
y/eoZVZ2Cc6A8kCoj9LaemKhxmb2hYOWXhUa1o/3fSXJW7+38j3RkM6jIGseNeSK
tdtVFsWv6Kx5RmoRC763UKYkCwEIOlJJYLHWzqXcLU4uRwbuYTWmGkLySIX+1u9Z
TPjoewz+c2oqZfNkty1cLYBaFGcwL6PxBaq0jg2IZa/fUOMFTsKNjT6604CXMpRd
760jaCzhz9vjBn31r7UqPkNZ7GNEf9CcBrKIKSHCZIBBLdUXvzPMmwI65mf5wzVH
c2ypHKXPCPAQNOzjZIJ3HNi4pOWx28O+qffG89thvU3XjNPaeIC8hqavx3CkOFQm
afhKefF5Lc7IFXtgkD0qfAMXc4EssDOfqb333GL8qoGVtlxsREpR0UKtLPhN03EU
gkZlE8oh3z1EHNcb1A3qmW3iw5GZQZZ+AG1646/h7D1dFtX81GptXZ+ta21QVCjH
vJQ1VrqRynJxHk0slurMYgCm/IL2Hg3B25Of9jMkOy9oxmIj9MpxaUTZd9hTUfzA
mZfFyyMxXQspYE6R1+gV+SDrff7fGCo+Mh0K1E6ySJRt/9rhdqj+oie/KQY4yvdT
3rpsK35RNsK/npYIUBotkHvI7pn9ouXfAGUfqnf1nObJUBIhI5IODKKLglpN1sXE
OSUjC25xIXbvmpWpmkvzpSOPtRKod0vppQAcoa/PqVxq2S09BiCxd/MtYoYj+9wy
T0xh7WxRRxdOGFS3uETYqqR/jrKYXYz0xNV+kSRKEtBbXPjcgGz+JIszou/2XdaU
ptMG2xCdh96ahOW21qy5Kw7+tGMru0tJzrMGflvJKlHVGCY02NdDxwWLm/PgqJCU
uhVcGK2+Sv3d/flD5fh0Bwv8/PF4sWLoK/DrrDBHFlZgQ42ITF+ozCcWbD/3b3um
at/g9sVau42ZIJUbE7ubmv0Tii3RuhITPLl5av4yYzA3y6+erYjUHr/Bm/w26hoA
rnlHhzl1mmgnDaLaK0cpqZtjYSL2LzgUssXqVVmj5NjtSUaIJy9sJ7NYZ0E+YQvt
lrXL4O9lv5Off2iBOjg3XzUnvNJUiQ/57PAIksi03EhE5oM5I78cVKdC8UaCmLq8
BeDtKZjfcXfWwtr5E85UyQ8cqJ3GjdC/TDf0FF1BJ2jqBoeobnvYCliGFT6oLQvf
3ELp/RNVjWzRQb4Z+AH3NJrQFv/GJXA/mS7M2QA1HdFXcCeSZsTqYPqOUCZZ4z5S
qIrGzj3J8OcQoDsXRhKw+NXfLfixVPyT+QtVv9Lp/m8CAE8W9hTfb+HaGB02kLik
vdi3hUEN5FHpY4au3rlhzqkZ7dkY49SBW0trRtNd8JZDV1ae16WTTA8oTXWpm0Un
+UXAa/BOeUS3voMMd9jX3bzCETahzoUNJsv7Yean3fsG+Y5EKfHP6SSdE7W4I5I3
M1AhuI2lPYAlxUqpsDAwseAlgQJlkDIbH339NkzypvyIBOJOzp0VFRz7nHtaHEFA
3lBVIOzmqyymEAE5InUnSk48cN4aVoik0NyF3wVQ4Xe050x4X63spD+GTDpC4u5J
lsHSqgfutlHm1j8CnYwtdIgLKDzvC+BomJEw6WhkpdOBem2j7vbjnVwZ7c66Q0jh
XiUon4dep/TAZaUA0BAzxEg7SQQH/wH8rnWo+1pzq6fFz/nH1nZVFh3LIIolzBGE
vE5BWkx5F8aLRnFEmGVyWZvf9ockmcgnC7Xh5bLI6C/7rEtIsXk5E4ydzKMaHL7y
lOfVngw63Vi3L5aO9YCn2pBzV3cbALnUgB4ol3BmvwsZsgbAG8I6BEu/eeAqctrb
vMkD4Ckfi1VcjcTg7endjcdv+7y8Kbejjywy3MBekmIZp6mZW7comALnNGq0n1bX
d2d3g1tN3/0hPpCnS8g1X0RLBtoC2IXDHUah7jdIVEIjn+KBAkLTUVaxshaqLWWp
OU700FyBX9HgYGGdrPYnhRutpqdRQFKHoV+RDTmZumtRu1UOID5jPt/iT/PxxTTj
vV3jBXX10AZBLYvNgEs7G/U3bY96PZXyeb8zMioBLr0zKGh0uWvjNCMa62HkHs/A
65Qbvk7b5+G9Gi+EmOEhN+ApJcenneCxNJQUuxDH1uuju3ggk7EAXxXJXbmO6+RH
jXcLiqEMc2/8fR3cIcLo1Q05afIAH8AfPRqDv5LShA5Dpu3j6ncIxzkiEJTj43MF
wiaeH/hhXoyoBVsHqKWSdgk7C2FVyFgWP/jpGZUWGAteb3fIlp7N5MbzO5uakTav
aIRNfwQCteEdkkYskmxIzuotjAZB2CFlOm/KzShKnn5mRyIQccxXDaI22mv2u37R
FTboB5JY0fpLAOGqxBneyPhiNBxspvAb2lPGmrzZAsWrzrPxbiu53sRqNrM9GWsw
i6rMC/FhmFLyeasogO9W9HSyZy3YTF8xY7N2Uy48hYktgaPBNElM1dIebPbjpTOy
6kkMuJbUCEMmT0BNZ81B4A1EaGMjEN3uMX0sALZn6/mI4Z8e9xhm7mGoRMeMkttG
a4demrbY35O6wNpeH02Axb0CWnYdICs+FjZ0nh+XRZ5hJQeIhtqKI132KFKQXnoU
ZBmhbNRUOGRy6UwX7DzyJYoeqDUuwQn3CNxMTGC6Jt4HnKJbe13iMTTAxcK1J+ic
liWYiYTEqf4mqzi4J1El9BIRBqZL+C+A1R8KnmS+2ZfOnWkjFiRQUSmiCD0MSVe5
pPBDKy/1vuKIV5ANMi97XC0gZihT3ApK3JflkYvG/ApU1hj4MsT06x3RWMit6H3F
8Bcf9ImhDQOezcfWs99sn6OHLGg7aDgV1aCE+k0zglt2arwONG1woYH2hm6Lmqln
EbnlNbWOh68qiREiOPny+74KEEtiNGtSy9BRd28yxXNSj8jB7fyopS4BIJeOnENp
rNDxuo6YaBvTP2z/85gf1cFM7/QTjRpH+lfslJdm+c/Xgm19qzR4VdneWggttLlg
/6tBALmJz+7a2FwJ9/2KLs+w+W6oTYAJ9zUroneLcWWlV5gend4EDFvTe6UcaXwr
CjKnhUpsQBTVY+c4m//CxXIWqBvv10RVB50hTnd0ZCSggOxT52wqPPpRz7uflFfe
/5KdwgAlRmeEIx15PgwmSpkajami++UDQbjt4krWzC2cP6MHrMsPDiespwysUxN/
Xxi5lZqz9uqMlz7Svk7X+F8pjIr8aVq3zSSeSunPcXq+FQE7K8P+6YfjwJTZpI0+
tXkEl3toPI82Edi/7uT03HquXrs9LcvU/bxDvmy9S9hBkVLFETC57eitS2WBX708
JBwMeQrRAMmcMQxPoJLlUK6U7UuVtrb2EjqvYMa/Fv8K4ZLkuGwZ5uhaYqObxoCJ
cqO1A5VY+mJOR7MRSp66qVuRFyaJXnHqe6dgQFinV4zqsM/s77poTb2zXwGzJOM0
DkM4lw0A+LX71lk5NfuTjpVO3fN1D2ukxsb0dOakOBSSLXqRqWN8TaXL2s/QbQ11
Jp+EkELi8EFhZE2aHPO8+Nh/zTtqOvEa73/yvLmwmxyH5tVC6fkU2530oAuEJQhS
s7mB/48MfhWu2sOcc+IuTf18WTLbnTy+xmrTbGu4PeuillWHCQyg+LLkuI2seprV
kQu63ky5wtV/JdxyDlwkOhkyh2f/6yQJewp7nkMoaK0MK2yluiqd0bQBPXnH/UYj
8/Ms4M5ggSoGQ9N1DJni6/gzW8gni0IBQ/L7hWPzJxyo0VYjZNDxNlMVtW/7xYEk
IS+q5VJB0r5YJ3cBvsF4G7yAo5LhZlXuBZeR7UVyloM6qHpdIx+15jHtRv47NPEh
CrdT9nbDLKp+za8wrUV0M0ClT8rLOfLwMGQlgu45I9TKLYmGIFMJySawQfHPtBnU
FuNuYF864zZyecPp8hgVYBobdapD37Ta2bQ4xcmFkK9Rwcc3tTkRMueuNmulCUMu
wayl6dq7LzQQzCNEsONRrnOKmoZ8AtEQrKqPWS8HHh+KJTHKl1oFXfAHKDFAqDRI
D9ddzl60sLhncAVbFm5fuKsq91Im5k1ZI8m/BoqYFLp7mSY+MsJFE1Wg3yvoRSeg
5Q8LZel2AO+fpMQ9x3dV/ezK8q67xhvT/7uhdDc84Q+Fwjz2I6lodpYxgkgsNm1N
VJrsxJZO3U/g/K5D1M0okUbzY3EpRVcNKT6d2FTD5PhyxnoacjhN5sYFPlAjpPbk
nBJx4nGuSn23RMQtJ+NPAIQ2qQr+SSGQh9m2Wmw+FGxS+35xO/j7ZkxdTM7YzYkY
r8ocDjaPzjPd/3OcHuN/XhGN5s/1FYhIcGaBn4KgR2ekT04oRJ8aE+kPAG0gcei+
0Pn6YzR44OLu7BhYzL+dS+cq1kkXoPp+NrqjlVlTSuez/AS+13gs953wBCzgAuT8
VJ/Zbh+bMVt/tLQmEBCR/6H5RIy7C9zi7NDmyIowWUbLNT9TBP8Yf/0iItJb7hMU
iKH+ZC2RFLkUHmlrl362FG9VhLGmnUaVmL1By8xZylRawwJWUEp11BrMhmO2Zr83
Fk12NN/bjVxmtX0ubltH4gkX5Jh8qwPs9FMXe9B3lBiGIuhyRoxrUFFrI/94danM
8sbdLgDr2hzA4Y0Z82mg04IU6zqwBJK5Hj30FreScD1Ha6w8TSI0Msq9mUU78PQZ
WY2vsrqdzuGCb/v2yHMryErWnxKtt2LU62L2TwTuyopaf/l44kyl0cHFL0BfbaXP
Wpx6o43vq5B9E2cxllmC9bNLiWHeuRW9XZhTgE3cSuBXiWP8cyX9Wf8qlGLP9Dca
owsInz0MpY1c5+qeC7rulFxmt9fYKkqOr8kzNHqTsa/xq2vGs/PQguLgCRX5O7BP
oj+0tqlwIozZS2i8jyORkI6HgSA7WwpyxiM3dcis02WdNdSEjcySSXRpxMnVjxO0
ycNibalrZg7HXdx3UUQLMCNnJ7HfvO9LEM2+GrPSzRxDAJVmlgXXovrvc2LuIzbX
M2FR2lqTlW+ua4YnoPYVeCWwh4rGtjL/G2nD+uiv0Yu+mjbyqX9Ilij3kQRTri8C
H9ZkgI/ut44Usc1yDSDuSg2v2lVIQom7Wi7nlyUolTO62E8bI3XTmmFlTrP4QaH1
QnbaO2r+uEC+UT5fipBoE+0Ev2lIbELGtI0QoWi3ErF5AMOPup0LYLOwesC8iCsq
pGc0oH8K34+wrBVLRkEe8B+evJnPYhVMw35G5O9xufVgjVXLpAL5NP1PdTA/8j5A
SPHPi4GEyOTqdlduMs5iGNEWV9jSyn3XhUnDG3ET3gZmgkvSmJJU1haural9lh+w
/NxCQX9nLljfD86jgaAJnf7dASstp2HW24kRMh+QGuKgmNKoPd4wAF4SB189BDkv
WyVhb4+0pylt/qHDqcTWqRndgBw6qTFFxMjuzjz+urjehpe3b181GrHjE9/t8U2P
KVT/zZ7Eh6+Jtuot5EpiC8QGNxMoYdDm5SD9Nh7mnR32RGrG/BcyoujX/bnMelhw
PyxtrHJs4SbA9b+f1+HYIhGLb0rqtOhkQwxdeQrVDj/g/ZwFa7czWmKWph+YOgqn
zuj/IXGbHcmDCpqXVL00n+04UTIhtQM5mL/Ix5x3lr9I6ELgnWFplwPYIAW4apfI
cMx6rjid+q5fJ8bVTvnzjWqHuVuDrNMCdYj8u6UKbppRikvp+wpAx6z3h4NVftw3
bYZ/496m3b2HUG2bdT2w4+Og2F0As1hLWucDsxAqcm10dKZIOlADZ7E8RsvjSYFO
HypXRuFVyLuvIqdzNBuDWPzxzFHf3kC0vi2lSeQdQErekQCPFxp0JE08OH1fWCB+
S88RtorKi71IpFEAobW7cOtS1rKw42wm/27J3/+KiehPBvew7U1RIdFBT7RHBb95
JPEq/RLEvJgBW9V7vb5CPCpe/5b2LLeAdnp7+U+98d5uNz3wSWuG/RloAYqKRaYz
+TolSN/uvtkKNAnqMDf1obyJNv6fd2So9NV/S1UL4qd3tSMLFWGUbWqRbEb7Qrkg
KLcFYchEtQAFYe1Ig6YwHWCaSUSmvOKB4lUZN/PQXSgXX1mOafD0IlSQTTzCWULz
7ecmYhIPCoGPldxGfPvVDPBe0/EgT8eg1v+LLxfgDQeZOz1lZbeTALc95YbORxmw
+b0C2jZ94Mo3G+gGMfA+e0iz0Npj4UvUS3bFuD+JsTfnueRmVEkaiF9UQwmpJR4Z
9tesnQyECVpC6ruL2/zaOZtA224/sUx+FkLlOrXCIKphkfPeTa3uRF1xXmpFKDMM
Ojr0+thEWmneiS1NlXfxiWJskKHoDS3LZ7Ak22+EP1rvgvxMUYYg1mJcFzgb2A2/
wAeMZ21KGI7JYhLkMV2zypho9yGXRf0OnHU18SAnhZdUo4fEeSKWtysxSovLhvFK
Os4Q0s8GOFKnTgO2U4NzQ143vt0JZIFquQ34vIt1FeGQ1EeTKCrHqFVzLPICIzG6
Yd9dB8Ykqmk6c9hyjxaf4oAqIo6TgBPPxb5Cjq51RL/AVKK8Dkw04G4z+mYnyNZi
t+v8ksCiYaab/VSbQY12U/vxvbsZA9+OZh3VZppHjr07Op9moYRKeagj11GbogVV
QAHDFxk85KnsHtw7cOLwM86SNbVt/9XtgpTSHWKIc4vXoQ8ORjWHFcpk8HaxcmA2
0CNipByUonOfIWDgFMhTSFfT4pTdd8bANOJ0IWE/CaCENBXmurnPdb57et8eKM3p
oQPRHzAPQqqf6+1sPNRPEi0lcRvNazb0t1BeSgy36xfNJ6kFDITr1rR/3Y3OypaP
6eghNhATh1IzIP5NbQKNPyOqARCWnwc7UE39gPAf+QIoDZ2pQmb07TpyMQqBS8FD
uTCY8QIkY1zfamcp17mI+a/iyWan3VB7B52SG86jR1ehekcplR2JzqJciFuD2f1m
w2i01SHtLFwrUuwb0o3ib/QSnXkrr4w9rLSrJDMoqWpe2fWJiWilTFqz9WgXOifR
dFOR41KLpZAIKR9HwoIQ7Md/BLi98V5lyWTOydm00NQ2oj1XzlqlACC5wwB0YHKL
ouTGKjXmmTD3/6QVEAgtZGKQRrr7mExlJV38MdQoNBdvsFi6apkad/1ywjFpeDwh
SP6G09tmZLCUvDJMiWjGrOsjULtYUhkzR8ZEWOcsMeB9wSwLkwQ5+jc9GDlijQwj
X7iMXxKZaqoSiXvcXDtDuusojzWT+8CdMYDTEXh4tinMEfT+GCBSRNePRhwsiUwg
fL0uwDAQp3wAfmOdxZLOlFMTIANuO8uZ6/WSsdllCcg2rSFTmyjfPtTIYQh0IvUJ
f7i1zmw6puXuFH8aseU+r3Ki5aRwOr1I3tnBIhGrA1zR77pQs8tqljkWv33O8t/0
9TW+3rd4TxOORwTi/CntfIo58LM0QX6TwGv+yAoOK265mYv9slTKBl/oSFVQO1zY
JuPrHVATcH5Rt9E+A9omWe59vxR2tXJAu8/DCVhH7n9SJTT2aj643JNUpj7L7oYq
Xfcj+tNOr3WwcgHqYL5tfi9yJ8yoC835uuXN1qDiIuT8n1W9a+z4epWGWSnvJnpb
3PB9Ij+Cq56ygICfn2KyQtCDMthvogpiGK6znVC6XjDDnNTBxCv1/rdMM56SO6le
x8iTRgphF/gVd/oiZnFFk/YhlE/Nc+c7NNZeVh0iySldQS00pAPYjoTYl7jYJaqJ
l2ilnPMvVfcbb2+eGJLdY2sb10ecYl7WG93I7HY/DeyQAKKu3dNPu9n9a1msw5yx
LaVH5hrJQnP6DG37VqmxWoI7IxZrDSde6LbWqBjSHxzns8ThNo514EQW5EZXEmIK
0jxfwgt6nYmDrrVBVDgBGOc27nRCXHu8JhVvSegdnk/n8pkrvMHH6eCZFLNlptAU
of0sBoL5wio045dlPKVFuMlVru27woCAekWV9Ft5auvhN9v53iwtPnXmUIRMXb1f
1MnaBNMMn9PK/fm/I5C9OU/eKm7RZ5B4eHp2n2EO84pGbSIh3Hq67LVgcoQBaglW
aqWKDROxQOJXAnK1RZXUWvmAtvtiZCJ2NCwi4t3OtD0fleewXMOoqraFSzn0Q3um
4N4SJd6/edbuG6TBZz67Bq4htDL1WTYBgWPvtoMbMyKsYKmNp9IqtwOoWJOZfHZE
vglxOT5OB9uv22g/KDzpzlZTzvc+DA7iMUYqnu6pfNv6h/9JbMAWo8zxrlO0fEsn
bdW+LIahP1fxQ8XmdEHtBwmqyNjPaAID4tsZYGsPnyEjYJrxelJqTX1dz8rNkhw1
34ygzagFQd6aLy+DEuxps2JYoGFKmdjfYFu+qNV053AHvnNSDVI2w0hJMZ5HM9pl
DUfvblBnPmbiWtC53GGVkzoRP94hOAR8/ZcNzA3tNswG9pxGI3FUbGoqh5PYGI2w
wOZeVuskNgJFkGbkhRA/wrTih1UjtaIHSJqqEShwTSZiHhPQGphpKh4QmSdx0Cd7
bZQ4RRkMbNZE6/wNN869Lk1kTu1f9ouQPR2jOXIDy81gk/ixpOSHf3goEiX98D3z
NQo+ietLFRrP9t7u31sfQCblkZ6lw4iQqMLEHe6+9OtZ8ia4H3Kv68T3feqdNoJd
BuJRfc8zd89qFT3gh0DBF73ZNBv1pOOTJCbHnlmlNuEaEOdJNGh2PP/PLXe8qRWV
tOJI8qk+bSU30En90uwuQcf6l8iY382gzx67yZZ3WkQgPcO5BpczgiiQmbYTPOY1
7rD9UKXEGnujaTV2B+Ln1ift5MnOH3SKH240qzxmfMjilxhJ6+/5pwUFgLj6DI7J
/kx7flXsDVeIhqUwCDOzgVxRJ84ZRlhvfQNGppIEguFsQZQBLR9XKzelNrdQCFqH
lXYslFeU89Nva7BSELcyVl14Sk4l+8IiU07vM1kBQ4r9QlH1Nl8EFVzaR2FH79hi
fGPzjVK91Ls10VJ5rBES7v+Y4ggn4dtScB6SVktiNRdEwFW5r4S234PdNGyDYxwx
t/1C+MbOFevcK50gjGD6EfPZO44b9oxRXHHtfcm/aQoZQbej1RUfTxIKveZV3La8
UVf7CxXbR08WGu0sEAtNOWb5WRPJwirZC6jWHtSRKqLMpmQbA/is8kZBqjoqyQGt
ynxKJEQRFUVeKMoehrR/yR3IWDfmHXizOedb9WqF0ser68sJr3H4ka+8ChKC3qkZ
YWdDrIhLJCwO6Kx4KTAexBWaS87377uXasGyBbNZ2AkjjgPIyKeMminn7J2QRtq0
2upokg64on2K737uYwjnBu7Qk+PveHUTIMStaUwvJWwicXmbEBBXOTZqNCp0B74T
g2VTbZxWBZpqZx4OJQV/TJKEMyZ4TKmFt41iFp9TFYN4PYoNkJZGF5r8EHO3AwDM
n0mAqjpQ6KyzrrGKPAOTlF2MnAftpEfBiaAL7zWrep2VdPdY8RV1N54hYWWEmK4b
+R8YLOQA501wQQ40RtbMh0lWeAVIp6f5N722RyliTX2lhi+5cvC21N6q/cz2kuGB
txsLvR5dWehOy8tThkPQnTLMsbDU/XfLXGFrPorhOHedr0AMIVxnknJrxthAvMcM
R40pVEOQfQkqd02uqq4vByXhoqf70MfszYryLHJVHYdTBcsqRMGkA3qtijQ68IfV
7ZAfSmPTdmENtctIgmsjh0O7ZmkfVJPfex3LY/r9GPWgvUDoUHu15XTvpSiWD7mb
AFJe0HLAMH7sQMBJAf0282dxDaLgzOukjROVHu1sgnp4jw1a8TwWYrP46aJYeruP
ktOB5GHWAOAGr1l/zrTZtT6GzqoRKdZgo1QSxaLERmKe5EYqcUbSPBli+j6wdc0P
xKNxncwtDMxeZAfWHIDYI7dqQYDBk3rGhSrGhP9lZDXrLQjDl7sPicRd6WmH1dr7
uuoHlQIKNKTHWHVgog0K4575NXYnUa+f1YUq8E68QkcM7QfOlX8XpPjgV1q/UWo1
doEHcGpuatUHUg0lJyf/YTnGUR2YmdNQnetq2FpuUjFcMmg0eMDSAZ0qAAXcWkk3
rKv8FEf7EzPObBYUtIqpqgt+YpNQ01oe7enGC+52670bEdNbHSLZf1N5umy1sx3n
DSKsPYPlwrRVNwwd2J+aoliNIzt4/oKO24wBU4/qzvqzYW0qINVU0a1FoQy/J7bJ
Kr1glHTQMCrDCM9uPTJlMq4NxGo9P5xdGUtKRrbcH9X1vBgp7BeBWJNRGtar2kDI
mwk5fi/ICNT9OCbnKmuS0+G1hEJ+37sZIorHnCrpTq3UQVCU9jGk+Y2Nhv8f9Cum
ofvCHA/JHWra9JS7P+g2e6JMPj0a9tpMNsQCUhdGJ5bOOYtYWtwZ46YEACp8eVhi
fR09aNFnS6HIZEyjzBZjy8G0oSnIDlVfA7Kv64mA1Ws2GE7qAhLTGhOCMcVgz4rm
ByDcHyqSt/hzBgO0/v+uS20lcGqr8QFLXZCh/gmsXnRKphLYFKrCs4h9uHJGvBNW
V2Ow9aNyyhWWSEt17i916Bqbc8WJcYobmbdeeU+rRU3cE8nIBDxTsIRIt09D74pV
RoagSqwZ6zcsnxpru6Rwcihvw/q3isPNAoWsinmlCnFG34c/SmEeonTYMn+HBPbl
+aKSEAbREhFFpN96l1xYDBBCJsMtNXqkvum+SyRTcn3ZHb48dbEICfwL3FPyZr4z
3JWcx51f0epxrH9LK2hLUoVF1PleD0+DxOOIUGmMQpNheIMYI0uZ+E7F6f2pm0m8
cCWqAqEz7k1Q3PgTerBOPVMwPkLdPmDjWjLcSnmeeUBc2H7m+K3G9PGJh5+MP4UD
YQ5IM0nDEMeaiBh/aBwDJXvYbXPKUS+uUTF6OBT/RLjUsGOiDzRuiPuj/wffOuPl
YZ1ZImQXleyQhAh28sUDRhUZsXAc3j0xt3nbi8V1KyEEmrvmEn8fYbqFTS2HFbYC
2BURZxMmuZaLlgoCFznX30gMHAkW+Jh7YoWsbobJ7MJIt+EdIv1wGsozfbLg8zJB
OJuWfwEx3b+zLozNVuQJG/fvXo8IdMbgVGH8ty6Pqg2qMc+UvUyd4myY8eKUaQVa
nJal8MH0AGEzwDbOMcFo+WA80JI+4Y9EyGDrUrcaF98nok8x1jemZn0gLD8nueA9
/R6k5o9XWWNGlkNRbaED2DO9/fsi+HNErowJQG7UraTlX+1uAJriyM+yJYgdz6Yz
AGLlADgNFcM0nblzaAG9amqlVRz7r+XZ9IhAcPYMWOfnMsDxZ9nUNfG14svudTyS
gxpV+JSqxJqpkbzFcxJmymDGXFcKyUenaLfw52Bs8vYQtUf2mWByx44K6qN1RXe4
b5OGOkChTShdN4F1M0jMemj/mkiEO6AWgUBZKn654o/F6t+RXT1zGey3Row+3Gw+
CeJqX+xZ1pag2yLrfiZ3ooHbgk/VvkEX/DxvZnGheWY+tQyreczV4qhgPgR1k78Q
3Bk/folrDNX8Q4DlqCq3s7X0eAd2yTLvYfNa52wWvROyoTy/9QuWYxoveTMyroVn
grk/FbXTmT7ZhbKldzEcbfgy2cjLmm4g3/AakZ/Ta0QU0qMg7eBcEI/3zgbaNhaj
oNR4P6FWf83t8C3H7BC8K6TSoTQoZGVUDfEvtsHYy/E81OKAF88dZCO59l9RQD4a
prAxYsIV9MAI3ZufbLryHSvWqXskGMPL/yx6bTrErPBvTuiJ3roa2uvTqABADf7i
kdStxMrGdK2QhAeROM0Ba6KWPKZD8EMu6yCBrw5iZW0hHuu4kJARMgPLSvROfTXb
XpervNLCSwPMZlc3RdtckIPGXbtaDRPwUWo3vw1VCXyKMvibmautYQKsnsRDYI9h
NCORLCKYSm6uOTvHKcl+Im4I9fQ7TfhkN9qywa9loC/gOKIefjq1CcLcePQgWCM4
0q+sW45LBSL2nzT7rBNkADjoq12Bw4v1T+kP3bjGmi2cGkkFXfRZP3I5jp19pRvo
O6IkDn41YP0XgD2Mqpg/WGoTfsCEZePUa7yuDdqHdPMjewumY+c95bW1lbJNo3jD
/wz2kzp9YMHTwJgQrqpAy3dJDe0xvDjBFLZ7rgw7kODvBEYfwlhkWhA0fpMWNEb7
2iV8q3WfOVcsdhvKmglouE7zqhDbkElyyc47DMfZwP+lEJgxwm66hYSmoMhoMfvL
jmaDyG67YuxrNxic6vrNr13CU6iD7gbjLIlTXcRnIxJj+hhe1KLjI2U64xg1gyii
ps+BdQeB92JIZf6sMqXx8GetDk5U2npH91KbnB/ItHQLK/v+NYf4bjV8GyGTmpJV
aLi5LZ8Zud8fNVEOe63PuJJOCKzl1LqL1EBr5xCR8Qxn0vZzxzvxFDmVb8r9vKjc
W7gFNJFLQ12Fqs9c9uHQhBTDaXEBrvtYI0RULUlZsp45lD2oZKCLfPZjr1+Bf2QH
lb2E3XhHHj9Czoe/plllU4P+Ate0MXoinfu34EV3z0y94L3y++XqVShc13YQPUy0
kqKPo7bYk8PYK2aLaFCIEs4zSxVlFm55U9z2GvjHA7MNytOhUlJeLmtsj445M2bo
JD8kFvx6brT4DvPlGCj450i4I22r31dJktoatu5pcLJ/Pyiz4+YtPiZ4AtUGsSAo
eCj6IHmaF/32eXZjzHhgY4EXu4q3/F67QCv6nhEdAam+wsjEwaXo5yObPxSatBCn
RvM0AOiTujb5WuMa4MBL6uMDNMswXUj1Fkd/s6ku9YIk8u1rSXpOkj7XA29WOKSO
MTPjEHb5hJrCdWZvvUBV+NtgMWyvq1G4MZxWP69DBc3vSP7Bt/zl/SO6NSOO8d16
NHah8726vO6iCZKgixX7qBnsqRtM3JRtP9xtC6wYDVrtzM+C4JELIu/uO+VxH3pJ
MS+eE8JI2nlpwm4AuVwFS6V/dwMQTgzt3GP5WLXDEdKfZMZzmO8eL+ve6Gzn2W73
fa2+kYAsHg2K0LjIaxzgZ7dNXN2VlxTGS3Dk/u3GDBQumlozdhY2R4TUEuppG26X
+d/sj71zZXLkFHACO2Jaj8wMwPa9eBFSrDqzgT+xh0z+r9Od9AaCmJfvXxXBW3e0
joYTxlWKugni2qyYKzoxP87rCDdfNShkoAnanyUn/fY0QEKInCuqaY/Lb6bXx+HW
qm2+Ilcq2J3xiGKlQ6pYwJnJpYoiSH26DzDnxKKJVZ06849l9MfuUQw88GB2qmCz
M/dB9n0h2ilcImpOdsCMWvkjTGfMNZ5SJ5xnbtWsJ57giB0PfWNUNU3vJjvbRcko
8rDlsScpwNkZni6tJbWl6SfBegWMDH+OUES9CSwsiLX9sATjqlKqMnjhN3NlTDou
4647eitMrq3n0T7dyrraqInBtTgDvUtDyUDwJMhWpscIXcto8+wAb++hU1eyRs3k
fn74GnfeGxZdn+VHtksXQ+8jXcfHmPoGMRONxG96h5xU7ipbYJ1Y84h+U2n69j3O
ED+FNv2KdP6miwcxDTDEkM7LfwjkIBfzJtFOKUyC+p/Im+7WZ4R7Wco3kQY22KJN
xSTfOGl+pD97smeNiCaxvWAxuaNx86MIxhUg0M72G49vOSCJ0dhXCN2SUeoBJIFN
6Mu0iUNHyfs4yje0WWEXvBkWiO1FsEy2heJgf+C3LJbn+H6XWfMAkXaLUbBu2WEL
10dlbm2bdruPxXkkxIs8rvdY/EtXCVCLxwnsYxG8aCfVNBqmh8paCjvW8f1KmYsC
qC8mgg9DyoyKfaGo9yHKDdkD5fjYFOvSF69EXUWeACTAKfBfutPY871UhCjzEgOH
NA+iPSQF/bai/Egld/T7XqDerdRLsYHPuScxZYG9zN4iCEmiLaiXFXpvBHeUjgO8
TQ4cWm2siOEbL1l7nJXrMPhQW9hetUp9E0fET/uEm8/HpacpCzD1cWJszuoIWcSK
B/ZKhV4dtXcSq7PqK778ypK2tpZIuKTTBm75zQuw/KCxnKP+a/P54VqoOFM4yUWV
QxRG8Q7yHdSdqBAjNRq21xqNL7H7c44GbklEVnSTmSNJzwStyHEaIM3YlQmjH8No
QRA4P4HcA5Trqio+y3B+1vWhsrlpZGyqJ1qlVyYLzZwss0dya358xAKkwhhxb670
2BqsN6RdaYNEgJlidTR2Hu5yvRWMuq1bQrE/KTcwjt1qlHjFGza1em6IRAb8PTrD
EhJbiJGj6ZnnTNqVpLnihUfTPVemHxHmT2cJMlxRTTobwWINA3oOaRicLmJ0REnp
hgKeHZZ3RI8QaSVEIbeQnhcny4sn/1KWo9PGdNn6NcMy6Vu7TGaq6yGH9Z5fMC4W
rCYy5n5scN672wpyxs13meAvb9e9cJvBIlevt6jBxWyq87rXjZyAAG+Wc93hfZG0
G2Z3qyRKhQA9qgMQmky/8O4hNqCE9DF1ZxvEq2lf/3YsHa5i8usOj76J/cJVya1o
8VSVLMkZTnaMV73RV4sW+f3H33Sd3SQK+ihsEPjLYqCR+ASDzH25QDszUsWyq4Yj
Gl/h/q7ZoTmn7NglJcorHjG+p9JTAjgDMcjm6CCs6gk56AIAVH7i3jDlW9SlFu2Y
mLU+gzuPjPn6JREojGcrRzm2IQrgOTEip7E0+USprqd+YucAbFLVStps0hvPghMM
Dpqd4hm9T46EJGKdwhFBr/ekFqCyoqZwWK4XwiuYPhxY/1urxOa+2P5sgMnQcH4L
2knDKvpngrZoETISnTPsjMB67i3Li5gdv/y9MMnz5PftoeOUFy65hKHxoJ4sLWAD
7Jd3kI1IdKT/0oMbrkBg4TL8GFBQc+U2HetBc735I60aVLUTVYAtd0Qc1Lkbf3Yi
zXHZ2tEwuuyn9z5bo3x3wjGMs6se/ky0TZWHRHRPS15PofJNozPG00EQfwIdLljM
hK8kyOBdusMWJN522C/47iv7Gt0vbGgwMq/xBxZLWI6Vz1joypu1dceDX3pzu3/Q
V5ttBpcXsCPVF8tYfIdV54tZ1sRw146BjDpPguL17k/uPCpKnJDHuNEGkCgt6e/t
b2AU9tF/etMH/BCvlhkutXqKT9P1cyjWHjdX85t1vE7zZ5Htl3hd6jB58OT9puNe
111Jx5th/M+SnlQWwXUUiXcsewKaAz7lb3ykBpgJLi+nvl9d7/pw8n/bMmn+p2mV
kWKAcbBlZgZImqUHNRl7pg+0gahbbO6Oey/kuiYDsr9+v0roQRwjSMzHckHFTIWl
QiFNN5j4hdDhYcPWda0ikN9esMOuF89DMP2nFCjh5DtQyFvEJnHsj/qK8U31RPZG
p/JyPM9NTw2YcvBmS3oNguCKA9PRyxS5Ec5HVdho9bZ2nh5lXmI27+ZPbQOsrF+v
5/Jo57/7d1lTAtB3ezjQ6Gvc76CWV9NcpeeQT2skzohKqDjtc158c9owOedEnXqe
8q5dIGaMMRsnqmmw0GaaJ9HpAcNoXrGE0l0HARcw5yitK9VDI2Y+WLK4SM1Sd6S8
ZUx+EgAlh5z6OUhyjmL9k7tsj2n2rv9ynydLCOZxOwxNUWOZl0AFv+MHnFMUE1z7
EZsfXRlxmyc2Q9ZLsG8zUxd0o4uWtBjrdn86GvQwZeCpHH71Y1KckD+AL75EPNCT
2ZOz4K8MVd7McxmE/Qg/EhKADsNJU9AmbJrBShzRlw7TY7rmnLMoxezR5/8EZ+/M
CYaLXY//dWqsXLsqlYlSCC4L5Cbiu8IYihNeG95RaVjVH1KnTOx8tr9tG373rz3T
jwt/4tXmilgDXoEdUW5BjW4asryClvFF4AtYivA2EvLWTGusqghm76lOLcmQywf1
fWssk6OY8nyRe+ouScK3ToGy619r3m44vOZK09tnfEo/DYSkjwPhz2/t0kCTMatL
0aNSRhO2Y/tnSfGY8djavwtxJz9kBNtl3oh+f3/8t7KU4MhXQsXMBNbVI87sFZmJ
m/pUib1rBRclDNBdMtVicxUCNjdE3pu5IiLowmgom2Nuj3Tpni/e7aEIVl5fcBC2
PvRFiocUGiVmIHdV3EvA7IbYfhCgaHgJfWeBuR0ztctfz4gfnFrB/UhSPD+C/ngl
Rm+j+FYzZkulfdok6g83+rCq7DWDeo1xZkS5w32APqiKqDijQQFOrhfKA/1qR6SZ
a49FR0TNK4vehv9nxYZLd8P2af28IiZsVDDukFh1DyI9HobYXz+tI0uKM+itHFrm
opX5pdi76DGqvtvDgS7ayIdIZ1Bw9r0jqiNy1Z9ShcP4c+iKyj6Hl4bnE8NHQ8uU
DCMrJDpKQisCwXh9fz8lvxOAW6+EC6yGoLU7+wUclIxL10ozVyiXXJEX3ToZd4WA
Nz0vIO4HHxYinKS9XCDdX0MXqGALr0vFTdCZWWLSo2m21is6gA3AvmGliY7PGdIx
/7z39P2sEtOrPLWYwtnx9v6ycAibDMhSF0OHOGJdA/+SbufAz9PghU1Tq/ErD2fs
avJyNjgRNNcvQ6b/mTn6SPuXuJNQlx+FilGh2gPzVmG4wzUlE0aM2POXPFXbrTIF
MA4fDvvyzPj2jGah1nhPaI19KgtjRBAYAKR+aZHv3QHjkdebSby9/C3X0cJd/41E
z2roXR818MYEicvfH9sosySjOB3KH23c9fQ01zNBCfHrm0YpaWBif+vgdEz+0zZA
7VLe52lR4WOc5fXCqLIzWYZZ9w/cKK9LsWRHPemVs6jx+5KQkKZRXEbEae6ckWUR
szxQpI1wk9Aki4a1ttoqAO9QwtX8AVXL6HERqCMAKFUOhnkmquyrcBn1HBQHERwn
EKy2HyxS9HTDXRRw/0bvDH+oEivEm/4t6ur4l33zB7N6VfA9uPwAC5vYiDIkZ0pX
k9fnMqI2TYg6Jo7x+qSJ/Qks0SmZGS+VzFDjlNU67DgkG2mHMFd13qYAV1fI+pQk
hYJ4zJRQOPu50nFKRt59dWTstJdvwNkcm7BcEVN/qSMJ8Ifgo/KeqbT1dfpFuipW
tiOE3MpUw6lNmxr0ZjudAHurrlL9BSJyuBwKKkbv967SMEoXv7XGPz3IwqOyDn6A
n9u3BHVaKRmsv+sGGQgs+8RPyKp/nR5MvsFZ7eZugz8JIEceHGAhFf6ABMn/y9LF
1fNcQPB/5mvHm5KlPBlkF4oO6GJ2iRtbg92hRd7OVKgolgI4UfEmxUTMbKga8Vub
r07vEbl4KWhGsLzpC1XKTdzf5dPVmzJWk2ztgaRwaVX2F76nti0+YMEfglQaue+n
ZcfuLQZP+4jXwjg6G/+uG7FvUqsbaYS6wE+3x+eip3iSHmU/xbGNNMbcTEyBdGVl
adqL4i6uVnojqnnOAjswf60y0FpS+qhcUZnyXwXlB2hED++DhkkPJdRKImbOichF
XtLxZohFQz/L07RAYroa4dWvOn1E7K0pxt+swwhhHvD/HYvYTaN6dLP7CzftF3d8
N8XoX6XrKKV7RIEh9h9o2uvBNQWEcgg6CiK9EnBwukhC0JEUyGJz8CUwXRik5yYN
jHfpnGqcOpQva92LE0lZ5Sh7Ic+ucxAV00IEFXHY2Fs0TXIPrdkg+Q5oRVDbHHnL
Gc5JB89TMNjQyiFPJ1Y/yUXTwrLn9nblj7/F4qcFqVmnlx1Lm2miftO856tEd9f3
2h12SioG4qSV7hyYoTthxXtpCkuSKXTEXEawtI3pCO7Xk+208M25/9Au7TpBlyq2
DlO9hsWU4Mlr2gv12m2VNB83aCXlY/B1IRDVr+VxUMIM5Npq/8JInjDxzT+NYFxY
hqq1D3drENSpIUt9maTUeI0cJkE/8ANOMj7m1BaJ4cDna51MC5HZIvN49xNoJm11
cajeZ8H8JLBrgRC68uIChCO10HuZ1nPNQIuLV3he16hYHdOCnli4m5MDozknGg7D
5k81pK7rFq8/MT/Tch0giFsANY8BRGKL9ucA0+YBRNurOFAmsjhlcO0xmaLMs19B
LGuuytn0iRSXKdMxru8FIKO1VtkHH6z9ln5Y14/6nP65vpdSHlM/IspwZHX76cB1
UGIMLS21gUq/3XJaZFLZGNSheHhxnSG/bJs8dQic09XRSWpq93oeXYdjkB4fsMX4
ICbSbpjXjHuoMZb+RVrRwFbig41sFf8lxO7Mq8/88ED2ePPoBsc8fkT6kKZF/fOb
2dOM8EXgZx81luqDRbKvdwNjbLIrvTdmH53Bj6gIURs/CEmSeZPSAVQCiYkCCd9J
mGssAS8COPjM39HMJwVRz8KrOS4n/YPc+oiEB75WdQfdhkmlHJFRBTWU7gAPvbPX
R1wQJqwtiQl3okZedk4yRJltc24NxhrYKPHLUPItYOM+tm6WIFrPOVeoFFKPRjHI
e3WL+WREqlSvsd3IPEwseS76VGNiOOa5O54EWE2/viyqdM9F2zOIwqTjcWKe08uI
o2hJVtpNK8ycZI1dE5Yg84yvayBQ3KnMVJ6VSDskWK/c6bWOAIQ0Qb6VLjEp3fEo
qr7b6MOP4imA4Mmy1sPCsVLBZarKeW8WXqftD1opCabH5hq55ZRgcKyhz1TTE3b6
KghGZMxnDWCqFmV8VQpMXIU+H7KxJGtrbsX+mjKM3Bp7UV6w4be9bd7Z25of8l/p
NuGz6SdhmzOjl1EDyrPChZ83ysCEhBcjhw4WolG5hoeaauc7NoAgc/qodCBPhQ0u
M79khKU6sLr6dombjJveS8RxQAKrLYMUANTi5R/NWmB2zFqbLtJTeqLFK6YQAnBq
W+QpwSjKZE8ufuru3gT8RBFYYIJR2ttqd9oF+Fuo4YMkp1wUsmATuSUT3IytjFqQ
7Nzj4/3Y0TNH8C6cwjepm70p2xMBeS00gRnvJ2RuEeb+qXLRUhYlJt6czX+r/oi/
7/hYWlKQVyE3UPl3VJmDr5/Cu29WXpIeZBbnZu6gZFH3xD0Z1wTggr/kfZLTACDY
takFHARzpRw9xXJcldrn/mgwSJPsfpGyYflQ+lQJBqCqG+L7I5H/7xn4T9h0F9p0
64V/1OG3lRyb9ZD0WIk6Jpf/FoyjEuzTs7uUL9ICjKKAY6X5GXWERBbOAYw3nF5O
TUpukkymqR7QkvOVBFlpYml9Cf+W604RySg2itj2TbPrzAqEnI5vH+AMN1WUbvIm
shYRoOMcQKqpKAfkX4IMiSaKNCtBgGTs+393qtklWoeLClaolYE7VNTYQ1+TCSM3
Uh6/i9olNaDZ2c1mbKyHsemffyG50vPt6XO2JdeF0NpQAAzvBDoYuKkDMYMxGbpn
n/65AaGXQTdVxWVKxwiLjQ1DibNkIAopju8SOaARbAPyE3ovOPDRP0BMoAzECmPT
aNzbUAtBTnS2sPzlyUq2MmtZcmV55LVY6UXgWhJ8x3SdQmgW3be38xHl2CyOoHko
V1pZNanjvctXprrodenYHDsAvrCXm+ueSA6RG+wZMHItzJhlRNHNp5CivRoIRUKy
07vd9UDKPkKiVbV8M9Ek2iOOpEj1QxbkcNy2hLPkCihr2bH1G2Esk8s5sl1GPuwK
dpnExQ5WfASqmWnTDjU3hzIxtL9V4aONfrA6ZTdLpj/88nOXif0ufHvxwi4z3dX2
jbetJX7BMyCs7fC1b9qZptdotMhz9ERsejd65hYDQYWEOrv8xRBHYQ2I4JFi1HKF
m95FO2vDTrCMBMvccWd9NqF4ilFps44ATLfBPM5t9bNQFDpV3GoDZvmMmhB2QeWr
yqQazf6pqc/d9Ofps0Yy9VTvxQR8pG9R6qOzlmtLKzkhCVsqtWm0j/IJZASCzLIy
f/iUVqrcGXz/R5kjx+bffk3JZx1wIq79eDwljVcLOeIcohL2+jXaqAUUQWmqAmzM
fmjpaL5D388frMJlzEYyu0Upi5dDbHn84t17lefwekbtvLDSn8zvQ1e+4MVz1qz4
hTNJNrvsd8mqvdAnNTLvB5jQWDHrTWW+/TtcfBWpMPALxykjPUmyP7omDuzxauxV
mcnm6FE8AfiPsGCKwzdllAntLGQGmIIYxUu4V745GbeBRLAecAdllreVgyWkRYLe
azkvbtooRAaKC26fkGC5P1mnXu3Y/L5wO/jNeNDNvKTOARH5bqtZs7aApNUYHz6k
CsvqXCWfq/SEo938o+OsMFBYlO0xJnlKbztxZEiULIBLTThbWZE3AvRQqLagUFmD
6OKWb07jfVFXB1CSDPHwWk59TfzN5hDLvgwf8p2QB6V1dmM+HvdCOjiUe/N+ikKs
hE8nS1yMlplIVO168OAz2N4QjyPVsEeqrQcehjLZcUHmZQeozJ5etjo8c1HL4RMn
lWYL/tTYyzw6eBjuNKMF2aJ0SzHzhpoLNRbPmmT25iw9Vvj9oLi0JJyF0r1PBUs1
C2zXgvqvzw2akBny3+zpzrp6QQqm63arwjEa86UK4GLfumbxHRIoeAIfhdXWIzAE
ZBjFoVN3qKfUwx0zjp61SR7UMQENm0yrWXlKIIdbz0VD0fEYQwMdqNEMhgv7Emvp
33Mq6izP12jqhd0xcSmLY/K5uwgFNoR2NYbLqstpRPwgTkoCYlRYAsIDW06uO5cR
e4ZSbpT0oXln7r80oPgAE4zDs96cCxk84L0annZU9ZxBp7xqRKrT2XMUhzuawEFP
/wkPJ/TODxpaM3XgO0lv6K31glxWwN2QqCU+50tG9S2jlCaPXvl7uO9Q8ZB0qZqD
LMzii02gUgYqOmuqi40FSbWlDT6TPLn25dsW7bJgmkeTmxKPvuHvLkJ+7Wkrfjk3
tH7yN+swQqAKI21ucHpB3+v5H6uRVcgVWzJf8kkZ9w4PsRNq4K+hzOi/ojcSUHvf
zjMT9DjlRA34viAlEZXiZX5Pjj3yTQDN8LeCIOQmmYiSNhGHVhZA0GSO0wW/vkHI
yh8RJvKIbgGPd+7KOKV5mgR2kbc0Pp7BQjFwmaJMCmxS45VNIgVjR1eIKtXfOSC5
cVNdx1YNyM5nIa5yKgnn7uDB3U9mdvFH2sTqNXswQ7Yc1NY1rj8LbiTDak7BWDjp
HTBLRMiXhk4GX8XWTXeHAB/fukT+yHTZZgICbafGg+bJKtJQPUgLv4VTUoLtpVSF
ZQ46/esDg1mVKPQCH9BUfm61T+56EgkLttCjciCF8fRNVeW5t9KNqeevbyIEuxC1
05CBS3pr9FIb/AMVjPDwZPszcWwDjikJ9cRFzJguxoHfEQWZihLhZ2RIRAEUnCL/
FkU7S1wNwficQIRiwmADhQDEu/WLD/VdVaNx+AQnkNI5t+COK+faPLUnj94eWdM0
X9cX24eHq7YGp1Gd0lB+h7F7g02J6R8rjJ7MPK6OfmTFbnjnlyQgASM/2n2An7bi
zY8B6PyVLuG+o/xRSAFi/Vg9b3BLQMcDQijz7CrSx8du5kzbwJ1J6ktBvv8akgh1
MDg+weu77xVKmPtkPFXjZHCx3sz9W1X6bN+QJnIrJThTEk3rFon+ztTwB5LMb66V
3y0JUYD4Y+F3rTTNgxb1KBGboEa+8OIiL/5Np6jZprUpk514gD2qpeRluKjkWJM4
IHl7IGmUpEgAyfbptfiE9bGlxaBwjhpde9zNhx07DLyq56jq4s1WjprqQb5yNMuf
8DeC21y6FcDV0LVl0u2g609jouQsgQeV6Rp533sh6KFMky+WjSzqQF88r8dFK1nL
nxnKyRT/oHxkbNPQ2s2OPjHT3NchmGb1n99OpJiUt1oLiOENye/16S8Y3Nfkv/fs
hJo1Qy7UrEiRaCU+6LZDInFhTy73plj0czany0uNMXj76dBMWx62SgElgUFncprF
dQL+dHA5mpkHc0UCy+4jpmZ/EGypRjptaSbXFwgc5Rm+/HeavQZ2ruYTWrFe5/JT
cX4DAgVyuvK6NlLtYpd2UoQj6CBVdoI8fksJa0tcFL+jC0Q8EbiXdP/klXncJXq2
0Vrqdu4hiAa5qnu4yevvmCBP3tet7v3qdahm+kzeb0eHnc0Weeqpw9JXKxUunIB9
1APt62mAVNd55Av5OP8dOVVcCGbzu9CVx2tIcQpHT39aw/AIirwqJjNi7TfjeOFq
zeUJAKKZHPxuIjx6bQeNMmxDMDExVEi8c+rcE7BC4wijJfncLlhI7H4s3ATLsh49
um7BSNVDqsUSBXjS0bnpWxJrC+gHfDptPJiw1rEEvjcDNmYBiPneENbTx03NE7yp
oQpXxcHQ6dkzrpIZFrnNmhypqvLhOs90EOWFxicjjHPhP/0U7RqDCRZUYM7RqbNg
GoFHO54tXjRu2w7vX9YsWx5cy83T6WE4gOj4GrPv6HefYeDAk+QETKAivzoeMWW2
4sbtsJLN/nNAu0sp8p5n8tj5Eba+q2O2yqx0UrVps9Z06MnInjgjwIEzeRv5ViFX
UKn4CBqO/3jFFGgY/ML7lEuEBHOQHGvvY3/QQsxhxZv8m/BQTAMIEn4F6lfVVKXD
0x/0v9Zh/JkJYqWbz2DZyocCMCNZMvFe8grG1poE5h+2F2RWUlJHjAykj52rIKhh
G3RAtgF3XGXs8PKAF2aCZEsXoq/mwgeUxlI1qoGnauq1EXh4F15gM948VIuTcK/m
TcMs1dZIsgb9soNE6IjQK5LSvyQ3O+/vAoGczJaj/uqsIubDHDZ6NKM2FN5aEnqv
YjXGKdb8YblCb3mnWF48pYSYrPHR4pCRKJz/Jbdfl1AUWTbwQfGXcMMj39ohf/W5
p8VHZSLLhgGFjEt96ZLZrm/aI0EzYxWupmXpakZ5WhI18Gn4f76u4SaBdZ/+EyoX
T2COZHAhTkynZzoHr7LMKXYAW6RlstBL8GK/3SYpCs1kKihJqfdQmSldvrlMOLDK
8AmouUfkyEqmN+dk94TQXpb68CVXWEDnHhHYdAPjqs3Avd6WjH/vMuQtJJn6NZEW
xNmVM54OH03BTZBY0Iy42m542uzw6YWhpoRSzgiy19/c0ADzLhsjYcSGWNdvSTeJ
iLDSE6dqQbm+Jb7DIl1cZdsvuZi3xKuNZRVvSwTgwjEAojKUd9Eg88k6OzsDmgiL
mrHaGKENd0zrUciQ+WLa16REjRRLxa0+mkB/akKY7+WiJ2GYyN88nQrKvWPLrwxx
xFMYtnKzS0tw4x/B4RZk4rxE7KOEPd8J+jgyQddfwqw9O2b+7fy2TibpCWVwCq1Y
VGnJBWmh7rBBYQW3r6x5a8+QDxJI2jRKicMrGGYtLcy65cyI8TFwvByfBdzEztnU
QYy/nJQI+z1tl0EDWq0Gizt2qjx0IKSHyyfEMWcDovwTdnZNJgHBo+zsOGL0pmbd
KeuH7AfosJa4l/V7Bd675YE82P/nuyj4Tsxh6puTydapggDZUJRS8KftfBAxcBcD
pdS7/5T75M2alusng0ReVykhBZcODfUlAM7Wjb7Dk70kuE9NHVMK2hxCNSWngcgN
A4RBD2qdAmy8GMciBAVGBQ7Lq7HkfE0PB07slPvs80V3DS6PJWg1huxIspeEUYyD
IXDOxB1G0Y7RBhQ1SSJud8OWycTd64qXGciowXitp9Kd5fCRvMIRYhCMQa3HWiLs
p0ixKI9/j4I4I/TjOrFwr4fAMldEgZ9rLW2h5EnhcAi28wErU1PJleqCrBJJkbWM
GsjwnBeuWrNQjNHga1k3VOWjLDz3Xminjrs5Z41IjiPmx6xnRHD/sdQi8ObKnahw
1DQwjAG3TKlaf8ggIF9qCaQZctb6xybMNBAQzeuqJvERZXmDoYLS9PklkteLLLnX
amfZdRJeMD5kv5G2Hiktuas6ARrPH0yEeXRRuvRryQDNTE4Tf6aALA2pmP0mUSzr
NqLqPV8+A9Lw3qS88Z3HJG76HlgS8aqD+j+v8uhKTYp3xCCm1zV1eNh/n96hAoVw
Y1Q1ckYjVo7rwxqm3RsP1gPy5hM5tNPZc4o8qXkNRf6BXiNMlj2wU8XA9SfaM9IG
95xAeT7x7Za73gmzQJMHIn56uGbHzEiWfNHEJn0vZM6sczp7K9E8A8VE8dG0vqKV
tv4riTR0cQVJ7/yNJoQnlFujZyaDYPjcSJ7MzCjEvaEdaeqTpFO2A/nRXzrLPWzt
WnlvTi66ilpMoocYg9zdRipe+efiJMwPCTIFWjRbUO2AUIHE7sA9G0+toXih0pjR
5neXLzgdTQWZIGTfFoaxsPT40bFVID3Arg9gFwyJRjvasnbH0RCCiTN4i5fJPYzi
D7sOG0nhBCgMsbfVESBeIB7gnokxXAo3pX6bvRGAL4n4kwCia3LX6GzN72/p6TnX
MrDFEOD0Qx83CpOaGYaiAYqBLcOhkVNDCtMnsv5Fa/tT8fVWc56YVPdsFVu2h2S2
zU4mbzr1vZhgkyBPy0eB+dCR8igYZrDx0v8M9iOB3fQtp/EgF3UsB9sLbQQXA5Pw
qDxqVTfB8MH2YtL9Bh7TEEhWl9rcOfwI9bDN/dsEqGtLbqGt+P0ZIomCrjOEIorn
sa/5lnG9dnwCsCkfgz3ghiRram9vZQXYmXmgdc0PUYlqgpPNklKzF7Upx0POdcM3
mf5CukEBuq4H5obC4nzCK9le1hatIBJaKtcEvmNnOYb5ZDriQjOLIxy6aiKrUssM
obbM1mm5dtkKVxDmgvtpXoO72CBYUdjXjcSWsBjO8lwphevMn9ww2KVTrL4JyTKg
hTk+P4GdGOXKq4HQNtaLZFgALXEQjKF1oqhvBziCuyi1XFdfFKdSlqstwE+kKbRZ
nIOZPHhPjBBuMYw1Ro3uGj286yoXNmBgjochRGboDvv3XCueI314p5ecCbkvp8sk
WGGeamgVRInsX9kxQMQo6zYFSJfY/hGtDDoDG5DR/UYZtD6pjxp27JgIzEq/ymJC
cxQktCzdNbHxOmKlmp6IN0UTlI6w0H8AUveMxX80it1G14Y7W/L8hccSem/nXvQZ
ea5I4l3Zo7+htPWcTJikvDqin9nLgVROIgSOIMJB6lsb/osktcn520k1rHo72Oov
24n3eRl/YVNizwqJK2azBJe/FqcMik+ge75C0DCCQXHvyqvi5j+HYvHVb9Zjq30d
nzW40hH4gaTcdVTPjcpY634DXVYr4agXlUFk52UZRKGcqlKoHn3hke0fa2XqU1xR
7nVL6uFG4hK7DKjT1Og3MvAjZ520EqUj5Gu/Vg14AFP3XHusJ0hdQOstmIpBM1az
JbFRM2HIy8SyoBXi1RUtjEiBoT51q09lOIkhTlqkEvV7cbWK2eqaTWS4gqnEI6w/
Az1101Aae/AUeU8HWac9Yluv9fHfEDy+oG8BQVMNmnQfTrjI6UAqGjeZPoZKAjn9
76tE2B+LeEwV1ho0Q6JcC6DGzxvCRQQUlbT9S4/uKN1TcTm+hEW/prYMkVoHi1/T
j16CH/zyeWeSm4zuMDjNr7ThcrmBYt1bOAFrtvXi+X/eDfCNT7zecs0NW1p8VxMq
9ONXOIbQus+I2eolCtFn6aT+DN07eRJQNfEtFoIFPL1K+vOHV+IHfOkazoJj1l4d
uY2clhMGrORfNEVKDjx8Ry8t0a8aoh1pWoC0i7ycjgPvDFI7nf+mv7bf/yFZBSqo
5aguL3rAx0bPzqsSkExKlr4rRnJltYZ49f/kGcyGl1TU6cmvgcMRFUlQX9aPENYh
1XtyXG+noHA49ANrsHrU/gThU9bRrFGEO+8o9fuPyhtvkC/ozpYpIwEPvD3VuHd9
PgBdLRUyPqFCZwJRUy1gEetsOc4Qbp5lE2Sc8NHOReR7M8sWuGl2aTSnWQYdrV2P
r0VCrW2icXj1iGXRi4zkSZBpCTBtW9E85EOIHB5yNs8S509o5TovAy0L41ueUMAk
/Q3haZV6kEFK1T6jqFZ9YTeGtjOip+4Ph9DxIJMwOBkexs6iXZ68jerbeE6rRlhL
IvN1O1wHq6EfMmA7rx0EdP6TSLBHI9ZQtG75G43h1S/cc/EAvBZzNhXRPfVFeT+p
xz5KxFtUC/PHUZuVOcYqEcSVmyRfLYsAPYq+kixgmvBGOKKc2n3iFRJV+kDw/xmH
cx9Sgs41jvcS7KLb47Aix2SiwShC68fmQkAZiGFDuLOTWWJdSWB9ygMKm1tPLuB1
8bjKqz5LtlIPGhuFbLDhzhbt0vYjVKsb/XAlpKruBasONKFLBx0b8rLu9xfUIDLt
/j/puCSTZLSM8tOIg98cCMP/I8Vmbu6dfJH18JzcO7zbIgEa8oQGSrNQl094jq7u
XMLfikCpKmfH5X/VnsiRLZnPGKwY3RMpvPKXmF90fhqqSg3YfdN7mRQm5aVEfKy9
pGBd9aY1Mgej0t6lv8UcXrD96CbVShsiqXuatJkNDOfsaW/gtqqwQwBTIYV/GWHz
Be7y1O024GYkKAaKcBALlpeJwemdOle5x8hXY/EPI4nGqtTjHaZIS5YJs3rxHBap
XLKIiVwR8o5GMv8KevXJTQZ8qQ6vpcE+VCH4fkKJSPeyZjtDbrfkMl+5dFepjV8y
JuNMIm4fW1CSG4KD/TBwHNAzKdlx2z9wvpiLSBwwFEoLJERpF7N1NpNDUf0SWDVa
0e4klhGzks/98IV0TOaG26a1nlIFwHkzr64tKovYqdmv8oAtI78NYJvcRy1Hix7c
upiuyITPjcaG3OovrPzknLKQ/GAAaGKIaFESPYASbb7EPWzeH72Jw6O5wy5OGwAk
6KBYB9M7UIAqXfZNNTxug48q0RimZuncSd45gcmo9+Cl1RMxoYEU2QiKbiEFKGET
zH89bsRo9piPkdMhmlDdnPjo/262q3pEWm3LgkmYs9FbkMmqLO0m1nLLkylERLr6
tEcvrFFSERTqKq63Ts9KRLCgeiWly1skRjLNvd5KbKEKZwbdN8D80vaRa3Y8iE+f
Xtr7ZHinZxTAaGtpH9GdH38IwD0b5Pk9u7Ktf0h4zprH2L3qdUfJaJs+tu9nAdcH
I3Xe49fZL6q1kK0CR49ULNsrkR74CzWd8SIclLPI8+/sJ1+M8i6knYnjV8sIrsp3
BEFeYPOgPRZO7saNrV4zlkiv3f4qzPT3+C5Og+x+jf7gORqEmgBXbjf0Y6e6V7De
C2IMormW5Ds/42vpC0x5gqNxkvaeDNlyhIEZdSm7wS1KQ9wgFu3VVSe2heyZ1/J+
Mpx6L1PLjjkZyjCJKCx8Ig75yC57CeD0L2gcsxPZUklqKxAsq0safgGlEBRiLjV0
MygyFJwWQydnjXBpBRQarEmbltTw6XcqmjJTCaEBflWfhVH9huRkyo30jxFMDp8g
1F7vJU5F1BPMp5LEpjXaE9zcTShFAAFcd1xXQM7K6I9+A7VzDMJCUQvwJsNzLUMd
CsD8TvrFKLNXxj/9tQi705qP+1x9WoU//TD1BhAZ2NfPoAk3gWV7Wo5POBKCgyJH
WFK0uT1khvdCd5mP4+srfqZke8d8hiFYZ7m84sZu576+6MwXmRm4pbVlkFIreYAS
GSaHZcjK0mB9FNvn6wE2tXBKO+lvV5Ieq0m0VyjHSrEL1YG9iS5XNmU1aT2r1syS
b3h8/wPHWji9urkWodD7M5TLD6143nK8B+yc93QYNejDa2V9XmokFR77d/2rBThm
W/UN/B/tPN1JPFkv40rD8i2vHTtsMuq3WWVXp/j0y1k7btsSx0M/kRKkAQIir1a6
2jlzYg+HPvLod7hYG1VqSn38ZyLbZy8Sszts/NY1K67Fj9VixtEISD0wrhE2ljcR
RqyCwMap26TDzrGaK7LE8YaDZ009q4hV5SbbFO44W1OXfAVdn8FcuxnWngJ+KQRG
Yiz6b58E/LdjutFWe9NIHcEiphtFMo47lPSZnHTHMD9TExtOHlq/2TZx2/AsB4a3
6xmNZsI9t9afu7QcoMrrcNQavXhaRcaGiSVua9P4Ux88VTqC/pCWsDwx4E5ktOsR
Uqe5dneM//KfJkMpnIfDJhszGpdB9dFHS3r+bef/STwCK4CYKd0EgFsLvF1vPbP1
uxl799AtecwG1a13jjge+jWOweGfE1n8yo3j+uzAFc8LCjKSqppNTeECPY/2woaf
jYZMYsn7SpTG2K1Nts76/FU+TFrvutigtsFSXmHvj3H/19S1yWIqyUHXCDUULGSH
FFWXOwHpIfzZnZPsyQbtSVagMv0uupIHrdkKgt4z0en3x6J0T2DmaL1eBNJhjmY4
cIJrnMtqSrtPAoKaMlYo+d4Nz+zJITVpVlA+fqh6kCe9JhRAN8bJ4FKGf+1skHcN
sqkam+co8ya1bQbDlUZwJZlbVRDjeJAHMOT6mMpP3zFCtyFaUtubFkDXppKUYIRu
DzqXgXntOqrnds4JYWpdyDsGBnV0n22v5H+DKgJ1qDYj2KAekea7Ms9iHY3+5IGt
iXpDm0mw0pzC9U20ifMyEz5WBsmlTrGUIFxziJ75Lh7Hru3JbqrxhpPALDzUmEmy
bOHv2VQs90WSnfs92BffvZe2IettiqDglge8t08cDOyXnc8MY3E0ZFQvpTVLjcLF
pvUv0BL16GTmM3VwZXsNB/sdh7xtgGhuOoYSB8FwlkwjSioRQ3BfUnvIhVJikyRM
pCYf1NWOa+JSMAHYoXdmH2Iz7FFUQeoRe94I8+ipR3h0sMcT4ojgKkIjVko4DWzC
I1tzLawvz917bn5SyyizMjTEcMmfQzRyQ7HyZns+rx+9TRheJLsZExUeEuPE0+09
o6a3TaeYdg+hKVQlICZe0b+w/bGl0HQt1Aec9dGJjdxwQoWPLt9vrflqYq5rGMQH
EiBceBAOKdjPmNd/17Y0UfiF/eQ8kdqjg+tOYU4WNfdj26NPkaLOJ5qukfn0BBYq
/lFbN3yC6V+7VF6y8i2TcS4PsbJSESheFItk6NVKPswCbgOEP4QsoJMR8Jf403p5
hTp+SSoArDuaJnkCLd/F9tQGrHncKDWgWMsZ4F7InoPou42WvnJLWRv+Nlp5Vny6
1vFCVEGhm/AdOtoguCkJkda1bwkEaOkMwNcTjrf/i7RIkY6LIWzU0jWcvEjd3KWe
9zG+qZHaF0lC4tcU7mNF6Z9fsSeKw7nkmSj/P6pEvyuLRBDZsLUwXs3VPYKD+RdK
cS9nQFpe4W6Z8QjIHlWLrSHtzfZlHCDfZ6VblWyRXJafowk/pLfStjJ/972CnFce
h47c6xT3X/3JfTZRZRWL+SXBpqvfii1RT4BOdKrayE3eqE/bqK0pSF5pB+CJWAGW
MtV8boZ2IKj/qei6SoY1w1VBYs3KE2nGtRmBHkQ2sTnsVArpeQCcjoFhOIWuSRcT
nO4kd1KTgCjoK/KK3xPIV8xY1Aej4OZGJL++Nv4goNt4DePCpav3rK7ukDZKBW+m
0p47IUa3+wKg4vuu/clRlZUVerKfefujNqVUGUYGZksG+Dt4694dEx5uD21M3aDu
CYSYMMkYaY7cl8rmMBbbjqFMQYF9RPQFtvLY8EDHIzi2jtEamM6XkVm78Jvz4dBR
3FXwFh7PjPjxMNJiLl00Jp6IxT4t8/Qqb5KuyxmhFtfBcECSfX+w5Sa6Lhn+9/19
2x+9PX9Lwbv3tf5i3syjDRSOB7yFt2u9UPcusMJcEf2z/DnzxA3oS3ySY0FiGHEK
emsBZN65/PJUkJluy1yqz/vFcUG2L2ROgaUv/qokgy+OSFnjjRhezGKv5bj1rNTa
E1wLUchmVR6u/yRgWEd9STXVSKST3Yxw+/xhNeEeI4HR7rDIfYp48DkPDTY8LqpK
aoOBDnlqafxpFch8tTNtuJb+RhteHWzaFA0xkSrrjFGauL7ahRK7wT/ILqSkmrjs
jldYX+mDQFJpvndn3kDklYlivKEWPTLRUcJio7yzstXYBcItuL4fYQhBrOBWLX8u
n4Fk1F+3ml+T0F5r1so+v/vmKN5RlLMH6z+YT6vFRHZGM9aivj5aaWLlSeWkxyL3
424NzSINWCbKfHaFtPIzF0kqiKrGGUdRrVeAT8XMgRCqzyOCggkTN0r22fWNtQpf
ZdBQDJppj+kwoo6cjFIsjYwmT9bUmj6eD2nrPaI2mu8K8MUA2Ve1uluPrVP8GCf3
0+vO3xIOdK4fbV/8kCm17fwxyc/4Ipgs6eccea5rKA0abqQMBHF8qB5vjZG1EDW0
j6aZRWdoXMxdt+XiYgMr3Jzg1nnY/7rQAlgwPKGGLS0DE+fIRqqlSn9daP3chg+3
JXNVP/DYqU2dxD3jXJ9bkCOyKrKlklg3mIp1R4qWyzC72soov0ZSfsTPCU4TC7yM
O4r68f5/EaDv9iF2w24WsJl+3VdIsLmrt5+3MRi1SRzZnYvjF9JuryfYlIBjSxnw
IewfaLYDOTElaPKeEW2YRY3sAUOAh2Wea2IFjhhcOW21L0nlgg4lPEJejYLLbxBD
hocLeiVU8q1JWbGHXSFpzRS2P3aQiUgh2vrpjZRMe+BEfHztzbvzVYGzunMuG37h
azcr1taLIrkE6upY5CIOSXgxgciQ4/iOHNExf7ZWEAnJp0PLOv9V5AYG5dR6QFn7
FpazExP+zw3toUt79dSyjtg/EehYs3fu/upHLhOSkmGwm0p5K9kjcCWjw075uNHk
P+Lm7cOrfBdM0Z89DXearkEGQrOP53xBtT+jX1t84NOSL/mvYNO3WYt/SL8bC+qL
id3GhQVFjR4vww2uKXDyul4CZiaJ+0QWhaXs0akSyG2CF04Uhv1npTQIxAfOx+IE
828g6b3A/uvaOXi6qQOtfMOTOqd9NVKxsFoaBkYPVaQQm1/684iJDS4r7VZ18DZ2
S0V7e+o19ou3v9GDyPaL8k1M5JRgZg8i2jxfdJL36W4HxDNJz5kkbVhhukvm/QCW
2vVAroQRRf2XpCTaG90lFxGEp2KB2q1EJAsCNJIyqqVTda+f0GYA5EvRB7uJF1CE
IPIHOwmgfGNyCVYAVljRfvcVe8JKpCIZepiCom7shUje/tdbufyQgWKxuge6cP7f
x1ZPtix59RRfiBAgV4t/AbV071DmxS0ygx3LUnD6tX14zuPd/B/w5HWZ9hYB3IHq
zSS4Vn0st9BQ92TPctthaQQJPmtK82Cha3uhnIv14zl/3mNmH+QRkRfZMunbFt38
8LAspk91oHE1MBEqtKtkpmRmcXRd/Epq9jgY/isJu3u1B7kxKkTR4tqUDrdYcRIP
9yF/vs1Uudq7ZBgx645StdPEnVCvaz7RKPz6aAvB7OUBdckAGnFrsQYL+7h4Ufo6
NbejwWiy6rbvrJwxFvqlylozxPtBlDX6KVmo5mnsTWKP6qN2KVVB4zFIH3Fo0nSL
tfl7S0KAnH8gbJcPUTDVMlarfziMu4UH2qELdBOlPdQlI4RsumtKdTFvu6VRy1oq
+Uv4xthjIjshkLk/+IJ3M1xLLjEKAEJtii4xt8dLoHLMqwq1Khas6+AtDdVw4GeJ
Q0paZO+k5F1AYa/yM+ljVyF2ga4gAP5mm1iAV+NvXaUVNYvAHP+1IpN1qNba6Es4
iXCQ5eDuQ32PHXgYIZwuSZk7qCLnhnyFuPKZW12v0lIehdo9MkbtQuaWLr3QCs4a
a4nkg8tFSUy7bQ+Nj/+0n6fWoHykrZi4KfZ7hR+suCN1oh2PMWSvYL+aFkmfmzze
ttIt0UwEnZAjcO1oZoD5LaObvGh8XloY8eAZIClkOpCY28BqRRPwTNvCG1p8Wxa4
C3pqHqifRaJL88EFuqtCWeaiR957rMemDIeFMxXF28LYzxrsaxd7ONzYkvxFu45H
ZtnEnhfc0yXEszkANN3MtDl0ONU8prUqJKt2I+OIJa6PJPgbOqIMlIrrz8vhP6X7
MPP4z1HbXcqXbzP6D77jE0T2dX118+Iy5UYYKxCTRToK8B+48UJP2YF2RXakGPHK
/Bk2y3gswP+WkBUS+ZadG/SIGLXzC8KCNFYcQmAuaMxgQoXmv8cDMfffPDVErM3b
u8AtVySLmG2HIm3sWSilrekLh7ToPfwTICKn3nFrUCeAJDqWYssPl12LsTQJltVN
cCHIZTLDCBvTWe+vnWOfYOzRPRP6x+i3In3cZhRGeh9ssZbISMSN2Hv7Dc0oFeBx
PUcW+vU9KLNnAqfoCFPdfiyW9W2/F+JY/4YcrT7OO0TPIHmriSkYWVuIJsFm3H2j
w6gmMRJ6X7fT/A5hAjgIQb5Sc4jYAzFwNm1GPP4kA0USnMvz3Gqi/OG/A+Ovwreo
lDlH7Arteq6Os5ZiAvWxlgGKyr8WuIXXa1xrv35JWD7Mg0Tbb5a2KxdFmem68kqP
ZYvehnPBKrWAE74cs/ke1ZZb0u864CE8rABtrT58Ehl5z5hj0dF05/fpxQG2BH3l
7klo1ksVpOYyVw3dobJ//LtWU0EtiXuxGjHqMLPYfd57GEYjr+Y/AX2i7um756S3
igOCYb6V1HNUFpJ6u8IMK1HSg8SioPYQqHu4qf8pE+yxGbgk5X3p8PTaM0hFg4RO
CmzXWox6DeP97GXxG+xWOxGGSIH9V5FQb2LtFFPDJtF0roWcIkResO9PxfflEfBk
fjQ56H2/lMqF1S9mSaoajuJQ9B1baTfBGppGoaC/KdQdJ/gToIholZjeJKHb+m8M
IpCKGdu+RZqT2jgoiQbnhkGr6NdP9hLtXpTu/69dnZ5DUSKtN16arr1kOoSx4XeO
H7369JSqPBC8SZlSO9ct046Qsn2brJdplXSem5rtwCX7JcYYM9M/F3bPEjIVONsq
D4nE2OLTrpvM8UCL4yFiJWMMzQC2EgLxW8J2A0J0S93aPSXawTk/8crz/ksOFAp1
gu11vbj1VzS0yAV9HWTg2OA0tyZPNZqd8o6MBGcI5QhdUgPKq2zbrqM1jTL41KuV
pNLk825ArCJ0soL56flWGU7WSj/0S/aPQgStLdH1LPKpog+K8kztZ4RKWSlKGqOR
tHHBUirRyK2QTGs5egTC9iP8JMg9oLLj8S88dmdgKZFI+R9We+8QRrY3Hzt/+1Ag
6Yn7ZDjZCDd76/lg7cl18caDKgCT4xzUrwsMEYWmH/xL/h/EOihq/2EvEoJ2sDXq
tLzcjcfy6gOYTmGOBziQvgoBhBO57YPooOPG1+VIVesr4KjVhMxPSI14H8XL1gT2
6miQsQRCCAEw/eRO3CkIkCDpJoW27dkfZffVY1dEr/cVFImZSvHDxA69dUEjiTb8
LHhcdH7DUBMK7JhE7IQq79qow7ow2z9Ynb/L33xe/FnwMZuFBBYifSdLQV46spi6
lsPi8BUJE4/7oUcaYWSuoIb92JXohYkWbfwqDZlTlCBg1qiwHoDdk214cR3FkoMK
rQUNg9jJ/A6yLlQorYPpmnjYo6xuQ/+TjrqBjrvs6DCMH03812WdzQ69nnygw5qc
JAOjs9tJisSZsdTpRjcC4vAYXBkLiHilfQ4UbZ+LEntlSSlIWIr2foib8TZ3OWJs
xFG/nme6ZquL55QKAGGEeTxb92by4/Z2+qQF2vjczA+QeIzJzOPQ58zlTnv2qtSD
Gpn5N1XtHlXbZ31Vk16GDBfMORomwD+YmiCltrmdDjPDA3Y3xC6Sn0fOK3KWnLPl
/kvaFE6U+q/svoJhcoKWNdbQMQJa3LirBGqWen5BViKrnAhbF+/xmk+PprSiqC7I
NgBvoAHH3clO3SqMfCQi30hAFvAjt2WLnpwVbcH1HNxm6a/OiE9nYwBJYNNAr4hf
TJFnRI0AuISzItD9S96tzZc8MOKPK2f9IomrMBcBd6fKrLx9PeL/PG5Tmo8ils4M
4dL4NNAzVR6d4YRcm9enaxvQEuyT9jOcNc3Tg1ke5RBTBW7fiN19NiMk1nR9MX+X
A0qFt9P58BX3aCnfe7kHNUq58HCPC+cxWOpGsvOFdW+Z89OqjOwdVPIRs32kTV/Y
i4mKK3owTxbgg5tL5r7b+sQGGIbukIaTnw2SMOIH+pr4SoMuxJLBn9OuQAtPqF1/
Ji0bmI1d0aEbbZoK5hGQlX7rpgDzrQJ2OX3ePUja7vQyVf/z3z0Pk1WXPMLfMeCx
yqn4a8pAzaHiZjld8nqrOKSohokYzx9VCnsLSfdjo+kjpWj8D1r86aUO5EurW6Wi
eTUAAD30/gsGxloESVFZmOVyFbN4IoQs3VEy4PBz0bMRX1MmqFerA6thTozFEtey
GuQnQrl72V82ahY4v/nUvt7TQFaBwTs38nM1r5pFOq1fv21BU9+PEVoYaFJd3qpk
yIz26VGzL7/C99PTK9TXRh02GmrdzLy55Ok5/AkskgivYtCyYJ4Tmak8SOFm2qBo
CYlLoefaij/W9G6rwPWbmb139O0sDO5V/0jHcBwayvPfzZGTIqtIbgExwzw73Qsn
bhfmesBe+OtDY8hPF8q2ievZxzG4k2sPXPMO91oWn7tjZ78jEhwhtpcMRPUQO4cn
6GE5+swZUb/q4MkFL5LktZXdHZGsj3Qs5b73yJTEa87E+kXWAjUCfS6HnQZu32DD
PBEW0OZ5/6fJnJ6H0Y/HIxW6Mb/0nI+P0+kZh6y5p7Mmr2yKVGaCeXtib6jnAITs
Yqz6RcenJE9CyjdZMnbjDPFH9evETW6Q+BI6X0LzbUrnWIblNhuFxoufSJ3jDnCP
sGgWdjyyYN4bglfL+3Mq994BPeoGlNUK9Y6TuuUGxYt5D29MYqMbxsfrMZzNPxUH
mn76bHDIy1iq8Eao2r4lWYEWixqwHNI4yiON2esAAuTM219ykxeqz/DY4QPOQF7g
7HPOJwlGG7eTNVvq9TgMg9zDiqS6G0Fw5mJLG3lsw4TR+nFqsAbtqb3PK3/x5Aka
5hZ3b4D9xGvw5PTTXG3xajayssrmjb1QkjbeaKC70llErvV65Fx6VKnlRAAk9pdP
2quQCr45XebwdZ3YGRxzG7XsHxep+i2KAztmBWjLCiqissxji55MB5cdByKigueV
xuu7vdrTbhW16kstbZVJZ1p4/3zKEHOZ8qvFNGIqobVL+xqjTa627cLbtqxIm5Y+
nKU9C5ZfSb6bA5JRG6YiT2v9ItQuQ9CJ93x9jyxip3qoDjS7lEc/FXHV1OCNg6qh
S7rek5ed56YUsioGu27pe2Ug3w+oHwwdVsN/89Hjn4DLfkgw92v5dN9DuFEWoXL2
8xhM9zIXYk+vAD/mjDoHM+RzA2XoMSNsoEdV9tSR2dFl5cHeFAXAoZSANuffbymn
WKoaoZozBYUcc+lcIj3N2EowKHZg4A3GC1MsQpZGEnzZoYtCRAjcnPYtbKrqvcSu
EMHlGP5XaG94NTcT7MVy76fbwwfy0hRpTCnffmyxSOMyRxk/Rfm5aSv1mnnzssFe
FxD8ctLMpY2eri71MMCs30eXE5nub/GTRdOrbhVubQq0XeZ4HzqqGfYemTZJu/xC
jhlLodxkZKHZxHy0lcCsoqpGoZexWC+dIPVf/xTcvQBXrTqiBiXtzN5PgBF5VG8G
J2BgPEOmq/Jgus5rHD5vKo36iJQdXhdhnTGtTRf/HrAotsy9aPPmsrMEIMIxBNzx
JOgTYEqIcdI+Pb9TmmOyoblJtwa+NqCrls1baA09Ez73huwasq3sSpsOr15iSr0n
YnZp+FcK7qj14qTg+roEBnSArccneO5stIjQRHxu007zM4vq4BQcfeIm7P+vU+7i
4HMzhDzoIs2+Y0tT0bJlfEzC7dqUF1oOPD6E5JrzApE7a3m8fo686MrI5x4nBH/W
WAPLF4jFbpjMvVu2gfX57Ax9KWK+2dVCjhM+k/FdnODaABIKzhQHRRAo1QYl0AVz
l7SESWFvHYrINl0q6md037pWAFcqdt7r7AdAUsCuU/ljSuik9tTlxpxpBOg4cX2I
W/ihbly2qfA9nHOLinIAuIAVnIpg45Q27gSl4Bt+vSOnl1vWUQPTB/LAff8psmuJ
rPXjebs169/UqXvZFwGRCmAJ/wITCXa7o9poP5E6TSjP7qJNyan2eRuFmIeudKra
jjFKHjRuGNDTTDkqRSg1awvHOzPNGK1Wjl9kYgZkDeo3upzihkf4cS/sGR0yIxwj
8lwljvam6tJSsPUp21EVu3IKjqPFNXYFGWaaVEM2Z7TmfruMHSi6OoZkfqb3SD2C
j1fXeEoBbfoK0js+hKVummijhyrOofG5ffuH0PLaquY3NvIKdnIwCpkVXI1ToTBZ
hT5rtoEjWNyeu6uVc1cwlscuskwwF8el5EK2TjNeMqwJX4mNnWsLyMy2it81gYRZ
5P0fd2pR9bNHHk2/V5f9AJ1czSaMKdHCY+9zswFDoi5VboFXR6+i92CJYfbWjcpp
yBZspDOxO3bEI+MptrNdqc4y+VTJzq6oOX0xyeGV+8vbPflmt16+qhoiwYZqrLup
040HzFWzpov4Q54Vhxbvdd5+x1DWkI0MlILn5UVYzUFBkPdL3jf27ekdyaeIFwax
RUm/kHIGRazynIlBlAkBdENrcOfIwVex/bbd4fbn+4DFp36EpP1Xk7FmjQWRDIwx
f8nFx7vdOlG5mqOT/j4zCBFla0ViMiNivYSSO3IXaNwFnzG2g+BHyposYdVyVlgW
knNeLZnKreFcbvKSJRZuLDb4tQ/axAJQxCsspFbzcnjLTqo5IqOzQVQ8GVCoTZ1M
TwcXN7xM2QYyUyZpXNbKRBZTaXli6dbN4mYoQoZ0mEQCAIxoVjuz9/ThJbq5/4pC
sDkQvIVyTpHVdNBkagk1MxhIo6/P1Qki5NPc8jqglYOTkJnSvMaTPhMAHypmWGYY
I0fprzeD9XPtgOTqsnTEH10Yq2kxSqYYrHxonXMLSCUVI4xx80BHWVkC35NI+tUz
J2QLzMdvsc7p6pFKQm7Heim+ZUUnPu9Z1tIEgE7FwSCm3o1CcA5vdeOQU3r4i44t
SpaoQu4bo0L2Jl9zQaGkTeHFhx8IWT4xEfeI4/WOWhecFP1whPHmd+GvsT4+8ryk
FAH6I2iSBUf4l7XsOSSQj0XcxbLC+DZsL8rnRdwzgFq6PEOT5xVFjF8Vf78gerb+
4P93/8C+L770RujgShrJewcnQx0p19mn+ycS9milwyTFQQ9jgAhnVHfpomnx6l7q
sM/6cB2px8i3IasbKh+QB3NPipXpZv7vldALeMxnsCXumqmvpBGyccoyvVfNhV3A
0TWzf1s0yq93jJ9MAkAMNYBC07Qr2/9pdm8JFaSp3gE0bs4XrKIUPa4WyIIH4sXr
mDQZWul3Q2h6sC7//ycF9YHnmoy2ZodlbxdiRlhBUmZ7BrXp9V6GQeLpqpFKxedB
F/8QnaD+1kJ0qhPrN3du7H+/0iXJccDAfsW9neMB0ud4X7fhjrD954YWgUeG915z
jPW9CF1LwK/hRCY/JcKnEsrh6clDA5Zx+xA/nvfcrDMn8UktXHzPofl4xej0RsMg
QBi9XP7FQd1cse6+gVly/bXGTJtfoBw3WpKQMchXWkPXx9QIkOuyQkYGvXs2O2PI
zF2kDN7yRAx0SLjJjI80IPaaaS9fnurrpGfuFRXdpfr+SCjpOkrBAMOw2aKHtFvM
Nw8KSGdCDqgIfEde60M6x0DkOMu85NY20Dn4VFWycoyYXlbWYGI0Mf9yAleuEG6O
h3Fftf4xE4Ux6c/ColEq2hr05XzN5AOP7nPYg6QKEIk2/hgxRLHr5ktncXKJpG6z
ucz1WcHN/e79HSLhgV0dJhYyJqaGoKIoYBa2u3MYnuBHOrhlcHf/otoxlRWnXINX
BYf8KORhkcro3YETUT2ctOh4cPMqhON6e9L0PVE1zeWd4LPc4acGjdm1831Yib1B
oWu2ZHaM+0KX8WAQ2XYHIolQHHjL/6xAsLYixzPRXYpQ3adKU6AByNRucsCn2TMV
eyQX/Q94ZdwpL7whKdFgv9Jf3O9OdG8i/elzJkAGe0S9zbDAUip9vi41rcWTj/9a
6ilBJY7Nx43dGye2OnxPYYgMrRaGyKW9LjQ44EhZgoNS9ocEKuYtf+J/CXISHy7o
16n4/l2yIo+FBn2ryyjqC+xhPaxJpd1hMbJiWH7ujJ8JS6EEQZWsAzF/qB+7ERYp
N31Ah+OnkrYmcxEBMsTW5YLqwCnAl9J1+QoxevAcHpPtKSOtBWkd51sQ/YygGGYt
gSztbZHWUMlfucabK/1i7QqES5QxcS5bmJcOH+5PW04BfOEUllaSKqIawa/3sXb1
p1AhYR3SPFVnBObFo2f+WdBsEuiALuGk+NSFA9msG/fqfBMkPdpdHxKXCeuIb2h9
RwcHEF9kJ15blQHJf/7DLle8Jq8E2Nroi2V6oHrstLBtMLHkOYbjlw/6fH4D0V41
kuNV5XBJg3dqIzRe9+BU3ohrW5+YpuG6q0a6sDdKsBVdmffp+kzjzW51kkHF616M
4sg4d93ygWgANapaNRjsGpBjf1MnUgrG6J5gahg+MYQQJ9tmAWIgRUKQClo/dKCr
sA1Jpe47KB3RVTipRRkZeJlx42skBXLgzVEBmmEzQkD/Dux5rxptKU1rY6ou54+S
rbLr6PYpgjtwC/5l6Zmna+MkB03JhsLSaoIDUlQ8KzUw0u/KRShRVfWgb49tHVcO
yquSFiZ/jWjx52fFfjjul/XvxEeSh8ogbI7Nuxt81QRmZO1FBCSd0jEPPZZR8LeE
0CJ4evqdGBBEW4sPfKIPGWfBl6fGZPe34CfWOzu8ZOALsDbvdh9NAQhRJgnlNk0C
gpldQZH50mSO1WHekEdoSNBPUxVzBJ1gKi2GBsxtD9gIn0AK2yWMBAs+NK2lHiDU
M0TP05miEzKPCQ0MKt1h26GMagSD27J4EbP7gxG6VX0pJZHOahZmr94Mi2mlvjhI
xAREmNq/mA7YW1koKfTq65bSKaFPiWsn+2G87Tt+34JbVWwW0B0kN/d1dGBbZId4
0Iq6as6mXuVJK+1FjzaJythBn2BFJtZg2hNQgOH/w3DRCVltjvIiX/lLdfMN63DO
EoxySs8DBqwiuDND3115/VumC7r0b5PoaZKGy7qKudaQ0KU/u03vNlyKWvKM0XgU
bHwKPfMTSdqjMaJrOrqjYA0XhcB/GPcaMKTp3rCnxH8g4uUBvw1tCVEN3cTN+8v3
dncfNt3ggTtCbFLBIlyTNUq+0TwsXMHCVhCX+WxrypogtGAqTvqXJfHNmWIih+rf
13d9xE9ipDH0RJgHlTDEQd5gZZWcFcnO/AKBTCNot43ctiTvH4HxKUV5+wqRNxoX
5zIiAJSfMAg9Hcusn4du1bfETkicQUKFN9CExLUQh3G+OHJJ5yZYdmJBSiP/NI3P
uDRvJRkQZ0jJgY1pcsUmEOuOWQSxdi2DPPZdcKzy6LmVIn44plPrDqpnl9aTUbxY
gY3dU3uUryykiXPQGDS96kuIqD2Z88AJTPDvICeTFT7NcmbutUAp5ok2A7YSL2B0
6vV9OApmamwlIMXBRXjBss77nMiEggXwbzPMbfIYkmUlN3PDX8lqKTzp0M/blwGN
QA0nCY4nMRcvPw3W2HmkhvDOmr87JrlaMXIlBpqT9frX8WIRIRg6mLiuwVZc9ugA
1UWyhe1kcfWpoBVGu6PLExec/ddbB1Jb6yPVZa3bnL2pLx3WwDXj55hxcgNuFVCD
d10vAm7wHQyA7rwpSSXVOXWgfVkMr3EFQ+Z/nacgxetSCu7FlIcMPuX70hUANOW2
HOsJnWVACfOnPxltftqoHKkI7PWby9KssonnU+rl0NJCZTi3ZNQhxDJKSUhszQ0K
Oi40ftvI019ms1eQZLY22FqDBqBxE3gpyPf1jQaGkHJ8r4hPb3MaRfUZ8pL27ICM
8ZPvYC7CjJjlZzKfU6/fSu9P2oGm3RPW9gFXayiMI/E/zSTyGGzMh4PNcrLiJKbT
0OWJaYFJjxvJXUWUR/nxLNt9zY+uClq6V0BhpXUsxQBa2U2wPZyKhEeNozaHq1Cs
7lF41K/P0Ukvggwe8tFGi/R3X+uKULa8bEJCLvhXGzRqp/5d10IvIqNPSp614sMO
xNYeWaMNvqSzublldlQW6d1VpwEloMJ8Io8NjZwilLdkkVVIuGt0cIreOYppo1fH
JtEv23L2LgkrVwfFVqpiyNCRAUBf0+Cddscb9u2v2jHkxtEo/s3mzmjEVfW7NU4m
gvjO2WO00GZHM+ji0NWiZTfmqw1O2N78+g8eFXwydmNIcOVlwZA4F81IExy9oX72
6rhcIUeM0RDDQRcuHyeNkQ6+76557WfScexv+6pilUxkqkaGvROiBl6CoQ1QV28X
LA6Apz1l3jtF0SdZd6AjeeUCuD+zJRjFpm3D8lQ9Eg0JMp3tzM6TbUEB8aNNaMq7
c60+N0bVU71+8dC8unF6uR0vPlDrFj4QCT7gk/ii74XClThZ6j5tFjGbgwrd5ZKu
lCMW6mreau2/ZdLZAsFOKNchkEi8jzkYk5/dK5mvXMZtSnxXHIjo+zm7EwMjDF5J
RPBiLgE5fjQaATgMQlAkGjEYaWi4BrYGqlElIhMF/12PJS0Kt4xSBljW3taaA64i
9js9I36U58f8HeE9DUdVRbzSGO3Vuq9kBFkS85fYpggqlvnffz+7gXK7566k9qzy
/PEQxZlhSaZfoPk4o+WB72pvGa7DzN8mWD3iqDr0v9tNA6zTxCen3gX5aZZgJoRf
jIElpx+qziHr8mrn99GczNI3E6pXOrU011DkvgmC4iFF/Gs6gqzbs+T/EkF7PGfI
QZFEX2nyoB2y+bx8HPzttI86mFjGYTDPRSL5kt669aVJddSk07DGFxwB5ivZ6weu
YMNt/AJfUqdRLW3LjPaX+KP+RBO6ci3vPfOyXc9RoVFv3D0be1FNdMyyXNu8npCS
n07XX1u+QneoePwdDK2QD9+3IyXQr0qSIdkFk7IDOdTc8t2gA4TTN/sDPVxXL71i
90fUZWY/XzUZWJnI8c3Zsd+3QGAgWBPJb3sq/UzLtq4wxSslDUdXRZ6jUQDYrWn+
IpDq7GMLP9BJoDjqb1BPTpxrgZKLd5nSo4HhDs9bbi07spaBOpA3Be+JrZTpM6Pa
L802G9WvftEgxtDWkusO9vgQnbi6W8W8Eg1doASS2ppbelQKGWHLdClBINNd7MC7
sTmhwCmV7Gcgc7hx5FxCQGKWf9KYPGT6iH1R6o7NLZxjC8a4my/liZgTliXJvdS2
w5r0Y0Rhzw5TnUZLEyQ4+lE25ii4m5M1U67SZR8+BCOuDd+4dtzMzNVhp5Fp4Llo
MUFPidjatU1MfvwQqCaRySrQQwx8N9UDOY6COImfLsmtP41jFQQnLYXuan6kU64g
FiYTaO4/lyupq8tqvyjqn/I+mmNXpDhdYmA7UwN+dWsePekSBXhOjqSG4kz+HhAN
dVaPMcfpxBB8Fs5/Z+ie1IzdIbXyPcNz3Jsm+1VzK4FPQUffjSVwnZIfOdcqAMrh
RN5T1HL4SM0gaKcaqnUYaliO4SGyrC04/4sGKRaeVNKVRpmNgs0/hqTXlAztrBIW
NBfxzjUJtx9bXzEKDK48qmBjMf3cAyznQDBUfR06Ge/m06BUu0bgofqD/Ci/+hTw
Zx62LvJQJw40T09DAhzOIPViWW0wZifaSpIinZAZCZT6QM9XCCi/mXO1BIoXIFUG
YWMvZNw+frbgtHJqdNDHRyhIvhDSZSaRAb4AhkpdvfCo1ERkXIUk4XINCxs2oYYj
UTbB0R+k0DHvT60Gq6YbA0fK90bic/yz4Z/BjLxwK63RdEK4kQY3ryH9BxS24hss
xw0OhfwZVa5zCJf+C5j1qKkckDcnZW/DM9sYW4jqJpFcUBYt79RjevtPZT0I7wvO
I0zx9ekS5iOQT+OuoWNMwOwM9CHKb5/ZDtaKwO6Z/KloHWUtyhCtDL4m6i2ckdGs
TxpVesYTiE2+U9jqYqPYipN+8nnMigLJM5JBHp0ioJFGkykr/li9yAzCm0SnCrhh
9imTxkGoQkFvN84HjLtyN6Fix6CQQo2NT/0qURPlru3vZRfYRdX5aZwxlURIWFxt
uXAFN3/sOFVsRT/29Eo/TzdiWVYekS8Dj9rzfagpTyofZGEUsWaYG3vLglqXDBTs
ccjSmMMtGXaUYBVGw+lCKNCcInj8LQeIZjZvSnBFDoROYKMGWEuzv+g0ocD2D2BV
AP4UP7s1kGAX7kVntWwyFeJpjg94Y4TfnHyr3AbD1czCeF+r3RRz5ohpzUCV5LXU
2dMopIl1hicdwuJIyIAb0MormN6UmsMXMcGT6egcpBvO8exyVRhqXWIJqAh3I5YY
hTQsLRaI6ChD7PUOGAA9JnUosvpPCdwxOyGZqs0ohMl8pwVBhV3NcQcqZK1fKCMb
hEuAUGzq0fAYj37HlcePdpo+X0d+U/F1Opn7XVM9n0/OlH227kDM7vbQn94CBB6y
tbOf35S27d4p6qVYxpNwuv4lOtGB/b7SuN6o0MqmXHbjgADnXA+1yXw+cpxO7tGN
/++X/UYAw0Jhfe2EBfohqDjPr9LGvxnxFspNbZ/UVRH08sHnz2hTvU/urLNZ7jvP
Jlw8fyqqOo36uhfuj/t6GrQM+qsiRT9YgSFagGSW7Ywf446XeEGcvbpg3+i1eVOq
BYntW+FS86hGSkvYxrxRXn6vwNOfsgGmTl9zuY8tX65e0tkWSuw4Yp36upSJ8PgK
EMAOhPe737q9HIVpRwiixHIuiR4oUEos7bFcncjfjItIN4z/5L8LXj7l2m2Dlr7w
1vA2AezRsuTiQBg066Z0xbITWP85HAtS7qbxqGPzcooOvSswj1ouhoT/kVuxmxQK
iQFaH7uoB7J2tTLixny6Udxri0/BKQxkxWe2N7yGY0Xvg93OvPnp9yG7AgrNR+vZ
ArKU10wb/IM/M0CZrPRfgTUTubZjtqSStYkmAOUcMoL61h3OkaoaB4GbtxOGctmS
jMXuztjsxCyBaV6ycn0zoWziBDEPx0yBRDfCHRuRGJpaXm93O9TJVAGHPIgUdnm2
eBdPjcxj35vwWwIi6VwZrcli+aRMDm46c2280M23uDf2Tx4/DXThWGbsoCdRNzQx
on0s1foxmFJdXXmIrb8CPofgeXdMXJ2Wa5KRjrTBEocpsMg6QfZTl1IlhE5ksT8j
7RPoWL3QY6g8cZl3le98puRjU4U+XP5ECscwOyKQoJZYRGalSWvfDaA8+VzQ8X0E
x+VI3+IL5Cz4CzmYy3uhP3i9EkIZk8axMLHOlbhbmQa1aKv8oxH3/KeqrMi2zTz9
GHP7cYsQmBL69zVFGkLwndu8nNqRH3hkGkeldjbvu2ba7vF8zGiD/+31174Ee4Em
t7CaJnOZxk80WBgrCvY3gySQTC7Kbzbq3qXsSdN6Dzwp6vrUs72dp9pUQGFCuOSa
ngh8GwtUq+l0SU3wgfqlKGtUqbIZAhrDTz02LcTExhBorOUv2EBo68Tc+YIW+kQv
3XnLqFZebWSpSZW2vaHsUF7LrjWJeO/Oxi/gC2Hl6IuGyPPe3zB7HA/jpw70PRRu
aoTLopA9LJ+VjVuNpCHytEH9jUVuD8TjCEKK7VlqUSZwleHmBdbzaF1+EQXebi6K
j6wb5oUQS6//Y1OmfqYOswDJKBxRum1eqDr3AGv3AUefqKjLMngZxfHWSoJZqo00
hga223dBB9djSD7wnbbJXPUEvw2P5GuXvhQG5nlMrNqCTnM6Wm8FbE88CfFe42Wj
N4Y3Fck8WCcGBvEGqYQyethGCn/wZ2mjSgAakXuD/n6B+2D4dg2M6R2J2PcR1GGW
MAI7NGXQTYYTLu2qvL53kQFQcJ4ctJwr7mXMJom5PLMVusnkcjvo3pBg3mUiLqxa
gqWaCSc2iXURFIHf30oM46/y8rT5GTKbaWgQ9tR4WFkq5CxTmb2aYftamUXiwRzb
bW7UCy6S+BUPGY21q62x9eLDQEcROilB3av97aL17s16MAwforNeVZTp9zit/RtK
/3Cq1LlfV9Yb7CQY7mjLPEzTbKABA/NnYfDnwEQd+/1+m6tmO/phdX3han1JvQPz
WOKGnHlHThojhY3XTlSihCziLvU/OdYBXQT9COoAEfAbMB/YwFScclFrJl0r7Ciw
c9IrRTNws8Pqu7q0eyit0G7oIOmvYE8pXfckRcbFNxz8LD3A2I9JrOWLIYJnsZUk
JpePLhivrOZ3344NtT/3hSh4Yci9XdNCzDstPp7nw2MRjIrG8KMQ8fh0evOT+hFb
r+sAH6WuEDt+izuKI1LA8OLetg9BlrFgb6OMx14NYqiVWedqyhWjvHc/MoAXZDpd
npak8lrYiLfGgjpByZjmWCuWWPEVdqRkTeLAW4qSmTszmWHmUNg8AdqZJ4q9q3JE
e38MGAifltgWvrZVrPnsfd817NakXVmRQqdc92I+G6lKe5Mp51BRhatlK07OCa8y
YFd2bBnZj+SeoTgXteOFFjkUPfgM/Qc0GFichpT46fXFS0+B2+FA/jWLxNTMuKyD
3HO6t52K3t5/eWMGJczlEKgrEC+m5bvIc7nD6yqCGa5bHYjIi6MRwJ+V7PUTmsMJ
Em+Hd7Liyt5brzpgDdx94Brma9IijtQCjYnd+HJRYrJOvIpyFI562fatpFSn9zqz
GRjM4EKoBeSriy6m0lKXVMHobFHcI49lp7JRPoQETQEI2ckhMLN3gELj5nlEQtRD
EAaFuLe5p+PQix4gPaoUYebtlkUw/F7qedxKh3AFYrye1y1apmmAj+K2Q0VYd9EU
aC0i2/XjfOl8F1BhX5f/R7uljA0q93QWAq2h36NrCTwcjyZ8WlnhHKfxHvZmTvZ6
TjhF2FmssBvCPwhmwT8wDVyEQk5sdvDyxzf7QFiF/JicAVloeQGBOgZ7cjJa3L4Q
7cmqV9bUDv8l2cm983lQzNSRK1sL1hn2eSpjmiXZyvc0HnnmK5CucRVQ02dth2z4
H4tDPb63UDcXUrteMcOvYSezXUy440g48YwR/DtvjEDk/BRGft2/TBa6zEopgWKu
OZM5pV7VsQqolAp5sWOKwnFZbIBoMrg5OPePhRQpBgXtECSvBAGjyiMfXCmzB99d
knA8lSQN3wd1ZvNjlQTCn1SVHjuRT3CBFMn/TQsRHAyoGpdkuEy89enEcZCIMjtR
kfDbSXw2WMcwz9JwuX89eLrsfqNgOdbWopy1m6mAbk+oqnXI47YpNN9/fr053Iz0
LhKAq1Eyje//EWkqWLmsKiTwLSOb8306j8RZbURAkHaszfkPAFFT0L1/yE9nWZcv
/ZrVNGMjHp1n3JT5iyLbE/ffycCteVxqayoMf80kw4zU57kJBx9QfPF9fQRa2aeZ
TfxlkQaY1mF3My6egcBGsY1IfDnWQiMp21f1PyyTQn72SmRzNKlHWg3pWHZrl9YZ
KXDkLmdSTtwtkqEH3zC9Ibvqb9wt4bNM5pHeQYJur05Vhyc+Mak54KbBvUFTFTAj
OKgkuXYYkEZGlIIiDyp8BYRifxX2bU19QZfy1kO+iNAeEEAR3qfSsT76Hp50M/VP
cixCo5Dkc4omVMlG8+lPszYlZ1YTDTMzqHC4zjE14uF95DKJUda3qRmt3zxsrzax
aIb6Am4aZQ751n8exobm4KCZTn2P0AV8qX/5kCrITCvLf6V1YnTqJs3FPIYFEaj1
ekW0hRCRpKgWfMH7ZxfgPOV5Qs5yuUkg4/fwbWxH4qVhEDWHUlFH4iKT+pV6UqU5
oRKopsfbkcKJf8iTAD1CEfOQObmIsUbk0kN18uVie+7lckHAKwO7dhn/1WLfkcJn
tCNJUvXSf6jyz6mNQH4SozLoHT07SHQQr2X/jeo5vfIGFoRBWeP6tQ0ouXwWu59n
0qep1N8ti25oV+vzlUgXK2jvlK5erqOloyzuSKdu4j55S/Vy2VyeTFiCqBxHU87T
H+00pLnnHX+8o9U7Ngud2EGinlyUU78/ZHEgM4YiKa2w4zU24hG9jTUVlAt1qLWq
IKt0KxjepGH9tGFQ1tbp0llxaRJPre5zimkOYIBrFfRQMzNexpTvlbnrdjEDm1zM
7/LvVDac09bLa8ympP+RE3o74hh/aP0v2my9667zNVtMBYgAKTrVT0h+vXGOTJoL
IgYXotSFDxBF/u6YSYrzpMHeq4uN4Yyyn/Zv4z52JZwC0Tkft/EmrFMZ2lIUtkEs
2cNySJXUpjIdneR1TPbqAX6081qB96RHdFx8xwjRG0k1qdYYRwT2pu7U3XkWt/lO
/oTmlhRE9KsQD/yWNasiC6S51o7edmjjngNR3PdbUV1HLjByeouZJkzbNaaRnq4k
IzEUqvMkzeOP9OxWevYrb9EsKgkwWR2U92/W6TfxvYd0OJzrQ7NUpWhbVPld+Xnb
0TlQMoKcXUKkbK9qStwubZe9c/rvR1EwAVIN2NLdCYJTEHApJMRLWIOezrtPU2V3
hklTIigYoWkChwqdVaMioB2kA+XOyLUCEcKl8WsXJtBLMDWAEJu5ufcGsLghdyMq
mMZ6TxrQNyv24+HAJb54+vFA2a/+WiWf5NmvQjpyYwnbWRq3Ed2regl9jFnm2g6a
ApQ0SE9TSFNqHv3ML//j9ZHAXDENPFxsSF6rpBYre6poRIBkikaFNzRzFEMsJhAr
gNASvH6IpqymL7aHq8QAQ3r/o5hgAmAdMnOe5xKLrqUXeJQgaV+oiAuKft3+xvEr
nrGcpW94D6zlmf1cSWmF8hONXAwJwc2uk9P/WM7izqShYivMOEQ+0mi/nbPQvn3m
/W4Xhp6QDTg1sUhiNoTMZkNA3drAvZLhSHDJxkZcgdGYyBhHN1UUEz3o2UlYG9SD
UuJFOKNZHm9HmCkdXGBHZRnE115owDcD2pB+KPnaS6TZOjXVPxtfO4CH9F21nbt+
SuEBjE8YgxhH6Ue53yTIGCfheJCsGn4hMlvXFko53shOTqK5eZzaLabGgFfynA4z
/4ymLEw2dHa9TDRq+9/YHiYbs532vHgoO5egodauIdb45g5/7PwAmK5GZyDjNWZ4
jRVUWEcXUIbvgJPZJ0+jUIzb+DvDOZPHdyjsQ2S5KjKzoZkCujADXsYFKGTrfTj8
i0Y44U0PChyTDVRda8MvGcJEYiKX5+v2kir7fLwsEUTedzABUTXc9XbBu+blb28y
BKrLov5GZIfLlu4k9GgmYjmATR66xu3CARzxxSyCY8JxL/usSb89mlsLVrTHqMMK
jXoKW2fX8wDyhKI5bRuSWLSw+PVAa+0wHzQsT4s/4pRvnf8f4ahVrKFggSawHw8t
MWTpJVPTGJBv+JP9KbrOWEmgUf/gyuc7FQGCPY3u8p6USmXr6XovKM41kHFCB9RK
xV6KRVxSijrPJzVwrfwRKOOzsuhuBHfW6jCONk9fJphHLDINp8ulmqy7kOWXTpt/
mRFa03W3nDrG4nalWdpt6TQTuoHJcnYmyTkwlLawusohGYFJTvN7U1eEgYUEGf5k
8X/jtBGSnpeFMr+6+lP6A+CHFhYurUM7zjGJnnf05In45G4s9RAi2N9WcIioTEFr
jNF5uap2jFn4Gn1QvMJTPczekOTCysiFfcga3Gn15L2E5MdnMo/UskvJF1JjGaIp
0Jp2zEq5XFExXsL7oLzO7jpc+lWk6gsfpzxK/tDfMrqxlIvVVGBQ15++NEAA4H9W
D8RIFe6hYroFRsfTmxsiWL/6hS/QYOmLA11lydBce20tt/Q13aJ6XO/H6YkHpEZf
XrW+CraGe2MxXdAIQdzjGzIVq73wQnays5wWFc0pmrqhOCbazZZ67muDAYMAC8WS
V7yeO08syow7XMVIYlRG95QgizN1+vSJPormkJwQO8q5MQ3Z1bY9pNpU6Ocva23B
tC4p8EfhFNTMmlpb1qyka84IddOVoD76RrQ/AMRVEA0l/57ZdhQuieDavISMzUN/
xLmcJzHjkD5vfjlTteUinN/QVug85CoiW2Mb/NitpMr+HEF45mucLubofvNEt5ed
pzCFY+nHdvzUTJTNoocZ+FUxBjb6ClloDQqdLdc702CiuMxt0l/aEdl75+GLScxe
rxZTPDEXXDTaZENB9DLVaMEpF+b0A/lMsXki48/s5GT9EeZWaG0G5nBGY1tGkiLR
dyEmVw1JkFuSFBLLW8H+CG1UqGfDCgyT98jjbHL/ljizN9PbogTWha3nxQMrNfZM
ki8sUEsVGs8rUYWSH0eTNwUo6krY1e7B2sg321qENvKwh52+5NB0iP1qKot3oxC5
LSfau1O+729ucQjU5nEDShnURs3KnmHp4Qd6JVUzrgKnAyghW8WhjqhMU1zrEY9j
+jj1dlZi5S68Q0BisS1NM4sdGZSU3WfWam5nfH6tHYNpkqifC5FE2K8TYAf1w3vM
ItE6hqTQuckLhriwjWbIDv/U/1x1/2+bDerMaTx8cr5RhJIqem4RbqNnR/RZjDi6
sOuW2u1ZDL+JxlPKnV0/P7qN7ln5cJfR/5NSVWaUz72042jYCXV3XmwVnrLuDzHB
3y3i43PfWCz904TDIlC/xccZPsrQLiV85NnYewSNCzNeeSMsj5X53YS73YS2Mrda
DSiSInxgMOsE61ot+lVVFrAGZn9m6mt8l2t3QMEm3Io882D9B7zilQu7ek9dkW2Q
CQPQ7TzUTNvztp1Pkpo7aaHf/Ngm3VFKe2UEFlui3TVvlnZv/0a5NK6kPyzvDQ8A
pV8S5Iyi/+zMAbaTS4Xo3RfAFG8sBQvdPPHakGl8N1/ht00cu3bckwiVd2vtsRsC
CHKuuSDe5jou6T9aKgb/mHx3SgZ+1FM7D/tbYiMZg9lSPPFaOmrrn4Hd1Aj8CnuF
m7MqFz/R79DYs/5qgy7+kF1DD6y72TjLT0FhIiP9ESs4T6LOExNd/ZADzIkKxf2g
JWrhPC9AOOruKyOBwRfoTjUwIqXBibOuIAep3TDMo7xizZMuUqCI6O0ql+ziYzFp
O49ftL73oAWyvP0e8JRNNEdcu9qExP8K57i7+r5xApA/c9CEdgzuwrAdCfinVEUZ
4VhtsHw9SrOtZDcVP2lDOIH9xmx6c2gwQb3PZ8blg6M+BR//xqgjqciTRQtyrd/H
RUyEl7d8uygzTJQUw8VffEI0NCBTR3VL3S1tSlKs/RzQ1D6n5puBfkEi6MtiAfJE
FDHw3bQCffvA2wA2MEyjTD0MWzh4PhDwsU5L6uu84IYLeHl1iNCbDPYBZ28Z6oMA
xjgG+2YKWadBrdrsclQG0HrJPOFQApI0lzVhOrCI1sr8Blt2JTctNikBzdCzs2MX
Qme93NjnuW+UiALaM6XNC680An5e2kG3+8xbG3m2M6npmtjmorNEk1HtBLKSMgif
peSE/HzE60IS2R0mxoibWkL5WCceLkz83qAhGaLYXqCXQrVbv9qHkD3DD4KKQoPn
cHIGhN1Z3Q9T/fV63jO3s9OiS2Irau/jPfmr9Dp3TMl4ZJgI7V/wcY9IkKj4YIi+
cBnEBfP4GTWOCIF5/JXeMRSRRmBv/2ePFLxR4mQs/mibFLIOe7NLsnEh2+nATOYQ
zFAcOLrAz1A1Ou6yejN6Gxk9fLf2x5toVF9WDhIslJDmcqG60Ers2SsXNEWe5DAx
NUs8fpP4kDUkYX/0ddTcFDdW4PaX2hiqoaMMw9Vu/OAX4tNa5jMGWrO+xs2p45Bj
gvzVjRTJRTzIFysUFqIpuMgQGQoHdPY2IQq2nJBCo3UvvGAOv6SkUC7txcJp/jn2
Cn7T2npoxKTOR7Fi7j6p+q5czWfyMCzGxMu7mcQuiJh6cuMJZcJ5+PSy+nbjOEgJ
XD4DvXTmvcCAhvUN+NRpG3QZc9iWdl8nkbpo0AE2gm7pBGpEwkThtzqSY4ocVlTM
Q2QyyUXVWClzuowc5uDIkFu7w6ntfLZiVTfplmKFV3KEgN9HWtZyz0B2eACSepHp
4z9m3lRjU2ykpHrnXzeDqfZBEBwj5YGWmRA2sw7wNjPFILwanmJCJZTi3Y45fWfE
nx6i4thECFEoyfVCigI2JT0kRuaVmDP+2k9FOD7y1F31h3zx5FKHTIkhN8XOGg1R
oPbE2EVTE3zGbP8O7lL69RBrTRSCMZbGR72dekmcDWzP7cR516V2X/QCWcPo7Xm1
gAuKp9e9ttyOiJMhUVRU35No0K5H2XomTH3yqrA3Gs7yoQAy0ZqcjzyLzS6z0PDt
CVDX4hELZ+m9yy0TFGE7jsHzrDrP99WEr30p/WzUiA1haibWi4lqUCXIWzmtt/LP
ksBTCyCQujNA8xOE+HadJR9P272PV04pf1nki/kdDih4NjAc/dHUjnELEhe3ZOQg
W/GBA2KDARgNqK1ggp22veH/kiM5CTb+qgJhjBgkZwFdpZlADq1FSQTElrE0/M+O
l3ihEejgAWefYRjH4eFh31fxh24ybzYAb5HtlDKD6oqgOnnCjNHKlCSbTbMxKJJY
zhG3XZDpFoIGUQ07+vqmpztB9Zn/RlJ0qmhQaUDsXaKxBwUvv2d6oF7Nobt/U/97
IO38LZGme/Kppyey/2ogEY/qy8atiLanwBtedZOtOUqBC1fRo3ew7Y6Sx9GghQ1K
5zeL+Mo+aCsEggRKoyJ/M+aMvbMRC5E2DZ8sqamuNCbDahvl2+ZHJopoOAR2eUz6
aZtRpVwa5cGdvbQ5uv5yhS2v/4ejEApPthmAZRgy9rBKpjrZeUD0DqCHTwPIHvyl
vPyM14IXowN24z6hoGktC43W3Z+QBLtcGxGoI0zoBut/fnOwAi/LUkGvjlLmMq6T
hTZ5b191RoUpwqVHulbuYv/wizdYRoTwErh4PMY4vqkYObSMYQW9D4SdOfvgJ5zs
TUIQi59qqnpAxoZEJhLNEIuhYbtE8kOmT0nT21TkhG41gVcYfNIx0wsIqMOoJYEE
0OE/mWiXizKa/b9HB5wJHHLXbSFk1Qq4hATfq3GvljXjc4W8gsr0BmwBbQekN45k
NAX/joUNaOddrO41Uhj5ZVAI3nli84GbY8KW9f5MHqvOxkkezmG1dPMepyuyiNbG
xREqjv5g7kdC6UgcdKAXaMEp/Qf/0FFsq/ggLWinWixWP5Pi41M/+E0xGqLPeOTt
/py1coSErTJdE3saAj5QEv5hbqcfD91ZwRxCrK/u2r54hGaVrVu8XSNPBjGr4FD/
amiJqYQ7Dii8zjAoZdn/DZvywk/MAmgMzwpN8+PrVYkpQtiGuwdmWdhaNXetaPZE
aOdqSF9oiqlU28fR0nHRlgdFJZNdQJTZVAkz8jrcmA2S3YdBBtBv52opcf5TuTZ2
27CVwYRj7Mx4skZNwkhexISY1RImxG3YOl5Dd1Kv2/GwdKcl/6sR71oZwXEzDIoi
9O9utqESAI4k7g+Pyj+mYAIQm8TW8w326T+FSK5DXjZ3aMnkmFpTRXIBqfPEHK19
IGJXhk3XhoLF1FZSiIyGCwbXyj7ze/UiCq3hiovY49dyU8OgMVkaLHGccGohnCUg
smWINTekyWW/JzJmtjn3k3/pd5bhKua+uBr+ad//ns9oduNIltCJikmucB0fLgcY
CCd8EqU5wQhVCTcfUeQBAAazvnbIzCe5t4KqfAwE0dvn+esgF+jCzruKxCkhmwfO
aip2MpIIZOY5QQWjDqn1MEOLVEXq3YgjJ/7qP638WPjShwerqtz90FzOFd5HRhZU
QlVaYVikyrbcglLLGmpk6MFoY2GTB2GrIbs47Qt7rw0rJIon+Ucp+/+/EiXyRxrc
9CqExAqz5iS8Ra/NsrVKSsxZx9UOrLoKSOCXoTLAm6UYYi9z5NCOcwbPXoVSg7UJ
8GfFN2LjsXY5TlmK65wC69tPm2MQuY9kS39wryC2WNRUPEhnLcVxGmBLwJ0+4OSS
lsUCIF+zgx9h49aQqJgg9OiRWb4Yxf466o6u4EId5IdQfH0HXjhi36xuHVrzgWJV
bdW2tRVUz9XOIRbLbRyfGpugp6AlUJRkKV6Xahn78PdpDYOX820E5nJ0aJPf+HxO
fzSSpL61+h4+zzzcYyMkCaq8Az3345cZV73AUn35z5ouN+ht3Pwm/2Kh0stwZTkN
MXJKdVlFdreja0O9Kzbd5qr2kC6E/70f0xDi4NFi1LEzaxWROh7FDkxxIJTBQ7Pa
g82L9AkOYtSX/0mceJVCpPQE3yiRzB11ubtt3W+hFYKvxQ85MaR1gu+w6kpabMXG
KHAn2ZfoBmVZMs1bWnZjVoBI8lF2eacTlLJYhhGyKlAUK7kRN3RV15s291jPHhf0
keoV/V+gfPSoL3K8cdgF2QNH5hM/c3PZSWORhYkNcbU3W2PhuEmPim383J9yQrLP
Rdia0i45Dz4vedQidxawjv4ycSYQh6iVFqtJbheNmoExqk7mwvvN/UlMFOYzoVYR
TgWL5HmCff1zu7hcOcy8wV7xJxSyFEzH0cxqYxJyBU5OJJ475SpzBFtJQ5YdiBmv
3IAzjb6PuCd2cgqf+kt9mcJhVRi3yyv8XvlzMdE46FOL4jyWVdNrIMLw5y/4Kcp4
gdKvrXV5JNpvVQPZ3RgXlRMFWosECO4gZQJFWj9RdCGSlv4AAKU01x4jwlTA+A7J
YgeEggLfvcwOAUwp8DoeGFzqnEEKB3xcynuyKgd+jUNINjpkX6/JuLd5Vzat/taX
Ws+4p8JCrGgPnyxeTV8qtnLfoUftwk8yBFPgQYJYzDwSRC5mD8Spec2buVze4wcZ
aAcoj5KvLp6OJUOWkJKNImGpoBDx81x2Q/E55lzolDc6yVh6EIyzlpGxrsL6Bj1k
AHw6bhyzI8F5lMUcIZuZrgCsRx1+rpRYea1k7OU3hxLsA+Eeg8gnybPqVKt672ck
Nwf9+0iKmdQRqcxwyE2Y4sp69NL1CU1RRodJ1Mm+hXa667EVGNkZirUOR896rGmv
LZrzc7r2jnNLeKwz6TEzYZSP4qVy8MleduMLJmNzmeTYrAN7VAjHs2aVhVsei95a
+oD4AQLEoFYLWI/EYRink83GNBUSbweokbqPb0K993PTG66wcWcde3naZMNOJyMY
O6cefOGQdNO2tSYIgMFNNVDI6vRD2ySoS2NGaZPfInfHYSQ8dv+DxHtiBEDQeckO
WzHPW9QKEdjxQLkRLtT8/gr4gYj3XshdPdSygQghv5Kb4VJCjZjakC/JDDLcXsWc
RP8XhuarUMrwzLvsbQ2/3KC6ziJZFuw0IXWGHnQE+8AdiwRBjY18pcrpwNjG8RRs
vQCwCiqiy4pU73SCqFrb2dD+dzAN4zUJrRoMLDtb86F3RSZ9Go0giLdHk62zGn/u
vzw63zfeOAGtHx2MLd/A0bmD327rW4XW5iXSyUU1rIqXTtkI1DK+G8d5lkuoxCjE
gCKvgO/0dhN/v4uDLtiRVkL+qGNu2D6HQpZTf1gIERKVoR7WTivtMD5oZo0CvBWx
fIjRkl8hDNPtoCNpopx+8hBu601THqWf8dXBscfMv0fuH6f7QpfB2ZLTerdjOED4
OoxjVzV6aWa938BXX8krNVyQ8QkjQz8LZsmWec61m7KwzxvhmKy3Yj04GlFTpx0N
pNnd0gEdXQ4P/YjXtrvD24Z1irMTVCfmgs5QEt2WOEDYum7vOPYHqhz/ng0BDljo
fgnC0a7/toU10O2YgIpFL6Q2DqNGwweP+ITtXupY1NI3kPMz5iOIEAoSNq7/024H
0o6EmrxCMYbKjmfocmWtiB5OP64V057qvDdxnbkOh5KGWykjnkD4JRI4o5D5TLCf
Hgf2nCb5oAXq+nNwXb1vP2zCrU7dQki4izq0TA4/G5N6Tfm1bH6uUC/tPY+8Z/nK
3kow6OkfjcfK1cLUiGc/pIfFjeXX8dFvldbkCWNmkWPvaXWQwZrCBjbf162dFEBZ
qDPgHzga5v3KEccnnE+PZ197OSWIaLs19Xh33lbmtxcxQYreaR/P1HdhI4/jvaJc
W3RkWNNpRXZrcNxPfZKD7DPdUd9yh2+J494ExvnEEhqm8ZGj+mDVOZJPQEhCnchX
vTZVJfz4xfyiWJ9PuWdIB0wdyQkLvUTuOyyr3ZxL8sxH3T8OoXHPSEYRarj574VC
XqraYs52xe4OmxVM/1W54mlGE2psH2xZZ68KYWivalB4kZopXc54l6t/9q4XtkdV
AedarJTa653d0WFSGH5dHoNWugXTuQFNjg9yq9S/AC4R1t1Ao9eKR9a/HifL9Bq0
71/WpedABkwwZZOBbQSRnaJ5H+B9hYJ+14fAt0ReKNoGZuwqAq/OsjRiWiShU/VW
M6E+qvbDrPuS2O5ceqG88JZMRS7RmeaBZ1a0fRIf+Is0gIDI1XRRj3+pZL5zZz9q
Rtg0KpAua3tczOzIjFIQNrAxH2o1K1qAu3oVuqaE4fJDQ2cHlF7QWQlogNWP6VLD
fOg88JHsfkVNJfRkyNqj46gOyL2tqrVaKrdjVELdur5lvj4TsVPJpntMGGJLfL2z
hAhuJK3FEr0Eh9aNbhibpmWRePZqiKlpt39YaGVtuT5Hv5tzYAxoeggY1UtGUjKa
FeyXNUsF6nYGoGx0Jq4hdiixhUDzGy1JywF+o1aPatdco/VNocaVgm4LIGuX3QRM
R8VEo7XZqpXEKYBhEVXVkOw2x8/TYd+5W8ZHDIp9VX+emdRf1+KKbdYpq/Y00kvB
5sHsY/c1iVJCSfFu/v2b1BkWScDieVxaP1/N76IZA0eYTWivUFkbDitWbPyT+rNX
qOSdeziVC1QIj5nIV/Sk1oOFziU2LPrtEfILXoYRTYr5dbWZmSCthZIymFB4ti1F
bdQ+kpstqDdv83wG5adgQJGEyKPULo//zpTMO5fCIJ4NNBx6yrOMbm80ukFbahXp
1/NQl/g4+zyHxj/T+52AMzfdOJW1FdH7CzW6Y5WIH2ZOzKBROgkrAGaGAWRwXNWv
5ggQVBwUy2du4VrOVNlQZYolgt5pOATSqJPGKHV6k1exauOHmejx53Uyntv/Q5Z5
Ev1RLRRsZvuINU2qBOw+DGSRrD6lsyjeQHhRbvhcTPQl/gmSic5XLjblftqvFNRf
/7YeGajkktnBYwzaN3L60Jt9Z1/AE20lfF6RZ/XEiH7wr5OfuNAwEIytYLiLSpCB
+eWO/oH6EZ5RusCxyZe6jreLPr6KYwJGJnY7t7h9pV2FlFewCj1U1e4VZ4UfnB7V
LNCJv2EoPQKpr1UmZ7rQJXH+HUCsBATRqIr5CZQAIX7MQdSZtMqUMrJaha8LS5Qu
EZhyGwJVq2tfSLe2ofHtI/OgpUjqq0e8fM9gIyJzb2Df9GAI0klishEZSSWQ+FVX
a/r0+1pj+L1hWkGRuL2ArC4cpPWxXtyWTp4JMl5lqBt5RoF4v93XQE5/nq2UIalp
dmkN098A93XCS6MOVIigRT0HD4L/ARg2t/xlv1osmIdgwWRYfV0Hgc8sjVnqwwYy
ijnyFI/GKwAtOM1l0CFoXCWePVoTpb7o7XuCpaxueXsMrde+JbMglHfpeiI1QWki
z/4EQDJQOCtnRlmnV4jR+LiY6o9uTcOEfiFJs/6vIna7sqRm6vCsbPSN4n+Gxuse
KOhqVl9ZrY7ZeajOthnW0ebmukVQH5EeitpVtDV4V+ZppaL5MLuXC0+N4JP6EDjN
JYg6Yl3EA8fdE21AQ3CXIN2/4LFNLcvm0B4b1CDfT7NndTftta0slbf8qfEBF6xa
EGxlpvFvwhpSThKMm2GYTi4ZVW8m47CXxVIUtdKJbttJqIloW3OH1x4Q5oIDThpI
b0l/R0cHAJxo2t6qTywUb1bvqKDRI/nS0kiFIk30BJmLRBHbjYw6edH3LNjE9OoB
vRFCcazSO667qCo3bG9UFZz2w9M5svl7SQW5RLdljy4LFHrZqj052E2Bfho75rQ/
LbQzoyRgPsRbo8qNkOrldbcmyISDqbT+r3n6Fj4vioh5IazQ0n76kwiFNYcEpTIJ
dW9phtK52SoWwUr3E1g2PIUj5aUaRz94WUtJmxQFj6Qx0sbPK6A6ugziDv+bO9e3
kAEqm8zcYutVURfyXUktw9i0E4H1JV4AF+wxfjOEzRZ/Fa0ahroI2xkPeyACR8Ui
HgdmL+VSnqR8usU7/5xoURBz8hIJJGTp55in8Av9HHa+cBkx3R/sxIATiNk7248s
EMSyS5NHaVvLENNy6dDWUymFQJYMEgFliHMjU/FwCk19ZyPqVwV1/klHI0ZtNzlk
X5661o3Nd6q61bcjCxJtPf6O5Ra4JKoH9vFq9XlV2VN9Rjvx7unghJZyu34eIRJ6
B3uhbBg6RnfAXHKkVCgPst+UgUz+RInasZWXPklgNaNEKtwfw5l+wgT3jgcdL1KW
Rx+9YSkGlHZ6kFDrATQwqqXkT+ld3kPLfaocZcEGzPcHo/5rhjcfgKhtb2xDCDHh
VdHx1IGpYVtqiBhuXS3nt2WkepxwJ+Sb2cyEYGn6wPQ35EjBzzQWEefNpaUnJyMT
rXNSOUH3PXhkaBcjY3DoE1P1ckRRWSGukLRKMkC9yh33ryvzzI9Lo+RicB9qP5z9
iGyYVokkP3bKw6lLj2EpRqt3oDYxjS6quQMQuO2WsuHkLUlUBl2Cdg/wMBi8pMat
bgdBQXwK3BL83/LEsNUSelY4P9d1+CLIZcLN3Dph+Hb7t0Zy+7iCeaPCVnYs31HH
t8nrKNRoLHCNm0cCFmrFPC7sg8N2JXg2s/DvKl3IUYW9kCsp/nrez7LF8sd4kyTR
4xCtq0sSVuM32cXjor+iNe/+4reFKcJVsbufIxLfIMbw/60/PmboEUaj/ckXb9F1
zbA+4XOhCZXBfUxbuDiNkcNsVLtLO7jpm9BUfK3yHhtCxBXp58nyDDqfbuxEO+L2
9PKD7VtMolwD+1kMyeMTPffFXbTS7nPsQLAteDbujqrvDMa3QsNDtgS/1BCMqiZx
kfl0nPdz9Kcfmph6eblM64pjDNznDd8/EfiI8iNBDd9GEn5agPEN52evkOirZiaw
pKjl0Vqs3QktVXSKthmh0QNq5j4jPiywxkkMNRsYw7VC/XWs/2BhjlT9TL3HHaOp
8OG5TKyEVCfuQYi/CXWOKOTQ41eEuAkHmxqI+DXf4Jc+53UfxN8WIgVFJ5/p3STU
oY1WSmQTA+/VH14MxQ5dkKSwTH9AqFPKuUo7MaNXz9duUd207XvAtmH53my7je11
+K2HqI1WQ59+NiI5t8rxUbTVRKyTZQMBAZ1uv04UrQV7tDXzn+sJbJcxA5mFrjdi
p3msEfzpFiqYqMqhDqsRmJlycI+4lJxr1bInkzYrHtXefagmH3hjCnRwjAetqRK8
xbkB9/bnUHdBsw+fFUOcxwDVBUP5p0WD1IuVJHj9AZEW1pyNsUU8RVJ/A1nt8aNX
5z8Eapk2emN6rjPTDOaAzhYhRfz4GeB9DOnihRy57qkfg3GOv4CeapikSgL22xcG
kncTmgarUGVY/QICXJlEm35662B7IMN5VMRqJWFd2Wqza6LMhsIHSUndJMH7m9h/
azvf/6AWKHWDDLszS6lSPRC5dSlZRLLry8o4A0jf8BvdPDdB9fIX5e6YVE6pPi51
f40zteA026LDO+Z6XE/UJk8ToYudsKsaYR9GxRPOMyaLgQdcqm39dNyydElxbFA6
sl8ddYn9vwvJPUIv6Thw6DPegjjnaTbOvtu34xWPIk6N4ZY1O4KcTwR9828Y+yCg
5mzMjxKI1VRTcH/faBLihUPkXdyVZuoDi4dHDXxWeHi0ldV/6sPSunwPPcx+79Ei
Wn9s+7IcHV7qHOvwIPxdAuFueXgpasyiejqeHBq9t8OtkntRMLg+3cGa1192kyUb
soFloqX2eTioBaEq+TwLZVL1hILcqjIdK/J6jiVlPkpgSjhbAWK+Akhs+ZJVRFw4
f4QZpiYfLDaRng68l7z5rAsClIpgklrcKgi7uQYaRH03lihHXgCT8RpHHxI0q7Sf
D+3Xv6fjf1uJLQAb4VorcQdoXNFwnEcmZ/ltRwXcM+XBGnCvw1kgm52rWmb9q6By
LDlo0Ok9nLzU15hBpWML9N5fKEhvDOg/AJsel4qBrCz07JMbE2jyKoWxF5p6ALtK
zm0XIm0qhFjvzRwb/yCdvcPYch4s80og/ypBOWfv7peDmMNIKPcQYbvT/KFM0NVB
du/4FNsTya676MpXknOXbUSw52ctcK2lgZeTPfNpxlPs8AwMQp3SiPfX7H4CJ0qN
JG23LfV3f4Ax549+wtjtHQeZsYQ7OVukGJqPTrK5AdGINET4+yAfvAtmqJYbFWI4
GmzaPTpv4/KMLGa2qpPFZtDX7ynb2EkSnJe7fARy0USwMyWgKH0Xfp964pOzDa9i
m7pggbMRmboxH18Tp8+09fJ/BZ666aM5iv4mhK3MqY/bJP/cFJSFKGE6RWf0KdAl
vL5xdtx6TA5Q83VlFpAS6hvEmLjOxFF4aY0zEkopFNXn8VXbaUSirPvy4Cmn1f2O
hVpfSPXAahGDfIJkVIDsesExEkv163rHGYxIr0rXvpGVBwjEIkyElefDPAomc21d
ybb9E7VhBSpvFyZQwHJVOKd8OIz4KiIAZX6PHmrIXLKiFczpdY0UdLHNas6S0Ftx
edKIe91OYj8/xHW28ooSTHjdSZSUwC/5vX1NTll0myFhiftCtWBw76dMSS6ZWZJn
HgUFgpwqtW8DlItjzGMWlMoCj7jt+rv7SkohKqTjFrJqByQZSJWAoW3t5s1Smful
jBy7TlJQ1YzNJlKVOOst0a3MP5HwiiS7xeaBVTgp/IaCOhcIcuxWBdLzYAzi0ja4
Vikd3uHJ6L9a86Y/X+RWWdlvSXRqQU/7zMA91fIGtJQdhiTa6uDYwfUz3OG2JqUt
NAzucrk2qeC0pnNXToD4JDCIIkyCPFjKHFCTKBRgYBfxd5Ikh2NlPvDuQ70GRFdL
EV4oyYxCyKbp1Bw5pJENCrNyNz8dtEDAv8sVB/SPAUUU++SMNRi6kSuEX9Ln8p5R
Y0vBTnRS+l4g3XvVVKL3W432C0dqdS+30wxA/3KOGGKmP61BqftNkoJB6m4jc1oY
YN1TMIjUmBfmvgd50nXQnR6aw78IF0fDLKNKP12gp6ZGZnH0XNU99jBGVn3JiOsi
5od78Ur5KNayQXOw7CWDILg3kZOuNRR+VkaQQ59xSNINaxggWroq/kaU5pJrwbra
EzDL0okNb/M6NKYlQAlqol6UfEAaaa3zMY8xwt1BUgaemzwfg3fmnrk+1OlfkLxU
TauxNslQa319rexYuOLZz+spHOe4dyOEmmSN1Wi75oAX5w/rTQ71fGaR1E/V0jcb
Kn+5ZapmkWPjhGNdKmFyI+xxEeuDfT/qnzpK/rvzEeEpoa0MFCFloJGmXUWi6Mi6
FVEKi8GjeVkuEN1dGR/bgoi8qEfG71y3x0ifQnWN83iiV83EgDmiAxbW1GfuTGiQ
g5S7Yn+Ro/kcaq1eT64LnrKVxdAXSHeRF6DpoUbK7bNFcUrZGjjjJ8jRs1tYU9N6
72be/jZT3jSShGuTFP0t3KN265NYz6DVxa9UpAuBWAzRNxtXfKCTa3RBeGybFeGZ
cC0kvHZGDeI+8GHqQz2SjiyiaPWAk4XWgaKbdEa1X3Nenwpnx/WK4rWgQkvwfg60
I0tcAUfWs0F9J0l3dm6jL835/7H1FUlqeCBN/n3xfzktuyIX4u1PHuwjQ7r+I76o
Ups8R7+4H0MH0LrJd48hY8kYfAAbgmvfqOxjF/2SKjT/GEOOWSSiMicyDIfj17j0
ObFxiFYYRTzAl6eWSZc08Dlqjjp5YLuYW7pye4MMYcgbfa+sajGZuvAD3q17QxHH
4q8WFfgZjrdg1Lec0lMhnSTZDHHslPT5TYSgxp/2G0FaXGll31tXcQ7+z2WLfNZg
g4mEUTQUDkrH72KH80mFEuU/waHjFMNxvZgm+X8oIH/jkrN7qN+RtGzyAM1xzKJM
1hSJWqU/8jrPWzd9gVGIj2Xq5rcsQ8eGoSYXrL0pQSsJIGndCGzqZvl9LobIiiM3
/xAs1I9S9/tJKiKfxgRrUvMuzBQOBF0h5YDIxBeUF5gKwueMWZsDl/gfp7hwnkLA
aKHkLPyqbW5cfchNDOjroKurwP3zmWpRIOjGy/YOF6Ov7W5jhf3E/pO9w4JmQyH4
oKetV9hb5DYrZDgbOTB3iJVwkPAc5beomwZf0a/IJ0XNfm5R8l8LaeYZe2hQEIWL
BLcdnw182enyBWNAf059fttc2ISLre4rPLWy76lmlndVuPvumqgDwUB+Ms2pDIv7
9JQBh05Ui+jss94C+50ahIQmCn8IPEf42ZVnYgvsVAwGFpnjPrQ9F0CKClKUTZT1
kboi+2xo2nHeZsOrBHRkdlzfKskFF/DlrOlucAM+R+cB6Uo83oU+6g+wmFXfGv4z
WVuqjBjcgGjAdrz0aoYL/IXpOIaaYEEzmzaMZEUIo0RSFZe+OsElRyPdTr+qkRgg
BRXpY54pdhwUKpdfEqbo3n3t7jkHv3wkHpaUOiBJ/hke7jsjzX6IKyQBoNqGtS9T
MG43R7mvgmp8eSEmowUnQpYDl916f3YnPyUmfXVo7jxCd+Bop5i1y7WOG1RA0dk5
FJOZlvBTd+29I9gFV0PmINANlku2zVdwKRairdsFmWi7aSnEgahsA6f/b2feew6A
sjFLHyzPCOxtuQzy2p7axzXqrgqYlAjK3jxiW9QKzoVsEHTcwLVgnxFoFk+Q9rpC
KppWWQYwRBjNMB1uW56orU0vRsfT1Jh0Xtt8K+L+43rhzR9Dpnr1T4hriZvAB5cU
tova4vhwk1LNcluNEz1hnV6zPBCmpHzezhTFFELDlsaWAyYfTesBWLy/CvKVUrAC
e4ejwvF1LpdFEdS6SqNz66uMMiMfFxLPbeTeMDsxjcOS1MN8r9ZTvlixluX5xEqb
Ehy1AAuyRyb45nAWHkjcek1tnOyVR9dEiXEs7fOJmoBeH8L361rTV3UpjEUEPxlp
mL2ohCQ3KOOg5ZrtnN19tFND9vMWFNnf3aS9N0QlP+aPbOPrYLR76vgirKtd412W
cMIRbun5+Ga2oSfSX05UDRIj7bUdDXaIdmwyMBr3Tw+BoIFPit8JOzUYeyCKAVaj
TwvSAJdfw6ep0vIIJQolvzyyxEkOz3/2plCDEq2eKdwISC4ILtdS7U242z+V2AZ0
SJPxIRHFQEE3ZeSapNeEIUKibeczyGGFDlr3jOhT45JXcEQ1gk7ACIjGOOyJa8Pa
UDOS3avSOcQbGy8+dE2767j/MydQPBDbulRtuSJ6HiR3vwtW0b0DTfy9vxsul15N
2hgSfspiFS4EYZ2W7FUIClh5dGlmBHhL1W0q10ebT8aNCbllhJwpr6z/3mo2IWBm
+ljU1RybmcPI0wN4oMUcNqM0jT/tPwuXho464Y8IDhWeqAeky7H/GuZ3hAPoVZ7o
+LYpzwI1Qv5KN5P1OX70jwBxO4JzW6Dm6caux9s/I4sWoKJdcNcE6km/SCtyfeKM
LKYyK8fN1ZMldeBK9+Ja5upFYH0h5kB9Wfh/G2UPHVswSuDlwO8OhlDjhqwGpj8M
k9EL4jbkDPwEItPUGZA8MfwJ+GDPG7WrZf9JVESkS1ruN67qt8xjAHn4bB6sZKQz
E/xt+E5zUDKbSfO2h+zK9b8unMjq5S/TCtOHAOAO61bO5jo8jTvrh7edoc8x2cKp
Yz8w5PB4x1t53bvIINDQh9TH1fBam6Y3uEH53+BlRntZGRFDad2n3tqkmtQ8pSeE
DGyW4fytxhp+j7Yjb+GlzxoC2Bk6ZmAlJpn40OdysG0RsyEqeJGdA4F+QrZHCLMK
o6CLJk8ovF5NTYldYGzC3HAj5BVLoxS+hnGOlYVQr0rYxVqmaP88w9FEwvuju4I6
1b1c0ZJ751XxLa6klU0oVaol28fL3vjN4mceG8/0ipk5x4aXcPrQ2lAWgwfloOus
3SIjlN5ZGTosUXyghOJTInok5op+pcoqTpySqPMUywfRRSf9QcwMJODbXVZoBrLL
Kr4KSYkpY348VqdWAAMT9zvK0I5uFKPxKzp02pw0exYt5uAAS33Q7RKovO3ZKKa+
Xpf67x+HLGQ45OIvIV3jExT4+L6ewsPDFTL1iw61EIUlAZLJKe4zHS2vQnZTfn7a
cyh4lwNigdH/h6/C+tL9iflao4dKkixvrLGUbYm3l2PbeJzmynaw5ojiBE4Tcus1
HSGfn7uyukvw+E0SmV1UfiKa+OfSRPxPnAZWwwm2IktFjxrMR5Kp3h7IF06C4hrl
pkYdsrz1Sc/B6YIea8dn/TqsTFQ6tb1vA1tPrzxPLOwy1OZHoSw7Cwpuvgu8pKhU
RYfaoIQtXuPbLu4ongsn7skqrHyHqMcaobAre8FFu6uNEKu5hmryt8MmpZuC0gSi
YhSRGSc0v7EkuUGoSdK4mZYWgAKcET5Lvbu7ryKi53IAMz7VsDpeDBaBxMBfMSRh
5D/gjxiFX8Ili5WEg6aA8KtzqlzTe0akaTalNziWHamOp9gNOZaGFD7HvLMQZgxl
9DW00z3OGAlOVfcfR7rDr7cLNqzsB5GMIBLjaQC8RDnVEtShaL/DmmSXMrO277nJ
e2MKkcQbqeKPoNlsAtaoLNQNKf+cPlbBsdAKbLYAt9b4FHzI3t/XGNx0Mvi/+lsw
xMSzL4D3Oq0UUkUahzQT7VNujdmaLBqRQPphWLEAommv6FmPKHSy7IvOacLHfsyj
J85B+YJF8YXpQgVpcJd/hx1YorFqVMjukc+JeUGrc8JcW1Q1Bj0UHsCjeBstYCmM
RDW6mNuE1i0a2crDyV0XXl55hPdSnoZqOq9i59KVrJZ1j7HN59aKJMCeKw3WFU2v
jdQGihw/e6nXosyjcDBOSHmTAOM7Zs7oqYWz15LSk21o72NjqLBDn4RRu0i0mPY/
+xsxRxUx5KSgYsZGHRIc71UugivBN1/Q4pdgWmfS8Wu74LEeriptzBtH5DBVxt0c
4xGx8KPPzTlNwBW4/NvMrjYV/5s5fBrfeNKG/PKzwz9Or0tal5pIyNFieFNOamf9
NKzOriCxuBK8ugAqZhqEOyvefCSTKUeFTwaqaNC+Yp8X7ptEfnmAvKq0wP7Lw24g
YkBgsuKatUDdDQeZgd//JQNYtbyxqOVNlv5g/uyTcp4wckYueP1cv05sdFZmZiFw
ZLFnALWt5vz9rTb+gzLbsKaKQ7NYVuGyIbGhmH++vIvYKLVS4AC6YytZu2kcD0xE
JWiPr6A6M4bYXK2Wlk42pBQNjruc6jyHBDADQDae88nZbxujrvZycYc91EK1/bD6
vjJH8/w6mggCZw05bknxz8wSIdaPkbmhMAnuY799Zb+8lkcmqZHN9mepBaZXuV3h
zuZCBnokCv8BkkZJD9GJl6VjIPLUZp99ngCXUmaoJCdfhx44X3D90keemq3S2RUM
VCKCZayK0mJcTahx0+2TQGWEDboMHm7vMRR/n/FIYYCmuhvPGpScFV6wBGfLWcd/
dtBp3xwUN/22S4QkrZfuXo+PCQDlQEOyC7aw3/JvdOjFxEfzW+OYatBj07w4dho6
Va5KEigReYMktVI6ZGDy6JL7lZ5vbAu6tWPz4a5ZxqBf8KqzC6HGaMxcFqB7OW60
xu5XKcKvXevCSt1E1LN0pDPuf0z5SOuvkAQC8lDNH7psynqNjiB1pT+JLZ/43APh
8m2YTjDOl9LYZX5pkzd+uubpBF5nifVnNSSdgt0IA+CLf6yVvFRP6QfPbbgGPQj6
92lZC7ooMbOOEsLaRYJVdKkriNg1jy16CcmsqqTlUK4MGiklskJxbyN4KZMRu3/a
MayW7kSbUBJWeeTbSvRv5Z/q2/xD1TlJ43qvWIRQwFp23sMOyso31Af+rG8BwHTe
U+phKXD5N1XzJ1D3HG9zUddGcR0Qf6d/W09kWSH8Yyp8nLMEA4aG7+xzLO7rCSG7
u90BBUwpy9Q2jq1OpL9vg5E1yR8Xw+PRm03YohLsJMT54qx7LqUCg9lb7gZ62Js+
3Y++87SZTOFztsTJ2rsutQStg64HTnM8o++zw0BI/VCK419CnwkjjwsftSk8RTeo
SKPSG5dnF85dE+4zMIa6/4cauFkNSbF/pe1c2IgvZT507enVV9hwt+wxtUBgPjtn
925/5BaHfpKSEVAhiL+WVIKf8+q6CwM3LnXmMHFGa4XIGeYN8ZZRYr5SDW8bjla7
1Y0rvmn6Qzf8mqS0va8sWqrg7g+GhZY2yMn/A1JFm5rcMWKMEnS5NpPTbqAY9qOh
/HM7kaWTbnqCCZGWewqZyrV278ewNQuvuqEPGARvynMycJWAETfg0xvDz+Yw8tY3
p1iFGOtowTxKvRIBBaVyzR2r1Y4OCSKfixeVFJmyTC+iqzVmbPqeCuG5T6yaxP+q
SKd3S07lGeIYQjX3Ukkzp3Ux8hbFxzNdHYk/aE9TPn4JdtmsSvOB37KDJOEnG/ET
NyV2hsWHAa/j/iSuMc/Gdlrtx/tto02yA4fhvKUzhiesKtFgWjoEtu/Wwkn98ulN
Spm/UwJ0SpGu97d3loAYkl1GjTVus/P/Lv6dkiUKT3CWgVEjnww4i4syR2a1/FA+
qrZXocKoMJaSWlwdG0otY65hxwY6OxP9IHtBMg9ITrR7HpovrVtTRBY6amKf9hDM
U8R0SM4ngC/fQHQBHv1s4I1I+e6q0CD2XcfV6Qkon7gQplqofF/2/BFtkqfF82wR
6ANZ+Se/c73EVvnZVi6wWCtIiWAMRis3Qpww5kgiTvIrkpWK+q+BUYaPmf465QvH
bgYODKxvuG6ygoMgzqaJzMxOZ3qzs8BsC3JTug0erXE3wMvAzgu4wLqdmtv1biEt
t6T7MNVDmh4NZlKfe91OnvX/pHXbnhSYg1ltyBU7ZmR+LKAqX1fV5P5MkmfHXBb/
Scj4qp4i5c7lV67ZVhXd1a042rk+wYw6TDSfQRfdsFJ/o0rUyN1k5SVQYypSlf0N
Y0CZXRGDEwd4sjD/u1BG1Ax6sS4TbeRVE8/DHSirpcG15vxO8zkimvvdJhI3b9bf
KR5yLRCSM+k7xlSJNZKxYj0OFT+dZcsfgkcXjZEZwH2voRY9WO+IcCWEl0pdWpLm
cspJrPbQcCYeiHnf6wftPb2oJPhmiYQIxjQ97uSwHY+EYqcqG0q1X4rFMSjFIssD
qJhQ3iNej/AOyLTvw2a50MAQw2aBHjUw5Z8SGQYsOBr9eunSJhoiZ+HDHHgHHKIj
lnOx9KxKdYnaaXE6BHgZeUXBrVpCkFZKHO6DdnBdZCvmZu3OA+30tnA2I9qxvNBQ
Uc1KT14YnIIkghwNt2IcnxlELLScE4aUslkH3QltsPOb8JBvibf7LyTvkKYS1fQx
OgC1/rhEa3a+jJk+6LmpCTPzzurTPVhWYpkizHYPGsjX+RhNp1ARygA+HdrOTJmL
lCOj8gl4o5FX3ZTJbUegdJwn6AEGNwJgS/iKccQ3iHYBMAxc9UwbcypAMhBeSBDI
1n8Zgpd+C31nRtH/T2mDZtNg/xKocLba/3iWx9utwaVOkVMwdhEZZ5Hn8n0rJrYl
4eeG0lN2KUIn42csxWzR9C5b1s7CJh0dxJjYbSFfpYb74mLX+LX3JgiNek/ne6DN
afOOZtIL7P0pK1wzKAFXJNNokJu/oZjuLykNvM2h9rDGrR54LWTtUSkceYyGJhLG
SvN6YH7KLE9EwuqvislrJlp60puIljlb4avc5Nn6qEKEQRsNyhjIne2zeppLvhka
ew4SzY63Uxj19vSOKCHjhcn9+fhrzWe9kGCvS5OEnmBTi8uD7Xkjfa2LYAVEiV3C
I440M1wvcOt2ZIzNkBlO4cZdyU6wB1Z8VccR2Z1ZCuI5IcEh0+IIcQHAdOKFw5pU
XWwj/USMOqwz8myW4STL2YclmHZNTvAE7p9qQ5qrzEmBeEBXuZ5T2rru5oGPfG6U
gFmImxemJXR9yCwrnecbjFX7VNdzBlDpdsWgoDoUaTafcez59jf2Wb+1kQB6fcfO
Ln//xRCa7CYAVx2gidxyjrKVT8XnkSm0/OY/doLdtCt3SVtdfKagFY91LvcLRpho
f0PinOPTwd25GtNO685gqxGt7v+0t8dN8frjXpqyMUSPLtDaqUSAq+P64yM6OZEM
KrQPpJ2FI5Wf8N25I/JP+OQHv9gHhyxBGMy7G0bAQ19VPJzfIQN7OajqgYVd/h+R
J99472PPD4CUmyUSRZhKQqyrCgp2y0PMzlnZHSB+Hroo8rh3EBs4BwuZCKCbxTRl
pyOoPpEQX30pG8MRzQ/TmVxBbgjcp/s7tGWT8cHDhNYBlHw1pTtaYt9qSj1gkTRV
P4eolT4bgsXcDbIT9irwUPQsHCH0iIE+QTVQYpf7AVjXJj4KQP59CUZUI2s4uisi
Hs2DTym52dWyRyeu3izsaFRNoBg2PB4/lJPp20D03QPEShOYoTDmiq2yyuYXCY0I
dAUVBxh3lsVcTpI327RI3je2EPvkt+u/YZhpVnjhqceYEdQEzsGnCffc3LGrSw8s
QepRZqZzdA5dhmrjL9b6AHCnOopGh93tDG4lsYyQYceTGo0AtNyKpLuKGdTV7YCJ
FhGOx6erkUzAv4pzTxydlIDtuUFMeOfXYrokzWPeBFfWwXy3n11DlOmzvZnndN/B
LYKcjNpB+RUwQTTsZDekibdM6nfPJWUe03s8+WCmIgReZuTd5vD8g8OwKj4T6+Hm
NA9OCX3aEitb3YnRamr6UHiOWQZHffb2GkVdlft1PTKfP74NTw4bxX5wdDdFsYic
47Xp/QzrIeKKP68tWTaT4+SRAvNgwL4cm+zccmHkWS7zv2jTfnSBhxXj6u7FKA3i
/UwRmdLgWSULgZbDLGM34r19u4OHwnm/oXyMYssb9bHJUCX1bW+cIzAswm8hkoRL
3uyqIaxoMG3ebnfxATzEgW91lIomtZhd54VI2NJ0tr7aGepscVudZa5KqX0GsJAT
w5M5/eVzhsWNKyu9tPOgvMsL80fyVUmH8Qll2oB0zC5xIWzhXNRp3QYgWBvhpHKS
OGa3zkXfzxNNjxwhG6Sr4N3MT+2kam8R0Ou+xjBQYB4KHIki+YTHNr3ERIVjYty2
ymzVNQaV0hLENuIMlCzKqVGlC4Ppi9l5+74U0uRQRYKEZQMC97jbQ1xA0Wef82zb
yM/uDPCpRrZgGsJYIjQal/S1Uc28NaA4uyQRVJzBW65G2dcOv35nkNc4ZXGJiNR1
E9w3rIUpseSnR2ezq0cS4/8Eg+0KnwBuEZbT92Iy7ZVHJ7hB3p3IQ6qlGBo3GPoZ
z2Rgiv7bIH9sroYzBDMu0y4U4bTGRy9UuTT3t1RHJfBSs4cwSB25TBVzikbYWFcz
DYxW11+jKILvOMINysJ9+TbDFlyjfLzkHigDjq0O67fmUUelixkk+qK03PZ1ITJK
yOC7RYCYimb3dXvI6Ha5ESRdE6xo/aI9S83pv65VPwwvNWd7UFpu2bxLJ8jgoN2Q
403YvnTZMJ0Lgr8BM44Lllm52YCyQi01EocEo4XgF/eoIaH9Exflzt2rRz+IQVf1
IHALxngmCwQPiJygTV7clKl0v0t8yqRsvNwSp7S2ladGzoipYKX3Rn4mARC4TUj+
ekzz5PiMcNrtbKVs4ec/FLHOMEuWa/7WVtU5gDFH6KEeHYlfdW2U4mPGqhmY4Wq5
QaYMANJ50OrKWaJxose7nfvhIRN15GQOua9lCWxmAJ0QFljqGPwdwTnMnUHwuikr
/qE3TQJytuiSnP3bc7HpZ6wMatKyez2GujJiNiCtcGfU4FAGxzbjsUu39SylvFcA
55xOvs8PlLn58x/MYF5YvzE5TJST8fAlx4wI5o6OE+NhSjZYZJ2kz3f2ttw2l5IN
E7aCiDqn8ZQtQ81+cEZtlrLtFU4xGJE1MqNE+QbIiqshmcjqXLB/q+OroUbIxExz
upbXDfiqHGf7Y/YKQd2ytzN/ZpcmaxGA41p2/Vn3HQox7HIgsYgaSPwzZAQVRFcp
xv3sQ20kR2AKJeuLSPW2ezwmY25TltOr6IeNzqk4L8QF4jHUw2um1Oi9evl26BP8
zm0Ox/tX6Ei0CKes9AvNw87V+y1MkEKibdojE79o2nUyKYpMpCivEcrJ1565FLhq
t6bPCshV0KXLYirMYWx3cA1El5QTFQfibG7dYIFo1dHuL5cxjAtaIWLwSN8TSHh8
dfzxfOflK9J5NDIWwu0gXnObETl7WN36Vu/vId4Qbhvq+sHiB8D/lW0tJnJnP3BI
CKfamBKxhWrhs17UnAvwL97mxPBFUm2DdCaffKmw26pOLSTZ968rXjjf4Vuqyxmn
ANFjnt8r4ji4XRyx/jZXlXLKmPbLPNhC9ToEsIWA94XZdrrYIDK9Emejtw5yGfha
++3GqewqJ9AdwebUSnKobslqD2GMWR3fqDbpw2TbCcu2OwKl4T2Fn6WrXKoIxgGq
DqW5KWBdhayqDP4BMarswXlOH5oKKVesOAcsiKCHpFNUVeITlXdPXZv+dCunYyL9
TjNQEfmgoxnqMue/MafqyYchwKHVpqMShni1RluH1862bvJZewlD9zPtA150064P
sw3xwpIt36geg9hBaoXDDxOKn+LU7B3dLRww9G52zaxr8TOikdO38z4/nPSzW0vB
O+i5eOCsslkdLqwynKnY7A/q/GIVdC+bCRZS7LycaxfZWXsMLb8OC9YxNB/H6942
Ad2JiKYUeGcLUJ7vdhG+I7Mo1Dfgy7DBwFQUlyVGa+LSy1y+4zr9w+KHV9MSNt8y
PSQ1FMGbpvWNwh4GI/nk50/bk+1G3EG1Zi8o2+eHrmFixmD8KcOTxFbzFROe6K9d
n97w6KKwUz3zz9HTy3/tNVYo0Ol+oZJfUYSeI2TLpxVxHHfWbmSnNsXBZU7vvrDU
+d8AkOL44/rdHIWDy4KDQbNZvgplfcN37u4yDqs5mhi8aN3j8fFwGm0WbOQBvWTy
4WhP2AXLBNECYPZPyGgtPwKqDhNyPGYmWJ78R3f1bB32XgUQ3nrRfTRjePpHwAu7
dTaAhtgM3uOQBc93wW198RTKqaURqbGpghsGg5BG3lak78NMuA6rfAR36o2LUJqe
mI3SctRNQXuarMILYrBn2pjhIkQHmF03rbUcvj0313qGEXrUpzD7vWZQxa0n0RO3
QADwRX/HPLtXVwRiNaZcSYkFaKMwOfaV/NDHzw/nMhtaROrRYpGsbG8VPcbkeBD4
YY0H5Iij4IJ7YMSL3G4n1HI/7ssGYlYp2+KB4NyTEygevW12nEQGyL4i+Hz6gBLL
32S0XQXdLeApU84VqjRub0JSZC9eakcGS5jpLD3w2yx6emeWz/KGGADuFlCLpNgq
ZXJy1m5igm0vt2XjnFiIGsot1Gb7V56PDEnS3TRpiJPZ1eYaxo0zRIX88NegCVlw
DLZNh0t3KRR80GBekzwsQY9vR7HDkICEXJ/kUgum20MiJRBZHDhRHTLzNIZBTzdH
50RpiPzMqswYpS7FZg4/Tw3dYf6v2oZw6UQm7N1OAC2n/Vn1o06IsWrJWS3urvDO
Xjm6q4i7fYqxtj5hbFcuR9r+x4ealvxeO1u/GPR6RFCwC9hsG0LWNB4GZStWeBev
NavzCp1x3l49liGXe5ic6Qrf6bAzi2lEvwa9aaIpWptLPpDvrB1mUwRt2RlvO6AE
eeET1aNC3jN+U13lps2YSMuDITxlMV02SZ4xC4i44NyOrC+xQiulIGQgZXHIdwip
WrQUimCkI1xqea9LFY4QMgM5Ulisqgj2WmtS6uPDuIo4Ax0oqUsMdgiuSskA25if
e3r5sRgpVpdnBScqyyGFHmHkqxto0/PoX4KSLxkggHeGv4EbyhIoZGL2L6iOwrRJ
czt2FrFStOX4Izn1dQFYr9xXYzOOl6hZ410h0Gjl/if3RCWbA70Qxi202Vi20l/S
y5FE4FyNMjYAYLepQcML4Fy4jJ/1v0h650ZAT5SN/yxrmNkKYeXF+vAKXAZA4gSV
6+uCPe2q++wvK8FdQ33uiCpOTXBbkgi9jGjNx4uuZwpWDieUwaOjx5qj4fctmNtb
I+vez3tY+YCz6SMjpqD64ciS+7q3MAvpA74zWTpYcNnMtv3wIeQvdnSGVctBlWVk
SlpIQiBAdKrO+kyqkOeUiwqlpStTv7Q60WIMyB2rwa8M+VwwXVN9EcCCiRxT0mlF
dJz8RYUcy8sOhxpaeSXQJo6PurmrWTdfr4AH25GXFhnPVA2JSmfT65CohLxxz43B
qUd3mkw0wZrBQKdEwtO35i8hgtv7Z1NG58rXh6pXC5uJ1Do5uuDHcUYmc18VvrIc
S2pnBpGW0Aca3j2ixx7I26O2QMmM1wt3cEMeq69ODO/M76mFvkSBNFkNyLcyvsAL
noDVPrjleGMSFv9l1M//mXfdpuSLH28Tot6rV69Oqc0Stt5leqTOcx2Esdyu1YOE
9z54GfQwy38mthYfyortBwc2bRs5at+8vzI602nbd+De9/Mmc4hXmd8wb7BYrkX8
Xy6jmFwGiyoTnq6HMJLUaTncjY0fPd+TplKBTrc3vNEE4wupk65u6X+/dB880j9p
Hsuz1+tD767gtnsnTSUFKF11hyNpHjNAUWtUvQL3o1Ow5LbjtN5KLhnp7A+wMG0c
6MHiWr2kXeUBttURNDsckJTcoHRsPLnV6gsJOzFKHmD6VeSCzKDN7hmtMeJX2v8x
OrVJDW/Jrmd+LT3fJu1n/AxpMShZaiLDsqE7Cq5jIJ0sHIHkuwrscCYLVrZ8f3T9
2Eqaz5uSm0IQAU5DZmH2OBiYMhSmKPvrdITWld9qcR9Ra7DN+Hs2AZ8n3JAxEU3e
lrCzs97EYvNI705n/SOcbYFqo4b+p5B/8F3Q7WUbQZLRogGF9VzSczyOqRmfc89X
sJPgAdJnMAximmQ53QXF7ZEJNxeeeG9y5I9VHJwjS0srNRP56HlMcjnXOlsFl5CW
sWHs0X3WzCAHHhDGg9CNfFwQJ02eMgEzyhetEH0vpeYuRF39itQ5t2y8MwgIVaEI
uB1ThcB7H8/VRFFUmlIZdvB2xXbAibAmTNGj7Ayx1ARIi6ix5Dkyvt8J6c10kTw/
VhPenGskCcXGRouZpi8Mn95g6F0PPM/PsGiT1u2h77PCoXtQVBr8TeyaEc3fqG1m
4Rc0Xh+VdcbZpdhGQ+y/bwzu2dbs2klWOwM+AmYcgUbLs4ZXUR++RDt+sfbuHW1c
W1u2qVrO0Es4MTuhh2YkL1wJmFSiMQ8jRPbvuYkwD4o94n+a4r+NLbhgA25EX0To
c7KAqsYfkV7aV9fTnX6kjH6WcM9fwY9CEvqCyA0nXW3nzxvdu+4CLNJGV87XD2rx
TlAVgrwMWACvMEaOBy1npo0k9XfZca75/Ixkp0ZeFwOjvTj4N71DiMFVdcsFq5Qe
YmNpirLNlwzxozwA/WmWUS+a45tDDKgxweQ4eTlD7ShzCovC8aNy6mfa9+d7JTmi
LNNIoyobga/D0P00Vf5AiYVL7sHaKcS1cvdQcPsrPYxsjvR8QfU83VBBD9FMUP3u
bOtEBb/n+numNVlfe4mYulL1JMmJylmpM1iBYkhxhGn4aBqIljaqzil1GbX9HWgQ
gIGtLA1bL2IpJI3nHWahk7vZkEiBv5JT66mapvmLNH/EBGmMeKVPyvRVtwXvbF9w
i7L86caVBBEUv7uXV+BtxV06g6ANCL6oPSH7N8qqGdOJHgq78HZwYZx21cIpjHlA
fUVFwWgnP83KPdrCyEqTswrGnarRaJpD7DgH/4lKbKqbeIWFzI3vW0c68ccRR5GA
w5MLBGb5oo9M3UyOSOBLFjqawcYi8YaPah33V7udRrG67GwiBBEuLIgN21W9lnpR
qDbOoycjxpRsjMHHGVyr1hILB5ZUVQfugY/l99NVmgol+qlkLX2usVV6Xdhttr0e
4UnPTjyt7xLBIcKLG7rAMxuWR+eeKG6FGL8GotwEyyhJGcz34hDR3HZYAOzq2fOd
PYFl0lyNpjx2HOKAqLw3dGlt9r62B66ryIann7G+9eHu8NtMZFyL62MuODmmcZOw
qIZWmMxcgiWTetrvNSxzr1MHeRCha0QNvMmx1jlncxG8ajoKJi0bkQmPrFwAFHpp
Yf8auaOhkhKwpu44FT6KUZDFr5wpGI+eFw6DEd15hAoiCJhXl6aiF21dFa/ipFL5
MTXgzyC4wixTdLkv/trAX0rBNFoyrWvLbjn0vNy09i1tbdzmO7HXnyzzu9seHlf0
7nAVkWKeRFxGgYbzIhEmoj3DZXl0x7MAdoi9eldhAzthxLZD4MCpx+iW1mWuaXCV
R1tY6sE6q5e11J2+aAeuS2oMfOyn+6ehdihgweazGlZc68HWhjaDHvQDb1V+C0RO
2LyxJYOhR3WJ9Etca2cUlRLMfXI35eQb5GLgGLG4AGvlrbtXtkqYaVbtYcNcf/O3
zZxYgjwM+StUgibzm3wzk0nPqNjgdlPTJVGFXJvUtncnMZHM6yyIjE6BzrRlWLh7
8sk+6DCEF8I3EUhXK10ECoipyzrCNonX5HChOhw74byRLQRYZjQ8TFYtKGcu7AXO
HDDQGidI/aDEIjMBe3/cbHSOP66IXvHXEeMGQv0JPlFKEs4S+++cu0NOCA9xZ2qg
XL78r+mmlQr/TSUGU8jkDFxcEGf/47hXEYbtNnHOIsrSRMwR9f16584+sAUlCS3n
ZNFrWmvvKPsNuunuLwwlbysSRHRaXKMC4byPCJSYxAkPCUWzGrlLtXeRIh5xnuLI
LUhItAaF21vlqo+Et5f96ElGk6480Hptx/6DMoL1ZKZmkXNFWcnCE3A2Vr6jf6oI
5iEdA6qEI05RBszslQ3BBTPzvtpfxajpoNWr2Tev42LhrecJ2JnVd1UhWyXJZVVX
BAI2pkl8udZn+T+fdu3Dzea5yF1QLJHP2FHVmY6wMjZn80Vgl2yIRG4JUMdiqWgv
CAcf1vyPoHmsOfaBaB2y4cNGkOkWySXWCE513ZI4DHLI9VIHDFHfo3m37uSKjSLq
j2JU6Yo36Xbh+J6nCmCKiCIDy5eRD13tMaU+vBwPQOfpUunyu4Pgexq4Tc2K4j9T
VlthSgusyjcQpb7loy/8SZdQwwDP6NHBiZKsB2wykt/V+fEVQRI/yqEwmVhJJzrW
QuMf1t05OTicCTOUDVeNZ0MaBUEPpF7SQ49FJuvGbmhSrfznPvaooN9olY4MlkzQ
DQFRju7X9EsXsgdBlZQ9XZKpEpB6ON11oyzKJl/n1UH+61rqDJgynFa0d7iafA4i
y2tkw6mQBGAl5/n5avIVlAcECcRV5VxKdH9B2eC4wP4SGLs+F7b8rPT00dm9fq4/
2NM0/5wEcrjTmOYwbpSG6VuGzQygoYblw8Iubh6/qGMisFgoN9wcgX0DBcCzA6df
U4qWQX1869dJxtynJUcPLJgZ6XWV7pUMKCP2aYvy1HR3Eyxlap6AWO/T2jYEqbFT
lWHMYwVE/2hye//ElH1zQipbTI0fMxLaoV9DRr65Oo0n2Pe2//dfX2nJFpcLTiPY
Ss0LZoC9Ue2b7rANfKH5MiaJr0B4JPq7S+5/5VlBlick875ajfVFmszmPNZ1ZEnc
1ElriMs9NGHiAgBKb3dZnJNTQzR3z0ipYaZWH15o/1glRGJUX35VLM+O6VqFyu+L
3FLqCkP5wGqrkS646o4uXSqpaG7wLKcV/YN+La7Kv1Dwn0+Fe98ge7vE726+HJ/M
IEQyv0eiNzfD30394zGQURLJdRXcgVhCZ3SujX4VOO/krnRlTkNEev3dCcobbnYs
lFtYs8vDVeA/72/OtDPDKrJvTZM7l3qUUJBHxu3bjCR4lGoFzXDA1VDDmk4XqsXU
ssrlrRVZgh38ZLEuUuJf2pv/NTUM+R02wsh444LBYQ22jgR9jiJZi4fAB9rSi67i
ocHnbWw4IE7h07+4r4LCIIwVsaniumKHmh2GNxzYzPTOd2VuBrkE3eh3mHgSJgBu
RCG6hFxcY1bPYyq5fTowPuZCG0bHI8N5On4KfbcnKU9H+RvfVdg9vvby9xjG1Vz2
cAG5KkEaSlu2C/C7WvRo83CKvNfpbTZ4gaWZNak5QQTMIO94mB5GNVBljDHEZJc6
k288PitAmK41ndjLHc2Rtp/pXb+K/gXEbmuyhWEE9PlJWrFzHqdebwTpal4dfwzB
yVBRVVirg3WpqCYu9l2llwBHrzLWcqNPoROVDMpyebrAPjr2l4njwIVxgJ3HSOBx
MLRHElj36IParVSnXA4qmARQVe0ccu1j2sspFfEM9l9vt2YeaDm39TvCxzWkYjcX
3VF9VwdCl2dwhnLqtJLha9F15wdPNIwDKZ+/MeKNCj7hdybIO7pVmgDyAmZ0nCca
z3bmxJPP20kM3moZ8kU86Ris0vu5NQMn0I7JB6BO6C+cNWzN4G6g4KuZ9rQLTBEA
yLsiED7GX00raL8V3NXRY7ZfXFAWt81qqy4ZT/fcCBK7SX2sZk5rN75G55dittuX
TboIQwpiwHu5TjjHf4EPRbiO0ovogBjeXB/Pe1+eQw6pm3Lo1rCW/wwnAvmcJ92w
sVJAle3wON+PjBTipwEUveqinG08lM2mgS1YBwdsNH3jTMDBrAlqMysWqlIvi5My
cuvP2Vty9YELGQtP366N/lT1KQf6PdNRJI0kG/vM16kReR7Z07WNQJRKR8tO0DP4
80ajfs8msQIeH7OLds7N0yVygiEauJGeYIaZeOSA/e0oqwriX3ZOHJ5MDlhYnkz2
zj+eD5tf6MTjy6eInaH4mLHEd9k5VzGvQJh/mupOSgliebjUFHg46rigJKPG6m+5
a0kqKPexSH/MypkfZ8HxoP2y4VoxbVstBT2XkdYZ0FR1dXeZNWOLXatHECgHu8Cm
grStvqRNuSClqVaeilKaY6fWdtpvscHMTUKZyNmh8WyXcqrXynWcexC9jcEVb47H
1csfZtqBKpHcJ0o+8ITRkeGJC+XbUqQ7rqseZqz55fVOFiLrxC4S1eLdV7PVW+wE
OG0XGNJB9MRNQtDWgc+rdxJpMaM4ijRi4xgXuTVUd6wnmyYLSRFOyX26FXdFQLK4
N8AHDg9WIggioMx+7756/ZKRzSST99lGJMyDAmB22/ymOtuUZpH6bjW4/Gus51KJ
qbQBtaVH9FA8psTjwWdG53j7eeSzAgLc0j/qG9nHNEPvpx4Gq3ln/kT2/CUyFaBs
FWhoeD27sVSGc3l4IbpsT0E/GAHcV0Sji7SqpjePrk8o2DfmWM2PeXigFCZGipPH
xqBR/g8J4kV8TKsHA2soKWPXnbJB+QUJtWf43eyUUFs0fVqVxPOEjWMrCeECbFQs
Nk/+PvTAEg6klLoatdCSY6z0mK8BulVWTNmNxi+fKyvOApG0CUYTtcOqHfq7HdvI
RNDCTOeMotnf2INW3WKPTHjSz2oOwvwflbuoO11GVvWMxbRvCNkBFNsxh2Jh4CRe
Xoxm9CD8XcB0dr3BWhrLLWsHciK+byxMzVV9pZlo+EdajydnaffEnsRCLta2JdhI
qtVBwu1SkHqBEnuEK+KLDnEjqIrLk4EHSsJQPJXXMYFNv93xtX0XlkxNi+G2szrs
0AfxpbMw9qPnQ1B5GAYG0YDGGMcI7ak6o0kdFlWl/TwDnhfTq+oZDIk9FJYbgNDT
38Fe9f77qznvDrQg46h/JXFE0KGa5tI4be8MvzoNJOw3ZyLqVI7+dgiLolfJV/vd
xjxzkMgRAkaNUT6ABAkI25x1zUVID19UbxmD7MWkOZeGPClWLx2UwO7brq/EG6J7
wpYlClCYDEMUjb+Yxkloab3Daz6tKX8OmESQCPOMuI2b5rZGPIoiUPLwrEG8LB42
qd/gEKynZlJJkAVQ5yDNVOc3eB04zqpkNt4HqjProDFwACiG4gfjxF8D4mX8Ruo7
7Y3cuDLM3GU5fGDcWFYKab3f5q7/kTXK1RFbJ4weCZQyVituz2tbn3ePvrHmgpUH
r0OnnEYuXuzZoSpYPY8gLWtSQyT94JQx4a9UOa0espwIVnyxiPlVhky5kW+basXN
dOrjozeJSDCUucmue33PG9gfOOfsd7Xir7bDpFK4ZQ9zJYHlIS6+UM3AVcXH3J/3
H7NstuL0AUDcYFYOPj64YfWr0Yldyhn8uvf6+kMVStPDOIhCdBTuf614S0mwz/Wa
wGvv2PHV3joU8Fe61By3jtF8+VZi8ZdnR++Unzu2E5E0nJlAynzkEosDdfjUB6dG
8btpTJt0T9dkWQZ+ctEtNpQEk4B61sFnFQQ7kxDUW9Zk+tnewMDqGu9KQLYNQmoA
t7se5F3X8rOJlu+uIeSZMTJjrMC6y+Z+2/3uSdgE2M8c9VRUhLkfoZCm3pL+NLkP
GLePLpYCw1xXu8ix1AGcM4oeXyHkYf4OUoVOd3ILQGHpnJO5DPMY9cRv2/V6wVfx
kC6hrAR0GMdqquE6vfx8gn+rpEEsbCQm3Is+p/0TPhaMH2R0idjpcP8FNl5gfnHs
PH6YfVO6JXUGD2jvC6IHRdwgj7cKCvFRvkyucpYgm2EMIn2obpm7o01Haj1PGoK5
aze1dN+8eI/dytZ+4apTQkeAe2gJ54abHySqehprVeG9drk2LDR0Hlh+2ZZUFyKc
k5pu4hwlGKA1E9eaZEI1HxWe2btOP5zG+n6QbIoWEvkGOZ8MWh0oViPm9V8yFbLk
f84LfKJdkAHTJXx7mlqi7w7qr8HuyuOb88oT2xehWzjPQc+nQMXmZ9Be6BBdtdUJ
jI2+x45d9i0lnoVhEhhrOh3D+nObbrEkab2urmL/uR7htbahzemGhfxJQJdWBHr2
uOpmAka+884H/MiHa3iiLOGihV55vOW7sN538t7JlgvOz15VsHG/Il2sBiN1pj1W
ZV3+Ls75C4eOB60qEtrV4vg4qVHBsX7WkvNp+xYwIKE8Yu+OyC05T5kIIZnhmTHF
hJtYIsiXxLUHcO2AXFB7dnf61o9W0BUufVJv1SRwBWjqJJLnTc3C5qMJ4AEjbhZ+
O3PST1j9GHPgERg8SMC431RIeviFbKEK/9wVqwviIKh1+qzkO/nuP3sLn0UCLT5I
yMK32ZoMIyHPaeP2H8AoGBbby7U1kQVmhfF7q4RpvEuU+BU2LS4ylAQXq7BaF9Mh
8ZC8qxtlwVJsaL0JXMVBMSyZotDud5D/mstpMWY5La5xENAXA/BWyLG296Qq2CtJ
UbghgGXbE9bIokVBJ3hN2ddk/eYSU1FFXirudAa3SfSqUzqF2tgVv/4dw45to8iN
eVFtP5PkU6wXgW3UkPQEUKfPWOnOOczWKVODd7dBg1xKudIuTeN6JWTi91ZkkIZU
bFZ9fIK7NH3lYqoMnW+BMvsnvvBxGiSY1TieqFKmD2tOhCZeh541sSBVKGAdPoPe
wCCr0APnzkXS1rIumveEZgqCi4pcjNv987Dz6XFrR6s5K71VBQ/seyFOnQKL0FZT
yDO6hfR1JbQKRmf5cvx6zRXHPr+peSEBWaOStgtbEA6TXBpzzGT3GfjO5m12/YE/
gKTSwNpOTs/5rBT6iWuR+8XU7j3Mee6vSBja3bDAWyVBOkkJaAq3e9kSofd3DQx4
c94AoqxUqVZouVHb5Cm+eHSLDac98OAoaL3VRSUtMCtCFTk9FWAIBytVa8wsSS34
ibvgNJVo+cwCMrbBLRkvn5u+bTtK3m6BPN77ukp7Ze1o/h6fPX17M8QB95R6gs9K
nfpVme8aLe2P9mZGud2z4Wy9jpcv64IThYJ2Ayzu5mMlkgs47ebEpwGeT7t9e0tH
9gZ9A5cDfXqJrJIi3XgM/zNaz8klmE3OgqoboQq3F2BfSS5kCSluocNKadIoLjhk
G8PFvi1GEw+UpIMEyCXMpBi7UBQTt6sxBvh1RCG9xOvhiH5+g6YrHOX49V5AM4SJ
PetnoBZxurRftVO8niFYdz8wK2j6uow/5ngmHH8STHOnP26NeCFWvHXwDnqNCrr2
r+9IxZqR6nmdrO6E5xFHNjQVXrQs1NT0ViLhfBdkd63mYvgc57VaYk9hqY1rNrMZ
HUGNW/1AqNuvyYxRIWdkZKSwg1GV8fQNqnh8sa3N4RtcdUgFSWUdnNnccjogZ6f7
IqzWn472y7mflkF+8dzj3bfgSbnidv9y1pbR/QM2mFeEfZGtGUkLOp1Jho5EJVN8
/kb87nu7oIQxnjkmnJnrE1ZyAKIFVj/ZYVU1L1PFyPm2zBzT/iQNpkw1uSI7eIsh
C3o7EDS0xbuGD/sPuY+upuYRkR8yVfeHOgEQ/CNl9tVqwy3EhVXABlX0y3EJYGH4
wtj5fnobzhQlHqo+E1uL6BIFXQn/nI5EAYP2oPZlbN5TUVmPu1zHAGyZJ9lkY5Mn
bGrDc/2gb8suwZH/VryP/zNneNnm9sNmHL0kTSV4xU+D5vVx4xEsS8QOQGvGTkNt
qC7gdHxdDgE8GNM23mEN9nEtapcAXkNlsGs31jBKhTqa/JfJzR7yR0VGoZG72wkk
lW7s1DksXbWZj5eGdQZlyFB4bdAsbbUsJMhiaKI6DEFIKX/32UcOTQ19UI8m0ew8
5ZZzDRFsCT2FA6XQEmOj1U4Q5q5BbIbis4JHdj5sqDXTM4xzUaO0w+KbVWMZrHoq
nryOk3A1Fr+NK/VNtSOcgfyLw6SNmjvCTx3BlcsyGFugHze5YHE6IVAE5gUNVJCS
IavSV7c3y+pdRcblrGVT04ydQRYjrTX64xS9CGhUqu9J6dcVIx5nhJQ9pwXPfrd2
YKYt+NmDAHws7z+je3TkMwfzUJKuh9MZwPfIhG2QVsvIwOzvQQAyl/sg8ZhE46nd
VBNY65q+lgAMPnIsEfTwijSzBjPKLwL/2W7gwUi35kfyijG+MDe5NNG7LAcD5Z80
o+PYc57bYYfLngb25MIPS/+htKSe8UP/4EuBhav8LOYY5qFJfutX3h82ot0FHm/E
RMPN5COvJ0+L8otIuVwO+nQIsmflgZCezKRHNYk0JhiIaFpIYTVt+dt1VhycnWLV
SHY4f5J86niVt2of//eoEw0mzzPhvpdP0HjSdGSlKWFuUAolyBK3vaj4ULjEF++X
dquwHwWbFwbiWkNiyL0O66okMzXM+gJuIcp6jMfGjiJ8HNPjdyOeMJ9bqIO+ut4t
3FXfcqv0lKJHzHYZoop/zSh0PqduWmV+Q0cGTovWIyPxtOoulOgMF0JFN0h8FsHO
KjZ6rNEBGaeCq9KHAVzXCv1A537zfd1t5PzWxpk6KgqgVpVII6S+IUUuYwsSKBBx
ef+nOIHi0tsJYL0iE8HlzyEcjyFmxKU05DaDYF7pkgUMXn50H0BdjDLsjkw4avXb
ImT+aMcXgtuYaayLF/7FnvhqfdoLx/34rnHElblTIS4p44lm48O1jZJF4ec3IZ+y
6mcH34WGa9BoaSls3l3LrarZ8zxNpwJMNS96pr/516U0IwAqpdM0HRWzi+MotvEU
i2TvgnjNjWlWhnulUhqDEwy38TWr4mlAlY7KPdsvwkXThhkyrbYabddnszaysnW3
ZlIiektKy+Es1s8D9MOaAalhlXwrwf0OeOvAgcm8REzf+85JJ40qbudjf7Dsz6Fv
UAn93nV3FgXzn4DpyPm/+A5koWgzuKDerBiiubC68WBuaOsKeaTNMxNaqOGnLyAU
hSFruThK3HPwB0QNGJeTVqinGvDDbVE2g7Xo38Tik/L6Wh9xxFEwJ99Faqwhazku
buhz12j/v4F/Fq60S/QcHWF/kRa/L5yJ8QGKTKkg/t1QXF2EQrx1ygFoGuXXE6dQ
N3snaEbgLXcxpDh2WuN9fPjHW/SV9e03K0YT3c0NTu/cLXTV9sgQSOJE722BE2Tn
jxsfUN86w0ehapovjCcIrXwwWxR+nl9jkK1eqCqdlY9WeJyPAswFCZpMQRRM9C2V
QW24qmKA9KCQOX/qMEAcg29EZ/cpHM2ZLgbSwHMOV8RR0XFm8p/Al8HVeE4hVPct
erNMqbGeUSEOUhfxRBzn62vVX6Myeo4U9AUu6IaDIP4AgRm58K3cuW7oXgGQQcfF
cJzK7N1vCOoHQfCV4w5tdcvsMfj5ptpJNTQUL3XvOPB0j4xqCuxtPLcQvTNmBoRS
Z8vdt+B4IMZcArTrbEBc1mIccCqCfKWd+z6L22UF/JvM/f4BT/bdWL2f9OqTswVa
oWCsSLTjpMoKXHgOVaFpcaU+PD0tk8emS4g0UP0yPGUFbXEBkqRx8MNqCv9jIBb3
gDd5R+pl+sulZdUn5xKKQMCxd929ne9TT4K0hJ9gsbkg+ij/Tk3flZHVOR02LLFT
zhTlHrcnlCWhTP1mAlYgK9M6z1lt1njxGv05TwF5Xd2C8eQvn3Kbj/BTsHNmxUei
zLb/BdKGvr+s6fVGP9Ma4UjFh2g+YBZCrKI+Sl79LFWGUUIKBM8iO9iMLTfwPSra
zYzgOJwxiFijXRHC4oNiRuovqNwJ0g2Q3vrl5Dconud3QeSC/iHT4kxfYKcfAwYm
xNQBFnN5tl2P4Hz9L5x+RpNUJab3bUsK3EhMUJA6b2MmrLgjR0gwQ7WeoVOZ8sFL
F5+QWzsAzYBiWiTELKeoIpQ557MgDPyJGzI2dLuon/T7PqN7Yz01mN85mfrOacE1
UtdqSh+Fz6Ekx8f9S4eGSWGr+kBq2WDZp6KXjE4k5/uGxV+R60LYiR0FZDhiy2JT
JYYIqZFQvjB/8sAm3zM8cpGfTmouOQYTHkcqA6BxNTtI0KpFGZTtXn6Ro4pz7rfk
kRwaMkh9pUEFtJZyAge0RDjjQaKbB092x80FT3/onQMhwaeIhDyOhm2kUxFMvl7Z
RZCMbSwvX0uofx1uPWQ15+OO76yJEQ17O+7O0GTAfTXYq7Y4h+l/nFijqrdQxAmk
C/WlV7+uP73zJgUcQVdmSe2T/wMpsPgz++rdTRYnNelS2PhyxFl1Kwib1WmzDaWB
27n3DKCpPdu7UriSJrR5ddKf0NsarFk9AcfASf5NPIORPtU7oVK21xnirXtDz+Wc
Hf7OPMDodNHvLE1xq1rEIfC8NZ9Avw221Pjg66z2OUG+FyV90huLg/1tWL+0elUE
lBjDuKwOvRdIuKmCLNdhQjCgEJg91t3SDWIt9HDFNBf68/MbMMxJriCEUIeTujxK
jpBJioiYWrtv+B4LskXFNm0NXw3tC8/TdbRVAkqcebzqgffgAlHzSfheOND8ZMj6
jb/m0nIhDgzAwTpi+DAEzLCHTsMLWdm7fhi6QnWAGGcePz+74kcSPra8Cl9pS58y
itMTs8pYJWrFK4Dw5wUNrnE0lHYAv/M0SbtXU2FnQKKmpbaY2X7YkkSNUCD1U2Uw
Py4JpBjv/JzdRIPJwleyM3WamrTjKdfWd6fgF58I+NxsfP7YRlsGfdRoQLqxmwNa
MINw3IsQHta1XAXkBFUZovUMi7rsxy+YM8pfZ9DGIlTU4eaFcEctKoa6uXp1Diaz
Z4iE+SEyWHNNikdheoIsYVVlFCdckl6YsJCtcDzIQ5DSMiHswk1YrpR+gPwFCyyJ
1uZg3JMQWGvVEAI5I472rD3ZXqtM0hgttMHolDEh3sABHVCkW51eiomTSITOQnA6
tPk8m0SrldneI/fEjuyF4DmvKbFppOybyCMdfjV078wEyE/rKnk9N6hSUgcTruGq
4ArjclMSO1XrX/n6/y6K9mu/cl7fbl2STgVIlxBMUk/xLpnVChgPavK4+ISSBFKM
HlNxgZa5AtZag0URco6qstFsztxR9tYUb9j4FEi7Y8zKOPTaji5TkTiXHHkDxOit
lxuYwS6S0KZedTPqLLJm8FrrkjEReBzTQh9Jmi2jzghXAoG3QEB3bV5Q99uFoIyl
B54ha5gXVhks388fl9M9Zr/03H0aQSnRxQhql3z5GHZ5q+pdxc9wSCq7QqglKQ+p
bOYfqCY2yAEASQnGk4z6CVfDpyzXiyMW3h4+2dXXga3+bAX1euKJvCM7If/osaf6
cbk99UJgyqMVR4jsnis/qH8JeifMR7nLQBU3eQ5cl4ZmSBz9nPzCx4jwyJHSPDcT
sFeU+xCi9WcUIBkHOIXmFJzgL+4GiSMWboB3wBQfqFolgsVh/AFNjWQO2inhCcWE
PsI0dsRlcEOnS4TvEIAeWGknqB9a2fp73kOZ2JJ4uWPxEYWdvAKgh4z2QiOvTmQW
uVauy/saTkFo1RfVfueZ6z4kxR975soeaIHeCKX2IWuZGXENmYB4ikNeM7mfJAVm
b+8wAbbc/SJpGXG5NtdpmaFbTV/TkPJMCw8PmD/ggmwltC25HUlvHu/TLtgTidbF
hmC+DuSSTYHv226qkG9QbdQbvHkKsv+0EP8A0pi/dgzqsimRrwa6zN7ccVU9Q0nC
mOlg5M7jh+kLF9pByMENnukl9zM+NuVD2QO/EEMoe92iVY73pHKbij140pbhQOQl
UXyppREDmPFd48b9MjHJmNVG55ecMDxnwtzt8NUFnp/J/rIzMeKyYxxTnKu1gI/C
c1MFsDdz10wH1PgXhBHNuSyOFBN1uM4SgQuE3hwAucbpEfQMGcGuXzU1uhKYWQGc
ZG7H3MleCK40VkIw97aqwZfQfBF91ne6Jo9XzNK9Ed8TklqpT75JTcHrGTv+Vk3G
nIEq0PoLpOV670TjjF3EzFWnidOCrcZzrMXkeo+nC8M959S0/kqS7qOo+3+9xBQc
3oN6IK3jQ6msZYvboAIqS3kcGdTDZyEwSEB40V5pfNuUyJIgq8KonopQf7mp/tPm
bsS5XEFjyNyHNBvncQ1iMJwfIUemKj1px7i8SNWjw5xB0aoiYQz94E4yzPm0MuQa
iNHAq2tTh4s908bolKfslklvJExjOYW5PPtsAziGMfmCeD2BZrKeMoPShXwy/oLc
7c4nK+1oEDTpbQcwa0fxRqR8DuDfxGMWkieo6LB0ssCQH/6YmTY5gbXblhgcoLrL
6XJtHBmRqgKoWvIG88Hg1W6mLfO8jFon9cK7WUN84hAtdahShBLFx+8Dls9s3Run
BjowoQXLnMS5GnpPUx6IA6ZNZLadNBWsKkhLzWq61lGh6dTcnTKbYURla5GZrOyp
+YXyDKvNG8P7iAGmxl3Wre0/Lu624eumc1h16UoI7fGeG+auk0lZh3SQ5FXi2NNX
9Rbt2Bu9B9EeGMerAIF1szlTY4aQMjv9beWpg+xi2VJ7qeU2uPRYIYSBfmbOh9uJ
1OgytIoiSD/TzViJX7rxGsINn2P9a3Q+Z66wZ1Sjb8squvCunCaZ4Zv3n8epe8t7
SdAmkRAE3o8Gqe0+lmaPL33fmewr+Ro8RMQefwU6z8Sxx71htfp4HvGrV6bWCOJ+
Y64n0roAE5CqKt79KXVGQu5z1XhGXwdcKVb1o4V4PfLhhBFLsAdqkfsjbBS4ytmb
213pj6B+nSRl4yvWZ4XWnwsxTXW0B/9RhbUz2ZpwLRlCj/mtEvaEdRodmw4nAKpa
9r+0X7Ozny8LnDJKvl0Bo37fBEJp6ed2Js0CypIx8sX7JKmfGuF++KIjtbKYr438
kdt0IzT41myw8PNHiZF91W6jJzLkT41otXexNSCofStRBA97a9//Bja6Bdk1wcWU
U9l0cyQpNznWQH9WIw724EsGFr7S0eLFl/9dIwgshUOgtWluNdGIT8mjWGwhgEvG
ISdFhBj+n9LgfQcadLQJnR0XvHH8SGLxE0XsZ9wo3nTSTQ0dzGZ+um4NGM+wFPFS
e6rw+dPlJZ5USYrOt8curaMFPBrWYRxd1v/FkmcjSx+4j+HdONuWqqUq/bULivAn
51phmlabAqGvurs9QF3xhzX8TUO6KDLniNjLnLJD2+PeRTK9Qh3C61iI2x1VNIBn
HrdBynR9Fd6A32AJ/g0PK9RR//YgEeOy7qiG5C6X2C1f4mMul7m6py+oRaeJ9mYf
p5MVIWre3kJNqtdvuP8ybxM9QrK+XLytbFZ9qBcJUTNqVYQIEeg3Vxhr2Zxl4ezV
qt9G1HfemNp0WDhhCgpxMJtwTJz1BCha3UAPAN8dStyZOdE05SKHnvMN21ttQ4LO
DQv5XIyC5RSHzJBa5X1Ivh+jrMspVmF2Oxwvfsl5vs7vuwvQ2mAoyDgBOyJ46baz
J7ps25ftMAuFbaRqWrDuizvzuDyw6GfqK8eUZjsZH88uWCt1Zy9bKmfIjDcAz9dP
45XcQbUizhxjG/EaxtXe4dBtkRMCDCoQxFrRgRnIC9IoBhkr9VEPN3UCe0MMMnWu
6EHFDrlUG/HxdHsdHS6BAPx1xLnVhHd/iPW9L8lmaTCTnyu+adLRXAxwTGN6k75g
Q8qgVtknjFitKSerqD+oPZc4swE6EeRMj9FBtzemsbJPl5qHKHcR47RxM4isi1S7
oc9sJ5XSIAoTGCpOzD693M3Ow6KODCuubDR9rLpMZA8GMJ5WQ/7j9xdlOIV2a+9q
wBKt/8VGoasDkwGRxNllPwmzNqskAxq0jq/40A7RuH5HbYuN3YhacXQJOzBkvDZl
5Wmx0YwmC4gzx16Y+DeLcVybhIyHYaiyIMHF+BS3IUq0U0g0FRQ8XJRiXYkfY3GP
ecMb79JR+svbZtSawGFke4aJnao7z9XUmjMjdnKANhDJ1V2/cDskAXG9El4SIqzk
/Z7qtsIQ01WOTkD47xO5XWZY9NCgORVQBBUt3y8G3Oajv3Jc4HBUFQHMrxyFQWr1
Ny7nESO0w1gxU9Ed+5y2C6h1OVH6YzbUBsf7yqdDqgkAJGO2zidlLz4YC+H4eRKW
++VHgq0qSpP8oAvArA9NNCJLse/oi/kliMOC+57KevttKMzA/QZ1lpC+3AsTycGz
Gttkd/Ot1Xx04H8MEIHAP3SWYm30q8dAjwDhCWHf70E8fQCgCoPumyzS/quw6KqJ
dmDbRQV/LX7A8jZHhs43gEEuYWMSgTdOSZdCYQQb6/iRbqetsb3YcDcdcY9LRjpN
ArAxWOwO1pbQo4f/R9WaW0xhULIKRUi0QOgVC1JVCdlb9+gcWJm4hV4v5qyd906w
ckDtIsYPIYiZGapVPhk1oOyi/QfIatRr1uhUkbe9MJKFOPol88Lus1EvsHiWQPma
AjO3+sxa02znEKIAHXiJkrsXH2U2/QxnfVwtA1+Ag/+4YuTQPbnun4PwSTdSpFxf
e0mseZpdhx/6p6CD4QLKdefDhr0Lz+ASJ1qWuOLqS2I4YWHsGijYTbTJ0k07PwhY
c1qTYjeEq7xWHwU4pzkFEvGqUm6wH5F3Nii59E7aniE3t82yUCe28xlpIrK0z4aX
1RsvkTNl0bd13lxtIzsNs/WmyuBeDyfpYZBA4T3ZILtb04T+x7H5r4Nnxp0GSFex
Y/WeAnc6rN9nR+MMrtVN31fwUS0dh9VMeeF4hgZIzfS3twnXnlaVaWaUysOEwZG6
+0hiKvWzi+9LhWgFIrOarRmBzi4uH+huY5CwVJSpe219inF1zd0daqtuib5TJNDc
oFTeGMV3aBK+OInuXZLnrQQCwTPRubUchC2fC0krz4BMrUg2qZ7LENy3TZDyPnfN
HcfGkcYKfrEEzVDvnORsysuPiZrL2KjRc7foED4ZQZx6uAPE69+gWOizVCmB6rPm
Bat37iTdvvF9V2z3WOGALqIaTiEna5au5r2fDuYjuT35RVO08zS3zhTajLANIGjw
bolLki6rymsYlhME+IkKUs0YECH7UQNfgQTQAyA75VtEU970kT7iZFaxtotD0BKq
6wsv1HzZis2ldbu3RnWz0kznJjCnk8rxsV7rABdHyLvGC+5p+fMw5J8AKw3UyHD+
f7AoS8ruE/KqQ6iRP3F/+xEfK2LGH4tNZK3AlHDbxHrakyNxL6IeAlhtSdRwSC32
HqQ1PrSRGfxSxvry5ZBIhV88Uz/rQKHpK7FZaoLDvxfS3BOILXMEf1uGfxWblcKt
cfm5thp9Ysaf8k3jHeG7J5KjCNV8xd7cT/mrhAz511hdfs9c8RA0y9pN532g5rmt
pKD+3d9uZeSnvJGqtykZkhEnQqszO150SxIa9SkreRzCRjDYJ5PaCflyl2M91r8V
YmhUKnX/gZHS6xcFusVju3iyRlDnw4F/o2ipzEDF0sN0+tuLfQVgeWJwRD2WdlkZ
LwK13Hpt7f1Js8kwmuJYH/7lQQMEjYcWn34Y7reLVYUuDLFreY4Mixf09kkRFTmX
PXOKtteol84W3Z0nH16X257zUXgWiVmPwngcLJ2+BOj5B1SR+vLnZMDGeg/SB3sB
FqMNUO1oBJ/IXqjgC5M8V7F9CQZjTWpZIBJM1uPct/2gFZZdLiZH4lYfrebhLP3u
rzs84pYJE5/s474vhq3wCEKe7e69/ehDTyz1gQ5rAFXyPxOXN16BtlfQ+BcnM6BV
pf0o0ji3iLxgm9fdAyubASitc1kucd/hYwhP3XDsnZA/nWpCr6p9aY/uBBQVg0zw
kZc9svXxflSwhLxLrHOq0TFIE28RYX83jOjac/qW2IwSFVm5KJCJ7gn0FBqSs4sJ
6ykhWPCjh7zFjGJLzpVKpS/MkqIMH23i94rQuBcwxkD/LGUEWlE4AOUfZB7diBGE
/GLqEA0IyvwGe4XkupPkBGN5+wHKMleYEWuIOUTkcAc5X0L+sbZ2E/1Fn+bX0TTA
w0iHQWhDNNF0kzeH1yb5QBDEX3bdj+XAS2HlHFsavOmjqruyF0IKPV5e4Tafm3PG
lOYVcjEqM4D6MQLbKlhBXFcMB2B1BNnZJbl1coVMsNZ4vSMDzoU8CwmuDA5F1Udx
RC9P/i5XyCeNzHQm4+aFnlbP4KF0T1L8jrAEuyEa5XD9kBO+9iyFnAH+i4WkbRld
UNZbfyLNZTCPoNxTz7t35jVEu4/xD+tFxUJ87B3AW7OaFUuk3vlxVMmrjEk1ztEM
p2XVbg+NEPp4lvsmlkuU2WsRBhYnbVNVZPVxI8pf8/cZJ9Tj8X6sOGFiLIQS+/9E
2vtJcU1IpmBmZ6xO6xocaiIq+EZhSmq/ehfYn+iaicEJUasSaquElsDDAmNwKJaJ
YpfBJliRlkgvG+XdJ8qvpaZPfD1KhGYQNflq8S+ENqaB9JuN7NXUa7P063SDwSm+
fgTQQLIgwnc1AhsleOkkUHNCQlDOOTpM4hQNMLiB6BfjNANnSWkCWxXJqUI2x8gA
mzWG3ccvi7HdrLbKmXsyqhAfs6lR+NciFdQ2hv0+Dd1VYUKM2fFAdDfsRHplBR4J
wz10BlqxBgbTPdqEYPKd1K32YibhnSvs8jDHVI6vgfH70t+0WCdJ0KQlkQE/M/xf
vqbYJDsaOGQZlh0OYUhwt/u0Q0g2KvyLRFDxFV7jkGgvQeYF3BB8czbuveYeyZ6h
5sNaonM1bTLmZAr1KnkIDl4MoOnq0pEU8iMcK4x6dzaOZJYG9zTkqIkBYjl57Iu7
XMqkbiqkXF8s161GlgVU5nyuC8V++JYshDFabA6iYbEZf/N8pMQl1HR0eV+BR7OV
kuLHnQdYZEdJkdgJy5m6wjY8KNIOuLxNE0T5N54yVY8JDtcK+tYSTkGqQlpFR1nA
8SEOJbPshM5l9ILJlDvLNfs/TZlJsamUR7KqSiXezjr1LvI8IzE3r7xGX7ZuUZiU
QfvblBiCseNi8oakpJH2Jn/9giUp6HUzS8HTvoL6H2xFn8YN1yvgVNTDIQ1JgXjf
ht3IefXHLxAlKj335BySKh7BHpNgA2B5R7lUs7mSG2kceiOsaGFOR4k5OLDqRm5F
Wi5maie83lHfnf4jjxZKmVWasVmuNFbdB7BfAqlAI/0gJQlW1gv7y22j3IjNsnXe
kll9BWCzE/YjqYc13N8UtaIAyJTOKFqmX2fkzkMvuxWSutL2794qTAyKRCZRRU2v
ZmtkO83nE2+dcPfPD8qktDVMCL2RrdDCOP5VkE/+bLNcnvEOctRnEjqaTUy6M6YZ
W/u+ZqbfSzq9vtO6byO7uh+wWDinA9dqbgPXJJsDEu/6XZHpEh4/uK9LwB9dH+La
NSbCnizx6tKgd5IcHQ9FbtAHMloYgHwhYPIFqKvpgU9+0+kQO3NMIWr6L/6nTjz4
htOeRpzVDmsb2qs7bpr/DUY4ShiQxszGy1qCufHO6hH0UxAbXnRWHnNEafvWpEnZ
7YYHLE94SHiA5RuVvLjuiGlKyGr/68Igj1ZMVw81rQ5mXQpByV8YHZqe8FH3IU+1
c0xY1R8M88r8ONvAZ1Ob5atuUJ6o01EDWi41+xh/9hR4kzF3b8un8UDbcCmGQw6q
p9hiFI9PecYn03QMHQs0zyiwEw9K+x3e7liuVebZQhVjs00qV2K9wFFGWbHA4hZB
95CCJZ+V5ftR4N/hnIfk5E5r2MtJhN/SlzHAeXFnQOHBvlFhF3+vlKxCkZ5TmX/0
GcdPpvafhmrT34jvU0e/RhM7byKZKOupKa5tW3/YY3k083GGxJg+SAewkrVbxlHI
4qgWBRP3C6M12pDgxhb9DU39f1wAXG+yfgfvYLWEluCz+VvUXtYB+uLkiCM54czR
njH12rQIebj99DEQqXtI/3aM54X+Smpy/9YX50WYcj5rtOsGluNba+9tMwaTXnrw
GNZM79kaMdf2pE50j07hdNtUn1qIzmo8+OwRVuaLAC67ew34kh3QfTR94FqQmFZZ
+os9NB0FUdktuLEK0rp3tfaH75k0Ww8PrtGNIuymwPIib0faFsebQMZnWi+/+Cxk
Lu3B7qB9L6TUN5ikXtoUdbWTY13ix9T84qu9p08m23RB2WDFmDnJL00eBXL4GNS/
ogA4tvh7SlzbxFnEphNFOPpArkCwrduH4HAlUwiUCX3oh8SCZN+AYp4jsdYzQkSz
/nXad8xPQ/5pMUwDZMQMarUMDab3GcelD1tKA3Di0L1yBHv9p87aqqaFHzL9D0Uw
i3jp+59iVaQIe/pR1SLfBFOOocpkC6Z0mM3L4soAAdmP2HEzggACIEwzHARRW7jl
VJ/vCRcbRs9nE43YSOjnv1GOVFqd3JHjhdoJYVWpz1EdRUdnfZvPzX4qzGI/I8Vb
9g0Sqx5M2v2eGAYL22/4NpqhRzXgPFeDdkMLhxEeVr4ItXy/uFVV72vT1R0YAXbn
jy7pTFsRcgZsZNPAJ3LEDyT6YXGlZNZ6SGiMETzbWGo+t1wryWs6rh3rBu24Zcri
qgf1PnRLHVW/RGG8g237uvrp2A5fnsEKHNw4I0vW8KPaJmZyeE7KDNiNv2qRu8GB
+gEjWFbvjoEfAcgr1guWcwrxrFoh+xD58rmAvwdLFMBdE2aXfaZDq0yjGnW3g5CN
hkmT0XU5p1LQhhQGIrEeLW+TZf0yUD/EvCtMsrl1WAkQjUCEDTEQEJurgjwvnAH8
aqhj3q4dqq8vqdcjcZmRrpaRAN7p5ky9SHwDr2jd5QYl7ArZkEMlzHJT1JemVQgS
BknQeRUcxqEL36XvXoBVdQ2BFcjo8IZX/wvfuZEuesQ6ffjadkzvfHXVhpCmhjTY
4QZ/5Ah/48kymD1EFd80J+i15iEZH93cC7gyuOGHfDqdJq3HIEgb+JbI/q+e6mc+
jGcRZvcob5GgkfEjLEk8nfxn5JCPoyqMEuSP2d3eM76Ha48/jQo40eNKlTQtj0GU
E8us1VBOxiQ9Lnt+AYi6Xt6A+r8xXNuVKAaoUbnHjYxYyDpmAHRIxALlRP3Y7P/F
ex4Z+ObzCSi41VqgLAo6AwkoA3JWO9LrXfQvtx4dgkWvoZ6q8i6p3oT7wbI55g3/
E4l3ESOc/bBtAJgSOBb64c0bX5WVYsBkjCN5wtoOuPLBLiq//dqoj1vIa+OXEOzO
b++T8/bxsVdxuCK5Jd6BlWqAtoso9K7SSTOyxBSkvGEaKZVSUzW1gllXRkDi+d6m
vVMFiJVXz3XciHyLa8AYfo28QO2rE7zscWKGLDZ4At7dtgu2HnyieJXNo9Jw/yjJ
Lz0E3TIzNWarAWQrS2mEV+MCEVsBApDGD0KSzKBhYlZ4h88R3CNhPYbS8VlwWUX/
vaaojO28Wc52MQT/ImIdTCTXmy1NX/k83CPVlXHFTi857qnxxj0dc/K/0oKZm5tF
wspQpUc90niKuvO3wx8o3Po74w07f9FzAnJ1T/qp+xYDLTtHJzNvJds3KLwzX5Fq
ZWRq88cjAlA4XslW+7Az+w4uOBcKLB4lGyUlMJXZwImlx/HfJo2CGFst06w7Vkkt
FDco1+mBKpDnzlaSx4HHsiGskqMWGwJYiFDetBL2+qQHwLWCTqP2+Nw30iM68WYz
ZNzMAbKMjmRYnoT8g43s3t66JSZ5y4PNaVj2Zvzjlki+qOFKlycxQY2QufV0mUWo
VwGCYZDd/H5vbeKQOdcdf1+KWRA1deU3aQBOCo2rb8mie/137meS0cuvvZv9rSuF
91y9CBsGaC7NjOx3j0CuZ0ZZF70VfEuHtsLRi4HnQtMEVspA7j+SXo8lwUHiUIpx
83dSb89zJbftnHUlPoIlosw43+Nwdn1kWn5up7lnEMr1Z1TkbkqEGGEPNn6ubP61
7r0GckV2LcmaGE05a1f63qoLx350GjV4epAS2ZiSgeZ+8hp9JNTs/iHBY7Bsfqbr
u2/wdmd+sf2bl/Fvl8C65UsBpVB3OLcOJHhJ73j6r9PUuBtfreynG75vH5WeDUc5
vSDdJkru3+y+lPH9wblJhhHt/PFJYpWChvWwpiGYCgsPA3BdBFFAp7rNqHkI+Fga
kvZNwspRg2yeGH88w90asDMjQSxmjvFF5GFJh0WCjsPuxwAyuOcQj3w5wfOsyIgh
RAK5qjvJt1EVQDqMLhcqOcTzZAX3/Z3X8AtOsmQmlZtTedGJndLLH1gbDaetfGLG
dCr4W17nopNs2AIKK+6FkgdXoHf+hPSdKgpY9K92aSmeHpr5O6QlqATFvOpSX1Rh
VdLIv0V6wwuI0STMb8DD9HjuOWGpfViD2xW8+CyhBwb1OUOaObTRqqN7toU5sVvi
SJFusQz4oZjwctTg1F8690w7khiSpgVVCt2BDF91E5yrz+5gqJ+Ezlx5TWs3ezW5
Vqgsk0oArUoGh7GD2X+G9yCli8+YiBzNErmZAvWSs4N4v/eAoKM6HIkcWwdr80EM
fG8sEpf3s9Sx11gSkmns1v9ys5ww9tZOZkBl2dgtBmCfB7Cj90UzNYUTR/T6jzTn
gD8t+hbrSc4EUPs0vRSOisnyOEhW+eeTr7QO4kFkJw6YzjDQsMrZG4A4KbtEx4MM
u/TukAA6LeTJf9yXHnJ9qbdghJb1ZvqfgSyFVwmyZbpyebIaXYr3N9CDBFqSlnns
I1AuQpH+/dXP+fKPJk5IFERtyTWj4Mg0QscYPkvoxHauoBmGG13EaO0JMGj52YDq
q4GA5Qiq1M4CYB0q10FDKTxgBl+GpqwccxNN6khXFh0bv61idXFrJzG3ai9Q+hyI
R8QoFi//L3lwserd8u75B4oABb2FEN3lmaGChNl1I/FapKdZh3eaNP6Keyi8IgIp
Ldkodq/zlslf1gGONclu94qj8/Lm0znOCUMR+rmLEkXqxPRQyXLKQrSjWFHKbd23
R6+ymI+S0QhAyrT9G6itaxwsV2eEYjddEiluBRoKFMr5qTexQ3UxIgqrVnYGiBtz
MzlE4gtr1jQlqal4pPMVYMPCGPiEmTsVypoZBgCWVa06i5ao6Skc0tpO0bVLIIRd
ly1r7OGN4vZ08VKeJCspSSIWrMNI27etnN7XzWICwwUyWi8DXKu7GE7vZBVXxx+O
sP9tVEh4mllsKXAN0bMlcpSpcvSpeQQBHmBkZZvl4SSK6lBcjpO9xitNDAKr7k5T
zQjwR7kXMyfYdM3MwrBrDR2KHZ3K3TjwXzBhk8FJsxboBRyVKNfU7GoF0M6rfO+U
ftK2MU78fAVF1iTXiP0hlZ49gNW26l+YApZQfnj7zYZawbUG/Wgy8Thb1clLws7x
kHYCZEihJbLRH5G2qUcr4k9wf3ioPytw8+RcNZi3q0YdS3bbwr/8YrB/5I9IwBX9
bcdEAtq80vCeFTGlTPYFTFjQ1ecGfvY8Qi8nQ9bhw6snZe9Dyu39liF+PaQ3EISV
ObqvdzIgHaGOuq2tOPLGdiYnnchDjkIbPqeoRRm21EDOcpxKvuTJEMS8iigBmdO8
IzKwd58OnOwlOoOtxy4rLC95kpySiq8vLNUuww1H6+bdClTfW9FOIHCG0LOpidnM
zFbZBEcOK0MmS0hGinx1Nr0R2W0UWYvY4oRKX5wLmJI0XHxDN7htLelsNdUwt7hU
Fb+UOFuZv2vdL0JAGlI42JcrWCSMiStpLDSDswZofxV9ioH22DpZZpG6N3FVCKkZ
tRCXYdKAOtw/k7gSwwsiB4nO2yobbzu9U/1ZepaNWuA0aw4ANQ5y8MOkE0O2UEIx
PASbBbVihM8R6aZyj7GBmUB2faLe00n06EzWaWUoot3zA6jlVLayrrx/487mqJgX
AVaHEJZ6CCNXbquVZwUABnLNGMgzd4f9BoRKgzkiD8NGT/SFIy3stk66r4nR5ClW
enDFYv5SSRmAJcqZG6ZvE4D0xxlOqe3UO9eajv/fqH5EN5yHW1judEhdbafCkobD
zbtv75oe39otOzVkRF+4jhnjtiL24Ji5t+RIMhY1OfCRlKVRgREh+OA5iGQpkSma
kQYUElccY0R5wzyZxp8Le8MgIHEYHiL3RiL4MwrZ3R+OZNTbfJ72051sA57cZ0LD
mNMKTJUh3uydmdbFHxrmG8rxMmIGcidyhnrIP8cbh29l7W8aE/6i+TWhME+911HQ
i9vq8u3ZlQH2Sj4hGFGh/YP1f32u75Ba6+d/nVjwudFPY5CJ4+AsmkJ0NkIG5/UR
TlpYVUc0mpalaTScuY15dlsc1ReJGWo53DVac3cbBzxFaqh6UxY6dNHtSGYl34Y2
PHy88nuK69JJzmgHpAdxtGLlM2S5JbijLr0s7Pz6BbfROlBNu9eHdOZW1IeqwPbW
mD45+XSwciCVpQ9YeEfHO0NkEggtuQYH8bR2Wrwbkr5MRdfX5+UwFnLQxqlH8fvd
OlkZHPTUxWZFN0/886+Fs0lgKUDb5selDyhuPJz7QccWJl2rwPFEtnJtABUoKmoO
gz56fDHlg1Mh5H6YXc4RlnZohcEr65JyUg77duuMA2WJsZ+RV3ru4uj3yH6kCuke
A2GTTy7/vshTtTIFRquX3p3Klm66JeuaCanCmRMzYXba/TgrOLfRx5CPxgM9T853
W+/rzlow67BA5RIh4DDhI02u5+TpL8dWyqES9JNiFvNGlF8SvQBlHHatfpVCv2AQ
aFqMv4l/88ieiFFsqhR9TCOXWt0cOrSfcervxn8eVo2mJx8i6obfJ9x0fGen5mP5
Zg9n2YzCTmR+3tsLMyoXyW8bnlHwsYmJSNszrZEy7XD9Ri8x3/gF6BWzA6ebidJh
OR46Ee/Mk/bcXo8h7S3qR4rqbW0TPTS1dOmZ93xHrAML2SxowIVcXLx9V6rbEoiM
YR40km2zfgSCr9x9ANAU4Pjy0VmhANwrl7Nsepmaww/0l0HtJJTOUn7iSoudF9q6
Aa2R6tcS61W1fTMv1+FaEjn4+stPkkWQnG3sF4b8D5cSqSGPCXtGxUkFV5uK5iEc
qNwnqbDuAzF75DwRvnpBbBng2f4UhZaodt59AfaajsMDG2cxBvqWkZbgZZ1mQp3N
oIhoCtaaoFlPJkwn9TpM8S4ACMbLGn60+NH9qmDw0T1OhJrj5T4o63Tzel3VkQvG
FQb3Q/ELRpZCtO4Q4GGo0Q4uRSKHBmLxdVSG/j9Un4xcmYSbK4o24Ydls7GLNGj/
tT41Zt+VWZlmiVfDOSoxY/awnouugI2QBTM6o3nWOWnBuWcbxoMpf4+QFKCyfRfp
btnRsgVAAD5jHv8FdcmPvafSEQd3jC39sJK/3R5bSk1AaQzr5/dAKTUSSODG7QDb
evDzicfd1sTV3pEaeNkCIhAovTg2mD8qc/kzE6WBdbAbugbzy5B1dsg5IkajP0ny
fEUwju2OqtIlTXVZ9izkeT1shGtm1A3CguNfSQtk4LID4Yo14V5G5OVeQUKL2gei
pS195bp//Hli2eMFDCaE7tEpFkkVk1K+Z4oYEtMgSNnW2rsdF9426FDLo5/Ls6So
aHaKms7r3FusyX6/hEeEy4w03tk5e/dzfvwX99kyOcFzLCe310DcCx4YUQbIWQ52
k8Tf6EkgvGUbD1Sf3jahxUfyYDUfAaNcjFM5vaa4sI+Lvs4n7417mCeIJrmGlzx1
3wcmckFBNF18D9DORL1kfA4uRPj038vEeo3DSpcauUjdomAzA8jd1JVDgj9jveUT
bsmY9uV/uH7oAkplIt/ptWTczhzcKRWmkyWXcUBCjaCaLCaWuP3XEV7ilD6C1YLu
t3jpvAqUpoEBlRas/barR3q3aUZzzEptKWFa6iiH9WfCUuxgqc3jphR8c3Ikup3D
8igPBy2RQr5XvYJ4IItajrUVqe0qxWkQfUynOGjI2lU1SFyJE69f54t9yLo5YaZB
SIS018w3rGeB64bYsk8YeYKADX+XKgPIgZWFyAATKZoC6OgHhlwnIQiZoiGNT7O6
my9VIZXsHT7rOXbm5QiBJcqlLG4RR6F1eK4WWbMI9yiFsZzqewheQfDB9QtbQNJ4
5qxWiFAryUx1Sw454CUnVbEUFbfV5+D2PoLEa7IupoB56q31Y28jXNkfGFu/32oJ
sRae0a1OjYRuuiAluojjQpzNH4TSv2+OH3IbihN6hUGJR6NN8Yn8MIjrcKi9kK17
AVxuco+IHHbgYoLVVo665lAVoRlZVTjmsqhu25n3wiZdfzwB3V7rkNw63gchR8f1
kgS2nj265GDLqs9HuDh/TCGvfFhQbAC9EwPA6UY+Szp1S4mnmvDx6Z/r6Qrbz2OK
unsKUZ3tbXLpeVAKmPDwobYo3p8B2IGQzmtcyKsP2hgzSFqaUJDU2G6z1wQa3GY6
JLgCUn/133BPpxaYJqQUIOXW7lOGj3/j53r2nJFwg3mqRucB6/CbMcFeKXCcmS6n
YXmRzBcbBvikqzKnf0INr4dZGtHNGan5dZiD/98LoGq8b56zuPUD9BINEyNOgC25
slMRa8raPHHN+YYcnhvUEFHtofZFV/GDOIjATLEUsh2T/XSI577t4dSg7dedereq
zHldcnrUD/I+d21QJLH59F01eCNY7biljLyewgWjFG0duifHakFCIrtFgB/Vb3Xn
BnlCv+bwn2PPcYYfaHLe4eCWS7L9D3j956cDXU9nVCSg6n0K+bpMBfr462Kr9zjO
+sZt8FSkhlWQltwfL4OX0FbnZIfUoVqqjPFNWWnBPkLrFGl5y8WRfLQ5cEnRJV8+
sYWH8XAm5+jPGgzX3/ff5jv0ZGe89wMNF9WcM4lWk1+IFk5GQAdU/6Wpi+e69YWj
CE9xcqKTik7LVYnHw07Z5mQY998d/jHGsxEeU/o7X80USTywZpIZutU67SAuL8op
7FlGSym98tuFVFSI4slg1ED+IqDRdXODF9mLyYD6P/DnbmXx7VP/9qLEtKFusQIv
E3VLa8/rWueEm3qmMSm5C/D4F1vmD4RSinLbqr7OwWAx5pZriJUF+rr8rmlK5oNg
R3DfR8HIxaK59rL5/kqjiphNbmMbZpMwIXzzOebRjYeNrGNPLIpSGnNkmiAQThlL
6aRK8CH4H7O4UCLpzw59Lipy18vMh40bGkA9jmroGYBW/9Ne3iAPW8AFBFET0FCM
Ekt4SekaUcHVTb1nC1XZs7hsYDze03ErOSrP7Xzwj374Qtfihrsf7NsnHLMUmsS6
TB7lkEEPpS4KQlQFGG7fEEx75yscIwX8SfCiCDc0qL8RIwvR3BfieXVT++yU2dB/
QlYqACjmt3hOnDxyUdyE1XLHXtcEr7TJIV3Lnto/E6Za8CCCRSKRBXZmTNiSMdSS
Lir5SVz0e5AgNmO8Wnn9IuugxyR513MWNUp6mvChflGKGAd5UPm5GV2MYes2/yM6
4M9uNHbQ69iaGYHr/rTrSY3jIpMul+0uFJCPbLHnu73ClfbYKJzZvDGWeDkVo9uk
Jk9Q2C0utKFEVofaij0iqTPO4rYeliVBPJmS60opPCo2KZGcRQL6RnFLrFfF2kk+
kZHWGmY5Ug327UwlbdhHoqvqm8Fiw5HU2ohJRtiVQR/oo9wYx/zYt31mToD48Op4
KAGoST/RVNVXzE7Al28cqafu1k5mwVG+lwqNo+zAHMdmlHD9gTNlXonuprYR4BpW
+Y4078d4OjPFlKjKq3zOg2Kug20vCwDl03ZysCMXpv6Qm6E87BlU48f+8DrL8PDN
1Q6VrnsuI+3cYGHN3hri3FRP6qxN4ccx33EEwbJ2vrU299dC638E4GDFP7jVM30p
mUVlseVapXBOSuDebYPlsV/ZAZTbVbtf/3+xEK5t7qJLt/O3QxuxrY0GkuKzR7Z/
zj8RTqqQdEyo4vIDwMYgFyXI3PYc5iSaKS4xIEU4nE2oGn6rvuX/iotKVqdCU3PK
4MDlV8bXJsqDCZP/t6FgT73mzG+DLXL54wtgbGrEGMzwwVglYyLmvCn6rFl9uea/
EiEdJp9D5lVgPmvlaq9P6y54tcbqHQMQmzAnbHtYnCbMF4czUjXAj+VkKrEE3ppu
SBmBj5BT62sY4U1OLWIgvj7tx2UZNfHQsIfzVlHHXKGCVvicTj+Zvklq8jC29kHE
RPHyO0QwmxkdA3L/h7eh1LiEqGxgQNxw+KOfTNXIcMOlAP2W4swEA9VLu3LKkVze
YHIH3fCbYM2D+Uw3ty/NeJH4PmgMgOmQycwIATwolD03cAXKc/4Dt1QEKfLzuJ/4
FDOQ5fm+ooZeObbl0k4JswjpzebE7TxjwRQS30NpMvkbv16tqg4KPs9V/LzRbDjv
MCZ+9Xzz1JWL3DavtwggfcFMD1a1gtLYVXQgJSq3/9/XwmMpDQ+Xrg5f99YI3W3Z
ghQ9MLQNZk91qSmSEOzRScVP6khDa1BntAlr6IbtoZf2Z8FHCTcHw6eTQC+t6Kzh
Urx1D6CfnOCQsqwwcD5J7CbjEbFM64K2siaTsVngUlBIIMWcoLLF+QausobwoNql
UteBgFbY8FCWBBAKfC2HQ/iS6Lo1RfDOfEO/3SQQW/712UIxFDPcTd8pyVDg/hNz
nzQN/l9d6vzFL2T1ZRMjVVNTMptnw3ijgf0yrG5Lczp8EVvP1+OOdOcEC4xlfGpu
Fy7t121FitCi73xM+qZbApkF6jVHzDPo98623lpPVvi3y4Gv/CP2yTZ8/BUPWA/1
JCUUxBYEwIb300zY0qeDiLQ8ECyQNFxyNGIQ0UGyVNA/EOsd4bstrnW3yM6qk09b
oAX64oPEH/W5RX8cr4dsKX2VZacNJQIqbrRu859nyyOrkQL+ZbE/Im96hwVoyM9a
K318V87+eQRDRk0Rkp9ELy3rVwRpeRFFhkCZvoPMTvNb8dN+2rR50tmm3FNvc8Ml
kXECxRnhrZK0o2LOzXAzji/XycujnDRa0wY6//AvUEavuQb3cHQBBrvFylvcMtGY
hy83zagHDU9xunBuB+eP6jqRuM6AueB1YomFx7CzfImnxt59LZmJ2WFfFf+xDeSI
dYTi+4+fJLvTtIu0q5dDoOLn7j95KNtnOfvWvgC+0ioFXbzsRYMsyrHyOo6Wx/OB
m3xZvz/6FMa/tJaIH0shu2qya7oN+jfH90BzPJtz9sjSzYWwAIaFQTL7US1i5VJK
T/8R+q9P8ph37VcAMpuf7V7TE2EAo/g2HmCWlEGnJ8530NjacRgRsmmE6ndIIAF5
sBgpAfvfCLmKp0mUtQNkq85pCjpcMsjHPB2byG1g8KTCG7K61VdNep50H3guJ6YS
vmT0nMeF8wpJMKKjR07QnIy3w/Gorx7XKgtMQCPjbDlVc2P16QgtUlnj0j0wY8Mw
yykuMasPGNrgFPWnH4I2aU/TYlh5toKwORgmDKiF98JavHSdRENvzdUNMljcMBuV
Q0r6tPBvyvyomtL34iHN/cJV3FHyAgvXUHsoJ2Gxgd+ww81O9UYsDjIDTLsXaaj8
K2orkKnwb1EEunSPr4237TiJiiv/vW9gVlRUhPf1a9ZkCCf4OJEcdNY6GTw4OcRF
9Jf1/5y/LvkaCRI3HEtQSI3wRfognjcgVnCRmQkpyneBGG2Vb1CsXLwaFq2C22GC
RA+jMU7QDvAwF/M3SEWq22EjS20Qg69xlg8jZhwZwidsAiPdsSaRDjqOygop45J1
zEvkp+BxS0kdI2lM4AZPXX4rhQg1NU5Hf79xcXYqrYgCN8pkqGIk3LGYFr5s8XHp
0lLmP2m9jrM9OM/PHawiOSJxY3w3y+38QEcos8/cCWnAzLZbz7N424Fqxa5jgVfa
sWd9zu88MTxti6n1XLYlvQFBVRVjc1Vtj+cKlQmOOlIai3JgHYw2oFpcyS27C8K6
k2LoEG/O7RqwWtJkiIdJEorSxngE+QEVUXU5Np+kSpEUIS/9+urIC4jHYPCRIZix
iQc5+jjp9kkWNKrbzTzsH+1MJkM0zfb2SidRzjThXndrAHpkXdHAR1YH2L+H6s6F
GYzZZJxhtbaU5FRFygKi+kN04AaON5kOLrMaYxq7KrcJDEqwnMqTpFdN4FcYpZCC
x2f7JVeWT6jzFN3c3f5zRpdjI1o3eMEW/03rSfxnnbg4TPyPU0aRiADeF9q+4aJz
FOnDn7FT2Xry8gyzo7GXMcSyYL9SO/6ZwrvdqE/o6mLO/0nlltB8K6Y/egCVkRw+
ukk9Bv149h3u/uAca2Cvarth/uoJpGhOVeGx7t0TrAcIbcKJvicf0a1oxfPTv+Ow
1YhJP0WWuyH6dmZY2TKuAWbzBwuzAurecT4gH1VUPs5XXV4X0TIgKA39/4DH87JR
KbR4XQcIpETJKLwVzrHlOSKavsnt/RMVUuFp00fQzCccsF1oxrOpc4VL6UHX5ATY
51meJ/9519wDlD9qu3aqjymEdT+uJOjEqB1YWZPpvtqCzSbP0nqBJC3ZeJwWlGNj
tmFOLCf6QU8rC3+h9i6cv5YZ/Uw1OEnjjbDX/NXNbSBxtYG7BVMIju/OqjFXYW/D
GqZrgK2XNn1Dxm1pejJJb4LsDVswkg1rEnYo2vGnBB59FW7wRXppSkNDTJW3BQeJ
LFVwO5hW3vnELMNZdxUQe3wzrDrhHTBZHeKQlzVFFse1KwuacVyMJf5YCGRRQRx0
Im67nTBU3lR09ET3SVsxl0/Dhn1IZTbUzrduTOumSAAVzUHL3icvg9nysXH2XhCu
L0zn5p5cs3F0W/lmb58YqlLCcAcigRqCaSO7S3ImJMDZ7D/svllvM624ufsnLHRm
Uo+c7gC3YjeS0Bg1IfzswXRiBffKOTa+duWtQECityUFW/WLe7g49BmYNRLOmKaB
3HXltT9oTRtANL3kbcfiiq1ZpGas3r0Egngx3bnTD++lPtwJqsvPAgBEEXOC2LWG
GYhsJWm0Yqbn0BBrVUJfLsuMLjfnr2sFKdvOC6+dFWyaF4DHHrdx/HXBJazNLLVv
heIaN5GLYXatkBmAR2kt7SXwOavmfJDAq3bKk4/TH0iYfWEfkmuNtNG/mWQn9k9g
Nalyg6ptqervY4MO7hgIwbtdHO6M9D59EpjR0IM4oHLQUpY0Gp6yEkS8UxWnwy9X
EOvezFaltc2FZ5LlDr10nWPmoUaiAAj7ApFJ4q90dr+bR6oipsiP+a/IefWbvvpo
/UDhMs7qjSPBpb7+FR3Ge0w+IJ7YsHI5LrL3yTZ3dDUYbRxLf4exig5lK9y6mtSq
hgxrY5OPkDvApkfPYdu/LEkwb7agIDdfU6X6gBhSZx0QENZusgF0j7utcrpf1ON+
bG8LlECrtOwxeXfyFv69Zdvsr33mOvHR5qM7naQYnhCmTDSQJq3NQbiY2cdcW0h7
9wn6H2wqhaySNHR2ZMx3AFi+0DFnayVIdg8usiYlJbmC5WH04G9wNDoN0dMGzxK2
Ta60HhIywTl+ufSndG+jeC/R2GuNNq1Z1Ab0pGVrWZglOFTZBp4NQNaf160+8Vjb
mArZQlxGXXcvN96tK9ANxHVW8VIs4Iknzo99F/ge5ACYrJ9fkgrrn7dLgGGfJK/r
BUGKZy0e5o3mUlzk6qAB9mOdhAvxT+kEhCbb6PmsCpSI+71AxHT/vrvUN10NDDZF
v25jPwqAlF9PPYwbpHBbCb1HWQC4TSkJ4th1WInEfM5M5MWlyIgG9pMmng0TPoG7
/fEOd+IDWvdREBZAA8gy9JDt2bnvQgfhKr9ekQ0k8o1c1QT21PldCRZjukJsceqt
ze5UD/iaee6/G+xURdkHrQJvaXkNZ8deVNtK1t2g8Lna3p75PXRo+kwfZ6UNI/7N
7CIxlgX6mcnjIZAWG5YwmRhlpAetVhlbhrBTTCuZ7EgbXx4z79EW0KzCjIzjJf9V
ZBjs29jU1XW0QSDfDG+PV13pFF05a1nE2jq5EIrplHo8mDRQ4c3Bc0ydtsQthhGn
xdGPad3SQB1dv8yviSBo3ZtRJ7C4WELmOVHeJfY7gbOy02ckgV5qXvYiBBQgrHRx
i54Z8pdmRsJnGXgogX0rNoMmPq+5U4yH5CoMWUmz8/s0X6SXQ8aRm27Kcf90tfU9
d9BXi9fpGMc/aMGLchMFP+vV92McggFyaNWbR+J0ea36XnsKU5T4py+74xS5S0/O
UHk3TE3kxsbvClWCwsqyPe5Nr5qgPxvuaLMl1chH+erOaSWhGd9hl0YAdHxJOpDG
vEMrVhWJgiXbNEHVZ/EOtxOw84sCFnfvLC0HCXvCUmgiULOrfVWX8TfDWqXN/svm
3rIUpNW5WVR3S0bOdFH4aZQtUArT2tiuGy8k06v2n8y9LvLftRZUUWMww+x+4O/D
JAoZVtediUbR5OEGcxExZkADR3DcWM/72H6IJwbC4dpcRlVbReamQbGyMpNqWcMd
prGBj8blaGH2X2Xkz5vODLiHVcoirqoAl7OLJ1eiD9/5SX2nbRcZBPwOMrbg7uuA
jbnpcrHQlzSAoIz9pr87+cz/1gDkQplD2SO42YpBQ+SydHmwesnglsHl6zUYurrc
ZY2sd1C9YfISCWzSLLEvB/eWVuyDXF7oMsLdVFWRpHf+yLBSd10uiEzZ0+H9/Ior
IUb41xwuiVhbdp7T8BgJvfmbQKKInjHsB8yPH/qOGdhPEoE9otM4WclbEwlBjbgB
AbRQCCDReB5i6HCBH16NynwZ8mP9x6+T2375H9CSCW2ldhhabQEpj5qbuuabSwnh
5XbGWKxiDuY87+pMfPLcSUP/xNCQH/4vfMpq6t5ZQApgaKF0GoFOFvAv+Dpq23bl
YKql75lckGJimXvY2E0YthGubU+5EVO0PqCi54mahw8pBcv987kILoPw3VBvOegH
oJEe5nXOIOZL8CF/HGLXGieMEa1hllt7YcjPK3JeRcaaZIqapAk5LowxfJNebcDF
+nK+JnyG/r5K330hu/jvEzlurc4G0pedH4GWyuQFR21Ac9DdTUBGSQ2h/21hfIbK
Nr6X/mPZwIsy1FpmSaDWrf7HVwGqBnDdeGUX1+BzjpRaXsEyP9xAwMAwx9jf40NS
ZtGJzAYEbxCsSSBlvGlmEDa7uFzK3PUdmaUlh6Q+mOigswypy3d+nm8TH9bpC2KZ
UNu7PjN7E9lCqeGV1Bw8AvQNbJaOcWzQ1jVZmjw1o01q1cTXgAbhZOMg3gBWXJWp
RZOGCXl62nZw6mLJfedqB++vqJjieIQVzD09tbBBJ6LIMfcjUC2e/gyyVkM75wed
fNUQ4BEmReaGYQyXmGdYBDJ4Xd9h1mfzfo1ERkwCOLkxN991hEN2guafJRNYTTBl
COr4IbAMKQigqLG5D8ry2zTQHSxKsh+HGDF1zEriT5d0d59GfPejhvZ7Vjo/74fw
TLnv4dg+Xnuwr/brjn5fopyAaKZUqQNJayxxiwKUz11CoyKHLwBZ7nTuPibEBPAQ
oTgtEZ4uUWaSGuV4h454tGQpVAW0IjAOURmeVr6gj6FD9cMf2NLOTZeA7skKMuIA
QTQRitruAROAvjmmHmlFnkwxrdQ57q+TLLsoEKLt1bOdrVm/jMV9tmFOtHKz2peo
3MduTeKnM1SdlgiT2kSGyIraxCuRfOYYG3dFh6s3pxWUQ0kT7CcAmEwlBk+2zzwt
q6yjTuAMJ27KqZNuKwDkbVtELiIedMRSQHEbh1vPj7z5+WsEIf1D4VkNxoueHzO/
afcvu8Nztq9PpbaNS9xMRlR2/MJtmnx+kECmyBcbF4sjyRUDQn10s4/GuMUcaKOG
m00foPdB2QPFZGI+RWdzkdVahokPPpcj3fHg8lyOnTxwLGR3bCmYH7MkiGU/KNVt
fpKXF/B231N6gpYLns8Qt1jg5r5MKDaPCIwjFT4mXm11e4qCcufy7ply7/p9BjYO
a7jqi+kp67qFnzsQc30gT/+XdXSLPVAZ7HqA+6aERps/uz0aTTmgfkHPEJTG5wkf
PTAW2qi/fBE24Qmo/LTvrEKXPbijE5URaqk/Ld5+pFJSZe+JwuVDEzjGkm9qXPTG
6HG5Di3+7dgAFDrbU7LaCCFpVTZlnp37pOPrQgu1PxPK4yiLZfyPi+TW1NQD8LYv
rCLrJrwpxtW3QlBHb3KwGpy5yYZ1eZCYK9L4vE9fuvVoOm+cAmZCUZAsAkqTF2OP
MwmC/WswgGIjpNbecvZq4zAQ3975IWiVO/tCwAKE0enC/e9e5T384fribClAsP2J
JPZQvC8TiOihx90U8b/L/3sWQV89TRTUt2ApGc/ZEox4RfhLpHCr6LFJ1ZybvBmy
IoCFauHfCeRTgadG8eq8KwEfTea4KrkmTe4WNmXZeRxV/840acxctijD2tMdbR30
OePBraWZpkgEXPPB1T/VDjpLjCwKobTQAYKlKoOwnD1fc1S1SUVse3wEfh+TIC4U
6y1j2W8ia6a4tp/N5PfpRuCnKyxA3PiS9tAsiuswapV+nGGarMfVG15j5tKFXhTl
AFMHfnyEG6SBQIEHZst0hGWovq4oEx7EeHFRl7Jssrbig1uNFvcRScZZFiHJ5Bh/
lAh2JFkGtxExwcefjUKBatpomMlumffK1amLTEODUCWvdpKl3O2vv7Q/UkaPjLYs
XBYM1+IW75nmidqRh3XKb6yXPdpPDRSSSpXChPFO4BihbiIXsn5IjX8n/09R5bwW
H26OkA4wxBsQE+K3Zcq5wPCVe7jO/i/8xJSGFdE4qWNtlgF3CUyPfb95coWMdXAy
EVyOs+x8U7cWDb0gusQ1XMyH7mUl8da/L9NIQBoGKGyUqo2Lhjq7E/I1NNRpJOVB
HlDM75pMsiuEcFiekU66ZgO4ldCvU1nAKYkxeNXfqDC4UJZmJ2zjQoleRJJUs085
3BOF2+F3APyUtxq2CKx4779XGu4b3mG0Y/9fdaBcPNZxmj4PDEqNhFik+9b0tKHu
XgUoNZh11A3j3Pa6XO2A2AalwWlxHQ+d3e02sgN0I8wRb7Hzu3exAI6bmYgij99K
UDLnuMa/6BUDm8w6n1/XdHbB7vBq0JzcGWMhHyeNf1vkYrd56CuvYAz4EerWkpEP
QqT12oZpLDx80N2oHRoggrKAGPJ30Vu9QOul/hLmR/iXJ6L2QYNvvggPFmQmHvja
QFqDjGA7Vh5Sgvlwomw54GHuLN4USHt2HIRRlCerQWMh5xe9rfpku1rVnd3vDO6b
jEIrx5EHsqFaJphMG2K24Sedf5iF1AXwrZ18bO2sXHsZEDhsTlaS4Q8FxYSwYvMN
XKVJzbH590Av0HTeMXhyVEYZiGdiXFEGTZuMUthbQHuvSVX1nZfq8B5nRAyedS1n
YAB8q6QA8p2Y4bUGEw2XiyTeyi2MdEjkIIo6b9HG4xZKGiopiVubIQK/JDcPBLQF
LqMUhrgv2k60wNBw0OyvYwwF9uZeJapU1wAatn8Nf5kAt2rvzgmjf4XbK6xDYGtv
17N6yngCr4T8IMzHnfgB6yBzHrNOeFyWORJ4GCTo7kAPpyUW3TYW9JAj9Ct1zrVo
kk89sQFO25U0dzUp6AhxREl13ssOJLTPd0SYjgnk/X7UGfazLhnxYj/c/hMmC84e
ErphcIxWc2Y6uyOqd4CH+K/7u85I9LS39EkgZWCz0iIrh/LJxgVFLFy4Qpr/FINJ
/RPFtVg7+6e0FrC7/ubWoAVNRjg4B0rF24V9POcaC4gJe/MxnuXIgu5WSabYtO6L
p20MnQhLoMO9ZVSW6osuyMnDh3Q6+4SXY8u35uH5hWXfEZyQ8HKECzJI5zjOCPyp
dVaY2CNrDnIIlTUBo04qNcYo/TB8HL6QU9L2keXuSsDZZNMZ+ztIOYD3nGJA4EFl
xituMH1NxHJa8KKl9/g/qa/mp4xm7yHZmTQezRl6MiFjB6wbBnn4NChfuzEK8Z7Q
OeeTMz19cg7kU8DIxr7PfvaVYqqAZhRbeBbVUknnuH2d+SHZHAVplF98duXDCeD3
vHZLZBOaFzPFaMGXDvSIIj35TycSUsxQZuWXCyatoqHMQ15dFfxo1aei/1IrqMCk
oZqOTo4dAVMFnZOfkaHzyc8DMmLymXuJjVqih++aTqxY4gVYuZ8oo7PA4pp03WVX
/rAB3khhKOyvYHkA9w4h0cxodwWYqX0pt7gmU1o7SoxIhz3Kb4MnubYc8kupD3JG
nurBvhGqSIHHrcckC7WOU2B3sauwJAfPyXtzN4rQ9HNM1IOid9NQptu2qAhOSNfg
um0YVs9kBn0aG4ctQdbHzYW/XCzB0Z2yws4nMyV4BthjkbDvfCnjd+d2j65tzO6a
CLbdbCgpQ6MfUEAu1LgD+rueaIKndyOi09FpbCJ0sUwcFQa9yg0c5LaanEqiPhia
r7zWPXGd6orE4OV7eAjai0hhR7xg3RGOWQcnVmBOD/7XGJ2vlf5bW2jXbcPUyFyL
rdq10wxRGWSvVPbUTprd9vB6DaOCJGO/1Y3rliA0gYb1uanyYxAKxUnBFuaKT6E5
RHQ7Ads2H7eZZKjK+VoL99q/XLPrDBhJfWps+mLGgIlKas/0sTppy1JuFJs1DyIm
pqsA5IpAk2ByHxllRHPy33FwkPpCyes2qmJF+cAY+Esyc3Rd+cr8mQxfCvh2Hu4i
m+0E2yU+pyBKI1eOLm5r4pTjpRkU1yM7zXUmbY8N9qzEVcWLv21ORQeGPEAnX2+x
E6NRiTTeUD6L4BawXDfOLmgGttDfhb9gRRc5VYNrpEgJcxgg08rQLzEdxLOY+mtT
4fwWG/QE50dk5vSEQyvTi1y/ErEpj4DffgOwmuJU5sF1OYxF3IYGwqbX2jvuFUEY
4BYe0ammTUzilB41SalXkqRRN7r77CQ1tTSoQchMCWYeG96tJNyOtVH2d4BSKgij
hwlQCuWrZPrLONC/Vq2v7xHRZkLr/fI9ZGidDehBqxkcpKlLbjpJyOVGQrNBy7om
fBowbmf5W2gnwuOccR89v0uzfc44hvc0io/mWfW2cWw0dIMdFJsxU8bOJvFl+aLz
5Rd4RXHOgjU25lr0oQTZjYxxC02zofqJ2ztCrqaSc4F9BTMVavycPr1iJYcoNqXT
YxmVXrFlnQBXbq7aAmawq6lEOGV/XKYptwpk7SdV2jrZYF8GBMv0iewylc593+YM
XQRBRUkFcmtYeMMQ0hRUUjW2OI3TsdSgMA9AZgR7pYZjHzLQzzWLsftOMhi4iBRk
4c8WuTFTg4DA5xAlXoaKfKXiJlB9NBsS7sdUx3R5sMIW5Cnf57wy66yDIeJI62QZ
cpHIUsgIQ7Y24zEtkZDfGWK2V75ReG4H/8S8g00FxnxSsLk93nWOTYPlS2sV3Ge/
XJl+KJmbwimR3SAtZwPF5YXq4mQKsMg6OtNe70B2OOyEMdZfbSJbQwK4yZNFiPG8
odtEH3E6bjY2bUt2wpdVNSgrd49blZ3I6scC0O6Lq3jKzvIVc/8KDA7Cg1Fq7Qxp
VyRfFbsr/r4h1Rjdv8kVn0r71C1V2uesUDNncJU1vqAiZPtQ/lmLKhQX7VBSWKYK
FinOgF6UUkLyvOr0FCU1ySfYEExS0O667tlgG9VoQrOBOmMfZRkxt5w4ggWUXgTQ
7SSsPuMWS4ME41GZTTmhr/49yUBbRNNxHwrTa1kKj6E+o8BIp8zuB8nGZRIolG2M
pJbg27wkAkioWitFKGSemDLtp6D8Aj6XJX1Wiebs6wK9m0xw0cdiEAbbEGPorRCj
Y+v9MtOBmjIK0+KDtQVuuSHEsYPspM+K7ts0gp5f6tWWucfctbylhlu8zxbmzx8y
kDCjO4QmoX5SEo/FS+XMskqphMjsEY1k2TxRMY4xHbaskK8LoDo8+/ie8WcTLv7R
sopp7aQLAJQfVNurh/QIr/Ps4kFVUFB36UJjbMc8xkfrjayUUzA8uYXBeFpUfUU4
WtXjT8FAGEdIdt+KASMloFRUn9Jro/bU2haigBcnDwaUyvYSUrl3dmlgkhW7ncn+
uhJl2gldGx3BHxGITqf9P1R/UfzwrtAxzfp4N4ssN6AiuLSTqg/vMs/UnWc1pYWL
S6KrI+aZUys2bVpBFXJl3ojfINZJbaadYayNWqXIccvLXdl6s2tMZCrNZscXm1Xn
b0QPEPI/DBwjSa/eMKXjQyHgI0Tht+OVqhlwAV3VqCrKOwpqBHwjZGG73WOgvQsZ
Fe/ogKF41Wpgw6NXaKK9IJN4p9W+T1UYq+mO6sxrwHhEgUH2RTXWYjs69GVaMMWH
jpzO/ugVDaXO7334PqzM8GRoOUnbK/uLL44r12mtairPtO593fsGrA/9ep3I1sxE
Oo/EWjqkRVsRGa/pkF8slabCxtl/v5iSUfoyH4bI16rlmcfhCac38iii8XrBYOIr
qB9uEjGazczrrY08tGRmAl0oRmTkBtWuyVaQsyovgGm4wXL2pxvbceN112hnSlAT
SoV+au1lVtHwb5VMUsPchaei62KcfgUQqDiPlpfKnwnynpUNmerLOizoPaBHS2jB
tXG+1k7frT971CMpmm5kc82jgVWkFDgqi97qYCLZPPvFUuZKbL+UxTVgdq2DHkGi
6cSbMRLyYxptpZ1YMl7WhmCAGN4gInkX10i6C/yWP12p73klOUHuLcGdKggC8uc1
ClwCd5DR8ymntP5oexvdETNzsaRYdx7qa1oNE8sQYPWV/vvz/cjEIMEE3ieMz2Xc
eL4zZrf3zzY+BIpOy6r/U2FVli1WZEIsegEtzyh1D+hpdWG+OGwFvnzTlAKtPg0x
lzAlfupM/0LVUyaIdsiOlFhMSFU1kA9UfA8YdU5jJnEA7FGjM6asu/YAOWn3v550
Mr+5fWBVgy4n4ABRxKnZS1HcVLqOhnJgBrtWl0WxMTfSVGHojxNCKMr5WX1QBRXr
LAviip8cJNCKb9Izgzk5xT/9oIPw8YanDWyyFXA5vkKxpQUDFkLCbnc0ZedcXi/7
yUHdMpbdXjWKlkj/5M83r0VKeQH9/Iw5Y1VeUgQzO7X2Qgrpj5BKgvHCFwP4AWqk
bVBCDd2J5PH1dyLe85uc7Kepwd2bNorPLBPWwgPgOXobNlhgHytn+3re7K1Z/vEs
vJxvyjMuISVSz+ST6bJfqV6ahmecWtf6ilNUmYYgXARpwLvKETpH3mCoCmVwrHTv
ffvY6Ac285GVkK1MWChRhBRHD0nGc85iPdBLVr4eSDsjIPmamqkP5ouUpor6IxOo
hFrkO1FSrUmfoyzTCl3Xeztj1EqKvDpYVTa1oAXb+0Bo5yh3k2cpPX2aHStICJ8e
GOf8gXaMJ26bW7grhLZVeSMrukjnon4V6w+MhccCy/xIxep0KUKSwGV4ed9OMmEs
XuwwJrBvY5bifFyjXNt5LSamAN8TaDPoTinb54l0NfEvNTTR5Lj6kFAEe9tsW6GE
pHxK32s8A3qFtClS9dLhjxwjmKbsLb3Nai5vDPMKZJI/squrtxwhc78WMmXog12C
4bUYx+xCrKuVrz/3XslsQY17z8neGZy7k3EM2piyZuAja2cIOTbCHNQO7U8ypMLv
UoDtfStagY7jZtCYNLoS+Zax5CIq8yt5QWk1RoMrt1u/re/YyCo0kw8o60c5SEX8
paV06wpCmTCnyb22AM9Jne7DN8g7GM6CN/9sz/4hkykBqQVyMqbvpkDxkWIvoZJs
QlieXxpiKO6Q4U2e5ViYIjhwpC7vMUcaBbHlRkeChIOfkQYVNdAlDrRBvGLHFdVi
pUHxV5f8JwkKNTDZa0yYASrXStwuPl5vpx8CFDFlOQvXzNxG2u1dP+SVuGSAC96p
3zGiW6QfRl2DLnP6MSNzcTqkG5Wh/AR3T1GXtToEMprodhWcRobdfwgZj5Bdmygt
aQSvSEuDPSGZa/urcuxT7Hkd6u8czyHyar8trS5J1QuIunwDAQSIweQYa7S3iddT
QlaeSJyfXhuCB4xiLnzum4DPVx2XQ3ehUygVl2Ocw6rto1ScvQiuGOlXfCkQ65iS
3ZByLHkqA4/e6m1TLpnpEusiKJeyo07heRzJVUlnkeeoCp5Fk8OX6oyQm0wGtxGC
Ux2DIEKVHc3Gm+buLK24DpIjd6FCAMs9vsbOzEMXLmR753ocNYr5408BL3OjAubu
2ZvOO9eNA9O1xL8qz9BvoHHsBexNnwle/kD6c+WkPhHE4eCMKV549plg/pJqEiV6
Gtzk7ggiY9BJjGRaZy30V1CouaZhBNlYua9F3tFcip3a102wFP2oGQ4qKAFV2gUT
zs9dgtk8PViUFJmkU8jkPzN6uAZ54E0ETpIXl5QNcFRyP/6ZM/9jCrWMSeAf6LgF
u6aAYnTWRebiHlj06H+8Jqcm7oa9hhvfU1Wjk6ZQOKcwoHKN+to0kNAXvg7ut7CN
mNPQ/rr40PG/66qUyOB5XPQ3MF46Zdoihd55d+8XJEfF7WX/U1d6mwvYMPM9s6Qe
EqxHmbop4L9z5mkRv02WPXuXypv1n6Bw0MU3Sog9z9mXWCr+5WnqM9Gdb12a6wlV
auIvp0s8oVISh2B6MuUQOH9OufvRMDcpTBO5D/O/ub07auXQ++kUncDYpVJpYuES
XjjwSzqSvp6yj/H5zzDIdN5avS8AZtqpXIi0V+KK2IFoDXVLDyuho714MlhCudab
u/0MuP4QDIbsenhhYSpxTrNYtPgoo8DnjWptfRI8Rf7L7phoVX7dBmOqp7eZsZe1
H/Ted9z1at6xft0Lp9udMBnXa2Dn5ByPUK+hm7nSImvj8vV128eVO0tQ/U/GEKuU
3yBbUni3nGQitEP6N9TXZAnmmoPlAr+T7XFVffa3NV++1UgZ8Tves3gYkqNx2pmi
3kZmSh+aVqd0Atk9mzaNLRxmFqHiecTfMFQA3bkQgpL4t0ZcD+H+uNC92SsnvL5E
JzBzviXW+dPoIQ412I0Nlrt0HKCdGxyBQsXEIwBkFzwVF0HAVXP8F5nLKQiEmGsL
mJXYx7tixidk1rIIuTzZ5O8Aliy6KBPGD4EBZ//JFHifMi0qvKB3mkm5uRMdcCma
2uNOvRSwpkgmEMk82HUwXU5d9lF1+u+4ubMJyopBS4UvrwGCUMNzuTFevNWTsShI
H5qyR6418dqWLRF/7rJrZUYHsWm56hjSgAs5n9bM9BUuuvviDhF4AwotRVhoxtHY
+9ZsZ0ERNXJztBtqVq8cs/C/fnM1Zn5O442CjTYuQ7Zaa1I2JwMGYAwlzsK62/WS
V55KI8mUTdAab+EeKF5QxRNpJBbeflx1nHXni/jKHuqUkJcdjjJh4seXfhvJiNAv
bgjI5lJOcBfglA52/JqArKlP8N8zYpmDQnoYW+T3IZXxBrGapGSC/F3G1UEZDQ/h
bEqbLdaAwE3Ve0QRoW4IeOoO2FbMbiHzylTzg8jpzGDIkh64MQ9vKw7vIXp4KCc9
LZJCA040IwzpnatQCQIwsIFYuLsOYNkyWxQKmREUPhIYqrtsATnUJYhMirdoXG0v
yoz+iFHaClhJwCOHQ+g7AnIsTO6mDW33sWWFLPrBjuu42vtQwpEcm79s9Mb62/oz
Tb/4kPGr+Ccqd6tLpwh039nBhuMbTbIHcEEqHLYnqcPvZ11AzwiCLFrdEU/6ayKg
s3CnOPU7NytxS19JnvPsDt1FFCU+/sCDU2TrtX8oTn4jF2YFbPI83sPNs4JU0jv+
j6J4OG/j4G2yLxwjD0QHiTKVMMa7uc0ualcnc4XQp4lsAbtmOLmTPR2+d6yXolgn
AjNj2g7pXG4HIsVcU3D4JycvmzU9wn3/Cdin4moRSr+7l+zP/6g8/w9aXZBMbkFZ
qlEEgtOPGsG/wgGud5k3KRIXCrPkCKb9uyNkU1tMiTY1T6fiuTIGUb99uTjMD568
7GTJgkFj5DpwO8xYt7Nkd1iGi8gTUP+QNdIcr0Ti9yKqy0yADCM47qmklzqS9ozM
E8k3DrVRpIKYZ/80IAIqgxbyaBLC878eLBuCSyV3X0pRU46LQxe8k9JcqaJDaHaK
nhYidtew71EodZx+W8K3hn1Y1J8ujMwdnraYlUFIpDNmJoftxC3GtKtisRNXqM4u
tVmKUFH7c+MIlrpmKeBWoPiKhJt3y1F/d7x0sJr+ktY2757b0/pJHL0A0pf08P8T
XP36dhWCNqZv4jxnUZxSiEsc9TBuMYlBeu7EXUUJ9hxS91ZMNF46pCX4igWnh2xq
xSkPmF6YUcfG4HeWIPa6O9Dm8rkVrVeNpHPvn0w+5OQyS2qEWD25mda69VofXY6k
uwKBMKc9G7iBPJbcL7emHkgmf4UHMePyOt4ehd0TemS+4JonQSiAm+6rFnX7u0xn
CwEQLrKCsepiVGlYAOud53EIIH+/GPihur5lOy/flQLhPrcg+EY+N0rOpGvPhsUz
eavQSXvJTqERvRsprBqGEYHP9AfrSjvrNPNQ9MhntO5N/9e1QkJcrXa0RB/uoMDW
Mw7OMo+IwH6Lu9pMHJc9F8hjOhWbvKeD32B8iOFDTiEFI4jwMen5ToWrcPiShDJx
29EVhOPoTnKxFcEC2nVqJHj5juEX9o8VFtkCM9xViMz6wSvHEPZ4n3T/nLL7IDCf
OXxF8i9e3ftcdoxSwlcLWjVAxfMKRn6DsHXHx40Px+Y+p/aPAxrTaNlJT2qm6LFa
tddZnciTQCa+hZre4XXQG35mjpIXQnubx9bJ84nhaeiyeIa9BSY1ejQDw4yZw/XE
dTAI1QZnZLLZeKbkEPf37t4eHloTL7mfvUBf4L22W1LPBvzQorAELSCTn9t2efc9
Z7tDL3ahcwwDgyl7rbgzmeA1YE5ykdPyIgpsB1D49fdIqAuCF7RNy5ug3y/a+hm4
7sH0e+9HBHGIrz2dX9ib5EaA5qSxMVzJZhIBCtS1aeT1kM3eKEsbxHk9+UYYzA26
I0XMWN2FhSd2fnDFZmJxEINteqRdFCcn+yfw06AxyHhxSfCfFmsgpDRtsPGoLVLT
sXUj/z8KBzikPnb0L9ERt3wzQQ5klQNjQV8LTrxXyjWoNj0118TaU8J/aJ9wuqse
e66ZDMPirZ4LMWKP9KDnIb5iY/rHY/MGXYkDppZnVcOmoUZekbA3FSNsvZer2cNO
AIXcZDcq0y1BeK53o6WE89D3L3+6r4MhL2dxjh+rRCwwDYzwXw4gR86gdOHyz4qR
HiRRgJ2f4R+lzUTueK8Rj5KozyERHlGoc35+EzITXKT1JYf/aLZUZ9aVVgCKxakY
RB8780dQJ0cExgutQV8nQkNEUllfZ4S1VJl7AXYXeWzZZAIEXEqAMVrXL0j+VP1Y
ww5pW4/RNUo8hxfMmmD4o965ky/+Qv2DDL2/MMGasjDP0iqvsTyCWKmSiS++a9uk
H+UUTMMDO2NmjZvoaAZfrHrMwVweVvdCinfYkOx9yuCf4WYKOFJzxbcJ0QbF9Igt
e5lZHJ3jRIYVQYMH6bx2lCWvDoN9Bjzo/d2PBCFrg6A2YvadMFxd85O72YDwl75L
tLtHqM3ydWCAgSsPfVETlLqyAVGxAPVswiphbBCoBaT/lw1+ZJHF4g2eSxpurtVX
PyPut9NLNMZqJ2FZqqHZFvCNbxNEsuUnnEVY9AuB26Y3D48+befmloXJEk7XSvOb
A8/J+TWtED/DP9Vq7pxgWKkW1mVN9lR2a1aayz/2Q/kYor9tHZXjuQAG9YcMRHy9
YkhK/IVZWjj5rcGzkGyZpeuDpNYacedKSSWkcAuLq4PDA4ZLIu1phfQCCAUmIs23
mSnSrgMaqpu5T4QF+gsy3xnB6DZ8e26qExes+4TEKoMMOLjnozuM3ZUWVcZNnMse
dlRIE5Eo+8h+/M8SpMWZNlPFq+KQJUAmMmL3abYHIVwKBBeW9WwW6CUUuOmkDIlS
mK4EPw2ny4EN19LHuAKSLV4GKPK7KgLfIJz3mHb89BKJRj6mcf6QzynvESJ+Grtg
hjWzXQ2WqecAt2KObEi4oQnzkogulg1x5MuhAQ2YqKX+X8cPFnNxZb/OhL/oybSH
2O1/bHRda28iksqXOrV21B1XBAn0dZOIjft+mMdqy0kNGpJsv4XBQZOzaa1dqsZq
pl9iXnvszKmelNiGpltegE5GuvDbk4gi9bGE9ah9VFUNe9kXkIUswJQirjB9rJ32
dirz/TuVS/HHcor/6sREn3a0YXeicHaycQk6nG0cnr5e8b0X7ie8kE4MnSl60flp
4cBz8Arlz1rQIMClwTMxjMwMmznY1MiYzmQPoXgViJpm5Q9n+8HqhbCouTZRRrk+
loTLfvUyXKAlm+YVBiCPB5Rta+lo2ux/PD+GLANHNf+sz4U3BbcRnUCtUfKnt9GI
9C1HQ/3veJvxTydhAvrVuwFJs8eTQTzbOZtZbb4GA9GW6ZvRc/zF8VWybJWVk7/T
8ghEGP0qM+vK//JEAjW0TIeJ4id2BU6vTcwMVNoNzQpJ70ck84do6teDxyAd0uvB
A+oRAWfKRWJY51SPOuINEp9dQDI9G4DArpp2B8ZF19iMb0SNcDUVX7T7A5K3d2Zw
pGO5RQp5VCoxY2m9fb9/QK8kFwF/9alRd4odIYK74ZW8dsyNym7/JAqzakf4hXH7
dqXLUyjZd5fO3YOG4kGWSV8jMfmEvM7DmNkol91SdZCMpl+E1G0VhkpaQ0AFVtQ4
qoeZugIYlVLVDh5B5+VyhWf+fl7vpL+jW4HNdpJoF0+a3zgSQQcRlmo5krRw4yrb
gcoztdPvBDraOz6BV0NCrnzd1CZE0Avg6aUoZOO06fY+pqBSEQ2FUARykWyQgp5+
RAVMOBaYi22L6nJDy18jEOqzdLwj/WAzDg5IOKnrPdy2wsTWMwdb7A0/yIBWVDas
JbLUVTGzGXmZw8jjJ8MQbHwTN5JLwEC3lrr5j7zod0ysw/6iNVlXwNo9Nz+V7OLF
6E6ilhm9nKFfK+HZVcpSdGCHc0ASBTMFFZqhDVWvjsQfFjgkFIDNDBJU8uBeVwmN
iBloi/xu2tDxcxAvgnS6yWTs9Z36XfxWVVticY/lRqziw/4U1LjG6EBmfItq+b+p
9a8Jj8z7Ial2vKRbJNJsLIOIYooOCr8rY/uGtyG7ig/KPRwxYg78HVVnVjTs5dTU
dCitAXutniTn9ReRntYPllOaURDiDZtsZ5JO/5YX8CWhsHISfCPWVwEr4V1HUCqo
Shbql4B0Vm3kmBu7FGkius8/uG4gZNP5v/CShYrRmVevDwWW9+Q8x7yO9nYtwTn+
hL04IYvKO0f4yY1XPZxdSOSfjebXnHVd5cTY0pb4yrENUQfDOONWRvqs3uPyWdw1
dOjF0ZDs2e7IZ0c1/XU14y4r/8FIxzaxK3Jfll7e2t+2rhsg+7fMZv4/dxzZozR+
S1pZDuOxgDdc06zDetdCwLcCcdeQHr47FOVvC22Fy7XVUT85KDQbTnKMJ9Jijd8j
0bDyal+KUuM3L3Awc70tZpnce91qmTWO9neO/eAD+MMRORfF/Q1xbgrG4YOONJ1h
ZxW0ggZ5rDc4XcxVGsncqlIZHBZjEQVJI7sho4WWSH0NeqoZcZCYMXdbftZeuRrt
m/q8FR8rgoXFmN269NsPHQDe/s+LvqJ49ixTMleMF/vt5cK2ifrkt1eoAZl4gdmp
jsz47idcd74mDXfKNGcaao6+6e7IJiBvLr9R/6QD6sgAuL/xaCandzbqmgyBSxGW
63W5cnllJ2PpnvGZf9McUq1Y1xli6uS1wylAB93V6sZW2nuUUgUTwM4MSPTITody
rCrNC4/9I3w14S3xnmeFV1+P9ASp4iOtTB5+eCd3m46XFtB+uAdE/G2HLw+ozC6i
QMv3lsQlHGsTyAKTcg7G4DXT2KkwKuD0rN0oXxiZAgksc/CJQ/uTSxuvOC4MZqps
ZJ4TBGRHPbF0hSXBZsPvf+RbYDAJMwrVQfe+SBxm5wMZnnaLAN7uoMWFITrAih0F
bZSSROvgmc8OgAusejLK8R8b2nRc1+pHAWE3cmUNaHWj3Xo+/yuowcoiA5TXQuSY
T2fyDYOl7DfuAteGVekodmE4ohtjycI5I85/NhR1UXNgBHdkOzkwkWwPuVZ9GmTi
jquConZZy/HNFDJtbgZ5VAPer4Ov7ZLaH0YJO4+fIBxmEQ+V49u6Wj7Wg02nymKT
RfKsu2OE6UIepvbgPWXBPzO7vsreOn4NM0rZTgpOfdB6GeRysMXc4m0OS1wSWkNu
QA2qR7Pemeh/WyPQRzFyHD0mx1VCmwPESSr7VASH0bwAu1VXqa54OB2L2RmTA92t
hM3rtxDEaHX+rh+v9wUHwM25S1/R6YyuxjR+LJYKyg6IoOFmUr8U9ZBbJEG3BKne
XCHqUpBfFNsZTx8qv2d8sYQoQ91/XP5DMpyiMr3a22CJRjNvu+o7Nrq1hrnwfNcT
Bx3EivyBbcZOMIVaksRP7+h/Q/AZPZZuBi3njjj76Yuk1wNDnaJyDB4BeW3r31Ni
lCd3yZ0jfrcOZc13d/Jt2IDueZOvXCoBsNFEbETB+JHjxXXzCE5QXfF/zI424+YD
2WJ6tEhwmbFh44OeWAu/WDPn7E4pwCgpOfyw0sDEEH7tKK0OOrUNXn8sD7TeTa5T
C29b02i5dHgaIMUMBKLeRbF1bN22jfpDU7/dfr/Tlp+S+fzDeCxmvhJeFu/egOGd
nI73n2Q75treCGa2t+jdMR0SnICGQ4zmUpsOsQPlaW/IBns0csRwpq872JcdzKg7
dt1a4vcxmWIgDapLBHBBFkxYq+tyDgyemy/waJw88VMoPibUloDGCtvhKDEPh+c7
gw4w0uHsPd24n9BZYtGphqNzQGNmF0REandy27y+ym7eJ9eo/Ohclki9O021BXkk
h5NXzwHX8qPt01s2ICb+5oI6aa7Wglzvz0milsgqvLjm2EQW1BbfCk5mWACQ8tjc
U8X/k/Wb3SUw+Xrn96O1aKuGLVqjWDFHCAcZFjtX8If4V5YKDEohEjb7QsP+E365
t8ECSoPPiWDn2AmPiWiYt++EuTACMzcbBYsjetlsG3xDiw5AZJVK3ySCABuk4y9V
Al9GLqSYDc81hwroMz/isR3cnc8ts14qT7oATs9OAWGimyeVoLQ4g0xjPvIZo0Xe
zAx0jJy20tVhIbBA4Qa4Zd9bP5JcQkwk9QChHYBDSoOZs+9bEIC0ZFZuMpx1KGtZ
A1KJHSrRHXHLE5bgByTshA1JDAmtDqnqMzCTz8C6jvTAzXlHU9pNq77OXQ3dzCxR
diJEObiMDBbIm5BIShpbFtqlnrAxyY6eOjvffbbP9ybVJTMIn1ct4i+GJpOIxZ9J
AVZXUYDkj2ykHOJYu6zAU1LhPApu1VfPKHsorDtKnV5MU8o+Ty5vUPU1soAtyGwa
haNSZVnc6SC+qhMRcc0IUSr6xLxk1Uyps5n/VS7f7rP/HgeIn5SrPH54Pcddg0sC
Bfz5G5oO3MTtmhLKd2SyP4KoUsUTCDbeEb4A6bC2mxSC5gtO3X7Lci5NnvMALQWV
ZFguKFNAEb1FGSWedhs9bZxjHlSSjkWFx0LfH/TKdBIO4a4xe0xkhI0i0X4ZyvaR
fqUyDv07/axvixK9hBk8lbgTZk9qBAxeXQPxJuNghzStMWP/Cla41DPRCsfcRFLM
TSfKCLW3d4JNBVE96bVrmzFZUpDsn/cVikeZkklD0hAhsWoNqgNIxIU1XrAvgTW6
HRK4D2OEC9cuHgW7aqSNloIXMBB974DiEomfInmoMxKdfWn5Ar6IVLzEkExyND93
Zm31HBXFyd54PbUj2Nj+Jk5GSTqHEfXjJojvt0tiYran05fVkr2Zd4WyBT5cUczl
jY7YQtmdhKh/0g+/cQu4IFT3E7Wpp3GTQimEJkgsxoCdFFMazwuttMjRK9e675fn
nFqwTkXmdbTIR+aJzjHIr3CFt+EjtdV0l4xumKyzpnDc10LNxpXYjd4mu+bCEgiK
st+J1NtHWmgxxEZA9F5AkU6LITsZN6zCEk73rYisnJ9cnp3kZr5VOkciT9V+wVv3
WpgqqSMMv69ejzNy1WYpyMlVfrV5tgVhrqPlVw3MId4mCXV5CSlo2j/Jjn15s7+r
l8u7mbuKJrJtaj6wTq4IF3CW0Oho/QklszaVnq1YS4eOea0qsEJh7+bNmoAFszuA
SN+sBNKgs+kNrIqw9nEmAz2q8qXQUasT/OHgzPDkhk5kScMpT6W+y+Si1fMH1eXZ
F/AU31r/Q9SfWgAoGEaska/hYJuMFMAycJDa869J7ktl211QF9EbR+JP3xACbw/9
jeP9gAjPsTtg7gyUACetFHLHF2Cgc4kqS0a0E1QweERilfJRGC1u01gLzTkCNULv
MrA2s3dkDgQtyDmzKL/qVlhTC0ACoSduIn3p4ABrf9kfqyPaXYlSWapZvl5/UQqc
APuNSpNyJ4Ez1KvdeYNgEK/bnrtSF4kQWbSx7Tv67VCjif9kLlUYfT7n5tRopO/s
7tf4XQnGGPHEPl7pHShhnvdcHnBCySPGPAfWJaYiM83py0toE4p+77z/guThopco
Mv9OqjCbzSpV91rdnirD/xD06D6WmhoJxTeja7f5yburJB/pMhhqU4wkoSr5vlIR
scOMXZx9X/jG/uh22l6bgXfZmxU6+FTotgha2pRS6zu+oFBedIFQJ6AQeW5kin2R
OHfyhN7uL8+HWHJrsoEQLmYEhKF6QzVjuI27GaRjyW9pvaQINaBXc86AEIBugRZM
ztPpTMXca+aLCCvtmYTqphcwhxbC5BWZsxj0Dob5Zfn2dQUE7tln401FQIwVy6mm
qj5pdJ/xPeOEOXZUoWaUE5imfQo9mG92I79FpxA3HVyyNoEn/q7kt/Z/tx3NiPlt
+YxNXmj8R0pdzchAehjwrAYL4RT/TLUnF8bSTYNoVT9QsbXEkz71pl/jLT0/IO7Q
RPaJSHhTdoi5IzDDNtCSUyb/Z7Ti/O2TsYDqcc1UNscKqZBeFAJBWoLrjG1aLiYq
E9ndqpLRnx2P9hbDA2QRidGKic8sHA9fR8zbv7lHofVaEoM7FdGXbOlv48DQq0/y
ZoBs8RzwqF+i8kbQtXTwCtrBDYXlijCzvrXsn4HLh5O5j6FHwCC90gAmQFAOMiAG
tNlvPUS3KUPb3V9193XoCfcvuUbHkl383XwNywqPctWG+Fl1wy9mD3JEhlNVQM/u
M9r9+tGiwAYy/YmnDxL92h+DVyVUSwkkavzAEuNivx0DU9m/NuU9eOo5Ca9coU2i
/iyZZbPTbSGGjCJqijDr09BAEbN6yH8Pm1nIlFe3/q2OvXFy1IiwNaf0wEit2PuQ
FAQ+cwcr/zsv18YlGc4O9ioQBgr55uM8dtR2ry4d5WLFJqcryVtzipsN3pGcgGgH
qH8Lv4SLpHib2tz/tEhK1riK2vCZ8713IEjxulxu/5lI+MO7LEBlCionoiKG05PC
3ERFh8TDO/GWsFgd3EV8//EMg7tc6Z9FdZtQVmyRKtLtfUL4RSVya6BFYPiwQ+LN
wZrWQ48a8XA5sFKMH4kvf3ETMA0deUA9m7Bvp2So8i7C0BosXoLFNsBrq6J7xie4
1pEtev4d6ge8hoT9jbk+io2u5leFqPKsn6pBxCvmN+0KkVX48FUHulw0Wu4Rb6Cq
i64hvz7tlRw+1ZYS6dM/NZELZWpRT7GeaRS060xNWld7kdEWiGxc/QL/Xn+x/ebu
Q5spvmtmovzqDPssg8EpJKGwyZoXFZ039KikUnLjjs7FQsU5d7vDTIcddwVITiyG
4Rn11zwNDF8ILzLOeU+y5oKgFFvDTM3iDj4mAZ2Q4xMdhm58no1jVAabtzbgHu2m
dF2sStesz5sETn6IGQVzyjo6VxQMmf/KvFQRWt8vtN2bQ+wyVa2ZT04gpZbh7U9r
HHJtaiwPOsQ/bL3qBGb4ER5rhWLk1X9/HinCdusZazN8huO+5Be96kqcJ+jclzBL
iu0BY4lhlAheucwP4UbGRW6je+ivOzo7IOjPKlBPOyQr/rPPhU60za9oSr4Pz4Gy
KFogRYSg8I5r3/91ssNKjUhg7eu3wQtLodlIUzOsZs6EFj82CpnL2rGzH8hJqRIL
3UcEg9yMm2MLt59MrYQFFVj1EakHL5c5dovuJ8tQxTaJJGqgajfn8RG6A9DgGcK4
1J9PqWYeparsOIcTBFL8muuxYT1+dAmXxJLk9323LaeOsbubllFIUfTkJuLYknse
OFN9alKf2HkNt6vv34DDEiAPgtLePtWjLG2xQHUhijvkfAD2FmXlYnW6zeMtEVV5
+YEc/i5yxsGGbR3b5zlVDq36EcJJnkAzsJfuNIDyCLJIUUhLMHuDJ6dTe1SnvVgW
zxzaTORilg2BkNxIrek25MBeqJvwQkLMKIXTTSsHKr2AFF9UJdoU3KtifGyeXs4u
hs/ASjWnQW73R9rcUe1fUqth9WosSWRk6AFpJBGlbxW4/zcaM3CnCvmSbnyV6YVr
LWrIOpinO2/Z99OHNEAQWLSA0cJPGp/kKWE8OTiOlqvWkPjL2OxfGb3W5vLsn0wB
bAxXuQLsUabj8NDeBaPdr1WDsXisHuk97dLA+Hd6Wr82oyXVlgfihGfVG9y0V2FV
FGT3mm0UEOAX5v+y+6JJvxmWV9fH1XoltYzsljC1TeNjJp3kys69gWcMbTkAEM0H
ns15xO0hmQy/NmdNxzr3qX8XL3/oAD9U8zVYLVUkNawmjxsRIT2XKc+40G5Lib9n
d/9DyRPe3KzN/5DVC8gU89CX84jT59HkH3Z8QSaPIUYZ9ZoCigKqotMAfeqMlUXo
FlXYGLopiObvSYuPs14GcMC+I+22vrw4hQbrlP5ImrnGZUwPJko8fYXRMGEiJnYi
pCWSHAqailRwkmc9J4hEgorjPuE2Ly37QddDYEyOGA2+yp0h5u8f4x5twQojeJcx
y01FGiZCdsJO2+awyYp/PdZt/cYl5eLKP969SMNcNiMhYTWa12PF4GfBzYjESdyb
tfg9Vm1wyGWRMeICILvt9gtrcyZHzO1g/fH2PuZK+5X/KhlmRz7hF1UvsGWwVFWd
FNY2/0IAMR/Iriyok6UR532HYqjtGzAX0jAXLUyg3fzA++z/WzEI3D7NPzJwO6EK
xmldAwv4ROwgq6P27v1lex7vR/+cHWdKlCX/t0IKYmb4wq2HExFH6YZ7F9TkKJyg
c1kklP91PZq2opeZ9DqhFiTtIta2n5OLOgUx4Mr1JumWa+PA7XOLioxccI8SkDs/
cg8k7cJ0DPZqFQDSfd4wnv3BMs/uOA/6uKcwZd1YdPwrGdBcXBQnUUjPkQNs8a3Q
/pMKdmzPbIAX+MevoAfvOZRSSynqlPhrA5c4ik5fXVr0a2Ez/A0qhab94jnqAe6L
Vv7GyMzqRdvYi5XuDukh2Xuor9OVxs/HiwwUYuV6XTvonvodSnkSLvdV86G6dxVc
dRtDgITJjjXJ5JRfvX16zR7dCRV26JbJuOnYe60mAUCZM7bG9wjEVNEz+q/GOlI2
wLyIHpRGoxelTMjNuunuaWK5ntPzZI7WlEztOkxFljaKFb4+MTpspRcgmFr/vyqV
Jj6V1C5eAvuK6tZnk9IgKkvIFXg3nl+z8G2OGoRtqUnnTDdmViamZRddZroHTUnm
3nhoyJSp6D6qlUwsy1JvqtxXnRwJBc8FOuEl1ER2dnpxdELVPiEGIOzyXozDUlFu
9qcK5MYWRilp4WLrNkeRCKhxo1EaRJ5WMOtclBpEw4eb0x7A3/dsiJ1nhVtlvcOa
3kTvDAbl+kwn1xsFwU0dbXL7s/SR9YtpWAnwOmU8CFUdq4I0Wpij5/lsWkps67Q1
S3qcf7l0+Q48JbVD4NhYHd/osdDKCKgKrMZY9obHG9XpvPK0UteBDkn+Aqqg0Urr
wxTVxQFgPONfWyfjx45bmwCwmi7hnQKTGMsChZoXScCU7qWlVB8sukl40tRhlJGC
rUafMyv4L2gd65JQ17aR8HTN2HE/qFp9lzcVZ9QCcsOIApOtdc1NUzqUmVEB0qqi
ITAg5T+mzbK87knxWsLrC3+6sQkoO7HG0T+vU0jYgL3pAiH829F9twezUFb6ulTo
I2Npx+72krI071nZ2DkMCAfq9POdPJIHP5/nq8Zohh+6ipEX3VlPv11uhFj3exqU
4S2STC1xrqECYE/tvFv2tQeNE4tEkLq4CErNdz1yMXS3jkS3ZmL5/CsJUMYz27aP
9dGTdHBW6snKA6DC8rfCBRnD+5LHckV79pAFQ1sTyqvQ648D7aFZ2sj7UDhfheus
sZM9JN4+H9IAE+C3xx2pi0TF0bq0P2kD8U1Leitl3O4MJQVou+eLi1Rc0G9vMKRS
qgHwAf7p0y70GzmSBgixcPBjne5Tj4KgnT9yfytLKyhVV/48CN6c3uZUhJ/MCO1M
V+f4ocqhd2f3NDVTm+5N0FGBM1Y9BjNoD3P827WoPSlPsfSaE9Ggbp5KfR+so8Sz
Su3JIdzZf5tFf8Oc2iAD1S31rFHYAGRnXhUfCTBGP09gpRW2kAVEz4IB8awuzcr1
rvfuGsVvERmgzIAK3MNljtM5Ogum56iJBmU/I7QNqqHWtvv+AICZZJjk6gLjw41S
thsRVS/zHFB/Vm2RH6V6Nuv2i8YkGhMda3LZSb/UbKgVnn2jW/xtTZB7hsfB56Rs
qS8VEV+ouZ0RtCyWHCdW87HzC8Th0y1emFMQ/cz14+qhIlgdqCyPfDJaVRB4TXrW
8kA4EovcLL4K0vFz2H2TagDc7fWg+vbR83LJbXxCge+oAN/G7bUG0u0fkPs92hLF
DKk5MgofG1f560m/5lusPROk9o+YJBE9P/T4tVC1LJ7/vmynSkWd0XoXuFs2gIUL
0SQb0+0ACp4m6o7oiqch6mtM2Z2rxL3pSErtAMnODJu11cqGZmeI7WrgZs2Ky4Ju
8Ui6LqCUhII/IJF+h/aI8W2CjLHcjUzlkTap1a9Ij9hpsB/aSgLAHDAblmeSQVi8
O/jYryApI1UxzFUyRrX/kalfHWPOdUhwdxXEAHbZFIMsFyWIuA4VYVoKmIcmODZy
4MsmMQhF6LuXzTYcTWMZSoBGnV/2FQS7K5b+XMFhiSWTNNHPkOfLuP8jp2Z0t1T3
PQ32qvozZYFfGPipv8fd3/x+y/uoVWqB1FfUNDON9cZphk4neDiUqnOUgecEmANQ
03Z3FwcER+iIlCt6xMvxfI2z76JfNlW19B+OhO7vi3CAMfNnA7u4KWESEzR2MH0t
5ggtiEymnurPBHpZJnkVo/uty4oqC67LcZYvaVMnjeSf1bDV4q0CoXXFwUeqJk5w
qCbypSWgoztEoYt/Ph50G+X13yL5Qoko6fnnjU8NLADXgwcmDiNSLJJyfCeuTYQd
oOrpgoW/6bW/LmS+HtG9JHfYMPDbQ540xMFGmaNN0XYqG3UL6GT+BYj15rZnk7ND
gmLRRT/7eDP9cNJFb0vD99QiSGxxjuR04xelWjQgw97WIoc37sHl9uxsFzRdwOwZ
9A6bW45MbUQBuQvg4KvylMFhLIqq2SFBbLY3k0f2/2AKbRIvGCx9Gp9X3Q1FfJ8L
X2deecZgwCyOn6gFD7WfZ/3S3bjz8B55nMh6kPLU7CMpYliJIrHOR5dcu14U8J0B
B+KB4NosB04OSwHR4feB4ew3PWS8COugKP6jRoKG4Xeqox8HDayJIJ2pt9pm/dQz
dLeXMbL4XZ/Lz/r+F8PwbNVspCoqskkCRhQk51BM5xWSxj3g/nPEcL/3iV5pZz9I
3NwVwN6W1wGtMSIjnW0SETHkLdO4R/SIMZCPcpgq1n+F+nQ4f9pJCwEWXQpdc8fK
3FeM7JyHmkW2bn4fNMxw8aL0IB46fBYvZENfUIOB3fdC8ucwOpUisigzJnRHvpSf
QtiXG2OUb+IL6eTAr0NkF/nLiq5yUOUlh651ytiy8gVup76sQxy3h0VI6RvBceml
VyBzCiUH/EaHJfykNJwiaQmG25S5v7V2mizbz7JSPW2D3CtCqSqPQp44fLCitgMe
k1gbrf0f9LWJR2ibr9+30lS4pWkwTskhByYXx2H2PZ6u96bCwHI3aADdqUtr83WY
2UFdcwdF1/Rf7rZq5UhVpZ4UqQGjIUoFUjcOMVoG26zn4CPoNksh7S4A3qIM6pG4
WHksvJlzPYpHqpw65H5a7hVOXwqILsV1QF4tdFRwRHcslFNk0znUiFP8ntJHzn9n
n6SNrvBrRBBOK/60Z0/DrNtPqa1JsTpZw5sAVU6pkaIT8h33X4k4sbN7QrRmvwvk
gPeev3GNSrpogt2uwTA0JuMpcDDmn+JhwSto90LtIEz2Iu1OMcP4KsBMKeAi2UHd
7+a4JY9eEhu2T5zOmDcZbiyo9gIfC1DsIyexCEI6aagK3ljAsGYylsEe6xdicnrs
gYt86IpyoVLdFyiBH/WnK31hXCGFDkoDxTXAc7/c/j3ZrtmMBqqchBhTdENmRCO9
n8QAjTm5QuPYIHBY/iFpc6dxey7WbpIUWotitYc+tUAzdA7KNUZTkH4IyRooK2pv
5LIsbTSs2JCRF1vtC0thJzp3jTlseUr+05F+NRRQusgiyONXs2XCJ+njfOo/+NAt
nOOn7Gxrogm565gyfmG8SsWSh3MyQyV4gqfZx2WQeA/fJCyd2O+21DlhNkS9+sum
zftwTReEKpbP7DfVGvi6/BzvxP45Bez+bb+GPerUrz4y1nRf7OUr6z0EhLHxTaCt
HY89vEZlbTHBreZd97CLgVx2HTVn0EU5nEwDp528cpjTEDlkZX3TzSCZIJCxw+zy
kKSdT6iqkTTfeUgWgs4c/uvag0AaHIhAPnNJbsolRp+scO7MppfYxgG/ulZGxoWd
itvZPFsvAE+Mqc3LKjmwVFgX69ZjUVqHnfnL26mhNnSEfvPI0Kgw/Ru7er1UBd7S
7PNpUx8nYd7Gmb/8mJvQiEv7JXWM9XqMFk2wXP2c4bUEF1w9OFKBBGqRM4ozaYVe
CXcSaKO5yLc0lID5Ks/zYXor6SjVd+ClIu2FBa9m0L0NxEvkCS1YXBkt0zrjbNwN
k6KX18NRxBkVJ39Muz+4grNL8gCjnAl4wmu/clnJ/a6DujLgspdZqydH43kieLEv
39VX5Vpw6P4iA5NP9DLBfJvIl0GVu/Ed/VqS1WwqvD0adcVBp60FItQxHrdTnRIb
jDhCBT8Xm8nZLV/hJEvTGQAzNUMcHbE5VIrZtoUWlocwVV7+aMSZKFgIXQkk66uE
lda1auZFN82BoUfUetGNMuZu0rc0SV12k7p/OgAnQ2imR3Ms4abtWPKbPm3p0i++
bl0hahzkV63WB7KTb5Rb5I3pAYYUihRH8zI8VyqcrPurvA+hGv967Gb09zUDa84x
RA2MdRlxmIGhe2Rzgbz/0BYV8lDuiNw+9A9g4x49o7oWmgIDOLkIwXbLRxNCM+7v
kcQ2ZESpBLKFFGHzt7cc1+hViPtNUiNdyy2TDEzREsZZY8Rl3P7wT5ymhxYT7QMH
aSyELidIu8XtIJxuSxBv9OLbQNNRypE+PVJSup8pl0dDH1uanz6dgC05jt14kceE
li/JIl3xaYZCnq3ADMGzddIX//mVnpBSqpa80twxPn9ZBDFSXA0A1+i0aKnSvqfG
srnNLw25DY4koke+WpZ72/5DDQOulKeTiC9Wa9zxLERx+ZDNwQ/Q5qf4Ne9AH3Cx
9B7eSDDfK5zmCdqn67xIPoxEZ9f57FB/xhDW0hmZKkl8hsVkMwHk3OCBQdaHtcQe
tdUGmEh61ZvVmxm8GgvaMrHwEKoJ8iATUG1enkF+b8G9i/6F0p7mB+FL9T4zZFQH
dnmHZzYRWn9sysmYjwlP4q+d/tBziaq7zoT/p6nJ1Fx6vW58CsUAQdajZNhMJF9F
GltF+vxRdffpT8clIgnBVgqVRQed/mlqIGCCElFJr/2GjyS87yU14Oi7primaxTV
REjVa/Y0hfO9E6TAhTVK3d18dJovstHs9GzHpUlizPDtgx3hPFutDSr71bDfBNeh
QEA3DpvzNHUJHxJGbIrusirLoZpUix2WaArejVUHOLmbT+8v9Mbat7KeL1pnxj4N
r1zezKYI8ffhXQekdhOLSeCpeprPIyWkg3laWb1JE0brRQ1mV+nzjCcTmJqYfpvw
+dwppFLmcMClB5TQ0XIEEgcllWT5ZzMn6GDWSzXtLdm0PUcym/X8mxhfo6+SCEXI
HWm+0nPCXB+OaNcGVW7xK/HSNmhAPi1uaif9nxJLmgPY3DoGLLUlcrMiFE2QyR3Y
xTUyYusPCJlNbZtXInEG6nRY2Mm+ViC+zIWiWTLAk6AyvUhGsXBGykAJmyzF8lC/
5r9SkwwpUmBQ99Q1hXQ07Y9zYUnslIQiyuaeGJIJzZNnyxgxxKQIeppZXNUuBL2Z
IrWyNsETIghCpzOTRhXqiqk8ncCs95HZUqeQNzgBS5EotOtet54/+W7IMNX7SxkL
fZZnyIS459JwE3uFaNF2uou3fu+0/DPC2kcRjKphKKx5tQSj8eRhsUtrEK+AqkZw
1mKd/+duqWfklAl9/y3HF56uWUe7u23MUB4DyFxzDhf40Pf1NN9zR1LWK9YG7njL
cwr6CENu/7fpP2MNiVhCLpD3PTEPwc+F+OuffWGsP+hewCWNzUZMEW3wUaQwyunw
YqBYIXDhp5B0Z8z5JUxgD4tWvbyiyDNiSa6YTTqPKxKya/qU4Lam1iEBp+0eIo3c
suvi58k/Cbn+cxVVLGqjU8sTWVcXnUd4pa/ugaMvAvDPhP2jnnPkTIGPOSW4W4ZA
Qwc5SFcIRVz3NU05C1X2xMTzXabbHFaHX99HAzrtO7GjBFqLC0jt7OYVD7mdInlG
AQieaGauO4WHklDKDhfYz/pZl+YJ+nsCAaYB41MdqSpYEF6PKJdUpEl2w7s7esZd
WRpno36p6oLG0rv0p6H/sbQ8uYBNjH4t8ycI+v32J0l6NcoitVsJkOkgfYUKvyzT
iQ4ztPg4oEsroIegpHdivIaZItU4yha/1nRj2N2/wODJFj2lxNDr0JcFzRAFKR87
KJcvSBhchr7pU5C4lXUvl0XPX4nFrkSIQxgfH5MDITWhPJkDNph7f4l0tr48fOHv
esH4lF6IBV5sj5h55C3BHbnhtjF+Ij4jfJ44YVu3xHzSB+cB5nJDoA9sSnhl+8zb
fI9DT9hZ+TpLoNNDyknnzPNARVq56WkCH7TLnabWRydKYJlnHBVU+1HSF6QoRZ7y
yfQCOKOcLHaSZtTtuAm7bHzP9I0sllz/DLDmaO/zusdtpj3ElGTrBs2v/YPn3l0t
ZUuXjCSz90DnW7mzUEc+jMzeEQSWhHQTVdAYYlnP2yhMQjVgkAYRlSqhXJQVEVpd
PCCXDfXeV5r5Vf1ry74YQkBBYN2zldRjXWAHdhpq7uWmBE/AzP9zaoEa/YipWRk4
dZoDU33PpohxH5XahedNpiXqDlRyr70qby2/hU0lqUUxtiBpsNMGiNYcedL5VcgZ
fJPM3MWZR2EZ0ynyKdMyBH5FP9i6LGAhQRHGJL9VnaKBfDgrsXp5f36FQmZJ7pNL
h0aVMYIfdHFH3bEYtSMCLVr2n6B2dYE9+VnUxhwg+42s9RtTArJk/L8P6L3VZzvV
NcT4LD1mbo6wf8yFBcD1mQetTywy9xgbl7Xk2ugVYQ4h8oLkFcGlkuOhNoIZc1NN
1WPwNJ9GhHiJdjhNucrQA3SGgK44UVRefO2yHnVa//MOLGVTiWUnpH6Rxdmel7PL
H8zRTB0lGarrCR51gXib4Ztc1N/b1RxK1aNnxLlmNCYlPcoOXxianz8UncfzWpYr
lwdeB9MS4uF48iL+XhvNchbMGszVCrutZzYUs3r8NmSJLi3kn8pa8B4E1fQ4NqdB
z0nDEzzTdeAZH46eanLqJAN8HnCG+Qwblic6SEDSduIXnGy+fsII4m0oHKH8OggA
Q2qhF02lxAslIwhSZarqF0VWroL0kLQSVEk8zGxMFrhDUCcWV0gbCVx/INVXa7b6
v8GDqTHAXGAiyg7StcnzsSOxcdTzShVGCzBCZU31z6sR0bQHOmODn5zN5u67rzT3
7YKwqXBln+WRPsc/wWGsdbTky+7WkKHrLisVim+tVQsgErBKwOvYfXGWn2YKnrgk
RC/TPbkBbtzUbr1N187E5oOQytMoNRAkFmrozp/dj90dgqhRKUgOb5Sh+HOUDwZy
0OwjFRxCGpkwX7AV6W1OcV/wPPQl3mHir8sievLBqumBCd436WqDEVzpuzQP92AP
1N0Om9VbUHpAn3LqZ9TBNy4SLnyA7qiFTqmUQv9ziP9fwinNoyvUNGhHW5m/xeAE
qn1aZFEXpv+TUq0/gUETqMgxFdUV6zBM6b+0LQnChTzI3BHaIcyV5b6jAKYjem2l
WjB30y3IFXJUrHf9KNE6yNL9UQHy+r2tTU0wnvRO8vcBO11LO59P/50IbGvgdU0D
VL+oCVgQeN30aRXAle4/7JEDMj+HI0JanHn10nrggZfaBDdkpTVCrj3OTSw4GO3c
b20Yqlyrj4s5e7iCTo/ROdx6AyKMns3dsTty321e7PJ7eA1URzSlUcbABYHyQ3X9
1AXGJbtJpj78ru6L1QCqWFy2g2c3cdHJp7iApKS9C9q4cZE4qqLpBH1oRHD+NWi+
5COtmKEY8tyhlcprEMNi3uLLYcGCg8avNsUjP0cPut6i25NtI0YeiHw9qqZnyszL
gTLRdIzzhunvS4ycdZxQimRG/41NBllhmnxaXU9QiUDuI61ytjZXilGlW6U6CgfL
hs2inQyLqIYJd7pbKa6TUi7Wn/gbPSjsTOi35V7cpNXS/D0a82b7afs5GJl8ypeG
BJSFKuONryOnPVGl3K6ghUydLgPwqHzl/irR+68gXmZTvhelujO6A3iuXsr3xcvT
/gbnhoScMn7T3GDqqjK0NvPmQJn9rXA4HhQ/PF/HuzCaJj9vvb6bdQfFsKi/t+VA
4PYx15ScxAhFWQXg/cj1T0PSwOpcS8Sr8G2WQBKgWdQ10KDWfOweclmZjN/tUJeW
GXYkQtIAG0+eyZBnWzLAY5RLLnxD663sDtF4Lu9pPL6MipiQ9WgcwWlTtIQSUyEL
T6G9tTtZQxZWR3L+IUA4kc+R+h3jTQ8RzpEV5vSJQI1SqbQAeiyFZdLReEx5bKn+
WtpJcjKaBUoFwZ0qq7dcUzW9Nh0wAmX5N4kYhDe7EPKFO0vuaiQDLXFAgnKFEL3/
ij/+nZKKa6djGCrYHVDnVvHwA0ChfNhu1Zn04f+xBWxbatIjl5mBTAOmFWd8OhNX
svm5y2UQoWFZ+oU+C+r1QEqK3G4w+oQPOCgWr2vO64wVA9Wx10Zdl2MJ1HS837zr
wCWbK75x7/BD3q3dCIkaLm+Yv+V6Ci0NISbMa+dH8erLObYrytHgrCLCfMndPkVQ
lSzG82se0WBTuYMN7KxgWF92pLkEY4lia7hQOke5gNVZn3UaEOwQh+0yUKVujl6X
zAYPZY+M5Qlq35XA+Ua8/f96S4zID1E1peqB9WK6k5GdcIc44BEKkz2lE8hSEOqm
GoNAqZrt2iSOihxTQiw1upVODtZKa7RMyAFHxWYoz2EyUsDZoM2pAaVj61ujg6gC
YLy9QbuCKe7+KJhgMUd+g1bi3gsLHUQ4Ol7bluLXL++3XDv3uTgyA4MA8Lz+fDm9
HtcZJwXIUSUH3SycVW53TuhBQkdHHoQpFZU7tRtmE8YThKC5GAd14pYRmkCFfiOr
kMEkD++C0lmP/6Y1kAzswxver/Kk9F2Y5IBzCksfBronptL0FR3zFwmgOX9vsOLP
eHpNTZmRWWq54wCzqkDZ4DVWk7S+J3ksLEEYbLyc5sSM703RfxG29jS+DIy0g6sn
SD6zIu1Rz2e3260fjP60Dk798vExbt6th4+u9xik3q3rFznMvi/11zOr8GMYWohk
RhWvvEk05YpG9R/RTYUZBlrwOcvCMd2tu7EDFXNRQCgi7qqsOB3KBxiOOwWTJNOy
wW4VKA+kwD3eEXL/N8nw83wExXCZgYTMVPPA+mrINP2CIpRym1kmcxsjqsJ1lW9D
wEDrTs3haP50keBewqykjmRBo+SePp0k8Hh1DpulfL1QnfDc1M1VZWLk6GGG251Y
G63xYeWcW9AJhh1segaL0Zha04Ccb65ac6/DfIpO4l+2HFu5ljP1OGOtNZaVPZIl
XMXX8WEEJ85eRAkrtDvKY+vf9ZB5Z05WGOyj6/PvAz5mAttYWjrOg1hLbCUqkuu/
63Ovg1vWihd+vM7i1uoLRfke4zwbOdmeutSmawuFAmjooAltFPzgk6RvAS8UPHBA
Bc8Kpj59L2YKqrQJWijOt8bBY9BOVOKPdK1jYsb42sC/bYu2btGmRJK5xCCUwoDz
8OObnroUvmfr31yKJr7bkeC35Mxb9pHhPplLagAGLLHlLrEDu4MlcOAAhQcZ5rDM
5yVM97mM+Ghbt8rz7kjfFwqTbg7ap8WB8K2Xu7twJJSBp9cxbzxGTJEJCSDDmN9Q
eh7aXzIXGZXxM1RhYKHj3KPeqBz0guF5PyhZYJNxh9Sk0AtXxOUoljVqxVKGk5Ww
87j37G6l0gJUv+ss1AC9saRTz1vZFUdz8bQwPbFSDL9+28u/zL2VFJK9uncubm1q
tpmcF+NBsGLyBHjeF7vsx3Rn1ic+y3LZ1QqgpaVY8YVNZ8V2u++bgEte+KA3eW2m
o//qV3GHaH1V2mo5V7Ud++cVF1wzJMZbwv4qyNuZYqMIhQ2kMN47lS/hUc7pZkW4
fPY886mcWePUfa2pUFwCICNfb6jJBy2509fpAII8cOV+37GO+dcSjQU99toA5dZ5
Acj8JcpYpflQnq5B4f4Rto18Vsq5ijSPbG6UPrREK6npfwMHvcsI0LfPbPXD6rS8
8p8/vPqJNGz0ruiqEgVOSwBdOFPZNo9IiiqSxyXdWK9vpF8hr18AOTQECs7BuukR
5ueXbWby3O15GOYVPQZJZPudWNhfoYqO7JNrL1vv3utADvJPTUXKfcbJ53R1iCMV
Nru1C46TUK3V+9CfX1UyURy7r1usFQAouKVHsayo/KILClxp79AQETqp7YhLUYKy
c/zyjGpTVIVPuWfhzcWpVKW9UiPsopFxz8y5S2Ko2n/bcefu0YqcX4K2ee3unDPT
LZurC3qUQWMQIbENem2ptYzTOs8zSOIx/SruTuTAoapzurZJb9P5hSY+3vP33+ai
XN4XxFO1yOXrmeiBj8PAC+6OiMaz1zAbKCbw3EsQztKPrVr1bsM9CLxUmQElEoDo
zorMF9MgeYIXm39KzATD0iFBIZE+5DqrERo0Qg6Z4/nNeIB7RwE9lwJgBH0GelMK
JOg4oKppBs+fegZNgT4y+sPDAP5RI3k6GLHZFojrOEf8Cjoczj3gv2hIatZh4mbY
FfA2U9B3/0Yw7tlVPkAXVa1X9M2lnnGFTUchts2tIDeHtORVA90FOkXCCkKA+mJs
m80GPWQdfqwYg+As6iD0Ge6Ni2Hzm7bVzrwQdb2sWGh9at1QfzIa1fajFChyuHDo
Sw81NBrVFKhaJjVvsvXrreyflIZGwSdd0iNnmgoXttHlxaNhcx3WVDpP2sLIfLQ2
jrJ6hO+eSL/sur9MNe/W2FOcb3T6Nc5DnfAB/qaHNO18dURDBlNPC2maNaU6ggDN
FVdEdx+YIzYRjBQWjIxO+zgr7rANHOWAEUsL4DFoU4jESt/3L1G3jMLNl4apaM5h
l5RYeDoHtRhCs0fHKbC9+WRj8aGEwmk3IMC+B1psYUgMvn/nDggJh64LBcAL1RQs
BdGxAtpRwjg08cXqcZStAzAkP7o5R0XwWZR9sXQsqOoxv2bHSJ9miKQgXE9r8EC6
J7evdC6i7+CFHNdvNiqXz1/ybzJJKhZe8CweJAzNPa25LdPB/ItkVu4/GTEPW1/I
5IDYMHfrUXtFNwiHygADNYV8YdCb7yb9vJT3+0LLW5bHRSGMYJes6FKtanJ0Q6cg
bdV0HvZ5bW/6ml6G6piSRdzjEE62lIRTzM760Bi0mZ72PhUZDRCy64e6ec99ZSct
ASAVHq6woKlhT21tv42ENuMzAEn7mAVy6SgJugcHgw0QngnWw6VR/Nd955tAvAYy
BYf8GBaBC68oHKyPhIENQIbYeJ5UOldWa2fARnsnnreU0RhemlMFkJrlF1LFI3bJ
n2C987WGM6c4YkVTjaLlShAVOoofVFz77pWxxmjfScBr+JPj/mpkxd9mKN2KvSJ4
AjiMcEeJdEQXM1dE23d5gA+sDV3gTcyAGEB1XHCOYiaDs4OHwke5qxstqzm5aC3N
LThs0PuCeXAH1Y3aAAoba2IJTZbvAW1lk6TF1XUPm7j3MTxHMAabdC7gpagw/8r0
k9HBnJ/EmwsCMUB/ZtbRcc9iFZNMrR18IjeQfXrZC4M5P0DQnDYTt4DSfXG/VnY5
Sl3qLGbnNw52YJITmNBKqIB/aOTglbFXeD6AJGs4AgCTnp2622U/DE4xCOE2So9S
44phXD/8LzmetyAQLdu/Xv34COmZJBwLzVMFdBEqqWTGyztpnTUBF8Xlm/XqVZdG
h6EqM5IZY1uano9iEV0xMynd0UxsVd7b3quhyew+o52+3p059rMkFDMkWF/hcaaw
mCRKTUoraSa9WC9JpBFDGcFBaBq7PTTw/FruGHJ0nOW26TkjnxzcVLBM/0pHlb/r
pSbRbB4J1KtVoyGFXL05XXLztr3QcgaqQDJygScGxnxrIKB8Inr3icN8ZeLUKOra
0OgngQK7Nlj0RI6JEgeuFxBG1D8mpEbNzLU6YtzB0Civimq1wcq76lWQJ9mM3PVh
A3WAmyJuLM0R6JCGK0lrJwXlyT26yLPl1EWITZPSTV6tdzySZlmKeOQdtI9VrRU9
4q5LFUBre7Wk4ForxjZeHwjpXS/ORpb5zmUooh87EpVpAFpvzK/6ePA49EiElB4a
na71rmTUU3sc4w6z+PVjZQ0oO0iMBQrkEP7nzMPB8F0sHbKT6dXVsgTF5kXrfZSa
kYUr/hiVRM6SyRM211OHqMmaVeSPNEJ85cXbhG0PtvcH3rO29gyzF6XZxk5lfEsC
zY1Fo83nE0x5wbNpo32de/iRyNVkhwETP7hYRH2T8a6Phveclhq1y7xIRMByRHaq
uqtj+J8YR7G1brrtKjmx2f1DUdlJ4JGfJvZvRFXhZp0v/e3xqRwvIcR0apnYntxc
ukdyNAGYu9psjkflZYugu/COvDQ8kQa592FsLUwkV5sAx3RoNYinKHKk7ZmDWwXB
0g0TrjSXw/tX/Go7xe4HxRI1tMoPrt43RH6rv7RAGIQiGKSSr19OQexowiey0y+J
5kmZ8YgNLvWjPzvqz+3jkPFpY3lq9+9GSFn69d/GtE5VXxVHYiIYrqZuVNTUrUji
thcx7XRqHDUFQQeg8KP9WdEQRAdob7em6URnn4ssg7rWuJEgLGnKKinCoFv5pkfu
At1GDOznjmEOpjaMiwfltYVe2C0mr4cPDxD1QmAuBm1V5yqGogJhWjZd2JsA2+JN
eqWg3inOW1qdQNnD8QqOttQkg2miT5nQBnPoT8GMw4Ji5V400xf5SQbKWzGD3GT8
/vcLOUeGw5ZTrDT5BgxnS+MX8oca2+dvBROi/NC/wM1G9de7P1gaqYL77JfccU98
DTi1L06dtLJqHEJgD1dRkPeW7HadWbwGmOGYDPuucj/9mY74wh+ryO5PfXnq5iPH
mrw3q30EnXg8TOxsANBA2zifCQvpzcZVZ8Zq+6LAmGA6RBD1AYxA1UBoBBiq98e9
4Bk/jl2VJk5mqH93XWqWAKXqJr7AxL7UT/YaOi5yjZNGUEu7ZcM3DKGgszvdGCwN
aoDzkkyTpaF9ZMk81zdtQNUkDiHBKBE+lJTtMN5hWzh5duUfYYCNJb/Wh+cBIlwj
pSjje4ed+207m34sFZmmxYb+5Lhu6BuR7luI+1z+6IQxn5eOb9Qn56vZwq+8WxdL
p9ZUAGtOYaYQSt3EJNyP7GHm0bvWcbIxape11DQbEP97N5YAoTufI1Az2BInaJuv
JdPHUgDPLvFLXPHJAdzmjoQm+7MrIqdjffsN+7VZIMy4iZu35H3ALttemwBxnoMB
/x4jSRTt+SPZjguCl//adnASBZY1NLW8mf7GQTbVNJV6eF6FmzIfTDHHVFB/uVfp
q4LE480LNcpGz3X0GBPFgHok5LD++hQ09oF/FFEy7gNIp6+cQlBmfAP2u7adIvFa
SZpDdbZEo/U9is/SFWOn6v2QkgCfB8fZHNnu9E6MD2L4xp+i2mFJCJemq+fNib8t
IkU2MNzDsdahbfAXdbczKInx9YdnnKNBJvd6kK3/TM+x/AatYxgkGAecI+C4Rfze
Dz2vau1Qdz0qbWaVhFRHmKAvmrHAvKC51HHMdYsYSn+8D3O05AWDGmZrYYi9LxL4
f2mn0H1+fpKRYDEEaZzyZi1QyXaq4u7irlZy1iHH9RYUo6vCkS8RchduvBeAm2zA
Dri+yZr86dWG1Np2UrbDWoKAKJj4ZdS23VyGXvI7QAutvh8FHe2Vg1QJxfPxn6ft
DfxYFhUqRuGMWwncQW8nnZ8INJDWLMOMA5tgTHR2GlcUOdBzUvXHJuDh8dp/a+gK
xgfmmOUAwyvyy22lJ9O2z2eAEAjGqzkeqItqXQrPkgeldfkhQbqVuzcnawBlwl2d
+CX0PBq4UITUN98CBnm6R/Dd4kxaytdFmJocphaReSCQ5tJ7Zc2W7hpJqfCqoJJQ
WeP76pW55TuJz6BDgfN4P5FnaQAOaSOWvcvMsH5qvahB5wEgWpKvLAg5zOHXly8f
9r5w32TKhASbdG47jzFXAw715xff2QUQEh+rD1lapQWJFaBH7NBR/hoC3gGMXXhZ
MjDrcrc/DWAg4Rb0PtAMIctPfg5mf4q3pjCFNPRMZJ6k0Dj5isq4Fe+JjXQVZRTn
Cu2ISk8KyZlF0DUBcIgQYzJmOis3YHD/kdQIxGJjtSvg9j7LGQnUFZkI1q1DmV43
WMBqSVU0sAbX2TOFl3Ke+XStl0eMZSZ7Khsh0CZBHvHRFxdd3XI4bWN5brREbAWV
8xdZ7PEClNphCeALPh2j0EdwctPeec+SxHRsyCUM9QQlKgLFi8Qwbn8xR9fdQwDP
0uiTJ4emWrwInguKhh963+5a/EfVYmlOdx5SdkX/pe07yfRE2koVA7zAuBS8S93A
HLmz1eN+EnxNQyMhEJ+pE/lC+1vNM4mDj7m40WLmITU1j1ON4gpG+XvP45N9FhmF
Gf2xQgFDihOekewvUCgO3uiO3R+QKxxiE/vtkblrm/6u1jykesjHmOp+Cztw5Ndh
d4+HVyrLilS3vkT/xlPPLV5o5BIrMN2m/HtTHUua3DcvT5qu53eXs6BF8FNjVlHl
XeZPC7VsQOga4ssZIZmlHxhVddX3SltBFA4w6t+XQVr+xMIjx2I0cHEq8yY03+R3
09V4Z065Nzq6ui1HEURLSabwZokPrjeKFlnybtdoZ9HjQIJLteIAZXNgIbw5Ye1Z
rtj8GGUC66C9COxOJxSDPUl2+BrYFFCgB6FTsAxVL/b+AQza9pfoNuh7qe3kHkcf
9p+1AuU+6arxGJXgm0LFTPgpA3BEIHx3q3OLbi17J/lYpkiOSkOckdEOzwV7e6DV
y7Y6vKhLz41t4GOGKaU8U84WlU0aXN0Hza5u4gH/0ZUTJVQff2W2943ahhM17H2R
LajUEAitNgeJEv0ttY4dTRFmGbpTlo6aDlTXfSM6MQbvMooiiWxxIJ4xypsAQwQr
KjhHhDzXRkaPggaEdH8RYM1H3hTSK+k+1efg7hq+SWHukWh+DhK24rSAWtbj7dZz
Mxpy16ARO6OQoO9+g65D7FN/U9zgO82c2gPHgxz5pfr1y275SvJfbOCi0u3LRZyi
nzSDgWNSiHjY/eN1cHD7vbZOIE1ZLqIxZsGskb9MbUnhkTQy7TgC0T0I5il1N9Ab
iZ6DsA7uoGycnfmEFjK5iv7F+/awDcJCFd/ig6nN8kKVcGz6nb6b/rMn1fQp3nn8
Fsq7+RH/ErSTcia9p09VOmLp1IfgzdeIWvnyk7L01udzYVvnmm+i2x/sLxFpF033
pfGO0762rbLFl0N6MvhnJB7Ft/qZ6QabCfc2nHHSUBD8b4Ei5aeEueeLK3R1AdS2
qlLVLM8dhsxVNexuwrNr6Nt/J55erVmHHPRZTy65cqpbghd+DtO6xvswcYpzy9Nv
nRO3D4+81UXekbmDRWJRgGQ04xeJREo7MuOm44mpQAvz8lcfjRZaz16giJ38wpLk
4nqhTLOamDeBrveFwhE8Hr8A8uX3o2a7swgrmHq06E6IkbIs6CP4Ycvi4/99wYdz
IKF6zOylO8uG4RArF9h4gAx4QOLYmYO5C8fY1/6gDnvcmuzjjuFFWq0ts3xZznmT
DiA0B8I6agegmjp/RJ4sIIfeo5B1vBOkHH2OJnxdyCXWqNtpfzWmTqxbVsxNOBUY
reFxhRtmpJ2JNlVz5gFuEXsYZyWQijYxlRShA90LWuwsA4ZxePtvyiVcrMkNBMr7
6Q8ikrpg3C22aMBO0znQJe5yKFhgX7HXp+0X6wQ4BOpvZEiRGbB5k9QzIYXfWngE
px2KHLPeEwxcjetFUXB7hP06I5nizFU4QgK6iweM+uGIYPVJ5hQXnvZshwzwxYRZ
2xlkl8NZ5fTE7udA+1gLArLurqodoZ5eHuPc1gfCr0b8V1G2jChl7qC1eweNwRL5
4Vppym/iaJFYwea9L5e3TwjEzEFTKFR/Qph0GK/hV7tvr0iJ4V9+Cg4XSqAxLrs2
mLT/SPpQGM9nKJjSN4WXC4J1SxiOC0ddVWTH+52A9Rev3ARwXi1X0L4odMgvOKr4
xJaNAP2iDETxCkQEEFH4obKGuSqLMxvFWmBijHbyw1NqCfdyiMoYi0qSrK7fXkCr
rNqkXK0i/s2ZtQzsdDy4AwIUFGWxPpzzKbute6muhZ+uGu8W0Al0cJdXU0YQ0ZWD
orzSQE94+BB/bb+u+poOGE8LbdkDRBc2cEASAHNSErJ5i8uWcCiqbKF/yaDUQjt0
95BS2HWrZMyrXjS5okheqvAe5dts5G5ZtX2GaVlUZcTmhcReDtYfYKJELwz1A3O5
i58IpAyVGGnPR27PKVo78OfR42at7lUjCilh0plCefFHI50TRg3L9fwcj7nbz03r
AJA5WgmdyBzl05iUnJAL25qKL2IFeMfbUKFunORJBck3gS3lF5hh/TZUKMBFNzze
g+gJ4KiPkjDM+ww771GN8Ijwmjc2yafMSaULfU26XC7awGTQTLM4SUUkAUiZhOzu
mC+Dhg/KAqXOyBrct7EjXOikc28F1ON6DFdgWoYjoxEtHotQj6JUn363PkZnCp4r
SQntybrcS3ix7FXhwZfw2HF934QdcoDSetwDMcokT106hpJKUmcqGYSKK6j2SXIa
Q2pvJdDjX5MnMi4/+BODNuEybx6k08hlsRzGSWkpmyCW8njUpna8sCSJacGX3aYN
FiNf7UarhtsrOfdzl7mrodaGF7RKRho9rh6h3lVHWH/A9ybDfWoc0PfKbiHfSS7d
F5qaPkwszDvC0D8wOO4tr+NwmifN8Z2AVkvLBxIETlg0WzvO9PoWae4U0LOZN+U2
m9H4+3tp+CqNz+UU23h9oBv5GPa+Ft6dZLeH+8XUca9twF5DifM93z98WETczv84
qP5WeLzJBhQzW70je8OmOILm9oG5IJPaYCzbVsqAC+thBFkhehOIAXD8r1vuBk91
i0ZKTbYnawBMPj06j/IKf1Uvbot+JYjBFiunCKSC8JDsN54O9fVIJaCXKr3NZIzJ
RciJsOUDwJ0NxeGMrEzgy57e5wmR/XG4Q7URsaem4aTqZ6KzA4/U7EJKq7cVFFwF
fkK6fw9HA4uwStnaOxCa09QOPiVNylAg2lhhlXLLhq5zAP7DWjyDR5bbi9P8YW4E
65JnL4vfWbu1h4mTTzE2rFV+8wLdZux9ErWqxJRpDvSL5INU0Wow+fZS37AKq3XR
R6b88pkDlq7BimGqpYbwqZLKDb23Huow6brxSzEjTYy4uG7xVen9Z7tm7HQ5kYCo
1hEA/WNlQNC7ABtj3l5V8xmYt1GVFVGhxdNk5Xy4jh3b1F80kSxQHt83GcnwJlhL
WBMHpPKgiRlK4qPGVTwjfkNoDXvT7MiZFm0CTbgFHmpjoow3RwcOwP9pq1k9eafT
YQVR8db4APUu0G7Ko5Cgi9cdjUQKB3JubdoSzDS7DhOE0QUHfOAe6E6n6qWbmg2C
AaErVZ1XsCgxqPrGD1EyTamsWqO13AdPZgMjSm6nB86Ldx6zAG9vwnppiEBv5VzK
+DKrOr29yRIA2FZyCCMnxnz81veDts7qm3YKXaIg+xheuN/ls6wYW4GbzbVGpu3U
lIGajFUqeah6bltrmHu9eBkjM9126dlEfYsY75YLmeu1rLXTLmmMAGhsqIPfV6Xc
520mQRohMMbZpTTu/Kbh7Zy/vuS9EaJ+nm0BjpErWlMdb522CF47g8vJViqkMxvb
2F0aqDVBpkY5llhrmSXdnxl/faKKAJ1HWzdb9DjtrCSGznlVICKLE0ChJkT6/rVD
FtCWsd6SrcYAKzAI5LimLi4CMwuDIJqMRjCI6SazQQTDq5K0QxwZhzz3MMRJURN2
BAODWVcuWrYkHkfU22QMI9Ev8l6twtlK/Cw0tbjwFTFkcRoeGv/SWfblKZ9/BVw5
hFs3ZBYOIqCzl3aXWcZ6tUZm6Tyoc4EKcv4jzSviw7hN9/RRBiVu0m1/hVtbOZNw
ETn3OEuFUGSvK5oyeHdkL9Gih5zprSa8RAfZb/JDau7Q9Z7NKb1NpWnNnGDlbGEW
Jnc8U5aA6tp6E7u3ZLjaWTlVVhzHJIFiC5kbEmG9v9+vHVIqlGNzQi6r3+UdLapC
T8h6SMMe4rE/I74+NUpt4K2ydDUMUCcDT9xLcSKviirOYm61PQ0HHpsiO1d1JIuY
J+ceMM4f10gQNwOE2D+D5N1rOGrHtcXmsiQ/mtmrz6ticVgU79bMUoefr8QQRo1Z
3WrbnDCIDlT2dEj+wAWu8T/7OqEkn8lNFUpmCdTGkaVirES33TLp1GxJnLOwt21u
mNfj6+NdPuIO886z7uqXCONreJF4gdtvScRUjG3ubAEC47895i4ph+f09+JfKyiv
BxxpNUCwzF+f1NBB8mjFsRPu/56YLu5tF0S/D/EhoXI5Hk0kLi6BIG1z13Wzrif3
ra3Nk3BsDYkbTSyo9QpP/z4tt4VceMSLyaWQSBe4ZjnKzPvCBp/NXgu2GgIK05VA
nBQIyNRuzWjAvyJ1G5NBU1VXoZljXsCaMEPS7TygDcNIQxLy5VfhibCIaFijlQoB
DstUkWoBL/TPOdi3cbln74W5EH2NoQU9ObtXJMsXHssiD8SBlxRQ7Ge0QOBJX4u4
Zbk/vKpGOVRlTGeUxeqZT591hIr2v+3/5UYsI3pTaZrH0ZEQRGfdQHW7aRW1JEzM
Qyyvbr3JiWCixpENEWrPOF3RDWQygxjDRt70ilcay1vdQTG6KUruK7GAd7Ot82HQ
n89uiaGituFwahk6vHLM8qA3torBodufvJYwsBMeVqMAEtuX58qWXSEIjUtK98iJ
W4iB2CVo3Dw7uGi1twNABqEreijB+9crWcay3JWY0bMPBm3LVJJfCwVvHdr2UpD2
Z5sEM5CdkLffHOsBJFtVONl6KCrszAZGRyOTX7L33om5IBIh6TZz6GvHfCCyM7QR
F8E5rI6A6SBPW3lwZ+Lt9ykuKMiP0sipglyKbh0wgvY0RGg13FNOepW49+MXP/V7
uR3U/MwyrpIXnZWIGWkUMSZ6EJ9ndiaIJcd2s4uX4ldR89XrSzuYBd33p1XAIF+/
HvsrGJ7bGsbN57UoyaV5tlhtCLZCw9gdakVP9iiI1+zrulzuQZYN8EoAG4II0pk+
2z0nR1DXqUoWysO3gpdd/ZbVUp8V2Y5xycoua0zR+MrsEuCIai6t1HlMYlmznQSy
9WB8OTyXU6ClqDaO57HnmUNzzvU95am7HkG8ES4GTPyfHXnPAF7Uv9/YTRTATJwa
Zm/UhX6YMBAdiYY5yDQxKln/0cdKm6LQ2/m6FtcVDao7d0yFapebikKzmjbq3o8O
+h5jHghnLBGvpnaiDmmrrlgspvdgIYffbI4EB/3b+vf9EwrChEryVHQbxIrj1d6p
0AoDtC6vlXmkGZPsd9CBXg9v7bQhft3vRMHbx+3qoHQS+HOutnEzgaEzxtshCblC
E73+MS7n3k6DDiN1GqIkg+oT538GsGddhjUthytkcaYDCGMxplrtilzMOtf61Hb6
P1BWSBPAg2lGB0TEsJ0twGQbzAK/hJQQTsXgslNvuLn22v3ZhcIBdah0icWrJxpn
r+BfSuG9itXHbxM7ZhPaQNJDtZs50cQXaNMVkNPxSAaJA/yN4rTYmVNacxuVIy2a
qBVknYwLd0MvYQ/IPmLKXzPVG2WG/uDMHdnJ4zSfh2ackAOMWVGgEHWh/PG1104N
MO/UobIRcVe//VUEy92xor7i53qkUeTGfQOlm1//Tw8AD1Vg5TRnIJiByyA7jLF9
MPv5288zzf7S+QvNOvkYC6p+rVz98Q1G6KRyMdnOB7An/X1942PB3cBbOi3ebjuL
0YvobLqnz+fCBxu8nuRCBOJsB0t7qc8nqiGCmm1/qZ1TZvnFeNUiecBCen7v3g7W
jl9Wp5tN/Yn7+RpJmBRGBtX2BuxcsH8D1agc7MspJg5qPH9nI/jY8CToFfdLW8DD
3kaSsD/3fi+RU/ZI6RW5lS3ow30yJ5hjopEyR5HP3h5ac5RZUVz/xuHxw7dgybdp
G0bCIwkLxJ4fL3tLS0OsqHozjLdCMqsZfZbe32s4UYOivbcn7J22scJ7R5ZITkSu
fMbH/kp/ekYld/HjMJpU8qwRUEhcn00MHjDmtj6PE7AqF/WBxnU3QNXmGlHmvb8/
1whooaf2/H2yW4Fi92rH0VoQWCT6m+VYYg/iDoPDgJJ8D0bW4mYfzNbQyFKBujh9
YZvOkeKIRgMjhFwMMupas9hHbnoeL9igGyN+dYtjakqIQTcgBQftmwAv9lJPQVgC
sLLkhfo4wGgyNKwlex5NUnU+BSIvJNf2QRmdQWb7zR5d9F+Z5bcDUQQqQyFigCsv
I7Ku+6Xdo/t6GzlX58PJFO0Z4NCMUCLTv2rSLr8j30Faq9qUbPa3ndHb6D33La6G
TbYQV91GTiM322giUH++Ruj+2Uvt5HIfBdJrsyH+B4SYx/zSrMKLld06IbqV/21g
1XhPjsFlKTKrzonT8SvAcHRMotNMQSbPSMflqTKGqQzjQSH72pqZz1Lsiqu+YSUq
fNL2T/+vJ90YIrXeu2eiF9UqR8VOnqo8TIjswPC3Mf98sbxvH144XxMb1VWqzsWL
S0/2kPI1xXpOPJVIV2Yu52wiNlK7JNTgZT+tZNBS3VGwuA098NCZfd5jgTPD0bxR
vUzNF3fuUhw6OCJJvPErt0ci98U5LT6V97oa7nCqM4gyFGYYxBiY6SFdngi7iCrd
avykxwWcjXeK6kWXabpCyNi28ks0mX0QROsP0pNWekqEyomEBZhG03jbqUHUElQ/
tKsJ8hF3cUoUPL0yJVMW/lu5XoLnWw7ufXYCvgi39BNVYsSElkRKtu8dLzbiArl5
IQyu2mvBhA5rLx+BEPJGFxCBmLFzeVKsA/ojRs+i+CD3O63QS6oRt++Co5gbuu2e
j4+7DOaOxpNH4kPCGYu5djrPcytoRMFxABunfQcoKhPGsD4pJf2/mwRCLwFxOHaJ
KPrXzh+aJ8B3xlzhXXTk/VMZY8FAfa5GiC8Z0vBQoYUU0HRvWbRB4XQBig0MCick
jDPJ0/Y6ZI2hgzP1LkMHABBwNiw4Q0CZwgpdr244uEjtoiN2fyBMv6ZIm0Kf+Wea
QwVF9Uwqfd9y0ZkKhPpmAyylRSPBJ1uDjRpzgS864lq0BTQeneEiVmLV2B0UU2ZR
5UHR4X2AvysS27ozrT26IFZpA/eBw4mPPYOoBCLCVBeVgzVMQ4/58duGjNFRYD3m
1xuWeoXOqlOd+SBxjBUzNX/iFcVjCpy9LsNORXaYbkVUD0vai1fJwHCRLO6y2efe
4gZvqMWzDW8WKuHp6P/liL6O2ja81Ly8tDUuZs6pPQOPxbS7TBTbTM1qcq1ARRGd
vDQ6n6xG7O1KpcSKSCVqeR+BcHDkQWZ3NmWiyNGtK7sMRTZagZnAURl/ZefgsBGL
EIA92SS77ORXav67Lwy/sgernMB3cyFqA9JnU2XHx4vQKMMjiqVQwNqdM4Xhp/GT
fUiTQb4Gwo1cD7g7G4oM/0Tnk9SN04vIcjsUgULcFWtidhsDZABtWSgwA4zrws2c
1qkf0X3giRVWZBU0tZFbu/CTkES/r+nGGS2ECQB/4ULWx4iqL1hNgf8s42IBTCjs
082uylPS4rhagNSy+wMejP4nfe1iGiCYutOePeSy+j8AyCsIIuxLZ7lWBGvPEEoU
IRqxkRVlLjezLvEtCoeRfcyIIPG6M9WVquUmffxigutxpcqF2FLO8N1Z9vcMsXlC
oNb3GA01Vd5lEpHp+Q8LslrG1NOWxhl5TOyNQhwVFojjQ4NBcbqputVe+S61lOTz
OlOP7skS5k4rT4V2BMXezX3GGPIIqXB88mfSz3mLgfZ3cFBqZrnU9dFK343nbNjA
pMJBWvYOWuIws40bBKSAZo3LsXdeJgdt/hEO66RwncSNQ8Nh8TY0HM2oBR77IqPh
VJflKS3ztUs54shGvapHKn0cMHLUfg0eUdE/CCNLE1VL7XMLr5mC5dIeoTUWoqbP
3tNlc0U22rX6CBUiMSHe69QmBEUyufNJezyCC9F9c0CGuDnh21ZsAj0PumChZCtN
j148kv+GNto0EYhzExV6smGZP8SweYPFzRsrGqNE7SWSt2Gd/123J0seXqVmcEa9
2KPX4DNdgK6SjU/63md5Li4uLjw8l7H3yOpyk/oE4yqlNOOeVOUImEAyIfUl2Ymn
SeT10CJZ47k8NWdonRenownxseNgIvJtwb73dOTIRR1NPv2HbvN/AQq9F8uYmz9H
iSs03dIWOFo43hb+6BD4wo/20PN3fyZXrSxd/HrgIc/XIa5WrPg4xl2fxRMET69A
41KmrSftv1EMoucjmX7kyNObxZjoXSU29N59wcPWwr3IwyQaBsJy10vtis1gfP3O
g5+kmOVqAla+cuL/YZxANIQ0gyRXvd1h9GLITRv9IIZiJHGy/b9oGWn8mQiHr22M
RnzSrVMiAzLnfwR1PBnbsmtJ1kqybynhpEhHrVaRA2FOzmPaDjFUyb6qXmUCy+Em
GLZg7U3UFIMFs1pMJGCIVwyI3SW4/2W2/jcm5QSczbl/bH6BmbjQ/qozV5y19y7e
kMUeNVvwmeTBTRpxXu54OUZWHAaKalubkwgUZV6k+/RQSqVRRpm9fjZbzgKTs48A
g3X6p7ZNgFUsUJD65OLKTfsEpmuCjIxgWHJ891jB/ly2N45oeRB+w6bTUleKRGd0
uXT2EFqPgTyMEix8ELGLfieR8URuqyu2Dd7G3sRZRSYG495TBy8nsLT3vYsdcyfw
LXPw8mJ+CqzDvFhDNLQ0Ng94PP9ft1AOzR3lFRoprChZAKLub3VVWjbyQnsSEhm1
j+z3A4hiAlkuuC1EoUXMeroH0Ti0LLWUNpuPlSkovoEBEKvK7MDVVMecYhdphFbn
TNAOo961rbk3w1i8MwaIZHM7HalFcCBzchsknS1Q45jFwCLeXKvJHnaHZ/gort1p
nzms+zeuP7Psk7Pk1pTW0jso2+TJAL6Gk8A4C7foVGf9jsMm3UUgZXkjbJsY5Ckw
nIRG1fgpMQFBjDcwAqbp2f5O9voGgUSpTDfcY3KBz4py0XYqCJ6sRhbIEbOzJKGg
049QoBQ9w3mL/M6pD4J1/le1ixWZ+JApkuFA72jwM1bdGR/XzkAcjerIZPagh5W0
kFPbd0kY69JKecKpMo7aFcx6pJG2kj2bUl9zy9u/DjV4gNmsxgi3p1OQhGxoIsxd
+5TiIPXEEvOMJFTciI1uusuISXmPdpocIv7jwh9AqnINFHjT9pMbToyfFjjcbSfP
bZL4jTfNm3k6Xvh7sWDjAdxFViMoZ+ZLUNWv1oMogy8aOa9fo2j/NekpQS7ATw/c
BwxInskOH59HnWwtsV6NFQSGqnWryzCdVlLroO/qVst2eEYm67/5kb9V4vxqa1Bd
j2jiXdrBBbDkntA/IftfpMAF0Vjp80iHr3ESDFuYNb9dOAJvK4Ugf8h8gIVKQWpj
IE8h5kThXOvcgkpD8qlM5G3visE9etSk34lpmzqs0qh+6Ds4ShFq7uGzxQS6vDif
/9FceO7w/pNH19LqcnW4wU8lmmemaFrElPK7kPfhkI25vWGNS//b1Wi4XBEXnPVr
RUaJHFDwBdsABFYbJEPib8DSCsdV+mQ+DIhCgMi6yHUa6OSY2FqYwqPjKY6ljYJr
/bs3ORg/tgDA+6upmRm4TDFcDnd+MD5E/wwGf0LFF3j5QJHGQdszKtHNRfa+ST+n
blNjXU5yYARQECNBQCrA1Dqtycxz3zqHYX0qL4fu48lOBhCGI0J4gmvCEjxfPS9N
9yOsiZW/9Mfyklk6KnTmHRxNaI/owdY/mijPAQhkMkxvvcPRuYFxXwkY0jj2RIch
8zKHrTMUrE5mFATATqt5rEXSc+Irf16gkd062VKqGJNmQpsrsoWr6dUbDubhJnDq
mpwM9IaN2y9GvHLIU/Unmhruct0lNw9pl2p6IdvgPL5q3Qn46n3nPpTvuqwZsSEX
mM38mVmkZOvRMfDMFc3Xpucr4e5IYrM+1BA0MmPrav/FivSFvx+3vsbWsr9sVIwZ
rHCeCgfCnMUau7mb1bY4szEw3pFw2bQ+6h94w/2KjarBv/zv4Z1ks/OXznTzkm/y
snh+j8atrYl660BjIQLaFgghNPveVlsKMtEVxuqcqdA0290kCeOKyB3jcSmOO5YJ
OrGcuAL6xpSLeQ9U9oZTLPbGSvcjh2IPoDp2eyJClLzdXz121IrFBReCQSFjEe3i
Sn/ZxmF3GoocANUCXpeZfXmtabUFnFGKbVjHTsb/9pd4zzOnrpJy6PaslylltAVW
NZ7tLpItf81pHFKHm4uRqSlD+uAbMl0yljIVFNJcHGuobvpHexNzt31fkBTBgLKc
iON/VBamekFO3xBAUeWHM7jYtUm3oj4jg2Yr7oIQsoOeKIE2zozQobz28fGUxscO
3txNfS/4+yVRzVY5IXColAWxU6JFg/5n6jLrAVpJUAOih4Hc6CViAgbqhYk8DiyE
t0e5Rq5p/y8yMYBPVNVFz78eqELl1SBgwu3ty1NV7j0Vk/h9xayS6dQob8njcvex
7iiXbVtewSqTZH1v+p3ZA0lDfkW2Q1TwEgfvdowoYxCul6yUhdMJKqeoPX53C82T
N/WxdN5GMBoLat3uBafWnDNNwIFDiv3qBMFgwnLecnshgDNoodCQhWWKyMWpb6LB
2NhgFt/5B/EGl0MV+mu9//Ik6LQAB2riyGDnaYFDdm6kIoTZrjNpZ5adii6fAk4f
Fdb6lJGuAALegs2mLdMfVPTkhLQQR+KKVMn1lbzXMFFz2tT0qJk9o6MHy10fzMEb
YXO5hSPDibKYtMMjPRLrMFZqaO9pW9Rvou4elT8K16M+WlAYiQooc7POfdy6r6sx
+BGcyB4FbwwG0/sZ1aig/Dh7Lnv5uz+ESuirQyzTtVRpuTY3xeNyWvn14GoJW1Tp
ugsGU7syRUncU/9M84jggjkcgLk8eOV2JL2zh2Tl26WYmyVmCgYrD16CPvfdJKXf
bV0qewGI6A9p0v82XI4cCFO6OAyX+gjSQDZoa7YhvSdR5vHxcXH+gPYdPpG/ldN0
aW98Ws9szxy3AfIa7FuBGEQ2zNQg931Q7ysXb2nF2bDh5+dRwYeYwbPLD2RQ6FZY
Xkjb0x7jGmMfEM8QVa7ZywdJkAR973uT4RnXoXrCyElQwlYiPibJ9jZZCH9zheQ1
DT/3brcmx/bHwN1BZY+pLyhyWn886VQ3qaqOPTVWBnpbGPZAajiHfGDGJUfwosBj
Try2HWcsCf2bmSkWP1SwHYVOyuHeLzZCHFMFPmaFVj76bxDtpkYAGeEsFOIRP01l
fp+ZN/82sU9RycStj4WwDeNB6Vo8QKcv00erk8MUXJjsFJodvbwHp3d8/+thW2ae
Xl92Obk6QSZiDpuc5QgJzYkfggsMK2jIB/MDNHm9y4e4TY5+fd6oljDnSL1M/8nA
nbl9bKt0A94/6a3BFbK6j4ZiARMbTsriHL09Ra09Kcun79AvKpeaxWxFOHfKcwvM
vjabGAzO360DJszNQXnP1c1Wdp64x8QmxPtcgQ5C1rhW4lgaZbty9ScOBwZm/rPk
v/Ys6ChoGGlI5a8GpG3WSKicEhfss+a1QImFK+QNAgxKF0Hz2RywrIoJrInPy+PI
FqdnxoDKS431eUtLXtsSTcLA/AzKFFo7QRUNjKalhRwShvnE8Z765UOojkCfUTWk
4bqezIlOATcj3aM2l+xS/pRA6BLcKnbCKOhBJiTvuDr8knstMfreZDwLqD47U/Tn
FypiWS8ynzr9GjFnRCQLdBGcURn5ALqnj/9iahu4M3xQuFYIx/leLqAOqrauetgQ
eIqlJqZAgNg15O0HbDK2HgMTCzDKFGZpgCxlT/G1N3LmD0gJ9IQ9/84QBJopjat6
7gmrJwZc0/A5J+w6KfRJnanzWUegrUyKGbszx6HlUnAU0Zad3mW/Dg2mtaLKgaax
WHhcsfNmo55lN/2GNCg/smAYAbmWsynJRw134nQ2jC984TZcuLpKWW5AIKpdl9kH
ao8P0XygO41SwD/TvBvp93FC4xZTku+N5bgcVMkKQEX0t9AIhO3DIk0jZjHXSuBY
DwR2d3PzP6cYtYW6OP4EwLYz3U6EXOCNzXW0fMpPDSi0rXg2SkoV8CX5JGKSlaEj
zqVwWPXPCFw4JS1Et85JTu8wxTdkdFImAyVGI11h3zSWGD7gQgjKBe1BYJm9+wPJ
cuZCRbVb1SfcIGZ0PrwIHwME59QaMaUgqZ8tGFi3vBs74/myyP7t6Fge7Dbbrt/Q
p9Ac3LRyVIUNb1BEqRpoXooDj8Py+tYb1aKGVbFtwBjK47yn1Yi3GGfM3XabbMhr
aGTuLj1upeV7RuOkpcN30oaGlitUd8LWjx6066b5vGZhQnllCOSERNOGGkkqcrck
hViIC9z30Reh/Rs0RK5MZoLeqcmSrSEJARQT09O2ModzAM9a6gFD3Txxv55aRrUc
ahsAhnFEnr3YAF1UhkUCQp2cOhUZXi83NmExtRE8yaQrJwnw+Wpa+SuWj0ckVqR7
wZvFFTeSUy8zhSHg+URZYgWxK4LC4I/ECFpUKKujqDBH/nuFsrm79PjWB9edtsED
wRLKG6HOv2JymTy7SDn2l02KfJtqRsnlFGoVY6KGFQQxEExS8c3EZGRj16kFjjIT
KgAnJZhj6uvGXrljHS0WZ8KW5fQUxCEIyaLqAkk+yrWJaar0vuchcafyZDB1LidS
jWbkXRVuBIqsDQjonMYcNNEUTs0iN2zjFt1i0RgS63ByByzAlf7COFK5Ylii4k7U
mTlLpSu2scSA3Q+ywqusHyJGjcp8F/AMg/J53uEYKbT8gG6S9AMLBuYoEaP/rJpo
sV3t2MSnDRSuFudm/oFpbGjPLTK/lWtzm3v6Cg23i21o0TQfEfHcpHXRHrvo8pcr
2SmZG3GYx2oi/hV4jIffxYDVGmGoIFnCmyxUfVszBv5mghUUjen57xGouS1t9ic7
qayho8LEp2AATZ4D7rwmkR6ucQn5VFtMGR1omHvygvOxgVYWfb0l2+0wFyhTl92J
PNxj69xAR5xq63WDIWc80HZIFS7hJQzMuU58YS2G0yTTDD1SSmC/gGO4sqt2aqpy
lsXOxylW6i4HcHczogyZppCePwhBOudVCwSb8H3NXaUzI3vlk1AxKsg7EZpLicAn
zdh3k+scRQkohOHnbXqeea1CeJXbRHbmzFBGrxyrw0abGjqc4TDsb2tXPLkpPNy2
YXuaTMMim6HrRoy98/KeT/FpQtecAUo8vF22JkJG1LyFQwGC/+9zbZL/lN8jtSeu
197JJuLCUzfGDSpZ6Wj1QxgtDAFiyJykBcTyydbTCmSgbvTaDuyML46vA8gSxfB0
crea5ZoWvwi69gite6TENtImS/3e9XYK5f4FVYeapT6VQsb0BuYYZS40UOzlWKYl
L7FH5rWy810G79x/S/1BANb/zaKHUYsHiC4xDIYBuzVadH9cDN6OVTsmGv8GjMXy
XuQltpoWpA2Ee84TzIXvtW971jMrXskQy3lcdxPisD0SthfOUKz8ntqXWH029VDs
HBE1TWk6xjGTIsadBYsnE09heSyuFVJ48v9CKdVU2KejcumOEWLSW24mQ+RwhyIQ
1YRyYCqxxxGg5uJjg+ppYJVqcTHV/SRRVfwWOB2aKsDLJSiCUG1DNltUFYQRmQNA
DoZ8IDjYDa7u7ztsmckVWbRC87mXUOPVb+5QNVn+9iCYz0RkWncQgMS3q09/Cj/L
6LCUFG8TTEIGjzuZeyIwzIJKHPhCrxRd6WWPwpjUiF88RqaxSu0uNEzZhQeumsfF
xm1D8ZEZVZLIUzsFEqEoij6hFYk/gm+hRBqEKO2TDlUe/Kl2jn2XbNdI7De/roaF
g36zYo9aYkcKC23HgPev/3BB0eCZbEjw11mcziRpmAVO36iuuPCc4urRGdL+f/BH
SZwu/UsUnQVMiQNR365BhI+JEZtPfNJuk3zCu9xikqCcIoJeZHsk0mAUK9OTkUWV
51ledTGjkc38fGrYjVvS7UTHm24QFMK3FiKm055Y+ij12x2UVgB1M5mI3UPMeEq8
UR2LOju+oJJfy+MpO3GszRc+G2T//e/QvburFZD4BSn4SgO0Ao97Vd3V9QMnLpWW
5vv6St5zp+cqY2ncVAZeGzhIoF+RCp3LMqDIRcRs6qwD7GIRvZRXbckLd0VFAPL1
ue6u3F2wQZ8Hp7HecMBbE6n1kaMSxpALbY6UaJfdvkuWBhS9Z+kqahU6o+agB9hs
RQm3r8ZdBqAMbY/ARrVfNvkPu6hh4D7r8g6k5eHJqDl7xfmmBXxY5JeS5h7d64b7
8qaF/CDFoRIYJq6wpGCClaSq1GCtQ+RZGlOciwPuoXcMsCzHZOuEm7fVuee9+Js2
Wk9aM7rT/+TlmUc0kL1GO/ykRYi/EZcVAB0FlTUZNjv+fM7jn/G7eAOtDB1E49dq
hKep7qUo2SOuityc2mqotv31cAhr0dfzBADz7rqetdcDWX02CkE9JcRcAuQeBr1b
KvlLSRJdCaR7W47SHS9nAvMkqGMUC7Efep+bdXJDlQSr42wjCWdAwTuRgxJkDevE
gJShQNIDLyUFThkN57oahYKkyUA69vhRjftjaWCx4ZTYfo62rGuzrKqquJCmMA0c
h5x2ZAZBg0P95WIQm9WHemYU8dBnS0xpxBUFWSBEqBXzNZkFCe2Pv0iIgTUUlGUj
qLSLwCP/J4S4lkOu/+yG3DdHKwCbrWf80tAuvgZJKHWoHAMmoJJ2WW0rcXE1AxJX
szeXPfVPRR7Jf1rcFkZo/YIWzuPn2ZcxGv0llctVlnuYYl1/KBgssEmlv290a1ZC
3AVk68ucaxRDR2oPV5FXpyANdaMwwcIep3bumLbwJBEU8D3qtzHzMJMWXYLORL8g
DROchfDyqVkkES/s6vdxUA1jSviWhw2k9uWvzS+lQdJZuSSgIIf2ptrdyiFASAlF
LAdVhtpv5t13HN0dLYFjmjERL3bVAfv7kvOFLvi0B5qPHH9gLWW4WiQdGFo9uMYW
dsv4542DQcWlkCjE2J/krZ/Wx/ebLFkRAsPXGpJ79wGg/cZyCSOh72lOdy3zU/2i
h1p5uILY1ImQWf9xUr4CUR35Bl2p3Wp5lat05q5UodrbaT1caPhnMJ0G5LlWqgoY
rhAlJfjjoajbaKwYKiA33wD7Q3bIZfcYzkpZtUZPpJR4g/yNDIOYl6AIp75ACaBs
OZgHEx4GjZ3n9sgTs52UWjAPtxOLhoJ5UAbSZHbtQCKjf7ZcAZpdAMWcwNytJHUH
xiQTkOR3aoxrZK3bjFZSJ8CeYnxr5pbouCU8MaLPUrWZLdVp+3uPPywUuYcNazsA
I/4bip+1G5d7q9pk3vgQsnCblS3PlERJU8AAUV+WECJHxsTQcZT/2mjRErnMKxNn
+rw4jomuC/PqwXD0i4PKqnbw1WZf1eaIkSFQ0yYFkv/QhuQWA3lkxhl7nWV8iug6
YO3Srs7bkRQpa3CeIGKl1hxvssNvBEIb6mgIwvJ5L5L+vGs1ZhJbW8wdheUHVQLL
IJdb2xj9HbWAzizTDUpcHf2nyCPGRCbVLx/7OxZ6DJRC1NE0JZI9BWBkfhF8nTAw
1jrClRAFnaxx/Z7kvQvvckelJx3qjKNwh4X5T09ZesYl8RK4WyvG7hXBJm8zIe+E
ykCpWucTLsHCHuUPAiTBWr7Q6hJJJX/KyWnZx2vbEqfAYVUYuU9RCj7W43sVZCgQ
JiOuOCYPsUwqLkIER6nnfBzWY8hxRQ/V9k1UsjSjpG3dthJg46P+Oe0yCJeeMMjQ
E6300LyVi6zU0SR4H1tr2FgIvHLvSkxaOTOS2raAHAIqGHQcAbRyd+DSiiHv875z
CTBESJlxN5Ilm2ENmCGn5n4qi9sfrlgRoId97FmYV279hsddk8ZGlkHDByhd9cfq
/wZSZfEzTy4I0Fp5PykClmWmlGKm11pIX0Sg3Bjgd9PJjsFeovib6uylO6D04KPo
hdN1V0z90+UXCxDpEV0dXBCU4xGUT+eAtmJl3w7U/LuNjaGADxRTyPDIZD8lxJst
kSkg770Zr0iXIPBSDHoCwF5oG+HY+7gLGgEvB1xdceEYGh1B4fAnZ1/Y6M9/O5eJ
zRgj7SFiSUFzRYUOhcBf2uo5fTvnPKON1fU4Y8cFQxqKuAe/SRGRAc3AUkrUPniR
KpjGabo7cmXHqxeadgB9SR8eq+sBX8MA/2tlUIoZfgK9e/wtKpGi3jFCWEtKJWGK
tsr1iHvI6EWNOmVblFijlK7+5vt2saAl8P1zun29Cfkl/6C9bqoh6Dnn6zUHDKqX
G7ZxzMbnX/8M7jtQnW5gPD7R6vZHz8Q8MwMXdLJKVgvlIKrPEwuHN2UBEnW4Xker
wxOzI4MxeXTgs0CNQ+Myt4le4+xtX+hRAWgQBnakP2vKHF+3ECVaEQreoM+Uq32D
JVXNoj8VLtZpTFzth5nBHHo2gbnhNeDddYLDSwf8B3mlv4uJu/0Qqqgnc1xvb3uK
iknBHDEfqcJahj3KT9t0VZGvYJxVUVmVb+/aadeKiJVmyjmpzU1jjJVB6WyJkHT4
g6XXcbPMyfBKtFW5Z06rMxcyOqmf/DbqEXggMZxUW8uFw7iKe21N6eeI0ZI5UhUE
j9fPwZSd26NAzWRLh+kOutZNaBoyISIgItMMeCAokJjepk9mgSLxEA79BDSqbDst
sQR9VtQUWdnu4BL+z557+t49YZOcs8uD6PDup2w6Ql17o4Oekb/ycC6bzC2TfkHT
E+Gkk75gdoEmmUWTUN1ywy0/v1Fq8+z0aEXHde1kCbY388Hv+2RympQcQD38ETmV
4BRI374zohXmaoW7XHwwDhESEyP+Fk+H+l2UMvdeKV8+vHeQ87Ocwu0KQZKUY4G1
9fTL9BxlLYkxMMRAXOVSZUoD5TzyTv0HpI4TTfGuf/a/rRejWaXMLgDcc0VzePV1
7DiUZBJBWLLkOQMknxMSN76cI8bl8Uy4Alm8PDSOVeltx+Zl4kAlnVBAnbiaA881
ItF1hP1st3UQ0O4pFxspgzh0JgSsOvzo3x4AhYRdB0YKmamiOMR8/d+NcMdBdpJf
NNKI6SJIXDEfAdZD+D/xjyhA52/9rrO8VBU7bRMsWY9N9U6UnGZw9u3crwkfDHKU
rw+wWijW1/s3SbMlTnblNqa5tm/F1n7z7dGcK40XThtQIRjvEg6VIPtIUIZAwC91
WUMXypiQuw1TEW8NjBvGm65+qEWXcFKeQ2oc2x3VoPYu4x4PrlsCRzCPnO8uek6G
/GXkjxllxYZeAUWzD0BiQDlX0tKPS/WxzRiwy3P4DsaWNTt5NHiUJ2Ug8TbbxKx7
9LRXzl2TVFK6W1w+BfhaIce24jKRuux9eX4Az5SwAKXlqiW0HlhQ5mkkGt64+LZe
tVZ6M9ufTedKBc5JmcTS3eJn2AG6+m6x4dxs4mc6pVDr0vylUF0hPSt/puv+s7Y2
gRj1icQAOcLt4dKfYYkqIonwyc900VA5g2SE8pBcj4pA/u0z+Or1Dhjr5yze5NCp
qJGz1S07PYrPbjhy9agV3lwogt6QKUj5MdSl/VN4t7diu13IKNcC68DFwKPnkjLE
wLVy7ddLF97HpOjgLNA4gBrniMCruE2Nn3WqWb7wzbnobF5p+drC7TQrQKTfWkST
SNmv8oBEM+DsfR5/Y4KglCB2oFd7LT4nhuXHrt0/ZFQj6gxbgyUs+TnPM1PKvCel
83HLSv7O5FnlCWOX5V0UWu/uFhVjCk9QNxgG8OKOj0RbAQvxUCwnaogjLX6RRGxI
ArKRGB0xZYDNm0ZPfoUm1DyZDuOlOZ7uJsJ+/rnOS32M3cpYJcDPE5dzAazxFrsB
4WEHSIYBfUEYGaEreVPhGIj8b+gw/dBZwMNJ3N42kOXi5nWH0ag5Soe6ePT+LMeO
sHUWjthabEHMVn8dG7r+SzwcNFdAamlKV81jNer+UuXS0HlyQ2djla0pGvs0s40A
53VYxmSsyx1LwPtwKn/qEVRKyvVsA3tuua0Hn7evTYJp/XBHkAzaMgxOcuUrynYU
LZLfTdqNajJE42hWxrehQ8hEvJUV8o3pMlBT6H9fznNr8OVX0FtW8EdvEjZJgRHI
qoQh5BQjP4URgVfzXEwz0kVpNfCJspJnsQghxvqfaujNaOc7tQ26klruzIUWiYap
OOJMDVtc+r/sIE/hsxbv6D40oXZC93TS/U6vbmQW6DcAoAEk0T874wyVJqihVI5v
dk27q/Sgm7HigtYhL7C57sB+cgs3LqaY1y2hx/O2DYqFdht5KAV5BpLE3mIztB2R
nAsOeanKjPogwgUXv8UnjceUBRGjv2yjS9xVdCOq/niD7zIEfAGr3ZIVHDg9MSgo
8Nn07PsQnsxY91vAb8YDs/VZyyeuGy0cGtkGaa2BXLFXLjNAnTaokkiqER9CpgO/
sEOKnTBIokd90WFSH/NKSIA6ACw5XKz6IqYEXhhho6q3DFVnkxSeqOf5IPoiWjyV
KRTmiaGeO0oiFE4WL/cFuJX146q5+4rHz81IkDjnB6VhVgWydkhQysT28dYdq40P
eGIaOuDvfKEMAw5Hg3wjO7PkeWBSe5hXQJXSIVLd4zBS8fyvbjCRfjL5vOizrjfo
QqDKaODhqp+oJAlx0YlDQlxNaj37IarAxY60uVZxzJn9m8SWPw4p0TtDoNkzeOzx
VLhnO7V6IueQgqbKxe8IgAeOW1151kqw+BXbKiX3LpPJDadsVW35b8lBZYc4m13S
zLLD0mRShpVl6EPmzmt19NvokHF7z9FYmXfrd0dgT6FDajsNgHAWA0e/0iq+dMj5
HogMhS9QlWmZQIjZOJPQdQ9WqZq4q8zPvY2/bodyZjgEkMOxAuEgm+5C48wKbfkq
ZZiQ6S8UY9xTdvCNI6rsTSq07SiKDMf66AwTnA1DWcnJw2CEp3HR99gSnweiOUA8
EEAzhfqLUWFEIKqebVcp2WVVAU714NDdNnYTD2/IvImt1jRWtLny7PVFLKSUvU2Y
wznpzc32WHLysybclfi7K4p5of7WGL1z3XYjxr29Fbohqc+xNjetpH2DzMsVWSRF
HfaHFdhoD1r2C+eD9+jK0RsKKD6c5HoXViFrAim2QKP+ctJPfbmOfNM5L8ra1kFL
+GrCEBr0os4g5UrlOM8SGitpsHUrcNOoUIu65io2FTZq60zhhLIJjAP3bizk4Awc
6plbV0KE9mq/lacEE1Xu/6uu0sI7RFoZ4w7iDFp8600mhwaS9cniytTrcXDEusu6
AOZRGs9ausOydSOpB4YuCblRtfVgA7nHoBPCkmVmP4o0x0C9puZ7F6z1Wcn8jknO
h0P5cbOss/jc3b2BVMXXuPVdCSV58ej+O4bVxQet49hnTYCNyarjDCxkgjsN/nDa
TtCFd8+Zipb3dvhgpZN2YKc5C8dGl6WJANlq4vePK+PuAxoybyqYJzrNsyFOTfmh
6+/CFSkC+dpPRxAxge0df8chfLi6oNLpLak58KBwyDwK+RymPNAEbHznasPgGfF3
miC+fg3HqhspxBqK+NfYw2zJL9rNAVP/XsD7QX3yTwa6JFopKMlBv6OLN2CzItk1
z/DjAU57fvRZEJTyHPvZXuM0CRiapDGYlHaFulgIejWvIZNtWP1JNatRUi3yLXhd
fHwt9KEqUAOzuIIF29YxRmGh+o1jOIa1f7WCrMCK2JnFszwdIG6zP2sKd2tCT3MC
VggagCLL/M89RIi/TWUH9HdmoTfl5M/jP9HMCSdymJq0QqP2DLnQJVourgZwCM/Y
wgBK9qwW/GabbMdV4MPvlB8V+Qv0FQxIe3geUmzjMim/6FnBEJBYjp8jv3hLW9l4
ueSi8S8PgSsi9ga6WTNVJv0wDEYgwcxKezIKJMrRQnZ9oNpvS5cm8b0u62xFXZAJ
C2ZBBy6sBvWevOQf6yxF1AsJ2kyzbUjXW3ZFB6InDucWSmAQPEBhxr0Nqd4BAC37
ECU1tuHYY59vAb7goRsE39Whd8RpF34wcBzZ/NnkIqkcrAK5v79ZxGxHhvGr1T9Z
a2ul8qYWCgWbZeKAv09PQgH9P1qpVgq6mrTl2zQVAFbNKmtkhewyC6++dLPiz/TY
G4cUbLExfh6MCix0f6XvE+nCfQ2SsEqTx3EtYaoZRS/PmD5uAd+YU1in1/ZOUY+0
C0MFOYmXu87indphaZTxbp18fsVUGaBRagwTftGdXHYTZK/fzFKo4QM/NOHk0sNR
5pqBAxA5vdxdLyMjIHJkKtA/PvFAmTIjqFcDqMSanEbqopDF/8vmAEIyVMbXzqam
mpGXc1goqp/YDHBb9CDvOu4wkjgv7EKOTJNN7KtAhuV9KX8oYr9xZvXuH3/rsZlU
SwE8S5fuOOlnPKBAXGitGvev5o/IirO9UVnTkI0YiHLnshI1pFQjoMGk7WYm4wB6
lNwT3pLQ2dFvzR+JZNaCg5iVZL5rRaAUrWlPYT402kkDDbnyB2f0/Ag3Niys0YRt
mlFJ4FNw8JljZgoyG1hzZ2ona7qge5MrP45f/vjyw46AyUz65JZuayUfmd9vlUhe
x1MJCLKDzCpTW8a9VUUn5+4cE3EYPYkL15PxL091RzIwuG5jR1rHToPDUmMt4qa7
2vwdaPgRiBwGtRhdQFx+CHAYIX+7C3bqrM6BgqxgZbC/UmHXfZB9okCIFOFnIGoW
bf/MpwQFXL5N6rLCmi4mwgh2/JNUe0koQOuov/2DXb06/0CfSgXW4itaL8eat09T
rg45Ek3b77vrZ0lxZYskgEGjnp6poTaSEMCOlFGoZRN5AjCGLw65FoNFJ624NVuA
c/9PYB7ml7l1BFO95D0cb/2NhrKTpqwJSYpL2mAPw27Hw3xstd9xzhL6vZC8kdka
IwMrcAHh1mD8GbiiFe+PVq7TMySw6111YK/TZ+SCS4Xk7JnKAN/eMmRZTUCgNi6a
GKBLtVKOiPx1EZ4ImNvI0uvKYIjtvh1ZUugiuMmzPn8XvaUARqFL/HqVRpJb/Km6
Sem7WOTzRHfJlk/MC9fPhhCvsIJ68Sp2ko1Hdk3gegJBD/zsYs9lZAaBys37MxFz
LynohPHV1utOwyY9koOw4LBqxE4IdrRTqwZAMSyljrqQ7j6Z9+ev7gxh6EzAp05G
ilOis7gcw0hJ5+LKUlZGaJHVrZ013/xgDpwGeLeMtW5BRe4IJMOAN1nK6oOerbqK
vTIL0B7F2u0QxPaLaq09MV6JdOB5KDFdStdITjYLNCKEgmSvKVivUEG07PzhyCrg
MtpIjQrilE+CODsb6rI7mfkSl/mZUStZtQFOMa7O35jdIU7/RJx6BslCn2qRUM0J
nYYGRgZepRZvneRQC9rrdmGPZZd7ePpK9eqHyIddZyAm3Jaki7+M9ixamTrMcx5e
YigpndVGQE3lW5z6Ztc/qNcG7AXYIrxclvJ5IzZnBfkW5sBo0EN5IPlwOYz17BKf
vdR5Yi62AbrkLeA1SA1hIsdEtA/il3sqg2mJZLhSvkIafsIxp2OED2YqntsugjUL
DmqU344icDlBV4enZIR/KxQwyBkrK3ccJ9DRCMsfAWVASnccebb7//hwdsGx2uqo
IeiBpFKPZBg/orAL7955AbAybXBmdUmsCw2haXZik1ZcrSxFnsfJkXGg+5AZGhkZ
Y/kJMWcsLY7g2QiM9Rh05FA9kJMKeYK1SJ//jsrjjUbLkWQsBOCQPMSxqgqiJ51Y
y9qiS7KO4Jm1U14a2rwQK/yC+5x6MWHyiU1B9CnJdRG7D6VuLTDnuwEvqGCo/aBs
+2A24VXbjjnDlr41fgp/o6VVbl+ytmDWQRZIisIi/pnziXlPPiw4TvFAq3BOceR8
7hlxUak2rYzVNyBHBZQYctMFmLyYdjBKGEhCFHViiGA7eOoD4IH2ZMB7wFAblr3x
b8YP5VIF/gnkVAXhE3WD3ROjfK3M+cvvvb9JzJSdGrpstZGiq4pdVvSkIWeXp121
REz2vfpjWkpm14npiKG0vXTE9ukH3LVNOQ8ROedLARoxoYBrR/KdYCxsP5kEjNOe
KsmVf8igPFqeuYVGC3xgFUSGoWexQtJZ0s6sofWjXjcf0qyARv5u45iWyGBPmNuj
agSH7XqGIkh+D1aqUeQm1cHeqhrdhivJX7jhHl2MVvstalt+vdpNnNWIQuKm7j3O
ugxiFFFQAm37vETrjtIdvU7HVXW9xW1c1V61rYtCIcmpJVm7w2tmJcpGUfptBOU3
T1V2rprTxxvNSCNaVtWxVJEWvt2QWLbPIy2ads/AIQayogA0IuzA4X155bfj97RE
ZWnlSL0PnmtASmxDCpv6X/a2ZuB1OS1uEczeHb442oaCj1nv14A01IjbkYiAMwGt
5dhqq27pbF5CCLkT0mMRYcufoJQdZd0GcUEjOH21QkGjq4wZap6cLOPQvKsjNEPd
zPJDEVctiVdN8IEeyKkLECvbIak6OLHE4q7uhKlClKNZdvdcwkG6o/Zx9HTn5bKO
ORMd+gFVXaUfM8131lDBPMOZbN9d7KK9NLiqu7n7fWDplF1aFNGSOfYtRiSDaCFN
t4nVaUcw5T9y5fXh6NtZUFszxOupVT1kTcnS4S/K1NccFC21MMFVi4ErNGFAYUVs
YfDaCJ5PQ81F+xoZpLEwjGMlhAaM10sV7zOayOKJ5fJjcg0CUt0dM1bm22G8FN8q
yRmH0bsWMQE3Lo/UX7353COF7+9EbugPG8Es47ow+6tG//NaBDNoYIjacTCLk08P
BGqdGd7dsb6/2xbyTrcWz3ZpsPLrnl+AaCgT/hPGg4oGIKMEz4b3R/ZkSq5ilJj8
dmbMe6unZIutZC1co0fCakF0O2jpeyG0tUJ1XpGub0qxIoFUgX65vLfcuqwztoS7
S6IB8sVOUgQt/YU6cUsnJycHLHb+Hvb33vvT9A8pGJExxtDUc2VB8lBD+fNpanX+
I4OQuufExLK9p/qFG3vN8PJ1w+tZausb2jX2UxW9oyyugJHlEPyUjZk0xLPBrZEj
ede5amKxyq6wqA/w6OhcrT7DROc8VthE6sJZzLd0/Qa97x5jUZP4M8FVikMpEzOI
Sw57T0QtXNNaK1B33qTxrYqXCTctHuZljV2YzwEPPkxMB6WJK8xog6uu2ujOXRNF
aHWiDhoGuEEWyS6ctEayEDORqt9QTbJopOWKEN4I2LYBOrJgouu4nkmay5R3+E4M
ZPYGzXe7J6Hrx5wqBiqWTuMs4sodOpX2R6yV2PeDOAZeYKbHSO1pV9rJkWjYODvG
z/tR3bW3MweXZmlwfV7Xx/KESGSMqk2NbX/cSY88YK051pmo81DUcgGk6D8O2N33
YD2T8b0oIxkkgAWO7TptKccsHW7luWbitvx9MJvjuThJYRv5Y8bdRR4QWa5J9ss6
Ni0KJNxNYNJ9NoOiM//CSfPV2QH9Ypgo1hq6LfRONAB2tiKu3YczELaCkZAmesH7
JIRwJo0WBtAGhl8kFSBJjWhLSkNTaK9P9u/V8UbnetytS6fctuLL7TgTWZkC7MiE
Tjlt+5amOWTo7X2uHy0ZCVBV2N2XoyQJF56bgOSz5BR5z810//vZpyo/WBK05kiX
GTKXucLetlg7OKEjt3/2BtoymHqjdijNOPdcW+7Vs+ZUXRqgqwBXPwaK8U/D/3jL
fDRp5fPtOARCDQyJzhFDOJczypLAJI/qORWCX+tI0W/Xpt/CSymsBfiZkO9GLpC2
WhndXjqJk3rgRmlQGprS2bVevJqIgDgVqCGuumyddUu0Q5HXVHB+KXmVI0G8yvDL
wMSXVek4jNo5srD5Gw89tdTJ0az69wHvkuZ0LL8626KKX9A6K7/BbyQ1DY4/5LfQ
lY1vjnLmSLlO6AxJPl5vQf/zhDa4qxtzN3O4w0OBD6hqNPmCxPMCXSmADsAsVFNr
X2qvbHjUutApfXRlhz88X9JXjwxpgbYDzOcO7Y3x/gNn7ODFHXmEtVuE2+4k6tLv
QoYVEIYOkuXcUxP6Zo9d9TplPCpiUlpQVkVDx4/jrr376gmppyXXL8E2jJ1fTb5m
HHapWWPoTJmYfoCPV/kb4jqE6Q4sF7YSkgeYwtnRJ8AylHQingE5pujmUUkNwTN4
H/XNNxegwYPMuOQzEIE8OBVUvYl5cydrkaIZSr0UJ7EA79uD/3G1Fue+k/7v8jSC
FrkqGVu2g+OAglrPoPvkCD8Ba8hry3u/puefbbmANsehF/q2faxFlh2g1rXHV/64
8R6n0Ew5MMwqKR2RUxJP3PzqR2wYJ734UtA1sCXTYD0wlVU1DfmbRse0jhl0Ar9T
/q3rEIXba8OYZvK/1hl4hV83aYnUHZ3guvSQUSmrKN920EM+eHlo2FUwc3t+o9Fg
R4zSmbSAXsfMwAwwfFynftSUFFF0CFDudGdfkuNnbCn4grF93LM5ZzrYJNIvfOBj
6gTjIxCFglYV3UyLSBkhwxIWkV0IUOHYMIKfrQdhE8HpUCbNwn3hJkVo+NlZSkVb
jF/yxKb1I05sruW7SmsL6cCh5Uqujn7nrFMRjHC2csVyqXzSeqluz+Wl0MBs5FlO
Lzhe5Cu4JQb76zF9FiQz6zRbqww/GZsirlZ+MJXUZmYeRIJ9VPsVrVppnQjrKOqu
Aaf1rSNXwTL4oNt5Y0cKVlSGNLmXkJeRLG4TMjQDhBljHZ4PKcn7AX5EI6poVByk
UdU8YfHIPJ5vcTypinHslrExcYld3ATnZjxpHblgW+o5n4uZqOM60s4zZli47GsT
91OXKZ4fQ+WSvn0vsfZH5EJxeNR7RunGNmoCL3EpmUIMmHPR3SiZkuklKvBWjVVZ
OEVAd1AxkOpPAIZcbtgzXUOEvGbq+HON31iSKnAOQGdtp3Tk6+QIZtd5cEc9C3c2
e0M5/FwA7Cj6a6dS47qieSJ+00h9LfHCOpmmok5g62DBXrHPx+Si+O0ltfRjn4fr
flCFI0MpoQGGJPXFdrpqCii0rapuksYcHgUf+ACkDOxATGNezKqs4QB8sXwDG8hv
JPjFlv81M9MPQd5dgB2k2GTyp4Wqey7bc1O8AG2LsZMnjXnLYI/SV6iD0o+F0Vmm
SGARDJhHlyYFaF/mbAOPwGwVevo5Nr0f28S741FHfsKER6ixYb4rkSNnuud2NbNd
ThgtJwCxA8n4f0e8UbnvP+BQfGgi7vs2Vb5E3rIYO+K2dWs1anCDY+INJd1PGGK0
6Is8sHZU/kdMdveTWng1Q2S8gdpwxdyl1o0sPFUXjn0BU+rY4VjWE05BXBsMjCoQ
HzHb3V9Z8LOI8+0K7r96HQN8ec7Nd4KWxW0fAc07ihzcjKmQUt3Hck+aJDGcd7gK
1JWPRxTyd2cVy3+ECZDL3n1fc4w0KPV9NWdwtEtgP7T28gI3mR9yVtKrugoibNFP
gLIwuOiJzlWRAh3KrKcX4FJxbSfUmBvQAVRznJh7QQn0GgjDIedWYGdLHRTRNghd
RgSkjNwdLzewkpk8xfJhzOx2k1ze7CT4cJaAcXd0a4tlFOYZ6gSHtvWivEJXsbGH
cDhsD3YJ0O1PSkx/llPWa54gBFbG+NwYKvD063gPQHXQZO3U9AKDp7e5bGQzBSAr
YwOvzdI+MbqePZKxatmBmlboCcIVRoHU2jQr0pkDUzDOaJjAy70CF2kp5YgCIznK
ftXO/I85QXCVq8JmscfnYr6hFwKh9zgs3BxbY1Q0MCJxSmYeo1YuiT0wE3AORLZe
lYCA27OZUMRzwGqcciye56y6y/b9r1zwdVNVttTu1WjCvuSt28WyhIBOUmcG+MFE
77HdzJRZkogrpKKq9APqZZf1Is86MPkXLlg5KebKfNBvJxBOdhwPt0PqaXRfPiy7
uksePU+QXrnSxL9KHnxIawAc1TJJB547Tce8boddJnpbX86Z7Gjjo3GnMlyz6nkh
jxI7KYwmJz455M9yOarrWDs9iEFCkvrPCMVqA2agyZ+xxz0optV/WDgLpA0uG42Y
V5pkuavn7U2eJHal7p+iApsdNKU+sYGUyrTBSb1gpIZ8M/gq4RoNjPVCWUuJHJuC
YjIlojncWSj5XmIIoZy8rYBzO65sNBP3ss8diGTwrAu1W+3G5bGCsXtkAHyX1y9i
ljSmqGcmOi3Mi0PdRkeq7KY7TYexYStsWMj/8fjFaeX3EObZABTqkxUsf0mnVUe5
yJoFz7tkW7zUyW5TOORuiDrJe7Y5/Up9L2N0Ze98YIAWWQZ6I9BnU2pIrAIhnyfA
WoUCVZ4OK30Az0eSt39lSgGxHA4Zq5vwRSzeRrytMFBTjH7+IHZS5JHo8i+71PMb
wICJt/UNqSC3KEeb3mDtmebcJcFodO7IUdwE1MpzC/so0gZCOcYI0XPUIhW0foX2
oQc/JwCnbiFO4JXnc4a7ZSfe/2n2t2+NlhlLdqFUm2uxJn2uI1e1/+RwsBwUMPPo
Rcw3sKDMsPWOUH6W6nzp6PzBIwKitOdj/ZPzb4XNENzeSl+9CViT19Tf0JzK054S
Im7iRS/kLmvBWo9dgs9eqZxgECFhy3HvlLLVPNOGbh/zieae07nVg2fIktjZvv+p
ABpyIPy7Huwe42BkTbaQXdUcUCRJFtlBXz0nSY+uoD0VTclZP10I4Kk9C0RLyAdz
uwncm+OPGXSj0pmNd74FyC/sucyZxAK50+SwFLVwekJ/AL7y0nx21t7CtvMowDtE
Hl4YkKAXcUmNV1HEbqVf9hZSLSXTcI0tfjjFRj7/VowFq13oFCPhxlMfM+4XP0Hp
0ITnn9FztNIB4IT3t/kpI/HSaa7AlcOolcYAxPsHsjU006w8vrZvindoTCh/TsWS
UofvN3odAoo9GJZwuVNO2GtybIi7P12a3gVFOwC83FuzuXamAvYlQk7zGYxw9d1d
l7x0FeyETYg+oOVplpazJiEDVeYF6xr4LioJ4u8iB15casCEnZYupwaF+uBsJX6U
7eHyeFW8vahdZnUxe1hf5xUHRizn13EUR0JIf8+Z3XqSGKPTgnfPzzc6TpXjMi+r
vW7A3dCbS/wN7riBcS0WSX6G9RujblLqVYyBsuxYVnptQQ20iKhpgsIQi2vtDW3c
IwfW7Z9CjcSg62M5TCcjYdJgYCRRSU7zrIIc+7+zXG3K9mdgSlkAIVElnti+MPfU
EySNRjcGztaERlw9blm1A/oUXd6FVSMUp6hFTDQYQD2Zn4HtuysRAFH1O1wb+lgm
vRsogH8lEdMXK1LYng7P0gHbuTiEE0aoOvk7FUhukcj7wWYdeEuj9nGdzM04kQ6N
O9X992arjIxwaC7pMvlbJ+7JNuGoxxJRGpL1mCSRFyziGTC2hUud13W2vUaVhcRv
55O9sX8CkCvGUg66ntB/jSng11sOkoHQKFpFKGxUxE27A7SXciQqblcMMcFZ+/XQ
A7EskrDNIg0t6pbRY29tRJONXm7J6G3Bg6IvW2p/XPl6TAdiJNA9DBc7dGcm42KA
9P3UjqHmG5iAx1e6FmxJ9/a2NpXoxqo31yxwyedDVYCjB14IW6sfjYUEwckMsBSG
sWH14ez9Q4feh9y5cHLdDGWrBhtsmZwRn2IHNsseKDuEIB/xwvWmpNchib5sZgvM
QZ9VRM3PC0SyB9v55KcVaD9WjwccoCZ5Gq5PBYToSnH2Q52UWGK1qaxSab0NB+8n
aJs4fBsJ9PlaNdkJodry4aGiML43xv7SsaJeGNgWM7Xf52H+eJT829/awkf2H/AT
Mujng1ebuQmj3FgQy1AZd8uBeno32Y9gOsA/ag1bMLSDJpLCBw3uHAAJZKhGpaWd
k1hdpAvhv8WPC8Re1LwiB9Ct44j45lR5VXlgsylq9xJ6+NOHcJUujAUQwRKn54xy
gygYFHERT1PwpvgF4778RCR+U3xuzGIt8yuNikBO9HgpFPiZIxKrwn15hnVX36Gi
wdOMfXeEDeXhSnaFBQsksKhe6q15goOHMuEf9hErhO17O2J+dai9zxjITAxRO2bb
ZXgsaJxdYTWyEfki0wDx83TtHa/ALIwDhUGxc6ukowDQa+yVow1H04HuMOqNaQEf
zFerNvf6QZEftJ2/hOSs5ISX4w2FkYnkVH0WbciakzkA2ngQdM/PWXTSB0TODUAR
cArSvUg4yyKt6JLfhpvljgj82Wg0c+9zhHruXhCZ9xmDWXnlPNQKn3Aytj9UPAe9
kesMeaee/V8QCOt/92lLhifQHiMU0FE+w2H74GCqb+bRaC1lakR9yTu2OwAqszN/
zZT0zzW3BlcAPkqZqTs3bran6OkXl0/16PSXJdqsm1YlHHV3onttE4k4bL/8rn8M
V/C40IHQB+nLJAOUIGOrToo1BFhRQXdYZNZPbBKSY6gOH2fLkzcsoG1faruxW/VS
ptJkvY4J6PH6l2EQi1FkIAImoHjc/CPN2ipBQOb0oS3meshtLaqYF7H6YvuIZgq8
Ie4lXDBAb/7K0CsSYroYayGD+NPRzWic6PEjhROf13MI0mssdakN8DdL8awknRiD
D97O4a/v2SLY/3fz1sInW2BJKw7uZBCpyInq+7jRp91cfOc+qILmuwAQakR7bwQG
e3kBH9h6v+QLBjTdIwSXdhQ6mQjG4ToLgDwYF7VZL3VQDnR6rbNSEpoxTthuqBc+
DLeytIHeqwu6V6bxv81/63AapW2ehWLovmArs79MsldatY7A+1GlFjFE9NLivCcG
XmatgJ+gd+adRzM9r8QVYxkn7Yy64fvsffODGNp7hEV9G0vyGWCrxu6o/RVq9jGD
j7NWrPwZ6hkylu2X+m58S1NZ4nx4Lw+fueRPXMdJRaY/4fs9yQsmxZ2HiLhXESBO
v+dvBHt/mZA4ePRG/X/svJycwM2oILTEH5wfIkrHi7uvzx41HhPn9sh+MSUQnA2a
W64qvaV1Tb8Bm9DALkeTy7pFjyIV3ozcNws4RkN1FPwCk0bqlnAvQnYQgV3pqCgw
s2cruMk7PexAxBi/uSBk1SsUqvv1tfqMhs9IqBts7BaoRZkTKVAwZBOdjnWV2J+/
OYAIicBLjaTSKlYvT5FwywHV/CEjzjpQYg3AIkARqyQv1c0YSUcecbxPWQ5DC3hC
YPDmzv/kjCnFcjNL/6oBnJFIcT0ZAgP7jnrYLR1KBr+6Dj09rvrvpmumIIo89AyE
qJ9h0GeU6/4yaooYjyiUsA5/ksaOfIHqsEKw/qBCWre0XXpFfXEm0blPmyWFXGeJ
KgBDPhUaLfBQhci/F8WtkvrQEJvf4ol0Tq0TWr3FEkSJsdn4hokVz64KNeoTbC7j
eye57Tkw90wdP+jRgkj2IOHfcvPR+WZjhDYtAOgq3ioLeGcMYjF5CRfOQWTzlgzB
Cept4k2F1QFl2YB8X5v+XjAseqgwjtJFMZbSCYiVsqsmjYwa8uvDSpVu/3+A25Nv
rc8LRSoqdc64Wfon4g6Pko7aM+0ovzpJeP9X5YFAiHCymKyFw+Q4FHyo/5niGFLs
a7i3qtM/wM1ytBkEFrUaWiiLF6iln2xyw7apKdUIGAegfOgtF6o2j2kj6tDZ56NR
jnI3E3CGD0hwSM1uhfFkEa6xB2EL1d7BUYmH+Z05CiEVHyNq4nT8piedchMiaqc7
7qSSrYfK0gAzJHlghJDcaMQRSZEpNXTEKMxnd2gAoIRc6A7/vJKW8jCyILVhtnqM
jM7gypxk4XkJW+t79kFzvgeEdmF/EXKHOYYLgjkdOrfKuF2h5fOEICZTHKBW9gwF
Cufq9Ozm/i9m8U99FWObsBDbJj/Ci7ADRL+rYSSluIsiaJDO20CQ5oQzTBKsn35J
sTMPdtw7OURSOk1ARv8WjJStCdpArgBVTZhwTq0Z3RSZ+JIyE1uN2o10sxbYrDZ0
lO7guka8nPg5stSOuJu7HRK8aKutY5MkI0ryPmJIixhe7VKSIqRSM4Dp67tfIEI0
0yRIEiRCz6AGom67INV0pKgjx5tjlEGpty4wMNIjRPJZThkTqW1HpZzE+y2HWWmQ
7rWoENtCp+WHkytCeQoZ67X7zfYEOIaiclIWlQQN552PFq+hPlHDCUekTvtF5EcV
6CJ3MWnQeaas1Xt18PtM8O7GIEFQmRfN9+aVYKsYXSOohnTYNiC5BTejyphEp1cg
Hr9aag0nxJIBHkhIwvRByhVzI8xoChTFGe8/XJttLVV4YlMpbZ2qBGZfy+6J8X23
TT0pKd8IYugpvnPBXRs3HowEYORN8B7mFv2jqJMCSsbiRYNuJ96GH/xsa9rlVGUM
R1/rpaG30Lis3+3iM81gZOI7aWViKOkQw6UZQd/skN/EzKMeYkDjYGN7y0Kk91IM
8EV6A65W0fBoQ7rvOGEFA4rB5tlHpjGcXQJmip5eCanaP7mlDZk2dH+iq3yX3q0b
e3vdBEBPn9ubIeqiCCAAW4NCfaVcymIwelFrcSls8SyY3o444JX4StQPXQZq+aK9
DxCb+wWfZw2mb+maVc3jedF6sI57OCCxKC/lnNVWY3TA2btQtTEEoZh8BHU9a40E
d7gzaQGt8AYHUaN4a9DmNuTjBZrFYY0kRlWD0HUiFLR3d8KhDhS+BUL2f6JfGewO
QP1KgMUl7SFDAc8fPYHwXg/zDgkW2rz1vCJWUfWrr6EqnrS8SEvlVAdNpzhQ68zZ
MpF4SJCqnqWZmusQAcBRsY7uXY+5nvAb3UbrgVs9c4Pa37zTW0JC1pvsP++LwMYx
VfUMRnhNnOtbi9wlSH9ygoWe+JjqmH9q771+eA4NvSySoUj86/KhnLe+4vPsCHs/
mByyT1veYvSG5jWl3scW0iYM0lGdvUd15g2PFzeBpKG8WF6wEUGY/OKAsZYW13QW
/EfMEsf1cFxS7QPE3mimDUiWFkjgmtdo7UdCIVhpU9Cdf6thFNv4ldw64lCRQe/U
L1sfp2fYK7uBzZ07CHSCVEjW2Rd34pU1FMdAqaN2nc2rlMIsB2C7z0DMu5n1i9eV
fdmhEmepEnVfSF9sgpYb8iKlFbTKDOakJi+rRbVrPAstBfp/x7Q8rJHduNi7R2K2
v6JO2ZAX5FMH8Id/771wUhU0NCNt4QUeIDu6n8WtKj5tij2cfnCl43Z7FXXOWcS/
assX89mPuPXgKLW0JDQTOAkX8yH6vSETfe3jfSYjtmLgkUdVub33dqveQ6PE+iHb
J1e3ASN4A1G1WFeCKJSauKCxXSTe5KYpJPcgOXzhqRBI+b6xsuwRyP7cjnkCzNaE
c58X4JqmLsQlzEMdAa+5cKr/+bJEx3htrCEjXC9hMcWSlTPA46OD3o4Z8o2pfexn
7A5TWwFiR67JHagSMsVPFxbYlJr9YCkxXEKkCCjlUKTMAy632sBFq35ltA1gXMGs
uWFwkExsK2gYqjfyAPb1Hj0BUqq3KYM9apbdewqrCrEMJ1ycb7tu+AYc35jdCjEe
zE3ouGGm3rx96lhN3QRrGzWmx5J3lQvpiTOzmkaapF9yeyjRev8P7yxCeoGJ9Nm5
nBUkPPQjP7vitsB2ptL3m+F5BJZQo8Usn9N/Aoy6OU3FPTK/T6gpI/zgOiAPnVSx
jXSKf0Oqz5XJVdPHGQaNDqabuSSgoRuwKahURdFP7uzeQWOXan4NSx/e/i5/JvMU
bKNw8fVDhCMf9gYZfrFjHzShji6ltjcPSDFpedhUagLlIoabc5DYrJhPqgGTJnSg
hUBGvd0fmdM3TXSrSfoK32L0RVnT0dmuS83V40zB+6DEMP6feazc4btw4peVuys3
KWxDdOrg1MWW3Koe4BuZ7TFB1j0N/AqEC6yIBnELmBAhhVtuWTgz9a7+Rs2CA6l0
QtCq6Dp4o230IenvYEAwhkdfdYneByHvRVcCza3LcpiZq+9JQ6ZobrpP14KM/2q+
W4zMDLQYkLkONql3OLpn9hKnAN/4aSH3JVqoMTeojj3dw98Sol3SOCrvsrfIjs8p
x2odymvvJDBUcn8etbNY/NAL14FM1Oi0GdWN6Kw4ftdb5EfoM+D4Xhzb+zblzqMw
R+pDNAp1yyviqAXWqI4a09u8tGBTvL/1e3vMEet9kAHLzl/kzAwnRV7Celaaa7tC
QmKLl1i1u5hm+qR9BtjCkghDhQtVSPoc7rHIq01gQEYr0kxkOnYjufyaYC4+GJ0d
3Fmz54i6HAHmYF1/QNCKjNY2UjBo2OgwU1NqfCvBLFanJtYNcr0o10Py5rYcVhlh
bgUzQr7UnTTEXtN/kensbxe9o5btg6KSmwD7aVwbmTnDwRJx4yZPmMUJWZ4MQqSc
28pMeunew4LbVCrGwm27shN8q8JmMYZMzku9hyTx9Xvgl35aC1EcTE736JE0UwdG
22Syv6MCzNIrPcrVue6vnnmkD3C3+HTZMaLXard9JMmC55EfjIjSfh/J6M5OFDKt
P6Fw6yMGt8KaOR3cWWv9nqJz82JGxG52O2CO9ZQ7nU5K1+2DxAN1oN+ASaYPnuk0
qvxWclSwophEDKTT4NKOy5n/UCpOoNVDKUz3NhqKdDgHW4jQW33/NRMc72u4mWJW
V8zEOET1mrEcWK3L/UeOnn10SLRinBNreCJAVEKNorwvh1LqIG4EdBF5OH+5zDdB
tOWsNeZM9h5PHOQH/fQG4MwfmgbwAC5znMSS0rxHCeCDL79sVvv9CEqxLfrBxnfM
UJMb2cqjAycWvQAazjChfvBFlUKX6w/tQ9iCDPvaCreMm00epl8s0DdddCcOf19B
ZOVFtdOE3fWA5LOdZyxc4bXkDekeuslTLRrnxqV422tiLz815Dhzw8ntJNNbU5ea
LSswOHrmzwLhndDF2SstQBbGBLM3z/q9i3KoKfkH72cUqxw9PAeTjRrI5z6C96f9
7OokDR4JSwcWS889Ig8lc3LDD5/KaHMIhJefWs5z6CpirlyDQzJ0sGyyFfEjO2f/
4W4ZlqGmADx/Q/T5d7kEBc7E2gbkn23dWsLP46O4gLi468pohtiuPmcrN9loK+g2
9zIl8uQwrlbvA1GOx25n3BBXakRj4GQb0Tk6uenmxHLQHqcZgb12qgnSScyYtcIr
Ox0v0cfS69suzYjEkt+FhqOnhnDKXqhKJa/MP2ps+leaBnWpmy0wCPCkgCCUDP02
oszuPTC/WCqnOa/X2cdAycpsuZeZ2jii+L7Hm74sDixz3o+e2HmFA1EOyN11n57t
VD5XogaQ2SezrZ62tL+wKl1hzM1gsvtRkQiy7wJahTaVUmjFMWqWOKIpJCHsxmK8
XCqGqIPIEOB67Qm3xjBFwwFk/gNe5qIKTNEwEc5ba9m0gFb7GZsjcyEr+xtNUonc
5iSJvFlLjv35MPxiiyzNG87Qlk/RACmXiYUWP/CIggGaBIrAyy9+kTMn3MDfM8Tc
UkK0yWNuWJpa72Ox9GnkYHPmMxGuLu6HyiJ9rz/FOczvufjrPMfxzRsKP7nt6udL
DGJ6Co0Z3bsE9kvGhsq8270sYAS6XvWzrIRCzQmgLa6rKDG6GXgHCQLdKbyDGmgn
YYh3PNa3X6+9BBLegE07oYiJVjk2bEpxMnN8lT5rS3/NmBNVC8eOgCJBfXYzR/MW
IPa7bY6YTcoQ7EzmAZ/Fs+yFiuyufBQFObWJoQDPlMspAcpBCVVfbDY/TkzXzEZ/
Lc8Ij0e/DtvrZNEN1HVKMLqiIlESmKBv9YVaHi3nZ3Lj6g/baVOGr5aaqZBf2R5f
80ntGfrG+VbB62cc3uJTQTlGCzaFKy0x9wtvKCK/wzY6rkMaL3zo25QbMrt34gUZ
XToADfLGTaBa04n+/zotFEKfXXayBNfGbpxq+pM1L/JgsYjYzV3PW5CCEkhW7kuZ
QK4ITSWQHkvl1tRrPRIvYS/UUgWdINIfI4JhT8ELNdBoi4flXDQrUH3MWYAWWJcj
no8duyBE4v4hoaqUnsnNSwTi3Z94fcRkRw7hMsMvhAj+KYsz//PIrgrga7WMQWiS
yWmwoRB16YhSUmxbFMyh3LGqx+O6rwMPYc8nP+PNynll8u+c/w/Xzgo2w9myW+6c
mUS60urgNAyKTfEHSYCcDF9ULL1wZpRyURau4EV53J5YKYSxxZOFHmTBI5zW5Pl2
nBXxwnrS/vxJJwskiaLSZ1Uc0y+1DlaJ1zDHqbyoIS3Vs0gi8Vn70b+A0psnKiCZ
640nbgckPS6/n0NnA89D4rdq1tqeK8/dxHzJwioDtqr5A2XKMkZWimTBjLh0IYpo
iJXpI79JNv+DMdQqHkZleey351lA5lHCuG/A5G4V8ZBY1Poqf118yiRxLC2HzIo6
upoOXPvh+xQa7+32jnLGMRXKwW5GwVVOHUFw7nWDCVtnq1IqBZp4hToNzI6lD0K2
RmYXFspMY3pHu/XIDLaT8AeblprChspKdIWPVJR4Q5tjrpJl7U9Nc9lHZT4R1s4F
kmIdGyIid1OxMs3Xn8oCI8ShEolMKPhEWGdr7dOSxbsOAIIZxFhe0HHW8wGBZXi4
olN0XVKMrB0dh8hNRtKXJ1USsprE4x8KG0VapMoRsJzJm/kn0w4ZkQyCps65Xz1i
5OjHHhMgiejIxlxqbgdWtBd7lLVyblbpobmr0d+JXC6PW4HtayhoJdEXkMAL0Xgi
tZ2DulBkzE007ZLQRvkRB/wHXAAWID709LHRxRk6oSZijSCEhw9SdP+Yap2ezvAQ
DBAUxE0Bop5MxrIkqXcf9SjxL9pN/04Epvho4WD5IkW/iBbdItFjBcdGwkHyP6/s
ThaOxXGePLcIsS5QEPTLDU7WIpgPTC8Bh3jJ0zvxiM6MPGfJAboiVWEuXZ3uc6Bj
qHTgVIj6bnlbPrPYVl5FecWwvXjUXU4HbgshUl2AlN2u0pz421TFWg03MD3ehl8O
9maN/LAVooDUQyy96Pohl7xcnUdG3F+MSIchqojb2OnWFZmhB9Vz67/uw6YJ/jMb
LlF2AkPry1dRNYxAaLNiu2Cqyoh4aXI4QDSMAFwBLXOpP+9aPpmaLMcLmI2D0MZi
caqMZIMMZqGyqHIJgtdIqotA0zxKKyJ+IB9kPG1Eb+X7gdJynquvJAVIo9s/o+mV
czapnnbYq0JymMSUp1Cy0KVkbhreIUfwVrGeRvcPsrNYJD2VGdOVvLaexCckQW2w
BOhgvuXuLyFnwSVaW0t5ix5DJY/jwAIetDtYaHBnq8fpLPh5mHu2ovZDIM+fofKz
J8klo9cdGXYkTa0YzjxigypHoWpRDeyNSvwjcEY4VRw1sXNEDApEYRYl43JAFsWl
AkaShfiJdBYndTh4jvgki+xqMzrBPsZO1M5PiQa7sM68XUUp9wBzvI+YHz9ttkmW
oQGmcDy2mV/Do/fTOjbJZsFP2kxrkr9sPm+2RdgwS+czkiexw/NTA/6wJLVdsN8Q
QdL9b/nG9aq/uIxH0HZ4ae4EYmgM2J7/zEaxO5aCYQmYRprWH2zdKyvhulcS3FMZ
wnZdlYBj/zQzEx4m+c/HmMbCw70NEfEJ6XubUcnha/akW1zSJqmr8Kat/WF4ZrOx
Durq/VR40m5MtQKfqdonFKxT1cAutxq0l52+LoCdbas5vzi/xB8MBD2ST9SMdgSC
aiyH7jhDgZAnECoBvVa3pw8kC4jvbIyu1zuXAbYSnNiIZvp1TlAOyDbrHJwwvCDp
9RH3WDvhJOJ2Cb5HP3XnWZE/QwH1TgBP+PORpaAMdLaEGss5bgQLGuHzTGU39UMG
XH+fkQsU7Xa6ujWf6d+8G/EK/71Lc86yJ3UoEPvLntrdt+Lvbr/uvOpwgbaGjLrW
M9TBTn6/W2qFpjj+LYei8Xbs0J7JL4DTJ80GQpwfbARZv72URwVdBdLCv6dK4FeT
q5kD+k6ywdfgcWyqWPSGtEBRr9iPdjFm8mRbu4qZj82clwAyXQtaAcGQ2bqVuI7J
6ZPlmwaCqlthRuY5vvo+YGKQWaUWayB5+Qym5AzUB8TPQsZgenxnsuDzWjTfvT0M
hy2DTyZxdmsjvvq5uP7lCySqY+o2eDfOCBa0NIZ0yLSWCd9wTl7xqoBmfMZDv+sR
oPQu2oYp9vlN8d/bFH0tMSxL8orfmuovF7RzOl0ufRoB8USLIsh71KW61cV+tuF5
MFTdfN/fGS0Z6hHK8iS5tdB/TGk391ltdaIdTscC39TWgA48YU6pxjwB8LmBiLmN
H2ta2B1ypmJeaHYp3+QAd0Qix2ttd2S9tNBMKr+rNH43DMOM1hhhTrEFQz3GF3/9
THv9SJeEnaEpPdKlXCN/1FqBTA7KfFnf9LFC4KWngA58JmbpNIQ22v+KSKJZGGJR
yxn9HZg1qr0/a2y0WygWbaLlC70Y/tY3uUgdMSTzFZFRcg/YsF3wcMhgUMnWAJrr
xWKxvBnqBHgiWvVc0RLI+dWfjg2fsE7S0LzVGK3djURIfydnmg0QdY076K6EhQBf
4Af4qWVNFRhTN7L3ofizHk9edbyt+3m7f2JXdienhSNYKyq77TkFOkAxSKA4Eh7J
Wrgywr3Z4tbAWroJGaaqmPi02sOGnE1HpQ2FKeufbrIJ6cOsbky/feBA41dWHIlZ
hP4zRqkr20fOrw6j2fzc3wldFePERz8GqMrtdIXsfjz3usm/oTwujzh6ixxR1uIN
Y1N6MXdlURWj3PoBGKEFTPNYnEYf+cRTBtUbX5Ktl8+gtx3nvllXzSOxy5FxzZW8
Dy6SeNUDfL4WNSHk16SR7wXzweIwB/E3w8izz38w7S+f1unTyeGfxf9Yf1jqqV2N
mHrfSfDosXMQixjdA98TaEmYTQO5INm9ch/Z5pKzRrFax2JqF+CDdoR2YFM97EUl
XgQA4V7P0cCX/ZwCePUR9P6eXby0LLcALgWYEuBQbicQ0zsErZjpqmLGhyqlY7e5
/T7MuNNzDNTa4E7i1L+ovXyTR/uS4EvlQIQ+fDq0EXYV773tIVOy2nJM3OxFGEyz
Ayr3TJ/v0t1yBWmhU1pQsIkNwTD9e8SLjSTXZDBOgGcinUmjm7Yc5IfnazgIyeKI
AWRAnLOyfD5hJsiYNETdx80ngU97wLU36WCBESLRTFL3LvpZ7R3IJE5Zz8BKCAyl
1/BtpexNsVRTq8q19kZZtgmcNEtCfQcfi1wEkioeSiEePjkh35m3Cg2bd+OAjNQf
zrgUcoyaGX1w/vvKAKBQ3UFchm5KGwvCSF9tfAX1KrBgemlLyGKqrz44r7aSZxpL
YFKRTkdRYRMHC7eJ/exhhSU2yGQYLd7v4Q6W+iLpnnq1faSY3rCDneUb4lu8WYuJ
lzMJR/Ovkm1FknA2Z0Rz9QTVOq5DB80bVn9dwUyhquOV84r516uCjNqJkre1uf5M
wM/tdSLe92pFf74WiPK7XhEJUychSM/yUFc9kSY/b3GDhuxDlu9vmI3PVONUXA9o
wO57X8MRt/1brLlr1bid9Kf+6AT9kyPasYo8at9YWDghFgK3bWL329p2Qq1Px3OA
uC9QJVg0e/XEaKVNFRqlGUF+Zn3Mow4NGedKNEvx6KyR7oRS75s0b15EM8RktCZP
EZDkZ0Yqq9iRtUlSaZ7TbXkKVnJQ/OP8OibMlgGgqW71HKrVV6T2ijj36Yy6IalZ
Y6LNY1ii4YKk3NZAjqljRy1/vPI7768AY8vnMd+ziJ7FObs/8ce1KhSwOCgGqZke
+gS8ZZmGszBSbw3DAEmPO/mr131edFiDvEa1veypEoLfXtdiGoybnNZXZz0uAaZ4
E/RGczgg2uPAOQj9O+PE5snodexYg6b5a1Pu/0Dkglbyv8L+I1/3EGdLbfaA7cgT
bfD9C5NgxCgTm7iYLV+8hfzNZpHD1W9WEFAEdzsf2x6LCwomblYQTwsbsFAGM3ls
6Qxh+yiiMhJxgFDdq4o2hH9IxP42IzsX18sYOOGCkn8WQqERO2Apjl6HMxiMaDPz
eGHkdZISj1HVNKieGg825XzBcVqyGRKNpZhyifHsjzzdsnVpcxJJhtcgMXhsPXu6
LTnb62gtq7EjZGcRMtN7rO4OVy5tJeq+hhnBO0TKgkcubXJ+FEiOx53KPxpRmxt7
5xKmW7/ghTZSNM3ssn9+TBQk68kU3hS5UsQFEFLbi44ek4ll1TkrO2rcwjNMCBmH
un/XS4dE+onULeubY+IuL9JzIxJ1LiMa0rQVknpKM3gfM8BF6DoXRNSICUTUXbJB
9VzKaSYdlf06fqAig2EmcCAdr3HvnmAKb3mhgFe+uD7TxQXcalAiXjoYD/IxHFcY
z08pPLt2lKV35KRVaCMDZR0DJa+VKr+TygyPDPyWEP69K6RYkIra/i3sDLcKoECr
AR3wExnxmPkAVSjBFajiMG/GVYXetNeHvr/7Nel+Q6x7ctaCSIP+5dr4XJGZRgc8
VbQj67f1UNm3Pvyp174uJsHU1jXojuBhtwrU2n75taeQFsW5HrM2r6MFKMC29L3S
cRHwtTXuvKoo2KsmRHjOU85pjd8MyLO17+nCjFKwtpueTwYBHKpv65WjeNCQmjGJ
vk9cAhRLcXgc/JsNtM7BqVklB7MeTDmk/jmSYTlVSYv/3kLpsrcxfC4HLjUO97DV
kHEOUy/oofHMwoi7DR66S4v2YfvWsTI9v2oMFk+psxuvvmOAZuJzwkXWK4W++SlB
FN7OFYMjNXxg9bUfz5q3DiP/FXAjI5mR+bAqtL7NQL+my6b2/MNN3qLfwVzQUGJC
P5HQBM2KtPPYFMiMVJRyxfc0of3jzGJZ/aA6Y81yARprN/b5G8IAKJtLAvEwxVdi
EtJh8bzW2uDn4iZCaKtftZbdT1eU4U6YnO6dWoExglPea2r8L8eVIYmLomP0pGI1
C0qdC7YVT6RIFdGKToT5MF/whibDVepMffesYvQAk5xrMulNMn2a5NpG3pCEGnz7
bkypl0Q1/JF+Z8PhsGEOEj+dP4ssHgPCcgnnrym3nNLDhtWdf4ZRlFFrzQ51QTMH
fnpUKqItWI0HPBjoeri1VtkZ2jM5njO0DXFHmbAeRpwswGsKUWoo/0+FOMeCo3LO
yLIbeogRBfxonUH9ldAL94LdKht8vwItrii7c349aTph3WkVJUUduQeFgP5OvPn0
44Omsy83+3CaQuKP75nCHBjfoyQriM+j13Hzi4S+Y9sctQE5t0t0MprLFt9SjZtj
odf2PJdJK9WYBEgP3l+0wH/YJ9rwvSLcr+LiSrtxVj/8eSx/qLoWK5HMaT4etQzk
Fcnn7blkgzk2Ukp8KiH1sduQ5btsJox6zfgXPEhpIOu9JhvU+sszd8wDG0+juClN
b5DmtoVtLZIFchtg22i6dZDHxIWIAPDs+8WdX8DM3xKjeLKiTRQ03sAy0Rnr6Yr4
cfhKYV0js3UhQnuf2D83nLEgdmmqAxfUaG1V9WKXdC9eCt7kH6aW+7rYtqwgasZ1
SRZsOlHLDycwTZZuQljxL9V99ZU2vmCNRbn63dYVKP0abZGYZImz/MrJ52vHcG9m
gdgb9JQIZUgfiW/NeJQbhx9TCVdc6EJykqIWf++KBw2M9tOLzhZWBTSzCwtFQ8wR
bRh4ilmEyfhzm2nQiBpVphgss3qkXRvWTvRFWa9cvVpulGnJJv7nDc1jK3hI5n+3
vEj/noe6FuAFnlUO4E4pul0/ntddk1xHrU4pi8WaDtic3njSFkyxb6nWpDKk1vUF
w3+JgORESXDbZGhyQkD/ZgUGXJ7Y8I7hJ6WbwCxhveTRFHBOk9SbtzUXnh8y1Yj/
22HAh4yIistba3NsaYwWWYbCA1dnv5tw3zoIWaRFs+OHPYDsOOYC1ok/D06IBMNq
drLjG1Sx7lasiEGkSIzV1nORTomAk3en2dBdgSKl1vuVNjf2dDIE1quGq8dPwquk
t15FTEF/VXKRf9GRCPmXqy4nyZ8nFh/WU+3p6s63M9Fm/Hw9XeNrYXvPpXAWRK+D
/3T9V5BO9so6PRNit08fRB21dybsW/ptzLBAJLcvwQqIp0tOtWkIsYQ/tn2T7xCp
VKvnICAWHY5nGFO8F6fgKRHdecuD0JMAItkpQsnEsSA8yK9bMCwtlXkRjQ/Lmxc4
kigfyz6BE6P4OjEftSM0s+T6grr1OSzFESQT3vKPXbTjQmyEGOos78nbiQtXoRBL
wgrawUPt2uU5QZJtBwqWQBQviRrVHXhefWMDu7ksdKMN1HrhkUw9YHBJGSjhNGMS
gHUUDDaNGDyv8cY5bGGbSyYLDv/BtPy45G5HI7Zbac9l/Hbh92O04DM0tMnvR14A
ypjTYLNUMJhwuRH6IDvrT/cHLq3Qgj9hq/QjtCcVcKEx8NVDunSC2RhZ3TJWZqBl
dB22pR4WZ6rJzNoJKxsOMQt9vxgzKDBgctNU02sE4YkicRGDqd5Qv36hiufZrbuc
Wk0Waam2mNBSrJDkOcKkLfsxHBM5osadXk1Sv4iR2mwMMJBtnoV3Zn5ybaA9/o58
MkxdqwqBvvkWSgTbUqVTLduEm+kMpRn+hgHVLIlESPTD9pt9LExI0GDfhRCi+6ji
LokvFa/dMlj50ychOca3B1J59Xk9DZZIC+vBEflbgG18uVbBE+ER6YqTsVktCgH8
LFS/YMB1dgzpH8CWxBYJSo76S8EVqEp9uj7c9WorucTPO3IRWjW2Ac0vzVBJ0wdc
pX86WicWSJxYJEtKDn+usD7K/noDaboMTu6HfQtNpqd88viz9+5Bnra0XtThS1u1
j5Zxl1erTGPOVbYqwF2g1o4fo1YWMIZYXPfgTYak9EqIXZTa1BkV7HQDX8whHRuO
mqH72QE8KECxRWYno8PODqjhcgMmLjmLm0DxH6+xFgfymdWP2DZTo/ew1A6MXxPj
uqiTEkBcusy8NV10qdRunbL9yRD0gTGWgh6xI0+t4GkGbx4CqlzNihl8j9S4HzY9
qSCTVT2GD/SJQZOc9DsBHxgBEy8ktpTChHzqddcOHtL2Syul5SVifBYrTO/cmq+r
wlRvg5dEE/n6O+ij9EtqykYvpoWHhXa0JPq2SjHbYvh2lIaNQEjVwXBI8NJA3aIp
P0bld+SGT5u0II5lWXU67GSh9IqCdPYWcwjJW9qN15HyQ50mLo8PkZboUip2x55N
JSyDTQ8zLdKolEvq0gttHnV2+vSSYDA97b58IurzLLqvcsWqxKHjAhy4nfVvFNRq
VqliqZqKMgzbKxRtMIX2/jnpSP/0JrK9HZryV5xWulErq4IKfs7wRbqnmYtRVhkN
yjd9OuvXkdp1MCWUdxptADY61Jjt7R+ngbHJmvLoqVnXGHbYfIB+2BmFk5hzdJUM
ywsukLPBI5Lf0Px6sZjl/6rkFJXW6U/RlzpSYX7ORCUiATHnnLJ8JS8o4rpGyECq
Rw+88QoAv+rG1PtDpBukB1apco9nJoJbCS5posvXnxCXJ8kl67F57V6T+7udHyAt
bBenf6gOHEpeIz8ykcOBfKKGIb6xiht+2PFkAumZg94eDQ7Ho6lMhAE9VJ7+IkTY
RPt71pzKsA2A4TohJwtSW1FFL15hgr85JVVuby54aDrwM3CVAzs3tJE626eeCa5d
EOCeVhfSKXYgecP4aFzLaX21g/d9x6kP/KFiv7aCUiomT8HFWcxBTXkhRf+RFBkj
Ok1L5pDsWi2d/rdLH0MBQcaOyCFBYJBo2e4gZCQgoDQzc1T3X1+1ROdPJ08nB2gh
2MmsomRrqSbqmU/w7GDr1TdYBkNPrBRebqI20IsaE38PnBfmBhNl/htao3dyYgiz
zzvlkslQA1lyJ4MXKbjbbr3FQq8CQkezXf4pLpCIb4L2uXE+zbkU9YCdQXdFmhxG
/EKhZr+Onfy++RKWFOTe0p4/s7M8Lzl0PFKlyMqMnFAt0dn31g1wprvBybi9aADO
JKky+caWBc5oyy24lWWT7uuoMy4oH+aC29ax/qg4RdWXc80E7OqtrO/ZkSilRDqz
3UDCzbpJm53MBOuoT6PQS+z68AucE8qVt8jgk2PtN0ytXjljRy7t1VZPjn4B6WW+
Nnbt+ey2Pq5gATBjRw9eHqb3Uez16ZYONzBzBd2pqoYCX3KVv12Il5ZF5OhD0YOd
tt0LTqpquuum+b/AGJUDAegDMbp4KEULNa/axeIJ8gnlL7siNYCicS5Vahhd9eUi
KiwzEZkgD8l1zpdPijMrQBvaxhrCUEa6lOGlLO6RA1itOyBZpeRmK17PKnh5cW1t
OKnpTCuLiUGR1TIjryvGKz7RyGqfgK4Zg3IAz+0Emm1cy/X9r8oIdBwx4TZyYQRN
c/JKeLY0AMpn95IKx0aQjDB/QxI5QtFLsuqH4WYwRzjj7PQvEmFFcVEy2hpd1Hew
p74OF9u078Bb9iQL9S28znB6qdYhKyqJivBfma23iOZSUWg3ILiUhx3ELdnhPKKO
nBwI7LYZg4OydnTxD6RCuLNQqPaghqY0cNooxAS6QuaJIx8lMy0/u8FdxwL/5mQO
I7pmuXvmsR8kin44KjIKv5ESICyqWl7xgOcl9zbgE+Tjt7WukuN8XFpUzXTnqU8P
I/XqTukKX1al13EHCz6NgDGRMVv0fg7D1pm9A6uKEvf011mysYMPCAXfuBXLD7iu
NlVjSFug9Y3V8WbCVf+c99Kc4W9fWLdwrVg3ic5rZ2WR/Kx6wtI33oFPuQXYBmpY
9kv1hxGwlbTQi/sBKPnnjS8JRUe4RxIVIKlarU9b3C5DFY5muYvC3J8rsimvNRtH
UQed7VImsKgA2sU+rEWpaXS6OorMEogjmxQl6IFfgc99UhwmeDax1Z9arnbw7+VB
pqlCt81wTOlVvweccsY9nMcCOSSPWH3XmEMK4564dmpGLGzgpmX9unODzbI2Ri6x
BaQ2uHOrYdWVbu48Ugdx/VUE8EQvm6WReUVqCab/wLfqHmdH+7ZLiB1rdISV35Yg
rpZlohyDnh59inKU3qG3dldj3YOsoKB+hs27AfqViEhhPPyIoMRKnGsyYAY4eaeN
/vka2L0ZXc0HzC3PVMJc74QoAS3lqgBN/saP2B5BPc8KVeTk5IBvh/se0F/UQhJd
UNeCAg8iAsH2KXLEIPrJrrmlULA7Ec5SWMLtoTBtE8Fz++/6FXG3zCrHEJbdA4ES
GqBqoO5QXswSSNHvQb1zxBdPj+0TdjfM+B85aUU0CKJQIeM2rcUclh+ghb9mp3B1
ct+Plx2GdlMi1Sbo1kzpLLD5vtaYCHvdU6671nHpUDIxzTrjiv1Tk6vQ/9Bo6+l+
bmDaXogwZy+5g1Gj4UOi9yJiXtfSYxEX86DSFBl9O3W8AzSxtRR9Lnpb9B2G4Fi9
DO/TjzfFXpNA1dslJ56GtHbESYJLJHxkfFnB6oqrdwYgjznhApW4ESKMAlwoL2+0
IpXCU7ADoyL2mqgT2cLGWgaIl5RYRyc1+47UI2tUu2yP7KLorFdcVnPqiC8dnPhR
guWmuCt0ipXISWzwgJnsDtrKUAhu7L6Egu8cxPMY02Eutr4avElCodvnDVjXSOHR
4byGak0sa2DI29cKlrRtuAUDS3R7M75/NNDvaEKG01uLcL5FaQggQWln1Gd3bBpk
asVZptMcdkClCH72nR0XpQBaCAjYLiq07Pk2/IovmE9Dbaxn/aH9uIW7ePiPBkEW
+dz3IAhO1ZEp8TbOayIggZgvXqH5MfIz93wdnBdRvf6txzlZU20lhyXBPkyRI0rv
VzWp8QkAeTf6aKdeXHEOsjiLMQ6eqmz/6NwfZ5C3TsLNv3U6WMK6QIDB/tndkHuk
fAXJtu5yGH8EDcszchkPaQbofxEB2kyiBRGyPxX8z+WpiR0Wis1Zik3xkgwM97bH
pglfAkDtvbt1pKPoYaLxuiAh1rdt80uvEJHGKdckBMEF0V24WicOUdmjaEHvXzag
3dCikKDOVfmWpKgAm9SQ8Z83+HAHaR9ZT6WoV8SlJxWiGSWV9lgc2HFAVj/S+wIK
GQB0SnWmk20kxLl36H/d81qb4SLTOomMYZt9pQEhdNXQg7EfGp/gsKG4tWeWY5Wb
oCSGVgW4YGK3aYmf2pEXa//FvMz54yGRFWJ7H3iNutJv/Qwqxq3g1MyBsoNj20lr
qN8ZUJs6u44oBVP/5P0K8059thBxPYELDHc8QEOzDZ3fxEvIENs7LXhLGpkPzDxI
XbBa1ErwKqpVBtAT1VnoZKkm5QuTdcLBfYK4Qc61i3SO6+bBi47Ixzr1EcVpnoEg
Blw5DoAlNJsse23o1lJhYhkMBpbp6LJ4czQLNUT2FBL0LJGPILrsifWk5s49voLK
3T6q/9ZHnVR5mIbNPvVwqhaCXZLRXhSQ/RALhXNGMAXcATylyH8i8pcGDodJKa6L
Hhu6OxhakpAeKnsIFbvN41bdWbr6M46Rl9lyZLxv4CEmZoj2FtAmWVUub+ZCrZo7
mfaldtlhjyRZkJzxGKQ2X0+y8ov6RWF59vi1EriCfZTckVU7zZ8euKSr+LGajULf
1+yajKBt4kSKenhYwx05ntXdcnDZVj4mJ75PX5Vdk9Qa8eweEW2Fj9HUvllUrA8x
z9e2yc2eHsaARM6VWJfif1hfExDsfPqAflEMOe2TLrKzQnos/90RkTVmDOtWoam7
7qsKmaXb3IJ7qELAvjtaKfCYAqxZ1wuOai7/0euan51JLerGc6gOy0CBkUumQbCu
OGd6YKMbeYbvdLPtCnrEVBuI0KF4lo+v9tPljZB4f8DNnWiMe2dCLllqr4zkOYTI
LlUh00dlbM+ZEf+a1HMZ/TZEFWvW2jzey4yikxOU/FdtDSzDdYrkNOHGga+xxBq5
mWg6n4i3MacBYPlxLFEZr8pECFlTUXnpeDXgr5BKB4zhzVw2UMuNVTr1qKacPUGj
/xzw9XVfZI98lWuQUkGObwE7q2Rzvnz5ebeylMqd+iykkdQaXfRXK+BXiBSMkYg4
Vlyp4A5XzZ5dKjYm9ze9lTvHt6FW7L7um1hyifThy79eDYt5To0jP4zA+3sDVqnQ
ZBBkcYPmrsq3FiHrl4eNsP+Yzl0KHBzzSW1MbXbZvu5tM+6YiT6k+uJtHkZ819D+
HY6mbY/U02YSHBgLkCu7ZIrY1BwOQZByV8FXYUcyrFyvDREKr601T3y7npNxvJp2
oNXFvCaQrMzezJxec5SYvk7jgaGtrzZLmNBAziguKihH860V3vDlPOWAbaxx59b3
+Cnk4A7U9pdxprsdZG/xiJvjs3fGNooEk7pmv+IBYGZrt526bFf2l62UkK27LC2o
PQLJHt3Ywn6RxVoLBX/PD0Jpet39hDbWb52K9nxlbwImJlMW24j49K7hjphoHzYO
VhXWHO19Jkdcubyx1FCaYbmNukft7p5grqFHiQSD1RybJvDxGxd+0giRyTcmzdoe
Kcavki0WgKZgw5RSMmpWrjwN7YeYRJpQd+OpKLKaAcQf9u35CE2cajAj12+iEjxE
IuhAcrMKMb2IfkzEHVHh3+UKknQEr0fAAlKTVVhR0hT9Dyy2Zz0phD4dCUkYkwbq
74CK3iNrPR1KdTcpk8FOgE4A+a3eQ3/Bw1pTslaVSx1ze0tEMFidnbDQLB7jsEQ+
TEF6rZok2g3bY0Yf97tTs0rDCkR1LOyq2S+dHepEB4giYzvcQIkECz6IQJPlpLkT
jwmOnCWl5NMrsp4cocuDJkPpNV7KKXaeFUt9J3bWQvovfGW21AcCY3iJ3iE9m3i7
N+4paPdfWkrsQIlJykJyg+9Pdpmntl7jggnJ46eKHYFU5bNCdQAKMF1ReJYFpKKQ
N7xRJMcjZEk2+AwhZQMIAuNog6lrcWnnzyPdA3KzKf0hYwPPa+OaK13znxfLzI9c
VeDA2Gyvu/MlTPCRORsHPkqrULC18vXQhM1ophBBbyB4KXokmfe8qe9FfYcgTF23
4E89YuqXjmzpiwvwC1043FfSO6IFXXqyuk+IwYsl13yZzXR7qu2JKryPwGrVxr9E
VCKsbS86huLdTB3Pg42/AyIFRVICmcQgeDLCGY4N2In3poDQchiMpc32zRt1TEN2
agc35JLfQauhwIWd/lsokJYKhnZTXwc+rJy3gdHp1WCgHJJ0XG/6ho6EAofCZ1j5
6m36ORLpJDsy6gPvLYA9vS5jqB1ifXbjNQjlDbjt+hY/Bn8BcbdGk/FxiA/Vonn3
Drx1Bu47Lh1f4+UPDSpI6iB6hmDo+RU37P5wp4/ICbo+bkNVcuJYN1vR7JiQlcWu
n0+Wj38PTKj/T8cTxOY6BIDFtVZKlU0EplxcfVFjh0A8NETxzAshAlE0xe575Pp7
dxPQkT0NopllsbHK7DxHCJDxx3Hg3e4vqZ8D/l9r2kqV6dRS2fui55zucweHDFf8
bLJPnoUy42i4HJhhV+t/9SKotaNwCPMOA3sT3y2P9rlHujZLfATItb1HabMj6bZN
GcVfVdBqJlgvIZ6DIvDFy+Q5cP68HdyjxpHIFjT8qINyP6m8mNqDdeGE/I90B41O
MtR0VxIblj6zDFnh9D8Mx9ccU0oCKz403qV42C2DQgkJxrry9fW3Kqkn7fwATEMB
Bijuzjb3hM5ZYKBRzaqaeXugrcG//WaN2/7VhfQA1XtyTc5AlXyp2n3rD8ue7DyV
hOEPgZPxB8XLYB48cH9YOoCWsAY0jPvER9ge8nZMqYOpg4GRb3l5NPh3CW5Xwn11
0pO47N0/ke7YSgWxMJomp4fMcwdFIOZzyMXb5jAtXLnAfCaTnuppKXE8UtEZ1/Lh
/7gtoFh7F7LWNGNDbZSzOvvTdtC2vMgtG4WsKo/QrVM4A79+MDfU14yTopUJ+Vro
0l5xffccgSvus8zVn1MuWqmXOm6trx+ZeGt43QEG5mvRQpWgUgfkjaVpMds/s60a
8BQKaaZWMHSFVEjUJuWO+7EL30aZlxR2oDUOlpu8zOBwGYTLB0fpmalY9LsoZZlw
hwamzDYv7WRKps7znj+8oygcq1SsHfyMjxnW3rwnt+YpziQRDqvZsG3qfwKWqqWa
ZB9VMD7rjemafSoquN29ojN6VDByT3S8dwC3OLN0ZXZLO4OLONHlrTR8ONny+qeE
i3eQPNr2/6WRbfNOykf59J+RHW61qcNlD/tY8LMQrPegrECGdyVS/3feH1EctLz6
VTkkM7a07msT+h+AjZLAAmGwdjyRCTvH5NVPIlhVkoJ3sMD5l8hnRhqBEG76j9QX
XUxIFyjfGcrVLAuijSPPXFqthpOenvCC2rlirujbBltd92jdWmoRsKCJFhgSH0sE
HwZCMX5+vdSBX5qx4OYpBiwiPZ6hbwoQPU/BSyox3HL2NL4Y9HR+64F+1tC7Qg1r
+9g1+CaOTWcllpUIlSbeCN4iYlqpFSBZ70VKbUlADLAMiSHwfw9w3WhUkfN7MSFA
FuWjjVvgZTCJfAx+3lpX5DW/UYs1TEafB5RvEecTJI+CVELHRa2OwXxuJAlnU59i
yggVV2HIVDf/1ezLYE3lJvJiE6tupAdgFt8TVGH1AAzUTUVr9+T/qalmdU9MMw6g
73ZsnuZPlWY23rsaFLhAhdmW9LgKOGohdHkkOo9yTyfQ6GHH622nNxHRP9PQpFKw
t/Oh7vZUX1gcM0RHbjh/rdvrPWeetny0DzGEfTrDPzT7F0+GARMMt6KZLCwIKbfY
b+Bsh+H4qZP7KjlM5EQpBIxtvgtM/l0TSV4cCWBcQNuC7HD7e+SEf3ZwT8g8swL0
mNzBvtUvDBhqXnxUMGYDftDljHfq76WKvqaujf5O9TRVWG+er35uMQZGPOB3m1yB
V0XgkNwjbevxWSvjZyNtjxK71ckzgJ2D7wMZJx+EDEJLMRm2KcCQ/+hFNulCxmds
Bvtj+GbMh2OIP1gw4B6RfqQGqybTZ9IEeAhxtF7jyCGAdWghTAlem7d4Z86CTmNi
FPO9DwiQHiHtgGy+qjUWLOGE/lO54/2ViuctQa6fIKyCWCBlnvENVt/BUTHwUncC
/My1uPpz2zAj9buKyXnQjRopE6GVHYkWV72P+JLjw50ccJqhSk+Yg2s5YIMfe+od
+nj11ASHUiKXp00TpnuMVLx0HQan5rjAseG4ekA8VgvrDku/mFloBRO1nwbfUr7L
bSkvj+aM8upvJkRmcP1Lvc2rpiygWoVoQD5MI9iVQdNBNXLbX/Cd2sRAkbvatvm3
HYBho+XH75hXQ5c9jqGlXVBMks/cuyGAbsGDRAdNUVoVgcCL6JDtpXWUR3YLGD0y
RU8rYt4894eRphXhcSmnCULJm/0YmyazioFjrEfZ5Uj4PK/lyWdQQ4yhInVVUSVx
y77Aab5dnUBVMaTzhDMvjzSIp13yGRgjRFVeIJaSKzKhCb/H6WrS+J52dnDWtEV5
Wq/Zbke6RSGmmFQbn0y+vucoBESP2gJ+TkEgv/HznByw4vES1BRdoBrKO7X+Wxgk
11y2o+q4ZdLJjqrhWYK3QnYG1NXBPAVvwVVkJmt/AF9Sjdfy5VTF6C1HmK7gJ2aO
XGn49pitogo7yFzk5uIumSrfi36vQU2GA+uV/9jVPefhffpkJGHVyitnrTGivYQ3
+77JekY0EMMubDZfuAuOaq8goVIBjIgqSsu/9tF3R9vXZzyEiyeHQoHcpu0K0iHd
XfYp1+F+4h5gW0eKy7M0/d1dxNXUp64w9obRtxTFn9W0E6Va61eDzzeJe7u9u6GH
cN8jwNXAMs+g5RNJKifvp7oj/xKjwvKWac/PnyB3E3q2AUdRVepDSyNT8KxQtVCp
jCrJCXoy+8eDRo4L0H9lffcv0NTaVaRTQBWSUgTN8rO97XERTQXKdNvYTsNBi32t
v5T9nEYH+tm4oqLfEXOGSWftgmVxJBdjDVR4GaTtBgicjX1tuxPu8g7quUcEsiPM
2iF/kIIojDRR3YqQBbzzG4bc4rai7373gXZCnyh7rOKLmZpqGtfgGLHO4h08uFup
liuH7gf739uqXAgOcl61lpneUJsQu6JgvVpPmQDpvZGXKzT3jtThNWvsJjfihPl3
p1rvBS+scbE1roE3bd9uGk58F1lHh64Hcji2N7fN/khYAvBSmvz4/N5iBSDfKZNZ
LQzAvzd82eDTLYO2xfVvqT2P8b8nIvPyl9YKb++TLWmGvyE0zk1uVZ7AtRinkbQY
7ItQTid+Jx/KKoY3thxls7SMOfZ5DLGK+df/Gvmsyf5d1fHgtrD22vK2MO4Yfgn8
2KpS0qlu6ZGfKwbt8EhQEMDZ80eA/3VHUpJH8h7siS9taRdBshNt0wCRp3gUVUfC
nTOc2KHDIdUg8W4HHRCovV6novpZszr6wD2ddmHLCf4KWz77Qdb5tA9Ou2fF84bP
RhHuqnIOeM1HKJdoJzd9B24Y5lea0nqTDATlM2XBdKU7+nVjK5DLKUjCQYWMrYYj
8cZ6s6OAo+/nKvgHamKAoKhDACl38NaCQaXREbvLZsBydD+dNz7WJVmRg6hbfT/l
oBSH0y3ce96CPWFMU658G1iGO6781oMf+W0l+FZrVw1ZEZgpHMm0Vd23aVjdo7Ao
G5QmzsAB/l6BJPZ1pcUEKw6fOhLcULb897l5/DPV6LVcoqORYwfJg3YJTpYYBNnG
ovpp/Sg7OfPalaafAaJSeLxxYGyQtBN3HaRCaqUel4sD37m8+cRy9pEijamyguvI
cn9UjU9a2UmH9nBKUQQD6hcbufYQhVWVya4csEEBFC2olebTPhMv/xJ9GlcX33LA
4gT/fmyQxe+4jomYfhr8OTMge/I4NALqJ3uQkcnyxbOKIrAL/jU0Aodr/fQnRe92
Ni1sXa1x65SRXXMF69YsfSYSoNCiLSXLIUUw3DZ0cXJnZkjdOwF1zbxYOxZjXBfr
r2kmadxdaHYOUPhXAyq60uv3zu6T/kvHGXRVKUHWg8y82j2qu4gsj0GfGUwpwn1j
Qlddp87edvxtiR8Ok2t21dowMOcntgsI65dT9Og9vgrbkO6sBC/IOR2/piouE/Ga
2bDkcNnqaeHA0znVrduLPGnEZlCv6+s/NTw+NURk5qxASFHczNruT59p3UtBNRRc
QBuxsJxNXuFK7K79L65oZtoX14A3PD4cMpK9SQ9XEXSINL9icNLCQxKpPadQcVQM
JaQYaDKl8NvD812TzOaQY7GxO4nQveT7qb2OaKLs1pQ0yfBRJBE+KNp6X09dDUqp
KaE0Ls6aCqnXA++bsD9AJOx0VE72Z+wP44c+Zf5KStValk/128Zqw9yp+YWojt4p
T9LVMliaS+jNCj9DHIzCAV3j1y9pVuQTyvqBYpaGnNGIT5tAI0sH9ZfnxNjl4Sxq
2aFduUcRX5hICV31qv6rt53wO06GtnKg684wZWgsBntaLd5C4m76wz1a+/LtY3V7
gFoiA4iTZBZnPVXgT5KDhKpzy42LxVzgiT8JXlIFUNkdnDxHLX1YQBS0Z8lK/4T2
d3OflUOh7Refq92VAp5MBPNvEZ1jHKf61pAfR5eKeI/HfyAdFvkkcJN+lL/slUMB
pEswTep+FZG/nAkY/9xJ5QrZhiyc/23Eg7RJ/OFxZCbyZqrOR3NVIlTkOwhFDuut
Ogc+CN68dEJBRkbOqZMXjBAtC2lOU08FwOseIaRZohXRZMsXQWIjsuCUW2/h6Bnk
WsX9foJcpe2MBRffmojWr5xnijUpzoiqWaPG2iN/lX3eLJ38oQHYRcslKDpI/+Le
JbgXuoPI4BhAo0qJpgdac4e/goCGJlcX7QN26zqDCEHbUL2XmeRnIuEh2y9TpIKT
K0k6xHYi/OTi+M6Euqb3+Y2lVPvBHyUBAlx1altBteX19dBOD2q+lZ00976aosiq
2SZGZHONoS7m5w2ssLTXAFRl0bd/dN9CJn8nJ0sRn0xpFM2GbVkyDdccv9ZhTTBF
EGkdfv+jcZEFn5o8ONNzRMrsa1TO7+efkVKQT7UkbNMKckM1X8tAnSInsLhJIImP
WFe2rGOI/2iq5evpWvM7KCyyx4NpksiOWPCMvRpsSVXPA2PTOpyVQuOq6IBLugl9
wL5aAuSfbxnKKzi+k0c91iDwM1TVkOxqTBmVxGPRFcFXRAbtaC8SxnVg0qttXSy7
d0eJsrWBuKQs1DWIKw2eEbopIJVVbxuLNA7tkAnckj6u9y6FYPApolfz+jSaVFzW
IM06uvFNTt/jurUox7OlgTfVglMjEphsSdan4uiDXTxeJywowVhQ2yQ8UALHV8wR
9PZ1VHVeiaiGENCbSLB6UwNP50oD7eLItmYa5UAGzdYcVuBbMsAVp/7APVyANKub
3b/usYaZtQBEa0qrxi1A+j7Upuj6h+AyqeG1/EbNgbYqSQheETZ1yZm8l+gVhbK1
gcu+/nQ5KpLvox9tnyJtmJ+sxSuVruAALgsswm40l6PraQ9Nz7bCR5+US2hKfaKC
bkEwnSvMj/RKv01LFRxEOTvR9nveCZbYo62K0NXvXjPoEOixwCxNF/UmqJg8r9K7
dNF85+a7PDpp7pHyrcgOYtsbAqaQ6dC8DZmyyAYfY6C0EcMzbWvPItrMVySMC4fn
dYpJfoUQL88w5lwooAY3FIkR6Mi9J3ThqHE4drrXvr+66kH/Em3/9SHEhQ4GJjcZ
B1U9lSgCQ9ccr6BeQT2BzVXQ926mabkR5kHb6rbt2g+5G4y4DQsIfnJPNwS24UyN
KfkXvQo4d/mDLfvkiLBNvguWaJgdPMnKYQO555ffZfmTKCbl0SQDqZO/+DUfYOQB
iE9LkZ7hjTp6Udh/i5Zu8wnYrCAMULtfVJK7u7ESiVLfNdV4p7GWhQiU0lmTyR7V
0yFyb/zOMIqq9n0XPajVkpPXm9BuBMyrlFbnX5I+baPK0rsr4SorgDL2JMXx8/m/
5VcGjnkKK3EQQUnDfHuaPOu79Wn0b85+pdfvU4e+7ZDNYtoC7825noqjvJXar0Mw
VTkg3fHRB6qsOKF0qxS9ESA6KAQBorTii72gudcGusjCLLzNC3UK/FX8C8JN9C4K
2Ibe17cAh+b1sXT4Na0etZKmlyk23CRK/WeVl4XHA4CA1t97O/AXHKFM5BfNgCsH
0ONmvaboLLoh7mGX1scnpCn4Qv+3sV6XuipqQskDQSEDK0ZuIXHX5+eqkbemFkco
Wu3usq94RiU0AiW0X0IiTyf7tP78MSmzuZfaC7YGL8nLJLRo8op3qjLC67No7eeK
nkTSQ7F2f6b0w4UxENGVhNM/ccvdyArKDSmsS98No5euhAEKA42AvaKJHzz1Fma7
PMBIZ5YYDyHi2fyklmtgLlV7bJmSx2b1bsTW5vdTPghUf6GeD5EBbSgzZ+4w8+U1
nJ+HhoD7FbZxI7fGJUSVYqhTr5ciDOgS9AQpVVsFry2ZaUo+Hq6KddZtZG/iO8gn
yLUbkuXTxSPJ2P8J/b3cfClVewInNhgfOBHXZnuLWrUe/XL/t7BT8qdstxPXt7CN
6wP+9Sd0OzH6X6e3C/0n4ypQosauhTdsqcNEpnkz/Wlea67qzGmN1lWx21loZs3D
SqHFaOXOSUP5QU5/aI2vk9EEYAG/Tfj5PpLhlGavCm7vwH1pN/t9/wg44CU527cv
RsXAKf+qqsHldTdtUP5qYFKHHjbd5PlNGJ7po4mnQ4vk9E8eSO3jmMU4SgY20VYx
1i9+AlxdntRQDlwEUbAcs9uVf5YiMujP4RjT9arLOwbrySvUv5LBqPJBrrOVNwpo
v9lyQmFm4IexQBowNviB6fCGW5vKNl4xwY8s7lzipQTdsiNEa9iiI1/X6IxyRM2T
EXkSnHSnP3wntg7cklV96do2ZycM3LUTn4ElXJ0v95N4hh4ZwzzfLuWrE8ec2hey
p7l43Mlj6Am42Xy/XmV5659f67cDiBfBhu0bCxQNwG1O89L/KXGxzMN48JTxZRjv
wrA29gQA+3WAwL96p6beQ24zWGdlJdeYfN7lvufdY7tfyF6opF6txnbXoCmZtvsL
lozJfbPTh9xn/8qG6+ipkeh2eZ5gRoptKR3J06YbACMf6I7ivPGGYggkOp34ulPz
poO/oFhKHFiSeQ8l4sfO18DGLeAKKl/Ss96jK7xY9X+TZkrDXreoZZ6iPow8H0Gl
FAWR1QQZwy09Bvg83aLHKvsYKIKYdocfu7EA+Da9lMMY1ntxjogWQ/fvXnCgpb0m
N0yxpRE/aydfav6Y/k1MqJBIaw1gxPk6uckYBEwMstDWkH9REnhFSkMhBucE5+g5
YcrZ9D3PiFAkdAH5Ut6pvT/Ps6mHv4jv9tXPn8Eh9Q/8FkLY9nOvc8RjJSWLb9kz
ADKtj4MA6vRSfIPVtcNddsLm7Xae/wpW+XgrzyD/0siO+bTSYT/lLru3bTpbZBs2
Uegcsjk7jqCyU9ab0OL+vvcMepEVTO1pu7IMn8URtc3PNONChpcPA4TDG+pt9v1k
n57pp8enFArLh6099l8jk+hm/RvsyT+5AogckF2yInOsIhqhM/2XJe3REVEThbyt
0P5KZHxK9NnGGo0mrj0VZxwMzkYeZ0axyjbV2ATPUWSvCXU21cyRcUaEMdoIW0x7
+q5rT4RHbloT4yegCWzYnlIJNJkSdpbDSYkBt8qvRDaYQaxqVbuz5QgqlCy0DdGa
WziHVmQrvRlmvm3YmRLhrkHlKffWRlJVsUQR0ybXHde2zWU3RiM2/Rbzoa5oHmOT
ACPdchZxrYpwZaFZ/SPFMG7O1IgqoM3nVg3DfFUGzdHOX07pwsCDWLugiyP06CHO
byCqz0Vmv1NPBw9gkyiOhq/5DuFCQ1c4R3TrlcQjRtQUlltVsWphQnI7r4QUybss
SiylS29oOszV0dxp2BWDLiIZhRUT20SmIvjs4upJjGL2Ot+ZRMR65rXB+eIObK5o
drG5jPV69dq+KKQkX2pWairg0fi1IKtmZyWHbpxxd02mH5PtKlq9Dm4ygdvVg8vr
Vk/e/1gEIV5yl88SmjQluhtvpTb67YQUggFbhJ8+MQsDedUG9/VIPOVsEMwq3lHa
QEWay7fr+g5CFeEIwIi7eUTGXJo80P3c+hzReh3my/VJBWk4392J2Qyd0qhVdaRc
PdA/S23ROX6MqcnvL3aohcy4EAoRoNClQjUS2xKNFw5eAiC8fU4uO/reTkbfRLbq
jQu4O1SSCUDdCDo6UtqUgblFJz3tr4CgqGJE6RFILLAcO23HfmC60LW7nNkuKBR7
o8DKzixXq3jm9u8D4mNc52a79EQQpZIAQQ063C0Pw1gtTM1o8y9gAYXhMNoDiFLU
RBn8vi6V/3+gORaTdzFsCE6snDJatFhwbXZkuUt+78NzRNR7jcwMyER1PjWOCtLm
Wa1OSVXCvPOMgbwHJ6tcHZQzUxzPTPmWn586msWDv3Nak82iVLyhDgIY+lqoiVR+
45ZeIsNTp4TPB1nXDySJNzcLdV2Vp39iKguMFA3Ob8EnktOnj54tn3nPOy8pd9aY
BIB4Ns0GZaXRYexGLszFlDTpPfkDkQ4GIF7oYDi20bzvOSZH6BI3qefRKli8AiQE
SlVyLVKgSs4BScQXMYiXiVimUZ84BK1GOBhaw1NltjD8vHl21i28ds6198mvA1Bp
xwn6v696U3eSwpCFkYHkDwcDlm49d85lOv8BqEL8kVwIbC9famqkGXPlb4uF9cYv
yBQ8CewFKomQWWYI7Ne5e784N9VElHsiBUBFnDtGSKRWia83p2aL4Cj22tr+WKiI
MuRMiFcTlEgRNKfCSrkSd+EulyIBt6+dtrdEOlUa509iCS1fINtBC7OoEfrU4Uja
6/YpEqJoenf6RQxDU6vH8oC1AdF4HsfkaNsdAukFzRS70ylKvE64WRyZJUxr9NPt
6maK2E27mAq32GTgqpg4frelQO7cxlyBqQa6KmC37CGJN2zTs8GYCRu9Uf3RVzu1
ghNp+hYEw4gCupusRNB9/b16f8uqJLSj0lQ3fnPgllz9kO478YQyI/shfc5uY1/j
8+Jv9098BveovU5tJ2/xR1JeY6H0DbQ0PzX6i4Y8HE6bzIyj8N0gKbCo0zc6ybN1
mJisLVz0FVWJ+BfS1hCz7yuFcMlNQqcm3yo28ID8axMCMqVu1uBQ/UBzWceENd/t
Yw2oj2JMZGzhCIXlUlcdrYMdBoI1/AudwTPoupSEmvUYTu0hx6EaQnWTYXBHWrqn
N493dqNs3txRp3UnjXp+M5dYxJ73kKyDgvGMx+BZ73DdaQ6Bwhl/gN0XpYD/BnNy
nrWxMOmO3LdxAQxZTuKz2+QL0O9XwIkK4hKMs4Yiz8usRsa7AsAgvlxTNt/nDwAM
EgG/NIm1m5JSiOzKzSieR+YsPUt5APEsGQtEk0VfYVQGdvDA0u4GB9n6OXjYbYUn
aJZgfaNb1pE//azuh1rJlOsz4jLw121Hqatkeh8XokYUxEcumpocEckioihYCSfe
NUyi8aD7nL59/pMOAzDv6uF/GIkArqllQT4kupX0TOjMkEnYKIj4QxiiKlCWh0DD
g+MtgMICCzIUe9zjyyPxqy0LWIVVP/Z/UggVQGCxFUGB8ddwgsR7GxVTQDcxz/KO
pFps31Toj7Brce9eu2wOL8cM6lJqPIgbgxiDcm4VxfsxIPRgayxEiuWa6K0Mlgbc
GO0ZhoAmnY4/iH2sA3fuut3MyQW1h/n3FVDpvwKusF5Ss7B6CMWShVWmqZjPVaic
Ls3vXE43NpSotBKX3tUzf1Qc8PPMGHau38Utc2sRCAPgBVx6txewpZ1ZKucKJIii
Jc4ac11g+aEMkhTWSywjWfnbtC3qSGWcjve14UgooD9kWi8SKOXT5FpFjkCKqLtw
qGyfXS1kVNLWlYykfj3EjZyI+zmPTrqjvL49CRu8WCMdhw+J9NwvJPKSpWTeR4ty
np2V/bJHdDLp5QnLM/FVQ2igu7UUoD6IgMaC1VMellMgeFaA5XJ8bkPjG2eviy13
p84MKuodqWhj3DIPceD13UDw5G0eIUfU49umuiLdqwpt0e9kQJwEpeMDWV9490rz
GislIAyE68wsFeCX41yD/5+RHYuLQ2byeqg0RojEVdLYO1Rac/VdVYLcl3qxaEwG
dbs3voWBNRD4IIrSToFNX3pR4/13ecKJ8P0K7beQDENCjtRedDgkebiLP5pp8/iE
H7Ue2YVThZ3wEmHuAoTsk5NKtOZuupNKTGExW8oqB22Oegxw6p414r5ejiOQ8I+E
9djAi7Gd6E4RfNknKyCMOXBrh6+3oHljW8smn+4BGudt5mfzd8yMdmvoY85l68Ib
gVUUHJs9+pKd5WTY79gHcOjjEBe91gJG0OSdgAGrKVL/wQCx49X5ZnPqbAPSjn10
4/o6pSvJAuSVa4453kC8ty+ZUoC7HMiw0KTkOo75VUfZIWsA6OIT53v8GkmxuRAJ
vnGih0vyCs8qLZXt7CSXsk9EQcTsKSoLOAYVPYhn8yOIgp8dzz3ByBELSvYMzKe2
6T5H4aE7hDx1u6JzucHGMPz/hghOK/f9RJe886Hvl35DtgIx4AdW/UpYK/jEUPKn
EZHR75Xyt5l2ysQPAZMf3w5l0RRAINvRY0kewXoZdy38VCHqd1v+LQg6mvGTZa9f
zIW20ziuokLSwdvAl/rBexAIj0psGl72FQZY+UlmHab8Zzm30CdfPEfwUMlEMjf0
sHqYLFbixCCchmHC80MITVL13Qnrxd5uo6kKQ+kdYKfanqD00AaV1lQMK2B1euYM
dx3Z0pXnBJWWbtfRXMvFF2f1Ine3lW9g8JODXdmlqE6Myu6TwyL3oNVOoNNY9U0b
XfjGJ/HnLMVCZiqYWAuAQflUVJICHiCOyg93bA4XR0Bj331HRh2GinReV3jk6Nbm
6EG3AY8BKFtCKWzzpkfCBqg/Kle4GPmKI83z1yECSP0YFZkNjuP7XRnahY81BIgN
1iEPYRH4b3O0XO4z8w1oDI5GMhYJwhU7iB7oKXD33IUK9MoscIZg+VOoMe7EQToc
gL2SuUXIr5HrXPxEgHqmxy3rxMy+4gHSOfZy25d2FK85hK99Q8Sx6jWb2RS7RjkR
9eVb9ryJQ78j/eVkGhRtiOLt3BgE8AADCDWInuXnQqAJKTfo9cAy+VG3OQl9aNY9
byCalZwbGTW9rRZbdnL2wcZRU6V/2qmNu/5bnEPOG++2xJVXf8UVyU1Yy6v0ZeH/
NvPXqxMW3bv2LZg6oU1bC3Eh7ZJtp6gWreFDbz7rVcajgoFHaDa+6vH/92b7eMcv
MsDMZD6JLX7YwZYKMIzAT+NSRYQ/Cib36o9kFnYYM/CGxxmHwGp9tXyRU2yeO+8c
goaYoCZEnO+noRNv9DJryQfArXCx+b11pZ56ujFGojvEbrgr75QpvjXWcZQtcqLW
BFA7yo3SmvAP3UW/zmVUEk+Qibpz6jNf67nVeW/N/lXuQie6VHQDa52M2IEKqYg+
UvBnyIKAVLk4s41zY1cFjKTTAL5/ONE38rR9YhFgjNzswTTE/s0O9i8fulRTbsiU
Q2ajsDYeaCcD9MzVWHOvGlY4+qd93mP4jgJ8ybUsdWW+x3B2O3irObtEsGfWyH7e
P+vx22WFyY6hABdl/UY8xVT4rmZwQ4gLnDMEU9LJFb1X94/mTeR5ygX0FlPkQ20z
LCshGl+1XGzrpMj90i64VbOV9/w+0mLJChLvVxcIzgLrt1jwvymCu+rmWuUalWl+
RhevGGMuvRcnn1dDIwH6ERFDHIC1p0RK+zuLqmXmtpjnOmO1Y9kAjrP7yewH6kF1
H+VzVEApOHOwFe/26+YEgNHtwv67xM4uVVempb8JNlA9YWDJqxGclNcj0vXR81vV
iAI/AP7OtvIULYRl6AzZ4QXC3ZoLxg+GVxbHVrbt7LWSy0Du/b5JvIh6Yq0QIwZR
UK5D8WBxnjGwowDX2mSWmvWM6Rg7ViAAALL7MPhbHgyoxtU64meeqRMiobmDyNVy
2ynKoJgruhoTCvQ5yyf/3kZgvWQSHtTZIW5VcBcSiGiuvEDxJczAIBlrQc5cCnD6
9CRHzKzrhsBr5KpYDERgX1ia/fQmkizdQz0cRqCDRyKolhGKv9pPk4AHSRJGOleo
EksyHsj0ONRiUycFRfsyoW544vj12B/RFi+zYy8FjgCr3ypSm5bqck5Jl29D1jmq
8tOIEVyXauct9twSUCwA29NqjA0V1TZS0TLSpp6nQluLpdTupaOL4a6R2Mwfx6He
ed74K81Fxgi1CvqZLKe1chYVf2eN8BocdyIfOzuLtm9KA46LpPsd7DiM0j/OlWxP
vtmWbcHnNkkWxc+BATGcTM3tS8NCAMWDpA8nnXoxgkR4e2ydi3kY37FEx3MyPtSD
qQrQF2IU6NE6y2navk261ml0Nj8nZS3AhZX3mZQitbiMiZH7QTTZkIqft9JqEh/Z
SVF/5p+GVFPqAto0gBFeJTjZHLsq+Kp3M5zx9bc2XSYnPaGBmQyNTCEWP42/1p8J
eZvNeC6giwU/HZ8v8g81Y2os6fl44eJXNGqqR1PT38bmkFHRPVFpftRRnKsTFd0i
ZqYcq9cnHpt5YiLG8my9RxOSjEDGV95BjrBs0If7xD3nge9e1opmhAo0JiOLbwHN
d3xlg4inUNwLQmvK6InlPyaxPZvB1KNAQeeI+7g/pJPo7IK8gKjcHhvUEGlWv3A5
iP/uNwFAv/hWKGmdKGtsdgRIH7887fz3AZ0e84IyGCs/Mp5WikOU/V6vNM4U479D
KGxohQURqgDy+fgKIYE8ceO0s+vL+djV2Vgi5HJSB7fM2XbW90qwh44KAdwkIKYv
OMg5trwY0KflOdqOj+t6F/Yt3lmwdErY7jDW1J8Xi9yzjvsHbiWksBk0WjuaJHkQ
avSctt3Gkq5C7iJudoEB3Oywa7Imypv92aOjVcRE3QlDfOfmty4CdpfrOu97KcEN
D81iINMs5T/j+bE3AgmB2I7zVb79kNY2109qOeEVRdnZRD4Ne5RymNvqKWogpwxy
lpum2wNagk9QU37rJ4NLfFwVpEE2wVhZID+ltkLHMsBzrf6Wzlp4zudXi2NIJhRI
ruZX/tBQx4jSTD5THNvGqq4935nWPO9FEVxJ+v0RGUke3pUxjckuvC7BGMfXzrwf
nmfcqIriATuxC6ZqoiRRQY/mtoVe0U/jUYWU+U+ipT8NkKSJbdH+W84PO163HwXl
7wotp1tUZXDg1nK6kPlgti2kzVRwZ/Pgmh4be/Y+o+QeZl3YCrCRb72/COQJktyH
U9ZIzskNYV7jto4I7STtXQ5yccdffpZ9u0uhqe8ywTVD0Fm7dWHCtuMUmd6Jz0Vq
/HVk2XxWdQd+6HZJefIUm3qoLteHgB1CXNZqv9+vJRirHBxLNnsjG0yVSE/ccxMr
N5DnrS119w94B5flvIqD+OS1KwlfIUBd7Dh7NS0mubgCKTVK/VUUAi9Is9qO2jJ8
UVq1k9rNckMZSKJAY4NGsTRHOdCbnrc0BB8rs03aLL9DPAsdUTv9s9KDnoux8cXX
4rtT6jLCGHCEUFsmrGGrNIijTySnC+UJpWTxH4QQISEz+UM/AhwbXxzoBggiTR0z
52YVZYTbGJO9s6dWXUCHQnZdk0Xpm9NyTsmawzbUSOdWhlhzX5Tv8itfMUCdX6bh
16/DEPcWi7IYGGpf2UXPsFeHr/qiXtnOhiX5fBIBSi0ET30+1TExi7jUIXlDmoYh
c39TNFpcxVou5B2xzRSaYUWcSZvsXBUzYBLCQyaK1xylvQgMFP93UDql4gQB+A1s
kGNBb/ic/sKXEeIG5Unrr3kBfcPky8K2LaJJcehYzgvjgsRn9hFJyfinhC704fgD
hMoY2Rj2vU4bqnHm0lbE74Ucvd6muu7M5Lbpj/tNYPVZGwhoidYkPIOeSjxTt0vY
8U2guR10x34Lt8xdo4U6EL12jsIfVhwHlgAi7XPAvZQj865fLKI5l0b2Nh68HOHn
tnmGDHLsnq7/sQEPJuVPeyEXSjyzg4S+iEWQF6tCjfuJcgT45RXAXdaFBknDD4y6
qQanTF2eCM3z1UN+prSspUGsFepgzLH8ffv36IjkDXN7rVdFsM4lvU40Uh/Z6dYL
sGCf3vdABC8zWS0vRLur5lbQ5+dhoVpga7naDEThjrexG6BE2gQb3xzf9HMsBtWw
WcOVo0YTt9HPQskL00SrBJtO0Z4vF/1IfuKmPztkBoe0VJyoHm1hXYz1m0m2sw45
huabpNKLCdFl+R/X3uk+yIjnShC4276tpBlYt5sz2RokUOA2NA0cpTbvPvghy8nV
HvWPxrvB0P7wTFWcHcl9iTuouP4w/EEyQu9OGCCGaAW/PsgLwb8KRC+D1V52vvzT
CTj7W1iNMbbmMuZqEWwjXAO7Ql3aqgalLgRD9QNNoAFxCAs5t+8S6XKYHvyqQRrj
1REj9ynpn0FTwTqirmdTBGr7CO0sRprCYUrW/Bn00Ni6VRcU6VXcjPC22yREevzn
Cd5MgMHTKIzkh5NcZ41WULJptaM8Hbhuj/65hXqOJ2Ax20xP5CmqsGPSWlyj3wUJ
E2+MGgJA6L+GgilCWqxhoWIeX5Ol0vuqUf0kxYZJSxyZ9MZ+d5HixfjwtR8vKlTJ
QrcG2iJOiwOLgIdrmvj8wVv9iKIQ1jzRhkXhOnOVfb/7aRftzRA5M+L7bgNsLJAa
TYazVbXOjqOQkWdDUJS+Q4a0AMtJx5DcLrM1kB0xrfY1+eNiUvGFUIQHlU6yBAF1
r0smEq3Swmv828fuNB6FMHAYE2VP7z5+N8u4Uiu1qtLAPSI2+Gnx/fxNsuQ5VOQW
+b9I8AEquPgsqfkECArAGNQZ9FTDSoOO63Mh+Hp8WkOjX6v5R2AK4p+xoomzoKYW
F20SxL4GmZc/EsvKsQiFpoN+vkmTcvz0i/pJ9g5U/zXoZTdazPpYYmqVgHOF+cxh
VumJJqj9PJN6+E4+eH0Ir7uFkIeh60zweRSr/ehxNuhVNHxJQYwLU5XP3utFE5ei
SByyPBnWCSIxMcnuT4YMdz5CHDEOaCeUD6+uHDK5JyWWd5akpxxcpEob1HONXHyp
Gt02urZK9VL4o1VNNE0eOVku3GRQjM8EpewWg2kfqy936XTTUKAUbVi0pqERFZ3x
rHvcJpR4xl4wkAFhE7gDI6iTKf1i1kQmjLyN1P0o4fANTeD5xcOhWZeAQ3XtMeXG
Pz4bwhpKBmLLm4hErJGNaVGMMrluU4VYYHKEMk6M129CMKNKIJDvs9uTiBo0CEnO
Jg78o1eMGKzu8qYh8RvZcyyPBZNM9835UzcNPgm8bKL6FCxgJ24Xac87qwKro4CR
qs2JAu2TcUI4Mtc2/YGlRJpvtTHBeEGzm0Issa5nY3S65d4w46iiCGm9EIIRDbOH
pT1FTJyuyeWJyuKflfYi6qkeWobKs3XyQj58cz+tQtiTnme06PnFRjFljN6vBj+M
1QwY91d6UQv5fLvrgRZnBIwWjnudjLMR0BvqmoRPMt7lVtq7dFbGjMdUJvA7j3TP
JVI32BDv2f9y8Av7ipnHGfBIfqnhgE/zHph6UxHOmZSZzLI8D88rfzoNUDoUIUC/
qKO5uR+NB7J/n9jddrmRoh2yqoArwh3LrJe9JRuvBzYJPz1zDwO2ORPT8/gzheeq
V60JIe9s4+HQBTeASJW0x4LyxLEiRDv5aHiM2PAT3W4/K12yBzGVfdiS2+RzHEzG
DgGYPLL+D88RTzKQGMnfaN3905mPksSgpP4SdoQMbNR8hQhFkOp+zzTker9MUC0y
gVY3nAvLbCPl8/1STszusyNJrYLsNCB5clG/2118nDvl15ipRq2eXBf+tISmHMgI
ye8dm6lhfZ3SvPJAcZIJUYwqeIMUfymSlgiMaT/VBaqPiMMgjRAKcCS+oZcBOTAX
v0sUGWZn422ziKKjnecK+W3NYeNycsnUHIgQfgXNd4lOER+TqHsm7dkpMf8MHqsC
xQFkigXUfBEbCyv+JUz/VgO97FDzSuKQIcrT+lTVhq53RPRXxEbUB7vPUbPuedTm
ExLPqZkFBTzfOEV3+GtkuxmFoq/x4V8WTCbrVgbhh5N9SEohYkNG99UlxzBxFT4G
U8MHC+dOQqoNwzu0FGSvbYocf/W9E+9aw4i0IT6401hw7Y2ICowkCysNHEZ8V0FY
n38biXz+Tvc8t3TiYt930KoNUlj07AuIK7MluxJXDhqtXNvjr4zYpYN9iVaiyLFq
ludaYPIUxNwrjny9toUmUkiQB9FoZe6QU8cxsXMce8vRVo2XniN9+ejnlV0ilRQA
09jqmRsZiz1xMbgGZxCsehoDiZaXxdO9wg+zSNy2s7+27Jyt2y61MHQ1ybyukR8/
QPIYvAY/ms3qXcZzEpydBKPOwBsMhAe03D2VEvYJgJob/MxNsZdbslKfN/pbE5Fg
DDStOrQDXgKPKlTdRjhJnsHu5reyOheq4flVY8iQGLN1ZwHxfIf/CiKoH1NeG1i3
87ldx4g5hxSmIeKX5LcPEQLpuNaIWHVUiZuWyyXryJn/Vw3/g8Zh65vxzk7jyHx1
7azzJescFWKJKmglpSLG4g9RDu8JnEUVtFkN0SaY2uI5PCRGCEMRJNk89dCaFD42
0xAXfenAKXaz2JdnRdpozLLztZj+KChnDfQfysVanFiaGxw9ZD6yTzanvtxYD4j7
AIwR0x6YjVb3TapnwlNcqZj+iKOOgtig0JZzuZUcf0aisuI18Hit/+wsQDgvUtB/
GR3Y36635bfilPCzdOehxR2iXH3IecVvCiBmuHt+2ACPQf5pXqOEtqoK74AJ/Yu0
6+1rooTLJghTx23Ic7AwOBDq9ZXMtRdWouwGOUJU4LeYxt1DULfv3uV2QB1Jqvt6
V04ICDIlJ0YR+18mpEzYUGL98SUUcGHs+rKVx/PyhDsQkWdc7MBe9cajtymK+PD3
RXPvX0c9hdSyAqIZvZMUk9m+eEEaeZdKylb65Wp9i0h8XPwuQKpndcIy1us4ecDV
JzdEGAAAoYtQCl7RWNH59qpCpyB9dV2Fyi0IhREtMjqS8KllrpQelkoMK6CyIhCd
XhMyFnt/ELYHLuY8GKDBYdES4eYiXYPwPv0l8Aj5f6djTV0XuJSLDLtbuxxmhC8/
Ro9DPIcswdg1+5Y0+H2PBr7RFXygReJodYG3beNFOZyoGAkvwrV6JOZIHblS++Qi
tD/wLduGXI1aVQs0/TzIorBk3nBF6Niw/3z57LFfLOqIDedXiSjnswi0Bit1tqMB
sfyn0PuB89gV2CeITg99BTrPy2cCz2innFboC91OqWuOO/IqRfRi6f8f9X2+t4Gd
VfvQAAEjlj9pJdCTZMa1L5JLD8cehXIA/Fd4lm63ubuMGuIbe/vghIASCrho24/i
zAZbV6rX1V8Grha/B/oWskazCuEzaTV/gfwHccBT2Bp9hGqMaEICDWp9jA3YRukT
pynGOvgwRDj9DF43w4uCw464b1HM0Z0m0dxDsRnymi1lu1V8M1wgis74QScTtwG5
sNJ4++JM/GayvkhkI9F7IcUwdfp6ku/2moPhlEnFF7ZaS9wiGO0qkoEaTR4Mc3Ii
noobmhmc7KcPWG2sLrvmdsVkem24L0cUO/dq9/tygLfZrqx5sngMIVynl2B6yAA5
ckNBvLi6FCqXCbpPNXylqhqSwWs+DsnW9GLsZRyjZTMZNLHPLuw+enBi6f5cJ6za
YMnWtaTT9RN99FoJ4/BVqMo/syDbUP6u6rf9nGJUqsP3ThZJ4x/B65j7Ux9l1FnX
0MRMU/4YAdMmNDu/MT1woVZ1Bie701/TFI/ivbffqAHbUX6ZnQw8kDPlAo2egdB2
wZD2b+E2rPk9vFNvpITDiLUJSrX3CQOqP+vn9tQTyiB7TTgVBd381SpPJ5LTihLG
ErMZV6yK/t3BXNLR43/BB05WDoBlxNXzQaCWmc2PV7+v0tsPulEWkNgoIJVZf4Zt
SU+0sXE04owRZrKOAXK8PpmWY5tL8KJ0fZFAZhKhjX026qFXw35wgL5Twh//b9aT
c18kb/O8mbxi2MI1YOLwwe7k8N81CayQG+OlHMuD0pYxXGh+d3Df/U92PPzCFmKQ
bS9ZnHzMOswAJFca4qoB1g1weso/efGmEwE2hwffHT0XaBHq1tI7FFZyZLEALnBm
c2oxDUPXe3ZjfFBx5EQXzkFGCFne527wsK8kKkF2CowIY8HhlaGStyZAbfODIxts
JhalcDLTN8D7TMyy8pjU9w2tfls5jDuwugcp+wzOtAKePWyWsenXcsUNSLXQOFJu
Tne7H1VcwpkzjvXW5ccWz4ByelmE/zWWclE9QFBcmvbAgbs06FD+mgIWukQmjvYA
G0Q+P1r0Hr76aTIfU5Z3M2pL5v+Oc77O74mSfqbLHapHA6ySoD/e5Utc5GoI400N
w5LWLdCmlvo2GCtGR14o97Yf7gG6s7wyC2CWUirm7uJAOcQsRe9EZai9MuynTOH5
fpHKEW7/tFI2S6MuI7AhvgbExbUXf7cNshqynYHvjO3lDCRaw+4TLrKZ5M/Y8fGA
QrYkmJWoI2e0mGWJUlJzS+0cNNN/UckGDkNWoNVRzUJemQFCWKnulC24jZNbO1km
dI/RbacQRsT3KjP3vXPYdWme/+qtpkksbLXM667agfBWFXh0FOfsTPRPY8yepx2z
LTO/O8ARBBisKoe8BMDNnE7SrBYXiYANb8Kg0IfrpVUD8KjHL9XmYUtYjFNGrGb5
/TQB44KzZjfop8KrohXvHBZ9AAy06Iq1H1ht+VJnfATjMioZ0+YPTlwotN8V/1MQ
2IFojVrIFbTEEntHA1CxBWHG0EpvWcH/D0cUrISQC6xDcKxm1FO5TaPSv1O4qrav
rD3ugP4cMEvzotllqqAMcwWaB+5pOuVPMgP3M4UveSe6esJqhYckqAJiKA6aIhhy
eMN9Py1T1VkXICA7JyBCNPlcwXmAFCto1c17gOR4oYr2FqnUpo/jhEhTtBUWULpg
YnkYyyUcYPxw6Tw+FzPo3c9kD5cbpVC7LMxslv/GwrJSb3gqe/MGFN5uC0yNdfyw
IzpWhKoTy411X2fa6N/n73tDmb4zKv/waH361C8MbJQ4b3f9Wzn7x7WqjBd8g//E
mtBwlPs/VObgBwy7GOT9d8UVH0JfhvgD9oTZwaQx8siyenXne3WbesaH0W+iJcPR
rdX+BSHOKTC9M6l4l02WOYG51EjtFOR9La+Un8PRZt+nkRtr8rKFijTV33ztj7G8
STPIhdms9bZpLrjdi3emxRcOS4AKy8vysrOOnRnZ7J3AyfK2ekJ+ctLi0rSdeEq4
rSXQ+oRi3Uq3ybk7jSapYWqKpC/8p2QTjrUftm6TJEyHCTlaK3PEIepi7hmExTpL
imsbnNGiHRPzvQ3Mmqn0ZWV+RkHbOvaexaIlOGV0tgjBPGiI4nEqFn4jv/elciHi
OG4JPm9psMbyBPED2MOhToNPHGXD+uGQxJJZPLryoXysz0aV+m8Z+N3xhU7qUkGt
Xq4LgZy4WjOeNVVW0hm+/fS0e595gHkZrtJP7HgYS7U+IEM6c8BO0EKKSsPhzwTt
WvcVZ/N3HSEWQY+ScQS9NNFrNQ9LwA9OgKbJgrdX6M9ePxowYj/nDsEp67ohnV3q
kmi0fGdz6wdHXrRs+nwMYv+atLgjfstgzeHdcnMh/msW1OQSAjqW0N0wJpVEgcyk
iZlfdmik300axLCHvaGToBFkVxvgWDlWt48I1z7lo8kOh4RRNN0jZim0UA6/oa0o
3ZwoLLsS1EpGyJhftjvPKfZ2NyvHY7lNnd5dZRM5ia4HED/ehb6i4wh85ZOxW0Ta
ZzM56sUjzaZhvJafuSWnyvZ23Adc+jeNuR076covYo7N3PRCST88qvrhmPcEgs5J
8EUorjrGl/3bgLQ/Dp0Lko7U0xA2BhoN8u9QmRSsxsK6BZxd4nBd94saUfmOJDVl
eBrMUMT+VPdR2Q3BdwjA5qd/BgwT+BD92Ak2GspGX98ShzssKy5qPUPU7OEM9O7Q
32UWQrIbWtIsO+Y1UgSwvSqjni3XUXF8JaCZxbmAwEXoDrIX9EVR7tDVcixE8r1q
V5OoVjnL9YnsJtc37FhWpgxbL0cWixnCN4d4fJjpyeHOiaKS9p3QdEfsEso5LEqh
ZJlqxHqZdIOON8hGitQ27Hqd+L5lzUXkjqugsKQfqUBS/SqzdtFUM/g/iIw9U43a
pu2LQL1PE8HaEvix+E9tMsEmgtV1r5k2Aw3fup4mx3EFvW9e2sQRShU6mi6whEUa
Ej1GPTZs1XTK/hRCLn/Rg07cMzW+d4scGghJLAE4qUJEBr9MIWjDSBi7INqrI57s
uUZovcG5GQfn6BJz7hKX/7rT/iGgAoqmJRUGSL0NlhZ8t/6QvGg+qoJUl+I+sxcG
07XuowT6Juw9/2Hd2hVQS9bjMu4SCaR5q3nSghu0ZaOhkNa8ztKwevJfP71k4N60
zJ4Eo7oz+sR3QPj2Gr6kjD5DOXzO0w60aDICS2oG6BzKFhrQAzwQ+BHya6jD264P
KUVWBl8t2AirwslB6BVVvl0UFFRwYdRc7tJ8deIbaH55BP40QP6iQekhBLj8BWFr
tU6bejZGhaScZ8mA0+EDTMf0c8iZrAjbF5zqM+v0kaauf/wmnHsLf8RXu/181iuN
hbnTDTzvYvdhxNZfINrCJVzILXeuw0MMFLn11lJq5OM0NKrDi31S062FpYTsS1Qv
Oq74Ps22vNgXK5F6QibxXt/01fSPqKDxcHNm3AUT1I+kTld0CMQJ2zFwqj2igB0P
jg+fUaP/EC4m+wm3mNu/7PNH4WoWoc9xWM26PjGyrgHkYFZf9R7yVxy9Qg1FWhVZ
PHHFqeGRB/cZ3VynPBqLNA6BqaXTQOZKZ/T/2R0SJbC9hSe3iynjAHYt50CaDiRo
nMkqdCGWLJkg+iFjEzcm+b3R6r6ezoXyHNnwN6V3S3HMroTgmvA7or9/77iKHfzC
g/UPK+7wXxWBIJcvBmUExue5OJiFAc7hToFno/TyRngW1lHtbIsnc6LQRPfrfK4S
evTlcaJ6VP9nyIh4+wu2YLNpQAu3YU/UB+jv74RtfG2ZRurPnnYnUNa/wyzEpGgN
4tP6/vlm9gulE+b7Qg6FRrg9gqSq1S+wOAb3XzS+sPtPoMzfzQGPoeoBchnaQ7sw
k/kyY9omUNsXyWs24Iac7B7ukc88ypIMzmpOnFahzqNVR18Mx25pWCDS9IHNhn14
wWivz6I2BPTh1jGAhQ/vEA65/Rbp7ogg2givaFlCsDZRkb0iO4IDlrnqUmToAFpH
LNF1ck4GBAINUuXM9SbE8NsoLfz1ZVm54ZQRJF8XLm6MQwTawOIXBBx0Gr/mD3oi
2tC/Rbt8rN8BV/P9Dyvzq0XnoJV4gZGu7XKsfvbwduLFKMS72lpcqsL+zeCDxcj3
z+5pv4fe67VpRv2xNuVAcw/SFV0pXVTd6j9qwPLv5qNtdKEiJnBR/Ym7wbY1MUC4
ACIuxRG8GfysSWszUigt3lRGwoCPusN5u1kNAQPx/B0PBxkWkohJxV5ymgHPpelW
iKExnd1/lw5HyvORhNddMv4T9y2RXAMxct9Vx0/8cmHPconcfitFfW8qnhr4t6Vg
vdV0laIl7JEeObbWj7OAvd+oSs9LwolO4hh5mQnyb9pJzADR1jKZmMt81ni+Gw6/
GcpuHMAU2lUIn+EPvYURLC1lMI0bepzm1ljmiKOubXlddLwvLgeI2hArSm7bjkoc
ezREBk25MhdhJg7mK4gTbu2QiG//3Dwep+2hSSnRPfUIcHRrysiBOrNLVTU4OQOX
GoHn4RPXSPQ/Mk8q/erLT9vAgA+piJkUaVWESdt7CG8EQiSxWQkPrdTbVd6MTcK+
ZdBtRR7p31ie1zXfcYl+UCEP2jnCvyQt0qO/BUDqOXccjIiihvHaXtJGSdWwrytO
ayHtFsg5s6lmJfMD5AC1k3mNQ5AfYewSBuTicSmxTQ4gOEEPI9CrSEW7lpSbUWoA
cpm5VjnyUqu9zvqRLPRhVjIJ1r542ZSL8+h+XXcBlbmFjfP95ig67PMdDV/gFLyd
S/tb/vSnOdzjt7vd8oGB9/rvjuKbIh/ftffbda5FM/MK62D9Yir5OvgnhzxFSxgT
yXbnGGm/Msobb5yF+Z/ucznADnvatjMD2lunG6eiYX82wV8NyNwE4v3C7f8f7mZF
iwPze8lofpgYLjMtdviuaglOP0YJSBgrtwoMEl8X0ZR60o8aXzynbXv9WouGTBpw
8ukvPWZoRiy/9tjZ5LB8XS06bLNMaD0431riSP9OzAbnhO77r26jq7F4HsAo/bQa
GlaRFCAWauD/ZIjL7wZCKsr8Ffc0ye66qNzwsh0aIu/KAoJR271+E1nFkE0UY2Tv
14FYxMxloUUmPM6+7ssbL/gO0GvbyoUQyjVmmgHy7JQ6Rem+/5Sg2OAWuD722Z7z
b6j09SkVgTyNQSd/g0UbvZm+YT5OBFz0pCqTFSRGCQaF3XkWERqCzGCdXITOrOst
JH5p2Fgmc+WrlQwm811YASd7pZyH8CsvCadjgUqA6hmfJ7U0XgczGoUcmNO/lTRg
Gf1t3U6yY6KGScaZlCY6kz5Zc+EqK8d2rKDf9Fp7C5Jct6kTMMlUDPyfKDyn8D+O
U4zsIozoSqWFdrsm0cg1ODBOUkji9gndxZKW4QBf3lJkC4hBidHHrso/KM0IiwZU
j+2ZA3y1Aq3ZUWJ8ebHIh3xSlbOumm8Kvbay3KhmTFKP0HS/ZbgG8mQB+Ucfc6Bz
JCGqSwsfnQCDsjnV5pSYj7l56Cj/JqBRvtrA9GXFZuNA8PlfzrWD4LBcA0cLheHj
tIr9HLS3ibsNQX+ziSpyoq7VwxBjOY8jQTwYgMrZNBJRALQtpzyf0FTBOyQatKxS
Ju+dgvu9qafgJPqp76qs76ZxrBv3j2ESyOwL4RsRywLTwJUsjVrN8aLsqFCsKkaP
LZA4/P0gVD/zhOPkJKNYAiom2CoMRV18oef26vFypLFTy51xoRJZOnNW+Z97y3GK
BG7OtrabOO60RygSQwdGvsqZU34+pjAWsLcFB4roHFoHyf4xku2GR0yEp+MtYPtC
IFQtFLmmHorMXFVKA+zGI5fNTlVE1W94ujh8XZ2AQ173GnpoVkERlbhMqwjtkjcd
YhbGsLcnuTEMlFzNm8ywYvLHZcuZiBcKAPn7P/pFH+56nWhLpZOf6x7kJu4eCnmk
SPpVwwiVcduY1wVKJJOh+AykV0zNSSlDz+eDdNkiSa71ICWVwYcJIowdq4YNX4jA
QjIbJvnA2mAGRFaOfNavGJDCbwmL9s9xHo4gAAwntTl/zM/oiyLAcQK1OswZm+Yp
iXs9AXBUACQfqRV980Jv3vi1bCQqIrhOD5bz/jQT1kpRgbp0G7OFWbafCWOa8Pyc
0aWfHOxBkFW3vlXqEbYC8sEfZ1mFp+Pan4+ene0Oy5+iCUdL5lVhpymOeCOQse6Y
oZIqGQZJBDOsZS3ySa5ycgTLWNm0qcBlz3GwYrEjlDwMpLozA6+Ua3EhXuX9aM8K
YJDcyN94sSKnSHAfSA59ZiP6CeUYrYOWR9e7pQjSJx/VeiLYgcG7Z2m4kgG7k0On
xPV0ibQbyqRL9HfJ5R3gmRHH2bmi9oVzPbq4FvgrzE3qsZJGguZAO+h1/40A8MUE
ET1QrrvJKedZwzp5WOnNt74tPVyWA3d6Lm4nwqT/jc9UzrXrP8XE+8agvvyHZKE1
ma5+VIDWEmdoiXrPKMW76UKQdqpFS+M16PL8+H9QdZJGkgzaDxPJQ8VQpjpKPHkL
VZ/fZeWLsdyqZfGzfJnJI6kpmdxMQr7QCPF/sSYVkPEdCmLuRxHWwiLsI8hZH/YD
yaP82yMYOPdYHb6sjxPrPADYFdsk6H9DLmpBz89k2FZ3CtJUAQTBGWzGclU1cLwB
oFO8u7KQ9M3QaGW1T4xYT1JjFGKR/R5b8BP1xQI8qlTSoy7utMleqAc1MQdFe5rf
PkpRYahL/JP2iDXoTPO6IFay4EEN09jT9tGLB+Q9IBrSa5psCWszNK4e5yRbFjNL
SVnUnH1hqKKCyC567XmUZJYeUedumQv1he0YgcSW0n9WbFo6aIY21oXequAXwDb6
flTw+shoRo5TGZDm53FnxtaGrGVszKHLe1jkehc7riFuoLXwUXVr8hi+d8HBJqNc
aSSSA6gzmk63HZ/fka+xtF4BUfhdd7//gGmd/xFpSs+acOeU+oY8T2UMrnwi+UZj
5QzKuX7D7t9GTjLjHcsYYs91WgH+I3Bzr3nOlRrDbJAxZLS1nsgzQFJZMa8bvs6A
7Cb6/4WptUwOruMxPNH0qd4cnQAhglFySfJjYb0wI/PRf0BA4b2+qeBXCnWqFoh5
/M5rK1UxqFwZl6Wj48xGBybpH4B5K15c6HCSyoxB3Dcc3Q7f448LPg3GgONlYKzP
ptYC9LUf95zwOMIY/wSRquSmcfcOk3MJmTLtxXF5oSvUBSR3MF+jwQcvjynY2WHl
bPHJXHm+Ao/DfSi9O9WsSMMXJYneXehJw4WT58vzuB9YfRJQCSKAxdw2txbz4yAa
wtyLoagzXZd97WjE4F5BwwFYPpCMHMGGAw8j0EyZX4Ch86/nwDx91Iss3fRcD+R8
/Nf2dPutxXFey5AEwjDa60Obi+ZHHO9NVyjaIiCMY+qrcBZU+RwDh1U4h9q+UZYE
9XSxAd18CREZSuUXwRq0VEq5lABla21Jpc8ezQLrBV+dvI+EwlulZ1TlWbZpzEot
AqgIJ+FvGU8Rmq97DH9gpbIiq2pxfyXccLkTLuSkdCXMOEbT+D3og4iPxNey+Rv7
/BgZHS633XxlDmSET3ZnvR/7UEd9vkA4F2LdtPbC2p+IeG1bIUkGxO+Eg+8x7s2w
BrdARzLWANmo8p725AA6T1KPa5FNB4umPDpXr/PEbhiO63zeW5N+wX35jmZHlfHW
dHlCHxz/Q02bw0ZmEWWPqMuWvdI8g9DRv7C4ZWdmoWp5D40AWrZT696sfwC6BwUT
SO/G9ZPXXtqTXNNcwsfoGRwkXgATOI8fEZ1hkwGgAaQCSTUTyR2WL9ItU392eVnx
biaxteAVao3JlAOd0Trs54JlJ8oJehJY4Emdkx1vDLLe2G6FMFlAObRO3h4BcM0q
dUwCIhJ7xLIeQu70EGaHx1LZmAvNaJTf2FgDmhd69VUo0hRLS1UBaXh/hA3u3bav
I8omc2JI/20O3M/5YcZTRBY6RuZgAVs3ScJKS4a03zVBMRGMUtR6QQt/E+ZUItCb
YZFSlgFeqDUucUI+e2q4pWUnshEbGebPWlvtYZw2uDVcYHmqmvlXCeI0ZQ1l0aqg
L/kKt6diG3o/EctztcpkNwVIEWAG0tXrADGvagbGpoltM9Q5MPKiRoFqTWgx79AC
he4a5rsJ38tOIeyb1ds4Qd+3OSJpFmt767MaIzkc99iZcmfKMlQPd3ZlaFgx9TY+
ahEnZwKvmkNLGAaiDPjqYgun1UEujx7rlbPBjenmgn2FIIBRK8rj9r2FiyYFGpuu
hTNTd3G4kUYpF9DB49Nal0pokpOTvGRSBUuf3pTxDkQbejTlMW4b1TCcEIeiGZhA
Hn3PwNTt1A0kTublxq1BAOy2ugNGXFMUV8WSVWNbDYCrJcKOyelOQLZ3JtXicoC+
g2JY+nLBIj05ucbaiR4AL++MmBJjgURPzHvvETPTIRdWk4fEp8e72RAbIycLuhlG
NHkWXEw+4Ze09/EYIT1+18qLs3YkYmZqylCbptiDv3By6ItPY2z6TyjimAggHiLb
jfXrVpGgDF5BYdt29V+yzGvpcWRmFAIs9sEB8gy9cqHY/JswtsKJqYIre/n3iHAS
u+EKPxNhkkLXn1AkEn6TtZZZpZFUYMZp3MPe5Q6cKDCHBRddD8HouFH5OvTgu/dK
+7e5btTd2UNgjZh9tQ3TrBrv/XmZgGFFmQ7Gxm5X+FKmveK0nlton2azw0X8MXyC
WIeldS79NBWOgNBOEkb0tHuTU3wdI6O6TGoqnBFQYGDiIk4KfKPByHq6dZpUGj3q
XrE8NEZnUerNly9TpYMYbyEImdFwiVdWTxrBxB7AG713Yltkt8z6jC/MMgpEqa24
C8xYjaqDAMnllzNCwFYkFc1OjrMA594J7USaVotRTUD7sQ/nIKj5Lw7/JVDCtMEL
EYcU2z9L6QeA1VTuJBciFvXSvcbOSyQobJuMHzRHP1a1wZGBYJvE+70Y8AQCeTi4
2ScpU+TQlZTOIR0T24qV29DdQRD6GRrxUEBhdJkIaho5KvHz1yP5OMMsUzoGTiNC
HU1iSB3HUvC0ULs2Y0t+Cv0i8iX61tg4I9hTKTCkMRkrc/jD6cdAi9ZTLLbtXUid
U8K8Cf7aK/Tz/jK6rkCri2/u4wgeG4WJPIW+b4aXBFV6BvAGfgSRG0o5TYjnXgEM
J+e4zwd4xwc2DK4vRj3NC7/wFFliU3UjnOk/QJY81Oaemp3UwLN+MoL2JS2Qs5hd
sWhNboyth+GC0vC04cSsTEa6YNYw2aPghEZPWh0I5t2Jg4CkIYp9FAsykAJI5L2/
cl5gmRcX568Vh1ZWZSMtaz58b5Aa3VUke3hgY7FOmPGcBtujcrA0HVPRuqZwpMmf
Ceg3MaMtg20Y5En68QV+mWmICX+ZaQKit4ne0EV/7bF98DsQlqrCDx2c/EQR+Zob
gVIGI+/GavhV+3MXJ10q7b6ra913h5nv+0pqnHRu4jGr+QohT5eolKk4wdaHNGux
vEJq0DjM+kZHAE29/rp3BmlD8WTxOP+AFMMLBQLSqUB2zDefrUlgdKpF4J/UTNiH
HqIydDqd0WmjRgz6VoYFP8aYvtHcYrd0CwVCekkHOx7620bWkURI6qYkxfoprfnh
KpMxqK8lnYdQIcZYRgVltWL91aPY3w62RK4XYBCnvJLWtI4DVzYUVTXJVIEb35bn
nGtff0q5+diFQvc7mwJasPfdE1URz6puDNbGj4HQg4sRsWPtPTq7rpRS0fJGgUuZ
MWpf7H83+6NVfeKly188kvl6zPsqSYYhGECBJHED0cB6N+kiSzPW1c7PbFWdfxUu
IvcDpZ1eoeELYuuA00OTeC3wgXm01PoPY/lJbquUU1P4Pg5ZvTBucbvBf4U4j0sf
DAA/l0wbcPnpMpHRmPc3rBq7EP1B5HmCLNEmwbDwJuK8hVsUG+VsCwGFSoSCqXdY
+/xIqRSA1r+G27+YBq7g9UO6GHZ7hIfHkH5rbyXiR55MYdSMkmv2o7V6biloWEfN
wcXcoj8NcR4kX9+si7UxDVp23pKDXY/8K2hy60tk6Lla6s4Mh9Eii5cSNiWrar9e
lVlChbmjEWxEzUVQOvkDyLMO23g+O5weC3+Hb54jrSaPnLdybgfpKZQBXe0E1YRd
AmtxjvBHzQRUksOh0gKq7yhTqxQZ6ERknvt/0h3jbNoAuR69U/BQNRKlRkxEOOq3
myffKqFL7JAgNjUAa6Lvw0LX6Os8J6VBRGhgFfj29bn4uaWzTRA8SC6mr7d9W49b
89xAPVfJb9nsnz4NoNCMcWGNbb8/EIDxls+vK6/iEApMHe3jr55GcMNlABF3Euun
1TrU7OQzwCAvmWGzVRI09yqtGPJmfKTqYc4NPuVQGegPZaKAfly0WVslTbjRoGak
rIE9lgsRA/zX40S5R4T8U5IuxKj/nbkuMARkXzj2WaZ2PmptIYukqQteBd8CA2gz
eQ5eq/XBNdlaw+gpST0Yce67c6+xg3dYcjrcJ34euAmHqQokdiEHOZDkRQjjy90a
HLP4fOthxENGoMRTGT6Ti+8AOII+YkNd3e4WWk8x5NaRgD9idYSsWtOvHYIWbCoS
ol2m1qBC0kMBnIpHn/l/sfL1GGj8wqIKtg4l6ieEv2zrtzgAgOmux2hpbC9+quTC
pX03ub0pyGYlbiywNTwvvrwQzNaR3O+4WoJbdh0Eh6u7tKy2XiaR9nVZv9bSfATi
yw7eCrtfVUswRTBYN2alemwBRK/Lmqqe24e39Qh0qZ1a1FnSnZpzzo2i7KtsgQH/
V6i0kldPJ9+fdUm+GlpIRGIs6N/J5l9Nkt5s4dO+SW/M1pUj3VJjhEhHcKYXGY6e
7jYnAS1i103S1P+IbEGm/ZzV71RHTuQK0GNRMSd4ExGmdunvyWDp2b8Z3/MYBs5p
ZEyPgqSouBRX9dHEM9Kt1inN3NuxK4vura/GBAxARAHMaidqSeSXulsrwxjk7jDX
vUbpdncSZ9W6pNSMy+hxNkc6+KtC8lLOckTNcGu4C/62YKkKtvfPxxi5ksFHeecs
iDrQG2hv9zHjba6zaXrmOvDv2mQXzRfDRtsLx5sSUZHJPiCjMJLfPSbtOW5zt94b
j756x7r2rtd4431yJzcrTfK+3sRAUoPa+3iGVPXpJ5yp3OkuOJMo0cC6+EqvVpo3
G8EcRbcVL5RmARSPoQukOqfX8AhpCDbBAFryZxEmEtmu9+6z0XAYt0h2ZrHnzSN8
kJzqzyBTpiHLybUU1lu11Cs4Gtw3LXWyxzcQAFN0Ll7nOwsd1Ddj+cT2G+nF4cvq
Uv5Jc/PSIz/21y1lIYiGe8YQNYOrHurXtNbwoZqp6hmMGoLxeY3bnvGjslGR/bP7
B+ZjNSHi0ZszzcjC8vVPlAYwc/qntyL0p2s8wtSh/AoeHI10K6OTzWTmO/me7oOc
yZnO2KeBdftLvHJgPhmafuNS9SliIEgsWEm5/HnmCTGIJ2hnv96BVDAdrMnhQnKi
OXVo6SwRqKNYrmkzLokU+oT6r3hDu8NAiacByvdxk2h9S/O9UaJK5YTWRYoKWCo8
mmm6VridcfI15OoctItsH5DYA/OdYvY0+1D+1g+a7N7fnMQfvYewQ70WAt1O6w5s
CHjCGdSPNK7n899D5Cgc/nJBg0H8vZcbqjAYtx2kLV1baopvjMuYef63UiaadIiM
iAJ4Mei3Hk+lscjqvVOokIIqh4EJOps+dOzB0lquOxwyCBQ/FdWyzdq2LH+jJXHJ
N9KVwo5jMjEWl7XgYXkBoFhlfzrMyqIcbjX6vEezeAlq16giKtlmopWb7lcbcUlJ
BJaJfS4MBjgkXSQverLRnfRLOBpCSw4rmiTIb/Y0gkTDjtpp3rLcutrXyKBsZIDm
H0DNzl2jGz8u1o3AHqpGGYuCB3H9e3xiJRMsWWPB9ZEVGVop1KXWZ42Slqn4yjK9
nUzY3T5bKPz0+CD5OGY9TuprEhowCuJ5hOZ7lY71rWedBXZUw7xZY0NqQnkxNSTt
QVbLRR//twyy48U80/Uz5tDKcTU/8VNelDopackXvuspUmkzXYPPn63jCCRJRxZQ
xVa4gpeAL2gD0iMmklT4PKzdGcW5gEKEYdxkDGLf8P0o+x1PR2lsgGflgeO2DUw8
19vZNMxlPeQSWG3O+77PiEweUcopyzESc2NpQaBG3a9ePYYaScCdBFYpvxwL7Da3
rg5UEhqLr7sh/qqebQo7CFCTF+qdmyiFFDCcQbylXh2/I2FY1h74mHRn9AKgU3DA
gykx+Lgk+7beRFjKtagFLNTeimXiqR3mq2c+Y38Uye9ur511rBFrwhtc4O5+fk1H
nZgihqyymFqiplZ4CsH6ygxLpNqwED6fkkT0I9YtcrO6aB8N3Ghz6LucSPkQm3xl
7BCfV4dbOzgFektQQVK2osZwGwP/ydSpuKt+P4zt1/v96x/Dg+hhyGd/8GXpVHDL
ZizTr1K5JA/xH0JF10Jamd+Ku/cUuK2FoAWwtsT1EDwGa+v11DYkkUEAXdVNbiFs
XBRJ7T4NbNcmuvcabFZvAMpz7P/JjI0qhIg0UmHbOcdGMEUwd1cx4q0Q/jSuW6VV
RwY6YkbDHFXzsXK5FRNTSTd0IcekWqN3QhZ95G63370zu/AVk8/21JdAs4vkYdjt
N4lHH3x0RES+14USAoc8Pwjrnv7pK5ob+TZC7ovLg/c8V7g5R/hra2R1sMnI0FIA
CqE25tIDxGclEQsXuzPi5OuJwgK4UIUH5b6cBVe+r2hjYaEt25yKifDxvL2mMP2n
V9MaY/E72p7QdAu3RbG5vsZnp0BHuDPUi6V7+FVCKMQGTUFgwctF8ZasEVT18hn7
aemonbwdaFLwPp03hZLaUR5xWR6KQGnGW/mMZNYS3dpCdDfG7qcLkZeyMPlqW4EU
q/p3vNBKcnw0TEZOtszxdEJgPLZ1keLz3+4j6GN33T/E367b0VOiCNd5Pgl6n6Q4
OKEO3Wl74XqouMYcJJsreObs1z2u8RNb+lVFjF+GzwaI31yQF15Ga30xLzlWBP+k
vpp+tKMpoCbKno/0F4vHvvYSydWn7CCTKmrqkSNk1cM3nTTIC3U7if+f8GUh5wxD
Fv0lqDfcpYhbkK+0kWItB0VV8SXkb0gpP870hZKdf22yQEvdmlLvIWCtu5bBBViM
1UBxvvA15EPcYBSjxmAVSx2nElg89IXHFVIG28W7Bi0ShRSUj+StZZw+CxHmzeUW
ZWbJOMJvqe5Gw7918gUEhSR82Rog/V+fxg4JxgokuxU042OHsISq9a3Pxq6J2ZvA
P8qOBftfFnTQ9IgXelunBgpecUYF1v9wha3ASUWw1THaiodLu2U5HvyscdN5r+Sw
Q0lo/j6mEB3KY0X9iJ/SJaFIv2kwnWe+y/3zYt3Uxard9ICPo4xUQwC30mTaKKSe
l1+QWhF3LbPyqxaX+VO5hOob8nRArDRWgsXgVPcvBztipZSwFp9zGWjoGQWet8UZ
xtWAxQkmYvyW4T9hkAReNFNS3CROKzW98jiugntwow7TQ9Qzdc15lpzi9Q+xr1Eq
wu8u0CGfUw78VLwzD5vZqLUWcPYY9gUCJdRXBAt5vOosKU+ufg3ILsZh/I294Yh9
KlM5zrlYNa2+QH91zXvKni5nxiMhlGuk/eCCXwIKanz39LtXT5QbVtB7B+1T7LWO
gSBk8d+2GhBqhwxR2c9VI/m0HoycNRWQzG8+yztcfhhrCkpXqMHSSoNXzL0myEs1
9GYtXE2zO3/zCU9LsiZZuY0tIF+UpmkV0kg/uwbHDG9s8iOjl4kjeJu9A4VNplAJ
YX0/TLrkoiYTmVDIwsMWLypM/BqGj7dqpv82eP5tJYvvCFtLmc35iaiqTFtBFKOb
FPLFcBg9468wfmtz5+86YiqPUYBol3HUytCIyL3LscpRZtXzTv1ItZlKQWnFMbcD
CJikuSfyghkVWE3+68lJ3vq7uzbE9hL8BYCpEohXlwsXr+QAsvth6HktzjQNVGzl
Ks5lYG5ecpZnL2sizr7mWFLdm1gnaHQDcf4eW0gkSWB474jHRoR0yMWXLdS6JzIY
yj7yN0V+oXSGfTHrpJnIap6Gj/ArowQ3eyythcemy4VM9Y0RciIVa1vKpTtprixG
SSxa/J3H/yaG+jd7TPWjTeS4inB9K/w5JUmNU6sflndYWftlbryddPHWBgL1PtjM
s3llj1hsSYP7pAZz1I6zSs2YdvaublSztyF8cUMn2mrk9oCPuYMYJX3P1leQyxO1
sKC6EDh6roYAPRrkCibO+dYIOde1rLl6mlltob+NYnN2r4lX89/F55g2VgJs09Lv
DqMUN3ysfkrEWulGjyKAC43LtUnMGoWIzpQx6KJTzwVdWVRA1/RvWnSmjL2+epr9
w2iIfMr7EtNNxOZUMGsicWH82OuqQdlWkXHaiCjmf45HPYBwxFf9s4cJku3GLYLI
4jiGxFzU0k68KwI/lshwweXJx/SwvI0x5og3OVaa7EMPQQNCKRZCweTIxvHxABpl
vjg51PNyKY/w8C0eLbQ+R8XlTAX9qQW6M3O9o8U3x3UtOvf7+ZeFmIEDV6Gzb1O0
YFsDpiF/kxX3djQDFeT6mVK5nXxtwN078xs488SBDqIn2ShJFtuEqETKjPObdHIU
qwl+jtgbe1Fv/mYFEIz1tIZhHok3P0dFMVI/+wNM+06qLQXWcSWMUQMnPDI/kkSC
XAr7Hzg2mtVFjJBiKdXN8T/z50trBCQLAZ/iKVe7mRj0GWvKKVmhr3yKdPmjC8cB
MclgaQ2fzzI63YQDgiroTxVA6bgodgPeMFNa8o+lYFKo0mAVr/ILm9M2qSuu5Jtd
3NEusWWUPc05JyaRRpsbXRKPo6ay0vUFOMq7fI771fwVq6gpQ7aofvhrEe/XnqLF
sJXiZBdZnth+tEbdYcAocmhp6ilpQwRV1Md9X80NMJjAJpw2zl0v6SffpZl82hmW
Lr42zJfheAcThFQs/ZSyBI/T1ODTclTGbwWX3Xn+RfC2ch3VF69INf6PTWEhvfCF
aB7FdAXMYB9t9tc8Wd7fesxPa3c1VLV0wGNvjnzootQa51Rdp1FPx47E1h6bVyqz
1xcBJy0RZIoT34TyIHDhmWjQYmlut7hXlkp8iakXgLXXIAul9WiA2YK4EAlASkFG
FhNvqajHS4r2HZl/zsoV82kBPdCylbH/DZETAVNDPy4L25HzvE4Sz/WHV8uy3b9o
9re7p6goTwyjnPY0JDe0rgi3K6XohojVoru9nAjwhGm1wkg1fJOzrA43cWeofKX7
Wvp3larbO2dZ5bnEcXjSh2qlIlc/pp5vD56HAgJ6WZj/iHwJzSIWaxa1Suc2rlXh
KtZuL5XkV+7jYgbZXI+1WHkbIXSbGNBLiE1FERKAcrfOWOnVz0+HzpNqvUf83Bon
oopdtzeo5ZLCccf8A3F719J72nulYvEGRWIR98V20/pmTUcF8aRQEVYss/aqMyNt
FV/fY5uVGmFzRKDOwsTr9wF87Arfgx9E9pu2uhr4SQ0C/qlaq4MO064X2ZV9f5QC
XLIuMhtu2lPzv02upCNGelhrPL8Tj4pYxKSFfv0DTqV3C1yQVARqXq3yfFuEO/j1
oXskeRG4h7aDYoj9oiwXRfs/vC4QLoMVL0o8KZ0MtQFm4l6FRQ3HceBPeQXDLin4
qWn/c4zPEAXR3SB+6yQD4NZgug2dkQd38ZaSNwVO/2+eFrwn7bYs3qe4lV1Bcbht
K46eqAIk4uk8ZpTJA7kxJh7mZQOWtJ5dYbforA7I0U5YDaAYVuBgmsW8vdsbExKr
DakRtELrM86eN4OFwK88TUPYGigutlwCr5NTC8O4RZ2MecYkNLFGKmYnLYQl54Pk
Y71VOn4cRD8ELpt1Q1OFU8pYIRxoquomBXQ8e248oTLXgFwkhFt6yOB/EfJ8xLeC
GuFWK1drt3xfjAcDSBQZsFG24IeAddzkSFC1hOZbWWH1tlCbeCJJoOEdyw5wmQzA
v5dvzk96rKExXPFka3za94C4TrYKsfzEhvcRPW0NScxK5avNNFsHLF1g8IgD6Y2Y
/u+wSqWGv56NrbtHk+6bQGFhCJsXTk71NI6Aax5Z9+Qj6Fcf58r8XT2R56X4o5Hn
BPiOFxB1TsxkWsFENbrMwVD9E/onEGLM9MN8S57qCiF25wnCCrd8FONHFTEHKhBQ
UhiEaGhRbZww3r6w7F7odllgFp/MGG4YBgf4cb78PPNRf32u6C/0p+0pkpQzuhs/
LsFHtEQdKds8uixo+Lb6XB5sc4xDPy6hUVSZf1yLvl7GDHxRKvL5ff/0bNRjeW4l
AJCHc16an4rcQo3C0oxaKtCt+rfbX23leMfPZmCq2lSTE5U9iXEjAVcZpS7GCMy1
bfF+BVPaLa6gYn+tkwA50ZApQfV3MiOE2oi868Qlvt196/bg6vJkwLC67GYdLzLn
7QwW+XZ6FobrkkFRKR5FUX5Y2OX24hJE3cJ1mFxagPrbaUMMFPvFhE7rmZ+ACYY+
rHUBlorDPkVzXkBL4mXlndcpumstpUCyOmnEedyYJHmdq+Q0jU1VAmxoK/xJjsBP
aXNrm+33nW98oW/okgkcQZdtSCsvdM227UtJ4b+P1d3m2hTqVVkC5o3EJOkGpx66
Xv0cjEpU2zI7nriPlKkJ20MrOOHvWfa3Ydwf0hrX4R95XySKic4s4s/p8OiGwrGJ
OX6A0kuvgVV43zusaZsfk0ggt+/RIuXV118etkDoHUff6U/m5HYVVsk9R/jj3yoH
J7omrWxQ0In/sRvjK0m3Knql4TOQLKMR7mrdj7k+lPYg/cQhwl/5Mh815RTB87FR
ceU48iSGlpjofal/jcEhWE4CRTx+I+Ae9D9DUOcsBtAq5UmO2JjGBBPXb09olnGs
kGteRD4hVTl/oInrO0jPyl1LBTdeyyoUJPwa0Xw1Iy7OJGAWWxt9zlalAInX34ZW
3CUAGq1d6w2DzBkUyswHhFxQzkl9XJliOy/lOXWfys9z6+hZNJpaXXUEmNS1aMsg
tEUB0nC7GM6PdwyogGL7hCW4tkYGJVaShU0u3FHNYy7Y7f9ejeadVdfEaWaFwSwp
CmGInYZdfe5Blc+PVOgAaNDR+bncW0FFDIuv8i5gUEb7kngw0I8Bh+THfnRWtM7z
p+RtsIYYpTOWg1uLsaO+BDh+62PxrQGf1guI1ZOFvCpOD9w/DXCpOR4EidBt1m8/
H8OnyYXQPvwi760g2n4w6tBCpdkfBPhUfkZNjrtSzUj9l9JKAh7yUZifsGXoOzoQ
CIrkYzPYCaSCc0YaC+skNHSGcx+uKdhCEzrqMEhgqjr7GnocDqPMWwcfN+BONN34
odMZysRUo/ZLQ30N3YBC9xFtcuRdqUaul4C7W+IomacAf2GsVIoj+rI0ae0AUHdP
nMCiFTMetTqZiIGt50wyvaKu2BKtAVoKgqtbgy+Mmhl04EhqjZrK+HH5vLaw0MY2
2uCnqlXbRbLvT5zAwcTkU3ht14QBqIw+t2QbS5DNYK5x6CF184z/r6ZUsZvzTCbq
EKJxRueMA1SY4OSRZHO7Py2oVjGAsTiyaB7X4QseaGUQ2apZARzY2tUuXmJOGQ7I
v3GkcFrbBmBLnEnWBvWRRl9jTAo8HTXSZUQwGG37gTMCnBpEu3/Vl4J8Xdynj9ek
dXTScWcbKJdZ/Urw0KQ7GX54ufDyEO5yOAW+gPhAS9cD5u9F+n9vhedcx0ucEi1d
pHT3Rh13sjkqEUg1067jG+Uco7c5fCrMbP4IomMlFWloX4EYmgVHQfU+2yGt3v8e
7gloNCOrt62qfsi6YMiwKIFxcUO36mAWNVKRRH+clgyzoM92wsxvaXlTR5HI04C2
giSn6+jlcQKCURoLZZdM9P/FFLk+rWLgsDKSfdag/mkoqToBye+ufCkibcV8R1Dk
Y6q5pMot+d08gFVClG1FMgn3u5lYHOZlg7wkojvfFNURu6gXrd/10tOOgnr6rThh
T1qo232flpZTSnLwqOxvNeh/eEsvWH6lLRTnpv8ahRNmJQI7KIeK+O/S/tUpYaHL
dQezPAfpHB4DFjujV/ZOd71mDrqI1W/Hd7cBjrEQxeI3Zij6IoupGXdF0N/atzJO
T8LKbAQGRnp/hAIRvi0FD3MJ6i7lo0lvkwQd3zTtFeSwxP4l3ZvhNcwSH9UoLHFB
fuZ+IFzZAfatTdv6XDsUlI8MJPz9nOxKY08SbUQP4QSdvV6tLUKuTD9OKeY+fqgW
4l+kAufKWPHefZfhnVOiFUq71Fo80fg+ljlFd3NW6TLs+Wz1aiHC+Nu4Ek9krpM4
xV2g+xrZs50gaJIfXvCyp946o0IVAAc7pt236dNa+2pYnciRlXJN2L/ObhrdN7s1
DSWakI+JF5rnd7wGCpLAeGTdeKj3Ho7+oA3j+pLe5t+2ryChUCpzzmltytUfAsZn
vjfTNAhs9/25BnqoT0dhczUiYCJ1/DLGxKpWcw3VGEuNG9rduaTjX80qaKZIgRen
q7jnY9sAVimY+DP6bnEhtvSinMl1kkvrXbBqIdRObsA08BdI+310AzvW7RLL/Koy
HX4FwP8jxIjJRz1SvK/oKhWzhSu5zjbJi0WDSuY9jkycloL1G+P57JPQDJ0m431u
R8qd8wwxrnuLVnlW7euNfdiOnzvD4noFMgBMCGM7Egs6UdjBziEiJR5ogg9nt12S
owU1QUMXThxCZJ38lmhFKCvYaDXfFk/Yuy6rHp/H1ktRXciEILY/tx7R6+SUup9F
nV/dRN/v6TQGTP5NjS1RL1GJM7iWWQC7bnuXM8PrViZSAswe5yIrOmoi+g8ozdMB
vclsp5CwUaX4WbpFppY57auNdtgyDEXYiF0BC3a5efKnxOErU+ZOEs1o3L5fLwuV
2MDzRf5Ey5kKSpDa8IhF8SM5JIzcdg9Of0hYgGTFJxsK5cnogfp7KdCZ2hIIqyZ5
thyNc1/8k3A4Ims6FGGLkEkFpY1jy2WfHtxQZEJfTI2CtH3DJ7sGEU1GdkHcP9i2
75vdUpAvNX5deDKlWAhFqhqfKeq2t97QJVKG+NZDmF7EHDAkOITRa6Po3c7O3qY0
Kj5jl2WrRmtLDDkX9f3VAlB0KS2chhguBiD52TYw7Poo6tPtvolcish7GAHBx8mn
WnpZBC+EtCL97larl0qxGCX9J98e5i2jhzMcRq9nP/CvLouUkwKyQknlUXE1J3y1
PVbuZv+JM0t774Kx8bhHfoDE6OOhHVkjuV0XJyo8T5xdcsnyNe6ZLMeZMVXmTt5b
on6rxZJSjR1UDbcjaNYNYi4lSiDuqJxjWklFsf4DGYLlKnYotprksqiyLsjACPzV
cnn3yz3S1Poe2THRu13g98w5td+CUQK38EM0Zb7fsZQXhKmH+TDcfoKHImo5FwGl
VKd9f+9i0gwvYyz0SOFJC28CR90xqELLJN5B7G3HYGFcUZXeP3DCCb+99TvjPFHA
kddKWb0q53drQltdA5FIYeZa/YP0dayYfA1HdsFRmpJc7RwrSFlItMHoy7Q0lJ0f
rbVBFKoAMV7nr0vwzZbIDnCQ1kWt/msibJqB+1p8/dNkzlvxycFqmqTC+I+oJTNK
9lXsWOC4Moca0OSUZQeZ5fY61FL94EuRNa1dXgzgvEGMFDKxsIDB5rz91o2rzazH
l0dwdvHxHmeYIEP/6BtW+wYVNC/WMmekoKKkzT23uzMpC+A9s17Y5EVmPSTuR3Lh
sDpTDhJbY+mmQYBt6HEMEa2jmHIdLHH5/4hC+OV61sl/WmqNy75I1wy9HShqkeJf
bbUfpv0B9ehnLvigseps1WishQjVRmR1TD0wpNaTtbiuaztbdWHsYCGKHgZYqVY+
9WUHY2PvssPcE3XPO6P40oZZ/vWNm5y73RoHd+pr9qEUxpCgHzbi4slEMNbbmB6d
2rLQ81bihWkwoUE4stB0aLDbun6DTRVskA5HP3yKhwoiZxwvZHOMWFPTDw6/zL6+
TwQsRVnWpA5/zMp+K0C894KbHD6dLtivKtL11JvxuyTJPWShf9B6AEYvRs9Zwewd
4X1ykWcyVPcSpp6gDB//uL+cFcSdsZKDHOaHJWg97CUjFUCt5jOPXIuvigvc2rkz
D713kuW8LjdbuyfKd1Fl/IXgNrTx4MMHU3N8uc0Krn9V/MvNFIDnFus3pyAVicNo
22P5m1XHwvph95W/46mO6XUDZRJjI0njxK/ja0twGAdD7xBBHS5KjALMZy+DZXSH
PjAWq+TcTxMdnF9LFDln4Ou9dLx40hM/DnfV8sdFijoqN3gSyt4OMiz/KhqtMc3q
VV/HrcGa8/xjgIz8vHq91RlpKj4F34TmX241AB5WF9d7BSSxStJDMaLhmC/1oLlM
c+jzyMvrOXgAR7CLYMW8gKZT2Uf/Ey8KJs++j6CT2cJYHEDI80MZ3Gu72uhIqUAi
bX0G7dhXfZZJ0B7M8DB9QEkxMWGhs04a403jgmhVmvGHB/JbBNg7H/t/+eWlyykC
+kqeu36ct5vbA/K6C5UOPUl99a1EBgVtKFPMtHzT/EJkZLNBvFyzDBogTGIkqOHx
Iq7N2TjDs08AL7luqeBw35GqTCnv65RCFo36AK6lQsCXM+6+mwtXePb0UgmymRqG
1I/QxuTqrWvRkaFRC4Yrg+szjVmwEWajQvXkefnvalRkpUpkfuaS1EZ4u7lkOpax
ZayKoyjI0AA4bbFyrYUJXfOuRnNa1X/9wQjq7fW0fqVlwaYPvy28QZllE10d+etf
GJXCX+UNeJVNouTBxb/7HqidMhmNAHMu+OGURERSytMQzaaK8VeoItfgiTkVjiD/
mWIKmhBvxfZ1Hr+G0ntOkoVaPPeEUREdKt0ocyiRyqiVo1eXZCKitE0WdTVyTiAV
w7Or/DqhqUI1j88UdfUnNUjP5jyr74IpaAzy/aNulr3bvNktTVUBYXfxm4nMvSLc
0EZsj+ZIheUVf/c+VyZdFQh4le5rkRqqITEt81zzflvmHSj1Dj6mtoxX7v2hvA/m
Wkd/NaActuGhM3W5+ScJbwG0OQbUZ0HCw27LuJ3y4SF98uZd2U/PtNd45DgQhAPn
WTiwr/DBVCq9sv+snbJ+b17/pqPPG4HeKO1Ux6lp0zR+zCvXp65ukR5XxNsrhg3Q
1+Nw4bRMPgyDsB1vsmhy3qM8/aT6Ikf4P0O0vWrfAGWHKE5StCtUoOsuozdKWala
VMQXCTO4qmAfJhK2TWnG+uaM97iJ5exlea7P6tpixqQezIJOX07oB++vNfPw+1cy
15Y8KmsnciNAoXe1lTS2CNvd91W6A0McR+rk2gKyD+XZxRgZq1H5Qjhfn9U1kigv
l50S7tRE9Uk65tI/6ixgaXvQR+nzWcBVIoaevEWajdfrZZGwh1Hzm1NJAnZqGCyJ
pJzDadPJSUKIj/Zag8Qo4z2bg49Ft6VBLxy4IydiJEqS22O7G1fUKu0f1YjML4XM
tehM0a/jE+I2eHaZvOF2GzESDkDSX4QuTaudRt0DZ2vXpQG0yvTMyUnREtkf3Eak
QBAJPTPSLGSjKAxREYwVfskZ3Kj76wYYukiBZ388sCCefo6buh6/2avo+h+O5WE5
GycJNZ8Gsj4pTXlcAlJkuFv37A241N2Lq87159ltuucfKYaKF6uod1Z26wiv4T+p
tbL6BiLu2vyntQrc+aEequj/nLc8buTKqAViJxL0WZHRyXpeLVpEYhOVLRsP+NLp
v9692yM2A4rdNaKoTS0DZYV4rtGQ0wkEN4UAU98554oQ8BrHOxmhXg/eo/XLeenu
H8BImfDEqyU7Rvs0FV9l34NJZaUhr++1JgJQCIMSOGS15t/Dq9NdTt76QfZhalYk
pOyaYhwcYbj40uVuK+m9w16/frW0apAuQOFzpOKmtCIV2aG833bW1nExkSo4mIaJ
2Gq/gAW6+pjZg16jFOCP00/11JZAA/DDjBJSHRi3hfd4rSHhySCokn2Ycl2YHbYW
hiOoKURSLk9hvFPnSuLDdkuy8Jmz5W30bD+w2daxKl1bB1fzC4QZbd4Ozfjj1MQm
0PxLT1nQfWGolAcGtlPvMxQKFHn+7iT9G2i/gvD0mqJVI6Iffn2Geu6KhPm/fwfK
WDAAGCmiaUqtwOQizvZfjB4yRXYs5hqWe4rkfhHVGClw6lMMNDUSr6IkT3WVKCYv
cJtBjm8F/uwj9lQJORBDHJYXiERhf0fTpntku9QnSy2SeBiq9i95RNLFJd818Y7t
h+4EFshlZM09PYFjahc6aAVokiEyJ7DmN04dDHu9Ew4IqegT+7imr1dcCdA3tO1r
+Wc2QFdDfofTAXAKc12xLt33EDFwLscNrd7kCu4XyHqGudymAa1pz4dVpp1tAOHn
legZT7Vn3fzX/zKsejhI4X+CrdmuGQefQux1agB2tMjVZD9iDAnXJX5TjNBgX2KU
K/M1i1nKmO0fBcv0WgzRVu/2hKuNvKhL0XMQoXIE2JKYRoXQ3SwFLPunWDqvsIYA
Bzn33uor03GCdStYcY2fyNDb9S9vyq+cc4a0KLuWnvwqiaCtB5+s1026GIPNmFj5
MxCtrKRY4UBTAQjkJrF4/di0D7IWS8CFy+tQqrI5frIBDiMzkZ2zFdzDa00gRHe2
ERR3opMKYIcvn9UlMU4TjipQbdT4Fr+k1V24+cVHFH+RdQYIrRR9e0be6DKhoHOs
l5q63Vx2Wt19PsTOjKPd164fiEPDpwMfc1eJ9m3kIytAWUh1xHOm3wKtxcuAzH0q
VslQUu1UQD2HFfR241m93Tu8FU1CiuDHtbkGcT971A+G6VYvHUdIhjgvcetPEa0P
2B4UBuJd3yB7ScLCjWKoCFCJv/aJBVtYne5r4VDppclG98IdzBCpiKCjmkrqGNQW
qytZFr1cm1I8mayq0SO6Fzmaz83JHAR0jw54HkDMOWZYB8X7+kBJuybFzOKq5qlE
kzO+CnUx1z8LSM85ryivtkuZ3mBmvC8E4uhyP/aiooIGJwZD8/0+wY+lfPqiNZAg
7wp2tLxCY+O9Xssvdm7Caa49fZSikHGabHqjD23qF24sbq6N9oOmCafv9LxHfjh6
3yFYtq8axnV8Dw7uuaF+n+xBi9g7F3EMOJzeWWxRMe346OpzolYyyPks0ZVJ2Wab
v6d7LPHtojiOLE4C7F/Le4OGYbLNKmzjkFBlpgIb35bPDn3QpDFSFr8Kf+ZJy9+U
CdPNRnsKOGHk4Rt50JqYuapaBp0zMQe86jP50QTQchp6PjZtA92ImecZ8pFzdiX1
pAfb9beAKLzbDX/VDf9NWMgIKATvLNqtfuImX5YWT4hik6JTAHgIyDMOj7DK2ykn
WwUcmOl1WGe2pLCaja3BCPzHRJJ8urLz3ViFBODLnCWKXWGt9So8JcxSNXc29+sO
UUgtPW6OM1CQ8x2NPkyEQFQ20LG2v3YdDWpCUZ8LCouB4EbGnJ7xJYdEoVlyc1No
B2plo8at+/lFIXFDDjAQX6dd55D4peCAdxGBKwrAxhpkEhdjw1jlRzZqk813vY6h
yRkVY/n7dyYcszk5haUc8gnVHoE7KD70YFiCfd0+STukixBYuCg5AnrLyZAaOjwV
KvZ3CCEQC3aZhdJk+rwFfQABZsRxQTXMD0UeuroRBFq5Le9rbO/6xzxYMDGYl8Uo
vPuuy0MpXqS+xq2t7hhgq/IDnpxBIi4DnuM5CMbqDTOybw+YxlK86E/tue2tCQWn
acJsOxf8+lRMvcRNIKnsVoENm7sr/YVxkZrXNyxeIx6oDAG84GCiQH1X3Yx4Zwo2
JibqIWgR1i597mWinIKx8PW1LaeMFs7N0ZJubV9lOdQ0u9+58GKYEbxWhO9sdb71
n62I6XpWpR1CwxY9MwvrygMQjHf4hdf6HQtloBvMcLlQ9S63s9mB2n+au1DVjA66
GYZu7B2q8XWXB6zijhpeCcInA04hTxCqVoAi7adh9uv0SM29NwRmedNN6nO2kJ2i
PhbEHzmY3FbegZEn3RsFGfchOmDZ0WUf1dGVPdgcj+5pAWWSPQM5yUoEeX2MzPfl
rL7ONxHWMHsg4FqjkzsM6ffGStuR89RfueSxMB1b921usMMnDjRdA5giEqFd6QxB
Nfvthl8ylzrkK94HT9ZnYz81vI+Iv4sn2x0pxuffn2RcuIfsTTBkP4ocRW4WUn6W
3md7cOGsRJWKfGMSKV2z7pOPi3vSrXRobExjyi0co684ELymouB/a6HkHsjhCct4
gSmUNnQ7R5Z6tISspmN/88UBr9l8mn8JZ0P5skJ3QZXgtCdozh9xJpdB4pFqhKrn
AnXYXb9biNQTj59q9aI+hiPLVJfxASbQBVdM4SQHtA5OuMf2nAiAmE2aBtSVs5Fj
aNc3gwI9CQGAu/LmWpCBJrXheX5Xv4DQXdKNX6htsD0NFWLA1Uqc2VaBJ1aiiqfI
Xo4G5C5yd9+At0xaAmjLE/P08yc3FethW8jvxms56hfXH5SNNmw22RDmfHe2D3zF
xl+3iYM7R6r8t4OFE5paovIRlkZG1iJbSTHVkvF5EnoMsjnBQ5uO/YUHkUtqSlsu
GquOeyZn3XM3nYqkS+r5d8zsRxj31NGJwe01rL9ez4DUgncC2nfxUokGTeM1QOqJ
nZkG2s6XxPOoP77P//oovssUHPIvMphHqJH+R/Z7BRm1LFUZU69qs44cJRmHvVYK
6V3NQa4slTJcvDXBvyMwIon2XLSB6XdYlpnjxidTj1Fnf7cv2GkeYsr9lWeJBqsG
ePPaigR6AMPtb/mCvQx1IR8zrNe3rDh1UyvizdiV+m8Ny0QQ1DbsbwjqxF7St/hG
skO4F+2oLJczZCrR8B5oHIyxuw4wqu57BcKav20zYLAGIr5hh30+LylaK9434IT4
Zs87yE0nmoc+GiuV5J1PevjPZO41PfLojhF7cMlXj32FzbLbTT/Z1mLB9Gq6LxnJ
oUPgFOeowb/YG/yQO54z/jbLzkHQTUse9lZOTEASEJOv3vKutkA4WDkaROyBjwO7
UMcknqqyO9QhRAsmFPg/dD1592tae9NvaxXOM4nrxa9YWcZy40IUb68AeDaeL7FD
eBnanYgz+7rhz6FVzZcZdJGz+gPY/3gWymIWtaI1fa5kgtK71s4/7aqhJC9xxXyC
0MIxKvd3FFV5W8+OqDMvDt5H+TDKQ6uZuiXKf58a/l65IZ3kNnDEZ0SJUGLYXBUs
ytOdvQVtfrhBfuXzaEFe/xV95UXASOffHfmT041CYHp+H4KUyePEFPyGqqtQf6T9
2FQzMM5DsOZ6gf5y+8ax9n102VTWn20FeS/6JxwKDNqNA4K63AczvxKilJJeEmPe
ZoYiqk+YQx6JLNZLAja94ogl8VvXLBjcbwIELGacB8uTbpucIdCt0fH5gpc6V6wz
45XvCt9bYj/W6yDfvtu7iuTqg3upK7tTdUcM8oFl5vD4nqX5XoxfI45+M2UDCt8i
2tEVQHnHAk7QxrQ8qnuKE1sWfrl1HVXTIO7FHvtPv48PgXafbi9iSFG3Ko64RYls
/SWZuIm43P3ddKrL3OtuU7hH6cBE105lzxFP5jtb44MebqYGJV3GnLepEnzjNmmV
mixmdjUv6xaehIHvl+AD2n20YDb5KO4O9Ewq+AcL32u+wsagvXbSa1u6ghIYxZQa
snBhvMCQV+FUDur3UX2hFgfpm9ZFJAo03al3okVmyCd1p2kxHNvzNQj95XZOC/Pv
l7Mwb3x0EPfJX1jINdXeBCApVyMRZ4JcpZ79FZQ0+C+VXpvBQlNhrXC5jLon9Qnq
KGj56/PlHglgyTMTM6fe2ZSCA9f/A5SY0NQ02epwg0hB7SeGexL626eh4M02SFFH
B7anFBK1HEtted62j8ojMGvsZfnKRAUcUoLVS7wOS/iWaSsWApWyhAp/9hFoDJx6
/h9mLYj1U+EO7C+bPowQ+FCctRsx4U8R+v1hBCBQlu2XJNs/9Laq6G1PgohmEoqg
bd+cPKTsL0JuN7lCWNbJ06F1zuMtkYujjFSrhPH1Bmlnzl3eod9DTXdEfnx4E3bb
eDgKCfGp3U9cEyea/xdPPI0D6DoQQ8fpkji84+49RR6T+liV2EFoMGQ2Sz6mTpnL
IoUEh54u9QC0hz3Sz+0PPz1A+uogvIMlb7COfLQJYfX80twScqbPnmfUI9TbUI+x
XoQU0uMiqwVQQL4GlQiZn4p7TJuBrVo6pjdMIEQ8ZA644ROfW01hVfFZHVrO0hOO
UH+agKtrS4ja1rh5YEvKLwKkAMUHHIicGQ3i9UzShyDfkDLkEwP2ece7g0UeZdVN
uLDfQwRLnL2bsjh52R1AXKbgxRtPJ2o1znt24yZLDQNLoCpzp+6DJgQYPpQO676T
0+k11QG6nEI7t1xWzyyVVLWAWUpLTHnccmO08lIXO6ZjnEw5mnei0jtrg4RvnEZa
tqLXVaCF1Bl3Yvm5e1qazRzg26+N5ldV+CT1LIyT+arzhI/sEUhm1wBwP0UwdrHG
FJFIx5AcRAKmQT172mZgcOoHqeFY/zdMeNmI51zm2cEE1kU19vxLVNdRCjpfSyuN
d0ZgyMdDqlP0EpUCzaOge9n6aEq2kD0vWg5fJaoMex2xUNPa1bmYGn9Tk93GfG9c
BGGugQ9620DtveLsDMU7r9IRIFgzmTXh67coOMorYmjVRk4Z6RcAO3gHE6QCsT82
2Wu+XcUHfeDHbVKzL9lM8tfoPmyULVVxJ4oHK3u8Nd8PPewSrqdfpZKYKD87nBuv
yCUoRg3uIfIocWhb8lH9AcL7xdGW92ZVNv6EJCt7Bo/TT98SbmsOKIh2lMKAF2Lj
DP2oueJvlv0M9tlLsiy4SFJieyqx+wGUWM50yS+1GlxKCI8o6uKMdpXy66iN9hEn
9lDmv6SvBARj6X13hjWlz4TJ1WlhHH6PTjG2hYNeB12ap+AdV0NDh2HqjIIx4J1m
kFhYVb2MRhaURFQrFn1wgSKpt9bhzG0gQGwHzwHjNgokleaXoPUfzK0KJz+PMcg2
U8LzB4hNtiOSJe4kC+CD24nLSNOH/DusgBPjvHAUnh9lsqFWJWG9O/3T5qb++uZB
09Z2Ip5AErfowDZ3GKMa/KxPZYDJlh0TrlJOcGwvql8oL4vYLkznKC/y7yYju1NH
weHpsbQM2ThOfG7LIVEH6odbDxvk1JOiofs3e1KZE6sAmkx8aJ2T/fzaHm/MrFSz
1QptNchQhf4ZIKbh7GlV+thN2V0rhYkljY1UXw6b3TxCvLiusC6ifMbzzby+OUYA
L4JO7Ck8dAIdOi1UZqhZ0HgjHQDVXGxgBUjEEF/sqcckUSnQSgBjDh0ebg1OZYBj
2eUZSyCAuo0ixrQXu/XwrjmNqqqR4DUKuae2LVnP0fXg3BZd8ULYPnvK5jDGAFi4
r4j8djle1DyAL9HjypaE/bxZ3vkOIxwkRONW9Gm3Oh+y4ijdItfhpQpmKPYtshLf
bGej0gCvO/A349gZKG2lhNt6KGXkupiuO9wdf4VCGMqJfA2szc7L/HvaeAGqR/sI
oPKjdrKo0sQWvlkbrri8y1bDvQNfCEjrJMs/N7rHDk8V4i31WaMCY43ZQ1yPKQx/
+k/EM9sIj+L/UCydev4IQn3voqYkbXkS3H9JzdKMWw7l9wqTCb20SwIGU62PzQcO
tsl3hS689/JsLtfqHBN0coUVNWZoxf2tW3Rt6I1/pYzfohnxjoKBg0TrcW8UNM/9
ppKqFnUlHbjfoZ/Lw5eHT2zyV3b0z8sUgXA3S39Abz/aYnUdKs+3bP/lYBBEqpYJ
k+Bj8/3OuahIbFgG10dFr0ZMRiMT6DaA1YXzmmRL4VdmJoDXA/OZf/eJ8SVMFyyS
3DY7OOuaIorNatEBTdLMn+acMlMwM66Rdp6Si/hWOW6syENZWEYyXZz6aJq2WCeS
zBNuRfHX63e1s3sEewQx01TUnI8/zGJcnOp8csMdwEaXfgpKy1koWpH/1dlNA4jV
JqsPUruoQ3VH6dvRypRSYEZ6kUWefp7Mbxoyg99IrjeLP/gNpx5/d+pdvxYl1KZz
cwBk+1RfeDzt/eUVNbIX3YokFxp4Fg+40je3KXKNX6naZEwLSwzgQS9FjUThDUlm
hJtOXA5Qk9M2bZ6GAwEC0+EJOAdkz0avzJliyGnKAIjTpEyibhkarh+uJxxkjtM5
Fk7eUCho7yrhJMmjdSbDxN22DaI/h/C/wApEw2/ttIoxTwYZR61jnwSiW0W0VIeD
Tj6GthovHQetKtH7ZEyW3JQz0XBDW4iaQxcTRZ0g46m/cj6/uH/MlRcWb48b5Np5
J9BAopX/TkCYT855zUCKoLKhtH/7ePWOevvj81iJpy22gPKUufD3twNSnPfjwfZU
KEluPYmMk4jv/GL75id7fVyPUOsd/+ZZT2zUm/+O4tU8HnBguUomdhiuTfxG7cXA
ukuvEG/xRKIZNZTNC6r3QkXvX1lOvle/GA+Cy34d7Eu/wegrS5jmPh0jIx0p5qiM
zP/Ym/aCFkR27V+Ksh3InPc1JFK6rEgBExn9kxvSHs3rGcqyPiosGCfqx7wI66Fa
EpAbAr9P/UFxmtBm1Tka3MH3P9xC6G+JUTgNUpyNHj+pOK7Muh6ZkQHg0Ohtbo1v
ZzdoHPDhuyRg97tMGxKOrNnOhrj+yFLbFv1hdWZw7iBbGvjleEHlpBKvB3nSwWNH
0LFHsqX1xK5IZ5kToSgMMGClKASf3YcKywQWJzGX/IkDAonQ1IhwxqSZYntqssC8
UUBx1tX9Nh0CLTFdM3ctk5a4v14hu0FupfLRfSQNVuTJorJW0coAD1vHE72Zhc3e
GQYSMpLWrQY62Sv6na38YKNqQC2xgKDE5imuJ/0Ds9i8mFN5wPbWIkGkk6sAAtll
31bf20ATFE+mCfr0Q1VxCBOboAd0vuHKTBywhSGmYzBscHoIwNmbqixRzbSkNFfg
xkWryX2JTsys0YbaLC3oXRYINu8vS+j6HZQ4PEF8osMcYNnhOFWyMtY8eeCkLuVU
hOQ5o0c9gEMmKy4ickMBlgT1mEQuVCDSvitZ5xJ1K/9qJ7KNYhBvhi/1VZQRFa4c
ai/uXOT18TD80PuBfm8QHaHUOXRXEGtbDWaKfm6LGX8rYsBZRomhT5+ecvyxt7E6
D/VyY9sHA+WEmzOsGcb+vU3caDoTaOPK8i2YKzKM9NBFslbWoR9nfQainqh2w0Ha
sduUAK1A046FJmKdWThgJCMKzut/Vs7uGwC4Ok2OphWPGDOgHbofH7wsZMTwYH5P
2hMSZrbPlM/9YlYA6R6psJ2LhMCi+7pDnD7XT/frxTV9fUwkmaZTRFfRFKJY1bzq
27VKqM9d419XVAVG/Hb20zzLaybrvjcwx/ajd3vruxqaxDo+YGtPcHiGkV8ebOcf
+iXGudKPiqV+4OHAkCya4cE6h6oegqTGHcGEkoPJUN4nN9feA7+FgUvR/auwW3SP
NU9ybrb8edqBJ1TzK4zO1WgOQNC4mX1PlyN0eIMidcZ8al6Z0A7LZtgn1P8W7rL+
ZQiwMnT8BxwUc6ZsBzVuUJIfLSIsaceUIrA28PuqVXgYF8900WkvnKCbnMZassN9
seJDdOVYW9ty2TLyr4ygnHh+1wi1Z7oAw0jDt8yacDpYXFsuMwdkOLhN2O0WA6Z4
3jMqDjZV4YjoECYMAeYhcT9hgw/LCCnotB97HYjvKp7UzSglSirkByxTzAtdOI3p
gzIcrsql8YHQ0emTFnENUzE/lEVJJaXDZ2LCe2xUbsKDK8Gm8krkNEa7qCpSjU6m
BdXJqsjANqng/D0URRb4HMeAaFIK7EIGAjUzp6tUh0P0sAt8eY4kwYJWKOzISpM/
LzsPefMkEZ1hJ0QcLBf96kGf5bTY9NxTUJGdM+wGfn6UQgY6SdjzRAR8yPu2iWFI
WPh9DDngmuB0oCEZJNULirnPgHoRnFFnbYJ21IaZR/uCYskrc4+C3dlQ9DL2zwNK
vn70fGrLtnP4vLQOYNRuTR824wnfX3iZHP6IojxtZoQb5zTzRWxtMIhG0+EBI5U2
TtKpVSEi3V0JOO30uShjlCEGWAOv2cZeHI1BmFXtCUHVTK5gl7XSMZbED6/RxWFT
+YFS91FejWXzWgpvPO47hHDADiPRr3C/gK0sPttzBvN0bBrZe77E+Td6U+MSGuRk
3ccX4SiGIeAnReawe9zcsUwow0726VLjb/Qz3IeHcmGmLCbc2C0UB/z5TWz63+l3
MZCIEKdRhUQepD8di9oD5C0UkKOfxXW/7tkWRbCUw4GpGjMFvszgVbUUhMSlprS4
omFJdmZPyr8SvFq4U9LXerZDEdLhD4IIt6u16IpaykRpOz9cA+bBmAouG89e3w9I
y7NOpSjCUjyjqH8y32DCkWlVsf4K+ybhWJ2NSqWw/ibw9OW3uogUXaz4AjyY7z3R
Qu+GP0aY1+p5xV/4Pa26+sxDQ5ZGEMw5WEC54vPfHjk9ak7Xm+H8TZ8ODO/ji/8I
Nj6WH38LbljFAs8JX4aBrOAebA4pYbM9PkXWWhKixDKy71yVvEds7aaPWHxRy0Mr
/XAVlZkOy/XbNJy4XgIARv95lzhGl3qKkciX/m/PsnB4YFQb7PY98PVT7A+GE5kZ
w8GDx+5cHg0BByIjiJUVsUUn0ytsWME4Fvf+oSLjUiNo9gboD4K+4sDbIEWpam+1
TUzrsYLKlW05qvbOUutxPXnXzDkRbc0j0MzC0RBOsEakfI5kMKOkosgX9/1CBbWm
KaAl68QwkjTnO2DFT2bl86tSdh5SUoRUlmHqbyuUYIfxUhqLbYtjObxM5fK00kRf
Dxyclb/jtWpTuQmfHYjmV9ep0nmhiIhlbfi0yaW/gEyQ+k3zeiktNurQ5FQ4GpGG
KK5TZHm8obV10mG9C96+ANd39Q9OvRnk0G3WCp44kLakjMpDeelRh7RBDp0xqDkK
IcnBaNm/33ciGzrp4CtTOdixdGZDE5sJKCw3UVLCKQtvmWIcTthbmjIjIWlUod3u
g65ECDIOhRzc9v5+wE2ksYjNPVVrKccfrsL+t7M4zvSy5YW0rIVBEY5HsM/KKYSg
g4Q2cs2Lj2tY9Cf+3jsR5j+btvTXaL0/fcRP1/BccFPX1BsbDVX21edN23OiAVw7
WDSKqxVXR5VK0yfBVO0KKQ+pRmeZtUgqprGMk762MSDhy1/LKP6mV4FEC0uOJC2T
hywtYEsirUVx4L3YcEKKQtA1Q35fwuLapeiwSMPzpt16dqMLPRDN1Yq3fGcK3z54
rkUR47j+LbI6oASb52RAF1FqxdcGDnkluF04Uh6verwH4SrsAXSx+9v7TbBlkNoL
prLlgtmUnTFAWfC8Rex3206AbinrFKAi3bBxG6YcJkG5UOm8LoTma2s5nmETTDrC
3F2GF0HNPayAZkTFB1G/dtis+wJ+kiNGwenZSX+q3eMPIOdMLjsqmsHpuksKZtij
UxIPu1/AFcOcxKYt4h317ZJfUD8Iyql3ZqbICjw52SPKp2CWm1ysSO6PGNvUkRis
FDr46bEbOahSa3n1/wg1A051aS3dr+Vr3vWu22gV60igyF0AWqpMgifp0WmPNQIg
GQtMYPEzpvWSCUpNgspElYmEd93T/zbNfhBh/XFntGKcIV+q0EzsTGpyvlw77EG7
5BFvs1PSILw8IP8VgMEnycgAw5/rg7Lpz2Qz0r7N4QajKCQiLlzYNviyeHKiQn8d
8dcW2VBTsfCKXKPdaDYygKMSdx2M/nfD2vBkuglETzGWbkvs1SqLFBRlXr3PiT6H
jGilDm+8801iJbT/TletfeRZWu/+Ccw+2Zotn8iTE+jA+DPc0L7ExpU0yNyyEoof
6tJ77JldFd1vQkao8/7HrKEuFktgPHnW2MpiPxV0U2OxBj6aDSkHxFruc7zwW12c
To9zNmwIOQfoBmMmr7p4j9ODp0Fvc/bppnum1Q2AlqQxIHeRFPbaoay8MClH4WOX
KDvkPmhaPHwgynDGuqzmI82SpcxZH2ZWUwsgOnYYrKyRMQ0o/aPeF06xnHdCWE35
3WS6TZw0q2C0FUkarraCVUOSZgAoveuBq0JXALEwnxkTCmIVHap3N3x4aOlNyn2Y
E7v0fckxPTgjX4yjD9TewecP7EmyJJwDkQ63hkrdHIwdgw8gswvbZH90BrCF150x
6SxVPLKRV/gKCuTrtTb4Gmnd2+iOPhLWkSJTYe0qnVj3w7PdXRxsXE2pb3oWB8Rz
kcHgDQgmRY/+34bS5m5QQ5zpaW6ge3akBsXrzPEWXXEtufk0U2AJTDF2QSYrQAU5
wjEM2s41ml3bseN99mmtae5/UBkL4Ty1WwplyNUh81EOcaJ/6vP0wzBfYSGPWp6R
E8hEfVqg8gkAaCBm1wTVfuIrZ8NW+M2cMJruNKE3jmd6N3JXr8j40+cCU1avbVg+
FMWt+ATUWxn3fDIU2yJitHUYHJlG52Wmi5APAnyKPomiZMiR1AoaijTdB6LoLZZk
PyKFxOib+HyowmObFNJS+i2CuUKWMm17AD4R+db7ePt19iC4qiFhtpxz9ydj/dVU
OCJkOvQPHyCVZ3eeH3kKjk9Osyp8poiXcqFb/xdu4hC21oHWiqw2VI7jlB1BUPGl
Je12ShFGh/hAfXVGI/Enss6zvsAlq3+4ZXMC9+eiRCST+qfKC1UUWxIzhjwPXHwV
TbNDTsf3UuIFlcDfitCkCr1eo0chh+w+RQGqENzj5FXhAnbpXJDIJbiYhoMTlHt3
HPXXqAvnCDuHu+dYWZHsObcViuvAuB9P8yMhK5BexqMJrhqxQzMq3Eg2nZGrmCoo
QHCGGTGCKa9os2fxBYdYeVdjIhQk3KXyhS4Ck9IXkA1K7vaCC6uoR1vBmztohodJ
XYszHRNywJjl+AFdD/fc0SQj79kNpklTOnGz1ethPJVQd1M+6g8IyoVrL2FdL4QL
kSvMJidDLri0mkmWGp+/7kNlGYupkZfq8Rtl6G2O02OP5TpCxxu4Q5Xpjs/5ohCQ
I9iRcfGzfNnIzC3r3jPrI3do3d2bebzNy8hFHEiZi1PFfNutjnPdDxTgqCd6sHcR
+fOekCol702scBy5Mg7DKO+I1dyeBmGyw9x+0x6Zr/s5sfqyyUofvbpxKqAn8853
GmKth50rTfl3Kq85Z7ZGxYZsnxVbPJLY0HdWEQ6LbIf9xX0xZbpOR3Z1jGcPirc4
PxQ0Ngkan+dcCmtl80ixekPXqrTbaJ3L5ZSQ/yxruRBqdN5d7ZNczXoOXyMbKs95
tXDzIjbvNP18zzYSX6FYHWO0XRMyYwOK6Ria0beilx9G6JEKxfephz8d+FPQAHvP
8XgaZWPCwp53qe5Qr/uTs4R5f3VSQuY40ngX9f16tNHdQX1L56kjAYts7K9xT0oh
5W37tKiob4939nL52hI+mGiX+2qOZeeaKFWjrXPOwXBrMAEayy1w51fbiG49onkz
/0jJ7uBKJAq5e/EPBslViaFhD364gmwlSqoUmEhnEXldpdlKVQdDkeqcdCDxEiri
jsVV2IneRTHSzjhkcqMZZRA5TifQJlFc0hQbF3TM7kB0zAD6NN6pO78w0vaenjV7
kcRMYL46/u20U89r5gO7GG+vzJCOowxLva2ImWNTKwLdtU+JIndH+qFupCK2xDDN
6nuF73jFaE/dFkRyslilHP/D6ybvePJ4X9FFmQ6P2nsGimtHNYfdmt2wPPgws53P
Kdgson1Uw910onmuqZaUCfvRWKF6T/2vPgLYGHKdi1r1KHCiKcCT8Kn5WYDXyfN7
9YBxglB/Dvo+JC1esSr5c37w9JYuGQBx05emRwX1ejkkpSQ45W9CHNjFUhKA7I9n
ZxbQ0lENALLvW44Hg/H3WFUq7c5QxXSbp3TDg9KTFR53wgSSWmgJYOIf1+XecDHh
PEg539tmXZFjX+QFU4LO/JTYoVh5tEcZxc10p+Y2ZSsCv/+K2aGHDz2SS9w6pSef
LEOPlXEppWEiYwjkz0LbhuRaqn5/zqX9IY/JXChRA3myNeE7QlJUufaBEXHx7uOf
AbawDlreV64MuBQbiSLEoveLpHvc2rBeWZ6C7qRPZZhsAj7F+ykctQpCxeyvXhvx
FKVyaimQIDnc2l+WAohhP8l9wqcp2/uYVpx+rbJ03x4K8IRWzn+XiltY05p9gxfo
ww/Z0qYu8H/yOVAHNkhY5k/EktBjnMaVTR9p3am3AJPlIXyV6n2LtGUP6REd92Z2
7gXRasWrMNhMlwadxlsdXPKe6eWCz5QaooyH8AHQR8hgx7TeCgd9JePFMHUjYaMb
/nfkBv6BfbmkAFyPynxxc+jrDF/g66sYZBpkda8DU3N5Y++mxfv/Ce95TRLUQIMw
J7QkOcYF1iR5MKELaFFECqBzAK27bnqG3G9suEc8xZOL0/z/EnrEgSahO6xXhXvD
oYCrZ+fSTl1zC10waoWzNQyfTYhc6xRVHOdHwi7et+qpqhLv24tTa8ScdrPvxtbN
offcUZzYOnerXMAlCoiVNjL+0O3Isg5S67LhNWIKkQVd0PwoPWz0xkC76ye/2eo5
oR8jwrOid7TwnDo2WjfHmFwP8Vdd56xQ1ylorHWqYkEZYhYippQN9lveLAhIbK4/
LKa3Y83P2chFETY05ON8RdWnqA/r+qFcsdXl3ObV5q2K1FqvwcE8kAwmNiIcLa3W
fAm2Mw8u0uQ8HAFcSNaEpsy5N2wuJM3wwkJ8AN5VoHG3H7Q8dtD2RaM6rGUaMHZq
VMzLGJx6dZj8uOdpN2kgQxmnL3mtNZRNKEvOSDtzD6ndhY03MVGcJSVwbentWTZQ
JozD379y/QNRAzxHbDfyTu5aX/yqufB9JN9HYHwjBUakwkxXs/0OD6WlyuspPoHz
EwbTCNIypC4ZIkWUoVKOcB4GKTOYfA0Agovu6PnFcj34M357uvCclirzLjCF8eXi
j96/Jp63NlYkFDoiug5nhlaR9GuEjXR0BbdLX2Mz9M5r1Q8WEKydu+nrE0w+/GYG
/sv/2UGbDB+h5XnbDLKRO3WG6q9X6ITkPpLCaUNsssXf8X6x0scK+Yz82vbiIe3d
s148L24H5wFEMFbgfOWROep0Vr+rLzIfkcXSRpeOqkanHl2rRQWRrgImkSDzgmej
EfcrC+/zG2eHAgFbYcZVnYSijKcLQn6QBscV+Av4LCrgm+6gPQwFoUsDw+sXCuYB
33FSmeOLTRtbtOKlLXaRtIJOL4KH/MR4jc42DEHhdC9hkdBzDAT2sq2T9o6lnxie
Kj+PDpI4dwud9hp3aICZlcxubstWwOdWcC03FnWdFPUkeuuFUuaVo5AEiDetMtfL
PaSo7Ye9QaTMSFCCLyr9HVS0x9SO3rdK+JGhax4g7EEwo5l8+BgdT2J3xGsmxWV0
xS+NU3HNqoinLdy4jYMHSUz/381BPUZ580IdWntukbh+39FUscx25NdGKvdgS8HP
iIJoIpBjm4SThdU0xiUVWRVEAI5fxUiv9oPQYzDzrnWhjO0LWMaea2u6dbkqKYgC
gp8DM5gqjVJuXnKo3UY1wK8nCaoK95ShY6R2rG11I9vo87NFEqdbcMpzGCLH7TTc
IDiexOq8ykYBYQM4Bk6G0m/u3rIC/dN0uvvQvyaKkDn/aeaEweFToRNyJmEjtMAo
35NKv7+CrS2Lkxb3DYt7vjrczv8PeSfvAL6MBn1PSDQK/AaPl4H08gGqk/53chuE
u4C2bXc7BPw2HWEaKcu/chiWGW0VNQ1QY5YIe9IlSGnawEAAX1Sez/rDgFG3x7gq
kWuA95b/fjXPtfpotkyNB7l5AZPzPkhycPazuQfD4a7Wbt7qx6Auinlex8gQ21kH
cVfO9ovTC1ykNbeYM798iePz2n20/0zFDcx7cIWRZ7R9pmNRyLatY2PkFQK1Iws3
Jva+cCEx/bhwM0QDCvZK0EQGKgtoySaAx0jqo5WP7wCbnrJtxPSLbQqtpef3tzOQ
BOus933NsuRs5yd2Povuc7Pr+yVPjIqpOSPzhWcVwqU/WkVFtteTlMZgYSUo2pMY
8r0Va3eEsBvchAm7bSToyCU6wGuR9v6KGBcRa8XnMR4RwvncatvAsUwXxIPDLZlt
TcTY3xTFJQp4oWp/7ok1kM0Im8CFvGq1Rzqlk9HqihX1xr3qAQUsSlVoE6mwo75/
Xx/geAPyV24UuyWuxDTffVxmHEMm8e1t/w3qD/UGgRbm5EDqxECTKmnq5eRtfCsR
NUJ5Tu+b7AoDUA7YwhKBWoG7KdiMyOTgzj61FdMD6Mje0t1BW1RGJuUGgEnS5MRW
ty/QLLb4ZufVflew6/6bAoAJ++cNiudC2ZbzDkEgPd/r6cQEkuA/M/xXdInidT/C
Up490SSnJqDzuLwJ6Qrg+koMs1x/L6z51JrkL31asOqobKh/xx3JMgIJL5DW39Af
cXwBOM7o9mIApDaIId2lYyXj1JC5QeHJPcHuEAzENDbXc82Vy6u5TvLS/9MCcBRn
y3abNK0LShjVUtxJyzbSxGKETv0/4BuZxRfUasPPQqY3KOjakBmfH/39pdHKEUuj
GJIJQ8orKZX78gjoc1ajmXIh6qppCqPCrvUTt0ggfUhxAjqcxVW+wh/J8MUslhXg
78yLaDbRNkbhmebN8IfY2lGiTICNAga+nsVlG5iKg25nVTZTGwMnORgvqwxdVupw
YzBiRbKH7Ta5UHTg4+EizyR7Mju4QD4hFIaowtp+OI+TfzoNpEBUSNG+LMDFqN1q
tlpdY4YxC2Sy/nTeW/VunlJIGCii5goPQ4AYOWOpeo2JJLz/SErxJmKLHy7T/Byr
AdcT9UieygdQccq3urAeqOCSPF6u+UcDXjv5eIg5PfPX3VT2Wzfx4462g3+Li7m9
KhQmLB3XpL5oYPxqpbwgEXypvM5q0rD56bwvuFI28QxNpus2UaNx9WuLWjGB5VdX
xDZwIwLE/Z/tH9V7qe3UjHd1JjuzSG2oWOQZfNIfE02ME+kavL1aVCJYLoFlHG8b
tm010A9m+3nFiP5fCzCYhjzME1L4OlSBnSJvDGb3udtOQxVPxDSI+o6lYIknuZnn
XzlihF6Go9qcr7eTFVBHTJDtokO5hnLyG8qTKIPRvx2B0UZizc8UoM0NXU9e+aQ5
iNeUiKa6Hf7ch8bBS0mIlZPjeTf1GQngW8XFV082OKJqOUelMD1vmo4TsfJuljJI
2lKDJ1Jaeg5EHPnIO3MBlxrNQ/4Su1wwAB3PPSfaTmS0ZpbS9arv4W5KwjLM0OB4
7bN6epqaeLMJhA6tuBifwpV86mq/RKFnI7yO4Ijvz/hRaT2t58+AtkeTRBEHTgwM
Z2Iv//Lty8XJre8NJv+diT0mG8CzxZyQma9OVDYeHu3LzCVGYvaanYDGGGfRudFn
JHBjH4WNy2ruabS5/h6sOlWsCHhvr20ull/l0aL8i198PaluTrw2Au70VuGSKYQa
2XpL7sOhje47ma36zl3nw1wd9ycgbksoaxe6qCZ8Atz2TgrneEMJ7iVD8MEjAzc9
U6X7cpHm4Rp3WSWHi5b2CxsWocc+vY9GQFMBdXQxrUNhc8SdlGbKTA477H3UwtSA
GYqY7/tRYzV0+SLcLZFtkleGyHmreNsmrvYaA3oy6vfMQT5BnKtvgPrVt6d3qVp0
xk7VO/jffc1x4PQgb2Fdrc6eggthZO2ZNLdRMkCxFVwn9os721sIe3yu9iHariU1
ehuoZTy4HkPSA2POilHlpIMYFmXW4h1/dUYUrHT59xxdd5rjL763uNteRgkKNck6
l9GRoxfECtjV7ken3mzFDECb+fiQET8+mnklheoXZgOBmeWe7h4cCFdvGude+ybi
gHgrDChAnlAv3tplvM8+QiMNWwOLRkQk5VX6VJA3T2JE8reRAkm1RbxfEDXOpSPw
pKfzRnPWDRb4WyHHWObhM+zXLn1ADRbG/mvCVBhU/WszJ2PwLXaPcaJV/dDx4qye
C43m2QFWkLPVDtuwaEjhpYHy1odX+qu2jMgfS+A6NDVLWkeMl3Szi+J0jD45iMO9
kCau9w9BsvFoj8hbaF6Q7c+sjvTYCWNlia6J97n9yzVQqf4Wm8cabRgIQwSrNE57
zXirFWAWAKJuR+NEiTdkmGRGInWPoGO3zHkKmV1K8w09PPFpjVWyovZJQxp+Y3Zl
PzyKZrP7VIAWfOnnEuthXWH/uvhRe8/GA5eldW+n7hU0hjk8eK/tFlcv9hKqUY9F
JwxdyqphHruN1JxzcUbTNy9zV+asF9dU9oErKbaYXcecn5b87fj2/XQg069YJnHs
bgCSuUnV8Z8Q9rCsG/QJI8AZyX5B4MVxR7PK+ihaaw/Z6Cl/36to28WWn7lRFPZP
pIuMQHqUdu4NLBjeEF1SYPTDPn14fsY1n4jSoSS59Mcm5Z8+gJsMDKHQjktwGy3D
oGSeUtiEAy69iDmA+WmZTcc/S/1KPSoFeHbblGyb9WqB1a9hpxMZPCj5T7tyH9k2
ibdrHJrG98RJtqYENKjmga1sHQoszzQ+e8uOX6OzoIdSiQaVn+RiMSsuRdbnObuY
+7+HIuVZd5tywk7+jG6TFfuoqjtqCF0amj+c2IkpchSZIGO/Cu7E4pklDXotVbAR
j4jjf7h5i+j8d85Qo5rlCnwhIh3H+L3h02Fc04qjeJoOi2LA4NpW+5P/cT+oCbgn
6omYkd+U2fWlp9B+EAwa0IGrzgKHKXnNZcvCi+kFW8/jC2Y3y8yxw9lsF7tfWN6U
IBAfO71UKqQZJ42/lF1+fI2XQmW7DJZIIVuE1A0uMBcXPr5upF97RO3TZupglpKt
NWsvvgVkUkJ3kdUPF2ApP4XtkvYOONtY7TBLamA8lkmIdr+qt47ry2bvhIn1SAKT
DgFySBftG7mX6w1sQMP2c+vrrskJbUXO26nWhMFruQwd1nveMjDFcxCeU0x/XITZ
ZmaTCiUDhCRgKmjOg6EMtRCC/2pTIGznevZxseW6K+2I57CzrBnWPrdmy3D7/Xty
SFb/SUWdVX/8WzJehsowAy3C+l4HUXTDsdwMQaJ98Kl/4BdiKgRgWZC73ZMGXz3I
YH7MkTfha10TheaAg2eLueRx7lE+oDY5TaX/BqINd2/inop2lj/Ki4ygXWZ73Si3
kTGFI04j+INhf8u0JYgQITjw+Vc8YhTwDVemu+gqQ+c2m4VodqhEymJgzUsXg5H3
N01azBeW1hrQqdL1VL2ydA5r1HyeqABrYFc0a+9fu8/OAfD7FSVMzaXGSABf8R1Y
9bn6IPkSACxpn0qV06Z0d4JmYMXdozC1ImIeDSgX9ZYNxmvQeMnGSDl/OqipXJoU
jpkwn6VDNtRCSbtHE4VKMyhiXeNTbD0aVw+la6H6bdnkKV83m6Gv1l3QsctXFlkL
LATMs85uFqFfYatjATCxPIblQQwSlOP+BqyyrBfH2ANxWgUSkdw0bPddVHBIvTA3
tIZFmUV4g1O0S80KHa6npkfMzOLxs+YPzgMJxur6F7FKlmPZhjxsuuHsQ5PauPer
NZJk99kRa8JQzrPkkalrztBk0YoKqwiG/EAK8UY5UPwDuB6a+3TQGA94HiBU7RTY
MGJao8UDNe+GSJCTJ7e/7zYHbH/8MRF5uVxSEuvl/n8xUAdve09Q5yy5OhZGO71l
f3DUdIvyod5VUwe/hh+Zs5e8MU2eD//aRel9sJYqfkk9MM1J7wMC2HJcebDNuQba
pMhehU1sB3G3fT1N+kutKK9qR0594cQOGDcOLx9ic+UhTLHzJAN90sRCmWWejV1R
PkBNzcNp373GVwK8vpix6HkSY7gxZTwtw2UaQri7FPIhLjg8YJL5ludaJQ3AZtVe
q19F4C2i1EHEEZi74uBkwTMLMdbSUN4RIPNE/T7/ZlslC9AMVdTMF4pLOykMrcgS
pAsSphFC5oBcR2CBLTE6cvpc6e971Lv/wcYwMX8G0pJY8AelcbFCIC/hhfbXjklT
IXUSQbwGNr0TUuOR9NlEz4Hq/VYwYiaYL9EfUHGh9YBKTXUWepPnKg6zeEpTerw0
zli+StBppcs6HnS0BMdmc/x7rlDmR0S//KtRYOeg5EyfEagVw8oUGRQS9k92+Eyz
LPX3rHgjFPi5qVaNPLE0+bZYfRqIeH3b5xQiegWWhMBK+Kjlunm5lTT4FiKkRuia
Gs1O95yKa5C4PTgEhu7e5gjhQQm0mqIJpBHgbNCW/uivMhGSyb5Aihoc1I3Ya2Ld
u6WPJl2KHiC/OoS5bhMSFDLDrm/XOreT0/DZDRCqN/zfNyzf7oe/XM9ME1Dzvynl
eYdhXxcqO2Fqhg79Ax4Mq6erS/OkHu1m7/h2CuPCTzu7Zk7ZeoW5IKmtS3KhNl1J
m0rvcKfut5nL2HQRtpTTVorOgIXPOqH6rL44Jx6+d4Ucb0GYQv2Q9Oi5P1CjevFp
k4P2pefYqo54TUfK3P3A2+cuyc1HYbYpWXmDnIhihci3LpnUdy6AahomCwccdcRP
4lPilNof06jUz/0eLlyKTsTFPGmTi+ujxLw+t8bOuaXglak1s6NhrmtxJ0kJUjRC
pHEWBjYYbhncBJ5m4SyvMO8DAjCh4uMf45VU39Nq4vaJluwNDrN17Pw1WctwwoK2
UwoDuNcszcaRdkhWnAkIKVWUM1E0iY4UQ0telrJNJJP78RmXu5IEFKljlSo3ZdVf
LZWVw9+tQrk1Ultnd0emn0qJtq5kadZKKU5BqLMisLgtsvNuYm4Xxg9p2UgLoZUk
nrdw0rLGcnwPr0Zc0HtnLxe5zTN7aX5CeceD/9lFWq0rIqsybXwI7ogKl35IAiKv
RsHRFTFJIZYm+gthd7heBfCUHfR4NmcBnPEKwACgHjNEVK96qd90um0VfR4gwTuz
KI1TmSa2oIcKXTXR425zQsKe2X44X78eCuMOeBSWlAbhIUUcFqT326jpDGfbEvgc
dqO0StSsk+ElER8Yvg6qgBi3YItSOBUG4qEh0ngimIn0kKLSPiLxYkS7Ndljg71w
NSLTs68bwodWLFfUVaFXRebawxHOHnbm5B9J2QMnfofGi2NL5mQ0LZttOsKHD2cX
aL9vLE3NkPo8Fca1xZm3n6vMcd8H+KN2pRzzxP4n6YQpUQCfXs36Jcr7TRVY14/5
Tmh9vyeRr0Wt4cULxPjrUSyn5trCKApI8M41T0Yh9LkRI9mCsfgk00Kibw9vNdvR
MxiPLgydNjhELkvgiNs8hwB3MIzMqM2aHccDPAAHvdPm821iMTTuCRLJs0pFWN/y
XTU2494K95pk9OVwGAIynK4WYBEK3gUzdSVpi75bXx+E+eZvGknxyW82t4M2xfuf
Ae3WrUa9b9FsYqDLWERiJBnrSSjDfJ7aa8kc7CRnWMI743rrAFr7wsL+/FF6wYE9
Q+MUf1/RPWf2oWRaacslAHkTGZBjwWBX/wA6h0qKH2kgVBAL4MZ0LzRwL1cA1O7v
e0Dx5TVbw2WkLus6FMDaMRTiXEIj1tqaCDkgFtnnowQxeRIiy/Q/JllABFvaXbvN
hOCK6bEKxadNrX+pNybhTwwPFFpiqQYBjL4LiELNPqhLdX52wlLaVgG/MMlWu0xi
eoUKUFn2z86lQ4HottVpX+tli4QSOmkCOgmqB74B0kjBSqbVG0zV0RnRSUAB7kId
ShjYw35UQ2SIMe2+9XJd0HiXGwL9hWBxng3tvvOViivAlKI6LKFgY1pSf2s/spCy
aSCX3wkIVgS8fK2E7Ac7DkMyzIRC5q/U8+Gs8wX9csW9X6wBDlZgfhnRjmIdPR//
uOEWq8d60gp93h6qe7UvHy/7AnKsGQl/fOsbr+dEuyqWgRHQwJWfk65Ul9465pAw
lv0OnIz7Es9CsIEY1S6qEWqnjszEFqCkV1MpDi1Ev87h35N/VpK+5FZIelRNfwWI
pnt5j/jIr9nOt1qAYaDpj15PSdjPrnZLOB8ZMzw6QFGvpySrQRpqrzQZh0QGhBGj
jumNQgPT5htUPhu8LUQ3VtSjIJdDmbDaeiS+2XWU4rzAzsJOl/6RAExMWgBEv3Ve
i9yQKE90/QwfnMx7qd4LTwFgosYXMaB4kii9LqZGGcuYCKBKFu5BARwe0pobNfiP
2TVLa66J2juL1EYCCP3ZBWAdYSfz3jc1rsdTV32nIte4xI+Cvf9iMuduQ1EM4i0x
FC+7Y1ZMDjWRzLIOvsmD3cCMIuSLWoGjUlX1/Db9rbVS2RVt3h9mtfGlKRe4saSM
+74Qu6Lv3WUM3pAyYqzt/AJLazlpu5aqBabBrfeLagNyffsT02cAsCbWEtu8YMVh
alpG5rNE4jJUJByrTezbEJXzEmOj/88a2zc88VUFOTPpb+lH+SQdWBpnHdk7aV+S
Bbpby3PgHgbbQDh5b7z7niq39Ft4mDb0If7taKoN3ihGm72K1ZUix5jFTxItqPWR
lTZ9t20dlhFrSIl8pK9LPzFB3SUyDXtY+1oc3n0vck4NPtsoRKlCdDpq1E7SQU//
xs7W0ty87nGFhP6ZQCynu/3DvJopp2/3fQICED1evSdmLFE7O19JShaPHZhMUWUq
Wo8xxPaxPzCVq7rrn4fczFiogMl7PLnA35XH8C3Hd5sUZSljCNEwBo97C7In+fnx
IpOk+QtAasMKf/r9zL7ylV/vBfTb+fSW8kKQsCCGBcxZFz6Xe3u2Wvoj6ZNOxXU/
ok7BW2M6tvPMOmktjNCuIVwipqiexg61Nx05HtJdRHCh8vEfsDwgHyL8rA9tReCO
bsEjlZ2rNSEKNY2h37/GQ4/nh5Qq7e2ZHh9syo5lA8XfnP59Nx8102baC1MZq6bA
kCyHBILYq2Q6HGGSfT9R3fDoy/WFRhelK7+76y7ZF+We4iIOJMZ8Z+DUJOK8YXgO
JjzXic2R0CMRCRP8myZoHfgzoytbmOaQKeqmFAyKYw5wQCe9pVpxchIgBwbOvrzY
CH6LVdcwKhVp1iI1jsLOOF4VRigdiDCqzgrj5XmBH8MC0SNfDm+gynB1nViNzbb3
CD+dQhaKGcfMj5aZac6te2YxSio+qqWNtyIrLzK6gqZ3MptgOp+VR9FpPfnz+qkz
CAPbjUdmWY3xeU4UVjFWVau8fHySY0R63wWqUnx3vj65vIYNOrxlOIXv20UDeSyu
ur5tlegd5iWyp5Iokq/XMpwRIYa5u6jCfDAYYBO2qm6XojMmeMePIKmh2AkSD1v1
iDUb1BHUh4SocztIfvJPSQayDDMYXNRW2DBhPgygEHIm9BbmdpfqEHMuWjOfdu56
3NbMUtMbQbA6828379TINKnjHwV+gNSmQRp8UYdVBK62RpWKfDqojNIuh7toXeaP
+4nZzUxeDmuqRE09JflsW0MMsvWCQTiwOlivG+ZSJg8ofDavpMnYuzpNhWTQSn8u
Ogg2VlofdHKW6D0XJ+bP+ieQfLF6pVp4/gL1M4AcrWHOqsppWWlKIB8tOANtUxCA
22ZaqFZxcSiN2XhDBdUWzH0aDQmHDkNNQlQToCsjF4oDocwa/9uV+ShMHNAzRFCu
PjfdB2lr9yxm8rkFpLfRpOcX72mMySDobdc8QGXed3kZuML0cBA3u0H+ESm+81w8
8dokuq3IrbJEB3a/BpST7SKZhk9PcGgADSA3TJwlKba8SL7HcVuJPejCgYOloO0d
fdPtKM9ug7wuqMwcmKbvQsEOxFx1B4AJjSahcbr9nMy1qerMoO+uuOHkL++a0Bbd
/wV5Ic6MeVAJJGLrssGEh5uIZT3H8zZn1cEKkjkVPgMvcglv+NK36adggejaZbCB
hUg95ytz+aP3SnDiiqzx80/5YPYnfWAKulTTqFZj8xniKSsqeCgk84iDr4wvHl8G
PXlT4kdE3Fg8eUZ01T3SKtSLRVxDUWkLheEkV7Vzuy3IcY+5YPcNEd7Lvmz4mWNR
e4ZKKxahYzg76pNI24WNwnm5T1Nd4muFnhtz1FI7LWea9T/Yd4AF1mXabQtM5h4j
4Gv+9ZnqG7rYWr2+d2Af1cL6O9v5OWlq/ggCKL7pSTB06O1GRdBi+HhYfp1ergsp
epJ98P4A+yt2H4CXSplnQHYQCBhxe7XHKMZ7dYEhRr3tV5JdsPenlQXrBj4ZdjU2
gE1m1w43huN6t48L3sOS4BklGBsPz0FwIwgH2PQgrLfjmv/ZgKsB6wzC3jf27lhK
XDO2Qwv2tqO64X9XgKmMpEZemxdt6kFaQzKEfO9UW28ENCDbx7rEkWspgcHoHmHt
l+xXzn5bkQy8OSFJTMC6ITa30UB2kzGhaYnmi2x8ncOpP3ev8vsRJE4SF9YNk4Ix
zJBZVXFyArO+6InAEicecimcb4xbLGOLA3fY3cjW1wAUt9sDiBy0WUImWsa7rAnZ
UYQtZ2ezknAhnzWxozwLY4TLGB/hJmnTvmAsJZtfhKsgay8RHh97SeyPoiilrSC/
VoLR1qOrMOX0Cnk2cnNYB0B8lt1DP/YYqbk4VTG75a91q8ighnR5S0mcdAXrAPrZ
OceXu/RHNVj0J5yZ80SAQrgWMQRhyja3BI6sYLWQYAqjtbUVbv/yRISuur28UUKO
A1bEO/DxgSboaGYNPDlf3CJllWVvNG4AFz+GTyJBditR9hI+OW0DvRYkO3NEgi1t
BCCohEe1didBl1qk0DfAmsprN8WoOZ+jA/dBgZ3RHASppz9w5VRvUC726eJi7bOl
/53WH5e8kW9efcuPsl1sx+MHmzIeXoN59AcQ8s3wZJHU9a7gZgb05QlImYY9K2xm
b4/cVs/so/hfSlqd98Epsu2XRxm4vEOZ7VBD3PMa+UOoCenPR4D9e+LpyQQy1aOC
+Erv8xymakzS/7qkrUgo65+dNRoHNSzyEpJgDSZ2UzLK/IidJ+KzpUYdH/vf3HmB
s0IP7Ck1sJkq0hGGn1aHBAE6u1wSi+KfK9Ab2U0isihqViYvoT5y7o77hlzP97CM
RDTDqFc5HxWLSkJlZ+PmPj5klXi6tnMRjJjgKzLZ441YwGjr8V85Eq21MO3CcNT9
i2bitoz9FVNM0sJjaX3sQIW9OzCQePwm6zM8I222O8ZTJuu2Es7spC837LR9K9ff
B1zZ8NomgI/dFoM3uLvyr6vwSSNgK8d8do0HPvJzkyhAws8mJd4q7yxsYTyxIbUD
Ytx2wNZpwDsiQ+2ACf0mtFiZhTK7dtCPrR0k0WvZ553zWW99MO8rYBj/HOe8yEOG
Vq6Gmlrm929/o//VmykqIAo4Oe1wWaTtfydwVcwueMtygheueOW4NQ14oL0PF0NI
80kPc0WDKPTFWWbc5lQ1iH5lRhgYqOgH/SLgj42++2PA9c56XgoO0LqpwxJoZHEN
UCgDp0ZZYYa5mxYn0GKN0rX3UVgN9Kyjtv0jG6Zz5TFIFtGtD2yOOhYjgJ6sofvU
E2QooJz5N7lc55xy+jB1cLfF5EkSJxW2aFw9YYRhVNZEfJo0rSpuZFxBaqDlglQC
Hi9ac3ZkqnHfMbN/i5f/49urUDIhir+K1dZL2nafplp9q6BhD7wF8sdlzdR/avCW
LAAtJ9EV6eFUwDc8+HCg8p11PyGBZzNYRIHGXYC2Moiwf4UZRIWm87x4Y+SGZnyX
vAb77gn90Yz9ZSrTgAhamSv8t1puqpUxg+NGgYFS1qdx1B95U1d3V6B6HOWiM48b
TA8m6bNL6Ce5lyc/RCOuxybIscpqjX462/CSDPHckPkiTSbz/6Go+NN1wKoVRfEX
BzuyIAeTN4w960PModZMaeh4502ikXbNak1upw+O/JltbXWf5WMNDSEAONRy4+Nl
ayVQkcyDQTSBJurgZ7topkwoTmYfLPAzh2ssICiGDN44M0FB/fmF5i4HK7Ci/DGC
yapGBV9zqtSAvrTuG+bofl7ypQFewZ7dEPxkR73LldDPSidPCbv7bQS+kIy1fh3t
M8j1yT3kZrI0QieBk/WdHX6x5+CLBQXWB2lWGaEBMFnL7hXJpRG/Rvzprp8rOVzs
e0YRBJNMNZDmjunVoXmvRNY5mOlZLVd2AeLXKgc6al3VrbrA4BIjCZMkBva++hrO
B7p3T65MiDE5xdhkHgqeYJsYEeA9GniP6e1weZwPBmnZzpDaU9kc1sjtZ1iIggBr
HfL25pTtQidZsAh+ldcFZTu3v0+6XRE1sk0S5QLAENw9m1i6YB7pABmbT1/ScJxj
hzwz/Idhr3RxePLFrsx8sA/ahzxHy51KJ7NG9BMZa/xXHy6JJoxY6iluUw3+Kbwf
5zeMZJ85JHPXIgrLdbwk/WfHOtLN5JbCc55oLjtw8eCkmdD1HhGM5lumiu4g2gAM
nA4NBH8Rdtm3T8qjgAN46SrVepsqBRO2T70vkTTl6oCaIMcbn+3uoJCU06gia7aN
A3QCBclpJyu3TiWhAo/HZZ7KVhGhQKQdpT3ZwPJLSZYjhrVc5BhG+131logbToNT
L4Q4fP25nLYHmnztME1jk6hkmN/TSDWfi58nbOzyqZEcAiPUR4MNHxImFOyP7FUF
e2Cehxg3HUhr32bU3TF3/3tu+zNO1erCh6MTCYB0RxERuHqiK5Fp3ARPnjhOsIHB
LS1pq69uat11fdMkoY1YWQNj6sEy+AQ122I2gX1Bn4hDvpaSe55jzi+vXv00yVfF
lG93Pc/34r1gRyhyZfBbSTxxLLgWJ29sB+TVQWbVubYpQUT3ZsbPfyedKtT3Gtzu
H/9V9l/+TvRAMns/tgzsc3qiJXSaggW6LZL1/CwR1rkELx6qwxaPsSE/ZWt+iRFz
3nIHrYulp9YBqqQGF8uecR7iA7fmWBkCSKzmsaELzhAdhJUR4o22ZwK7HJlY0bZJ
mYEyhhhdmOC2M0Em7aGJkfNR1vbrwD+ge80/VoV1XeIG//n507OwpupIvyWS4cKA
hLC5tHQvOKlTiQ47DW2Nm43PtdF+siTdFEP31J8n5tlmhUBse6i5UKifkyiCnvn2
KA6DBo2zPe/ShguW2OAy9cF/jDToV71YobDVPof8EnKy0Ej2IpDsasyvc1YyIW0t
e7/2QK/7JvV3kSUhNytbkdSma8OJxXBxDSqxSK+5bwGmKczuPhryZ6e5o5Gsk2W+
fonxdUNveU4tVmPP+oGIBnTZM+38+IIb8xN112/HYC3FDxiqdkZs0VE1+MdzmJi4
KCmm9zk330crSanFdHpZAm8JLSUamitw/l1W9AhbAs23KTdFAOszNmrXIb0UjnLm
mPVFXD5DnB/5OiaxjAOwGyI/GIBBqKUnnN70ozRuKrpJK1/EKPn6F0bfvsjsCguz
u7rF8ptWFK2fh+V1+ZTtIQJocDPnadIjJqaUQ+fpnS9r85OaqY7H6nLCewMfnGdF
Yf3ShwGLNOh89BILT0x9Q6/WtoNK6kRkFjQnR0NM780FRLB9hqDymj2udaq3bih9
Kq+Q197ADHlBcGUQMw3sWunVzWF5DR9L81gCwktOKgTmDdlZBqSXhaOjGQwiq/86
GzQgDE7h/SwlDCPV3HDqprNF9aH/A49LTSLFijMlBNFS40f7KbcWWKZ2T25jemwC
ag41ePuPzI9oMmrRgTkKdgDgvFhw/6NYxMN9p2wtgcrYXps+zC+3VxatUNa84CoQ
IwcQ04xpk/lrAK8VBFs2xFUAXCbrZjUBajCe1ZQWw4uaVjRVAq4M8/0soXuA/lon
Vfwi/Ji+zeFQWiYVWebz2uAfC2BWI4KrrzYDvcYxhGeh2+S5LL8YOxLmhVqioIEY
Gdgvw6wQeA3hRV+h4R7lX3K0Rn0XuzEIMEtFa93y4tD0vN59dKp/+dQpG08sTj7M
WyS9YEJB57QO0pWccCXysxpF0I1ppX41JZcoeid9tTIDO6KcpiQcjawnUN0n85v7
IrZLU4Hdikq5AJ3wRhf5XgsJpuqLMXaN2q4n6pv07ipVIGJTkRmeGRut6wLofOBc
rYzRa+2/vPP62nKId0Wi9zefe1SatHMuES7IxoltVk/FfkRziwGXbKotyYqgmYmX
fKJYs0gZgQRupQBUY9EWe326248/KCSBm+oWppMQBfhQoF2wtaATnTXLWLXq818q
sr0y/dLQ5BzbGDncsb003MYlOdB2HA2u/yaLwRxa2Wsez6fL7hG2JKLWwCWUL5dg
M9myEtbkoTt0H/1+xmay5TvtNzAoBER1jGiTVIIVjxA0/ZXged+5MkV/Rqc/5u9p
jQB2EFY7xd8IlKu8glOlRjctk8BSQxRcfPnMpIJ/6wRa0mV3cI3wSl3xvVbPSPrE
sovzZOxOiI9D6ySInJWt1GjGyWGwLvilMmTz75fEflg1xLmfPa6C9FydyIyPPKeS
e0KBbDpr4qYC8rtkOVJKlZVrh41p34Khr3EZVPwMCDbtPhAuDDAhiZRGTiS/3XJW
5Y01w7WSJp3MisCnOFA/YBE1eUS1KIUZsC7p7KEFtrb3v7LSKSFG4zn/bLhAHs+X
lSin1wUYz18cbiG468oKimZW2qWCl4tBT9XtPBqOgixhlTHocJyTIkdZHuOrYjqe
NXUvA+qbafENQs3q1874MmNdy11b1D9dQ589M46y1xLRYsCoGD/vapDPGE31fUvu
ZgqBDcc+AWHLJg5Upha9F5PNo7FnMt/PvByMc/g7gOykytccOYSgHgMMg9V8bzx9
5vUjJmay5ZK6dMeK6w1Q7OTY3s77EaXsp3f5b6KWnEOXvwp7MH5UddrNi2ZsQajF
eajpsLghyI8IT2CHO2+PKSTAM5VEIztmvue+Hi9Fv19vt8qi0z4VUcHafPLX86F+
fugu7iEKf4BJ/UJsDjqqGGpDKZDuO6Sj/wLgIXXgB2qfjQVIsMYw55c4A/iFA8T1
4FHjNqUkFcBhgkAmQUL/0kO4GCz/U+SMyvczB6pxKPbnLklnngNg9LeLnZfB6wf6
MKcQ1K6AeTi/Fh7hCarUfa9kmSTHbqRROUK+ukU43QklSW49pC9KcH0g2qjvsoYn
81JXLdUnqL0zgDKULYoJrw1Xgm3erOe+b3uobQFkx+rVaCkZS4JkAgz3/TtEPO5p
k1WMAN74e4z78+t8HVamvnWM0BVrTqp68rP+1JM9yaeOAKEJE/y+inNheBORHrBH
xvHoUFsWqSrL7XpptafRPNphs8W9AmsXhd8KWxDAZ5m8hE8S1MMXzAhsKJmvol7L
pnpm9BD94h/RvUHbAXsA6nTP7gJ7e+1ATmo3r+pz/k8cjv5xdaWlyyl5G+IdGvyx
p5QQztVy3Do/UUq25hlKsh14WfzIE3RvgxWot1gkG3fObzX1nMeK6P3eRPw5Nxre
LCU4gBGYGBY8CSvMkpicWZf7mg2WgVTUKDi1EUo0jL7QlosN6SvZmcbzL/8W42BV
VQs9S26ZA5/+D39w9hL7a8VLgtWeiP+hq5fUV7Mzjq8gXbuteUWMQcGI6+nJvctd
7UWFmcKL+eeM/wgE28aac00xPsC/xU0nRn29YBM91Lgb+qMDmF3V6nQTXo1dkpI3
p2o3PQS9TArfpJb98+Y2oFljuFZZcJWgdvSa59q46B6VC5StoECGvQy7993+r35/
FfjKpQVA2h0vIJbJBUlB2wgPXQdBrQCPsW4QVQgTRo3poDvApwUaVOD4ek1SdeKn
x38Exw+vQvjZvxm9C22xYPlHd6Pehu0lshANQFL1bhOOsT9zB9vVhvaABcY1suXs
IvsWWjYr52X96uUtGXwZw61cAE8Ob8lX5KGl38VYRDbkSe5jHXeFVmg2dRyvyVA+
a2f3pzAab+dvjA5mbkVDoCYN4Nt1cyMiV5ApHg8su+Amql71I/G74Zl5plP0bbwP
HJzbYB8E+q6XasZoNEN0EkG1Sn3qEP9MDxnoIs94Ab55NDpEchc9Kcb0GoNTlx6c
NZXcVSZLjAcEM34a53NBxZQQaDs/BTQb/L+uCgzGRwiTFHUvhRMP5vsJ8VfPPu4R
BsC0I8ZSYpq2ch+N7MX+H3eOk/inngcyjBzuYN3Mh9N8iZB8F6YuX5xzecNyiM7j
WshwEvNUmVlG93dmW/qn8KQUx7fgA8V0YbzHH3odcEC9AsdaHZ6jcejwQVaaLAUC
pAVshUHxeanJ3fXIwIOIrzXd9TJUxNPBjg6B/Svz1oXoDZzTm6RNsUujPCyxAOZl
VXQ1t9mahmnWgbWBkMsoOMFOCMqzG6ySa6Ep26hgv8w3bwHN7iWGYcPNGXNX/U5T
bzt+YoAf7py/oJzmTDGF25dFrkUpyrdHloZ+3q2rIjiwrHY1wjwCa1LAUfo8K6hU
QU0nGfvHbaxqL3Uit6++RLidgUQUQu5eTjmslteOwvxSu0JOEZlF64X6RmImDyfI
v/DZEqgOj1fgO/P90Uh1C6AplpxScy+WKXgb99Mi3OOZuwFcVHGLKFf7RPWDId6t
/BDSzgN2hJSXuiwOJDprMSMKjOmnVX0Db8cDzj3Ulu1FKekr+vF0T7NbkgDRaOFG
A6QsBnR3P4nATZ39y81zu17fX3fu/0tbit5vCHuPULnkoSQ8N9d3jpwrgU0l6XbU
4hjLbXdNF77GFBptb7NBSttdSurMYcIh3Rd6wy7QesmEnfuipScV8jFxPTbpE8Kx
XTBTOqgQ9piQwTfx5ka/795t680BtKheRuw6QLDxHFcx+vK8xZwD/0RFGPelpcK3
FGIFrPVU+cJyDumnJIkK825G5rX9cWoKbI+RqY00TF8dwDZRg6kh1XIdnB9ZE7Go
Efi9h0DTppxUdkz+U+PBLr8u/pBMv61Sfo7ZxSxB6QTkGZzB9g5XL15YWqAObBNG
i1yc6MqjsSsHTmkJmz6QzCy/W1aJtTlCEhpRw4zdDT4HndPE0nhx4tOuGOTaK8wz
gY5IRh+avZ4cVAWFUZqHG12oUi60yN077xTbwfQ7PhI9LMHVjr8QXdqmq5MWclXA
ilqKxUVM5tvL7281YiKp5v4ld+DNOKwWV2AKqPwV+uNq3ViSmbwdU0Wyia/l3PP+
hhERYOVn6mdAfkz/QHNXe9n3J3djE8A0H+EpqE7sHwgcgEA7PrV2HSy31svhrKGA
ysWgV+ZKD9s0OiuoD4UvzQLSlH/AWIoweiWSowxV+uHqP3DaYPFTwExQTo4xCQHA
d0CHTmxWpcNJvwC2AO/VZ5IjczL8+PGAuL9HLp/hjSau9vhRgT6G61DMPMLQwyCi
Y+A3/6HPcD+W4M5ZdV9o2+qLcUps1NAo0p8pz4K/RZNTMKxhl0FBRGVcU1pmHNXM
sIC+8Epc4joxgDtWP1el54F6m7Z4twAF1n57PU/nEKj3WpU87Q0PKZRAPnGkTyTS
Uk0XdbVelystn9t6s9yHbDnRUX9R+a4RbFKijJ6NXOkhzfaQBEPGksi8gWzFy/QK
rV4aH9igbIr1RdY3xIAhwIDJByoPjqXIorQ0wKeCNo8jBrW/vis4L7GHGxEmMeJM
L2liwXekY/rrhwrlYR+7+rO8SjTRRszUWhiG3vvH2J64JnRRXQavFRCAAX62dcRF
xeWe3O4RrJgk/eEXUtvFunoyhUTHUnnVd0Q+B0Wr5wMX5AvFP4x17XhDwFh2nkF/
bofwsnhbiVlUkHBuKhxT7kdyArUWqfOnWBnyJ8yWWYZC9CXH8hahwg1fB24kpkrF
e/7LPN+Am3gBeyxd98a7/8xC+dDJT8jN92c2N8P/9C9uSnHRPJghfT2lIXmH+P/a
u0/fyt4CmQIy0njgt9ZWqLZ667pR4yM9aR6D8SjFKYMbJoZCduzhEmL/KdilLng4
HRrJLM4AYEbbv07IrpfEWKYKug8+fownPz1u7w1j+NWq9arFU79wgp9JsW2IUMnl
ebi8HWIKFXdqU0qhjiqDm/AZPk+UedqMdd3/5U7x36VdkiCiYDnStXDDl9HmnBlD
55WLzLULrafxCXUCGI/+5wzmJhjhObjGFIC7apyWpFnq3fqYM3VB7+WnH0Wgr4l8
eYHG+szGb9bZzRRjFGy9QNW11XXK0cotQEI0ZYAtrGG21hBN52XHo2MDOSf2p36L
s4e7Q22kxRzuutzCIocY4o0Dv4dVBMZ2vAsxvAkpHLKZjJmfAZOx72Ab5LOelx75
oeywW7TivigZhW7w0wN40BhXDlTIbx6muQLspuC/Wdu8rltABYNr7uwWp7QKTozg
RL49kfNABgbdqrTM0ViXhJbXAo7U/4qexoy7p2/WY2lVKEPB4WN+SY8ZFynLh63X
TreFt1ttT/iefOheF0KohsE0g/9GoeGufiVwLIf67vqawgMitWhrKIN6V+zLDqWR
ZHlZ0jWNQL/9HrmKrN246eacVvRuX4mXwLxy2uajRxBeadgOL4REJ6uR4rDM/RBt
2rweIZNfAKHioZ+sil+topMDO6+8spDkw36d9wfBrW66Hi65TcaTYa+KKKQKR/W0
poRX5e9He0a0gyJSSf9txiYuI429AVX7V6giZ86yLgzG+K45rXnvL3ydDrGYKUBI
v34s4mQ3vnpdNWGwOM+RJAC1HbDTJb1j3i2ZBqloVo63rO/ySi2p3q0UvAfbPUaN
ZDjHdekBVknnQoIVKiBJs89ulMKZEF8heHOXh+8y+oeeJ1Ozs3V3gQDFZDbsX4c9
wXli5mfHdRwdF1TuZxdXDfDzVDrF79RPgk54pHEa+oiyvg7Wi6VsnadkLZbTcqac
+dmCNEJGp6o2uW/hNk+jBf16MhCAwOKhJxLlb2AZm1VkCBrmdT+uv5ll9nOctb0I
95pao8pQfxiq/nIqBGm08Jb0WdClUXSYz3vV2hh2SBU0JY7kXHeIERlgWF+bsB5u
po4kEKG2d3ysgu/mm6a/KXmgu7rYQ0ZpT8W57eDJMd1J1OyDU+ivTUMDHW4PcnsK
n+dw57IBUD6t/+dp840+v9zfnRpyMtZ8KCUb9ufvwEwhfOS6rcZhEDucA3LxeR21
Y/Evv3SxhgnThlWQyW6aA5IQsYM4xp/xNmyBnEvxqNmSF3ggg6q+95bWT0bRCDPB
gzvbdKhMd1sm9ZbA9StffX4zVC9tblccLu/Z82Y1xc2vPSACHrOQCXZRuhf6A1Xm
RnZ2qzStXLuDoIaYkIGvrjF0FsocVGDuvAIA0Aukz/ZvKPkk+rM2A/tpLQrjMTgz
cYRNiN+Pse3CcC8J3iFG3Epuv1To1v2oV7/DqcsjtAUNwTpaUOkMCUNvZDWFftIp
4/308TkVlsjZby6ZCO9ZDEU//Fvn/pM9v9O4wpFuvfwaAyste28kXFaje38hokqx
jLIH/mIojO+RvvNvlbHO02uDmxCzs9Z4g5CIgG0A+rk15qhIDf+cXf/aE/8XJZ3q
U/hP+OaTjmBQh0nqgWmnura5VqprUuhZIcDrkCF1tccSFIvdmC4Z+1VzTbYGmm0u
vwonA7xdyKZdV+b/7cdBTXdAvP8BcsHUvfhDpVtoKcj1taz7hqVEa7vlYsBha5GX
hPLBizsdy3F5ZhDIpINUcjerI/4fztNSSHUNuQeYT2AxJTTKJTZguVsKHjvdfOkP
6hh833nlVwtSYiZOmNN/gqGWCA+EZHhDeCViCJhhSpENq67d2gYvFEa9abJSy0Mo
ivUjzN8+GSab8sqIeX/Trb3byzBebZhEoMsI7ipsQwD/9pBUvSyf96ZHt1clq1iZ
Nm+gM373X8QKXa/KStglqdUJUYl3VAWqLms95cBIBs4LzyT0gjr0BenfMvYFRz/V
Kt3HvFCWQ+44dnjphrkySBqtQu6ipTvovI+/SuI3wh6b1ZCm4z3t7z0aOyzmlyOO
NISBW+zhJIA3h7TGhNoNSKQo5bN6qxLAKZJQ9KQJN4XrQoRAEh3+ypUw8+J+mala
bqBmqFgpx+avc3yEROCAe8BCERKI6nItE4YXxI0854kNGRjZREpxvT6ehdCp0zHh
0mKCantWXhiPkxRSSMlVfpuEm6kESxuqUI9BnwwNV8RB3ubUeNa3pTPhwicesDrR
D5iJVRuc1HxRqyGXQHK14Xz16nXKtmFEGV7iMwC+QYbBaTaNtKsVQTXrKj+mGL/N
1L3Ti8dAAqHwcDcTTKLkL3uqePc0xoOBpE107bqYH0bznEMLhOC0mmSbEBEY5qRk
NYIuD9vUswO0XFXYyLFdEBkrD2S6qofAKqwXIXo+xcE1xS4mcpPDDLB3eFkaxu2z
czAH1UYh6MKsajKqZ0RdrZNFgQOR27eEklISlrnxJ5dfbTw3LZG7XvE9do8TyjSx
ceyZFh652H3V8QQK4RZJi/DhrNyiwU3r5/VdUsCzGpVV2RDLrn9f9tHrKMjQFcnn
Gj9FXguxZnfjKMn6IbWWkU+gGWlAFGSLfns2eUJ62lQFICeBi8kTV+4oZfq+U9me
Q6kStGSTncqyXwbc86pDmFuPSSULCxJExjeJ+IO7tMBk6SG9i9+6xf7Fmb6pfsg/
LHW+WNw1u8UigEj2AEeTTQeTPfAc33MWEwe+Is07VzFMGApcJrrWdb1vj/HL39RG
cXtvVTkrzfgtQ9gXOYthogBvCEz4kkfiaDZZvC/ASrEZcPAz93PUk3984ezw93+h
Yi2TAv94bBQvHxzYV94DZC3xeqS1EWBW4ejWDBocGvLw4MZZxvHfR6nqProxvAiD
pPApP4H1hDhrgaOLcwGNPyzf6ynuQ2YDVA7CQSUd3XfDg6SvJytncNwTSGhF33x4
0mgxs9wreLIpWP04ClYdmFFzd5CQHlk7wVSIfhp3F3G9YZo0InQehfb+n/uKNSmP
Y1fV2wVZp4jd7Daahb8JYObGfJqVnWMsDQfvFLJimACP0Y/Phjog67WXcmEjSUgn
f9F/WGIbJvZJ2CbmzmobORqnoWy9OZGjx9OPpFmfmanWvVDXqym+nNvgIqWNnc0s
F2jfb4w+sahuZhz3Ivp8Bjw0RhFxaA0XryI0wVG8jmaDonrhZmYYGiYb7C/gMXBW
gsFMWIHzZV3dv0jpR82FhLWnpKEKBYIFzehnMj+lg7S07pReLp2XFiZr9LYDxp4d
ggM8as1mQ1eEjUo1JEvIYxntoofg3aUzo993W5KhDhVifhKpdMXE1MGcyFmwWwnM
yfldqwhjO19Y6P6fiz0Ec8vCclHUEMpuWDIiRxWvSRj+bATF46bhZelnuPH8J7H5
IVP7wAZRPeDDbMXfN26pk49zqG0YvTdiBBJ5XaFbn1cxWDm88udIXoFqMzYD2/8e
I5xL/cy08eJIgifLFI3SplU2poP6rKJC032zeLCIIMnkSPhM9Qm0wIFf2ocMyAA0
QcTwOWP6/U7c+n8FeCrzBJR5Wxe/6LtCTGeeMYnDsGScpqZi67qEo65bIUhbTpCX
QxZEJk/97XQnbj2P0dQ6VJhOyXCb/uuSfz6nlKSxPGC/jOOm2/gFHn3zuGp3WFxd
+OHIrxB2JN9KahZ2BOofeiHE8tR0cSeqLab+VJCKzYL5EU571gf5Y8+OI0E7bm9P
wd55XpWHp9ATBvgsH8wkUg0vXGvzxJCMKDcjuo3CFmUAciHj76zwS3mVvL/NUpq/
R8qVsztyqi21OVxOEwWLho/1iFmzXbgRoGQ0X6Z0jzO/YSHb1/hsO/tIBgtt3NB6
CuKe7gFYf7AIBSQexp305mEX/Sz6ZrGmJpPugj1pgocOcDRMvVwjRvKACSDEzA20
FHluABmpS2IZT378VRqErumzxQ0ExFTVLqYUW4Xy4YNtZeIwb4s6D07Ad+ceLc7A
yrBr8qp6wRrYICUhEUu5jQcdbGmKu2kd2r3KLEnfMKJwFX9sjvCVZzqeFlFbf997
n8Y6Pbn79d82cbSH3+GNkV5B0swvL91td/lIVeWVRSc84IFboApQHJnW7RzfZaDe
TMg96jH+6v/EYizG/q0bzSAUhA6Bq9SuP4rjSceOlxwIzwnwx4R4yuYY5H6zAZCh
W857cZrpUDJ6EXx+1NsqRqj5m0FPYS6HxH4SFrRlTwKV6VOnZOkQF9xxBjL3Hfsf
cdHvFCYpd0SmyPqbWyz+ENxbOkHPhBx0WaMGsi49HMfRzY1HCg4+jQFycXqlVHDI
pM/5x1BArMo/ODRrmi+ERtOTNN5QBPV3i+ZXJ+AZ+6RHBgkHpvMZH/7RlWeav81d
aF6Ht2w33De3k1YoGB8AFfrCbtDYe4/VTPv/lPB00zX27pKPbctFXtwPPtJOeTAj
cwdbDpUbYWKl0+2nItZ3pC8EqWHycXPhwDOnKR/FSAP0wJhnysHGlhGk9r9aaMCG
dDqAD7W75CSNSwWf5GUsbdiYQVsEy6wPdY7JOD80hmrSxjvlPoAsMOtssB6WDw8A
xpN9GV2jkZVZhMCmCM4sTpv6usuX2TCkyqt4jHEIluxtj4NiEc1sVitpFpD+R7XZ
fidIGsliaQr+wX5A4/81gvBFCfXV1aHU+lqPyhx5MIwNeL30TXsCSouYq6nMe350
EqHRzLyVj/A8la8El83NbaHoWWV70FbAGEDFzUr+t+BAYJon+wC3pZqoI0hSBiZC
Z4rxlsx+BZ/urlC0aknMq5XlwxD1kqAb1sLhNBs+Pio6TQwUmTm9Q+ZJkblN8Kno
12urPm3orvXfSPc8nIbWxZT9iaf0Qisi4o+W9WEMZ5m+BebxlyXGV2nwnlupFr5z
IHdSbUpw99m3Ib0lrAUoBDOGxtJBzyXVvHPa0cqPjhdKeFZ+hDd4U3keqs5dzyYg
gQetp22+U6W2nmhSTpIjmpSLv93R5GAflxavq0OAV8TeTNLXTIpTdiG1J4pcqhdV
gMjBvbAZgFJ9MSjk4tFEdJhjLljg2DMStaE+JmzuyqxR+nQiuyOiIgtdOLGzu74p
4thTON7Cyk9o2UTHx0Ry+nuzvQnIny+ipBvD1fHgGduS1Juw3Wnnz06OaixuPtpy
E5J9CP2NvG2c1iAsWTr7tcQlxOulP1MqiFxBbdZtwDsyg5Q4on+6Q13RaiwJ2Qut
nj9DhSQAgdeTKeEA5o4mHH+wtLIPnlqMYckX/j6OMmbiDoXz7LJ8aMT8+0M2KwkG
QQZM78r1uvl1N2U7xBwKWSxy8ZmkleftwLfpTpKKuhKXKXDPMHe9g+4u/y9Cyn60
BkLKrkdJh+dN02w9pqJcRWn2jdodxoSksptT500LjssKzzRCRR/1h59I4INvbCU5
Z2tNC0NOgU/jyuhMgZsidrjTRv6IXjnzUC9MjiQjtZ8dY1CsILbK53rxy8idoXCS
HjnYqsKVZYNbL4BK+CZXRQit6+lpZLTejiU9EIdyTqG6z19j3J3jcuTqfm0UWPT+
9UcuB5S56nFZE/Y03gB5ORji16Zi1FuxcEwHGDDRgCK/LikLRnIq6f6yeDhAG1xC
E45mTb2ikiUEcB9IVNMaf8IwNaeoq1yWqeMjtfHKb1wpjV0zoLxXFkcP51oyIX+W
tcZ9HRay7drQq1u7fhO5P0dwQWFM2qiYawDJr0IHwBYautOrljEa5OTi0nONxJne
lH8ipLjPDGGt91b2Ja4DuWiEQwJaIKbHjAghL4Y7zNDZqjzj/ynMR/v0sc9K1t0u
foPPWtaYwaIQwV/GIn9es2lNusZlaRZqqGiT5un6NFjPGAwWYFx1ij1dmSHLxDkw
mL852mevudNv4Rj7CyUXKR4iUcyZbAnUNUTTwFQLdFsc+nUrNQ+osj71D/la+eo1
QHMUDur7qlHqoKijs43XsvH0D9/0b7r+HV0fpuxa5cHYKYBbdp7dnAG28/f2Uf1u
33J8cLr7a5mv2HH6QUrBDKLA5YVvlc8idOE9RbW6bbqnG13ouFMMGTV2W3YMmCvg
IAxnJ7p6ruELiE8TSnoQh54r9uxZZdfunsHZOlXPXTF5j8cDJbHbbb1vpBilUNzO
0MN5p9Na6xz9GyJuMIzVvNjLtpI6qvDuuI5XJQ6lLllhCjzgAl2/Wx1xqybAATmw
nd7CaEoMu6lx8Ey5iiaT2f575O5VQe+U4zGwB4Kva3xC30jUlf/Z0aahDw4/f5jI
Lxdud7NpoX7aGz62zFYbEBGasfvdN/OqAXHabp6YH5GbBi66JvgAAb2l7d2KpIbz
lgsg1N51KYsXIZ06e4D4lO9jb6e1rxHk7cJjdlEhZxcAfCdSi5Z+28qzksfM9Bin
tkM0EG8USeXy/1OONlz2/MuxZOFtEfgPGqSzGaIPz9soP/NkYYbEa8GU50v32jzo
dODwuMJG040ZAiktRj0cbnh4xpWUAUzJbZCY3EY/r1l0X7XYA3ECVB9GnGFxMZf+
S31VsLLWhtXa8X6LmslINz3V9rf4m0Zu6TmKmGFK2CDuDQzfMb/BgGePhBTvr6hK
s459lee17fM+OXEKZEzt08ZdOgnQTLkMR0HMQSQcBsAECFp9CKgrWOTlR9ZRypoF
+N0znYCUQvvDzL8+vE5MyCUb0PhXxesl5bX8L9q/zG5dSKZ9VAWu4wh+mCU0poAh
iGcFCMdtkSUUqO6aHhLbESquOs6BV9uAarD/AtWW5FGPqZsQFvn40kPYJH1/q24E
ea1fUNe7HIHXm9vMHlPficsCxG36M1Z1yyXuPyNbGigneiyrQwj4aBaQ1va9YzOu
EFx6/6820akvbafDC9BbYo4Py7Ytmx+8ESGMzr5/mS1mgowYcwFSvL2Kl2vA+jI0
b//EhwEjcyi3QIHnEyeDBidia3x4jV3DZ7BWrnlSYu8wDZmdfb2OTzGv3w8Dv4zV
3OxE7AfOILJe3gR/KeYl33kEf20a5ytHo8As7ySKeejbYB7WGhNuifQciO4yqQBV
OqWp5C37t6/XyqzCHEB1HjQ/2OX45CldEmogHrsxNCAt8EW7Xcgr87C+AiAlwTL5
0UVwtFGdzqDLojVo6GZnt3O81a61/oCj7ImwGgyufwtUaq8txi8fBkOiOccEjWBo
jjij3ANQX9gNc++ZI1pvKWFIABLbkZdXsdDpHy0CMCxdeF59sUc/eTzIsLroIrxf
jJt3DI/uHL//14e5McrCxg2cs5y71JfAoStJJsoPRtccAsNH3KAhiZK3IJ4rZB+E
qsbHPHpRm6o0H8piBPNmEDIhV9r3eBt5fAS3Reh52QX5keE9bSpoocNF5XQpzIvj
HW1cDijDKCu+l7mIy0gEkpb31SBUxYZYGTAB772NJRj7s5PnR/YUz13MjUts7q2Z
LS+Xzaer4sB7j/isfHgJzE3ZvkHZt+ROxcYwdz5/Jl8VSMaYtoXi2vvCqhwWyYnG
rsa55uJMk6VAH8Rmlej4Vldggl0I6X8wuBxRhaGjx/VLUTZoEr4QWHvElr/j9haj
BYVDxyX/vs47QcJVbEX4xn3zK5zqUQTPa7X3ZkW4uF8PeZR8V3ZeeffVjoBcbEE3
CamZtMYP81WBDT+SPum0/0Z9RMVgLK+yjhJFKGmCpb9ATnegdFizAyY2ocAzWzcS
Ayzkrq+DU7LaVnMv2R3bHjZNcPG0QgmxJQeo2sVTImH34VauzuJz/PzoQ69ntlPa
u/JVay/vsjHNce2KZh/QQ9S9BphmFSbtZWG2Maiijy1nyG22izxO13OlhApSyYj1
E3IcKdT1pMEi5mSlUQaRWCZ6rBQ+ULNGjsgtNJ0qxVrO0csrnnYXnFfAyru/OLRq
OfhTesFYRGTuJmTPaOLb3m6VoWBVcns92BR71yAyUEJq6srJvIlVdSU8J5GkoluV
jSK5t57kuddREcwUC0RZ1ZXPLesQG32+mQi/KApaSz4K3rc7TUOvUZ6Xyajmb2dj
MQAEDGQQjqhC86jxcOVKuVJM2fpzA2+LdxBpghD67JTqTchDr1ZWAcBFeQUX8bU0
U/wJ4gQLaF/XrsIjx2lnYMnp8cesU6x8TMpUAfJCw40+0U0/V3QW2Ei9e7H0Fsm/
LW3lzk7W5o/dmS0JXuNyAatWr0URiXYIhp8NR/gChqFLUOg5eHL+lw8NHB75w+EA
Zg+5ygWdKDo1JkV03c0zTb7X45UWq4BjIE8NmdVBMXDGcCsn9FLH1gxPUUh9ZpEn
g1777QPKC6mabRbMA0GHblafisJ8SvNOEm5xCaT9gLHX7iMleLrBIL0abwlvVcae
ZpbiS+mfaDjKBe0Fcg+ZkvD6s/A9EzY4LGx+3IICGwsj49/8nY0mfaNnqFJB2Dca
RO2qkZX3ZtE93+CeqT3tnemvblPm7eKrpxe7Edh4C8mMZBIuUukhKd8W3NcVOAQR
6jhCgKR3Rr0HaeLFrGXRqiuJxqa8Gr4rdVVdgvfOxqUPJ/vDyMCkPY/VAwWVuron
0JSImZmpHF2miX22kK+sqdQkTJFbxCJf5HQlmWiByrzFlp5auAe2+Vodea1Ap82e
gSi0jmS7CYdKVMzHMRrPs5MPUtSqpMSya74VtUA5Ca3NJpE/1ZkH7X9L7MH/0gwp
BucTNVSPEPKhdJqxfDb0TrnpVIE8hxjchcno+P+odFQ3fXC87lSuPUEwvAmMdiCS
JRGtszHYjBSfXY8ab0zXbMmYOw7NDSGeg8I4Rc1CqO0ILu8tfkkKjVsHRl0CfQT7
hea4TxAMRHltgtuR8/woecWySecn4HfKLQ8yvRJAoQW0lzFFtlmNgHyLqseagthN
+QfN2iMXtCqhkk0sciuy9kSx1IhtmUsdfwV121UOPNunVAtj9Mgy5UvsuyQhSEnQ
djQwNkSLQWyy2qEm67+aWOEBAhx4Hi7je3ZEAIY1rDQl7Xrtu/bOceIdf/eXMQwg
o3cDWbXmqi+cAxw//W1OTyayZ8eTwDDrs/U2v34PsOlojoC688l/jO0DaoQcMNkO
5hxaFVYLkWVcQvEMnfc0TCWcSZX3+OM0Fd3qCWAReFSFBgkyAzNFAv2ke9lJJE3R
8TpFTq1P1bEX8oDXKDDnauKfzYNHVF2/sG2i1zDYNEs7ZITK7HAliPtYT4SWKR/j
IhHi5lW4XVt5IVeLLdAsmQ2Q1jezIN5fFw4g/p5GyiNqnkDM7wsmqzQCoisLEvPF
g3JrqomSiYQ7HWTfdfds4A3GSsl4IYFg0DJxuH4ACf+KgeeiNaCUT20QdrNTPLFY
xKe79lquop/0H6Erszz2QYCJ5pPyb5Y8mP9UEwPvbOoBw3HT0THuCoCmDvsaft2m
+LyEwCbPUIQd7T1fY5wrHf/QqGINnRIMM6HUccSO/a05d9ILjLXLSUWiM9G4j8oN
TUGVqJCoWWT2t7NzGiFviKTEsAHNNp6GTDydM58RGLhP+NdWUzAn2e1E+vGMTzO5
5COJ795dSRVAVaCu10LzvMaluhzh/DDeQ8CS5SOIYEeKUVSXhm6zN3oQC8Imb9pZ
UGCWWzgTfgcG6F32xxRZUJK9SYw5ekca6WMBCTp06Be4mMaIGZZgs6h6poux2V1F
jsgh5Jzcrwq/Hlr9igN95Qd7olp/Coan4xDhrm0TkpvCfqhAwQO7h4SwBgxKvKbL
EVpHOPFM7uhz9dhCGrh8ez9TYohRrjtBmx+yauNb/RGONXh397MEllibTonJtKhc
Ljy2H8+ebiPVtndb6lFEgLYvTsNbQhFVQu6rftuq3nNaNo/+N9+oN/zr+v63iZJQ
3nJNcdJgsrmRV/OfmM3HG+4yINyNdZaPwNRxgLgbVFpBB50zytLpSfDL4wHQzL2v
EZ5dTRJehY5/Tq6AkdjCd+oBbrcJXRRTpx4VRM6BC2QU4hL7CPyWWaUqwfF7HTy7
358AQlhDCBz/LtKuKIeaSgLCoF4JMeqSqCX0TgOQrXlzsfDbIFuy0h46Ici+blPb
FUv5jrAJhPbcZIuBtVwleDtReH7qYPf20jSPBIFAy76rmmC7V9Qy2j1CLW3xxPZR
Rwr1Xgun5YAdebZdcNJDUZ420FWD7ysiMuRaTrs1KO7PK1jCP7pHZLocOAMjcDxU
hG7lV5Ltnn5j+rjdT+xfs1TMGjzOW7hX2SnQR77IofU9lznKNNpzaxlzOled1Tq7
aQ7kt2cPNp0vnAlGzqIa9PPTod1neipcNim/RPlGw4k/seAMJ4Dldx5AHA9lQDUQ
tfh/c+0Mp1JFcWsFOFSJi7KNgk73MTDEiBojBzGT6d/K/HYRnJX3csdnZKepVqkM
bo9s0kSpxFSY9j0rHGUjk/R/ROtJhANcRh72xlaEDLnJBBmm3nhkSOxcIDL+W3lV
S6wtv3pcWTb5TImBfJ2uaPMbgvvMpl+V4+sRPeJZsa0veCDbPhxqorFP5x6yR08p
LPo+RQ+UKVrjHFd2DvJa6U5Fag8vcA/3ZNCta/+JWCKVrHxmTB0BlQF7sXsWvZbf
aCp2U5BQ0ohWym7EY2Pdn+K5oAU//OZhdxoC2Kaw0q5jaRjAyIC1d+9ETmf3PFCM
wHx2cG+ugKEC+PBoPamL21rROgng+yz1GBa+uB1SawAZhPPRBde6y0hlaGUCnDCN
FYDZwnvNlU48YCuUQpf0yKCnY+8tglN97C50jv9glGZA2urS7BH5yGoznEBpJ+TH
9WnKqS+Axcdr4zEJcpisx8ElzKNVcaG+1cxvyqFZty8lpOS/2g2nUGb3vvR+twCr
EPBf0A/YCgn6c138Hr+SgSoSDJN9otIx89GWxHL79iRCYkrzw4woHLlb55Akc22w
ZfbkSl4o47HnLhtzgZTgyyB3vArHx6lJ99U6dSoYPX/QHe/YY0Nd5Foq7AvZbXYu
8AvnL+BCsUlufHIvOjGMxrwsILk/K99VN2oVAnDmeIo/bFepRKwuqmqBx9yOC0U4
P0MGrmPyPIrXuWZeiMp7LmMZZ56vQroZ/vR3dkUsgpABCz25g8YYmzeeZHmM2ITj
BUAOO2+5wEo9CQ0MFT+y/Rp/JEtmgFb+hV9ANfl3uK96KnxOXyxlVf6NNpYP/Snx
+x4K5jiG2sFCW7jtDwd9j+RsVwwj2J1oPzS7yBsBizEqUF/KOWjHkmAd9y194hmv
6f6IxXWotI4vxfTppS7TI7NltnMlJYLqfKXtLXOM8VkUGQJ10LuInG+5lTANFUt8
dPcfjcAlFPS/5wcMz6ojDuDoRLgeCzAKzydR7A1j73f4YxdgCx2JmDLPAtCdDIKs
kzW9AQYtMc/9hDSQAy2TVCLG/CSo/6x49NPQwP/4Y1L4esPBxwdz35jMOIHizm8B
gYxYl+v4DGNInjijYaxTdab/8fxe4w/yciF+9uWh1nX7OysNvmWy4VuCocn0jtGj
5xcRjTBAGPOIRIzlcydf1FDAQlRVvfg+SkQFYCMPEf08zH/G0Y98qqmp/y0uXczm
RyBZlhMgAxQks4pkyqrKD+zbjHhb/bfaDxdo2WDIQNxdRjilUr1Q7wkFt7sNc4fi
e7+J95wBZnwcTdgnBBzGCJc6w1kCO4uDiXxkMwPZZW7Z1Pp8iDYiIP5/EmUckqyM
cnJCOIeg6jRmgMilpP+vT5ECy51ZWlB3YqTjIIiiJ8FnadIz8d28tk1a2du3OJCH
Ygwd1hAAx93yaLXqjoTe3F3Ujg6p2hwguOuc8eKopENJMM/22pp8OQ1YiI9g9+yQ
7oc4XhANGhmjG/DFPtSN2SF8rnNMg/WnKm8YZk8ofN1rpYvPgB95KT5CZ4wzbgVe
6VvggzG9CT6cedVrrufbqKFHkxnbZ4EoIL3JZpa36EoQ3xMaa4RQAh+ly6n30QLi
Z0gmljU8046CI9rlWlpjv3cBwpO0ZfXCX5h6yZarifQ8Ui7sGpBW3REz+5i7eRnV
zo1HnGiLPpMMRyrbc950tND4io4csbFgo9N2r2vmGdGK85ew5/R1NhhquqjMvkEi
KqM/Ou3iSosMWur8leP5IjHJKIxMfghU27EOpHo3yBwrSp0GBFUeUxLRBM1v7Ayg
o6loDoBtlxzFwrN/0cAA9DAtmklsmppnINnStR8+94tSsMmg0sTUlK4Aq/m952Oh
HSnS3Z5eWPX8/y7vOF46Xsw/rp+yz6pbm+olFXKh5hUmDW8g+A2C3m+WVxxHr8i7
zhR980xxwQVpvWkeYsJ0YOG657oo7Fu1+tLhmB4gKMBFORtTwrPb03AEjuLQAgVy
4fPt7kZz8Uoop1VFSriq7mZ4RvZOA2ye3RjLBjxBcq5XOxfTxubHVuX/mb7hgH/8
xRU8vnNgI8GqOKlhtyExo/zOcmShgy8s7JZnNsG2rLGTn3Y9eADZL1+8SBUj8caW
qroHetMTBsxFHZBgPI/ZKivZ1JbCevd0ix8uT023V8xu8rHwnYEwxns0KkcJ9hbL
RRPUWjkqv3oU66ARH+KZ1UOkOG8Qldg2XG2GypWXe/wMolyJ72S9e/pODbdQerxX
vWbzwDpZJYfaKs/i7yxPdzmNYT2IFbIJdfadnnnFcf8h4jW6qv9PvsjlZmD3M9xb
T0dWb4d/ZYcKchuiK/8ejkj9e8WgMyQ3y9B3TLX+mHJxMUlOOb+Y274G8o+ndxKb
CzbKpldUAuN181q1GxLN5Aurdcu/jXoVmRDMqqzP4mxLsPxL389VKwofgATqR1l6
dAjD5KYXRt2d5OkbNYtG+olYKuF+1m/FQaucnxElIop0hiWNN8UIqTwU80Gh+hGN
59vfvUPRAc53g2hPYcs5G39LkFypvvUR4PeCGZsGpphSLd3UjBHS5CbXjfyGgRf5
q9WIkbkHAH84vWMKkLu3OZbtGzu4iSHg0A5/DsKXc9n8tM505U/Z2bMKAieJNUoO
wGJqE0iPCAFeHkoGn2B6j7oAF8JmB4a+bqzOiLQ8j5sBF3OnEMcDpx2Nf+Coy2C8
L56eA3WixFIJm9A1p8sXO4UG/QLIYvBCkCKHXW7OQzuDddgUjR5D8m0+4SwzDekP
HNdKg7KWGDkMVCx/XUYLxS9NC4zLL3ss8al/8I8dinEVOIQwLiUBEZmjqhJ37Tzf
XfW+A//XrSEde7Mr+lic8Ywe2TstPcYvm2dDM6JaxJa+wVELaNk6wxeCdBMob2pJ
jMwQ9FLI+LB6UEa5rZeVvZKaCWBLCfENyV41noCIlV47i+V72h1JFORAHRUt5M3w
GEpGWbFtMXCEAsCnUnBV/ClqNhlw2lGd+DWlTxsS+O2gPNCH3OWYnu0mSltFsIQ7
eHdzgl4gGm6bis0wH+QuRBkoGYvwmblXQEX8ix+44kK4ZkHvVtFAZepeMAC8Q1HB
Z18mqHymyR1GOLS5NdOQ0rwc+u7wYh0tjaR1iKu5fV7IoSLM8+Vgl8znQVrvVfgx
iAJagnDeajCBoWrVOeb+cralEzshhFsKpbGsP7nZY1R8eLxn7ieQx2Gh17l77vUo
FPzOpbKY0ZOlMIXAxu85S2flcGCcW78JDd2JGUtkNrPtE0wBsgY7fnKF/XWsJHh/
6jAfmPne+yv9n6lS7uK5aGHUBZzYVWn3oe4bvofqN5Gkhy6BunraSyVZx0DaQCxt
+aVo79sIHmWnRHEJdPkhxZemzGmT3jRJyoxRVUj2kAeiM5LWk7U6M+JBLLj8hKgG
J25LIJydx9n3EOQ/JA26EiQZ8GC0VNzVy7nEbObIyrd5Pdp+mYaMRbFmNJuHgKaM
DD/U5upGcAGmzKypKMfSCAPxkl183KF2CraVowRU+x462q1IX/tGkJWDrQYXwjgy
DO2m5H3tyxHU+2un31tA/PMchhITPA/HOkcYyb4UWn7/SeeVTLKe/XK0sp4NW+LK
6ifh5B35Xdq5dCziG/TdlWbmhH7BMsu9641v5N2J4vZJA1lH18E5LJe0+wXGHNRf
xY/GT6ZmpjoO4uQuz0aD8dBbezVs7PEdEkoLGEIJy0Qjcai9Sqb1T8yiwfnGYa07
rFXcmG4cCDDZXCStqorHNeu1rqTvvSOQiccHqIGUwrm6NrXqWphNpMCn6naWsJzh
Dxm+e7Y38L3SPLHKGIhd9tgaqpceobiAwW2iQQ/LRVULH6WdGKGEhPJ2pvW3VP77
WmLZztEUowG5iuUpBvPISDPquBKJlvFOAHTwxFV1gwzBUx2hyn3iLd8bmiLSZK7J
ZdidF80NCONBhEybCDSID6H8Az+uags45OASyRteAW2AXphsfph/R2XzaVv6De2T
ZAmQWuryXu1n4cwc7dqW1T575ajjDRqbQ2yYhmJYF8GYGRCkiXHSdexvypGJSdUi
LX6IiNJRn0Hklt1HNBz4ZuV7dTM/a5QY2XuFfUSzSEYtMe8IC70gaaT1JgljfBRu
lFSNsuaM4eFe1+srUrCu9Am0uBNXLFR0+RpD7rheC1uNUHrxnP7S3hhT1Okn6iai
JGgjMU61IvVX6tOAf63rHpDemLs0bG+sNAxNiPJoHvpbQrkkW9xa0xn/BUkaOzAS
97DATUgbJJtG+1ojfn8FtC/7d8McRqi3yAlluLmBQvUG/ujJJVI0DQfs24uJrNOR
Vs5vCKO88bq3vPfgVRlUCqVhV4nFAD/3mifO3ocG84X9nJqV+uShx9aKpBU5KVUf
eHI86DUVBykWVPYeji/2nJOp+WcZOzuimY/VTZ0Y5C1RdynEnW4Uo06TipUa+Z/4
gnJZpVRyGwdsM3cHWkIpGKkD1DpRnScrkWz8Ncs3/+Iwvkh0F86MshP538Mujevz
m0K1ZSPrfoDu1AdbyQ6u7hgYhAcV3cR5PR6TwrZbVX9Y8Wb0VoLY87AHFGM0wbC5
41IH+i1Vt6d8qIp6c+AC+w0Ma2NaQQgHV/NbK0V4M0rQ97RlBWgmM8WachfsUehN
AEdZdEhDiBMb6D7sjS3ha63Ky7sUI8T6LmotlW+KdY68yBhwqGnQLbIVwRmVpgd3
3t1s0z9NO7rpbzkf7KSW4e1PqYpIZqToVlXpdFYGNCvALbtTEA9eOAhv2HWYdSlC
dOPVPwZGoFn598arshWKisjEj9dZpA1W6J2YrRj4V2sZuvGD37+H1FGZ4/h18TeT
nrVpeC2oOysWK3gLvNPa7ZDwBPcN0O0cjDw0IH+o5TShiWUXYTgXM8PxviTckLuo
6AqJJTwRtm1NANMxN/hET4K2A9PA/MDb+StrUxUHEvwXK1Yx/hVFjKb9OFZbWwOY
9hpMsSDtj8XbdNc9tFz52W2ek03kFMfffN2vPe4DC3AEbJ0t4AC5omM30NGewb23
d9WdW3qN0eA7yBkMuG0xauvFvFOPSe7FH7AjKuT6tg4Q1yjxUV82SLqlNeB/u0fz
Y93or68iS3g4gekedzgS6Kd49iYp4BNK4VQ74V6FUCWxkXQGmTzj9CjeOMwBy8mI
7fRHjqsF1T1G4VHiBxoprQ+8EPkZ+brQfczo9dmQgBH4x3UND9ecunKXeVthv2m4
h7KqJt7w2V7bv7UHGvHYz7Tg0Sa8XFbsnWsal6PAXcyORpNBossoAiFpzYehsaOv
JOfM+wOHEuNJHnL7lTnho3WsibByM7WCJuiFHjBTz4AL8csbblc+S2pft+ZBC/9t
2neM/ZzYFKCDXdtfVz8tB4xAAtpFIed/pW8xxmu7SAcoxin9RFw6VrQWMGPkq7sq
4hsEXhuwga74oed0j/OoRW0wLSDeYzfoQHLURlxQ0uAeT0x8tUB2qQ5kf1n9uqHg
GKc/tsyDqjGLpU3819HYvXnurSiw3ADaFgNiJy7vyYqRwjPvzP7klLrM60X2PMG9
v0nKEPRkjzb5KNKgGtmim84SJvhkC/XABqRNiA9IX2gwEvuJ+Lr0tEYz4WsEOgOt
jIayf6ypHSwYVt/pi6zecZ5y6YeaCqUtKni+AvfFFWYSwCtm8RS/i8T268ACuddT
i9GWPrkwQMFpQuR2L3HDg/uhF7JRW75zV1FuIdtkuqW8zBWmo9UjxFdcvad2AID3
iQe0NLyapDTdnDGssBEXN/XNgTH7LQzTd6eLuvAYoI0XE9oaIJ5bUDBJeYDdPoMI
NybLGPaG7iGJllLg9gY6MCtdXhx8P1lTA8qtPNGr3fm1K8PU2Ho/MhTqV0ZldGMo
0VGhItS93WWlfoNnHsrcZA8+mf+xSzAvD74W4HJgbHF+VKK6MA154jGIiAb6Y3dD
LcebMvpvxtNcpSQCyys5ziPLEjyAI5YoPse4EWtWiv4ccsWBVESTc/VfdhHhtGIV
eh+sR684OUVLK73/89VV71TzejxbBHc4fcx7XbnOm5R965HI9lhBZfv92J0RqVQ5
45ew76Az/AQm9ZTQ3Kl+ra/ma5JpLXmLwZMeUS2D6HMwKSFYAv37epEVZPbjVS4D
jJuatePPSn2G2B3WUkVLdeDilh2jXBOErJSqIgZbsCs//9WfTTyRjde3FqEyBrYr
HOTYBgwq4Pmy7JFqTC5luweArm4EDp3GT4PftzWijZOktsrZ/IJZh7WsuMkwXk4A
lIxyjV4Me6qfxeqDfmpNF8u5qis5gzKog+/vbDuWTM/0mFdomaM9j4XGer55B4rM
N7NJFsw/95OF/PREcic23gWLqoLsESVEQjUUdRy9+aMIATqPv/DXX00ed6mbnT3X
i+vLDfvw2RtajxFeYsLim66X7+eyoXFg3nW536JpbSL06xpqpWFZvEDRO/UseWb/
X/550Lka0lIfvr4hc4DWBxm9ixvAOz95RUeJS3gJmAwdkT9JPNS8jX4/4loBH+Uj
Wazwbs8CUNBkG09pmHkz8vKqc/T7zrBJ58vWyNSrI+RUILNVo3DgxaAepsJPyZkE
EjqJutt3VN5KJPzDhRA2x0SvK3NQAEiX3jDhMNu5yhQL/4jCukH6G1AKrxn+wXdW
hNrGXq1kQHQ4h/Gu2n4c/ePf5/PsJcWxugmYsXfnTqG1GDlX5FFpK6ZBOGUwBQkt
jGD37Nf9yOe3J6meGNk0QWoNutO3PjVgqcCgQLUf5JkEAyxo5IsIT+yW5lKhKosZ
ap0qIchM+VY/DTXvcoyl8AfFS+4xL/i+fFI8EnAbstIDCnaHXbcIfvScHnXq3OL1
nKJHC12gPCjX+Ifpq3+3ONSwkdVWhQcnTflBMnkErIh8JaH/dNldjcFS+mrQv+VS
Pb9bm2MVidS2ciAG6hempd/Jtxqt7Et4Uhjyg8S2KrVAKKMwuITzXdKs9jf9CMai
nI/qYaVRciXONJW5gg6Qbr7hM6nqaXZqMBDiwScuQjc/jSrSbo/y5wUqUbUKIeGC
vcFC9rP95rAvhH9lfR6egIHhUJBPpUKh3gPiRPNV+v8Ke2LvyhkI9wow7oLzDj1Z
TbAZqupb1uoq0r3USt8W2FzZgRZ6RhJKERdRek8SRshQTvAXi+PAgJCYWMBzQd/T
jgvBx8izT66jg5qh3oj3C0sTZwjQ6Y/3Si0pA2RrIuRLfC4ZdgEDbeEC3ykxp4BN
ovXMpM/9CCNnhVGXwctlnUs3jsTj7++6nRfppIuCvWewMGz9J3WEsSgR/w+NtunO
TapBJa7V8bp6ctM6L2U3MtgfsdH2cIw31qEq4+jc6SGxGUFCMlhBa7v5KsFu9weV
qGn/nwkekfqhUTI2fkfxfGBMyYnwqzCPBM/jm83OE8SPCzv6Dhcwyj+/GJl9/8kX
3MJ8wVsRjMsbGjpIx43HosgbbI2Eueuh34BVy5ZQTEAwcD8C8CAkwRYMp9kbz+ZR
w79PaQpYKdL5EqTVeLdhliaVVhgqgioUrxm/SOAUBg/rwqFjc5yxy2x4V26nTU8c
ISQK4hvghsZtqcpYyO28yzRifHvKZmgZHhQYoUERsZ42dNE9e7MHmf2B6GJ0TEix
38y8itIZKMVGZCdbKxaabDe9eGBBmQ2cRcZLgdobnP2qZaLhoxYRWZrSfcoa4RCb
Ktzxx57OSmslRoL5BJC0B/j80L+dsOmUaoSuORCJPLqngcfjPbNwNmK5EpNiPATu
MgcG3snGrlpWnKEZSisHER+nr+1TOPigAdQXX2zDvIGAK7yJtoEOfY4iq1PP1yYY
BSOVDpOfXpueuNlRVWtyM3hfbtTnTGVOh4wHb8nMyd2P/WsGuw53fS91kGpTSPH4
Tc9cUGDsI0cDgHt8llzxzKeLO/hRssZ4fVKsYj0lCa7TJLk+AIGe4xuE06sOj9w0
6wCMqIRskQq6WvWhil+i4Irjy3amKCiLmedfBu8KC+aG/rLXKiF2y9DkDjbuqv8I
NKkOoy3QG6GOt61K84eXRcdY656XXLhwvIzWiTAyOw+nWxOL4FXs4eZcOIneQz1X
LSGCFZLVtuTqL763U0XkX0A2jIdxtg8te5wAdkgkADMbpoXQJT/TdKmpCawVUXbi
ixNyfMU9GNjqnXFPofnhaweQooxwmSntIUKwD6AsJmVMBLFlt8ZWSd0SMQDOGcFS
oz6TKgXxuukkq4yFT1ZnqkMFKLb47KYXkRi3N9rsMkhLl341dfWXDMfwqg3DxBS4
TbhLVjAcJi+A4JyUnAbEUKkVA2IGJJUEXfg0jcj02K4GI0oKLk2sVIi81u8wBUy3
pIfGtOxIJikCj/x/Zo1C9+Xp4gU3BopEshw46GVFiyRj12wMF/PGwvBiplFlIChZ
px8N0Mfr1rkZNU4EOyD883TtLBVZma3sAOTpAMkrnMvtD5jb5fgB0NLmXyVmVOmo
lze7E1yp+WBDq54H2y2JhZksKKitlnDkFr6wm/N8ze0j3KYQJcKQTky6V7lu5O7j
Qd2XQpatNIAAo57UK5V0HlAAlhhXpUOsOYmhm87clzXvhMWzWuLgMmxQ1QCHg2Wr
EqTikijLv6yktrqHSKTL5nSgF5yx/SO9IifW3dz9UdJuzXU60MV3qegsRp6TqAZ5
1XS/KKSx0WNFordAYO8qINNxCl1ZNRemoi6lZ0p8AXoN1fDjO1KyMrxMumMKebb+
foh4PqlRgbhBPvbKw8YUXpmNnIOAoNG3Eg8/QFJkrhsXz8aiZuFgQtSr9GyihUIG
ebOJ7Wd4K0LzNjwoZwV+6hssl55CulexGet5aDGWKwwlcy6t8UJMR+e4C9BZAWpg
5yeIbmPaLVYLCDPPCanrXnBGRbzmj7eirjZgCjGAScoSiA/kW8gfraOKfBwSqqSi
atnz6ULCFc9xwOw5LhQt7862PSuc/5TxW8YSA4nzW36l9L4EOd2sKYBi99GC+y0P
LPBS2So2I4/+/FdWoOSlEE8BupOF9WjXmcwc9T2KsvIBMN3Dl+IACNl1tIjG/o/z
Tc+EZFP/zlUHQb7IQKwRWdTAlP9kMR3qMb/m2W9UlDG2eXYepGUjBydKnZwDKXn0
oavH0V4s3s15/IgNHWXco35aMUxN72aiCY1KCh76LjUgozf4tzyji94t4op0Ia+Q
QSCQWyTNMs9nE3vlKQCbFY0f3JGEAT9wUXnaduN1nsbCCUjJwJFpe6mMnVeF1O0w
m3jG5k0IIuzhmfQgdlQL60kyC+p6dXwjs9vX17SSJddksxx6d/ipg+5iXA+7IEo2
7h6YlRo3vHDDYvgP3dE1A8uojdlqaD7ubZRErmfPd30+cavDaxDM12GIne/FHpdq
n628IiXeMh7pSFYv5G4l3PZzYg7OV7AqJhdgErxk0IJO+gylMlwZn0nL/BOib/gL
daX1UZ10dSZFKt5oDCevjsV2az1BN66FejXTYoCEXyAV2c/PUOEzTBysvjUef50m
ZGfLBWdzrx8CWQOYmhFZKl/AQQ7OoBqb7V+rDXALOxPRaA6sPEBaSQqO7jXOoS1c
aF1bPidGInyK3hdVBJo5jdJFoNAr/nRt8rw0Ea7YVuQmAC0Qiy1ZTFlJ8AcB6yyu
PnWRCYt3pVmNl2dTHO/NvZcFD/uiWVpP8okBG5k7Zo6ihthz4y14ldgRM4AVdWZh
llF+ZxSduk7g7Rx2fYG0qXTMO82uad7FeIE2uCY9S+LGps3QQba8ULaqiucsEzDG
ddB8iXSXmxtDL3g4R6xuNmMZxx5RvxyMBfXp5R5nEtHJEoFTJ6qPKFTVA94Oz7cR
w1HvRNyCJzD89wgP8egpx3VtvtfyrYe5VqNzBFPtlCJh7ZxOUKBrw1NxM3Y6RKSu
ad8mvIs+p7iNLW+Yp/vbIUC8vueCaSbBbmEuG/EFrwo1wMO4DLeb0DXySbex2BeD
c/t9AwDGN1lOs4TxN/2YUEEmJcMN+NnnLHEA39wNpZNUTbpRd6IAPEIpw1dEXRQ7
XX+KOxw8LOVh6ieT95mqeYf7AoNcWCAvNBRUzx8s7WDYbGVqIS3l/9lURZkyu+Wg
RhU6JYWcSa4PveHKfmhEyrt7cZiGp+hKgMwMGIjd8sxjipE6CLAan+sEq4ou6fHA
OCObJKikwdDmH9OzEBW3YmZn3lkGUCoQgb6RdHIpg+UJf8NnnWGEhxLsIy1rAk8w
4XRGZxyLEC6mYKZdBDsiYzyiFpjFLsvdY8YVwG8a4ioIKuk1tD2goIWIM+3R53Y7
rq/J3l5tI58zVSYECLX7ukHDZ6p5vhKcr11S2CLcLELhwgz4K2y6Oy+wtYDUfrUf
HgDTq8KasNy+9lqx0q5BvwD3s2PdMAeZQ+3kCUGayxLiEgQ6agnZ+D6B/ryvriqv
nj1TXx0smKKGuObF0Vp776ECA3kDngx8NoQScnuKf6qQ2yuAfdUD6bpH/r3UAe6g
gVC9IwmF/NLTZJIZz0giYZwR6PsGb/qhthNkPivPEpNCk95GPSWJU10xOncsacGF
onwbhj/ozxDnqS124MChZpp1XtrJuHoT2YdKboBwfU1TWRBr6Nu8lMmYNQgW0Rd4
wnLWEaPQs3+FVdGLbfXlbKqEBcjt2rcUsePeLmhh11eg2caVGxpy9/so3Lf3VpDm
JfAcofK1LtbyIPpJP2LDjFi+onSTj7dCjQNCdHdXf/xJLq0KSCJxFboUcoxj3Rde
Mj2+lah1FvjxyiLO1xxYtUb85M2PzYiPDTnGumEu65Y9UIWAcUainO1uQc+TXHuL
ESlszqJH+o0Augyp27Hcq1JDibG0BJWK3lvq8ZulxZuXLvRqur5jV3g4JvPS9hAs
iWdbMdalGH+1JEe8ns8Ob/YiJ3tFY9Z7cBA1ZikGubTcIwGxnEqo57PU7soeJ4tv
sX+gqrtAsWXN2+FxgPSznUIJA7uBCMuaYQflqOD1XJUIdQgM58bOm+hPDkLDlVF6
6MXAEvQtcuBc80qfTsIpWvt+P+/wsh/7Z+XVGI5UPQZKWmwdzpG2mMeY2Xtulllh
gYjC1FT1kTxokAsWHud+792PohkJas0CMKYHd8oNRlNmS5Uu/9s06EzocwfBT1Jx
HYoL9r7a5FunWhm6+8K05+mtbx3bwM+qoL95Hxoj4uMxdh5b5E/Rdu5G+tzefCyf
8hLv2nAkOaHZzN2L3a/mEyV4k9EefiDo2Buzk+im58WfnvbtEeuJpYJNlrGF0+nw
3d1FOhprinNzWIp7m1LD81ahFTNjxUB+bW13wW/cy+rwyD/wonQPwfJLMwqzVBvl
dydW0NTMFk7r3hMnZ3C2prO0tpLq9MpFu4zAiT8S+L5TEzl90hlrfVLJfxn7T/ff
AmoAL32bY3QozQUdTzzi/o/T4caZvJjUbP2v8eyfLUXiQ0g/DVd6AFnEJicDSLOa
XmsdxfL5BnQuzq/qU9sfoi5spb5R0cHArfKojNMaQ8Sl/5zkoXwN0uiCTl+JZpGP
ITU/1oGbs7YWmrfc6H5R1qUrjbG6LRSyQ5WROIWTNe/QNpjTxCAlBL5lNmZ5G8XK
T2MvkG9qeLIsVpSdDa/Cn9cuzF1j8IDSH0e/8FcjoXKKxkeyl9itCftnfOwjlSgY
DaJAh3abhvz30q6Sa3qjE0lM2FWDwpU+XiOScAs/mJq9g619YZUweyjjn83Lp8QD
/JjeuJAnIyQSHLqxEqcm2AbDxGMi6UVsxUG0knTWaXKoAwSwbvPDvW4iWav0Lf7F
H6+Dnl6yE9ghuOon4Vk8JWLOjUyWBOUSU9fLGjbrmSWNQaOQJomoEpIKSUwO/jSs
tqZzOu2LdQfXaAO+Ee8Png9v3vg0zh2zzSHzbVY+S+pXu8GVngFzntoTKNEijVY7
Ov4+nuFWCS5KBZMq2g6MWjmvRlaqxDLw18fdOtpMc0JR1nBxZefpsqc1IVTdRejX
NRx7eNd7/3Ec19kThNcQ5ZXb0mDVV0p0GBN9j8KMuIpX8H7+fT8VolNPlzRndzJS
Rj0n6C4RNlj+kk7ZZghFeV1KSvFo2wVgIK0s2FCe1qgmQvTccsWUztCqxKzX2ccf
a94Xei4z46FwunNarMNYpsyR/zc3Q+HAEf7T421TH0IOZssdZQmel6iXac36D3+b
qJPTDy3M2GodvPmGuGQQE7w4PlGL3n+yiMriWGyHNg0Yc5PwDoOO2Q1ZO8m4ZOW1
gc6fIQ+O8QldAqfHxM2V0xE3Tve0Y2ZCMDAaL4KDRkKfn+2nQxiLx7YiTeM+bDrV
zGy6Dn04V7MJnkfi5cwvV3sJBWhzbssXnYu8xESORlnFehx1vSKgHGXLB8mGwPOf
eVWk1xt/mMeD0G/pkBJ57BZIMoD5Q24ApQ58Yr6WZYGen7KcBoBGwFbo7Uq9XEn9
9rhQFSYE0My7O4Ux4Aew1uu/eaH/V6ltOirBEaKIXeQ5Eq2OGc5e+FdTUquM37e4
uFdVqwpdtoq0rvVtGPuOOSPx0fCDayKfrrDupVEJoaxpp++udTWJam6F/z26aFsm
w+FHWSzJ/LhBHWhM4N68/tU0mAsKgU/k2sy7y8bSh3oMisrdX4dhFhyEiNXa8DAL
/uKyorPbJRsnrNpG3T7eMnaEf0mvsuaaArRaAQ33OzXwVzfyfnKw6vV9tnjeZXIu
CLTPZpFo9511zlMahNzmtZJsntZnAZ69Ytnadf781wQQ+8D9OtFmucMcb5I7KJLK
hPJCt+qWLo52XxAXrysFvnXditKN0vDdpHWSO/9sPKdZUiCDkX/twNUbfdhRMJUV
5eMscjqiJdaJZ5d850Mc5wBE1SDF3AjTQZTHaOYszz3DWUfcERgmIuQrtUWKZUjB
714Lkm3yEacd7I9BeM/D2u8HNL7Mv3i8/HPUWpr4a4aXxL08K7Tgj9pAsn9HHh5o
BZlN8NHMtE3t7nABYwgg8/sJumDPDlx8etJkh6FvRxmsyxAqfCBAb4UR7qqMsPky
TFgB864SG9vSFoDHVEeUCGbSM5PPljlC/HzBsU5a7+T+78ymVHtLrTvk5qVZIN6Z
VhwPc+mbvmu8AQ/Qp7mZD0GNP1USetmsoXRi2di5f+1OMvEph1q9/MFN1+P0Tgah
pjWRjb5BG8qEXU1XG7tzoIb/1hxm+3zWI1zq7jvVNDeezf51dqBvD9ZdvQqRJiZR
XuMhIEZQSvoz8stRr5eYvRxQN6D5uW9y0gF3gb5uhzsIOL5zrqKpJkTZ4W3c3BXJ
k2FPZLPhDG0GAjq7zc9HiY9cA0lvJHjB/DdFCvbiH6kKrL+IJZOdmR10/RT1Sons
3xLG38OLI3xDBjhWVWZmU7FF4UomCBRWRr7FnV7I0ZvpceVxeRitbgrg9rDK5/68
ZOW79KMwt/tH2tqlNBfZGseWPdUdxd4NoMMtZVg81O6u5Bj1Q9nqVQB1nkdGtW7z
OFlT5BLdoWHSYwZQwUt7eC4Z5dIrns2hpR79bvwBOQrWCgqUOwTuOwiBs2WpmPd4
qXV2fi2H7/yjLHhTmBA0DuYElndWP1Az8mR6+Kbyy90DzhTjqcMjBru+XqMhHDh6
HkRKii36yS0nyAPR7c8Ku5mCo0FMqTJDKn8LbFre1r6NBmlK3UW6TDieJzByHBwD
a983ZeyoEODXt05TRCocdkllYlYOdX0FMwASGIPGbtpvJBfPL75DPsyoFGyhDGky
2/LZ67uHjFZFTkPnQlWRYcA+7JSoeh8yo9fB1qMvoezTtA0S1X/zaw9vhHaiwKYe
T9l/BGIfbBY5an34LZU88aOjRO0u+oMfMy0uXRQ+IgNbLFRqvapIuywZuqlMD6/W
ie5W4R30vcL/KGNNwjo3t7Sud4nTxwhZHgdf97TjCc1auOnSBzu3BAaP0jtYm40g
QCzTErMP/b3vwOTpNi7w+t1XWGGe/SsQrPbfzVc35aW/tZbrXU15ummgUQ6aSqpO
slTG83nXX6Kw+ViYgvu2Ien4IarDTKtmUwtomyrp/GryCqgnpIpOJNAMJ6S8XZ19
5GT3VPxMT+MQyt9iIEBBGoqRbeBKxkqpeNGr1f7hg5B3KqFexh0c6ZI1yRDt7/qm
TUJMPn2l0Q59zT9ygj0K41fgFFYzjY/M3Ay9R32gIF/LbQs0fogdO0mVnE3wRR1d
g8Nh4cqWoN9uG9DEMVm0EmiVVA/vh26GIbVzO3slYilP+6zsFGezyjEFK7qGSTDI
SR9/2lA+Nh9jn4/4s04xBZPyETTEun/9hRRvLuReascWr/wGEdLAwLlCHqiOG8PJ
L+WQ4zZOjNm5YKIU6YIEG2NjBpnKhZQzRhqidsTuY8N1Su5+Caw80GKvcancG5Gk
qbCH+9LWx8G76XjtXD+R0Ex3kNF7kDoR9HF1d+CSr9AZ0A5noFYBnpESJ6EoV4Mk
Ef7P2KgjkLE/69gHthVT3xbfUHppWx86/UJ5Vy9wWOiPw6wGif87AW8720OCA+Xb
kq3Y0TbKAUE57uhvLZcaduF6oej6Ga6w6pWhenopCaiCMCJzryNaq9iN0opHhbaK
qrMss/acm/wWdUT9dYQBK4MyAKXxpm5A8EtmhX1Fjx9GM5VUlkFOpLCpqArCoDRt
je6pmCV+Ywzjcfwf88cEbp7Pq1klpf1jchSWYVu/2BXJluQ2LZ4XqOnl025V/5oJ
NX4AeOUR5gnfwaMZEkzhe/rzJOI0lF4j7CKTuzosrFuKQVm8GLNJLdiFDDwGZcVU
nfruGqQdG5OBXTg8eVMiBq0LqK1GFC1efhWdlhhl79fzN9mUujqS8PFfXKbjp7kC
aVqjdH48p5gP1iPBAJWtUFO64qvreTIMSqltiCCiqcnvLDh1SfaMn0uXAdTkK6hJ
btheePDIGkDc3oitzxvi+nmQbouLldVLMCu8xjDfJh7Rb2FW7Pa/radxnYixU8fQ
g/bJlIQTPTY1q64IjdokzUrWP3MEpkc3nZyE7rttoRiI3MwVOzdNDEjK4RQxWxbk
IDqQE10ohpb8wypJWdcB7d5M8T9Kn/GAj3AwyOP5qfkgEJdPmohkggy2b2rk/4Cq
UM4K4kzs0+XLHZaX7FmsJbp2zW7r02i7BKp1innypgsYwLjdkPRY5x8yH88+1Inp
o9JKSXamuUcvHqngsk8JnLM8lEoBejJCXX2y/TcI4vYkC2lGRh0Fb8W4ccoEZnGV
8pTqp873nHLGRd/3qO6yyHgn6kQowfeK+ULlOFcxjOCKOH1GyjENpc+SJIBDxVUs
G96s6JT1CNXxZYhgJXy+KRm8ejyOLUoo6HcMk0SwWP+Umv/JmMqYgoZYGuFd1nbs
+VZA12fSuHS2P8beBMa7I9UHCItCI2X3BjtVl72sQ/4dDvr9wvUhzEYCjZpUWdTE
7mwEUHVvcFLOjO+ZgEQucb0hbMO15rHC+gwbjrCkY9wWY5ZPwHBYgKdPRuiXZZ8V
TpltXNTc8EGexaM6B0U3Nruz7e4r61RX9zt9+pM7Bq6wzDz8OqjNiR5iEvueUJZW
7/mAEDByFZ0VW+9PyPhGZ4gC7beP3F9FlIbfYzNEdiXcdlI5Eha9isHMW7U5tyz9
2dpe5/05+Ui1S8kkCywR08q8vVQ2P3nZNt93oY2OtRSmn4S503vmd6iIPkfdo5VL
f4TNIZMv/pT0RxxiKHxL6VSPRINsOapJKF1fBCLfpcV60pdTMAPvQLwtGNLCP6Zk
MJsWZSXJI7QMF9/kgiCVzTp/gp1j+xXvpA7vWWy7OFN8j0J0ByxrbXdeYmgOtjAE
+oTuz16fTn/D1jwW8SBnUUvn3BxzICW3zxatL1HwSRlR95ECVBukArIKpaxqEdXi
PykPcoJfFwxYaIsSfPjAbeXJywDZZwUOx0jpPsOEChcB3+C+1cyRFHHn9FBXyC+c
WQbO0xu9WcjK122X0SxqhWQipZcm0vUV7Cs7R6BgKfxR9MxQt8QOi9VhPSl95D9H
Z8DiURv+AIorgVzE4k0PM3os+kpSg/fI8b2xobvPd5snElC8itX2gFDb5sRve20B
xZf41smyxHGsb1ZdDfzOSoY/2MsT9TRueOBY5kqsuIrjH6gB4jJy4LgOnsR2Uwqj
hiU42tA44zoA68vDG2HA1Pt6cQww2IsbwdObZRYVONYnNbNXUE+sLbRb+sFddu9b
RsDFw+2vMpoXDEsCp8CaGP/xzFDWI2qKiGKJwt2jx5f9PjEDnF+dFuDeau8ci5yK
6jvSsWMOICCTUs0eSFRy8WggB8EZ/gKbQwssEI8Y91RmKAQnedcsiNSSMonOG6/5
K7LlVBDRuHvBXCDeYlKgjQou4KkjWPeS8dds5CCoyS6nAEwuQy4kR6JJfK3v7oBA
N2ue6IObrK6QSZtPJgNsm+G2A5b6eWP0YHNgqADQ/xSitkLZMo5pLfHQeOVo4p4A
6xYwmaZYZcj6ZD/D0uEhVq8nJV/Hl9EOpD8+6yQtvB9A5T67dj6bBNljnF91FVaO
LSURGkSYVIN+1fe0t2ou8Mqw7IQa3WcHMgNsPL9j7WF0NKlsPcq0ipaS6AHM3bnj
5f1ARH3GgY+2oB1gM6nIbZnD7C5XRcK5SOM05mNidWYUynd7yvKIvFxXzsjmP0mk
bGBLhefFNDe0AskHHj+OyjlNJfhFDnGRmeUi9emXe6x9R4aL2R5Z82gKKAykbAyz
F9oDPqMGsQ0bbLISQjvwS7GR0t1ksuZ88hpavaFGlRyz7YHZ5Vb9hn3zW48uW5/M
2bvXE8ovSBZFUnUKmTZhQaipzNv8MsEEUczzs2HbpxSlLilfvzWyuV9qk2TLjGek
5ZdY0xXOlh8zaG16qbzPUdvASxTakz2Ecp3Z4DLATN3ZULdzezOUT7xFsIq/I/qQ
mIwVk7+p+52MdQiwIiVICj31z2UYaf03BIZEaSzIMC+GMYfNyI/84nff8y0NPXFY
P4DkU68QCYohnwE8LXS/LcO626GXU8QKAnf6QtifHC9Bpfbl4AGTXTKdDNgXIYqa
5Hs97HV0wuNhdW5vhoRmQfH7fFfUM5P9FzVGjXGxSKN6aA0IEtSM3FzQGNC3udVq
4q51GXgI5cQNoh2PsnPExK931AizT8WnNLGipzL78NKDiszZFKoiAXQ1DzWP2/EL
YY9GdTY1CRRRmocBkIuk7ZkqxFc/DybYjBZJQ2+qLpgE3sY4uoXes9yBuM5r12f6
zS3n9cdBq5h1rvqpB3qh9vpVetRLPWFwsxIi4U53uFDPY5HUDT2tjo4z1AVtgt57
abOdmtXUJ3ShLv5W7+YvuEH85e7rjJOKBIa5LGKTHnaaoAC/doToea1pOMkhAXxw
950jx8+jN6Ywsbxtuxg8AC+YkA88LkSpDW5OlfgTOhFzb/zSf/1W+VcoH94SEzoO
537hT82nJfhiKG0VeHhC/lWgPoClgxN4vAwOYf8W0jk/jRW08Et/B7oBbo2pHU1c
/zVcKHtBaDlhYxpqi8oDAznSlgOIDgF/wAKTSaC6r8IOZr5guAtG0O4/PaMgQBUr
h30YIv6U/7DHYkkuI2QfNvxgBp8mpMIyaKKaLmtG7q/q9gxpXMGHGWUiEpAq53z1
045urb8DMCg0Pm8PfU4IQTfda0M7hcYdeCeDRJZEIB79zjtacaUzxyU8HLO5C63x
gTv2SYIazn+u7e9AeC1N8Lg0RiJRjx8A5+vwS3dm/npuqZAHs3mK3lme2qpYa9Tg
+oEEeSxDHkyq7QmHKx0QkUAQ1AuJNL0vZLVAhKth49esfJKeMNEYqSSR6Cz5u+wm
j2Vqv6I7ixGIUJ0C5Mc64fnbEpWx5jEMpEFIe6y2/e/kjGkDZM2FDzEuBU+9f7DH
MuBqYIgfJkC4h5i3edOELcK1bVwl7EgNCHGYzysvxI/ICn3cdiLA2AbqgWSjBtcM
8N/bmGHqr4Mkj+hNUCmbRVJOHRzMUOBfDRBPrYxoGWwYI2917bPlR/t7oP8pzuDC
SKDhWjSs6Mje3tu/BBNmQSLBH2I5T570it6dJf+PwxNHbThPVZWqayfusg5rsOrp
1rzDuVz7U+qT6jgwrPnXpHXLMlGAQCq88uEdbvq7tlRYHKH1DJhj8/scjHxWj6ng
TfquGMH+wsSCol5gBLMPxnXD89vI9kFjUVXoVyc1B4MjKXPbdsvu6vloV0DCn8zN
duP0PglOx2OGjHxF8MSrSSKNiZTwhvjn4aAuhccuJUjCH5PZMCUePz5tvwNkLFRw
3/IZ2f8XmMZB3GAvDC9Bq0znbTsDeGulD5d4qUIXiBycg0GxyUqUCWRHLcQLJhgp
RlRViJVqIj7eXT/fsOK19akM2cQ3WLoNo8SjaHZGYq7Lw6/+937HG23nEEF2CNjX
561zlj2oFCTi1AeYLTTCfmx7nMWiToC1Y4LfoVTQV77veUTiz3DW/gyFhaSPqMcl
BDtiJZ28s8QG15W0tcCda8djxnAarOJfRUv9MKH8Dr2PIS+kMzyNu1+hER7SnfQm
uMOjBeIr40gHJDCUsHOufGfdcbX+/oOaAquatp7Kcb6MciId7mhfjchh4xAPgDqd
RkPm9aKHJG4lnfiV6WFUQ3NChujxkCEV2xlgvWzPIFy1iLTnGO8ifbs1rHQr9X57
wvD1CVfStIkvf4sNI2gVLxmGpsQpVGaxfzIoi1kEPD0KK6RtbF8FExAfQ3x4ntVB
7ES1oQ3p0LXY71iz2R2WtX2r+kuvZ0biREiv8I3a5648gShn2Y6qmtu0Tc7MMvFF
3VSv530RWBVNkVbk/YL/vNIAY6oZogScT/N3nEp5APf6fMz7squzOv6TZKcaXv4J
bPxF1v0rzTABVYn+tnnp+9F4d2hp/zCEjTTegsNbnxlQrQSx66XJrfJdze9i7HP2
ELO57kADTd6eZQpb5JLSlmjo9Mg6YHKepBdAEoH7uqhmiGn2C2RYMiNRRDIMeQCy
PV+foX6UviMylZi8SeautopK/9mDUnJKbUHdNauXYdYCiA2EAzBpBmxxvA5DRz8c
ikidBolnDX2wMAlDXAaCKJWzb0D+IphPfyo8rLBdLtXgVE9BAIl938xKwha4BVbM
pM7cMqxYFjqS5i33b1MIc/fah1keJ3dUDXubj8nFIb3SrwTlUWdUZsKBHARdVA1J
q1MUOnUWQyw8eF7q11Tug0w2Rgy2FCL1Z3wQzKnsvIo8z7CUUmhFGNWrfi17yUEN
iM85xusiXKvqrMEFcK3wl6o5Xm4SEFDgJssKfTYNg4kymSrfPFPKsR1vZZGrhKeM
pKpdQ909L+8wGHc9Q8mVmdS0I/15LyMDuILb/cnbTf3NnPiK4GXiF1NTpc261d7W
3RAHnQqPbXL7rusYn9u509GAMG3RKt7n8EV+c5iwK6a0lJzDccC7kYHJKSYTNy8V
H7Zo8rgiP9DLiAUL2s1gQAz/LyZnuMrGUCiW0HqlD67sJlNECHTaLd08zBqo7saO
GcvkFoTkQg+RAsxhoPJ+94+1gGT4qIZyNxy95N/uH/Yt4ZMmWqZ/ffRa+i1T5aTZ
kH7MpNXuPm0xa/OEmmylHo77GxPG5OiD4Q9691aFa8GnCL1iClfMCZM/Yq/vV240
+v/DHqjOzWrejIqp+jpkN/iR5elu6EG3O0lMkm8JQNAqRVanRxjvvRJJ+999VIgU
LEGmY2XrmjbkTGUuBwuvIj1IscBCm2271/TZjDR+970v/ym/25/LUVT9DtusVm7+
n1Zq/nkEtd1Viv9GXnU4I9V+v+zn2Jxl0dVdhSd377CIXqqusgIZO2cOhUoiarBf
ikTxequbJ5+oGBxCx7zxNdGwTsawlLyb9tEsi1joN27FhZll8YtH8qTdkJVItPhZ
MqvvjmqZRWvK4pPzA8n6QCRyO4sQdlEh1eufc2sn/U0UKFekdvzLz9Cre+Ls6jTH
346/K8HUT1yFHoXcGHfvXnkcRlucWai7gqqePsVNenaoHWJGmHTR3T651FcoI6Hf
SnCQNhsnsBKEmKF3gMzk6P7Ce7PilSrKFvHouvF440MlimeRTusVnWCaP7lfqiRb
WLcF7CdcZE44KgZqV/E25p9VHM7DlCAIbgy31F3I7SmeMvrW3NzOTItu8M2gCbtr
XIlKvVpD35MYifuF8OC0DIyegsSLK5jROtqepkzzsWi5kqOLK6w5wnVI6nddJFy5
+Iy3BsPJg3G7Wx/g1kblrFnSq2ux4IPPWG5saPx3J1DcbNPH0Krr9HIhJuWXD2FG
WfCJC0C2EcHgb2OsGiAqrAos9Y4x1wFuFHk6gdoorLfzQW5ujJd1AsOUf4SejRZI
UcFDxnQzbW+Fnn21JTqgsDzcuyDmIQ5kJGnzftmK25XCrxtkMGwqqGXNns6cFdxC
xPZgxbL5EMGcz4FclxeuTVfXhMbGgHF+UCobs4S/anspzJ8Axeado9SB4G/gZecV
rCkceht18AKZR62t+cHAIZ84vTeJn9zIHXF7AuHBeuPPJqM+MmV7aD1Mhmxj/ug+
Wi6cy0MINBtQarJHbGYLzl6ih8V/p3UiwiGFyuBQlErmRNC7i2NdSJi0130Zri0Y
k9kuAlJDlfrDwz19GzM6GCPYIJ7eyibx1fVB+01S0V9l4JfX9Mndgy7T88r54MtH
exr4Rv9r22hkvL7+gjNVme4mjE8BSFTk+jvcMgysWr+pXezWq+e+jWgQvLVo/m/e
wOdbILJ4aHQ/+SNNKQa4VzOz3S4F+X2TXomREg3HpZMrymOYxTPKuCTeqs7BlHVt
QGNQjSx9MajSwY4lMasFS9PEPZyMWDGAQ89Hv81FznyE4ve7Ok5yAjcv7cz+ErZm
VHPoeMTV4qIuAzAzqLCyx/uPCY4mW1UvPd8Wb+GotLV4y5Ynu6vGBmhjwz4dGKGN
GA77WyiQPC0PySpPEg0T8u5pW2ML1XK+U+MCMCq8sAAxXPlctjMcG0q8LzMRLG3f
yXC2yC44u4RNj96vhNRgnmQnU2LnIyFJLDe3ueUaBJMqhAV98Kh0oNs6gzV3Cw5e
1wNlBx1A1IRBgrqFvvowj2ye/ZsGBcQLzdhByOxxjDqlr+U1tinqMyKexNn81Sic
F7+4RaGu9VQLWNAeOJVYhO0LJfmS2kbnTTLmEw+CZAL7+jHrZhwpeqLWDoQN/Dva
j2EmnEa8Mog9EToJ952pV8rZ0wnqdhXLSa4EHDlQgjaB0HoeykfVeO9ZpCHnVtXE
zkefmyhH86f5KOZ0ZBolCdQdufxeBur222la+5374Ia2J43JONxSKfTjFpwxrMS/
BYjlCW52yIATI2vsHcH0ba5y7gPUmYcwpZXoYl4j7x2NFcalCJ8Lzjlzwn8pkKET
7ojvy/vwXQUC4G42ZQzGU9S4brAiJNgXd4IS0IvZqMAUz8NwehZb6RoL/unRo4aM
8FfCce7lmdsQc6qLYstoOpN5Wwm/CxcVmwf3v6WtwgMHkYDztW4tSRchzZxku3IB
Oh/mfnMjOOl0TbGh4zsX7UNQ1xjl6S/lWzetj/D3r3SCBo/b64ABkRJwT0J7qiXL
HwdGuX4OwXNE5xb+Mp1O4QIlBeoHIlsbCFiZEtkgPth7lejjPvbnwWsRhD89avK/
pSBWb6BIqTq05gW/1/vgmFu3GFaU7Ig3mlyV6DeMN8v7wuGJU2rrpOmb84wReHom
yRBo3yMPS8ybWQ5BdqXLc+eHsZYu9Bu0oAm8IUYVinZfstrhHLXJpefhKdcCaH3I
bO0dvJqh09Ad4wEshqDZjHjqHUj41lkpn1kiJLD8e1gNI5UXH5Tba8T2dMnAMP5d
LpI53Je2q/cf+YZmYGXZpO21flftrZx7j2bXJzOpV1x/nFeuwzfn1jNGlzvY0nIO
x2cJkZv4pujFT6XBENaIvY70b+7UVp5DHDMnMc5/kbhk0SspbSqA00t3/e01JsWG
NLXosRXod88xkYeggj+dXqS4nH5IN54DiEIND6OyDGjXI6lDzQdEw9Au66gWGxmI
98LhPCUtpOkXQuhDYjk0KnilRAUNeqhuWE7VRCgOVpcTwaiQ6yClUPtoka6pTumj
ciPXHC1sroe6CNE2QpR0iEo2Xch3V7kflRxdwGcBpEy6lSJJIH5Wt5DcGqOoxiiL
WJMcbJlabjeSSLdHK1vdEaJnn/rVDfNBuQvsFoZCU9MO60ZQlIOu9lh5eZm9oEtP
do+ZFYET9/+DvHuRFp7Km8YdRqouiJOJb5jXLd9MgLuDa8YAZuemCM0jtMr92Wte
SG+E3MeNK7K6VyEaCV5h1AFVIULGblz3TPtHOYO942wCd/dykPCWCu6RNbme6fy/
ffXH5tv2iZQTSLmrlMxQ19wp+gL8IyFy1jil6GkYgKUn/VPlYbDHI1OAQHocTVNJ
X29+M6rw5FrFI4dsvJXDhDOsooU8yVC+d9IcJzXQYgoEfOUXZjeCl2j5vrVB9X4N
CF2jR5iqJscgJ2wofFSSO02a0s0tlsd7KGfIy8FGw48GYZBupxm2hYPLKfBKuvuL
ux/A1fRJevVTbLEx/loewJcdirkFs1TwkM/VMV3teea6UIWROjmWvkAVGJgoQQ8z
3biu3l5Bjl7zjOpIy/TPbYDIJRdfOqnkP/xWrkb7Dq8GQCluuf2wg1UqSYZLlEIH
PZq41/omtS2nE3IAFnpCLEMvknrx4/ovKTb8DE1VTRcxRlXFkzpXyGZ9IE2X8nKB
ookvSFN6ReoN0rygnLglTO/p2H6TjPlsULvNXY4bUyFbTjydGrq+4++MGJ8nW+Dv
KTY3KuEKKrn5/DMuSLZhXmq4ZQYJVwyKE6qx/EQmftZyHA8zXpSPCmbSH6qR/Ebh
01wU+xkHJ1NKyKb0xb0wjCzS1qEVEtUL0Egn359QLULRnWBzxwTzJ196W+bzv4UU
te8Dwu218/o/SDqNZhwl9W5XACSnw23UobC3+IFlNprX0QbcLeO+hEW1Da1wwktI
VBPSvi8cN1XXCcwn7cXfJvuhvm9ed0EXU20rGVrfLMzxr7pSQA2xfNHuCTv2eMdc
t0I4BcfyZdNH0BXDN3qN3nz+myNwWB/LBuWAbdObg6Gv3J7PJxvmGsuTEjPOIFBt
VwxTton4wvlv3jMoSYVTwn3Hy9QOZh1/V17WjTcAGTaN4lPZMbeIEaUL/6xZW/49
f2s8EnDkiIMVncxa5CKOIGc/WDHVmBGbBzyI8I2eeB5F6yGUOeXgjmSQ5uN58i8o
Qvv8BYj6rBvNYNYPLfaGgqfW91ZtHcgtoROCOkEHCFysIwduPV8xsbMXYL/oGZwn
TjdB+Vx6f3w/tnDrOLSg9eKzD74n6yP55+zq23EpgXGgjcK1f1rEVtzYBObsT5sA
oIZTpXvXG9Tnw32IEk4brvjIKCMJsS/wllGCWq+W7ZAsRTRLDoxWZqo+6StzBLjo
3G0lOiXjDi7OE/rSxCqCOzpqEs9nULtNEisbcTQWawib5M1+BHm1ZkMNzkrBCba+
bQd5VAPB0oARL10LMn9afdWN94yVA/BhjO0OTk/FsfBifbJxdzEGhqCR5Q67em9o
WUUqcX1OQvnK/uMD/7mEsJEirXR51l5wS/oi4CiwWfZLmINl7qnBluaif9gEG1yI
xiZZENIj1MH1jRx6GIWVLaVDvRx3z1wsGzQ4NuwU2ltfNQepVdW2rHxwhVBdVAqT
TJr62UZq4yAlNksGYe0HoQ6UO7Yju8aGHOPIb5qd/SzYhcrPrimsYVpNmYMdnpp8
PDCqZOn2J0peUCVSrANS9rOZU+EG0JWAQqvUp7ZNMrKiLzu2Kk5LNmqjVMJdz9om
PaAkq5YxFY02HSkZ38bzFbW3R9iIGYRlWNotHzKT4ip9qYmAMELMV6Od19yQc7rF
ygzzOrH+kJ3mSYxlrQM+0VePOxkIV6SIFFpveUgsc0BNMJ71xERqHoE5eL5ptP4t
xp6E7oK1CTCyc1u2i87WV7IzE0U+dDSmP/ZQwAiS5oaf1qJUyBBJBAOaox/Fe9AB
epl8wiC5P35Cz/aIGnJ1+AgzuUdsRY54JLhu3J9YOW15jXdTJF8h86ozYPlLLBus
qkgBFR2qCV/2zneO8JIW0JqArfYZZ0VZxzfFpnYCiLAGiv6XPrj4s0395MNx20nr
6CHSNp3fNGM93+3f9OgEsBpppa6Ve5gLl8s+AbEoXF24y+JvbrtseYZqMI7uFIFk
LD/n4x3Ln8+gE/tSdslgONcSI0AK/+vDHEDuUuDTApsBv/o9fjlKjYrMBJndMaHc
HShVR97Z9kmuvAS1I7fTBsnsnBSNaIR8+rYKy1NvqIroh74QGGVuQ73WObC07KQ9
jcKvPUQ3BpAXekIA1V/+EvmqkbZ6YOy2i4oP4Zgtm4AzgBmAK7nTvz1eG3JlvmCY
FJVuPguHkiuVwSqL2MNLCYaFDtqMqV5cCQUopSBBSnsiz1KkEnTRGYS9G1KotTGR
JhVjh1me6PevwB2OI3wC1UQoRlgylPowpXH5rGaorYfD7HjCPlgaP1lnNGcfZbMr
P/0bOBM0tUpmnUdCCayfiBuBFSq7Adq0BsuXjIEa8VcJm4MH7n750/jawcMhh+EW
4naSpn7DWn1Q4bQLvB+8+G7D0d3Nf3/CVT15t3/SEZmTkH2K7tj+FoKpUtcmfw1e
lT1UFb6U1V2zO2ViQkbP5D8H6bQprzwTOmcQXKN0KR1F56yD3bpv9pRldg6FWhF9
7sCt6HqsSHxVzkQNu1Gezwy16nzM7ZmsbbTltD+DEpiavBN/AEUvDHNQy7w3gJP1
ObdkU7PVvynWsrQwoKjqj54KqE9Gw1Z9T1jnEOJMz/vRN0zZo+ajkPRKrNZ1D5t4
IFl4HdqTPERuUIBdJwJTwqnsNsv7TDu8QNLXH358+B9B8mgd5i+ApSAxf1rAjzhD
Q+v9Aiq2BCT5hqdu4sevUgoYGAZbPq4uib3MWupPnyaWsd+vvFTK8xCTbyCaL37I
i4ADM7hsywUQOPYZWQzKxyPmNIE17Pz+APpRSuqPiI4XcmLXDgKxn7ur/mog7fpg
rlTx2d/AErc93I1Pan3o8NeNSyoO+X/7jI6BImc1WZnXgOCvCMRHre94zq5RCH+X
cPaeyQrhwPFwJEsn6z0hPWuIM54503Vw6fYbDvU8NYpBn721mw5TxhCRHLAUque1
LVdw+hihpEhKEj80FbszrUhPQ7wXkd+2QU70d7+RKBrQc1Sju3ROBGEUHyb5x8TB
gmXWmEsI8hLoqqGt+16BX7F1trV+fANwzLllV/DU1tbA55rOdRNTruFleQX9alIv
dpDtYYLvY23D7V8PPz1f4IVyq7OxXAkWtIM6QRyVY/1z7wgzZvnVjQEGI6/ArPqK
Tw26jesC2lJEhrxFpdKL0RBgZlZkaLYKLZusViSuZVsXbCPZd5/hBjnZxWyikjHJ
N6Bl1+h+zRoFSBcScY/1oJvpN4QjRFIaqW2xXly/t7KoRL/HvSa4NqwnqXtxWn/W
G1f3MdlJCcg0Fjgr0D+6clTzzI5AkcGHwaheabb/O6tdsgLAM1eq/OrKCUPfr2vR
tcjKTkCDfdmSnj8rd8zoKOE3fmh7On6kqFBSXoGY+YgkIA2PCRSi4blDV2YXfZwG
m6/gcQ1jy0+eEyzYNjdKVyIWgk+2KQj+fF6M+fKj2xNn+sjc7XatRVkLzwreIfQd
HCGsNeI+SViM/JLJb+ZrfKG2Cs5n+rA1zmMWEwt/Tky4MOkm0JfV0c2oESQ9X4cO
nqDHrNc/4+Txhl5q47tCV32sIlRaJWNg1RV7uZzlUqwLlOqmveT+SgZMrcYkD0jF
WWHlQfOg0EYL874rkSBBl6VqoqBn5/bVUKzsAAtNvdyHKgkqZxF7jVUSYv0sA4l5
bNmnUcocEYltZkpuiEtS/hNW65mTX07dFcq9rzGTm5BpVH7hdY8OTZCTsdEs89uH
I6biYwb6VcI22lEmMuNqY7ipOrgXh91jX5YqtgKK+AcW5u3DFGh6+LRdoOQBUX2h
Ioa4+/zyrno09gXyixbCfnQn4nBbmNApfNExJVFgMqU0yBNPWLhWwoSPQl4PIbyh
2NfBRxibOwerxqFMe/QbyzwvkfIAUbSYeAUH6dFGwMRS9Cgb6/9zLUSMFxckeLwT
w1E4q91zEl1/JzVjaO63GaUdpzrNiBB4I11dyxOp+2j36YOKRUqp285q7sDyj40D
Jw4w5lrDDC4+OWaQYhjz1kq60hb7zIFCFsh+Dvi1xVE7gg7XtOFXKexFDYZuFt95
LJ24IV7+N/vwJftSlWwFkpm686/fj6E7NBuyWWlfASLwBmm3OOXeHHwDiFlT93+m
hHkZkf1+pWK44XGQcZMNDL/V/Hn95t2nseTFx+70+Xs27edEHClpafCCbliUjObi
OWSGSzA3odWhQ/S7nySstceufs06+K4NI64/8LK0U8/NoBh6NYDLn6RBQxwYPnqW
YJ8JljEMfUxp4Hqry6vmYgu7x2LWGhQn5xS7VOlbzhbP0heEl5mzEIoQ4wWiAUk8
woRnDYY32UYLC9kURJz5zNaBX6j3SBUwz0vUjbBEWk+N7pisPnQa/6Ia318Lx1ov
JftZTOHfU9obVGcur4x2iREtfaMHQSQuXvSuC6XFbJU/SkGk3ldkNMmac649xkMI
vn4DDvCNaXK5/ckkSSASYwR33FzsLh7DJGt1kVZpaU1/r5l2C+4Hv83zt52Y5mm1
WNEia7T2qpLX+LUZBvVLlPYlNo+/XZblduHposX3MqeE5PDT22QE5LOqB05XMcVL
LrgfSdVHHiZ3hyzpHiHzliXNyByCJDA3c+Ro+QI89EH94umzVGm/bGLcNUYW+L0E
M2RsMUovnnEMPjm/TjuGXmT+apLLL84DF6N2Q8cd5TVVxttBI6uas7VT7S+CjBYX
WmMyoTnXXQQNN2GcEbWCk4nhZR9uDXLQ3TTmwJSf1fVs3a74bN+aAM1aKsFS4+VR
Oe1aWCe/k7W6VfA6hhTRqe61aaGR6TyymRI59sO9RVIhY4TPJOGxizVZWWy0GYf8
3VsjFZpNlW2UTnTGGFHKAvIDTDxmg3BJhBdy+Mo1ZkwemtGDiq7q/vt6DyMWT8zS
Gz0ZsvrD+fUIi5kvzp+2fTEB275J6bqa4fcw6xubJqLCDGrbVh2YaFeey4s5OOGB
ermMzXK62K/6YyT3S+2tNFaQQXLxySnUgqhKBR8YS9MPm/hmSZdfEc2VeUJgBjcC
sqGWR5B72kn/PBTUhluE719f4+WMdHyctXS84+j9QmOVAStZpK5EVLiM5gXNLtAL
Z/TiXthUW9JCbBTxrOp7jTWKXWEOqDm+VJzzGBFZnKuftPBN+b6fvmUTtBkSguio
ICShyRyFigXAkTdwAHI8aNBDm2jhFOrZedtzi6jGujuvJPCczadPak9oXzF08O17
ONkiaXF+q9X1Zt247AOoH9T7UU6bVokfT/67wxA6IC9zdQMHo/QV2R1AqpUdVV47
M+WJ2nTsSex5BPAJNuQQQViDb2Eoc6eFbWnG9s8S/czf9w271/p2Bjw4B15ep1AO
NA5/dxc1PFaMrsGpaRTxO5oHA6IQpJ6aptPLN6ymHi3aPCmqRkDrjPG1qvQPvIM+
6vHAGfnb/Ah/4TjAPV4SYaJGxAZLs1TgNNo+TQl/Z+TUnCzXCTYE70l0EtEeH2zz
PRbjfXdwOdEUQbJst6vbpsKI6mKhUsZvOi64Dv/Whj8D2AnTmeWax7jz7W3MKOGf
pFW6TPFjI/y3uWEMO0oi/0wuQN7RKFxsTw3braIaUX/5QmermgPfPsQxoxe33uCJ
Rm2gceHTv3rFfJFwbVNnmwH4JF0yhcBuDdYFh5yLFe/qpb9QJuaNOhzuz5RGVtop
yadMSxd0CjVa/jLItIXcYH7BlT7y6eGblD9PywFWDbUhaZsQqIM9JCuha9VKJTxr
t5lS/MQoCCoVgYHK3G4EEeyEiSFgqZ3oq9UIbJlCipELfYExf/COXTM1Gt+R9pnw
qcGpfE/li7BMmINeOnAto+4j26Wv16daqMn3y3p97aS+wLBQcNzbFQxTKQ1Q3lZr
JPdDkrYcCiRbmYxdzGCS0nzIeKMprUeDB3SynWTxE2Vu8gQa3hN6NBIy8hW1t8aT
rPor7TSsrChtGQqeqdcGyAs+waVwadLk3oeJ8v8jUmtnfdaj9XE19NV3cTksVn9n
E3EJVh/93gWwPfEaQ9X0LxyFjLNvLUVZuWynNqhJMUeXYaZXkMGKZl3lymuQZsGN
9dTfy5Ro/iEN8H0Vspg4IYwxDA7NYXLU/slhzBqVXRkHfDBaKfynxYqoWecvq8zu
dNMchWS496BNeXUGsIhl9BAvsFC4WeXKdIxMbRqKGCvGoVeApiYzRUP6/FkhTNQU
02Qo7kSpAYX2TGHefRSlgkAoo4aqLAU3ff6JMflrMofwQWL0qgUINIJd0O9EZext
gxRUlpmvzb+HCUnAoE685D0ho01Gck6FM8nt6SQoplyjhyckNT5578X29MMTyv5C
xsjeOfSTT8x5+r1A+kE77chJFHnIGKcRsXFYqrF6shGp49ZFTC59RXbryJCTFmf0
8PiJ7Om1qBLoutQzlb2diRagOVYzES9B9Hlpc/USsUap5Ln4LO3L4iEa6+qD3uAU
05mc9LyFYUZoBRNsZ8eZHIMZdnV+/qn0CGpmUqfii08N246WImIH2eBWvDJ1gUNs
LG9+KN7fzipMWTl2T53BdR7MNoisJgMcFbuNptm3if+gA7ObU2i5/JSLDS9pHKyS
iDk4xpDmXBuuzJmV2ZqOtIAP9arSkJs9SlXaNIvOehHgJ59YpG8kx0psR5CA5jl3
NCVw79xu3GOfPTTH+jG05jJcaayRgqUtsYa91buEI3L5EWH4lRt4PTcU8qap61wY
75h2xoksAxxO0KJRzhohOjtgge+LyYvPby+67wJmn1D/ghnYVI4aLeGdJ3W56NRM
0nBa4xzEmVqhwnzTV7vtD1l2VN9DCcFJNk251cYzt258r1xchee9dJKoBq2cQJmG
HqC1Y/AuJK6gQ34YP5ylxRkU/4aJClvwBgQe8s08P8ghC93e1rnUBU1NlKqr+HAd
6ltBt08nLb1QG26PFJEzaKO0Y5sM+TUIY/dDJXuZMNsTVx/zE6PF6pS0VZtpFrjc
nsmArj4Dqb4LHoCgk21h4qLba48SrpV8MHfWNdHelZ5/Sfy4wzd3hkv95S5SJpYm
a5z+pMV+qFNMmPWjsaG3WHYQV31DO/YLYpX1vfHz0Dyyiq8GO+SNF5de3w/MFLAq
OI0WTiKs1P470a8Pm6Va5WRCUvmgpqg0G9UOuDmHV42GPZl7jQLsHP9oIwqQ3OeX
IanSM0tb8TKguHysrfExNOMON2e/2fTDsHPYVoQ52cp8//OqIzYO9OWqq2UyjRxa
8CRe8c7yh6WVWtM8ZN/Hm4eodS4e2eQXWZu6Y1WU6XHa4/mKTUAHw7kslnShb9zA
JMgn2KIRMtTwz6TFEvX5aTY+qFG7BrXUsZJyWpNp3hTWi3D+XRvfeo+dlK6ptodL
yX3Fbof407UJGWClZtPKeVcIl4bDyl062Rq4NAKyvlI7AakY8P2M5vSGRgdRD+al
2yUtGwMn2DCw89bRc8J2PLYQcx3B0g61TA4q7pS98+/8jjxJNwgs+d28PfmlQr++
O75H/o9wI7Ic7/vUrZCLlcMkRNLKvNv1+VsEvLe+H+GPi2cqstqgSPSzu7wi+NKN
CdeBgUdPjAFVt35qqdcDTtg/bDHisHQO8cUrJ0HxicYBomq44NL5wWdF81RkggKi
PjWPxe0oqcYSEB59g4TxnPXENUAN/ZIlh8dPfcDIoNK9iZCppgnX8bQG1Jl5ewxg
6oXohtdVFaBI9Jhq3Ete4XJBp0BT+Q4OirTs2bsK6i5jg6V25BQa+QFNBAReGKoZ
N5QXhkHZCnTd+YkN8J7lbjFy/7UDiOY3+E/DvcbenYFxl2NCxFgSAPltKP4FAgcU
pmK7TUTXn8n2z9duFP2qHnQpxSKOfvbvnq+iEONj3CD0n3W8XcEAzKwQY3kaHwXV
Zon2wk7CVcZQIDvkGLlMucWaQhkWqzyXGgJ9pV360f5jqY3JhK5b8SSotK0C7w76
aVkwvX4roKjwaHtQTpKtjwKLHAiiyzKm9wEBQVsU9ajjOBf2SlnGYVgwLSo3ur2D
BhQxMrujd5Wi1LShZBUyQXVNINkoGoCdvhhp/uf/ca80/PoLyguEhHtMksGeVMxd
6ngPuzPMt4pf/3ySxJNPkbGAk0zLHVyenlWlqwXHqK/dVnZ1TGOtmV4TzOUJ8KM9
Y4KwD77N+jHjMn+6zrSyIMuyIO2OrzHzVWm+cr6QqbfIofcFHK7f9IeboHsP0TOy
gdK3U5hA9lwLBf4S6XC/2BElrjgkDHzGFbapPiFtl96lYwRRIJ2JpqT4aSp2yLRL
gdD1gHriUN96wSwvzTJo5HcYlmHR+Vteto6nSarMavie8BLPK93z2tYdvHndgjKp
NYC/9Lny3BaUUX43bXsAUTrMUD39OYH/dX/+0nC7JnGVjHuRp6clW0/gxnhQX5Te
4uG2c4lasheUZm3ks9F8STZ2RrWY+aLgSLU3G1PL9jZqv07+ub/IipN1qx5k+i+9
vvsSk6c6C2cajcK4keIWf4A6IFGta57cd4shM3uzgrZxGawn5LbA9fzBYFDPZIQQ
zxk/ASzMf1zP9ir0/8nNh7/l7yhFl47/L2FTs2aM0fFVMy6dPVLcfBD7cqomXc7z
iwmsxvaHuJ0zGsdE6dEKIdbl9LYFCn2qcklZp2X87z50dflEfVloAMNPB64yhV1y
fHMvsg1/8Mwg2gohV9cdvH3FHXMFksJAle8es3MTcD2Ns+3O8xsptH1yw7GqVpif
Tv112rpqf0myDOQTIHUJN/ufHOGRlg595waKB6t5yR04geJqTD8Vk+l23DQcLCar
j0P4+6ACOIgEigaEDJmsdPLRuLQTGmmG/DoFs+HMVyLr9jypCQ3nCGcQT8+AOcxm
fW+7lEbROJjwB03gYmUgKVTJO0eMXxsXWcbdpQ3XNzIJL9F364zGZYH9aJ+nubFa
/56vk+KIGsvphXDrz5FZpXJitY8yLyNKcscnMHVjRbFtuq2x5yD2sB7v26dEq3h1
h5I/CVK4KoeGf22QEogdXoCNpP6PEyQtsjeR6RnAcM2doWgBxwBXj92RL/5RNjqg
ZQHViDxrRChqvK0U291Zuf2QFqbJ1oPzjJn+mdCUPOSDUTDIr/884LkuEuGM0Jvv
afZdezwKkICAqh7YltXSMBXwu/vBRFV1yfHRewM6MFxEby98UVTxPQ4BIZzr/DL4
PLEjOStYt7OB6/zFAQ2/MBQPyZhd3JrzoxVbKJbsot0jyAl5fD2DcUz+JMcNMg+c
f2aXJhDvl44bTe2VfunE5bwRojzVFjuaK3boa8sr2oDCnf8ufXNQyiqZLkkNY2Pr
+ZpQkA7kmYL90Lo2dJghLG1b74ouNeE35fMIlXI+n0rqtM1GmNJhrx6OA1jiu2IR
MYjl320sY8a3bIjydML4GpGoJbwIKPJfVppEYVeaKlDEcQIbTzMIuxz5XPSIHVHM
BUUfWivuYZul8PCHhfdDv+2cU4KJcL6hWM65dzNlnZ7dY1yX9KFI8JiWlJqouw3/
NSgM7Xj1T+EM/Mnr7yzklzvG6XcR81b+4n3mTF3UOi/9IIiL/k4I1BkGY7rL3U5D
GHWnsLU8sLER+GRw9N+uAjfVsvWFCqnFWp2lyBrEt+wE7hpnepqi+UOsLS1Lnd3J
bJn4Wzpfkq/+8/exzEIB23DsMtIUwflxnHa6KBdkuyFY5gWsleeZRng55fbni8El
vhhxOL4RRdoUwCn1T53H8xIVA8rrshx0PG0+Cb3Mwz72SRQthrp6Vt48x32DdPf/
Wm3uxAgOwKHjcwYcS75vM0ACk4SQUiwJINs77kAy9ZDSWjuLbHPv32CH1aSIzy0T
gzMo826f3A6ZkJtWs/RWEWCesYGr5N3B5t6udVmExUEdlD+qok8GMbGMPb3MI2U/
CS4mjR5UnzbYUgRobpK/vOC6F70AfmVnsFqwCuJV4FDT++Tmrn+WcFGIdlvbgdmS
XiTdx21HSvAjJ2qtgxjlA7OEyC9CPmeJpQi1mSdTkcXxGoS0f8mSKidteaLSj18H
Sthzgt468p1T2ey1Jzmr6cSTp4MtA/UtbGUSpKX3wQ+ZroYhVyWgCyXxPX6fmOfo
9FW2lHaXQHq3wrwjbDaZDihsI/agCk+prTSCB6cunw5+s8R9NfKpT4I9V0zUfz8I
yVP24kAJmHs50dkMhHlkUruHEbAZ9h8fuAVqe3TKBnkUNriXkg080CSpCLeDfO1d
N6zeKd5RTgYyOVlYAlnvx8YoDrRF01vzQmEfVOBpnXKd8o4VUe+7cJyupZIXYxVh
DSLeR0BxXWJHxsPu53Of6qYh92GRXcXrM4Hy10DAQ38RF/E10MFszkv+6TfkyASX
ComSNf2KyF6WTx71JZVEAKGHsO1iQZ7MF89N9lQyyvdxhkEFyaRTc5y2Egn27umh
0IjVdh9hZcZvt0OzBi9yjtOspRr6lOeMMDfwTxNoRmqpDlYTazc5NeKfDlXyaPYX
5QkXZvkUHk8FEdwt60OvEcaIpTMTUJyv/z3hmOR9oE42VmcLm3EG/v0lAMPYWBTh
wRgNE65tdkmsuKYE/waJcRCzf1VZ7Yd0vMrDKEKqJlXU/cxH1h5f8BSi1QAHiY+B
fyFsy6zFM9zdy5lHyYqFyHl/QpBsr9u+zZodOLa6Cqb/WPDDaT3IqapEcwkMnR0y
fTLz0MHCJeuMKsELmCByRp8wUiPqu3LpipugM+P0viL9l3dtphanZw77G7Go+Zop
9j/J/F6jWg53VLTsH4l5nyLejIL8APzxNc+pY2hVP8rPclDYthB+tbvw/TkzQGxC
ixX8Z8Diz2sewvXGB3xsQrWc32jOuOZO0ILk/2TUH8UW27fAa8JBKGhuF19uWQd4
6z+xFUtRljONEbfxics8ikr8X6HAO93WbQDOwSpvra9hWUO0fwEA9TVqgXsjcydT
ZgflgUXWj/mULS6LCWvARDG+gvznZ6jVlI4pLgjlnWIsr+oFitMNhq/o0yTvjydM
WgGu/DiIwQdQdrAdDQyLsH5zjZ1axVyGCf/SvUkuXhlqRZcNOtZ21Edy9tyrvdVT
FpYMaHTxiH0ibFjYZxlVISj+JR0aMacfCDdpCsHHR9T+CjhC+WsP5AIx8czG77g+
A0etanqwnbH4SDctLL+9reYvi6e4qwyKxK5QdJ/WbuG3CZg9+SlH0nDNg8/Z7FdF
zVM96IehU5leMImCzJwcKR3rXxvN2UxvoXxG+8H4FV0jEPhdNoXEY5pf6haNlLBG
LKVzH9RYL+vVmuXAnkS56yQglbfnTvSkG5sQbo0KEQeZIQcTerctdnbl+hM1T3Qr
XiwyIg6y4g+h3B86X8nkLBUzjAgdGG/N+90FVDVlhW1o/spw1+suuH+hJN0EOsAS
e89JvSK+btKRVC1AXDUg6mb8uDtWNOCZoEsO4Y9IJfD3qDHzSQVyFbFSe26gQWFu
eRjUI9dSktf9OoOPauMQv6A5zpES+vYmCy4RZWG/4Km02tGu5ZXyFRczwLrJ4wBi
jQj3kK4BoYcfBeT30oKLc6n6byobKhaD9qMQm8/nScbY60k1B5l98S6GxkGYPMD+
d5phfES6m1KLbaJiToGszVMMvqCWQyLDD3UGobXvicQp/5fJSgIoDB3T0UxteRcc
eivS5rqewNPVCdNdFmZVWZAsXJRzB7zM88uv0UdBUy/OQrgxKXldFpT+mwJ+jC0c
5fjETy6RPMfjz2NZr0EU0WviB4nExfkShrhNAcG97/NeREq7eGExALwnU9iuQTtV
bYaheQp3atup98g9XPje2XBogePfaK5Y0qunztz2mTGI7XUOicv+kD4z6jt3zPQb
m6v1T3kLhF1wVQZP2TUdXQkie9zba/C6BdG3ldCYKwWWSkLwMLecqcnSnyNfvNiG
6gy0FcHmXZabNzXDUKorlzr/VF5N39lKTxa9CNNBQnjw3jylVuG4TgFvpmwl7ovi
WGeca4fKKR5I2CFl5qotHIB2vG7Uq27Iin1v635Wq2mCP+I8LkNCkvLOaM6WTvRP
PbEh+9QpyF04j7/sLKvLShqkhUGEJ0R3ZxCJDY9mAEp316DifKJ7R7PVi3II4SGA
3zNDEIy424TQ6YIgHH8ghOMf6mKjHlP8y8L2zgyrw5rYIVnTmR2I1BcBFC/RsLx8
nQNJ+GJWSDtG2aWJnNXkeiQhiZJoxhoFLkPCLuzzR5MVyrKJlvDgkXOZD+jNS74d
iqE4S/C7SbE54wcGeUj0dYVZcBsetBOcYD/zYEOVmbUCLrPOWohodnLKyf+l0Ba1
xvD+uR+cHwP7k0p6oeu0kX0iS6ViqoSCH3O22hQmbDDxz/rOsyNm1A/EWQwRu2bC
mtw5ZCip7+zIUf/ltz5JBPkf82U+GwbbkB6AlUX1sBOXj9U02aK1fEDsO6aEvK2H
6qr64dtfq6/QGDGXd5EZ9AoeY77o4jxmYYMnjWwafWHU+c383Pi0CKL9NusgnqHZ
i5KFPC94e0AqB2Kzz4sQX7h7fMcZZ9SDnOqIsc/jsvN9Z+xrFR/ByNdE6WHtFBYw
sstdKmOkumFfT5mvY3cIBSm7ug5J2UugynndZhJLpZb7p4I6tfYWHAQ/3kjqejj+
kqN8W7sxDhSv/pb5trQPmBD7Bs7b8wo/8dU8SBcOpzsq1sFG+fWTTONnv1B83v6M
JnesOO8Cyrel9Tlt1YNN0KnpZiAOEPJICo02ipsGlbJy3pE5fxiT3cmTgPDVucE/
NMFSkmJ/WwQ+qOoncbYlyandGbjADMG/lBRk31GvJFYKr/WEQjWnvQASpMVUwxPY
CAE2xvUpQ5EhCecmLaVc73rhsWlmeWo0juj9YZEKOI0RB1E2Cqlip/Nmrwp1Yopn
CTAf/KmhOceUOODLB1Y2qAW0n4EVqoeoxZIJ8ucSQw9Aur8ljt8fkkM8vFWaTVo8
59lVb0zGuPE+l6zosoFynuW9m6ln6a+hKji8WSVfmdFvFAC9cHEekEMmRErJPVhg
Q2kugwFwW+SpDvKnfG3k8QBuz1ATOMiDfksRyytn4ahIIbNdUKePquwRLgLjIOa/
c9ygkvoBz7/YLG11lM4EDHBT7iJuk8hegKMgegh3dmGoieySa9wvMxNMS1VQfFO6
6OQ7tjqXP9CloFPiPQ6kTAbu4CnpEtSiL5umPJZGemzLftwHHu4i9lFgSnRBZCTI
Bjn0EGH2gQzVvjrdmH4miIyNkmiLHuvd5gSVrKSdVDgFI2iiJonIq95Lx6sv9AFP
9dS9xLeqKHXEy8Sj/Wxcfk0/gH57kUgEEJkAAEQwnz/nDiRqJFuxG7VyzRyMy9KR
9mNLzU2XOORBiwSHFcqhf2eepHfrmlg3kN/JQ3aKKWeRqeYcvp6bKCWC5ykJSIO4
kHucLuMR561AsRr4YqPV7q6es924FS8gYxXW+OI8/YCpXbDyrssyMxZfX5bHWIaz
UDlvI/qeYoTECVZW04uKNGlHOlIX8YzqaejYS1Z5ye6t83QISviO/71mSmKRmxPF
TIx3jrSLYgQ6FOulxQXb3tg4Jn9bNXSaxAXASzXB89mN+pjid8RicO9XIN1jI0mv
O2W8KV45OqzYSEMtB7A6y9hzaogZq/X5UI1/KHdSbHMTXeQ07Ky3INVvPUQ9G21p
zwIB3Ks1ZW/j2+T8MCCqorczvIEWqpxwX6m2dG2T6vkPiY2ueXXicy2mFZbZ844U
mUROXCWFNqT7Jk2UhzvyvEB9HJRXdyKxsnSRHooiJWydttlBTgCrVMCikUdtfBxt
afPhcInW5CumuFtmQr/eoB1VbDN+xkmQK9tDncbbKTQRQ7XUc/gMvMxnVf4OUBFM
SLiUfzJ6h/eELvNA9jdkxFei5KWtYJiSA7j78btNNB6VKEZWpjkbAWXTORIsYbLM
E008hidUn4zo76m3O0KOq17y9MQPm3MqX6UIh3lfyxgbHPTWKejSk6t0Ap4Jv2TH
PGHF5x3KxrdRphVVltDnUVs+PYSPeYK+NR6H9NfN8nBnRTmmDsQ8mcztIn1f3ks5
dXl+xLF5GJpSLRQQieZGpLY2HjuUvBEUfCSpSxqEDJ8vtforew+ldcF2QAEHgc5V
ELVClIcz/BSeMct8vN478lMFTUx4QmDiZnHmNuWDEqzpm7VBbW4hOVY+D0dM9rO9
PxsUt5b33BW+VPDEqvHrTiYVQ3nDahAeHN+TsLUnHjzGGu2EYoTQZ2d5rxGlL40k
h4GgbQQk3NQau15OHhUwcoMnbNqkvNbjctDQ4kqxV2JbNwUETzbgJvePWLPkKgLq
x9L/fdM9EqZYVq4lrgbf5pxVhxMgiplPaY4+xziHW0J65qRsAW562shiPlc+Qfo4
+I0WKDfNqt/YgamfXhfXsR4az/5mrgk6mazMN3JD4hD0bk0FrWwcst1tPlFBwreI
07+4LL2fC9XjkKcQKQNVPvb6YVG/B3+wiSnyEOVztqTvhUhL3MSNL+2bmqbaTu/x
F0ignMyLJagjvUhoC4Jm+MR+OZAnXG8kpN8pX/44TMuXHIbHNJHyn9nLM9LlP8vS
efcdL1ASm5yZseu6OwA9CkhY62Sn4CMkXlupbIvAniBfLqAOt8cG4s0kDBDfUJgH
uKvi9UreRVIglAperZHAM9cf8LhLbEUXfGnJWP9jN+YMCK/0qk6+0X/+kp9+MtI6
WTbAEyGg55sSg8Q7pOsjuu8ERQ245NYUtqM3Zx1lmrnEY7PzrPXOYq+U2SikO/Uw
OguzurVJdNFrw1GSMO/SvIU2BLgbnciuhlXy1HqyFxxJfpzLDiXQ7sOEjP8KnyFE
FNXVPdOi0EPU/tqsNcgN41Ezy0fzCAjLP4jssSviudAgH8NGqwPJj4jZ/5JYrlTi
EGRi2Y3SQ941iHxHuyow91u4o6DZz83e7rCimT/SNX9qU+41MGUrUmny+STw7FID
GnLqxANLYeHBexSIHPIJNzu7S3BE9Lq5zZU90ZQ6veIVFNsKHBb2mN7jJC3ga3rA
+I6x2n9eYchNbcw/f1U5lgXbEJJU6iL5C2ujdLa1Nka+SLoNz1INhosYsYf6jdUm
CzhbYIUDyDbt2hlYjP3YEG2+ClCXC3C2/ZjYjK6SDsY5zJ2rNZtWzq+Ayv4hROx1
p3nKVqyLzBYft87dFcoZ+WMGgoVFkpJWeBE5o7hRue1baVnbfbhJzrIY2dtODnd2
AfSMu4rlkQT9Qoyu3ikNGjtzVcEV+jc7kJtt7F96mh/KmQAstwKZz6D1NtDEa9mo
GZXl910P+VCzCGsyDXPvc1WCRHz7xSfct+M6G2IAGHxFUlO6AfXE6dsq80CDN5bc
xDQ07TeeJpxI5D2EYoi5U8jqbiMa8HYY9poK2B9WR1+y3LxnFDpaK3SUbj0FEQO8
fQO3fvdvk4CF9L8qEVqZKDiS4RYoON/SMFrhDY68BaCyyG9Zjmyi81xa2yNWII1l
0trDeDKWkbYTREEdG+gpPxMLr7hY7Y4Fhf05zQeVfqXEgAQbDTKPxM96/2MCimF6
cVzr5f+8UUuU0GkgcKGFCLQ/MJrlkrym+8LlX8EDIelE3few6NSgNRAla77Gc+Zf
gIFwBodrJ28qAD6Fu1ztN5ANZf5uvKnefQXb5dORjp9xJFj9NKedoCVQ+ZTN+cmX
e+Mle1iq7GuDWqRWk+hH7FY5bLBqwMc3V3el8HQxh6Bno47av1wHNs709aFdyuS9
2uh5ThXl8gSmYQxBBKzoFnbdTmKQupZ//qjRT+++y20NLFcLqCNq8hWRAi8qzUVF
S1awE2sQcVl9Hx7biYOZOQXIbbEQ8ltVAjRnvmnCry6ttmjQAV2tBy5ACJKynBOI
ZXpkNINfGnFWlaXPtfiLJxXLNDOrVQa3E1ncet5EvA0FRLM2fI1BO6JpP0D1Ymvp
ov/Hagr4znMnnAYwkM4Y/u7Y1SlDv6YIUi7R5AD6WhY4LyqPOROSh6IhgGq7qYXo
C81XH9Vw+6jGtVAqGyZ4R3tqjHIVrnLlwC2Fls7kNITraHMIsWCq4TDRjIGIVcah
wSJGj47kK6HT1UXbhILUvw7l/MA3ZhLBFAxFfTNsciCTWLHtUXLi9eLDERXKKez3
qFniooFTBq1kFm6wcSen0JNJW5NQN5PIokBZ1ojVmQE0Bbyw7pJ3zCInk62atAGS
XOO9VEl+d3Lec1tVeFvGvhzfnBrsoichMITGFFT2PimI2bWiq0dTzyEkE/FiTcVn
IHu7fiRU8cWSQ848LqmvJKsG3SFeJHXlIVd7vdcJuHXP5buSu4uoo8sp+GdaJ7u5
ef88zKaW7jhuqzwo5kdIgAdJDRIPmipvnnGjxbTQ12OM4M3AInrJAInNmiFkjXNw
RIfUQsgl0Evpq9LFr9dGD3J7j9Ez9qJSslf/X/gABj8lbMBodWwtf2LtsNJr5wIz
s7H1LN08YyH3jlqliqZPhu79wKjmM8jBKrFW9qcE05HI2mow9XWiZPUZYIk/+A0x
ehbcJm/VMP0YqFFumikYSCc+rX9nzr9hEshWRcCwxh1n9MZxBKi/8bI7O2vJLrUs
ZBdP03nOsWwrNg7Jm8lkIk1giFBcPQT8Ti6f3H6PuH7HQOrJ3Dql8JeUkqKQlqQk
C8QlHzsoA3bJGOYpBovQYq6W3e6vkpx68QnBCFK/JLS8n66YlkwCYwiX3IesWO6s
lu5u0Lqgwna66h4EtW03G0PAk4Xq0uIJTs0sEHmwU1dvaRsNqS+bvjgP3McKTFzs
lwmesfTVKqAnG96GySuTzX0D/QZVIA0BSOJVBhTy5SI7zEgrSwJJ5T4iK+wpDrHs
6NvbtYWvBdMH7mXpd3MGZ+Bvuty62gHqEsnMOJB4517LUyCLRfl8hXZaWIVAEfja
tXF0Ley6BFZ1yx+86zfNLbnmDS/hcfKk8Xap3xsOxbrr+d3bgKyScNESp/2prn6e
V15HwBMpz2BSyUMjN7Ni29HAiTwP7SRmag0xQ0IfZWEbKoORfBh9MzGtfgYKK451
dwgf2ibBXJT0OT17cwFGf79zI0ak4GcNfiazaKwpzE1P6D2INzzYDqVFpb9OZ3jr
kFMIJrxJKObIqoskAZKTJHdFsz67QymWcR0DGJW2yN0XZRI0baxJvy8wt9VnJYg8
GotWhy2HGjvDUyZ6I4PxqSOr9ZooP3XdA0lyF5ACfXeXjwtrzgi0xE9aGhIc4Wq1
4zhdkyLE+f7EvCORUFeMCgd6alg7dBmLWRzdMl03eVFLxmuWKtUzR3uNJW3VX74H
1rBvyd7JXmTsPSNmwF+oBRd0WyApVDxtBYvz5AxS2rLOuIdqwMYrcTxGJjn+cAKm
tmoXpLSvHl1PRAEhyNJZ/EVmlxbjpOD5h83Dmu35pUSIo/IgXIrTrGvV5ocxa9eR
+QmiwoGzzvgcTGlVaz8zQEFJZ1MyFRNKFGM7cKTvsegXLNKo1AVYQk9Fc/vo75tg
/OhM/aLIWfK/uPuHdXpmqCK+wbI5vjsd5oKGX0ipxU6X5DbLL8JCqQUj+D6Ol5c4
V2FTL9M7EjD3gflmd3wWaSLSvNxKnoVZHxO9VdfvinhqVtbHiPApEZjNVPX6azrY
qsWrJQDs0tuqoLQhtzCnXXVtQwWtdj0MhJRZFxPB7+qMQ01IOySxk0p9l/3KRJva
X4viU0tdPCBB72cDuhhw8qQfESOAmCGryhvBDBXAWJ64uZMh4oH7ym7AZAR75NXd
zXej+VZl6SG8Wgtm3ozht1BfYZE7NRcj2mtEurvFicoli0Q0QFuWdtjpPGPpbCN+
jCcd7dPFuE+bMzJzvy9FSbQ9PT0lqDnkzuuI7a/5KIzny+ckarcmU6vFIGfq/pQs
ufihh2NISG5qVf7A56tV/JzoZohpJxHVwqyl3ixKZwZhcLL1IW+sTBVOCcKAnjR+
EyKz0QrKpwkmisuVTTHnK8fn7kCdULa3P7P45abG1P287dT448F0tCQT5U9EnV6i
Ssp9yDbakB8xP+fMpMnbNcViesf2n9AaYLc0YlhozQiZINg9jkLeXInvS4WWfwgT
UQ6SX73J3ku2Kv5ktgdJvpB77tNorIcOLgzg7T8f5GqOIoo9tB+OVVeW0FlnFIRZ
DYC6nzLY0RPRkjBrCt8ZtnNa6BaYgkVuqntpTo4xHBZzglOvgz/pCN7TEQPTpOwZ
7lTq2d8VEdttTVc4+FUj4836hGjwKQUzmHdrS5aAGx9i2qUbfP8uyG2yk57eG2VU
tRbhucI2hn7wSOywF0p+QVZaJH9gM/XCcWf9vhIUN28FXI/oDiSgkwXWBxBDcBGn
WpjEwphtnV0t4Ov1A/WMWaqEdg+tfjeewx8T1dPIwuVXrsaPXn9tQlAQXEAJAtwj
BzdulPjrA0Znd+TJGrXCgEdK8hBWu/BV1XbkpMrj2JZf2XNXwzcwC0DvkDmtpHz3
CQGTl01tZKqNQQJ32lrT1kd4WmYPS1ObH9mgQ+yWXBxRSoxqihZ9chO5SNcVxmgt
P/nTdoQ51k56rBAxMhrfb1Fs1h6oE7vE0lA4CdNWLOaL+TLfE405AH2SlcjFAxL6
T2WlPDUL/HZwmgqNvKoQiYqaIL/V9PhNayVCBX6NN80T1vTlIsQ8ysQx4o7/lVcN
vdk6Pl9HMQ1WZiZ1GAGkXYt/EnPlm7ISuBJ37n8/rLW1qCtbP84XJS5gaYkfQLD5
5JY4loMa2OuxpNVZlXjaGIEfgmXfTcCw5CissAvqBcnQu9VmSQlcwav9DDCgiSH2
ZtlCjHGM2Pyw00AFBVPdkVBqisEbgz/aXxkYM3FR7fpCBZGK3qHc/C1tSC7OpZMf
K+gL+Pzh2ektOhp4mn4x2AhLZR1WpV1nMtH8JcKyk1/vH6XGmoI64aV3rFSRSC8z
RbhjwG5uHV8xyi7mZN4G4LXpbWErWeTzFFI9pljceZSUWDR6Zu3Q6WS4JT/UM1iW
kt7Oc0CHAl8wQ820Z46+9xVOV6zat5AcDhdhv5pCzgVrIWkMEGNplL2EslqKiq9b
/LOuf9yQabq/GUY2frT0vW71D8FsNNr8/vjvrkTG6e+gUMvOL4IHp6k5MbgeoSOi
tcrD8L4KMm2/cHpe05+mRGAtmG9I9jPMZLLzhBmj4UMqqJ+YASeTnTS1o3QAwaVY
0NxScOY3TF6sXaGMbGLNGa2PG3EeRd2o2Kq5ZmNZKsqKRxW+5mjCs5YIMcxDFwWQ
MMiaG09rYONVi3VzeGxKeh0h4c+xHIEtxrawRkq6NUGEwbTX7BSLOdHt5vfBNcNe
nwgvOXs3iPFMTkB6kVp1qRhUWqLHPsYDd2Y2SfJ6KEWaHyYcLFL9VqPY/MYX8QEC
Mo1wXuCRY/D1X5xCwEYJgSByy5FgcmWH4Q6jDiXbRg624Pk4xxwRVvQPmnxZY9zU
XFnaIGsIWDfOAnNcq5t2OjDoKWvLeCrIBv3tUUoVP00LBeo3vOQ8T7MtbmvEcSWq
XUGSEniZZWO+9UpgCylqAu9rpADLEW3UAMv/c4xLtW9V/Pi9rSx0p6Fl09RwFv7p
/hrX4Glj3vWv6BxPX/kv1jlo3LwJPb31esAlhv0s3MdanhSNWwjTRji88/MasCzh
y+AKu8MUuTSdl/gSOYj6eW1hrAw452Pvjn0lgNbBF4R/HL+hyhcnAg8Gbdf2SN52
S0QJg548zlmKd/fm0/dhOY9X/J+A0+3ZEe+9NeuHsT84pZsfRK4fghOnEKvoXQf5
hCNtUFMHuHDzSBwmjOBaHeGDEtuCp4tkO5iUEpwkn5J4XXsL1cZ3OYTp5sbWw+lj
hO3nmXKvYwYr0NizwpOJpAZqG2tpNSu6FXHy6DVPiW5SubvAQt9EVG0YlYY2Zy/6
2Tpt5tRT3GZVUgpF7w13NI18IQtE3O5KR51uS8nLD7iqL8jR5CCsmR9xzR/8NNLL
XwV+tBQVo8GAAI1Ll+MQgQzy5OBEHIxN8Ytrm/tlbhh48P9/horBfvloisU4i3pq
2TYLKG79k1gsha78Sj+cGYHqeg+aaRRGdYw8ECoxKzMbo3GgVfn/eQ05sy/VqxGM
cTQLQeWNcHiIuqmF0spc5HM1z2ITqY0U3r1A+ONuaQ8njRrV6Ti3yUJby7L6Y6e7
gnVtecV3UCcqFYc4HgfxvrRkAc0A068ZLLgs0XBBx8IbmGrbWQYx7bcXvYbsnaIQ
5TYJYQx2iRdEGXGwArZaQpIEBKVXB3MugV7yZcsS5Z3ukwmP2zfcJwCeHObjLO8z
y1p16PvNRsmQDcwgJDkAnLS1MThl8kjYjeKP/xMmvLLMyi4+RAzU3sFOxiAibLXm
NQPNtTnJgW4h2xZBki91Lox68KlVH/lvMpZCY3fdTDaVy2FhTsXB9u566cJiJ9Yg
Ir24N8G1SUaOOzyspsbjUA/qhKrz2HIBapljOHyT4Tj6N6M/Z9CoBu716lPnFAb1
YVXJ5Tc7KF8bGKUpMcCEaWvVw927IgcwRGNSySr00tV1Kqv+wClA1m77xlNlgKGf
Rmh01unN/DQe0hNnGDJW1qW6BBLDqDp0q4Ii1WkO9u2UzlFO0mrOzZBgDIJsTey9
+0A8Pe2myC9HWEbPFKJOTtHgFARo7/Zw3nH8VaBLGaYX19WxhUSv22bLy832K3+J
aydhkKhgErORtR7kaRzID3WH8p41+NGu6/+UhT3qM39+s1VeHBtHhwAIAsMo2BFU
M9ZqgL+Sp71rusw99yKQJhkRUPsWO7jsHGDweLboW78evoTY+jjat13p6QuC7v+6
zeK7+TBpbbmZGnbBw2ciw/I/5UVjBwrnpWmft4OidFPdQulyUZ4dZ/4KbE8iB5kW
j8CsZNXbC4/3AmKhZ+JcVtMEFx4oObUY0mdsIxmdVrkAZttrJcSUUhPjd2H0GIQM
GrgQVdw87EE/v4K8BquoSPcyFgGdj8G+J4ZiWZlKCgYXzzMXpmZnl0HBvSIKw426
5TxrC4QWS3xyrCiEcv3jcivyaS95fw7JwnkkWAsMWm1D4GDK+kgTnyi8HwwiAqM3
al9OQzpycbQEAtUySKkENXDfknZUkJjivUOgMqyOFlSB3Mb09fpqckEcAmOpFdVt
DXNLvZOeMYzpTQ53S7dtM0ig1FdcTyAm70LHCDLPvZLajlDbQgQ/hGWhkbonZuRn
4lVtp0cqkRpJb/suqtbom/wi/haPkDl7vMvkfYkGHR3UvD/mH7amVqlU9IzkKvWC
YSBnnOz+gRl1OR0T7oJIG2mKSAPXjysjfl3CBYfixVW3ctmkLTxEADQ75WkNlox7
pd9pNLp9Z0VmFJDsJwT5qww7bHkb93F4bwgyN3VUWF8qY1AK05wdu0QkoP9uiUd9
17upjUQcOLcSA8E7AiIPx8uHfEgELp+CBp37AHwcprQG7YP5tgSDWwHwPQMKtHQ+
cc8v7HsGV0steDlYEExMkhFq+aRUVV5a0bRmvWi3Vm+9fA2y/lAcFbApYdEmL5L+
cZbGn8pkb2+jPNqXYRZQYb2zM4Am8sZB2xOfvS7Xv3lbJPfONFDZyeWE/9uAjTDe
YrUhWwiiiJgoBjHm52pRpFBKcA8a1/frtJh993LX2gvWK/JuzMfDs137B3KU8nUx
MwjfwC4Whxz2VouDYXeNmAc+b4E9ctakGhhNDc8ujvywHeMmsFDnci/XjlFbGaja
U1FemEyiDL6sPFJWhyxtrTSCWNQ83y/Fe+pMBSqOiw4HLgAa9LJ6N1+SRaLLk/ft
ZwEWFGHwROfUdG7VS6lNSHdbD2g4ojD/hCQ++IcsxM7IAayVi5fvGIITetH/OJx6
0nDDDCNT118FTSZZZwTaHHzwfqw6KaQTcyzYUOUKn+uMvmosxAsdVeotwhfkvZ9M
zzrYDVZYjVP7zFJoQQEENocUaSS+kgmV5bhRGZeDh85EbORm2bJN9ZdOxKPMXmQt
EF3fqsXEARRvFlIJkVgOX/Wj66lp+2fy52i0Yas51sxvczMRzBQyau+8idwmTNGa
xLUi+7MICvuTvs34wI5FicPlviCDRiVKnMIGg96ei8UBwO2B39juvb8SH8LzIEOC
YyTDbSTfDXQPNezYxvAL1UM4pBUOuYpVcY1noXFCAAgN4Vkm3xTk1PdkD9cssxYa
7w9/zkN/U3HAEmuej1uq9UOT9qrwRDbWxqrTQMrr35NbN4CTxPhoa2Oumq1uT0NK
h9u56vAIIJ+7pJdgKZaCy81LBd59LPShCVb3ilgI57jT6YBR/umXIAYA6Yhauy6e
quU+uJDbTpFSdbgIHI1DVypQwZZ4G7cwN3GnhXLa+WGbRx5D827rYhtn2igSSiS4
r1cfj/enW9PVaxTp7g5XOPo3wuY7QEcaTwji40N93rUN+4imnrK7nIxTs5css3e0
K/x1y3cdizHVWELXNEBb7SvoGpNsJLs8Q9eif8RreqZialaF0aIebN6Rcgjcj1u3
79IPTgcN4vsRRzhxLvSzmL7gNxnz/fWbqnw6I9Il9pwJ+mRal0/Ic7GID5lhu96O
p75xMeVfn+heSint/Rage/N2awS1jQzbn9r09y8OEyCm6kk68hIDK+yzUpnQkY83
mwFlQCa9Yk/J4bqDVKjyv3eR3/n+55N2z7G4CVQgXsXzlO9CfnUQxJx4UnilUyPT
538LonXLvymODk+ytOA5OYBFeEWkmUZ8TlcWTHUbxENXU92YQS8bi7O24k09JKgq
GHx2oMunK3YOlkcH504He5Cntp6bVQtZbTQpggj2rx1hBKviZolmqHLtcNAaSIxX
jiZ19knCE7dTay6cEMH0HwR4w8CJ8VhfgMSTM+6J1LF0rZ3t5yDMcUkSNIDX6OcF
JNh2FUjjJDTCNu7n63UAv+IQYmcfzEKqx8yskOParSm13cKnR7iZfezku+yxwslc
iMSCwy/+RxOHqiUjGcGi9uW/LXp8dAcgIdYkpiayt7bqw8VVFaUOY2A/02CpWjEP
bMMRABEXY8xw4BwCK+CkMjyfgpb9LbljKIyHj6vHbFIIFkoye792lTC0eFhYHVlt
+Id/4+tgmUnNGrTrPVtQP6xIS6p7A613gaI9IKpJD+SNd2atSAJkr3k+VTlwQ+uM
4RRk4XCm6sbw6492/FCWPwpTMC+97+GpkSUNCO/DqEyJmTgm4NPt03NN2SUzJE9k
uSkiDqU+GFoCOca4eavmKb1ECmiyeaD0++2uIv92B8VgK7HrS5px25QZb1ZBveas
N5GVS96Vk9Fs2BrIpAeyKEjp6Xb6Ib0KZgFOeCckF3assPLkAkFofiHS14OkMnrK
8RqsiQnNadOIiLWKOn4JQoLnFIL1ORGlnL1AIkV0mQyLimuS9/A1kQ3dncoRNzLl
27dVpAoiIQRCUNSKHAQeBYPcDpTSWTI0rne/16ipvkrf07thVc0wbFWkoG2jT37/
zhMd07y/CfNLSaKyR6yDbFHjzg2cgLdlN/mcnhJeV+Cdd8/kuO3Cb2PyHuZmawRv
RPIL2WTGSDgehFZNvLfZ92vUjJkP5R1Z8ILUhlvD0u/5jfwbWErl4YrLoQ0laiYF
V4iEjLgAB8obiGINDipug2YcZ9vEBHOeDEBa6B2ibONdadZLBsDcX1bx8mWCpXUX
oHt+rsJWCM7ZG1lBJUb29SglTfaLOnVEK2F8H9KIy+/ckjnHRwXLcRLEC+hrHRJ6
ZokcOQA36UqwWZoHRoktK5o56NtLIiJO3VecPKQA78Qa0Zk6MNY6enE4UKaO5Wd2
gr4ZMNtPYXU6tlEMnFnmeh3ihUNc7dhgFeZG62bXVxtiHBcVTq1oa7tsZfRpfWKI
ijS02HlyJcAuiEKV0Jw0QH2FUU4nLR6UHLRn4dkjj6BpoF0v3c4v6VoOyzmOFBTK
NIZdCwricIWp4bLCF7+Pqct9U4T7aPCEqijZQd8pwm4/uBPJmJWdaQNegLmLXuw3
lDzCB5UC32kWz1yxZ5+AFeAuWqxjtaq8/NtYHEXrzvl1Mlx4ux5IPhqipQ191rPX
NoiynT8tWij5piTAgKH6AI24eZJoe0SmOoSj3IzOjyYAesi2CR1OA7tEqUQNoC/8
tbRfY5Tm0j9IbKk9ZAVmYoXDUi2PXJ+/7Q0RDzfLv79rh/al05aVq1L/p3nQaiP1
l5UfqIjhulAP9sxz4Zl/qoPh4tYXh5TcXcI0yefoMTTcgguQ0g+teWNCXmbqPmwQ
YAUqAnIwLZfUPHmaDsaleedjw6c+9B1+ToWMt4uCHfEo1IefYJrfvlYzxvTKvZSC
wXxN4zazngQIUxeZDrws75JK+ipJJ7LDC7ZWcglm3u/b0w5goEO0hZBv5dwID+G/
3BGZFrrGJ+3UL9JxGjwerchxFfZTKJ4LdPJahCOhTw/dojX8lu03rrC7NLMwo73m
Hkz2s9c+Mx285QfXV0b5mcPZR2wNdHfoM9B+O40+A+DUW7Xufq5Tkys5NcmEFvSE
L7Jku2xaWM+qAs3F8JULXHFDha1remuLKISeeDNtUAX5aeHfjbVEXbGb9/Cdffk+
1L4zQ/fDQKSFzAHMr4Y78M+V7CDxBVdVAvGde2ntq/iQSLdDW8Xidz5vcVG24fjp
U4UeMceF+/N/IBl0YkxgJMNHQFmB4bj10Eq3yaUWhSg+gVJxbqnji3C0bIYi8GsW
Tev4gR9LbsLpoyZvx+hJxM710gvqs9sRIJog/NwRQRqlghPUStiqRiwahX3ZcGP5
rH+Hhwyob8y2DNZS5jZ1qPQ0j7e1p71bawRWM7ZnQsXtRki4kKot4LUTuVK3syNz
B8UJxsog3p+kwjcUo3rnvcM1yLfpVzHqnjyvwLavJ+OGo/f/7yQ3WniOL1sdlfZ8
x23dYUIDcDLHCYXkeXKsvfHQN8D/YQ2LZcmXerNMBVvjHXowAHpnNy2WzyIVhDPS
ruaeD0pLkyMOzcIIYzsFo4frnxUydwnZpSWY1SeQ5tq/a5Z0cYogAoXnqosR+yI1
2NUCKYN/aeGSbNuLC7Xd1ILtezT8TjNctBlN8962tmIB2fcZYp+lqJARj8spUiF9
CDxFMZvuJim/fptDUCSNl8hK2qFzWM8NF9T01ycg5QHNh5XHnrQM4O4m8q35xpi1
EYyDriXl9NS4bg92ZaAKi/BrUmuUlFC+vjHhmmTg1TWmK1/Toa8U9MwpASEFNBrM
fcAzg72tBRL5Z+TPP6lb/fz5V0mj5oz7T1hamWuiJvldNkrNvPTnIaLy9fnHf2cO
a3T7EuTsOi7bQiG/bI9gAHG2ozugBJgCKn196mSPRyd8N/tvlZEyoFWyrnQ4fHWY
rfJZ3wiVTdQRhQ2FMap3PzCFOuhxErWxiTRykhP5wElTLHJKYeq8gGsYeepWnpDh
K0zKuo3xPeEl3ksvctt3YUztAkP5ORoDyOHfBjQeO5KIEXvAufrpwtQ8a6BUXmmf
DR9G6wMjiHvViX7KmlD3GFOi83SItX22IrifDiYNXn/6tDITCj04hycAavQzkEZi
gVvoLzzcxfYK24bYdhEbbEChc7Sk64Kfc5pn2p40fFH0uHujd12uzUkFHOwZdLft
l4b46uD5fYPzPbeQnYnWDGbdk/NnrVzgpWtlWVpNyUhJzeUwkHOuLVEhEmKnvfK4
IHPgmBu0gEJrydQ2wf/6/AOln3r+lqTbkv6ymgS0fGLwgrmAjBYnCow4Ze2oksPF
A5tAPNvgXQP80ZaNRgfOW3XQE0eg3AFWiF7b5ZOYqW7uRkQXb0zQVk9uQsWO8EAc
1bVUiHQGAnEIL1qpZ2/eJYobpo0y2TTHYNxlOfax9Wcn5JXVRZ+PQDKHWNRWZAH+
Ptyq4/JlWd2zfHT4dWjYNYUzFzqTTkNoevE8uwPpz7gyK3dIvw73jKp5Ejq0tNcl
qIh2dCm/xSAxXkCLGCS9vxMM3T9BAft8Y9aVl2iWMzHYpYoh7kz5bob25dZ0qtvx
f/pZzI58BYtA/LrlF2hoaopNFhyZSKn0S13T22rXOJ1m+7Cl8lyTuCLECFAnC9Ji
jHulh/tmGK56xpAq0EcY0w57U50Q6jJ20iDQBJTbrUMuKLWsnDY1ckG7BjIwTKWS
RnfcP+Ivl8qNmysBTOMHwol9b9+Q5EmDzLlCcsMhFa+/q8f2948m6AbnwA63S/oV
N6efzptI5wMqyEpQJ00juttsMkNl2ziJ8Tdj60EPjKK7fRinIqrMDcgiCw+lvryP
Hb4Txon4gyZhtorF/D8kmXF+HjPtule3eImqOfKWRqDrDOhlagUX+SFeMDloCDHr
4ZMqk8vMiOvTh6cT5CoonsLbeGSLJVR7RcPQTqk+2u8+c9Y4LNPCF3I8qS3FVByK
9nkATkg3zn/HaIJq85yPnbC51t/uJRWO+85XP1Dvpb8/GmW/LXxua+aldV4Repz2
BM65362sEMREIYGc2KKOqz6fHLBVhIyWFm8FEe+O/by24AWW5odTVnHQ79ZkKrSd
NVJQMSGX1dteYqHG6VMS5WztBtNrbCSmbSjmlP0SUAliIEC8o9JwAwEeWA9MTnKa
hifuZLNqfWEmMEL2xFZ5SOHg+rbgtqTJJqJOQU9TRtXlDd0YEJhBl7y1y7tTEyA/
3+47gnNwMFc+EpaC6/qdjhz42bHDwT4iODD1AG+26VRHG0aQDHtQDsD7qJ81gbv9
9ugEiVDCn1p3zA9/Yp/a2mJtQrTyieKCkK97jGBYjpa4O58vFEBe9kK8DiFv/jbc
JqUfGGfWAHL0uOxZuWEvRh7fRjI0tmMfKmpEPUCBRazldoMVgHyFdzNmxWn3i7Y7
hfHVs1Dj7GsyEu+9hXAbjiNhxzgRZxIbuzjB70mzWANWZIOnhoqsCAk+0syfJYoa
slYINtqSRF9ZHNEcAyWXT7OSnlHHIimdtN6GZKbapMYNqASXVWWJQ8J6G8HR6tte
2dZrKI+BDNSq77q+anPPv+R8gpRmvchSegilUImU4kX/Ld0h5C/ZbVt94PMeLr8W
JnUQjRH7538TcoSDKF00WpNwvn6m9h3RVvLaycKzaqm8jQd578QJD0T/z4jJhQTT
5bjqsJjyJ6v2E+WigR1w8nNWisEt0R+inEsVG2bqY0+o3+aP5GnGl+apupw67SBt
NPgYNVhfnXfoOTlpwdzczXgiCo8DhIfM5f8BNCFcT0RYpe8HuEvq6xqEj74HDOW8
x7KyiQxMS4BZNaog1hwp77zWLRsz2E5siE3yCBEsUUoj0NdAQ/e3Y4SOdiS6ND6D
YbJnMOTLAcQ8a7X1eLcSst8RyE5cwNPBEaGQ9LueGzMkfo2FqKq6HnBtKh1Hnm7G
s78TcOY+c1k5vQRCVH6Sfm2A8Q2Wpg8a4O5xJ7dZ23OMWg//i6xcUb8K7PfngqOF
K9RYMWCW+OvqeeEfqAhbFvPCco2WiEIRWobabA6+V+OQFDA/jMWrEDLUFtRUMGrr
smG63Nk8gbaFF052+TtChf+AqPwpIwZw5QwtwWDC+enJf68XxFF7UGkXjUfgP+dw
y/pWZxI8l5g5O5h0MtoYSpYfTYsMNTxgBnUBvLeyNafbJ4yX1IzXaOqZC6iN1rcn
xoCW6cQBn+0hitElVjsUwHRtGASbut8vSQNZKOE2yvUJoyISXT/XMYNBRHb3PzTZ
0dpqPs6BcAyncgMA9Wzts3b0Smzv21vZSdgWfj3axo+BKjjKoenu8e1HaCGt3tAd
GHqBPM+eR6KRV/GDjAo5G/qrA9xULRVMlGtCLkfDNzUTr1alpvPHAnR2uVpWeL70
jprPRqEAkfica17jCuNmXuMB7bqRjYwAvpxgN8o8HzdiA4BDHUWGExQ2OZaDkfXa
IUk6irWCu7OHRmVt2YNF49/F0j0gtnpVHtwW63C9wYh8KRMPS3U7/9GCYtXE9zJA
r2PJM0z8susmSyIzxuAhrI4i1nV+eyQ16hoDnC5W/CUGcQtNufFoM1Fnlf6bVAL8
4EbK2esFtvqpjIOS0uUolWwRZiMWHBVS9V3urUGiJ+d1oA0M9H/gK7jroL6hUf7h
OQDko8SBiCKWgt+GiqE29GD6hW6RUpoPFCO3hgexp2UABO5xD9JzEzx+nuENXtqf
8sM25125HKhFjmYPKvvvYESozA99W9PP3INXlLE9rm+erfdZ/twwXrb41UOdY4yU
XgOD+NlmrJVICW2HipOqVe7oR5g+ZaX5TzS8YXAt1u1c6b2YqiffX4tmXHLu2w3/
3yEh1QcAgtP4P+JBGqfgb7BqWseaiurQQwxWxWmwIzRhGAdovBv+HevcrUDT6aWG
GBkTPitq0Ah1QL2bmvw0Bfv3UXwRh3RD3yFFgkeQ12LJYmBSnpr11z5SiNnlVXO/
vUOpITTdB8JfRrh2oKsshT1M8AKa0mWhMqVtbgQN8Ja0AJ/zshtDiaBT9WAnSZm5
igO8XUeJOAgFnGK7vrpC81PXXK1235b2CGQMU7wMivhypwOQW3exsjAWEEnXMhzB
3sQ5r2uf6Ehw6o72zx8DrATyjD7mAT+Gd6aICdw8f1S3Wq93k3nT9X0/o1qyllbb
r1we5t20JWOzzZQcRR/KOnPDBchr+qa/qj9oWPVG3Lr4MF8fto26Oe+Te1DqsYDV
R0cGKgCddG4vU84P98lh4VpmAX17IGUrPHTjpjyVtSUaB+I4a7zlmyKey+Pwe7vQ
VzreRtBtYh9JZfwkVq9jJo8M2071eGLQwuhmTbNiVjF5mHecTdAbCnhPkOdAMJU/
8+oWYOBHp9EVyGSt0uy2auLRZuvIxuw0tRd4hN+Q2KZrppc3qpbrsAkob4HYZuad
DqiRrnSHbyaQm3hkNOWPns2kenSyMl2MammAnDKIeFfZnQa966WemaL9izgfd+85
vRIvn1m+YMYCKF7ywT7sqjmEOC8FP2m2khQpeN1d+lOOm6X6DymquYSb3N+KvJj5
FIxEFG5d50Kf4O9LsWUvSV6pHWlwzy9xrWOOLAt7rGL0RaBqojOx4rnGB+pVyfps
DFWszHIyEO4hzpA1aajCMKvZiGF001yGf6njcKIXVTqKtbcF/SBVchsWjy86w+iV
XNENBojmU59XegQpgSUvw3XfijSMer6ZkjC+NgLXL8h8YIlLyR+E7XJZxcn61GSI
cE293v/yUKSxQO7rKAzkb1WdTM8fFR14GgOEGtx3efrw4WiMETQrv9xQBVAWRkWM
n76yXl2P0Og+vsDo9y7dkkckScH/k2kDN5oCavUbXV6hhUNEbYauDUqRAOxyVP5E
qLRUYaP/9Pum7BQ5C4DLn6NLSY3MD8szvL9aMgBEVmwnvqNmvFAscwGM7H1uKXXQ
3kTkyLkJjTN5IqkAzbAXkCnzXU8/tzOV2Wsy2hTPa/0O9y8y/pjxfb2nYeAIxt4y
7aMrvdgklmNa0/Esi4ULde6N9gpZ0pOi6KGyMgHXON5d0plBottrbOiy9su+FArv
ZEjuzGPJuTCym5wmU9jrux9JXPG+OdYt6btRmIG89rX+BIpOasela7QWUQzh7I+M
NXCG5Q6QBuZ/aOKzPsTGJpzSMT6vLaEmxoFjxPM9pzZwj76IQOCjzyjkYyJqKIgR
hdurtIE/WBea9JUeUv4uzIovYIMzokgZ3BuLebEORk8QIFr1GS74BOpEN+MtjrFI
dGl4QlDA4v+x4vUHqPEI7ekEDhVkEi6SSGfBwpnqC/b9sN4MngK9oCI7Uogb1TJd
/j42PLH8A/xipICnlh2uT9IIk5ymEyT+7PqXPxFF+8K8XuZAPOe4mXMyrhoJ4ftx
HEL28lQCvaUqBkhCqRvE2n9au/HSN3Ej9QTvoRptHxriTS00+tM8+XKRZpj4ec8+
uzDneDSnK98K67SuhrTklnaI7GaKPbcwXDzAk6fHNXfVhLPHOZcdOvC1pMG3fO6C
aGRMY5C404ZLgtZroBrxeL9yRXRifWAF5C/N4mSLCYRUoh5c3SCDyX7Wo1F+k8H3
W44czRvHcuI8sND0nQ+SMe54WRdUFsB7PUoznDyc4wDAKJiepTqeBPmzzqz+QCVW
JHm6FjK+xpBwkRv6U57vnfp5HblMF9WEAOie7D8hXx169bsIuy0bd05BjGX1RIr9
lFohLJplFF57T1Derqq1RLEjwNb8z8wDzEn2hnnYhN3MZ0O/bZ5uTK0oIkT6LL+g
sHfiYuD5d+31UKLj1Ghz+rxuG9z4uAvxGMkP4CJCg9lT9yOqdhMqc2rptxv+5Zyj
B4ieQrX2PN9pwvc3qHYiI3y4/MPg1mzxJJsluQgVPeOXD2HStruGQd2r+dtE3eFr
rVmFiI/2U7YDC+dm46ApEOHzELEdDOp/klbyEGXjRSQiLxVgczQTtYl9I0yQ1kyD
GduNoWGQjNP4GnXcJ9H2kqMYK45qZ5AG94l5oKD+hXjL2VdaSaKDMA8B1ndJkYB3
bYGhMK/nXqd5NdUqR/dQSWhDAHKDRgK2Pm2ItosVLA8JW1eYolh8Dki9tP8+PU5Q
V0blXiHYLiHGrke+kLu/FzCLeeE+v8gpCNc4kXfzbhFDqsM2pdG+MOjLD/bwUZET
d7E+M6Ffy27AcKtLTzlS7uxyJvlflbfRdSAU5NojKctZmdZyuHzm5KI5C1AwrE2v
K5n92waY5tlfQmWagN2A2Z0twQPuy7IbdRHVYSl5xeKqGA7XRJ3QpsHfYTB45XHv
N/8HMfNJFCYqLTtN2nX2DRftg8TDKhXulGGpmaDQRVdTv0fF7AK541VuH8yUqih3
kc5i4LHMACPQV/h+0QcknCvQzmModSMB12zMVSqoaBR448YDiSyMVOt+d3vrxaIR
u7qRfR/fNOkVF0phVhjlfG7Fd7sbGJLnT/b9Uyj5XFfbX9lHo5hYpXlosC/jkVWe
ktJHmhcPKqAtlGey0E+mEU2DZkW5hfzID6/IN7cCnZ+fvGgZf8sg2LbSUCLkztN+
nXtYWEUBCkMb0kP7r+2CqmE1u96+LD/dZSpd5L0jdqrJgJMuoI+3Y9b7nowebYC/
NeuumVtffAnTlVMxUFwDF6epkfqOFXfIUcdjpGXJG/X9wNi6xMI4Qr2/9BVKHyzE
Hh7wZCVG7FkfBFCuQrx5WiF2oijE1H3mGZrxO+C/a6gJPaElCq0InHHifpAugr7o
7g6pqWfdTu3gZxd8fgYEFEhGX4qfmiHGUGqXWWd3HyT/5q3l5/8I/ify0PIH0Ryf
pgGU2j8eGYVDHUKu35G/LFkHPvI9rjUzHftdbUWiQYMG0wede3DTRvCa0EVGUOWx
TPw5P4LeW8fQdTwNPZzfXcOIyH51BR2DC0n7X8NDwJVH2e7MfsVYb+ssqQus8gWw
zLIsYo4T+9bhwgi2h2rvA+JFSrL+Hszu5wauHlrXImISHD48YO0lwk8B2cGwma1W
HXzI9anCk3XUJrRJ4KgR9vFO34joS8irZZ79WDMbsEgibOGeLNg+iuFc1WhOr9+y
CpfPRdfn7uNApykw2kGjOEZDRju+O6wsDhM8iPHpuAdRAQg7lDpCloLpj/Z0IQmV
7T/NCdaZwug5pZrNo0uoNF68+4ohkr7DslSZlAgY7zIF/j7k5ZHOQ6EFL5Qg86sa
2cU0aO10IAMR8znS0GMeMDBJfsN/OoYbvKW3NVQH0S0cFgpaTsefITTe1bDqRN8Z
HEEC1sz8OnJtfu+W6xLW3UPKS8DM89q1KmLxsOmGu4/XtlpCG9ENE7WkLJqWgT9x
/MsF2CISwZhegJymlqHqSagL6VvCk0KSov47VEc6IXBc1QNgqbMELJvJtIUtCecR
EBi6K8/pUVMum8aWa5vTrxJWAzcwfNGkH0UfGCkyjHVaKoUhgJ/Xd01mIdZbdvf4
PHZb5Ru7GcY1Ma/EdSNix8zQ+yJb7upRIwrgu1L2sVtD2ov8HZyB/iqZPIy/6vv5
WoEnx82ybH2QABmNe+4xv+KU/oIrNlKj4Y19CQd2mef14bHeXQfHdCkTiOCfEwXh
tT3NTCUk6jn3OQ66QRvwOggkGalsvOz6N0xYaH9DZfj7qWmrndLhD7WXKQQ2k6Yh
VC45idOxZWex1OxQe1P9crr0f2P6XLKWU3Kicdbx2aXPUTFIhgW+4E2aCkRpAXyR
30FZAmEcgikLH8rkzv5BEY4KzIUhDYCuUol089UagI3Z+hNFMaFH8ojkEK0FnjOT
IO6/ttZgeLPUj/7F6eU72LTQy1FlzXVtCFRJ+HlWnv4NYZTJggC9QVZF4kB51JTg
+bt/bB/bJNQ3jr8xn6lYwMa5IBjAE6lRy9fTZ/rb7AAsSVeqwwkgJaxHqx+17c/8
B06uHw0a0EQK1OSQDDkTcM/c+tg2ieVHoDjw7B+LnHlNb6YdGmmLWcmQ0hD4xYBH
ri4XyNe+WUWW5TXsUXhZY7mDB9+tUP1W3zVN5UAwAmf93kLYoKQ5YrCr2EQ/VAlt
j6AmcXoO9c7Si+UtgJ31fLr0/Kvo3GRNlhnAM/SmzyZ2MjofA/lciRvRlUaxC1q3
e3+BaJ/wtlhzYf73ZEy1mBfDg6PFHsAUykTVLVPXFUsE0DC9SvqkvdbOtsSDPSel
r8nvyqhqro89gX5JC9AXFXP7Y0JDThyhRTknfM011Fic+TdxqDJl/cZx1OfI9NbI
sTOlX/xBRf9iMeVKyB94ZML75S9fN1A3AlzS63P1/EqddAhxYJxdBjPdQ7RG6y6c
P4LAtCpPpBJEBsqQsTceWTre30TVSKojabhvGnmF/TnM68nFyUlaZReYG47tjUVx
+0QSyTuUFyVTzLA3VHEMCpDKpUynMqloIFM9WWp8qSNAsMWo4SDhy27gPS123Eef
JdO64Ohl7aiihPAoaYoitldPVh8bHpR069E5cyrrcXCdphN00YZKJr76o7tGafmT
p4Iq5WLmsVAQpQ2DOJvj0/kvNGExzvMJUUrLVrD+AZpisESW1WOWOP7zhfMpxNh7
LxO+WFMjO5caMZ7qBelFXoby2Krp5XkEDOz/Uem7V7O+W72kwIYVdg0mszgoHPZC
77XBClEtlkJUhlkz2IWprlFDOXiMv7Y3w2ZHB2Zk7SSctIbzl4XPIRrj6F7qmmhz
TIOwdRkhdak1zlmzE6EVm0ESudoku7IyExW7pINMfWjSptnwYw7wYW+C4S6nmWFm
3wueJgt+8/o9d+YmAGw/3C42ARqjHv0DQL2iLABDD9I+wyVl0CVqibw3bEer4r5X
j63S4toagdAA/Lz4aiYInaHo5dp4GCebDSIjdPmeHAr5NzZbxN4BqIXFxb78P1Oi
Iotuwr/xBrKJ9PYZOVI6xGHSyuEX70fh6MqkeElNXQ4Vh7JjRkKIXXucYNC9DoPV
WmnV543GSjEp4XTFYYoydyEcWTG8mH+MU9WCkFLrDB/Zbrql8Mg9F+3s9D4qyVwR
tWO0x6xcQn5saZbYgWuBq0tjxZuVhv1SP4EH37aO9RsC8hQsBVxo1sLjW/lgsI4Q
SGK+pptzphI6YF2l4Q15nqRBAwZ16yWq9dCDI6VF0FiuECDMBlRlsvTvJUtku1ep
jx2zmbza1SLO/jRnBztVMliQmvegqGw1VrPUJw4mUVhXNfVSbb0aqnIIWIYKlApY
eMQoLFKLr4iK/I74M5n8BUntMlHmBG7gTnA3Xtr4Agwq+K5NNAQt7+3Q49ZdIlPU
T+N/v99BHOdlHVQ+VJwFV9QCYjCPQP/AeNRSyckmVJ+SDacEC4Aegnm1V1SalMsc
WOQPPeDoM8Afv7JBQfbSJ8HjXvWkyjfm1mCkhEsXwVQAzkjQ9MLuQqNjmemoLPZU
3rO1Uq19J37eYW6/YGhoXPx0hMYxXmmizAaQthJt7b+9aKqPO1DAngdCLRUmDtqf
oLuqH8RrTQuR7nRdMh5M3CE6v7M6DB87Pg7HVfzrq1DS7wi8ovaWFJNbNdhMcWLY
xcTH3uAJPw46IUaAZl+DDgG/cS9+piaf9HtgipjlMjinJPBkHRRRvuQ5lMLypHcV
Feixmr1mYkGkaMe+AEti6gj1iyQIpFS161JT2Zjuja37iy/p6/msUZuWeFrlYnkc
E51v0jMfExXUXl4R5SUTpERiHldbT9qOlFnA7YNbkgi12SaSChQMUZZrZc1KfceJ
86iIbmYEtVQ/W7GivHkELNgbrbYubVx2yuAl0SkJcqNusbKwoLpm+3IYqqwEVlKA
rGzSHc+NlSQ0sHAem5fTAttPxGWe/Ic8+SyofuxNRDMqQdu1sLzhFZrZbB/uUcUu
pi8X4+cVSS6dAWw3KoHn9ZoxdHmBCNnOrkZdgEVn9Hngu5iAEpM+zNpEciTqca1M
4BZH1pNkB5yfw2HNaYUNpQOkJ6xKUszuGRW0Db2c2y9xhE+gWBDV7ZeUzVZSHFXL
iiYwFwUQD9nbBid5WwcmFJkacgqMkPxHIqODJcezxRJBWGLzn6K8g8uH2440ZY2+
GrQpTfVfd9lcqM84C7ZDtorr+Ahzhkyb/SPJHdXw0vExLqJucV5ykYescSzgIO3j
4HSz+W3mtdvVCXhmN5e1VhZa3H8Op2wqdQyGSLQfD6Ick+G4n7sZfGo3XbepL1vO
wZBIQTeBcamTn36JvhQDRh3dXZgwwF/j4i/gZ8GQrzhBgkh3gdl2idCGklJngKFC
CLv6pi2jFMfbOqqCM09UUMJTTMoR8UY/jr4WyL7Fe3kH1Ip/hKAiswfdAkmer+bx
SFYXynFd9JF8kqUWSjmhL4HgHpGIRoCWyPsKGsvP1UJ3nksPaDHUki2t/xAoN6ub
Yuao+XO0pIvijmbOXMm14k1jMzoWGnTsBfYwZ5raZm+Lsth0YZu64EMYjuKFX2hb
dkJsAvODrBQqb6jdL1bfv9+xzzSdHv6FE7DkV7AmquzFH9kb4sBmnjBuLIMSwx19
+CQxlJeyQWa7kWAnXsHcU44DMRVNvZ9+M1zn0TeCzyiZGUfHL08cSr7sT8YEwtik
0WQBknMtxCND0yO0Nue4o5U1GxMOkYWEhlUa6J5vxTnMehShCTZwZmXhc0u8vU6i
MKfYOG21VMaGSkEsBKgVPCeeAlqKDMLapeicZxCmd+U/wnWGnttyACxDKjpRXQsM
ARCNjCrZk7r94EEeWuiampFR9wJo5reingxFO2o1Go8Z2z7j2cW5PC8H7g24vMEx
g5DKbx9rFDawwtiJRoESENtZ4IXeRxBD3mfO6VlJfjhwavf2nCmyYObbXkNWj2m+
zPaLiqb5IMonouNQM3Yzqy04gqnD4tg7+a5Z1iOZsIEWCkaYGSNvNkd6aomOZItE
jlLkj2PosjxyNUjpFrKTIPRQin12ZG6SVjGC1L/sgCQz9IgnyLBU5u3J6K3sGR6n
hhEMKe14GI2f4Y10q0y96M/Sh+2ADSmsBRU+riauDvEJTodDxtISuqAH9Sx/ZaVi
+T7jF2MCkLu0OgrNxPGsm5HT122PYRx24RnIqblwbKU2qjagwG4Bv41/y9NWG25i
tAPW6g1cqV6gsHaF1vYe4kEvhHwTMj6n+2jenSohnTox1Hv/jCEdfUxp1ZuTfNZH
CGZkMHj1Z2LPkErzF6Db+z3qRv/sT10Qgl0vT2h46+y0Vdllo9IIijRZE6vE4J80
02/aTrm0Zw42NKpqylGG46ep6e9AB13MgHeXB5E9Lzobg+sgBtiz5VBlxB7rId3/
YsAhE9Ylb6aU94HwTrShBbpue+3XHXM4oiw0NrBG6IIB8/2OQssRM3VFOaZA7tXH
n41GGP8jEHn+vo+kepGQzalTgjLeABFAkY2PpgCFGGTgg1b9ZvCjhM0U5Db2QLgW
4GTd68V4mFpwgXCA+TJ6js1iH4cMd/y6fTDY3XJqTO2XzW0RN/cq/HxJlKhRy4/M
XJTPgwTYEmvP/kHLD0DsUkhC1R5VZZCx8WSh0/glYLxUasxQWnikeH7tjsn1mzhi
A+UvdEb6bDT9jX46jmZcnJ19N0y7RdZb9RBHcZ9U3GJunQoCoHPgKkkH72wwWMXb
bam72vIX6kslYt62Tpj48nID6fc++C9xRn/PYGGAUA2kLUd4Jky3Zgj1DjuyNTuy
aymWxcG8f5Q8JelJ+IxGsIDCD22VdSszi3asq5NomvG7CaQBFWFCd1qco6yre7mp
0gAR0SR9Y1BsloPdPCnw2+5KhWafm+o5MW1zx6Tu4JbLuKQnF6Ogr+DcwAaPs1mw
N1c1OsTOSnGGQbFgqGxZp3LnoYknwahNged6Vbzt6mLrHOZW9PGRkBRQADYFIrti
nSO5I4WVHZ5aAhuQAZ14HQ2zYDnkInxeu2J/3XsCMLZNIYxUF1B961jbL9b/Kfqj
i4tjqCkanz0qEkEN201sXicw+3E7veXKZDmLyF9u1FqTqpdapYNScYfE7zQFrKiv
3vhHtMAQISHRu84dRzfnUpm2vDKnIlU3U7+9qV568uZhrV8qrtHadDigkWHUyjC7
HLM+lqxIholJD2kTR8JURfWzvRlnz55qd6sP3G4+Qt4nZ1gJq99lk/UqRG3NKYBc
CTNrE6Nyv2SrdVfaBamzbeib73oCWvahgbba1wf4J8cMSxlZ3v6jW8EapcELct5t
bgBXlDyJ6iq8pLly9T2olr/WhyPKfIhrAjtyABPB9Gds1sNerDFJ6Ow84s7xyo2l
gAqFgaYlARiX1m7x0dd+YzgtBNOqrCmUcZouvgIiig3qnOkxIsbiR9gkc6V8hDcG
rizJuee4E851j9ez6Ez7cwpkpjkzTeTaok1IoaJ4dap503HF/Er4BqoWUSoiXQsM
CGcsMt9b3HokhBE2FymmBKBRHBm8PPs+N/6WstDqOO1ktV+ZOauI2R7y6URMYqQX
mekwLIDlwaJXWObmu33hDdyQh49CIlSRBOgqxAoXSQVLbA2grJVbqfhjshLD/vl2
UtAVFlrOHgO7Ku3ig+Qb5QjguSjnzTHbiexY2QBWS9YAskOyEeEDKPKn9IftLliW
8/dmgimahWjmNivzm7VBzvu3U4ZEDCnrzaz+DVR4fndvE+7zyb9e+Rk8Y10aNyy8
BlZg+gId66aFqI1dQiYybKiFAfoOf9XzjsV+0yIbzsfQeEYjiP6mOLwfvJWVQ6cp
tXS2OCypJFWkeZqNIEDVstJNMNFOybkqlTOPso0bCLK3u9JG50w8xMNcDl01TUKc
bUxWkIqocexipt5J+cQJtLMy6Bkywwx9sZcUlzVpkEt4nvw04HV2cayfrzw624KT
XL0Xt/7OFG40AlsWBevrWpDqAETgLhMjIzPnSkr0kWHS5zh7Ys1DxhLuWD68BQXA
B8nBl/5s8QIuun/gYgW1+MHmrcJU4zeO/wfii3DcrwX4nu62nexJSyKDt9PhpKk9
HnPoXK/Jk/MR4AwEefbFG5KAgBgooWyHGb3ujs/Y+DOZyszU5fQpYqUrF2t1eZFK
VWw3L5jVSX47mW/rBv1BGKl5mlZFGw/esfxz7eAzOMZpl9Io7BMq2SqdMH3oV7V5
jsDaNzKHe51fJ8lxE3YHLHQVzJilBzcadtRdJJZluuzwSf/ETMlr2arwfSbZCfvq
QSf5STdRHMu8sz0hLBOzTYmGf/Td5TvIs5CXRWdnfxl3bZulByWq/ENYPQbkjQkc
sLLPWKKC+/zGQQaBZLUyhQY4KQexjX5lcZrEzvzdpl65uaTiZXfhlyMNyd3WOFHX
J8yvom39/rXNlNOU05e3C659LI3Tl0KBNKjE7L3rGyVIqiNoaH/25lm8zbc4KV2c
JOCxDvcNDmapLwhO52k7o+zhq9kzqrARxmQLacaf1PqOp9O3ifWghl0mfV0g+u01
nHYf8Kw1Qgb+QcixKePDPdteCS1/p4gyuUWxUWbOBVY88H6dLf0627eUM3HCXpf+
1PXZm0U6vq89kY4236w4+jap9urqHtdVrC2xKSuKC0xZ8BMsuficV9h1PrO6WlqB
qhhpGbJiy7oIQZ8xEvvKRiNqLn3aCQEokYMyU4m7bwWUwvUYTafYWxYdcZiap5MP
cFj/jk/ihe65HzosfN82UQtqkjZfY6bAanoD1/gVEtJL8U90D3IffiXV/rEBapqD
ytPzGhjoko2Smsfmp08mAK7ukG/q0TRA7b5HLFwFKDZhIGckNaPL7uImH0GJI43+
74N4cYly4FiqgsizB7iTQJ/GG7l0EoyeY9zsG3danNTY6BNnViEa21RaTMUQ+TsE
zfQDzgS6URvOkAD+TYaYZycREk1MUw5Vj6tut1IqmmDO5zJBMBxco5vKiv2hWP3z
sN32IO3OtD8R5hxcQjIZRSCxLG2D9OLhe6An003vlDBCZWPjCJ/DWfGmIQFG7LqC
mbsWemJ0rf2k/+I4BXeHFEPD875r0NJ6NSujLnQo1hy6bxYc4GlZxK49ZxNKourI
RpVZn2BkZmRIypYeiANf1f4Ctv00Li/+9kZbB2ut2GGKONwkcdIi3b3gv06XO8CY
mZMR+yqtiE15YZE6LjCG9a0gf2n/ZMHANJSMfnKQFhJanjugj7EJFNvMAvFYB+k0
YOeVXGHX9IugT+dKv0idYnnXYp0JrOGrP+qk2LF6tFny3TLuU20vg1aH+8VkF2zv
+zVD81DnfqLkRvyL0m2BlQleuSVzEEmvk9rFIr9MYjiM2eOvGLHhp7pfcL0BdZNE
1mRMxB2NvHDvhFM2kjCt2Z0jRB4FxSTEGGcbSI45GOIH+0y6K4iYBjOIUCt6awo8
KT8HlhFGodW4W3ejbEeX5n/d6Onol8QwkzFdleLjbqU8P/njVzhY5UcmidBawwGD
pFqLGPjV2NeIt8Thl4/Yk1vsTuWbyqTyK+Aupg29sAFWJgoyDPb3Pu6JpwvKkNwm
0f7iL8Af+dRMMXrzcAc09hwSIz7cBjWYC3jQgK6AZJu6IQLyWPiczoOsoINy4y3d
yVGijHPHreRSN2PDNpZHgrS8yLBspVIEznUtO10h40BdYGljJwRlUdaasQoA+EhS
kRIRmyD45CYNe+auMp17NtNt9ZdotQauXUjySNA9AzUFDk2/AEb89+Rzd7IhsNb4
Ej6aXG1+oY8+MiLrNAOfdFN6DoEXvrl2NmF7R2uMqRs58ze0v4w0SVVwPsGT7yGj
brBobSHuIpGiej+cGb0EftOMElzjDofVNfBywmSBILuEeNirNobqADMUT8oot7cO
XLp19yUDiVoJLXs/bHuSsGj68I12X0biVct0uMrOoYZAE03//OlVHGlpt8WqzDFB
d7V0WDePlDAhf1opvyWxwTUvJxd9iINIMgTuww9cF39KV5/842Mkkxswgjl6I8YH
JUghVMKCJ4RkCoo0pg1fNXmaNoOOslMh0JDjw2JGQ1M9/cb3pXVn5+2A8Lx9wsv1
/wCOPjK1mJL+gC8pikS1c1W6j+DTOr+ByQS7UnLt4gxVnhaeLWfJbmfhgYbwXoED
toP8T4TzGFuM9J01EXJG98xUtqsSc1b4pbTiV3TKwyX7a0LDkrQgiSrMzOvCBjxQ
zv4ZqQ6dbOewT+Q/5EgiIaCked3S6zjvjZ3liXEhG/lWtZoXuRJMfiiaWtkU+Jkd
ZTQbgC7TeGow+555VEx/9XS9+3TFo+QMYeMSJjCOwkLlxB1YcL96cJ4KaQMnsWpo
3AbePqCdZ/P9KI52Qbri9XhedI5gPQT9AqB+sbT+heavXAaG41MHZngW1NqE+xd1
h2gTJX0/dDsFgo2yvhdZJ/6kbm5J1d9FqNEFcg4pBzgOjrcJjA44H2XG07vynZlY
cLXZch1KlHM1On6ZsQs0IBZijpr0igh+d98Nzs+ZUb9W6QJ1BUtLD6UdJZ8TuCyS
bXOCdRqmRWncPSBE02dYi4v8gpvzNDvubzKp7PGcpFWNeHDk06eMlvKYpg0JJPH7
/J2axS4U8MU4Q0sjMBtPRyZb4hFMFafi1io+qOPJoqFr1E9VYLeCIRJrxiBL+exT
B4F2YCQnPeRcOFhZ1Xg3zEOyvcceatLUbcLJoc7DUxsaAvWJnMZoaYhVuhxmnpdZ
2XNCODXPbC1E9dhb5/n9gBKi8pRUXQ+XE9tP3mK3AprS77W2mBza0FDWGSawgZyu
tvzy654DyyEePf7XsIGQfp9WZ7U+MDh9NrJiKtpl4doH57iDGbKBA0Va3d6gym95
pnQ5s0S3lG/cpZdmZUSnaOhymaKbyF1E7kuggD+4TM3I9ehbNUUx+28JbeoeoFWl
s/VQEgZZ3t+gxARQV+e7NeTUZR8L8CnDLcpPYY2bHy5rMXNsfh0nae84TIX7DwA+
pukLo+HO35F1h5JoEclqzB0LwTZLINX/GyRe7Vg+B8fK1XJm8yTLQZvOQOXldXoi
ZIgvH+u/RLE7pU6Q6xlfD1WJeya9ubXjwl58N4xlumkTCTjC05AEIJUybJUSI+Eq
J3ymZkoSUiDxVRDgf4L2peDbhveO2n4kwGxHcpfKs674CjNS5UAnRANwTU48UE9E
VrrRACzjtrrKYJZ0lJtb/26sr7EvCewENrvrm26ZpmCIuT5DUGArLLMkEmfsY1RX
a4d4Olwogg7U6++OAciNgxGbBHtqUA5h6Zs3cb56IypJodcf3hpEQoB7hNYJ1Xz7
u6+wtO3VZ/KolcBUGTzZ+DmKeof2MJuBiFVqjEQ9ImSJiqnrVl0Mpg1CsbRCcmH8
TX0ZToNOxQaVp2XUAFXT+7InRrWc2nIBjUDow5m/T072nTGSgMCUCobW5uDjWyC2
yTwNSsMpkWUpEaDw/YzrCuq2XLh42PD2g1ypdYrqgX3Ukj9VzgiaTRggesRv9cL5
YbDpzFQYmIXjJofu4/bfDLX2x4nT5sm8ikbZ+iTeuayEALTRi/tlux8TPrRzlyUf
KU0v0TbMJtvADWHU981NQd4bLJhxJjxXrQrDaHD7/KuYiyDsCvIh8bI0QkBX2K/X
A87+nWHSF4c00YPVW+h9yobhGydpygCl/WVRO9uNuhACKAkfaPjyfoh3ePXsVhtH
99zwWxsxB0h88NZ7/8jT94J6xdnU34Q9dk+/rx4HfaKeDoTapK5Ay+NtYQ9qUtEe
NROV/CwLZFq5Q61KrlcgcetVp6CODq0xIshzrlxw6NG3J6B9je9kq7MDWpvimUgA
u+At/RMFC17yrRrIx6T9peI6cCr95gK1kbvOa2YIZwFuyLpyu/tY5PSEhB0Ttmvk
PG7FjxVsYzWeORFsdu9kbO3vHLFe/eNGsl1WRXFHE0gPlx9JkUim0TEkwBexzocu
zqKrbQLppy8gcRhoMXBYMV7fKlW1la40VeXxnkNWLlb7LxQRODdecmjRx5d7jZV5
bpfhczakqqF6TIX2ceKJKKwJfalMySoby6BqoShlKWBssFC9O0sMw4rbjjx4NKhA
KXHBDABpFoRX0rCxDsk0heAOTazq9ES8C9RFTl148a0XefA6dnSyyisB2N5/NSRh
Q7fxa55ngkjv8uUPQxkxUKS/x1MY6JaArsMJlzHREumFmMHT7d2izlE1dNEgbylm
7JP4zr5GHDjTGlhAOwGuiHiny7dBER38Wvv2I15tpfTK4IMz/0lKufD6YPe24foG
te1cevXSZuemG/NpaVStFTheqmrSGafXuoOWRN8HvuWLjdgNi4h78zKLExlFLiYq
7dE0RRJQQsIBMfwhCLHWmSpLqU5r2DOQ8+Obv+8bAf2ax/G1d0re1bHEXDl8jWiQ
wAHAUkOAZ85XcFjizxNs+DOWqXAkZ/bOJdhteY3c6vpx57V2JruiiyIuW5b6Kkkz
ArunVB66m7s8coI4kPmyw1ldEfgGSWTYdVjvmAKwyeP07M4sTrc1RIbiExEux8A5
vaToULmSbkFR8ENbD7t5y7YczUXVtiKMDcx/7vNzb8U5ATIXf3NbOP3fAa1TgpJc
AiGzmO1HxyzbMjECnJnrtGJDJAwh0eQETx31b7b5OLmXij4Mt7jtlxI0kAKqJLMS
9KehpGQJ7KdubWQghs3NW504LNatQ/4dp3TmarH7f/i+AGScGgIpEtFU7mTB52tg
pfi9wb6/+UKmfFAr309xbP70jA7yGlS20dviS6WS4n7573GEndJaakvuxexuHJKl
WoaVQhhxmDzO6Lp6RRx2yi4HyKY7bP8O4bhpNSIYgsi8pDA69Zv7UlO1/qqOZP9U
Bsggbrg8iPd6Wlr5nrMzsboMuxxr2c2ldnM7D/reISX25ZO5RpzSWNLNPEYLlC3Q
+6zvOmdTpqb3KDOZPD9t4xNo4jQBuwfxfqX/e/odVu+twhuJ9kHcAFge6sjMmRuM
g06XNNbGXz/rvbsnSeTpCjedOXlBqICtMY4qPEWHoqv53yn0EU1jxg1dkd3xDzqB
dUotjCxP9f4bJYWtKSp9/kaCEH37bUKnY5es2wzkZQsvjIkghJDP2W4p0Mh+EBqi
Lbob4oxKdM/RyrPGAJ5WdoEk7dT8SO3FwaFVy3/rKnpj6h1reCL/3ickwSOFycfI
ncxR/32A00ZLNe0FLijpnNcQIezyKx9eZVVAAFPBHL3faryiCIwPJUDfEb9oOVUS
9I+7l9sTKRD5LWbjYWnxNSBcp0QI79WVrGMiZkCsVj1/WWrU0xyiry9xneArdlI/
5i4xibTGIWTZ6z4GVEOSqM7jvhObbL251zfI9dYFdeKNxVpnlu5MAvw0mtHZbX4/
0vPukjStAXXboHEMwwf2yheiRs/QUDRfYnmJgPBfaiBHLSBmtLQUAFMbUKHvPJgy
g4dVsT3odTrR3b0QK0XSuQlVnE/XYmW/QmWCVcYYxyNUFKFMmw9WOIU7twToMKCQ
qG5JyOb/3Z0OcaHH7NXyxxB97DArT/ULWoff4zAMRvgSqvk+ZOQkDjDn7w21VGiJ
L7y4PStu2FMgBDgczcqevL8OTqqbvycORVH0HZAfP6KLqyK8fsDBi3f40cL4j8p3
ix/74jDWd9hWw6hfq1DvvyLUxUJF+PcBNggZpdW/43Pi9diBgy6QW0NI943Czxyg
E9C+FmbgE42HOXKfrc/C56Xk3ZLlkUw9XYOql5HQJkAFVk0/j7xPNDkpgQatwvGc
UGWqytpGbkmB46i5PFFlVGI54c4mAqNgQSd3fyL3hmCL1rWUlVCpc7QLC9GdiDxW
XayZ+AaS+sNa2dRJTrq58546AxoAeof+2+VRwgUc9wgIbjyyXGrvAa1sJySlCQ2d
VBYf4PQ97Ghn3ZqvpThzmAjWEPSNCTAj2ZK0kjMTp0N6HRjcsFOgH1bcIMA0EDXJ
AZE8iy3HOBdL8YAz0xQ/HBfUkC6/LrFV6fUtItMUOdCg7tS2pVtYhtMnpcyfee2e
nMc77X+UDkb3h24cCqcnJbDik680z/t/EmdHa8PIqKDhpQ4oUyYfpiOOzKRGDj7F
tT/X7+dUjLF+la/ZkAmX8PzXUnCMBUP4x3qRMx3dMXEGemMv5uYJ/kKA7fJntg6R
5kE2iDNVLlFVepPkWr2fHPuQ+QIEnAjTx9qBfj8TqK+/sdlHVSgi8qM1iKowTG9J
dQanK7ZYvk/lzNqsN2yP49IIThQcjb589W6Ql18foco75svJD4XHh3reMg407hph
LBy+8A66d/usSBQ9PC1PnqGwRrbmSGxKgnBxCjE5fGwiUSVVbD5cSnWj4JxueiiO
2yI7w5FJosZTKgoKswXJKtJMp8oS4wmUNKx0GtH/VyerACQ3EGfJ2X9RudaNhbEJ
aaGI/yysvQsxzh9yWdw7EGOYY6XllXQX2sxxFd/XLNN9xRZjnMySu5Jnscl5SOpE
e9BtM/zZIT+bWLg2eIdgtJhp7Q9sN8xh+n8wiySZNYbUbSoEE9o4/IU5GH5NOJPw
wxUtZ6r69XGr55Pq9uv/U5OfYaMOCD14g9M9vJScDMXbE2JdGFmhnLLPjQs6N9d1
1HergAc3NBUOrsyKVrJ2oOz16y/EN2bR/D4Dy00I1Zdafmm2sf9tR8HeAMfPi+oC
teSRJHTsf9AZ5o8b37Sfbt7qKpzTJ+JT4Og4cLUQ8Z8WYFbqnxMJFtu3LPHrvMHD
6ULTACHBCdaNXnPV7luJQ21lvTSEHNwNumBcXbnED1yddRvt8JWvMv2cScgaDLfh
wkZWnE6+SrQP/YernYRQW7+TZ+8iQwAb/LHxge6Kp4j21JD/z6NXU8eqpeQeyqOV
L4boxhd///PS0SCM8ZQgPoP3n+CMYm/dsKGwwQf6sGF3gjBi74yewRToff4mZKQh
BdaxPl5gkslYSyvvO1cHQYqGc7Yg0dvHhjzN5TqLpZ/nIECDIQt2G/4k/Vm1xDug
zlYsrCatyBTgfsNvG0vN/0oYr2bpas6Fbq+FIJKbd+AVynfFrZLh56EBhBghP3Yo
s/VdS4wOLw15VDpyKZzvmq6fOulr60MZAlBTqz4w9fiml8qcZvOEzT0fIH5goaar
m+pAm514ccIH9ranCUFRXsbs27+SXsM3b6TgB41nGQ1OlcMOkYfzCKp6S9SY4nvq
6AES7/TQBCTlsrgtoGeb+funKLdsa7ra1om72mQ5++/NRRIQ/HbnAQThtnGc9LRg
ihbIf1XxcLvkJVcQnga/aj/IyK1ktHteZ+KT04Zv2/LRnthRKfGZRVmsos0cQjnW
cEiXacFQSzRDXmsBvdan5Zrngwn6+MbvpJt04B6EHuLcuQ2S0VRAGTQus7JGz4G4
+707E9R33FWKbZh1vCjoRaSTH69pHXxCgyLYICNrG14xEdkC1xQwH6i7dBrGb3zl
O1bx9HtLFJ9tvPbkpj9iDe/gXD9ll59WBcQLexGOEdIB5MUWJlxipBO3Iu3yV3wu
cbFA37i82Gqph3d7sJVaSMAIh9xgB67mzeHjeMBbeVNiFfQHMXVoLx3PuWjY7IyF
mtCeIVFonEh3uLbWep9Cyu1oCwB/7mcdYWwxURa5VhinyMzeraAXLTda4NdrXxkW
h16/h4xH0cTnTolFw56N7DEOjgNHU/VSxD28lSBXDWADYRdkPGF42yTtCOKQkGrL
xy8h1ODXmCzGMR9PJHwKzeVLPE9ftastbzh/1ToUggP99CC8dR3NIjthBBK05Fwt
wSroqZ+VlgOz9/u7sn850O6gUHcUNWL8Si90jUxe77rVTqZWS3AvRK5666da5iVx
udtFLQofYuvOKK6tGR/r68OnvD3h8KYnYrcAlly6BBJPw1XStdfOSPj0JNI/SXCJ
YAtqLmBNY3XiTbqJ3bfAiMlpiOg2eWbYJoFWEHVHK+BEb08BNbDONSb8Yd9iUHcD
vc1vAOGIp2CZifYQBRT83Q/1dkdXPypIyWpXximNxDYIIDwlw0ofI/jDabPHhI0j
L1Fk4OHvH3vnu/1WSfMbXgYTFn5ZtEtWc68Kyz1S1jGrSO+h07BNaW7hwj3dgWyw
9FwsPC/Z5eHKmV+gK+HsWjFnoCS+mus6WHOjmk12JAqxr1mpJ0/ixninF8p99rQw
IGGl6YHuia++Z3fKRg3lRPMGS3H/LNBCiWlXxB/v8FKy2IMnCjzhd6UTIJyYctc5
cJG2A12BZMlLRH+XCf+cOAtNScoeRRTLBBF+TXIRs68ZuFt8Oih8gsG/RqFUvMxs
1jbS6WxAzlNtkcBVTCmapLWmrKA7RnI8573vbfr5Xz7rswT6k1Ye3T7MDS/NE09W
CYr80gTTe3Hm0r5xDW9ibRZzhioq7uytHjp014ZRA1ow0OnEDaORPFoLgoGFgqNY
KfqhRJBP42muj2re5qormECQRipWoFrjEje/3BmZIJj65QtlADUIO9aIQ/xVpsRc
7kjLig8TOoQP2m/7xbwep6IT/lLWEyJixQ1UpVrzHUEX/jGevGET5OpYpbOw02QU
3P1weLLDprJUP0CfpjrkGUo2A+BrU/QBCZvN8D3ia1xAJLQzS0BXFwDb+R5VbwQZ
3LlJMHiymB50uZgREPiI4azB8qcEiDRWOR5lI44IpOnjaJhW8lW2f+wxq3iw5idu
ZqYVBrKbtwxb/hSqUD0TfYp03fUaeK1im8OBC+cc0dbjg3kyaAPAVZdG7QpVkGVz
s4X2NVcJxbDZb7N1KwIZgEV0B0qFm3RiFY/RWwimDAwy3NHxwAUs8idRK5vnbCWd
vcmkX3ng5z1KpTdc1oTD5CQzN2rOBnaDwoY1YLTqfHWtMUC82arZpPVcjscM1py7
/zkK2fmlIjgUCeH1JSqgccr9zcl5ocsLXC9oKamSX0yw44TMVohf1v99b6kv+odC
bjtBWuHYsZbWtqj70cQquBvI6+Err3LCLFRCzInao0usJmziEWuclWyJ9R5Mg9WF
YpzcvNq38mz7xjomwSITe2blX631A2hGFRh4RHs94zla8MzdifToHVqPY2bO5C+P
+AGo6d7eTZfVnmrE5HmwEhTuPKhSN2hU5V0Kz8xh0R9N96DOv09e4Ez/9ryIvjAa
KyBBuF0O4ft1OCJEho1+qqdqast5n5jgLyORFr5JvSQgetSr7gR2GVVALraVmcRH
gbaUjp7eoB4eRgrfPGiSg15MguyD+UsYb+xJ8nGwwcp0Nts6117ZONrDnEXzj+NO
1nidfPU5b5/sFoIbcRBXCSWgelrH01HQjjV8f2tOiEey8xiHEpqzr/CUKBZZl/OU
+yLPyvJUK1NC7nCUFYQ6Qy51tcgaY/iGRNPbhAaegsU8UjNQMbLt6LWXmpwMITh/
G+tCK6vK/kUS733jKmpK7JZ16toxUab+oCXbrUaoz6JpqqbGuiZ0wtIEm1GgCE5X
qUvcHYid0RRgDjQQI+y/M5ylPGWiRSF36yAJRSZAFGuArgQZfbXVdNv59JpYVsNU
l7MshDcFM/LFhSfAUPeSddOCavDZ6gvqyY8XshILT9IjFCAfqJQ+dxm1pnW3fL06
OdkJ6LmXx2VqvzpabZH1FX1QWfiBdo1MngMwHDJDw4Ra/uJBc0tmo23+qu3s1OaY
mfy7Z/qPV834CGQ57BXRCunZ08rsxZgFBqQM5UBS3KurOrRMNPZnul9hiP66aFdh
z7CgrAOqkzfXX3qfHFUVGSTMKh0E8/63lSYKXl5Wjyg91Fctr4Fuo/p6yAGabS/h
1GQzinklFl4QgJA8RzCKFcPpYZTeldQTrNf6BKWNOy1qi0MSYlbFgRDr9y+CMsl5
l8kiBi09oohMwyhjZbHQ/tdWuhlkjVJ0H/vQhLMmUqKp3wQJzXQNA6jn4CdliVWk
zlYYStgc/X2QJUjjryI0WS7dp8uKhZSMmK70aPVDkgb8FhnjJ1wN9T4ELKWG6uUI
Gbj33bK8EZp1hPMI89T1DZZO5JguJN5WoytKFgSXK1v4HD3ys6dpgMqLEcXdZsxM
ppNOCwiW9YWCh0KelclyWWwYMoiLrDZg0fLMRBB/MjQ2Xzx1UAdKRqEuDCVA+jQH
rLAlSKC+pZ0TGdZFy99YovCFtgoipg3PEPH0mSRbBnZJNrishM54AIZcU3j3o2DM
phCOUbIkWSdj3JNBGnWw/tTXza9tnVwMc7DqjvrZ8oHwEJEzIkKy9QgAPG98vvMX
WcUxAnVDGUukW5USGy0UMtIbjGH1VPYLTYTVQNPHJriOkDBaxZKc0D9+WBSueP6/
fxopvR9BxnCgN4y4adbwk5qz/YMEaaFT2+aj9p4GSHKqGmzc1kd8HJM7/MX4rJMO
9w/nGXwj1wptO20bcxTxhcOMsJ30TJCqYpo5x0YfuAMGfyXUO2/IjCwR/c4+zeVP
8+9/vnVshAjUaZJ40ihUROdDZEm8sRSLfxc+/6Yc7iYqPoL++3Jr73eVi7NlfbOs
vWsarF7Zb74A/uNQI+921gaNQE0MGKI7YQklUEq6GJMAmcde/zOikQK9M4czvH3c
LrDbIbU5prYa0N1fyxWcoSMcKn3j9Jv9w7+nTC/sQK8y/V5IlkNGatop/FRtpvwv
+P6uWXy1eq2rFyYEcSB4iOVnZnQW11xHHdnGTDKuGHZBdgSAcbWyBB6l3KTpMhD/
tK1A3tVe13sjJs8nHlgNjCOvdcDt8OXCra9eMjW1NNTda1R/LzXWEzUMgEPY2BBZ
UOAIs5tde1KcPy25pT2/Gu3Coh+9v1Pnqq41h8t7Fi38XPxhLKgKgJXOYZCjzsKz
mgwt+HiXjv8gekbIQ5FF2BLqrJrJ4Q3iInF1SCHUbzatccovDA4FUsAfV9KQVvDx
yVel0KH0sVO8+7KsDYhNaV++g2IiHAUePEFyed34ZVuhNe1upLktO2pfPk0aAMkk
CprOL3ulxzi1VtslVQhiR2KfDz6W4UCowIXl9Sz4r/UPncOJzzSGvepHpAMiTLpy
HOvDWgi593SMkOZ8YFpU/pvLSyPj8L7p5NTMvHSk2ibRn8M4dosMg+wvgv7454dc
etaWTIKhbiVwD4D9CRSn6aB/iULv5XZZLNZG0L59pr2bi9VlaV9R70t/Ji+wvxkr
cPMAicESuz4Hs3qXTWNq0GC3mIM1jzhpgfvp0gx1SlpBZf+nCIc6ZgZ6ld/ixTcN
6qitiFgBVHwOqrI87qWA5UrUV8azn61texN5fPfKl3JxQZDhFe9y5mfU8Gu/OkkP
jc/fCb1Vo6ftO5u3Ee21yv2fmQfXa1bGO6DUT7P+rcZO+aLi82aN0cqj67qmTUpF
CkG7BHScF5whoL9QVxEXGkhoe82sr3l8q61jQe5+5Fn8n+M7ebUUBNT2W9rFq9Uv
MSDu3Qs5EIlYEyuyrNzgFaqNumCz4IqP7guO9G+uLu/mSCT/PCjDyGeYcjNIExX5
1t+Vqa6IkgmQPPJE9d2x4MLGbr8MnWlL4vTL6mCdCImEvjZ9K18fB07B8+flUOGd
k87MR6Q3K5LfZgGaPg84zDR/7CNJ5uFUBW5PnzIONKXrl5FxcDh6g0dWNVDulu3m
LD24vF98TfSqR9eyrGZCeu7gMC+KDCCcZXKv77a8GY9hGQGKYW4NcVQdelK5Cqg1
4yEE8HsBPxkJmrWlCO9MFOYNslGXWiWJfR2gCNndoWeDNhSkpYHx/3btL2nhYTol
L6ToWrOxKOBHphp9Ra+tPahelsJZN+vFjEe3fEburnZVph5CgVFC26GrVwOqDVKI
YPHHkUYYQXISdTnAwb/PuHeoJy5AHAjUiLVXhiqwcCusHBredl3sMCADZucB3gqg
+GzbB1UhUhFKKv6nTYog90CIsaY/ihJrg5Foa8bFHuZv40HsoZ2EYyCCXNQhWAM9
ucX69o1m/xoYxJRRkabMiTy7uCudBDdhuWBI8WDF7/EKXb5IC3aooDz3yvnRZ7Yj
s+aqZ+j6EV5mrhUxrQFe195vL4cPwMmbHCJt8S+LOKgLSspj98msIlouQVsufXFf
G1zPmbJ9PEyjDyeasycrcZDuYeHeZ/vvz8iSkKnsODmfA0LO+o2zLWhRXh76dTDH
/N6nfC3JjspDWCmmB0ZQ2LgW8Otc7sRud0C5pwg+pwOPwlJTq/O+8SN3gC4L2Tsk
mf7QPqJhVQoqbKC6EEkQd5BadmKHbqLVLAm7edQFDlvpTupocAF8dK0OLPkCzU5x
veiIOzyEvFMdd/ZzXFxfekhk3gjmGysPVF2EZvmkpowiMFkl6Iul3oxM/Vq9odr1
jKyv2H/PZ03VZCZJj1FONgjd5IZ+0dr1ZEhE+IJSNTzp17NmGBHA6fLONkM9Mcfk
OB2ATGoOM+G2OrXQJYvV5QOHSweIx1uX7T8XqE8m12EhU8tzAVMRezc9vbtOyHwN
Ozxz76OzUDYiI6bNWM8usfM70uMSfvtwigxivlLK21nIwKh6MPlyYw605ii5najc
DTWwUU/LMLT3rsg94BDQ1WzKzu6TXbk8CDrSFqkrc9ysc4XGVkt1AJDOQK6Moxtc
71rh+hnj+d/vibnCbPELrP1tsfWZPAZtrO2/1+WasLKUbRXY3O+8oNPzmdjYry9r
u8Hsp2ZDKP8uy8aeBdtnDb1/z+GP4D0d31/NK8eqQsi6+5AjAxKlqbNZhY3y6uer
vbs5KLX7mkrpPzJ96757LTvt0dn5im3rz639C67nSl653HE3bILkXdP/Q0K2qR3C
sknaNsZsbjGJ6eWuJM8Gp8BwKYHlsOCdGnJtP62cs6JaIuXYss1bph85rMwTTJmU
TWrblB7dqyh0M1anZAP8JtlndODpilTilORs4uItaA6S4n5HYT6Y0M3a7A9n5bFv
HRpsql5Uid4RJJqzUb/1TqOMnODm/EXN+Wf61aHh4KxDWmqupwdumHjpBoq5tl7s
dRupGlv6xehS3UC5u7JqwXSdsKt+Tk4ruTrqdn05ApLOKecMg50w+/RmLcBUnqyZ
OHs/hohT28XpP9/bjrlnIZYR//bNL+Vgeqd8fZqoGv7y6R4vFDHazTDNgB9DymE8
JXu4l0fBLjfo79xqkvdCAk8qoHoRCs2vJJG7IztplaZXxShb4+9R2MSg4UdGlfkP
+VxP/+ZUpzpenuMY2xNTlqRza6SxDY2vJbufZ9/XfYj7ROjgFcOoj7P24U9WWtAk
Lk374z0Gr5dxfflffWuFqk7vQOsRssjd0phUYEGNoS/qtWSWwSJ+PatNAHLwcsyD
LIFx1Il6lz9mGdAhJA62hPvAzGEWi/7s0d75TBMmDYBRGoKONFMFdH9hTBXDLX+T
WQEHSvrhGeG9u9xh/EN8sli+hd2pFjZzDE0AYYjQHA6tNdnFu+YWznhi+8q3NEMp
rJozLBpqvB/yIkoSuPu4APjpTRGeWqXJw9STKgmEdLvYC57lNmZ36AWBYAh1cQqB
85OzxKWvK6nFkAUrZoNyXCaM69484nbQaIBb7m8hC3lpXC8YhNXVTpdtM+u8k91g
9ciEA2qhhWgFLNUIY2Zcl2Sfj6cTw3DTeV8FTm9Ri4fChqRN+jz4uhPVzukhvAa0
A/ixZqhMG2h0yY4njFpukVSF7r1z6uLkHtyrGivuJ7nrNTsS06tr1LL1BU/P8iqR
dtrR0XptrxRloBjnRVfI7EzWYzK06pPvXlU8zYSyDpX3eAZVL068FoLSOMOEWuyW
9ryLtyyDl1PNTSeD2yBitpXxjNERjTbJdElxeoQvzQo7TD3244ADkNnBuSujrkZz
Wrx3t2mAW4SSbVOm9dx97RMFxeErTIso9mr8p1O/dXxCk2QlHxCPk3jKoAINxuxq
Psmcu5SH3M5KasviK2PnsiZZ8pOaV2sY+3ntdVVUr1S/J26r/wnTmtFHYK3p0YT1
pRclPHFJPi+ShvQBjveb/5zgV4fxKdpoLJONu5JhPq46DqdGgleKIeKhLEDBCkmA
EJYUL1isNiS5t9k4t/b+vaypUEoyq4wY7lplt+kvkQmnTK4kkHa6lkaGz7oE1EWG
0aHDRasfwKIh8FyqkyQGtZCu51pvVN5tSRMYQi8/kLGJtjH6Fwp3Mva0HgoxKmjU
0/TxRmZW+4VTLEdlPZO4nLPOA/RIpPnuzQqQvOqgGTjxW8leOuf+MFNXPuEgKTFB
v3fV1tc4xq27HLR7TX69w+IlcTd9jpVVmrqyiLIdKYBPWCNN71EX6FF9/E/iVQ17
S6aSDgN6zcJW51A1t35MTcKGa3+6tStOjxfqrXKlkkp3iM6LtIaSDBH8ZFKk9LX3
mh/B7THEzGeEBP7jfP63vqjnyyUiAxNlwZ/s9wDN0PlyGgUbFUJkVAF1doXd5EPe
dp/TG93OXd7GPAX5s3z5jTfeA+RbYF8rykuO5CUutW0T4rIrrBIkgD6ufR8h8tcL
nLBS6TMo/IsypT5F3zWFu5O/sPcyxJR+wIeVydvKSzBormubLq8Ev6Nwgqihdjou
L3E18SUOgWUiIqPOFlCr1A4Xs1lwyImwwZ7g1+Dh4LUre6mKi4+BW7F+S/4rSTbE
9Xqm7XIHRE6W6PkOTjt4bedwxwafqYswO2jNsG00OG8Mfpkpwy8Wa2eoUonsdVEI
fHnlzcjmIZ3+8YBqHKRw78UPfd1SJtNbwq6I1bf9GNyXORffwbn25qUMsfZRrv15
JRcHOio7aOkVvlZ9+zvlqwvnGA+G/LH8oY0T1QkslBAjDeSFkbjhpsf9R56OaLGi
AUSo5azZY11/B9AXAFYfXnxPZW0JhiZcsHn+Vl+i+ZHGKV7EUj6ydOBcsU68hH+N
UayXPrtYowdOaEiKiZ3OavSFL1mykFaAr6iOCb/CXzIbhzs2q7MMZi4XVxwVUZsg
Zdp7AGqlBJesIP0T45ktWirOgULx8tHL5iUEhXcw9OOAWFJ4SNXRNEK1RwQc+SB7
xTf/3zICHTgGQuQn8U8R+Lo4aovZne34j8UW0DTo/YFvb0E7DOE8iTRStQw+6tYZ
2H3OKZ/MrOvfGN3VX9I4AB79rfjuBWTsimkcGB5Z5dsPLE/GUfDzQsQ9RT44KGek
tG5FAeBG4oj3x9cGz7Fad3T2h1Sbzd9fx4/PCRXCj5bUNPk+J4wkmS6bHPx7xNrd
+WTfSxeGCJv89WdToocwUHHRsLNICjUDd/OCT6N9RX9ZxhzKam3j6ImOh5q0EQtF
ZMyD4fQ/LloM31jpRBxX5uIw6Qrm40W03kEUcA/0cBcK+3nRuKpx6pG+jUhJIzKR
Kbl7nXf7C04QQnGbtMS7uvUSETlPs0f7JOLukoWSg0L3l1vdotJdJVlbwkcUO+YE
jaI3CDKToebzwbH5bBOunfi4n4U6sbI6y15VyGTz4w0SOndw3IyQSDQq3PqtFmUR
iBQCrC5VebGje72My0kBjFL32b4e+6g4IRODD+/C7lqAS7ZXg7NOd8mk1P5Og4d/
Eg6aV/Me6ze3bFb3GN4GMH1yMkTsdJ+pWZnNqopCB59Gb6RR6zLgvKeq4OyU093u
rwQeM26UmwDiEdoHKqC0HXax4yCGYNrepyJForg7fVyb32LU11TV2PwG0bwzZFFt
iI2pBlfirkyVfUqR6o6md55vQl6/tleUhhZYfbN6ePu6XaglfE2HvcKwB7LYS/Eu
VqkATfHWvFNq8pOnCFWJQckFxU/SsdZAb+0LBEwxRo2nHU0oYkREYzyPAVnLAR9z
MkMMLZrRRQO6prqTpzgo0RBVAQe/YU9e1WqcELTeunIhZrpAg82iYPiMx9FC0iKR
G50/Y68WLRCBQEQHQhgZSu//Icgqj/3j9q1thR3LhAU4W8aYBhuRYzaHG45PxgcZ
1eqBHdrDiY3SlQqnHqU2utvF2YwY5gX37DoLq7aBj/Lb12zGmF+aD/QKMHcoEckB
C94BjxT16dgwhDMda3F1G64knB4/YMQgUxMgvZlXKHdchB1zh+VJvuTFev7pYNkU
H2EBJc/0FYTI3ghwyF0WcVPFbm8Q8XyZnjSusl6ZmSUThzT5FLfxKx9/NzbvWWsL
F73Y49sUxTVCnSCZWO2hO+amkFsYYzOESrolSxcL+plLiI+uQG9dLW9HV4pywbdj
p9cv8GhTXZDOX97zujQjfZ/PjWzASx4Sog6nJlaBXvBQUX9GlFS5UtFqsuMod5Ad
4Z6IKHDaSs0HJcM1NxQYwwbj8Ekw1h5uHykRsPe3rvBmofQ3KTjgYeq+9o8pZWEC
VdEI07eim2nnnjRk7VaHzUJeaee8m5sgVqcQpPze+LOinUKsZjtLfFlbNDgZ+mOk
lqOqawnIMZ38PZIyJjUWsf2ppGXHkJr9lXtnXAm9od/NpIjjBUe+sx5SZhdpmfaB
bJf4OKtjtWCeTqhaCotdYXkigOtUwlEk+JQ8IeFVrfWHkUp0ZGSADq3PLg0tSp5v
EDvC/e+DvnP+AsL+yZMd1cplwr7E7lMZ8jzskSU6hkWWr8AJ/gl3D1l6XoJLrNz1
7RKR/lHAlC6dUAQRMxV0ABqauDw22YPlLkF59p17AprUVLcwqL8v6B843KgEHRgv
9GOX4ZA73TP1FIyWd+8W+vbY0exOfI6OEZgBcnLSIzVU47DRVTCJzo1EFLUxPcuA
Yf8hhPQ9S4ppzpEIYedskfTi6HaskaSMCSfm8UkmObC10wpRnFzkNfvWBj/JPTMR
15fuvNAWmNjd3imvmf2Okyd+VNiHYQv8+gfmgOGbSiimnZ3Kf7tN2mx0tjjBtk49
YKgq4xQl3V5CsuGBbnZhSmpGJ5D3wRSQz9qqqNwmJq0b+cPIw1g/1g9iSOVudfx3
aWOfh8Dd0Jhp9p6O/YSwR8brmZ7reZWUNhLE4oLZxTqvQ0tCgRK5O8+do4UOKwWa
hsC3gZhqIWGDnodkvRrpxud4F/AS2gYs2J5PeUYbPoCCGrHAwlwoSfo7yIUG7wGZ
uwjNdEseRNX6SJdUGdIkMJQ+5rGs0uVV13qx4GFbwczjaiL5DwUPnjdALhf4sb13
VZPLUmt86noKJr1cmSo4fDCD//22HGf075ez7O4/nCutWdtPpgUGzCaQKoAU9u7K
NXIubZySW+c0ttg80K1U0VarFh4wr8ekOOrgINqAIu/xkjE/XdomxPJShDCE/8vQ
T3fivXhYU6NhRraPjDW7PF31jyxcI4hpBRvlyEaOPm22lTOC5DH7eYyrdisesOrs
vT4z3LKkSm8B87nLaDp2PAutiz/ZKwSM/ISvSzURHJKnvpc3cAK/9T88waVnhVBI
/KmXW/wJxWzJv/rnnknq22jzEUMYUbnCKTKD6tlfEgsssdngcwMq6iiu8NpUc0fs
eScWVnfpQwuMeLGhQN+xvjnmMzIiYYueN9DhRON4lRHOXQYgd6RoTgZRniNjy4I1
JoooOIJ2kaaSjXWlNmKahBwSifQPKuOQam4zuknBNCXCGyVmro/FiJI/8MsXd7uU
fm7+eGapnO9Jdcb9dnv0h6LscME3HeyzTtOW8YUt1oLqVJfPWXdjq02lzHb4Y48g
wqLquMMgHeyxQEq5n4FJWi8UQrABGzQoxsWQLouHAazsO2vLySjUej7DCbrga/2X
UpirCmJoR/hPlreFLL/TKYIyHMEbkdNTV+pIwcVrwzW8A2rejY1TcOCooFt8q54+
nwCmKXeZBVQ6gc5dE6LSO5eT4r3CVESb5aJ1MgwRRB7vRjPKPV9LuldvgJtM1xym
lz+n7Wi2RxHko1OPtFrVz+vBaU4Q1Urig45Z4bPg/iFjNhWqpMFr2UezyqwyHTg8
hymGVhV3aMCBB7GfRTao/diRZFSQ4KsOkkXuNhFTD7MvJqiBtIEtmhFaM34IbMbM
fF4kiFmf0bmUfikkMYMK+E5JTfJnN+1sx2eCamQzeoDQw7BAxjkPFshDyIEOuuCL
uZMcG0MWJdHq6z0M+XBmk5S7Xip9bj5GrA8LauyVnWbePmVj6jFt3yt8pkz/I81F
cFZXeUGozh8Em1BwuHTpBfcANbkc1mrGl4ufVw2Kq28sYnL20m/kJsJDTprnEbjE
nJQ3AqD9006ja/TQYREXgVeFMTcSsmMXAzt6eChPxOurxlF+MNqY4/YS4r21hI1F
KO9vtmhbnG9EsAIZqwzVQHRkTM9s7wAqz/v3g4vDaGDVnisLIl3lRFprOMrHQ2wY
rNTifoD4Q7AiJF8JFJ2+7tBqspQ/QsdJ6Oy5RyBBpbGyfWg3eu0+Deww3y49BdqU
MKm8rRf4i03c0ePBbiBTwy5Ht65v1XMWloX/lb8u68B+bLK/aiWfhfsSVUm2agNW
G/4IuW7tdt3BO56/HCWunU5Vm4uzAq6SWZNu5n76DyX7hpZ7a81LuataSa2X4Nnp
Zfjym/nIoqIte/Z3h9GJALxmAj6adS0PelJdiuKz3NZDpZB57Po7WOXSzpy06NHj
9QatljeqrqDHGbhFy3MMhqZ80Dy6bOTxdvfdIsbKQzWBqr4iKjLkn8LQHmexJyRB
MgoNaaNiRyw98r1htThi3Ku5vNXLeedSqk+10rdkonWOLPBW3ScR7kVptaQ8tuSU
T3fbSNUw/nibct4PAaIApoZdL6dT7/H4BAs0dp2zSVb4XwAXMVlfPhwYtQy+wiD+
4end31OMcOnAeBEWbJyPd7L1EfDg7Q+E1oaB8yMGIC/uvp6wSPilRFklASC62nI3
3UoLDYYERlkoycGzRXnjGhtvIPoMqbAmCCaaE4/5Rz6P7SBZhKFJlCdDSb6HN2MN
LcXMdxuawomZh8Gf32iCMqsHSSUDEUiTalAOMysFuGjcs0cZO24TZBwnd++U98va
6I9GsQVlw2t4HYw1oDZ+O1pmuqQesuObltbLEO1FHpYG0mj4e3z7FzsgMr69k3//
jq2Cn6tuAu0953k1eqvuNx/NoVo/EvSQTNUet6kiCRJRozR1Loenp0PNq6oWpgYL
GPlSjd1iJcz7Cd1pNyUGPF4vyMQDkcefady0kG2MKHHcdDms0bs5IrdE+cOxcMLM
TO0ckiK8tahC4kG3JpebPGHT8pIawepGk1QunXwM0GTKCRfRQX4waVST0YUni5Lh
cCv1jBRfdt+mMnMHxpZTdn9pg5YA3DOiqOXeT1dnJgasUeinlBvz0LfJezk2DqLb
NxiTiNVtp4iLgHHYc5NR2VjcqikPG4qmetK8Z3LkWosEC4n9JR3CzCxe2L3Dg0vq
FdmIUACfKFgsZFJZkansAS9M72B+LOu09sxzgWyr7XirYBt/qD8BmUm7vkSjXk/B
rIM3djfPG4mjecrV9VmgxJtFLLbCXHAZ1eGk5keKBEhwnmG/ZfV0oQJ961RvLzP1
sYWXhOG8Re2mvSD0Ybp9AMdpLZZO8eoKvyUEiJf27rhnVT9wNfm59wznfnyq07MT
Utg6DdgcA21g1J3G0IDZG3eYhtE68ml6r9UiF9QPnziFADon3HGd4GqM7eHp7Foo
s9zv9akdbyS4QVgISk5pMg/y4k3CwNwtxuyfdQZhpSSDzMhUPu7O8SiohnFqlBK4
UenGMl9zVCi9LXHeB+Marw5FDkmhxlZQjmG1qopCQPm2vN51lGWFESLsjR9i/wcu
8bYDfrCAC4tXUeaDsAGlpQY0qPZWqQmcLMaB6zCZq3hXhIxWFr8H7SseGTHUy70o
i3DHSVKPTG8DXtzJMjiUkWQTCmFLrTpihIaEWNL1CDhRKAK5OoYul6nk8ljZp98c
olvidsN6H3g2t9AFRbRx3zta/CfKkS/mznHc9b5uqnQS4QtQgnECsqsfbNTJu+iW
cJIlCCsB3hHTzSM1OhDQM2215zLDrkX0WYH3AJhWXvfm/w8SI8O8NMtLqdFEnkL5
jjF58l/t8ky70ML/6bcPkMFten3M4EGxGeccmuDYWkidv6ZJ3KKJImg8+a8kG/Lq
+4OUk5FTkr+VOCBLnK3azgNH6z3X3LzxSuPOFFQUA2BgNd7IL0tCKIvzUaf7ehnE
ox6+kOrE0yJrG/qHzpHnybjK3PRfcLP42fHEKZsGSB8PVEckKgR+WPC277lM34Zi
HWIX4LnhmuUZZiwNPlnFUowNZoYmHtxGQLuqVqTPeiwVYT3t3vFQUqS7MlRdXQuf
e/NLwFHSm4Dun8M2IQyvXFOgP8MY0ACD/YyoPhv9bd9KQie9Q/e/nqjG+MPT77Mg
PC4fyyPoR5k+9HVUXahXwPrlzuuBY9sd6Js5aCHN+AcbtyvDtWJGV/LZ4tYt7jYp
Blb6i+afrKoMYfXBgwCCQbANCJ6YIqPMzJS6NBiVCAb12rw2AZL3c5ThKi8CpfvW
/mWwO2Zl3I9GrYHulHojYxWm2j7/H1A0YwLBn9aJru9ZkmN8B0jkOblcucfCGFdQ
sGnh2vVpyTUbk9qWv4pMilzjBUo9tGv1W5QDsO2rwqasB5vRRNOt20YjjlVcpzI5
PB+WARv7cEYd7yCOh6CvGXc2DwKjUyPZ1e26DqTNelR+SxjLQy8rZ/xUkJ9SojII
EsPAaofZkEfx04usyjWVKWa87BAnD/WIYSS0vDjYqNg1RTJjJTqeIGojsA5Rnbu2
NH4wOL1wv44xa+f6OqNMZJiMUQ2kAUGjKRteBocZKuWpak13cL2Vew3EkJ4DUvQ1
qHZq2zvJs08RbI1+Lfgd/y61q2AMPreL5MRq+tOq3ZOGldfNo1WQGILzpTGM3pf8
BTR3zFxxlRR8sCZDmi2L8ljaK5PviQmr8ZJpPJYw2/zCDFMqqcL340iUJMN3uXzP
joVay7eOC99SA8g1j1QOx1LkN8IdeWei6gD6JvSaQ3I7k/m6wVJh4EXIRYGAoLPd
8D++ekB/1bK5LdbtKUt1aGhNwHphmup4A9bGQ1b19SWxHryBhucHID/HztiuP2Py
fFa+LIG494V76vepcLWJIiE5FkptM2+amYPGxEIrs3bLT6Eev0wljRBH5pxSbsl9
3gg61qxoO0Z6SBk5rlbN2e7sqq2Htua1Va1YFMYapap1lmcZVeHOZ6LkRUYYINUy
u1hy3d3cGyeFydpPbQRl134b021RkvTqnQ+o1DUO0YuF4+WbzztGzNuOFTtzUxDa
omVEndCunWysffRxVLEUJBLb41G5wDQYNZ5JaZJe/9DvSUyAXdDLtdCJKIaDDh57
RtOdeTUvhVY66S9PQhGZq4ZUYpNTaCe8dP6n51ho1alGDD+tWCBiTL1VVb+JZWlL
HhNQYrOHDWpbHah9FrWa55ZSjxLFohMmoJTnJ9CyzOlhm6qPlI/h6BRwC0k8a4Cs
I36HmYcThZ51bw5lMK50CUW4AIuyoDAsst/VQUwzM4HN2Z0548Tgrk+N5/gPcxvj
bMmKV3CJRq8zaFjwWfW29RRehXDmf4AEaAgHdH4mBPyaaz0+8EF/lca68v8GwKFm
gstJ/zvln1VggjfbEg0MNUZmeCJiedt145GAqJG30IGdO7S5OAKsW2p7d+SoSxK0
e0LGU8dp8+FUkpB3CnHGyvvzXRJY4Buez6oz8ZM7N4a2ZP0eXJsS1gKdTCR/UfHj
NekCRba9THBw+mYla9nJUWY+7EgZGJyLGlWvHhPuQ7R/PnhypvsmV0WXxfhQ4N2D
9Ab5xWw0+YPSuN4wg6Xk9JoKBuoy+0wxG41Ykg98ubPGRsypE8SDLGcadd9EoZI6
ZyL2nXB8OpCcpDQi7aGknnxBym2sD4wxZSrrqCFs/xeEoE2egMk5vBJTdr0lJj9h
sDAnBmi4siUUbzaTKd0tPBENcuaDXjWfzp1mqsiN8COZrh/viZ76BRBK+Juwi3Q9
Bf5OFeC6E2ZKRO58IvqnrBZkPhYNlp66UctBml55kBfznRLO1owUJl6LyKPSQ9TZ
YxY0GUGhoUZFE570Z1OAtCMf8YqwDKCv2a0o+K6LQOUTA7++6ZvA0hnqUys43ffI
wWEUdlr4KMgZAZFAShYC63S3tWPZlt725ODOI6qOZ6VnHcs0YeETDsmi84Deg+eS
y1iZB9Fz8lPMbwRoSOnnYQvtvdgpP4EPt1FdvczQnIW23BppKyBnZdOnBbVRbhha
z2OHkGHJpYxEGzA97BWx8bHnvOav4ImE1o7eDp3AU3eLEmL7WPwz1J+01mFDex56
Q1lsqDuAb2RV0ER+KQsOpSC2RqoQi2NjQljetoQOIvXzGWu4plFzQCYzZYKmViFZ
TnyJStbYHJNAmUrYpWlc+WT/XH/oemWGytHym7u6q43P7sMZ17IBeVqDmLhtrw2i
ms9Zq4W+XU3rgvjtFcCCGkAq/I5ZBViqc7ibGtG16JmiZNj5+9bBtlZoxRXC4hUX
xyfDdU4CcyBtfZIkkbYxAz0mDRM6S94TuyPIUZVIMCxB4UWFtqH3Bbsz0GCAw38g
oJPctc3+Pp1jpyks4/Zi/HuK58Ak+jikr9PpBMRKuBjIbKazCICbNx2RxAk1Gfrv
yvxETirSym630R7f5OjpwwPyAW++yG6ArPDwAryi9YvdkEVjHwPO7xJnrWBsaLlS
D3BIBlio5OMN5dugozJbvE4OBgKn1J8yg/rvJzjPj0T1QMfqSeVKhfs+q//kvgP6
33wPp5UMmepLbOdz4f55ye1RlmVNeg9QHIhXdIsLp4wy1vbmy+M0HojH/XMBdxEa
qdpVFlf2sfLJU7VMF6YIDTgEasUSxKfvzfiWsvB1TQraRpAEqAddqqOP3UG20nQs
FMEkBsDpB2NLdzp3YQZmWW6UYs5KYwEKyKHPat6l5SW18tHu+yva0DBfenYqMTIL
Mcas170H6OLe/o5KFmDKHj0lpo27roLtiuoRlVgbF8q8q/zLz4GMKXHh9eGSD+4a
wKtldN+UwPb20SsEp5eEZz5yiuRE6sZ33FjZZmWnG+yV/l9qYj0FUQkSFM5U7hWS
PTB5PNCgZ4czUabYzWqYV7zQONgObQhrl0xjzE2KFktzDHIefBS8XqHVCd28wh7x
kdToskWPPqugBbkVGXHjgDTCZ/YaIpxz9KxmphTr4/fusUYRNjSUDnBHLxLzUH+t
0ILVZrMuVoEbzcjIhAnE0Qb7B8dMGxnXd4GpdsOaXjIFJOcWXaE9CjjSpC6kTUUR
2D1JmfZGA64dTdCT5taEhz3fk9Zza1tLeARre5tgLoWX6qQombzyS/JDJQYGBMjL
rrma36J/1ZkXfj3tqkqsilDmNGkh0hBOT9qzfizozRZdp5cX8Qie6QwpnFc8utRC
bz2fJq9hpEA4ds04xHXXZ6ss+twd+ggmtY5ugSpg5t/g+A/4X3vWVj2dDdsitz2Q
z+HXAAMtWrKEDSGSyeLd4iv4cMYbhTOxX6pBlt6Ko0+vgxQaJTkxZ56YzcKGXDwk
cPQ5qey8icmUmTjpr1nGAzjD7JZ3BzRwmv9WF4EwtOJWoJEGXG8oFAdDatimed4g
XNlp+T98xi55hawHjR3pLJRj3qrO4v9AB2d6igd7qIL5RDghVS61e77yWW6nZ7v5
axm+NgS1gnqzavyqJLC9qlqDgWHb2xZ7dSJKFzFE7TKQfNI1yLW1XsZZqwPLyTGA
rjXVN/e2WUDwNFH3lNZKJScvUugBeDs1jTZVNJtOSUwuuVoyeuUqB9St4iqM1918
s3Gk0pj/CHes/TjzNBP8z8oYQDfek8SippM8TcuarTYE+OPq6X8HfRJVgiSUPo65
dcw0LAWaVqO4BCBVp0lbZs0+LUMAb1baRvskioYsMbjgkd3ltCEaNuZ9nwLDygak
V/mm3R9R7wmth/z6Kheo/vC/8jlCvymma4JHwlHSXLdNCk51OxYgQiAAxIcakhHq
NMQzNkRFiEvJMhKTogH7DrA/soo5pychrGC9xBGMf/0wlppf4J8DEhTKdKH4OzCB
2mVX7Yh1RQp4F2VZt8KCiUG3s+8YHb2nluLRVTSHVTr/P4oSlcXMY1JFtglxHnTy
fdWRHBgfL7EJ9E8dMvJB0z5JyCxfSY5UX6DyTFocO5F+hBad4/SEj1unhkXlXpfQ
JZSOJksbojKW4r9n2Qmtw/lMWTILjxrWZYFeqF9JyXzWeOPVyA6deF8wibWY89pk
sSmCskJus68m9mghyfLtL14adJ38/fishzDiL9abCA8c4bTz3Z7JE+UW+zAbRpUe
bxxBbbUR4Mx7eVBYE2fnhiWTg3rbwQXijsOSgDCvU++C4IEJRD327Ig5Se2eOQpc
IAcbmwfKUvzcz5p7jcAQaUhdRRCfeloHY94URJb2SUXrUZpPbJ/JGI2MrcSTg5kx
x2sSKy72ZiMxs0gaQho11bLa3/g/WFy82pvyTRNEnz4LYQ9rNtKRakF7teFfO8IK
FEtFDMZ5f/J/07YA+iFIyOvpJm1cO2/FPC8/au8TxwQ6x5pPHvNkW6ub4L2nSPLn
XMoK8f9EfEbvPuG5gdcThrFuKvBICaf4YzmBHrWr7PlPe62hoGSCrvf7IBpJygUN
M98FDepVWE3okHmCb8bj5mizgqYvHT6UxjB4AgZZGJp70xUzUQoNEa5v+p2mqecS
YKBvcp3r/NqTpnl/q4HDcg/pMokPRGMUQkv8MFOCo+S0WrnQEh1WI0G4H8WZtUpY
7OKNd0XAAFWZ0enndqXSc2Li4qFK4fP0Vwqhkl8BLT/dTREF2Gbzs6c137f+mNVS
j+MC+0TwAEdTFHbt9Ry0bHH4gRWpyVaE1f3OEFHMDViwXGLHeYBRGtL4lMeXCeJ+
O7xZngm6CXd6btdamkJSg1DXkUDRmLN7aeycbIVGO7N/aciREQEQ015Ppn67x+u5
9Gtu2KZFD9WrU/5iyXM+29fI94CK5PsLqQmgmMxwezfJIqUFg55r9WvX8ZRJoUEX
zEFgkqm+K5ZbzwHvkl11lgLvsOUgk4P8UP5kCWiVdfLIZEJdTc76ntRwqS+IBHht
EeBnCS1SHfctbTujxtBEMNxMMs8SrWOuKi2+ta66rhotRkJl//JxwgjtBK3HY7Vp
1VsG9uuR6p2zQDCDiuTkgkpvLvtJxUPKKAabqX/+bHAInak9nyi4vg9P35jp+MK8
y1KGAuNctXm8O3fKFy0kDNaVSPo4VIgEYPPxT4pfhTlZ8jEbDpRVTAFAYXH9Xhws
Z656OfVKtHx2Acm2I9hn0YHdnptrg5EO5c76Oj176TeZoZjK786MYTCOUTFuKIKG
d+xTv963IhSnLV9JaK7+sUc6zQ1IjnbVBWamOoMGgfYMr9Kr17D7HUOM2YbJpDTM
utuOuP5jAJajAsGK7/cWWlQGZtSpfDot6DhA+I3ydCQQVS661iOa7wgpeDpbSMME
s1kg986wPi0iS48v/ClLa2/VrkwNbrBpSNbkYNg3BN897a6xAlbMvyrMm8EjD9NG
IO2C9uu76Ni80YBo3UJPzglii83aKmf596sLH0NfWNbwyFZGK63o2EFRQnc1MqV/
mLIoa97TQVYHbm1WzRQm14Vs5lcJZlrN/vSgHDsTyFyhKk+YAII0wOG5v0Y7muYs
k83WS74CoLKPqE2QxRnZnG2LPHK1O3+xkYBVCZWuseL1ZGKKJg1CCLsN5sYAL+vr
mQddeoj3hpnsVdqFf7j4rEgLka3BuD/v3TKGbZo9vOfiAIRoTWGD+ycT3o8M85Pl
yMrayxAEmL+DMzgxPMjNVdWP5OlRGBPeRnm527h005Q7+egw49kG2RV/XTEDGMsQ
bJJPy2ZVznehH0Qcm2rwn8B3qKE6Ju8UbW2gbuds6HbRqSgJyx/WoR1xlmjlU3FT
maIiqnq39grZcuL4puqeaVX/aSNgcNv23XfoZtUJrJxmWEh5cTj9m0MQLzUeIsTK
vmzGrSZ3XgB2mySHEuh2viox3mawWhs9bFrlphRlk5jNo20D9xgZ+IweZW+VhWJA
TXKzTfwVuaizSa+4O78mClx5vFcS4rKqxhB1tfgnlTDRR1ILnfD2LmbbkMwHtpce
iwaxML7ahyD3yGAbv+ZS0pYW0SVSknB+/lEwlgo8R2hGpcv8dZQ9SvS1+dxdMAP9
5dCoW+6DxcQ9+IA8fGkIgHUsPHuVIkw1LxLMbstSA4xMWei17i1TlF/VjiWeaAxG
HEtHD4bJtO1RaLDAAf6FR2+qO9LmkSpIPJQkLWuda/nhiMweFeqR/jhsl9wp7qEu
bBxYrAsJVyCY9W5/51kQSuMz0gxPJN01AyWU/VagdHl+NCsE2xbQ3L2pilqVUd7/
g4PuwIIOZoluqMietzgX5MCBX1Yf84pictQeEyrzSU4jNEAdzngMO0WWKliryyK2
Pp8/VCdoKOk/tyLKj6eY0Km61WPe5vPgvQxBL4E5SEpGHxx1KZT6tLyK7WU4RbV7
dKK8W50AsHMntrWSyLJlk+AF6jScjGMZAbF3MPRlbLCr6d+JBuSMlCMcdEubMP0v
5BedLEKU/7Re1eNV45kFgyao4wyOaQFeET0L4NuBUMFWnWmk2x/yjY8glrMAqyIV
PWH1SuQZrxSz6HTCtf/XUaUu5sFDW95Q8wfMjg8ikEqK1GF18MUeM6rzHdcJ0X4Q
OA8W8/KO2XkNh3t6aXRKRVQK8+jiMOWfbtCU+gHa+uPDf1eaXUciPnOXtcWvK9sW
5VFlFAdgnKrFJgKRn9z9VR0YqZQRtVPGJwEH5KQwQOh/FZQ5xjlvEq+FTJUni5HT
GN9FhEgORcm2PjXhpk9aDy6NmXFmfeSJrFHIYcSADZbNArcSnD1KKGnhR7d2HGpA
lOIKZ3F5oUt+Kh6IFneb9vPfCbysdt1uoTvfVGaHkih7CZnDFjeLqS3Xur+y3dIH
iRLR8ItqcX2HnDZqFb2ujmwiBRwddyriZqe/FH1RNs3VdkHM0jdRvLDmVdMcu6xV
EFjxCFfG1Cjh8tKsIES3WVIytj/y8MZuDFsZYlPt5cEv6l+hldpauPxUXfInuzyH
hT114roCqZNU0l4FjbYWZ7wXeHuPuUJkEaliTFTnc3z7epwyU+gfB8qp8ksXCAuh
D+xtrxokgqxbkquyyN50M5Mwlu0GmpRNce25KTorHPsnW4WAhww0oA80LvWJv3J7
0zvFYmGkRnzK54nCfbtcYslMlDUJi3WEr/z9EdCQr9+eYlOp+py4seQgL61+ZR+G
yzBlUajpl11031NHEFAWQxyrCoCXnjtv4VER6ePTLz1hc2hicIUeDOMQVnzzwGf7
VVGCORBmqItWKSJcwoLKZDD1dX+V5KjbjsculUPS8RUxBTnuTOLMowk+K0VAb511
eHD6pTw2FtOBk7O6yH+sfjd0dZi09naEVDX/LqUKQB3plG8ghkMhN5Y1A4mEolO9
5RHk/VT1mQ6DD9EfexMefj3o7wyaRVjUGRf2erBLZwvSW5YYj7IViOPlcToCMmVW
hRQuelaQxNFCB+PpVX971/4aUhaPBf/r+xcVVsistF5F3My0/t1beFJcUdKMgocj
N0zJ0aOjfV0Id94VEcTEn/dUVNXp01kJ6uQeDcsaJyX/j1KDGuEWdjF20peNcGe/
L9N3j0KEXZyDGVeqNuXzcbdRXtaGM1CtDOnEU0hjkuCSyqbwmp6p6ubiSV5ceVPJ
5F1edDUKJPk5nwtUTM5X5N2g4FRqgft66eTjEHBtT3Txh1ULIdeAD+gA2U4l606L
yN0PeC3SZkODbJPzWS+64TdekHHkttC03+jJq1FfEiUv+xyxZdsBSa53ziOtjOIQ
Oi2eUwzZ+eIiU8ceYPXJZ8L6uGGBN3RmYAChO23yhksLRZswWRjUaOLyChQvg2jH
W/Yap0UMvogL5VzRpWqVHpi3wGahW/0EUdLD2KwM1LARTfikMPGtA8D9cFcJEF5v
phsvYsZdcE+g+7s/8xnZNbDVPTIQA5xJZ6C7n9VVdzTFWn2ekdVZ8UrTXRKzO4Yh
yBpNGt4jXCd5y7TwAtHX6TfZk1wWJbP2H3se9UOqD2MXxC7rFg5l1wVjCWVZFvTw
ZdoiJlTko7485rfL/i4O/9jJOQbtWDMfkOOjn1WeY8ZHofSY/kOYd6La85DPRqlg
5yh7qtK4Ntr1yEzMi/LtOIHcgfRjlljoJfgt4Y+B0RTN4gNkP2Cl2HL1OMtT3FtO
7IRpnaRE0gQPa3ifYCzCmsRb0wVkKFUpMNjjSHzpVLNiFzHEhZUDKuT2RC0nhfAD
MgklQSJjRMKrGV6PJA96w53pjzKke/n5sbgO/2+Rsz3sCeU78BjnGbpyCenK806Q
pohY3NXliq7PBZCyYF49D2iAFDD9xRwpIhoJNpcKsv4n61xA1Bzg9+XrQGdn6NRA
fc8SlcVBDQBTsqnfx/c6U52/E+pFk/hfMOKrGGYYL7QCEIMzs0G+Ylw79ZskBGVN
Ac2CvaK4Ky9/9KInZjfkLYw0bTfXpnh5ZmePSxKqtgoVc5abxJ6RND5lwqAw5LxX
iVSAlif6Cfh3LGzwnkVp1BqUOfR+fp6hdvuuDRSCG0kot8s36S5cszuOPRtIzTv/
/fc2hLe/TFJ5oAUy3YE/aL7/krIYIyX7FtTRdUx8mzcWttwKTXjXjh7cwSDbCele
Rnubmx1y7ExWTpK1gDalz4HMZEkge49xN9hdMFJBenuj2XiBcAnHgXqgE1oUbghr
pgstsjIUBz5he1qpJG8hiYwO+DJL0mNO76ibFvIIIoAjAj7ppbEdi+o6MUqEKLGQ
wUqW5eQkrbhifZj/PKimfxPateAmHoPJ/oBjLcVyKy/tdDAf6oj40RJcU4ie/BuP
nwruk85KIeVz/q3ZDYcEJCvGC6/+QhQzr7Ximtdl7/qPzc28VmXp2vbPThvWl1th
25FisA/int3upejuTtKelGJdfo+tup2UoMXM6YDoAfWZX963zUkNqexnizwQVymz
zzn9CmLtavg4SWgfRpCzRQZmh7dluWhFoS2lsxKmte5yJkV8Fo7bC6drk6p3Dx2h
k+hFCXU5VeY/skG/654DHzcKWdCdv/W97rEbTiCj4X5IkbGu86K9HNN1dCKunz7L
U0sP2CPO66QN8sL6+5RusfL+bdFGiDBzy9/mHmLlwAW7tQz2uVFOZTNuuUCtdBvT
H1L+YIq3EWCjduliEjeNzpE5D7b4YtnFuNkNQWacVDYAIyG32iLv2QtHZgA1+NgQ
2H3Z9tvXOdZzqC2w4SDbWWHI4HPrfcO6Ewd0RgoPB4v3C1veIGaz6pGITENa3R3W
FdXC1gc30ZXLkcwT//fUJHghsPu82SkT0F/vQ9NKrNQY7fTdoykm+JpyUv1e70d1
TsdaHowrhgQ1mmn0xPD2aq0PpqEXeSmJnkwOtxj61no4dxGkmWUelw0v0i9OQgEH
nyxGL0r4ET+MrXtjWkukqA3UGN4cDa+PVXvnQILP0kc8d1fJt7HmKB/+nQVmfQJ0
9dJPQFFdsPKIuB+Fj25wz4JXaOx7WZForlqShYZcZL7wz87hPvdEaeJh5LYZFp5f
YoxWrml9+o7Q6nVG1rsA4lZ6KYCqI356vq6Ncb0Z4RwhGQRYMiouBGm9MlPK3ZrV
C5mjC68R7W4pLcPu3ucQvN4eg9orlxFiEw+MtEqrUAtdaJT1Rd/SGtp+X/ajR29F
AZpUU+pSYXc5rOAXH/isLiC7F0BK68NqRa/2B8HanZaFqBWiweO6T570oS7MbOBX
BTjdANf5KciRo9I4wM/kcb7zyFzcN5u+IIR9TE4bz74Ib5DyLPDD3jfxRVsZIqpJ
sCu5AJQb3wGypFMk0V+VSjCC6XUCgvKceQtBSQuwYodagDCtoPAjO9teHm6T/gIg
IAmULrmCOzewp2SCQ0FOvCn37eZikZvFpMgQHpfjjupnlcreI4Ff1+2dZktzDY7J
jTKfoXkpJC2fSapzUwZy2DbvJQlNF4lBetjNAl2L/688tqrwyQglPnGxydc0ctLi
rfct8JSA7du/3Iilkp6ik6waHL7+orGqZ4zLdT0FERAXY59J1iIXRa9TMMRqoRuU
LccVb7VvuvlzzUO4ftSOR8UJHmBFKb5/zzjbr0+GNs6UFLHeZMP4PNILR+kqf9cz
1VOIFGv6wVbhTvkSiD0yqX9fX4fbucqyl2xVWR0VReMVNcA4Ft0+sBFPt9g+242j
8bokRjnqBgAnF9hVjeaNiaNsijJDyTE22eXE9s6M4ZhBjZrAIQy72YVWN4FPOW4z
g4SpWGJYNup3qYjtwng5PN53JgCxEIsWBxAXU+tOg/2baezVwC6CIQgdZYCrHuf3
2vAH+9tzkysZeR+e4Eo9sdIw0rzWJIRfWEIrzzh4759urOEVVtBt1hfSlvXBUS/1
ERIKLJzu4TQT0rgyoe6O6RQILGJietqeb5rKSFdDdvCl0NqRiNdv11SqiLtJ9tYe
5DU5Tba36kdbL+THx7AYZwzbVGqOdAZIta1sgvRkw455i7VocbN4/28XhgqTz8A0
+xY4Bcmpyvobh5z6GqXAH6ZerZ4JxfVjzclQRLRdTHt9JDyEyeHn8ozhzRU2dwV9
GRXPq9zwckFoulZcRrEcUepTDnxSr7c7uR2kQ52W3pRWXwuyq/YzRB1tcz++crX/
R9nOrORb7VggL4jK0+kmVb9NN9ahgpnq5CoMK3603ffZqd2AAWSo5tD/wrTmAhoS
AVxm5d4+oboOef1MZObEAeItsgF3PJQ6JK8coRdQgsgPgvZ8oGu8JKYVawpnfy9s
u05+u0IJSWtj9sMmV+PfXW9K3SY8zMcpcWUZWFzlLfYn1DHGqq6EKbmOsupWQdmk
b5oMbOnkoVf93syeFcA02ei6f2b33waUQzUtc+1Tp7V3SDK+1LMSJNDKgf9Rr3cQ
XRUXLXSp5203M4BzjqezT1OFaB56L+mIsEdwy2iy2/87q+FzJ3aDYknnDWe5OgCK
PUx9RgrRPA06LSypQt4niw8NsOVYy6lt4zNZtKqgncxxBKawa3jCIcNgYq+52gmI
CyeLid3Jclt/Anez+6g6BHawF6eByj4zbvndR6+UkzA8X8dxjw/8o1Lb0AP3/TAc
bFtnxPRDWAULgrIlvoMsXGoiAxAhO5GyWHzzhtSsp0e/zN1aLnGRJaQd22rFsYKH
7uFlZwKyefCLXCiLHl0tkL1S7TnGBpsD7tNK0DL6FlQgvUTXsQhIpOQKUirHJRc7
mf851lVAofjtJsk8LCp3m+oB4yZT/ec2Mu5YhgFcPCVERhmTCUYtvU/ArkdZ1QMM
yxmAfDZ89bO0QS+yw6z8qZt2oqqy6Oc4qFt6M/p2hHfhorPgdaiG+kX4toLlxZh6
ug7hJ1yVAUuAo7/wp+z47zymh2DO1V9nAeOLvRllvNsBA4bKZuAZ7diAoku+30wb
HNaWpIr9lgZTSGWF8Wnv7BRFP2OSBAxVafYbgnKBGkGdqgTqPVkKKiyHJn+vXfoM
n5QvHGDXe+UrNpt1ZRpBn9hViws0EpNA7ZW5gBUJF1L65kseEJClo7Gk3/h+72ir
y/PVufpJqqzZ6/QWZN+X+hr4ZiKefDQZicD6l/Zz4y3egkttT7WFm9qReHGN3tZs
49LSmKDuG806ZBP7etDgS9Alazy3EGGZW7ZPZcK3VUxwaV14b/+cu5xl7idOc9BX
B1vB3SNt57w2P64k/AfwkCaxmGpVdaZKrwdGbPaB8SFVxTLBomsxlT+MKtrWO38/
xxjZI+dPrMGc11OhLgv89UHZeSEQUaLdV8gYkRn1HXiscv2kUKLp+COn6w3+rEs1
PZ8WP1WNbZS2h2LGh303RY2b/uXMmmcGzaw1OqvH+DQCSKSNlkxzv4v19Kx1VEcr
71n8YPEOCPGdsfdzS3wMt6mvY5HPrtWlSIcHkrzhjfjBNM6j3qYhIQU5tniU0f5S
5zEy7W114eDmtl6y48FOqYmKYqQ42N83jkLQRDZyvGg+k31k3CuUho7jJm/3T2Wf
NNf7/7ylCWD5ozb6Bzjm6JsNU2B7IogdCFBGQ28do2aml9vXF3qyn42COASYd8Qs
8C0ArWwjD0OG0fTi04AKFB0UgKz5cbswNfir+BRE2RBqYGqJ7BsK7qK1gHN36ob0
1K2TjiKlu+M/XGtSU+DKopusfWcD5Et7A8DROnNaRSh+bEbBC0FMVAbKwoiaHRIq
L4q4iEOhHmUNRbz6oyBwSHQfpFvVDK4gfEcrWEHnMLwgdG+X4Cxc2MC5HTRW85Sn
4QlzSi4RXf1Iy0kRJ8avxUXek/+RZmz1L5I3VtYoI7Q2Jucpw8W8rmQJeIEZ7cNe
VcgEqqJLcCk5N48dUf88J6k2zZHkjFWRXhqTb/tPqmGPbUcwE+D0QwtyslytJ0h7
3hiSJpOFEL9+tRpZOlTn1uKXnJZPZuF4Mb9TZd5DsfcmocdV+cJM4UcrKJKERKxq
dcalueMVY+WOaHk/j34ldvLPRYlGQJTnKfeAW3B9OEunFDtbLz8/OkCtjul1yaeX
RSM4WyMvAQWR76gl+tLR0kYyfRJAfjCJ/kVwDdFSt+CnUDCNgMgi4w3zutYONP7S
9QGi3ri+Pt0Ni1WKVlxJkHnlV16njvGKk2s6Cq3/oTijoy6meCb3UAr4xxBLtq3Z
SUkSgbPVNxbH5x0OA/Y56OLlRR+yrvk+u0e/T/Om55qxIs4AYdKE63Xg09nhWVCJ
ae/Xep/nV8NfqxhG9TXd9rWhTEaOPs8BRZS8/ZmzziUt5sVR6fVfiPfZoAaYc9JM
EA2cwWzcE0or49gfK+9Gu1vvqGCMRydBklsRVhaTduazjlPXj6JgVmHSVlo1DWDf
jvc+VhoxKccNSNeCVt/11CwnM2cIh9j6WERW9XMby1DuV+XoXeaINLPITjRRdNls
GqqJ5djJjvuJvHDx6JdnyTXS0NZY7eO5R3V8WLQFmtpESYq3iVy1yF0pzRkZurS0
rj/QlVIRL59x47oYua7/DhCSPPLDkt5DDWYUYiStp9s+7PyCnkIchj+2e7kNxY2k
fv/TqsX62N1OxaTUczDQl0KwTwaCZpFQ5Vk8pYosenCx80pJFzC8ndz4gT+Ds9+Z
1LosspI73ssw5LO99RQ6kKeTuzTd8+UPhzvGAHN/M9+2odFidV7Mxrb6zE81yOaX
xcAPjMmbhItNV7H54W5UZTzMoF11JV8OtLYdK2JL8YykjmaOCKzR8ROlVucEdTmV
jiv7bRUNFiGfEPQn78aa7yBRwCDO7xz0bKWYDLHapONTQ8nScDyE6JrTmgKpu3gL
w8As72LBguDa+jO6bbrhmcizLuTKxTGvwVqDc0OVwW9hXUQcYX30JHzrYevNPqWE
J46WFUc72iKE74VnT2JBJRHFx72aqstXHSsJksvWHkEYqbHpXQq+UrmaFlkfNog0
HlXydrI+nqVV67DxxsxxvIToqWB+VMET6fHyxX/CG+2VhUdPFpLgrnjwd7j7eKw8
uXyXplOcx43JJeVeFmclmyhlCcbgIg2mdeyL7TtneEq7Y89eN6FeOHdlSwqArXdx
FCvhB6hd0cQTloXhSklVFszz9ARkcjH8PSL7Z4elhSbQnGgC5nHmfzgK2P1I8uHz
+baHCER0SxI2Brvmui6C5JPU+kSOt4N3EEisFHbgfv7hCjucmkg0y6WWnFm67dw2
/IeUrw7TEMBAO/ABdo6sWGEu4IdUUKgWQ6VSI9F+KMIkNSSNhwvbBEMMJseJIfWg
fBAOVMvep9/lK6l84pXX3jGSW7M5wVjzD+L562JN+OuYMLJszpyUVOFMWZ87vECs
R2I3+PJqcWavVxk3x6R/HpFmH4zL8uAIOI/max0j0AxiFKZT0rpRgLFn1nm8iG8Q
OiUlhoWU/XzIt0KFxDiAebpZSA4fFGer2UpP8eoR8hJWdq4fTzfyUDwPTYYe0DzK
kPc4G+5pCCMDCxhesiN2LwdL70095rsp8emT75CaB/GMz4Iwm3JhknozzlFBqCBM
heYtEDKYzsu07c+gSPuHLNITYXjIpD+EBDw6WPOrcU8vn20xybO3mvUSNsN41myd
j1/nRK8ISiNUln9LJ1AafeWycF+M4XjodJC0EfjdrjLkbIJcyBfqQUPav8lJFD94
Pg75WUBuntfQ/graMG6AEtKhSSV8IpO/SJwyZcp91mJDqYD5lqqSeV6eBgsVrszq
SdFiCAeCaDu4Dr5Pd0KwgVWz3wyoT5yK37VQ3BPYVw/M94cJxp/FTEQfRiQIcEJS
thyZ/54e3vQGqmAcp2K2KW38TeXCrLHfVPNO0hwgBD7WLPlyVhXzLSE4rm4GPbyF
hR/mlekofe4vPWAb9g9Mav2Wsvz3A3BNs4itu2blwLbevLtBESMOWBngHv+2AVmu
NGXwE133p+ome7CEjaW1eFWzWeI1dxjKZU1BDbl8zDkdH99D+32+mg1NpM+z4Kow
q3HLVW9RpIuyufEgsG/VTOz3uyIFekHubLr04kwR+V/ft1OedupT4twHZ/ktZbNW
zkJuYd7LC5qRhbhRl5/+tIiOTk7hEwTpPb3V2cpvSGI73mQScVE5yM+RzZbBzPmz
6tPPeZXchB9UuaGL3bQ6fwvZVFG11Otp7MIvhE3x0pCx+zkgJhgnasM39y7bvhV+
divwMZ+iCZSa9+v2r1QyvguybwHBulRROiIkVbgob359wEKxKh9Igc48fQd3EmYP
O01o97B2xl43E1JqeCI8uh6hLeoz4mMNCdfXEe09CyamsF+I1sTyipji0lKb4Y8h
kjp2hJse14wXAwXdje5L2JZIudpblZCffbRP2Y6tUnp25MknjsY08pnoEx7HDUpI
EBmZLSnejkN5+1brRo/Ri1ojjxkMp43JOaSq+dagC284UNMByLNDFdAknpKbnraq
ct9MAiKiEkmJKt7r17XHEQji9l2HESJ3v+ghxjMGZG+eX4ovH6bWIFl2GsSrtc92
u00LQF7wIuS+EuBEJ/tz+AayBC3lYHbQpuxQ7vMWfgnX/XNhLfrwwWQIWvH0BEx5
tq4tTL9wBi0unz3IfJ3DoTGco3plORqe+Zr5ExTq+P+NLEDKeQtWRCCMZ781XQvH
66K7V7/ngCNw4+uYR19S0PBNEmEWxOlXoYZWFsPvozSvrMg2IhVyXZA80NCjZ0yA
m3MW/F48oZ71LEvDYLN3O6mJPxCHhu9bmexeCFz/Cl93n+cT8tg9EsbFy6aFzQsT
aShkHxmVJ6owRkAFR6kp33CWG78IE7tmngdVqC4hUubVWgBmuz8BTqP8A5zxXwaR
iGAwgj2IwXqFqfS3jC2UyLHCfQIgBQa35CNCuLd22m1aD6NglYrX84uA6OIY7Dv+
L9AHwQI6e+XDBRQVbqTr2WpQ1ztxpiTfELJS9iBcWmhaDl2OFc4gKjfqeMD1TS6h
E42RaboirX6L5BxlNn03iRYsQqOzZAouV5xZK76iOIISbMvS1NfkwxMYQDh8407p
NAyrhHpKgbd5cdhs+J8ak8OgQ6iiWqg1W2Z9dg9MevIRXNbGMaK26AZxCbiH2777
TjXA8D3bTHvzxyb6yDfbMsXpTp7Nl+5gM12qVC+DBvugQJFjfab+mtqpxZddvCzz
UFtcaSqkGGBeq/pUl/tMxj7q2krozZWQfgbw9RxTOIpbrXQiMxH5vLU9FbhVcXsU
NyAArk/M7LRgD5oiGITzhSatZ9muFnP2OmKXWT2+vgR6i3Z2sSc/4JvTB88ESE1h
IKIMRG8Hgqk3rEo4Lv/qvoPTt9OO+1pe2hXVIoDoOLD7tPPFNZiFlviZMb/ZlCHh
owLLX/JO0qCG7PFuodyc9QHNhigrHmkCtO+zEUIAMdS9xdao5GGWKCU4/YuWbyqe
dIU4JYW1gKfqy7Zr1YGi7l2x8x6pXnlUxm1TzGZuNvYyVWS39n308yLUW+qK6FKg
X4MwHGMNtj+sfzDj4q+WFv3sccHUEp3dmxXBFR3N1sxoenr3sIr07iGUmB4/RyPv
uKUgmw1yBzPS03h32KqSj8x3+qRPxmxJgWuQgsgLWmFfWF6koIxPWPSkoAmXTf3+
nMH6RQfmF8OwY7lqmhSzkSu5Q/drD1I6OA6Kyzm2zeEJzjvRe/GC+l+7nDPflz9u
jQgJIKfWRc9kC3/ax4BiZI/iTinsad/LvPK5oEp4V7bzAxc1UW3ypZuAcuh+NMEq
JID8yqr5sO1UzVaahfbxM73xWs2vefx3XOV/rXnXCSwnxs4kp+2cEiJirYEbaxgb
Bxbt7Oas4XIaXHK8Zbil8SHfLhnOt5EcF3Yko3WypHUZNfbfTHGapnw2+swq/hWe
seKdJIajW2A3mdoGq9khAiSOFEcsIGboRRf1u1wU2SqOLLWGYQ+8AbcH+b5cb5xN
m5HS1djQeotQa2YwrVGVo3IuuojFFdQbal0R+b/NXPqdi8wwudYDDTor9moaXtWF
8YJCAeA2hJOjc8qTrxTDVm2g5Vtr7P21nSectpumaYcwU5dAhvwxu1GnJcMnPiXQ
v+r8RPM73BW9kzPKzA6Jf399hEmQhngG6hBd1s3wvNVaKiu4TUCLyOgk9tdlDzkk
HWUUbYpuInP14fk2/DbL67VbdAcgvaP4W7EYREM9fBaifh6umDVlR2baEoG/A3b/
30kjs6cqLyzX4EC9PBvcUxz3qijOiVeLXuDUTWqSHzaF9V9MnEFI56/YY5bwR9O/
rdxg35epyfjQwk+H+SiAVBYWnX735YsHEFDI8AmPbjH5EFKFGXURsPHSaUhZI9zK
zQhDtoemZBE9zOvUVn7flQSM04ea4inkfJyD4m3iVpdNnxNTWmN7Py+7nzCxfPeg
rRnqSIk4igcnsB3LwBQBoTdPLOAZvczIMzPx2lEta0RlvT2F1xEZrdOhxzSDPz0I
RcXej2wcb56UpIMGIx3WpimFtHQrP4owlyKxAkQ/EGR0ezlFeMFhB4A6sD/xUj87
W3xrxcPZJTVE3UTVXycKH7f0Y4LxGA92cyevIY6Z0bGJGVYwU5TPDHue1eRt9eWK
kbu7IPipVkmO5O41LNIYHZP3D1Zu4pS2ja40CD5pWr6HzB8yMXi84Hs6BdFcgiG5
d2hfZvk3C0GPoL3tPHnIN7o0ryJrXvH5O0o5MoMxUIS4xWLiJnogM1f0bliFHAoj
IKOHpDjd/G3MgP8SN0d6CvKJMns6Qs71finXayB1tpi2AtibMAsR41eXo4NRFJ+W
wYV80mZZjCT1O5MC1AhAbLLdJ82X26Umr1kPjWXjyh8XbTihOO1WKwL/GavlQ8ua
prqUSQCIQHhaz/WeKBdbpqxNdIExOVYQLtB5wFI9gYG066KOGqKME3V8DoP4pDqP
kBQ8TL5yGuAKZGhupchUrKW/eOVguJw6BwtWuNITsHvLYLv/LWdhXxJ8Ag6pMJuC
tZZR2l/cDzd1yE7ctd+BaS4uBP5fk5zlXn0EA1i7xGCvvLXNjS5dJlivAOUsTgfD
YtJwlIfC2RTxb4iBiNZLQKwQyi+91i/UM93EDB8Nj5woF5DSbMvX5k3HSsSZBRnn
VtO7FTpu2Qi46wOezAfQY6T4Stxgt+Vzht3R8GMKN17FNcbTzJ2MH3QoBtis2Vdh
SGOzbqDHVesra64RzX4WSSXcn4Lyz/HFuVnENbvs//JiVj3bfVjj28khkxnYHyET
G/wmn5LTPkCcdJLyDnDXaWKIAsl721wcuR3GeSAuNpMk7WWsZ9Y8O5UH38uVEc80
lTqIfmJXXVsjBNITGns73wdg67t9TsPxw+0wcGUGPFjEwkcvb7WD+XTLS0obPkSK
lafcJdZpBYdYtRc3PeFgAK29BZifh0WeiAN5k6c92ub1cBMsJODVEf/nl+gH8zH9
jluG9gSmmWbxzURLLP2A9pew220tRVDYkKpwCSBL2sc0mv0lWsP9oQ+K1zWUcFNk
3OZowoJzYjA3x8hTc77pinzHQBUc16Y8bjktMzuugjCPhzuoLFQeO7MDi99YddFL
1lGMWEZ5rQoOtIoAzVncJeUXik8WO230NDrV/TW7gsc6RPogRWJXLlJ8EQEklr8R
V6gSQ/kJy3qw+XAWvHEDL3nkeH5LSNeZozUFG70qoM3j9owm6jQmJ6mGZWxHZcJe
X5U8JEuX+Q+PNTeoji/scGhqjiKq7G+/C2leq5QQZtTyaK7IgYqCltFKRNeMzjaD
PDsIQITJBAP8WW5UeX9sDLnXly+qki3JXxmWT2WVoHa15RXgTwjIK+pRzXESWTia
j+mDOXaDUMd88/7U+WPbHmBZE6isGdYq6vydw03pZDN4NCt7hDxrG4a/ftZMAHai
BbbfHhmu3SBkowQwOV5zUis+gSwEVsHz7BBDfyRSjBXmZlWmy+nlHTfZ4/oYmAT/
Etz20eDMXSGY63BNpm1txA0RXJ5XyxIsacCMPRXwiXGSAlnYM9LBGJtTPQdZYUrI
1auxHEw3WXpnSdnHZgbql7Iro4I70F7kfM/+I5gJTfswfGqXd4IvGpKClCs6Ngey
TQpKtoDNKWAHmgr/Ksm/SmA0V0Sxwu6uB5OBBuVhzPCmH58mEOmA7XYUFDIdgtWF
4GzjBS6w4b7JgupdEdqamMFuxosUqRrFgTzyA01bHb33Unx+qWn0tm+kK+6amlmb
MMeASW3V49OBngtYG6J84O5Gwi8PLGlEeqmmAyUM3ovWBWthBdq4zOIkDYKweyLp
jgFdtYO6XYz56QjjZ8d5seboVzpfm082oLHsw4kr7Ru424J5WhNfXgvtF8K5V1r2
R/G9ffbHC/ci3zzoHC6RQ38I6zoqdjxjKdqHrfqWMvnn6O7UzHfEuib42gT0YqLm
EA3ASLG9O+FqkDXp1MQ3RDfRt6vfdzhq10jMd8MkDJuj8Afwr1ERozvteB0PDgA3
rMugvnrX2VNWAe/jXbi3SLxFEwVJ/Sma48ffXVCD8lUDI4Y4AfDCxHTrPr02ilpJ
OO3Mj9PSYS+Qqx8HvJ4dF9Tept2kmZ4107cveJu1LvPBRjOmgUuu/c5I6n434z+L
6m7DMj2Rnbsg+ThbVc9pmvAsi6evnUXMbximecPUEmwhhfYq1g7f8LLQgR5bLzid
KAnz/43aOSDe1YykJnVCyQQFh27OgeIuf1NFMLw3MAuES51gJaH5cLhQ7VV44+VO
i6/ZybzHD6cE+aCENLyqPdND+Gxwq5Hgc/8kdRhQqH4q+8iKkbHsidJYabUvyNvH
7vZb6aDF60FjmtmXqnQfL9Sq+j8byfP8EKayqxhvOpzVgRXQtU/oc7JoKGMjKjya
sb3sM+TlqYMJlZgew/pQNy10XW7ch6X1vL6kximKbAsV0nkJw8Oa5GaNcvpoE+lP
HgkcruCueqmRsuUw21mYvUZzPse7Zo8lElERA/+iV3xLhIyqHP5My55XkM5I7Hqz
zYzgkBZ998V85bwM1fGi5Speg+5NlZY7F3jzbrmdBkjJs7YKDvwvrwrHYRcxBtKp
zaFhiOU7KVtdFN58O9DWk3dg44EYWXPAc2ZAiAQUVrCieOw9GpaAAzfCh35A8AXe
Xm0i17qgpjAC6qctvbS/HTacDCEZt9f4d80HSBFFiwq7+PGVYjcO6uiWUA6qQC5W
l5d6pUUmdRGHZdLAHdq8/6ZNit/Ueuc/3Y0bUdvh0VoQLcSS64pWQBGHeTm3m8z7
2t7FQNJsfQiqZmGtG9w3UOl+H4qgVjOx+VRkIl3CvfIiupapOE5tXpKSSf+R3ojR
Jm43lwf46kaaz0YjWMyrjbZX6acK9pV/dE0PqAYv60wWhW+yzsdLUz34FObXcdGh
uqzFNkaZSlGKAmKcgkLXT9bWGeW41Hj3Fg/HmhyAifB69aiYZQyN3Ek7E+FlDOtp
BRFHvKMzC/bkt3lJL7RLcd9Atz8Rp81E4Ht3ZgRLCismHMDQTfNWAYCUKH6n4lnf
2Yd484BgjdHJ1dzlPeM3rKyEv98yYzPmdI0+HGeS+TLcfSRtQDTkU9RD8mUF0n2o
HhoTdbfUoHqSuWV4RsGPi8ikfk0eBJFQlEohLCrUYSZ+5N1hFYxxTKNfpncJoxtX
GrgCutuxh2sxB+v9ntVm1i7rk2X/MetQM8C+qmp6b66K0E/c4GlSQBQatMptkcP6
WDoIxNExnS4qR+uaJz9t4LGOU/CAlOWfkk6a9JiNRahB4N1Q83nLL8xGGSAn55dF
iUr03RTR+1SvbSx1apX4nRDA6iAiq7fqKdh60f3463IZfBVbzsfmGmMRTDKBn50y
jfEtQ1OAZGeIXrwSABLvJbNv25bnGwcsUjgiMojiEgP2J+8sMJCEPo2zi8n+oHyZ
RCAbN6F56WYc2eLfjFSWp3XvrVMr+9h9KoPpAp34dqP4OFJBHn6pkxD8aH5b5I4C
EtcAyFPdBquNWdwNQtMw/sPdyJ7SQHtyuaqJOY5w4jM1eK717vxLxH/yre2qEa/m
ACqHkCLF8ZBnfIGFH0MKhcVZHFwuRS1O9eec0XetppojHK+QbgN5YS6VZA1gF2ZV
QHIX4Nm+AKr3e8BnkWbeDM+ezXl7+ldMi7vjbpvEyZn1M9vzB7bXyvo0zzGmGBqP
IzMWBiO2O/FSBUlJnn1meoObpfAfdfgY+wmY5TitejTUC21pGxv+HBLZrUFQbt2B
C4SEOM8fhNmaozNUMKn4CTD0yKgHbYRs+7BF9ete32v8sfPUkL0I2W2JBDVyNnUu
62B6CViaSI/mqJkjOTkRjEh4kt3KFCvoxeOFSurzWMOkvsWeP2P+mjquyaL+AzCy
OJfssqJPbeU9pbmTXC8TOcwy5iwDbPHy6IelVUlZuFI1oBkavd09XB/+IcT/E3k+
jotpCdUhkKunJ16lk8lRCJQsbY9K/OXJHwtwaqQ9Hpq0sEL2y1ACj0kcii6XR/Zl
ilGhmw3bIXYSaV/HmwPxuQRc9quHoNBenLRBRNoEQjIafyQLR7xbFmOomlwgi+C4
wtOjs/yKVkLN3zeGTNBftXga/17c/rAqHPjyN4uyCbDKuWnJkjBkap4Xxr+1hIID
u6DimdRAuL56nm6+sVWOMtoxOoS0b78LAYoVHvHKPJOzEMhyzstdsipFVQW9Ibjf
FAfLaqJiy7rNSXgup1uZjz7mBuCaN1PrmeSFjdXRHpYht5Ie9vZygoUjOwHG6Tgs
RAmbANkjAn/jKPYcu92yuROf+8EKwJCIPv/0W0eDVk8pTP03h4O5FyW7eyElNRGp
uUpZWcAc1XNNxjvF+ziilIX8fRC+0ObQYRAYWrDs5uqYgsN76rrFcWIH+02S7pYd
PdoQVwo4Pc3caCg2nZWmhv7nr3QbZiLowAULdOkPsvGQ8RkokyF/50BibeZMbFL3
Uw4m4Z6ALrrottOk+/QtDVP+yPfYXFIHppvJQuaOhZqKjZmcdmdYzrrH3vYpB23/
59+rDRe9lOxcwsXVhrfqpXWLCZTUKmsF/dPOxGASCcDKZg5GL1aLIiq3LhgWIRWQ
vEETpiPIWLaG5eHgR3rm2G4rmRJGh+w67cpx60WH45wdfSGA28SRHbYvOBHSGJ9H
wDJ38EUgKo+CVBBabgGR/FrX2wSsEJvXpoaFdbHIk1qP+ku9eHVug431+jRzB5yo
/59DH4Kv/NZVxrE1ivAMRo6vlIN/HoorK9PTYOWTOilIe6OzzB0cRItdXSDiDpR9
TB5AbThiBnEZ2veoQSuWYaKDOc1Hp/fe/rESA+gW0thKImYEDAo8kqpWiUkrk7b4
fm/zMttqSAm4Z1rcB/z35K5IjtDCE8EIjtPHs7a7UCjS+Uez0Q9H2vxUnGzNs/tf
wWkNWbmzwIzoaMMBkAP7/sq0PYDt3JYTlLQnFDBm4r4pkQ1kDSwM2Ww9+zWD3GqE
lto9KTdcs3F/2AQ0UCu1rG6d4+5w0IFvkxzoJ0EjeoNyy7LGr0naUwbiS7Eri1LJ
kBFB67hjjAqHx+5H36TAC1GLjDBxml8UDB0VQcWoSy5ZIyR5yebps2PXgfYyyE0m
DKT4EKCazbhPEOTpRBvF4ySYbOWGIB5xuE/k+E8kxLfXm+ZlV35rS4pwwBtonFmO
TYd1xRFOi3PatEwrpUIVsa2gA71LDC6bmchg8LmOSKXw++CgblCRLt414LztAIoA
Jig7cLFPDPRIMueocxRKrJGQHZO4ZzDoYHjrLR8Mw+4a1JzlswoD9uzElXMxGWi6
ZQooLeg0LMRY8kSK5jGiiO4RWKU0wvqAvbwlqE8s/l4ykr9e+FQQqgLH74Rlfg3T
02LdMdJpnf2GoIDM2aSHER0XRF+6CJvcvdIpsL9GBC9lfuMGeQT6yI55xbst6s6w
K85fp9YoLhqF3wrK8W7UXT9Wf07Gn03Mvisdq0MbQVDebJCTfAGHn3E2iy/wSi6k
7XyE9WSqccHrzKXU4FZPZTO91ILfwHSjc1yorgmrNg/+O1vW14yxNH5JkIwoOaBf
xSWrlcTBAvTULGI+j1pH2uygiEp/pdMRFFT5DsnbCNnIvyLhURY/uQZHz+k9N9v6
x5606YuhRrxwoz8b9CPt85UQrY5kx/mTXxwMtIR21/0rXXWppa0EU7r+80MHDyE8
PC5n5b7nTnI/ztN8bO9Udw8ZH0ykUvzoCt4NEFTx4MmZrEKQvPxqm/cdY7TfBRvE
ggEv16oLS49UdcWbSyhhExx3ThkZZ9AqMT24mZ9a37iIoaH0h+aduNPbx3XQGeRO
HZwJN+M4Wxo8q1sRBSjuygrH+utfwuNEK/Co/9NLv+HLxAuojHrzB7NPJ3bq3dDq
QQs/P3tpfynMU/Urdxa19Vu1i5PMnYjWq9QwBd91SstWQri+W7WtXmT+TXa5jZKN
GIxzHn5db7SFBwj9iKl43uoWZ/DaKKAByO/fM9j6lZ5S8qYdSlpH2sc+IJ5uoOkd
LQd4TwanZIhP7nPP1a9ruRrjd8IHh92/wQkzegpKhI3V+UjmTA/4/PmscW3tTQOT
ievruZZg2TSnDogMGWCHgH8lFhJS5dweMm49hcPsy3/9yLq+sxe/3GL5NYumlHwc
PMMkp3EwZOyHYRBnITaN0ZeZZEnRN37ZQizPUWfI07wwjN11uTmhB4FA0hltHDwa
7+UtBdtwcq6cCuS56tM+2p+/iPoDRpIUBO8/wQWqwF7ZhQj73KCcVklNhZQ+LBwT
mC8odIPEgSecqE90zSWuBSH3XEyOFPGOAcAtmPfPf/iYKqPISNMOVM5bZCfSz7ST
2SRkzxM6id3CRs9PPNi/OjsZNE7FxyZ6OdqaXW2nptXwtAOwsnCnMlN9oTIYki/s
FHPOa5AwdsrWve7ceKP1ketN3/nHfjnlBRVUvbxStUG9zP/o3LUIiM2Bk0DpM2IR
b2/G7wJCLad/0cN3w47gXAUggIo8UHzCi8sXU9sxoG+IEcJuWGctJ6dqVjNwUpvN
fAG4PZPQZWK6rO9wNXQa4s3dR82CU1biQCJ5JZyWWucKQwOaAbIiugqaSz9I+2TY
jKow4D3puvvs8ZzGK00r8mWG7L0p1v9bYaLdbVDFRU/1IEcF4gkg9VJTDeTOQeIZ
yzMdIL3mSAH5/1bxhz7zXabXUzKjCFsBfFe3igh9aaoVKWr0RfWFLgVAUTrsC+Kb
XK/10kiAF/aOnhbHXb9Y8MMeki/TsHFnIkX412QwqG/O996VscKQzM6/MYKsqiSs
pPDuUllm98lTXuZZpvGDF2EvbyZnn37A/SEgPlq7ycl/C+SoBRMKqgwQ+mrCcIJU
M+nDy4wWvBkA9jGNXLLdoPr4+AEe8saHQWqVq987YyBCbgvN2l8ZTTCZ3NB1ggZM
rGKpRruv13ZrgJWt3VM4ksng3+8uMLZGp5pcU5hsbTL12XaawyZtHcyIcTguomWg
/TJTTy5M24tUvjK3XDiiZSQmyxPgVZ/b5L0H2hmW/uYSmOhFGpxcnScUVqMas7El
8In3IXVq6TMQu3OraGPHNqnr5Pr0TswgmZj381PzR+Nyf548GmK3GWB2aC4u5C8b
OoZOKsts/gWsKUKHreCJTsVzc3FZlVVa3wNJ2QAHiuZWpJ2e20aLSzoQITW4ZW7F
yOPfuW7qAjszAVfXq8cix4BEzXZC5GFcFO5yzkZWezghrhc+wpZDBsehh9dvTCye
3kt2ErGyshbkfShD1RcHPnJ57WvVyPHRh+2Rof/hKlGixUCpnkSMiut+3Qwk5z3A
Xhe3iGCLmxITv277m3VMJHh5jlrxDtGSdarih3yew4P28P9H9+ToG0P7hyQNPqGb
4DDA1tk6CUjC0U7bczQCmQCjOUlg7XQ0QLo2ZAkxq9FI/tdJ6NM1MF/fZZG6nwXz
2yWsdqGKBa45LSasryEacfMhB2GjFYKKGH8vUhXjcz7S5wb/Rbr2j4Qiw7dVQgOt
GoQbbdIcWzxBitICNyORYr9zFqb+IUAmJPZ2+jXsadLuH1pEdRj1STTowWqEMNO9
scf+qv1sdw1CXGXDr0pwawuNGL/458Kkk+p+TIqkXGw6YnIUn1IowKmjHTP1uamq
cPzM9NCi2lmwkTjK5N3PhQAX9is7Qrux56neLo1U8X2HxVkEekYYI31kTeMFXIpb
Ch2SREosv11xyJExYrpGdoePdhJ0TFXJ7vfXBHzInB1Hv1MT96mRvfC31UbNbISY
gmt8CouKi5Mvns3C1nczrjHQ/ILnj5jMAAPhoSnHKADhC/P/8qd3T8ExPdCgm1Lv
hItFfXd9UTs8zpuQ2fQwCknUm/kTYIH2zjFd+WIWS/c1bmkvh9G4w173ClyUQiaY
hn1F7liyUA3Odw3mQCtJAqI2yDcCneAAMSEjDDLAYM7wIC7aPQG8nUSiwV1jqQE1
8S2+bmWu4zZlfIz1B8xI0sbwx7WuIv+SwREWRViHcukK+QuoBsjbCWoimGWGy8j+
w7B8ax470kOoPf1xjA35hZyVOu/K/DTSuTCtvqXj0X6KNPjueQhD6OswYL++xLzz
MTTuzKYNaT/U+pudZ5cP5++fyVHo+K2spDS9J/ovAmDIuTAy80X0JN62J2N2gBNf
v3/gkvn06yyGEePOfP0TZeSQbiJ8xIaczNxyUC9jcF+1Zgz9NBvx5xW5j05yauyH
pSlsvLEo1ROKaoYTW1w7U2DeFnmyWTe/YSvX5bydfe5Y26tS586kC3CN1PhdOAI9
7OZ4W/xLrPngShpj/sk8W9KD0agNhvBCk1ORSs1yc3jQC/2E0Z4YgPPBXu2H7H1a
97cBwpOWZdCtwqvbzrWk8Zr4avxq9OENgehx1kRGDHahP8xFUWXJgLwrkD/eSR7Z
YffkWzn10kUcMZT7bZWd0+ysU8gYsi6QHLFRDmZ1GmZTBcjPb4nIATCwTADht2EV
ETTDE6voU+MuD+OkeMdQTN5L4PkyZD2+IX2DUdhm6EOsQ9k/sranfzwcRHGkcrhH
QHuG0dBvbcq0p3JHDSFVe17VgLYqeTjZcZ6ZknDzod6XfeGlfPpboIUEX9XAzISF
CP2QZRLDtxlC6RFzmRTkUHPrzcJOLe5zzHN/goX3buqhPx6UAAXYVFVXI5kpThX5
kpvBF3OWYM/qwrXGyIo7JcL8XlfO13GLtjF4ysmyH26Y5hcMeAzJ1iVrL+r6mb/P
KPGwt/WRtV5ASLfbTcV3VejOyr+8PHiRr//Tt4AfWYbLdB/nsyMc6JrDtHHFwFQa
ZVq5LcPPWxN8sQU7IO4t2WpjM9gtGEfXg9nhwwy0aEDWNu/VYYyu/n3m0DbH1AGf
r+EKhLHUNSTFvGVidyImVRbDyXm1u7p98xWW7DUYvOMaN3dX8o6uzptHRNPkC3Y2
kGdxP3apUKf/ljAdMo8Dv/sfJBemMkfVeZhjBr/usHeFTctqbZAvbDGCx6ur9VAm
iyvlrXO963FyR1gTGTFOvbhAocw8tkwp9bgNhzL1YjCjCOtIE4qtAtbc1ztTEVXE
0/Zvrr3bOm6JK18MvK2bM7+hXZojQb4UOlJrqWNT9Z+UJR08tzi1j3xuHXPRoS2H
WxFJi1/x9PVhCL1ZuBlHCNZtIu1i9kARdNjHfPMPVov83pTHpfEXpFvDxIMjLNzL
eulLww3dzUGyrtm16nmjvFiWvo38fPZo3zQp092QLUkh2IHoyAaDnI7ScQb5PWfp
3d+NJNuOky3vNnsWz4wWlZCOBFpgWyISJD0iEtytEMvyD+ckWNkKRWFyoQI6Uq5U
kxSajjBvYmTiflx2R6x+pnxtAHaE0D3ZxOwY0YYIIwgvhhkh5pIsW2HTR8xQo/Gd
yw6ntK8YMmaxOhpr30x4hCniVs4PVz4BUxRzTZ1Onc+P+ByZGxNTVfWy80gnf0tz
Mi4kQcJe3XLYPCZIZq3/tKdPK2dmXvmLyiO5IJ3qa4lGM8k1F8iUEaviogPY8XOa
ET303Zebi8YZl55xXOoD4Y7M7OMbWCuEJW8ak63dWDKRRmsGzCluN8SmCeD9N68b
N3lzGqgbtxAiGEgMFV5Hg5XVfP1fKNq6eK58EoXUY607AWO5/S5ZQZYvC7zfA49X
ZcImks8XO/fusXTkZBE2RZE9r8NydQuPC2xGy2g98WLszj62RQ89aa2GkrvQzhem
l2RyvXAEvSGGSWJZ8YsLkYIh0+fhnMYxJlQd+3bVoKr1oZFbcwQTT1VgO/nvNyJF
PLGzNzmNe/J4+vBH37JMjK/GHadSaVchxLvrCnVeuibGGVl0vU3/2CD1gvVf76bG
+XwDHQbrI5tRpjY7VzFPTb0J/QgB4G2QxyUu4K2l60myfcIg1CaO2UxLNsc6K5S5
hg5c/MR8Edtz/q3Z9p5g7urPyBVbc+2xNHaUlGLWdqTDX+htbZus5qo5cSAhFqpI
AR+6JQvdgk9fQg4+h8OMA2CXP1RRcLYsqrzIJvpQyzbTU96A9Fk+zdc3i4ecp0KE
IV1spayc7tLG749O/YE5sHJ3CelQan7zD3cEMzD5pE8jhBYs8PTC+fNIodHC+n/D
65OXKifFmGeFA+RyQQjpFwnzVQGGCUsMnrm+Bmx7vZy/zZFiVjpFZG6E37VUDDSP
sIVlZgekRhyH5PtHsq4RzcSjx8JHN1FJghFcVI40+5Ob/baEdKJoTIm4QkZ9d4Wk
0GupGNUbr+rvyw6SltYUkJa5Iew2dcc1dbAC5YzgilhwX/LqDzw7w+dbjcb19YWZ
R7yh6DI9SGPlsGx2hcLK0W0LLWlozCpM3qHHF2A242qGZjLFM/lN9vBGsWELddxg
TCWO3X9mK4PofpV6vYRFgbrfuUiReAkAKjFWA+5FgyQV9JSupsg8J/kJf8ZU3J0S
zsMMv/w+uzzmqlntTrlXYKC8/sLhfqIx87jMQ9DXrElhnIMNtIS9bk06PM2jgtP4
sIHqGAx2/C50wTnOBvBmWqyABsKXXmfl/vMtp0ha/Y8+h1DKd5AuQBau3yGYkRr4
XfCqXxbKdVAELOtCWWx/UjQalVIsF5GplpUjuBtrh9ED5b/oCU+RYnL+6UqDNFoI
82LVq+0doqwVRasxBZEWEkl280lt4XSReJ5A/I3xGgBP/HVQ5jYSw5wK5FgD8tsl
NkIhPfvsbu+c99A5a53vGnNyHrCgLHQYTAx9gFcpXlS9x3k4hgXv7FnuqUqdHT61
RHD8X6AZKvHA+E+22oFc/YQ2Q6n22DBOjw7m5XBoYsWyTwBch16FkHLj14g49avq
OsOzMBUhsc6O3I+tzDXQ7ikmk/eJBm8PCNmfz8FvoSx3fudjh0QgN2BDof+64DMD
zEAwd2UACktr++NGAJ+VcMErzZACvJTN3s6mRaREl/FOYDPtWtEt9bhxypWIcqjb
U4J2yQzTJdplvxK2+zZiCTZbM/xby4KX0vRRC07RmPKFv+J1ak0gwgceMNZ7nVWa
wlX6GD+0T2E+DNVnwXw1nnnGCeZcJYL0dTeRmOYbAE0fFEjtyBgQYklI7cNK0GFb
f7UjVcdiNvvvIZ09l7M/ejezq4o3KN4PKvShsRDt7T63qMKJA3AAlnxy4LU3h/Pq
VVKo3xVSUVdgLkWBoJAmE2hXXYmJKcuj/B6qmBXjETPjSyExYeW0rlUnjIkkXRkq
FUGljXH/yAEqQUSf0fgBfvWyPbuqwkqCd1E9Nq2dpBeAPvCOizHC5IEFhJ1lfRHp
qZ6MmmYnbBwAR1ItFAyz/vigt5xBgi/tZWmr4QCrIux1G4+8COIU34wjOZENDj1T
3x9IS+Ml981sc8tmiFJz4hVu+ja6nv/lHOFrrwSB0qwMmXr1phRRokHcnXOHe0k2
a8+t/7dWpX3gw5VzwCW1SP++exEThjPNOqVEZmao7shwI7zmE8wAmoAJok1oTT0s
mUkjVkuCxykPKqy5yZDB/bv+lkBpf0jyvgLqlBm9LA93Jg5EKLOHGlbxlTwmGQyc
yGmJ0NYKEo6sfiIqCOkSazUSTKJFYypGGvhWJjHUUDgLnuCKDFPtgpX962g/Vcy4
HNtvzY4puvClvj9Phg7D2rvYBuPWUUlp3b0bqFRhXr3ENfooCthIaDh7I9TS9Ikd
GwZGEwQV9hIomo6PvCYlHbuw425Z/yyyRR5gaA5rcjIJ9eBf+jjNvZI/esWiD2n/
OD1O3mIFtRf//wWZ/lSD8MKsRBlGmE/eaHe/18UBwcbGOJq49JwVsUPMWYK9IuOu
XS4Yund/lK38LOBdpvJf1pgU+iij+rmvq1ZTWv/lxQNgbDYemVXASFUJnLIrOS/c
ZD1zqU1aN9mShM+QE4N1lbRH7A7DCKvTfHsXlPGBYZOrmMk9bbpaAJUU0uA3zBHS
GF4Z5tp6lvMIb2C/LGMrEScppgwyxHz4MxEUmwLIhi9C1+Weeap8T1r0ZhN+9qID
nxqW1dGJjsyF7yKQv5X7L3Jo/rRyeIoevVFcOmCZASIDsw9P4+L2/UdBonKnhJjq
VWDhVyZ5NqlPtQQYBvxxdG973usdMCDoAp+cbcx9nzz28pc23WmhqpUwqyv3EEsk
MTRezfTUAfhEGd2ZdLCSosVmkKP7+ChwMhZLFLWeHW2RiLT5Yz8HyNpD1yJtOBVh
I5UQu0PCjOqJN3ya0zoMgF81qQue/ciRf7xpOeFBXTXcPXVTvlVuaYLme2sq94md
pRA+R7KcO6sCuc0CPOAJZNhfa0AXbo/I3pG/lh+jhjc1JTuwSGicOgz1Ke19ImLG
jbuL0gKUbPKdKgAZC0T9lo62nKbCuudXlGCT/uuJlt4NAfrwlZseUax6cCX4lYVi
KmO4miljYNig1hO8sPeiKdQEE+ixLVy6bBW5PJ7v+jNeWm65KfUjYxsGcV+nPBe6
su1jAvTIOLTrVnOBwZlX7FVBRuvLndaGekYfpeotOAE53XH+070pkExugX8TlEv5
+H3spi3xlsjGYiADWBj/2lEQmlqg7TlxihVWLinucPhwY8bST3RwM1PBBq7AxKtd
l8r+k44Ck1IwepQ9C5KFrP9r/j+iOIEeYiYk1HJ8cTVHX+DbiPe6OltC8ww31A9E
REiSN4qTzhULOoEpaQesv696U1KhJ2bxLYacICi4qp+MCBjmdASdLaCCcOXlZJ/0
1D0n3V6bhkzbZEHLas/VfGhdlpOj/wmHCn+CzsascGveeaQ7Gp7N87Bgo4v6S1wm
R9ThcKIwSCpFJ0JBM+tXQCSdO0J9SsmA7idAdcLu65enafe9Ty3TxkfIt6bWfvto
GJszNcopXNYsbSebvjfmi5YES+ySAt+l3SNVdF/tMZp/3lITy+N56D5/t3UPG7h3
noMBE54qh2jCJBJtQEVrOzXkLxCxRpNfunyibqKtyh9xWM38puJTMkNeJCmxmRNz
jY2RUzKHfUVapo5dAinuPCVOyinbyq2MK4hM85yGtxyyNISgZpjPsPjsM3OS2zGo
aGcXH7/O4gx9IQDnPodnevv53thLFur7Bj7psCzH5kyTuG7eG48lCrVnIFy2cf3m
GX8vAQ2PkNKU2tuX3EOGSHWbe/WUuLgDDCgMCEd06OCR1GbAZASXT/6vt4KvH5/M
A8M6g34pIeAlMEKkV4MlIRdegGDEiCsZFen+L/YExGgN6Pkt4tcxL5/a9weiTZLi
RsbGYyLFdrmqSIjSPI67Tlmk/nvwQb3uyDBLVkuPRKoKGg7M396HR84XAQTItA0F
F5yjpB96oxOhb7CarD6bw3xcwZRJMutRx20DzrWVJDt84iV0mJXKDPtf2mW+8Qv0
40TKIeXErXSTX8jDgm7c45xn49jwekEnHUyk0E9P1qkUeNNa6iHNZhZRBYyV36a+
rF8XfS61F2zL725s9hW9E08+Kf/s/7W8YveydqWW/BfEHQwe4zngKodGmr3B63EQ
KXdF+GDxY4nOgKFsuKZ/RVReG4Tt01KkaulwaBuwSBczOR/DlePW6LDiJ3LtIQ2b
O0vYoncUkWKkgaPYu8sxJaQepHK+56SioPoDEWBk2CBfKx8zfOWDIirmn27BtMoq
Vws5FKuFE8r5l7Yh+JjBDKFNyU0O9w09cds9UkbMvijkm1Yx+EfNj99jy2uYe5al
b/RLIHYJTuq+oZ2Gn1LKLBqj6MhMGg1yehyxw3MQt6WfpK+QKiQ2VX2brYjVXKOP
EwcBdfltYlWUvxm+al/P7JqAI56TCVEc8yRtxaQqaK/YUNToNJk7aqlRDxy+F/lW
g/oKhmE5/sFPbYoTgBEzVkqkTDHnxE9Kgylc/VSV/cliqCI/hh/M18bIN7U21i7g
QK3m/2og2c23Kfshk7+i6xdALsRXolA7jjicegnRQIcAzwzl8SnAc1kFgXsBFzZy
AWflGyv/c4yr0OxTkHOzr+5+0bBmrmhpqSJCoaOTb53RFmlpxbCotFrpwjMgMbsi
As+wu0QKbLUbidqtJprlwRKKnGDtMI78/Vg7DZk6qJpiqiM2qD63z60rSmZ5yQ5s
6fUx2OKtYI+mxvwA0fKcpszi1uMqAuW5/LzyJgay1Ovun4mMUEFEuBPtyfwDobBY
V8Sg7/xDzXHWJcVdm6IFnaPmuq7C1lLRIinHTt/tC0GKsQPKQYbP8VE+k/rq7dCk
KYzi2vBbbIrI2szQ3TSw7cT8049s2GgVp6rwokJu4DyZ2fuNhaJnHdC9p6fQMlS3
nF0k61Jm0iInCU3AI/fgkAGf0D9e8pEMPrCJo4xXRLpxu9KOX2//Gp1LN7G+xWc+
5eQ93vCV/YnluyiMnnoaDS8BfCSP00N1HUa8+XGshTR5zTPeH1hMjQj/0kRiJVTq
MWh14vSMo3XztHGoZg+BnK5qnedxRHJxKLQgx9DJryyLuu8X5IY1LZSpSrva+nn1
51HrImrTsfainyhk5SB+o4UoP640bORRNTCi4SAqDTO2OeboNBF6WHg22buz45gq
uU4P4YIZGvDqjvhYSdJ1OR9tCA6Ez3D0kU6VE2e0Zvo4r3mtM5l9Dx207zlCsBlQ
Zf92M+ZELUJvAaQGxImd/kc7TSm9/vjDmJl1+Xo1HYsX1qQyNG0VFifSndfgXNS1
TTHcJDucUK8i+7F4fwP4yQCJcHRdIvO6MiKs4mrGjGxHygk4hmKheNjBei+Ukyfv
DHPCuEvsZ9RBj9PV3tNKbVF0ZNSAldOIZ3cvHIiytcOTfTBaXOfrP/RDsy0daj79
bEx7VRb16L6rRVQyknOmpCkiaQ00TJHrQs7Jtx758QzgPKrO1vRnIg5B3uip4gnP
rgeunV+6xMDL5+ighM74f4q6VDtiKL70yAkWDksJi8X9ZULve4IimYo8KZHAMuYF
6KcWOnDoUdvvBe5chQRerXKW3J92gDe7Rn14bAKhDhBXB01KOJztJrGmk1fZjWKX
n9C+SXTXKNCDSEEE7IcLHqQKRF12A8mRix5GjkkS/zOLQCWdgX8qUUx9ouBHnckZ
H/gms0FxJh96oWzos8XSahPsECQVw733xFiyJmwwTUf2ImtHYX+dBUnIWQl4BOzS
fEt23eS2KSHfNtuBQubafbmhVUFYxBSyaozTPtBD8aZl67zxfOVTU6Q0KU6OxC9q
r1Ym+ezv6N0OXQuC0ct07ZvFsTp8z5sXDj7bVOK7eVHtfrsbNH/F0qwvL4ZlyRGM
N/qBVSA9PA/95l+aJXNVlui3MEkX2bjTtDV+AkfVtP4BUYv6bP8fgQqWq8OwD0eI
ytw3qx9SQBtSSRJiBT7Qjf9cA/p56SXvsLdgyEUkOy4vv5n/7sPzoeKzeGmZVVEQ
m3srau+iqYvM3i6UfDYVUkceVAbteKynkenh8mMeEpSOujPsuGjYPSCF06fGlxNr
oAx1+wbayeneAQ7z500pcKueLiT2gT7t9O3v67hcrlF9+cLpbN+rea683XbgcHAf
k1Liq8gY4DiamWGQ2UKU0BFkNhHSwUksDvTSwjleViZMSWjJdNoxJ9jIRrlVnXO3
zSHg5fTERq3ifue9519CHOybhFDLf0loF+m4shkPELEk3Pddl2iJTaZoec5Y0I/k
ht0aaD0Eu0GP8Hu/LnTa6Dn9fdQO+xHxZEdIz66oBWYO24XQOdKYRu2s64MqmWQU
vJa9A/U49ijcigildHwvJ02Q9tVpWFmDW6nJhTBwp5Vra9qBpXb4QCUXqWMKoSiO
tqtKcZjPZFqh7PfV/Kn5lHbFZwSahO3ZCp+eMg34bVMKFzwQH9e7fmqGETp/m44s
aOcTmy1HoesXd8hdb9DvwuVVWblAE+uSFmr1u16byOmjKE9ynt192Yw1HFRmT7ws
6wLBaSZPXd1FeFhtlG2/HX85/WrT8ljUK0VVXvex7fdR4sqiv/CHUbzHWbFKDWgS
bbdrC4xKs4VEODRJXUamk7f9R8QlxcSyIICZmcNa+0db6hEYXq/kyqwMkcaeE6KB
w59fL2rgggIzAXkUPU3NZuIXsbMH76o2pcvGrSWwrZCKb7LajSLvjpEBj9zfziRr
+U0IVb2U4Zo0FzYE9UUpNhaN/rDm6gcBqKwlKlD4oV+xAq0zzXLdAmlxGQYHzH+5
v+NafPkkC6p2aVEAy9F6A0wrpW51+RftmCh1wX9mOEccv3DsIfJRU9MzFcEdUbRf
0bRunDnAErI05hB22LhTZnrMndx4++2nV4j+o4WLqbZcy+S/eLUByWiOpwS2QE0e
eDjiH39OqBhO3TVAWaf6Q5X5mWFA64r3HJon1x04bWuKjDbtR6UEYkfcscXvqLER
1Id7Irxt2ZzElrDsbLBcI+RU63/XKa6fFVutH5+TUGoKqUgvvvsX13WnRSLEq1YG
vfdlOM577Oo4JdRG68BBr+Ri0p4Qeophtkuia5l4ji0V7D/5iqa6W15Pt29CNfLG
APJ9/R/IrNH6GFlgTtj0p9FIYN1p9pbBsceeaxKnEgD40ZTYsCmcBD23G8q9+45y
ye7Hn7d3lUnzmjdLVtYxOFP6pfhDunifRwOJFv8qUQGJfWVQ3iZ1YLoD+nOIMss2
Qn1dswLFrA+ahVwBpdfQL6uMU0NUuPRKzdtbtdpt7vBNoShNrRh12AT72ATWe7lu
V2fXrXsY3FWNoRQe2i+3hPPqIwbXha4weUTuuGhalihSpuf86xf5NlogJICkTjyn
ie70UMSsMzGM3mkTYTWIHCnfc51a3Wi6INKgabnzumHU3eGNJAzvWV7UdrNF6WJb
dqoFL9/tqT8uDsX7XB5/v/c1OpEQ759AuJf5THOMkkPe0o6W1ysfogw2zA5rhjit
8O9cftBju77XLRQcBPD7lmpUugKM3z/KLKZfQ3gR5buJS25G5Qx90gwtlyOzsxaw
EpRuBGBy7qqQpRo8o9nTJMz1NbXJjxBX3w2Hr5hZVA2ZAYzU5llxMXmRcL90Yxea
PY/YRdfh2C4mMmPw4+nUPbcataYIfAKYVJuC9SKFJiif2Wm3FfBwrJq+0FlXYDO+
ga/CMbZhcPpNqGbe/YH2jJUbuoGtmIseK9tgHlcfwjMjuj/R6I6kMNb9JC350DOV
Z4amjU3cCcZbXBM4fNRXinSg5wbOv6kMyFzXZb2RCMHMDDvnZOO7SGK3Uu4TSucv
KUOxw7gADQ7/e7tAiFb1BbwXLhPdekgph3PZ9MgbXbmQV9A0tfGMvSybzfhvD8o5
A/l+d9qxu9LdtImK6S3o6R/z1sbiK2xoKtXA0tybQzHT/5EJfjLYapgyNmYPxOeU
IVVphRHjaRS0ZkV7gElNQFZYN1mCDsg6f7kmTNR/uLJFHmkDAoha4Q0dH20dJJY6
L8W+w2YRcaj/6vWDRenI1gwwyvOvhT2vdlazWocoAPVj4pbG/mrwllYIFgSIg6if
d8Y774xtMMN/IZDxx8urCv5QbqMzDxn75/h3q/NzelNsgXfpw4u1QyWBhjZL2z/Q
08IB+8AC/frxDoULWtlqNllidDAVSJ2LhbdY6rdI91vprVq78jIa2NXRt8tsz112
r2wZzgI/3riS1qjpQO19Ehr9Bbam6tml79id2OvVdheZuAXlzmWEjG7kmXeQ5tR9
YJz0mzrmue1spri5XeDe5SX8D0oFhgtJUuC38U/xTNUn3nTIzdXLHD9seQDiFaMT
3mCZ69Xj7c5xSjcy0g0jWSI8Kb7W6qpkYwjTsKtFwuHmpCJoSFr4HzqxTycxGb1G
pylz7AhA5qWXKqCj9LEQA1s1ARkji1UWb3ygedVrFBLwGWbqMxGcFahuF2rVXdyz
rG+VomY2nOrRFexPEPFouwkM0ZT9Ak0P/I/3A+tfIpaO0G9CH22WVvDAPzw4GNtb
MQtKZH/xfDc2nXpIwPlDqzKIfQdltkePHMQUvOQZziFXbdYHNSIoSWOytvFK0kqh
4AmJLYKVRLTt8KMRV6CLffWuUnyblKEEHScumnZ+U4TN2B89pvfCexO3rSqiJ4qD
N7xmwhB8HhQtrUZ+vcdNiaB+NhKhy08hGzJ9LZ0giqUnrgdBSCknTfxFcIDSaYl0
dGdSGQzB/9zNGOSDXb+a8qYSx6emcQXIM3K2dc/fGDHvmDfpLyWwnmGRecxvK4za
nFtfopDy0Mo1AdE/C+NCm32+fzXNlt0wXO2NUsIYvMCkZW17lQdWmvdAuNRiktck
5mBew1qnWETcq+uHtrXNrfbuq9s5lNZSQsB2vmH1gNIrQ7EPuaC/TryxehKI+skl
X2cFPhVyXi2umjMZeBtwGu/5u+8N1vjjv6/xUQ5t6Mu3fidU2zHCRyJpeFRUkzr7
oWU2zsl7ZF/MxK73Pbm2aETje+XlXDY7qHXSvSpAdkvulEbkZ+MrbRe37MScJpsp
V23OzMoLffkzHwd4+AVGBTXO283ZoMNlUE0FAWxnA6g68gqRTL+bk08H6eoMVj9I
CSMnCqzyuf5OKI2UufkKi7pXvbfSv6wsxH0+z96C0gdK5HBXXEIpg66XBBNuQb+c
nz/QOXNVp8UZr7HDi/41vFd9Ucjuv/w68f5GHNioxyC3OU/q8ZqMCObTlN07y1ZY
vfFkL6znfRQ7IjKruq1zvAF4ia/yC9mjlMEoftNpavJvLAYKZso/y8CQNU2kTweD
z4jo5p6FMJfUbBfL73qWrLpqhVLyihTQ2W6zhDHYv8weSztOVsRjhaKAsOToWG3p
75J7nXCk3rru7zge6fF1gwLbCuPo4XcQiMFGw6kXnMo6J+NfZNYjVVFEpb0x2+0Q
YsG/Y/410S4QRLXHUZJrQYl/gjWZtwx3S0qllwDGHowEYR6XaXVK1rUrfZGXbZxW
qWNCY926gC7kpBPuj9QOSTRG0xuG26bUTIlLR10SEBomWzcHJoNnLs8bZLZa62nW
wRsaIbMkSAOBai4HDT2IylP2QluoLAoLGDGL3YbLA6Ca1beeCcWqCtiFBMz+Lk5U
Z3oG4zwC0p+uZgFcVxxqUwJsbxn3P3YOBCSamAyDLnmyyzwz2jhO6bG4Hx7BbbQp
WaXFK3W90nexm93FxTMJWKtgm1TE36foi2S7iyp2IcMFwNueToin+dwY5eKH//zO
8Llb+6ErlpHrQmwL7Hb/jgfQor6z+zYvtbgl88UKlX5gekWUs4bqeRtHXhhGDcs1
pyqx6ImhQy0YF06+ImKyQ1FZP47qJMZa/4JQEEYheuo3ulfp8dNh0CldXqEvfx/4
CVifgioGN0gF35J20rNP12NRADmNDMYku0xpQaN/AJ6MRI72foWP/mZRvdeqVWs+
twOb5fAOA4rIwDd3/phf0mQN7p36jakezca0oUIRh5T+v6c13IsemqDLUMFUD3YL
GBYpQVM8vuLcaj7RlxV/w3ksVqMzTb3esxFfcnzD34oHf/p+BjgWdoAOCZ6NJ1CC
LdSeqk0KOxjO48EHZSzCrInqxQXVFQuSXWZUP6YiT2dIPXWfKbvxPhIcm12abgKN
Co+DWnUxX+Fp1fJYxW3Op4aGRKz3kO9E1tRv5mIDqJq5rvkLBM3CU4lJX3jxGA1a
tntRjBf/yqrlNzd8ICyE46h0zD7FOo4U+Fkn9/L0a38qfT7gujDItVohWR6Tz/tE
5smJR+fiZF8+AghaymNeascEAFj4DNMb6sHjUwMXZFX+WJEI5E0tJ2zRsOc46LgO
bDSKqsabZbZ6+/cL3c7+HD0XiqNBEmp0dNHkgg2QEcDRYoId4bg2z8EdRY5Kmmhi
hUTZG5iXYIIB+ridw9ssXwOlVm0Sle3ahUdo5Km2DZJtgCOtyy9v3LRieEar7wNH
RveSo+7UIjg9lO/Nx3ReaZIOT8o2GUynizB6VfAa4GPHJE8oLcQsqGz0VMfshdjs
fR1M0OgNnOQYUTWRBvdgHq4HCxlC1dgxd2CRxR+F8Zq6jveZQ4zSkJlheUKcFZPa
e2ZvOWjDt55+sGygnfhiBuqIo3kQQuy5ZEtDLhQ2DW6QGrLTjvmIyRkkdac/n108
w3wBRRHMsYaoeXGfc+x81aGtSz4dMFn2TWcYTwmbWf5tA/9+UBLTR+3LIYmag+wd
jMoFxsVukuj/ifF+7gPy6qc8mJFLMu8gh/b5gTJ8q+J6gnM4uCIixslxmxoTNMtS
rEqan6lNmCoW26tcmZuM4HvOx+i3UY27IKXqlW1q6+UQbTaqkxVHwRD5WCFafZx2
9vCGBZKkYDQmW18pDUULaguaN3Usd5aeKszVv99pGPaycu6iJc3YncM16V8f4zCh
2TxEa8Ll5eucNxZjqdx/r0ymy0Pk0+Rnb2WbZqLh22aCfu+gnwA7akA8DjAfe/n5
scZLrUigf360v5dmkQ5w3InGBEEyTL/4X99YyeM7CeZ/mtgZomlO53XNj2mWRRfU
c4BTinXbsiXAPS8L6r2y3QQx1s5YTnZJ2OTN1jsl2IGN6M9BoL0Gc+dcGp8uvle5
aeiLsdSlzhbkqTPRE9rkeRrPaVsFVhhCjNcJO8am1KlLLXijWVinh1f/F6NLz+Es
JTnPB/0JVNIGBnl8JcXO043epNe7ULBuzSyJbWdfdp/CmlT58KsNy8IwHz1bpwYX
0KORtYLnTPn439dxkdv5tNR94TKwV2pAuZ3v5SL1j6eHUNSEVom59K50me5TQ1ch
hgSN7rm9k0rmADv+SHhVaXRgPj4w9pxauoTIOsP1/OztI4dR4XQzwrcbb9ZuGBp/
aBdl1om+1WdOGWczF7RYZ2XBszSAedJ9GVO6+w+7UD3PFZ1Si+HcYTeo8hAAdrzb
JTgS77Q9v/0LcJGy4f6KqMebLKsWEPbkdCv9mFNcKiZURcXfLZhq/wc5OzX+wc31
3oRTpCfhe1GJd9AB2TVcuXBpix/sYiLc6KQB3uuDGkm7yggsWKf1AIiZ3I/rAsgL
JMSc7B5PTuFwhdTERJl3NxaHbSFYCGwvxi3qsdFEGC1wJrs2OdUOSjHtu7zg8Fji
EyjxIvTvrNbx59s2CKlto+j69VtneUsbMjkF449lllVcc3o05VXoxWhb8uPCIzgN
jGd8DRtyzFU4MggVzcA3gQ2925FPawvA4sbtpLwHN0iRWIVVNlhMFmoT/f1wCmWL
uFqzChO9UD6B9mRbQ/m0hq+ocL7SXV3Sb21rLVxDmNbS5VjvNOQWD9sk/rTCnOkI
ntomuFpotqmaAtNrU7MvSpLJFXGmDQXj7CJU4QeC204c0l0HjbnN9Zm2W4heYG4R
4HHVDiIjFRrZPLAnKRLdnF2+X7PystxkkZie4yX6Q6pm/ROzS+CESEMz8aUtFaoy
Rwf3IPOEdDPMf6ybRAOZ6w9I2W183Yt/NC6rzRLIeCsngltOkdx9iXaXuzu1F+iN
/L7pqJXJYwFAgbxewXj+sGjlve+4GUrDB6fXoh2+yBsGWCWaq4SpuUkJmIl25le9
rv2NFP5MFSk1qfGG3qSmq6Q6J/35UZEj+0NGFIxkMEC8WtwfL+4/S2XhpS7LFgyy
HyslmxO/KwycGQgDrmPq/UlvSUq/174vmx6e6tKilriu1RdqRP9UDaIX0zZdxsGA
Y+zcvWy5AVdOxrkOs/cYt+w+wxxSPLmtLqNbeVdAxZM/8BTHqNdvXs24ZxHMn7hK
i0iaLt7vF5Hg/Y2ZidK8yRoNRf7Ci+TVkGKQZoUgNzJ7bGkxU9UFtA1V5I7/Vzho
NdAwy9q4PobEmYmYL3Al8FqV1y5/YUQx5ez7aUS54EsLboZlkMGFxnUuIVbgtSYC
2VqR17tFyoc+15HFBCFLakmt9PSysC+JUVEM0s7KXFvy6/jwhDRxF7T0WmWdQY9Q
t5RXHhTMyjyMoepCJa1a081HH7LnhCbZBb1wluXYXR0WGRSJedwUCU1X0/VmpgeU
aqIWYXDsBRyJqm0wDVs+dAfof6X5AGcjcWPKMR/CSjaRNNf/iViXUfShzsMslURO
IEOgcAEdy3YlBwGgT60bBUWvuCy0VwGY9ShBQ3eq8Ce3602Aw728vp3Rg1ZYMK5e
wPOTjAKb4vRq9P+8TAvjTdqtoqtjgfZm+lTV0PiGs2W3HhTy0XSAy1qkbQKGjLo5
XCTF5RGU+HJUf/JW9hgTfqfTvH1wxAG1nfBBoV6MOmkS1vzf5k+6UM9qXqY4vFn8
uQINNa5ZHuKjJPefHcv/vUE6ilPvnsmN6WzfVlVfmkw1yK7MGHyzUypzmVoBMO6x
bpaeDLjeAOyFuSr9pMfGU6kRGQmHqXyj72gM8+oDpQVVSquI33y7hyVkNDOgKRK0
k2OATFIA74DUxFvdpaWrYOXTinxSY3S6d/SW8bpCnrqjH5b37APWbos5G+sAlkT9
np5ikwf2l+U9CjMtMb1h0hbTBNbPL0zpXVDO91rAoFBrtvnfrQ146JpCzRq37Gmm
Qsaelgi16maPlkO50z4udykwSehnisgf4w2hTGaYOWdfEHHFM57cPBODHt+QdG7y
y2ITnFA0+QA6gjXoTJi24n4SNjvgtfi6wueMYet/8vxtkH2/Qzx8f8RIANIDAOIo
/jTAry5dscehWM4u6gERy0cyVsvrc5OFI81AEcCS0n3k+RzHHAqML8Y5rhtvDnl/
bnP4wRNN+L7SASJo+LmztFVYNCKjALGLZ6C3n8BnUqFyNoPhsPxyYblceBnxfgP5
AJvsBi/Fd6zRWuWak2FRFM4EuuTItDIIHFq8Kx/EVjKGH8XYY/W6jqaq7ut1U7a9
ONAngQMJfw974pcl9DJSCavKTfFna1AkaOvMFnYtjXHYEIzC0s209CKfbT5VlHZq
fY9gFTZuteqlxkZU9tSWtwevkGWBhhQxF64rRQkwncta1idPNuMQa5yxFqeC3b6J
Y1pSl6PC6LVg8quptaqQVDZ9mS9NWYx/lW5FESQQGgDTaIOW2leYwfTMrRKkeBDM
kjFw67TOvZQQCBOfx48EqW0WXXSGEjD/DUCqrAXAnISenaw0rtN9JkOPrBiGCsTr
ZEQJPG9HV9oJ3Vib5E5/07TIxgwClcqRepzmRIXrZEX6nPWelOk6YXSlfnyT1x3f
/69nMhVzHfS36C8qlCbUT7vsU8VuUrRmHt0W7uMqfefHB4qmAWALkfiCopUOzw2E
CmDKP0XfP2LqfXsVuIx4H4xKF8y4qlNEeFHcAXWjyfFUPS4b1CvOsdMFG9V1kMOx
rblmXSFRX8pNbKNBrBRt4EemZPjwzXkPF851eY6+bmjCpRGv44dWcRKDmV3CzRwi
CsLlY3Tc6uhpDUTQzlQfp5wxwuzw3LCDfiDhavl/f6c861IIW36hLzXbxKsDWbGA
67IAU/l5baV+gitHTLgttQZOJzy2YkGEHVpRsHNPAFFYn+P+KVAY435SuJ1LZu2Y
5te+C0YVym9bu3EiOH1KP5mcjalpagzrzE3BdHQ77nSGU51LXwG0Am1++Hipt/o2
QsUEJcRePkgq9sh1aW4MyLabLZRi42evTSUAGyFw/kyBFKyh/6DB+m/r1x/Q7Omn
ce+Zro7sN/m0e2OFuXla/kwk5nYj+9lfHbLTmY5giO4pSj32u/rWV3ZwBny+sZri
GFZ3L9FNpZaDDOTs0EyEnWKsOx+xMiD+CIeZIgJYo8EZqgkeka5OKVzgrxMtrGJN
SY0mEY6Tb8rl+zdY471njHpdOKgbMnZ/trN8NlnAcdIQye/HUc9fn0jis9lyDYeh
F/3Vu/SKlgA/FPYdxrfsKEFjhzeiNSJ32RPLxgnHTJRiKq0/xQruQELGX4fwwrb0
aoSS7GcsMaPEjBdKEcL9RFwpRtbVvKrF6haCW4OLzb0RHwviBv4nQ06V9bA/eMvs
snQT92r6rfqHtLviRNVsXUOjwthzp3DQYdRITwYIN8XSm4bxojepNYaBm0jJaXGQ
7gMwrebT3FYunl9xzP3hsOtrFiwDq5VF/8M1DKakdQJJ+25P/KNzJr4r9cW3jdYf
KXR8JecDxsWB9NAZmN8kw9p6A8qWIS0M60s/bLe4RCN8AuzkHVOG5MgY+t+tIkRE
bt2dZhrNn4vg4wj1UIHUs0IqdO2SIN9OrE6xOmmymEBM7HwBNDXP/ngx0i6vH25Z
SwIA5tzh8mJixnJYTNKfrMuXIKPZDCfJ3ZUc2ZQtCQdUozAZG64yWOuXMp1wDr4o
ICEfWuTj7NtOlJZbuXEo5xuGIA3xzQqtV368FB4P2FGInn6dfiOTJOyp4cKCIHVC
cDJtzF4HTVrlgZqMcu43aBNCmUpIk3WZuMtrNjD8WXX7qWAFV//wtyQpPLNVfD71
dfoV2vmBbCoaCt1m0TUDtDH3zQQatfLZBhg8D6f6q7wfgUIWLTXKNbFo3aDxy4pG
Vs6fGikOdior3LWYgi4LCfJZsBBaFQekklSZA7sLwQnVktDC7RRAnpDu7MmbMsJQ
TqSZSQl6nq8nhQcLl6bMhhnHWGij5bwhFyDVGvB+8Aqidx9GibKb6kI5mM9o6IdB
3P5PhtDHPCtOKDyBnjpSffAMLRHDf/QKaAaYOJhRHNTDILjevoI5hm1r8+a61rx8
zynBfX3xTHvQFoWQaZYVKhJgMJTiPXLQKWGfQ3zLRwHJ5QpDefa0bJrFklz2aQUS
3PMtMJjW7KTJWxEnCOy1zQxYuy2IWz45I/X8Hx4SCkcO4uLlwzqygeHALI7bq/Vb
MNHJ0BOBRw+a4a/8YvoGICwo/egmruPzWJtw3M1hYfxyzpSynSX2HOwfpi+O8fKe
l8vz5i8tkEthfpzdeC4s3+hTddCmYHmIL7i0IkG1pMmXaR13NWPjGoDHQrF034jF
Qb0ViLrbvT6rgf6myp7+wDxZ/9TZLn8EulJkV+Mhlqi7jU4CLJJWftITa81zGfrL
4lweogbo2UPw/7sS1BMZEa4R8v2VF9J7I1v+zofx/hDkg4WIaUKnI/LXUA3Uezt1
KZIa5kamdWz/DexTTs9Y6WDd2MzOoj6VVe7Or2fK0PlDv8yP6pjGW3H+Wfxd5Mne
dslk9/hfowGShxEZpMwhol26uF1G2WTEBj2Rxz4eYaIQwchFQvNNeTj7CGvWMQkZ
Ucjy4ZmWH9D397knFW7PSgVU0ZFX9NmAGL1tTxp1xYa7nfDWT8mb1ZUFHsHxmIGZ
S9LO0U7flVKf85uve2pROyY9LGk383qPiHOk5uHtIwGhNyvV+Pf06fZH2X5wfkE3
QaNO8P4Ii2mzKJpVg3be12DmauMac69cELYUhlX+4juWTv3tTwP3KMS59xHiCWGb
lrTA1Tb4auxi87YP116iGgxVNgqY4DrEZv0RytZ1O7Uq+SsupI5EjfBjW3ZrBGMI
Hd/wGB4zSlUJn/V0eD3GcZdZyOdcSJjZ7Zsq2A7ffrTEIsA3u8pl5L+Lz58V8lF9
a1J8ATfIMaSFlqDgjF5pZfp0WohG6zYZZXwcrdfPeuEZEOb/9un2FhcS7/zukMIG
Jj3weKKXp4UJsImpfYYre1IkwlJbnk1T/hs5cjm+qBtuXUyNFZW7xmT+kFsCtVRa
gxlmcGdDlX97KjcZFfBcUVzeHe3YA10bLGKFXm5ZjxwVbM7gpsvbKX5RQ3ePjusY
3RpZzZwmwIIdN95CWyZkUsIgqLk7Sr0lUSi8GiXYMhUbX3aFvOLdvcxTycyMjdBq
IY7fK2a3BHFWyS4rTbrrMzMRspl2HNIVP9aiPeMIy3FDE/ZvWoQjvGssu2n1ox7k
MxaO397nAZVMrsJ4goGnchiSiQI5it9jQzI6sBdlk21SB5bjCxDsOP85KX2y47zy
QsyhD2KUSyJv2uh4pysiOZ3SYUH6j2xCTTqrcE8DCykTViikYHrjyIwZo86T9x07
svInKVL27Nks4orMGUwnXPhxqL0BX/TJl/G/Y+36dwGwa/VPex6+m0V/sLbObfU7
nh5smUGBdTYlYPdbs19ewg+wx6ni45iadsclRwR8MeapEqj/URjowHb8KgMW2mn6
NQ3ZkDRrXTzPW1qLvns0pT3L+ONYzMtSUPm9ZgcrPwAvrxSQlGJ80d4ucETUaSWA
preK0KDppeYflv4TYbgkIwO6Qshq8sePWgFNRtNRupfoACIyTlFHbw0q5ZRL6Ztj
wFKALSxaGi0c+iYjfF3Lr95RUjNhWjm/fed46IGy9wjJFr6/hIYw6d1NGfzbOVab
i0aHEyXCfNzG3sJtK3AKCZ6nZCFGRWEhWssako+stT2tFKRlLFlVqV3mi3v/3SHA
p0+LuFBFDMg2qImvMJReFZ+ITAFHBhNmFj7Ce9OOCyBNBSSfmsR/sZJ14CB3oOAx
fhfgs1ITXeSYGMfTAGZ0K4tw3lfRVLjl4dtKmyAuBrAWee2Z3Skumj0S3lKgR3bv
N6BSAwM+7MykXUxpP+qDgZm8g+Inx/8vYasS0tN6R+Nufb01VWGA88vuUPvAaqCZ
rrssP09yHUvZsmM68hhvWO36c2Jv6aXK3wSY5xIZP7QbZXnx0ds8Va4sWoVTHIxZ
T3/CMaiVmigS86Z8rC4o+8lC7s3CPd/QLpE1W+OYx/VsK+pfo/mQ0i5uU2rRBcFN
cfD8cZAlL+BdD4/I5u7XDzlvfhS3WM6wQ5cP6G3JmZHHDpNSkOP6weLnm8I3qG7K
BCMoT1aNCNjufHGBsJoTFxzSJIGCMjXWjC3lYnYxjyg+bxEi2UN7Rg3Brqih7vXW
osey/2wVdcECvbA1v/C5/JBwsfeagBmix8ecMGGBS4WtPpHe8474WMlld0NIZueX
7BV9YzzSYYT8iUxWXXwZJBAgdRNC5T0EryeGaZnyPBa1bjCKSOVJOk5UPP0ETb4n
rEPts0TjxUu5hLNf0063B07XC+AE9JUwtY2EGllKMy47ISoWxxerosFN8IHHPX3j
5iPVyFQFYZGru2r4hIbngxN9qSl8I7owK3Oq9M37dPdNAJmC958Tr/2/CPH1o4NF
Jmts9BLDORVGzllxAuxdNLyqxzU1AS4EDHmP1gB4/O3SBP7IUAkO0R+9tE3whnGx
7qpOBGOeQqYGc7oeRONcxl9JeNw90i/H07GywdRIi/jBxGhLgQBtekjiMg/sKnnE
x/aGClKXvgYbMEvR5iFNJ8s+kowb1l7pCxBnVv0InB5FU0PEhxVzQ2TCGdvBLXHW
xrIEOzcK+wguTe+pH9OfzZoOr0OVwpy7VkWO9nn5nlO9PU5n3WHHHRT82ykG1y/F
vscJxI3nwNQOAA9DLCZXYocmqnZ4t0B3DcHWjYb7Zf0+yd4Au+/Su18l+ePPec6P
zlDxbQYMvC57jwAoWupm1oPDZmWTSQ0/srSRZLx0R11UYPHf6TINsHltFuMiBNeE
dmqOFSyxPQ99yZf2Ha5/31Br0p0iCFy2wqIR6+JME/fLZqga80fClfqyMylVW2BC
R6ZfAe+u0He1IxDeFau9NEMrgOQayhZYSxfzHH6xbAh0RzDLkkOGrXNr3Ccwa2fv
lo665hXMwfNdf76jazKhQG91tT1qsk5GBxprvVfuL1wE0keLk0WHZI48NDeXclRW
eITXbh3l09cKsK9nBcAV5PNl1Sqn7KYeUIJxTTYgZSjHZmi26dOjV7ANy23zMZ/T
vxtKkDL5HyijVncQuFKw8hgnBAO5iVpJ+suMwdkgkVMasNi7ojh8nmKUnMz+TLQK
yUreBjltMi8ZR5vyoUqeB107jA+FqChwsx1dEVF9jsz4M7kKSRM6DbC0etaDL8m3
cRUWGOqqdC5J6YW16K0AM3jbEuxhCjmH6cmRhFnAWb7yM6mA/n5uOYGZwSZvEFZk
Ccx8VTscXlKKcsymr46MLPGwyk9W1R5cXo2sUaMkvXQpJ06wBhbXniKJ5Hl1tG+b
6WnW64pIbLq57wkpHuyfSIaHH2wtXJUlKWHjIJqw7Zdaw8Kw14SqSqxoRIT+9T3U
C1RkO/85NSd/HqG5cn8gHs2h76HuGKr0algmrbAkDJjDyRTG9L4qT5hLuBB+n5IQ
pzhhaKqeVrnabooUewiaGx/Cba/93/jWCVHwyUGIK+erf3ond/Z5KYUCd42xoaPD
mSFbh5vsseTql4pNklCH8WdkqKsyHLkmfiRBqT1/ubBIXua36tLrxt87tosFa1Go
NuzXeCoS30nfR3uZvP6uG4U9lZzfoco7VnylKUZAhwaReVSonJlA4TXFPMdjlIUq
y15JCVLuqQi8WD5aS5uyukyGVmryZ5/Ii8zA63jnZUAXy5ygHvt7Rr96ojSkCbbJ
hphoV8jY+HW3BVrnhc/C3JfHhnqZAMZ7psIDGsfanyzoieix9q4TMdJEml2MEmux
QrGkGtDgXvnAlmJof1bA7WbMl1evxa5/njb72eewBPxyHtO0gsX+CdLVTD8VN5Q8
8QlvCDEGNvzPnN6LGC7IwQMlBVifaHXMm0gqywB7yA6g3IE0VEmE3xggA4R8A7xj
GM6SSkILpClkgG+mGIDan/rWnkH/ghT+F//h6RsqnQlXmwvEo/6krPHciY1ABfoF
SQKkZPKRt9mVUq9d5WnYo6lyXYMoN85e//YTLJTNRE7NhaDpxpVp2yni3v9aA8q3
tREeIU6cSYSTQII2oeAmVI+vMkX/xW+vWN6TSobAJteUhmuZ/DIZqIUEY1C+U+cZ
DE7EKxZNLdtUSK7ipguVaevxvUh8pUeNidWLN2SRzQZfs9+Y3kL55Z+Pe24odvmK
ar8+4RZXsvUSuEXA1tWSQRPOR7MnFFQaulFajOxcF0yjhOlCoeUZFET4bEKE/3Sj
yd56cIUpMxolvwx9PnodWTh34r+3RyjMRsWmZyUY4/bvGqGDzhJDm3GB/liGDaRa
okpwJRJ2yiKL8VzfJuc4EUZvrTynd2c9KaUVrF0H/E9Tx1k/a88Z+9D4hzKiz1V2
WjUEU3zJsXS/CKxKp3aj+nR3WgAAUUfoMz5jVyxNeetFe7wPVkfrXaiOPbZ43Y4+
dm3ET+vKBbnyHKDppW12ZUeCaxjQjEkSX3s0NlrbTC+tCB889om9akefqA3hldYm
Fs+HjUoRASsjJFtGVdMuAGd0knoVfinkIuLv0HxmeSo0hX9qN4vPNjA7PifoGZ/c
dMV7ox91caZfugesr9H5m+553LjjKrA9Bb2aTPCuLkYRkZBzWLn7CXRs1vU/avCe
3mSN2+FpNvEhixA35j4a6xKDrvjTlV5srNz//O7F2JcVpqGZattryjJqfpeg1K/T
Gg54w44FxjmoJMOvQ0F03GN8Ja/hCW6V6Z5U8BYQALpRzirFLkcYjb5Yq7lVrM4I
DB2HS+/1h67DOzhwA9PJ5s0Ty26XBDFsvFMHVrXBCQ5qVUU42XgFwab5K5DQ2IJ4
THEeCTR+ZRabpUoZIjFuV5IgL5Vvhc/pKiovNhCwRfYLKTI+I5ROXz/q42cnyEho
m7LwsHvR7z3uCtV9pyxYW2WR2s4xtXM25pqRF7YYMBeonQLDt5qIPSM+RoPYnP+N
4wqVr0IwAfS5yCDLH3g2Rb4M4XSBrT9BtgcIn/MErkxIbywO+c2m6BbW8zGDB00x
Yn41BRjlaQ86xXJYdfS4IZQnwtWYI5KdpaTsT4wVUqpLKuU89Z0+QCr48zTCyGtU
tmOfKvgk8nfDX8lOFP3K9TUpAAKlEgsCIrq/s5/If+hXBr9C2Tu3j37TuPKUj+zX
aYGW72mA5RzZlZnpgUuW8XN2mg52bMKUeckXJzSkXo+8FFn0eWmkLeyjhkpSgEPi
JIAi+Q5RkirVD2DLTY3LQSo9X7LD/EVOLlP3S6Cglw4wkZPOYpewGVc2TnMnIain
ozhSMV/1J0edc/Xv0pMg/0AGFHopY2u8qVVptKNxy45lrNfjy5z+/mA4iEOqaVbD
ghfoC1q4+Az7XHNQLDTuzeGPqt6QwSD19nFYd/12b0H7x/x/HkFFRComYebeV0zv
PLPnDU8Lemvm7PxF0DNpkOXmUQplquWc/FbUY1KW/vFQ3fCmocmcsFoCFR07XxG1
G+vLsoFLJ1PIDlxPOpXvheNxUWk9UGAaPTlasfzujrTTPmzEy/JTFk25lyiPBZd6
GZCDWrUO0vMln+qdI5X8kWBu2Uewotb9EI1uqZzcWNteGfGubiIA3SC5k0QQibBp
+Lwgm4jEOHYcUSgrIj2azOGY8NI+LnTuoUqoSnM+aVc7NXGLjAbC+dY1q2xlqepm
O56rmsfjgbQ3UWxZCGthGJ3rdzPPnjzeNVmelLVMcVXpn7QuCCdFgFZnD0VrkDHk
ocH93/v9glVgyo5P+DZyexQvXcERcrwycBBHfOgCIvPydTMD/+L0GALopMfFxXbq
I8DxRxuug6Gl2DpdP9yZUYO6n/1F+dgkhMzv7fV/N0VvjQ9jwmtHBiOZV8Ev3gVx
hcxJOf7bYegPN5AKACp75F3890UTdfPJkKcbUSjZ2tCGktPG744DsJGaloB+58kC
pTqglvr0psSsxlsFgEeg0fEEpfSpyiXuT+7KI02Nd96th1nHHTG78KjIKN0jCa5x
+VuTrjJte3D0E5cPkhQv7axUgRwXY/XxEBx9mQJRkSw1eYoolv2tTY4dO5TQ5SQY
hrzYajcmPnWLKc79SmP2aG697//daAkmLOxbM2dvIG8dtDA3U5bLm7MQQazFwBIp
ry8M4Ir67gdPJgqtiVGLFsNplXxtuBV2ISIWpjcREXpTtYfAl5sMnGpRpJ6GMVsE
Zh9IdGwM2vA30cotj5+uDunZinqmc/bXWx+1hAoL6Egw9tD8HXReOEGaUbau/hE1
umR/l+HthL9LlHnloMxyphFvKBgpA+Lu853eqIxwmHYELmj+kRL/EPsRY617RltV
vA/NftpcrTNvzqMAzvvX0ZuxyL9So5Hlb4S243R366f6TYRjFI+YgmvjFw1KQmeX
iG431Nflha4Fu7KqlmRLD5R0pjiiNXzvgd4dDdm2FQugqxtYH/7qWkaEp5GTPQbU
kKBs2pI+k3rjkuTBbcE7PbTfW+PYgaD9OOV8b+km6g8ND/2oNafZnRoQJdZQAMAA
87IKC4eEuqk7Y7LR4hJr++I6QOccZVToQpYMlWz1LjsDPqRDIFls9YdFsrBxxEFt
jWQguZy6GTWhmSWCTZcOaw4GJQWqpWxMiyfiX9Yci2vn3TTMIeP4xhXLhQQxAW7o
9V8Uy4qHPVsS1hRa4DxosfPVBC+RSL94t6iiXYPUzuf0tI3VmlAYz/4xFq2ENSaS
mnpYaDteyTQE40TOBj6fFhdnqEjPGq8XAcl4eveTZp35pwFA61bdssUrHgei0n+W
ySnQd3uryrf70fmgHJmZbVPnMoew/o7eiSOw9Kkw0CKG5Ho7tf8fvIOxqwD1uGWu
CAgcjM29USRT8vVmBnw5yTHlLhqBgCa7Kwv++Rsd583ZvQ4b9f3768srgS4QFiCZ
ETgmt4IDxBla77dwBeLQkxJwkKJCmRKbHoaYFPIgBVDNlbL8+Zi4ydgGlMcxV5VQ
E6C11nWnYDi/QQseJYl/fWEyIa7w+ElegtQws4bASmq3948QqB92Lq3LGR8fc4Kx
5CrmWMkH7XPr8DuPWStJTuVwJHPwlgRHER47dbBpP7gvTHSCibcs/TqqkEXM4qIU
ZdboXd+Sy3qCKlbu5lyaZhNzgkbVp8hpHjkWhwHWuxb1Ph7i3PLaQQWAov+t9hvt
1b0I1nczciM9FwMCBgK7IApkNk8rkCbgdLGWrGz6lEOsBl45JcNkhxlye5IaHuL4
vDsE7lGwu+0BuyepWYN18GRgFGwIOhKW77rWaOXR4GQ205DQoa0oJLcZS2r56E1m
+U39xmtxnfIr2Rgvtj/UyKeHiKYh82Z+YuNQkilzz5V+N8VjjDy0WNYBMFrZByiB
ASUzK18GOxEgQmWv8gLk7yxNRGf80dG986n54aBsfOgljPV14srIxTvvVY5VsyMl
m9z37AExE4fWnzSSYkb289XptM45uBHlVWjhPUKDtWyuBGPg4XduyCZK0JyodeF4
14n7UZyopqkkXub/xvSlW2a56lW8335UvYNgyFzZzwtla5a+wdIArHWdZAtbUDFJ
AxjKCeNVMUXGKtLqNT+//eHQ8mSyKEJfAZXx2iUAJN2lmMs3sX3nrDpTjUPaYkzU
ajA9GNP9GqD0Ccdu6u/E2NoA4vMEwHl6cseNMPB2Ig+PTcWKQO2mNZdsTTr1Rx8f
J8swDRxpRXRXZxZ8TzElsYau+rbVGk3gO6HqFecsyljkuvIkM/dixdGA88yr7S/S
Ix4K3qFNprI5wHrzTQqxAKLUEErkr16purAShesb6c8pKrZPh+DBHZFjNUqBhPHI
r4ntyjC1IGN00+EZBWbCHH+n6Ows9PMedjLqbqIhc5+eE4ARKQ972xheqxyA5Wne
UdvPnpklNwWHGp4AX60oeEkUsjvOaM2QV4NKYH6upT3/zVcHJdICEYYnTE60SwAn
5aGvM6WV32FklPMV0amYCC5EupxLMNLLGZbQS6scTS4bLTHL1Fa3WgM3ho1ZfK0C
VVEXa1D/t1L9gt66KlDWd/0lNvQ2yVaobB1qH9i1bj5ojUhP3vkGq1qMDlrcpNUI
JGjBJ68r8s8BqG53agXoZPKQ2LZ8AfEfqx/sr9Enm3fgLwVSvZ7ajlnffivZ5pmI
d457MTCjj0+tZprho8FeqGL7kuncl7qUJcdPWifZIe29JPO14sOSc5A3iT/4zNda
7x2FSu8X6EkP8BWreJgnfcE7X6HIBZh/9fgzxmllCdZHc4TgqD+KWrsUYYf/yIRO
UGNDdF77QnHzMxI5ifB/iFGH4IhUdZwNGB7B6CP7rgos8dTaj/XUZ7RpNa78ymFH
VYyzKMesgU0TaLpiaZntwgldEh8Nrx3zVqlutWUbXIR/ZCTPVzDEJoziaFp0fBwo
5rX1L9Hi5u6Wk5o5QgSNwi7cst7mwd7KmyljhVn8X3y6mOv+IB8tzl54GSw1OOxL
Va3B5Kjd92Bbq7bIE1iYw0V/wvLY7FYgL9QXN6cgQLtzKhyY+hISzRRB4IC+OKQx
7R3E5Rr4C/pPw+yUNdbJOYrhBTRvaAhR5dDJqaBjlqqXM/L4/BSxaXV0wgNTd4dr
Ao4JIPbrloqxHev+Vbc7sKBFfvPQHEj6ordfPIggoXuzRXMoLKnpm7+WBOI01tNc
8FDrnuwj/fAn9MdFtIUU0vBfkEhOS6HRiJx9sp2cMNuF9JOw21efU3VK5rgQWq2Q
cHLkSZ46VP6BrTxqZkg/62cPPy0b6bDtleZ9yIV0wMmAk8I1Vo9f1sCMpBmgdW8n
UwnJ2AJdh/dti2gfJOVDvbrRnK7h/d5FHsav0pRdduMVPdYLF99miMSwCyq6uEhu
33Gx0qC6QQQqs57oVuVsDKbNf1KHeJbDv+Di36oHsCIgjBw5fsqZLkS0Bk1YqF9g
Gdqfypd2PQS47hto9tgBEZ/RC9ceWo8PjXTeEtoWxMEhGD6v9uLHSy0VuI1HaM1b
7EIwJs7UZTx+BsIH3vnOUmqS3G4eVqBuf1Q3fI+U5vE0TMg3P8GZdQFBBbY/9eKs
X7TgoEc5z7XxhbNVS3CoTvGHp4F8WvbBB2LzVZfMgBDEk9CsGQqe74XK0xKru6i5
8+/LQhtGlNWQ1HFU2WgC/csoxD0PColRkxRMfVdXbL8WygE0BC9dpDUWd0KDhxEd
bMATU4AyVUIhL9Ac3Py+w6YcD6SKbPtZqsFMhrYRoldQx2UeNG2VmU5+hbkl0Cbe
Ar3+0NpgDXwmekED9hencRMulNy4c3244g182wvK1m/hNWZcOAYNTpdgPFmKDG2k
Uw+X42SMAm/PiJn+uTuAGM89cfk7obK4zIZS0D6hvNpv+q26ZAvh5ShlT94KwCop
XshAwZwqjok9x3Q9eYyPeeWOdr4Gpz8XKJD1ZVKqHCPedviyWDgP1usV3zcA7GWe
pEkLwK6EFpCIPYxPj7+chpBAXPftYbjw3VrRzMbEBMedxqT1DlxiaNC7+Ufky3Oy
S1T8/Mn7zN5lwlH+8lfb1olczYf5syvoSUMrjV8yJqnBJw+7/76Rmu63oRTZ4Rsf
YfzDfD+cuPDg4Lbx3XXIHdwcZuA1UHjZlbRrf1iLvqxkFM+a8q5e2fJmQd5waXRX
vUe7w/S5wXJDO7q9FgMsbmdpEef4VFv+ja/Qq//SlKQiZA64RYfyQ8HuFCjExV8S
8ivtReSgENlWymhPBTGd5V48RPEANY43gYI3PEYisNCNWDhnbwlG1CjVNbX8jjxz
gRf/VEJNOeDufwpul07FkNFBxFPFhpWqnp1RjbwMiCV+u2+3x9zbW/Tux42rnCxj
yEyprBcqA+B3xN5UtcxhgHbLuvowIANhERJMgD/PhlhuJ4X1fT0dV1htT2cFsDnW
z1E8eYgJLOYrbHsq+C0XuzEAtWFJHrai6HKJ6tW0wNuz1nhndA1bsdOc05UpxgDu
xq/gu/SYR0fQ/xAuh4VRtnzfAnlBrI4hLuaSkt9zKyEC3U2p/7RFVOq0p//t9aCq
Krm8+KV07MMOKAXZTDPc9PVexkgiaf3biGdPycP7m85E1kUZ9O8zGG/5utvo7W19
zMyfrQ2Z5S9IowzYCPbJXbEkAwYjOrCrNecCKTZ+v43MvoDkp4obO7htxZpVezPA
Yqf9PewTHttaS85ge6AqR2D+NW/PT+3rd8gEXF8OWKp5grC7QN4vM55XUKhuQv1M
aLMgpxv78K7goRiYQTymkJYjMj30mY6w6CmX54UJchnkX85wpwRMiStsX5Tu1FtL
ASeYplIakcKHUbnt2z8NBe/byeMJlPF19sUXdjxNPYjEB4jxYM7wwCoJNItQsY6D
LthH/TLsR5tO7lVwGT2nplx8T9zvkfFB/tJ+mU2HJeen8Td1GY2h7dwzlEsAOxGR
klfRbOEdL6RsQn6bMW7y46s4/iGRHrWnx7eESDfLFyQwHo/pYPu2jdE7PCLee54S
1EI9qCJPIsc0s2cVQmvAtyQ4cgpl1AUgbw+ey7voM/jlEptglQNPY1tiyc/pNQzS
f0FBekKJB0sBUH47mCv3s0QLIlCXUHsP0aPuYIqE8CxrttEGQFwLrPK/UKUeZGXc
bGxYzGHV31jY29Ekq5PuKd3se5Ycdfq04AQaVleS5/4L76j7I94nNNXBkqqvpTcl
RD3cUU1jOLdyxFI1t+QILUC91Fy+Fxfo43jNICtHdh4GbLf+9UZVCWZtyceQon4X
L9N2/4OLuGKBc46bHSCcdaU6mSNjdV2bzUxo0wT6ZCRmLOvM8urSR3t+twBkkQhn
oQ5QadTQxK48/lxR2fairdrJ8gLi95ETfJ17NfjgnD339MUkqcoMtib+hESwdfUf
i2TwErdlfAueRLUeIcvluIlJOFLHjVQ8OeS9+5H90nMQkxyEA+PK1WihY/3Qrfdv
DtWE5FQNa9tLuq+TUlxQDi/Biqjt8ruNe6MTa2rKbNOVR+GPxEvnUOnpxq0v3H13
+0rRvvbJr5/a/N9ip7ExIDnpr7j/aPMWnfAv5pzMMI4dAe3M7fV6YL5fhpOyaDoy
vNIUkzey2Xs+oxXtBaEMp7Hk27Tg/yvQVPuw9uBYL/WENPPaB/3nkSZfD+BBFfGR
LRI06QEQDuBcACBwQpbRzlvaLeekl8/wjLv/bL7rAfbQr0/borL9r01VonvX2GyP
Am/x7L7uq/c13PKoos73LtbETMFhNkE+n3pmI/UUR0KofuZuZf6ZDtYS+fuKJE/s
P4cjR64pkKC9G3KYtVKk96I5xSi8BEH8BRP3T2RaRJw+D7pL+mKY4+3vxGqN+BE9
0gkOAf+PtGEQnT21kVPCTnQoiZE3DVhTXcczy0wyFGMW4ud57WoSOI1Ba9FZNJjJ
OdAS9EOEYv6ftauICFOgPaTMBq8u74TLNdWUSzua3MyqNDGRPShLjVADvYcBlAY8
bkDUY0OdCV9HTK5RceZ6FEajmyhcmuR7W6bwEuxAIBqPQr7OXQPKoDoTrIMzvgQs
LvoaFM157HUdmYqdzkz5yQ5DSXOfal9R7hN+/vHxBBOYoUJkUfkE4Nx0SH+iFy3b
ROw2NiU9VFv8sadqYb/PX3bycEy3cGe5Lm0fi1DAj8AFkYkLDYv1N6GcngdH7447
WrkhZSrY1WQ42F0Ln8zt+QvAB7mRoR9oi2sq940UdipkBbn+TXlg3WPA9eYz/tFf
pz/Cn87t0tCzScsxsUbmTUtKcECF8X/uwXrNQQI1faQo8jx3SgQnH4LX3T/ASoNl
exYbjpcE5anD5WTVpmJOiTkQ2wEhs8Sn9P1Tjhbh31TQHNSSDUNyr60/7153ix1Y
yVHJFMU7bdtJpzfHV3wdx2AYnqE3PopfL0EC1wZIv+11cExYl1nXOVY4+bUWy3+b
yldR5I/yjmFIkzA5i+Yp48C2BIhW1bpjMQTaEPT2si6zsM/+e2y0F5ryuWO3FnnY
lBBj5xIuJsdV4JOKkgeceGF59bAc9PkcPklSFpw7A6sFWuEr+wv+3bviI3MSTwYJ
REDA1opju0xXSIgyB12HbITxGTbWC9DI+Di/BJW5F6IojKGgg2ubkkyuxMrV9e3G
bFpaNnOSKQ0QZvv+959L+EodfQ52jWKvCTZOBMOmoTB75wKV4ipt8Uxo8aIPmNhH
cLIx3NPdDfSwZjZ8VES4mlMdMaBxuv3TMqdQE3hXmpvPEWrdZvuXrSWEAwAOvQF2
oVfWQjCmbGLmMnNhXQPsnj8ayfBPWNIceDRQDfPoGTzvCGzdAVip/WBxN32Pm5oh
PUyF2giJtk/xV066RuwqclC1umhJW0zCgW5WQXX9OiSoMzjb1gFCxMDD7DwxK4vN
UJgddpUvxcX8V7Yq+buC8G/+2bxYe+RmTia+CviQ3Qwai946wFfPmtIsbd+0WRwG
t++HIrJ0W6YntJhpgkOMOOr91ooEwW/lo1lG5N7KcwDIl1leys9JJSKj7BWsi0Gp
Ed9XcEF86KicHvePSwxheE89O4o/kQKvNNIomlKZX7ZRR/CWHN3VwPlUUPeQXjY0
/7N9W4s5kaaQ5loWFoohG5SjPCGDEQBeaxW8+F6ZgDGAlMoXiK715z6qFNCMz6z2
RXklWszJfiEibRkmDYVzKGTiGqm+SXTLY8yIFZOsBqqK4h0jLtOiziu6aLN1clrg
scoLYibqen8QQ113h8Du0y7QglqXJOtRXNR89zWQlkglQi81QZwVFgxkwjX4gI1C
lgJTV0D2onwNBu3gH3HYXXz0b1EhBoGHMXoTPKf8U4WCdb79FxsmhtXW/1I+JTgY
mxlhwFhappKaIQ427pqCnW7vLtcSNb/OlFHFErD2NxvPMox18o5rUAc/G/lyjUME
sjDoHMR9Z61MoLL9As9Hvjyc3kHd5/jDpInzRcT2EL5S6BRUgQsmk0njBNP5+h3l
/iIJkQbcy5gEayssF0oDIIVbCAcryvcYuiurXaaywIc/NcKAMs173sk78Y0iHILV
S9Kc7cfE3hA0mOEtnT5U2Dt8kOoWaPmiFuNKLKDNxw0UBHQHvJFf3HHuOe+/bWQs
d6nEZbpyt/fEvWvKz2N/q2pfPoi2YdSE/G4LfubzcBHFG1jW2bt8TLtEu5JUKhgG
sRgcJ/dlYF8JQuQQMpbNVM0qCwgPfOL030BgSJXO/j0KMxebLeBPfbKqYIQkHArZ
46R2AkM0Idd6Hp0YMwkvrrRveZbGPBX3Id9iMmLGJk/jFMyCtwVtmLbZRR8CWLL0
3RTlJCSPMXalYIGF4qR3VAdx20RrTG6zPJQ7TlNrFnG2dVSwqI2xt1eJTrZyjJdk
lZY1h1NCh/2VXVvt+PLpy0Jx4j34m0W7UB5IjuzerrwiG/wuRmkSoD+bS62MYkNk
gZcfpyBT31UbvdBdp0sP3YbXT2K7Ai1N7/ZitYIXYtq0xeOsmzl9fWWBgs+cGkay
XVJk5vgA9E8QelkjGWzGyCva6FWzn1lD5B9h+i/E77J7N3zuKnHePtU2DcaDOWtB
iNv6h4lcsaQ35j8zTR+iQIrm1OYTgh1XhQvp5reSGGciJHjl2WJVuL1uGVpB5yWe
t+t6oAMTNHK8l4dGLp/VB4TNxoBMFCKOeIOcz7ZOrUNzVE2sfBGeQe7bWZDUFcID
fXH3tbrzQ5+weJQk1dSGLYRmVaGSfKelIaOqGbSO24webz/cBw6tt/Txbh3YnNH1
zdmd5sl6mSQQaqRHUWB1dtRlaheiGj8H0//kp0BUSlmglf6VloK46Lpm99S+/DUK
JwX2HxyCx4sbZEYvqv/XaoeaoXFpLiAbaSMAzjXeVjpj8RaSQLItf9oUph7L4LRS
+z/8WhMkYPO+ctt71q2PaK3uy7r+8/gUeextbhBFhoiM6eD8abF6Bl2Y/db2p+dz
Rn1WPjBb/5EVGigNIgUnXSVikuH1dSCeZhIg922u7xSVi9lxVC2CB3WTJ6Obau3l
p5w8HZBHJz88EJVH0axzDvG64pDZV5oRBKW1Z88IWGc9XhiJTR+uxQPGozg4zLNv
3kC4JU7+U+ijilZTctB4S3r2RXHfkvu3N9n8QcyogsEau6uzrFCNQjLvlp0MOmrv
k4+hnl/OLPBi4lCa7LHgDP/U+XGV6GLA0ZiyHpbDBg239vCwO6q+H62ItXPum+rf
60fKG3UVdZYTj10Ptbq4KBouf8a2mDcE2bMANBFcx+Q/EGSg2o9K/KhzXWLxnz8a
fy6fYLunuZcSf8JX6HMkeAlehWlOma6LDyokABfZtS8ljSd9ih9OYpFXywAO1TtF
cCmrDrXHaAXzg02EZGN/juE/L5gqlFfqZ0Lr5yBtSjeK/rhEypEayeUCYyfYh9ij
En3jLW+1Dd8HC/XIddrtq00dwsFAZtqTUXB5eBMQR9rLfzaA4WBBemntHnUxcBn+
fdho7BI2fdu1JYTWHAJ/5tLcx/MMSsyaAJZHrm64hLyGhGbUh/adE64keeN0L6qu
qK+uhSM1K3+AJkLQb3S68mip7hOaa9PouWNwC+GvsVrhnFDqcrtw35+FSUZaPViu
CpsciQ18JrVMz6Zihcbb/19pNz5Y+n5ONOln/HBkqkfxS9rM5hq7GJ3XGdXGMN8z
zAlTvcms+D1Me6seY8ANgxY4rC1yaRdTy294UE0WdQFcC/2kLdBUhquV374uwYXU
BkjlH/qvOsUpVvK8774QPHRT4cCc1ubsrEIyJclLEMP2YyRjvjbUHU/2ncK2bdp2
8qK6Wn2jonPoDIPJeF6NOn5W4PEqL067DbAPxwnfNv4/Yk0al2JCGmRRuDJ2R0Ra
cdVeyVcZ0cS0AryUaNN5oQ0IXkbbew1nUOwP+X64TDJB4ti4woqy8X16rx0bcrKN
YjM7vus7X3u4T6geR+ihpmistOE/jtmktfsFCDTzMKW+qhMG8DOaDdfvsAv9nccS
4DPQUMt5XFEux9eh4xAfuBAm+aEOEPxCJxZRboacEIrpFcq6VHwdG721kWHyUlzJ
MZjJ4ZRLC0wakWTdIvz3nbaOQ+xyztQeHDkMUlMG/iy2y5ADq2pDTM1eQ2QqMKsN
8UkCgREX6LQ0HtojEElKQAvnwMR9gvA9vfEVtI/sBhgpo7pRzloeCl+oy75f8pMI
b6jkS+6KHDm5iDAao072rZ9IXCTsSdc4QgFJoVbgjzzdfI5hF0niDKqS+K/CTGOy
iKZhW5nrylpdGfo29UAQgluYIcrojJlo+8xInb0giW/vw39O2nHpvQii+P2PE1qA
PMRWYrisS7eQfLvZvH4N5baI1JcRnO/N5mO0d7KyLJE8g7gsvQAYxVrRdsCv8Xxa
U4Mvh08lsfbO1fL6z0Obdbqn9sKMMIQyeUxL1GvEYaxNh2fvZaXa4dhcrluAAzwA
Sq14XkFG88vopmA+B+JUXI0Psc0mbbLGJLf9cUxQBbIfDL0v2+65AKmkpYIiiL/Q
zCpPysVaOPY46lVyPFcTxIddH0iQjYJ8tkfSBSnxzVreh0x8VDRorImIe83ccLa8
WDBVMqQPKMKlk194q0e62milkTZkqMpaBE8SSHSpVR3STSUAJVyqP7idNSPK1Ftn
M6SQ/wne5VQmnyzFYaTkPMhxyE5kmHxRGDBACR1ejkID5rHCl/0tS4VYcCqqsnNP
FA9pvkpwPT3eLrWINiv2fbFVhrzCBTkyJamHmr9b+PAGtWJttuGOrp9crUWtRaD/
hxJ3jF4/dFrfHwXlZOFRqdFjvh6T9TCTSVnGAlZ/U6YdAyv0qdXY2JRI8Tgt9PO4
6CfUhzTXMyKRpvhvdRjapzV8QEgWCHPjZrNMwSoCRgzpVZXwBqJY+yj5GBXnYARX
DlAZQkYMGjRFNidvW+9GJtnA5YUkPcPHrgBm3lEkR8qAQQWZ00qgcK4sKqcwZNs+
EkhJB6cW0KWja3bmzizdCoEquP6Im/T0xffQUv4LY+M0BwAwNRYM8Y6LxEOAMq3N
lcDvjPD02glQ9TTq/hbrmI2pdqcqjOshcBK7q6mhmT5hIAuzXt/YfYmj+oTMUx9U
fKLjHEus1uyQW7rwozEoW+XLnLgwIBszhsNJcRnTAUuD2n3+sPAMdbE+/YWzi8M0
7NDCycfEuKuT2fA1Ozq/4JxsVIexN8FA8Bj0q9HC7qoML0MWSw+g0Wd2iccMoiXn
yJqsyjY8H9zdOO2X439mZ8s+CDjZIbx7ukSAFiDEjMGhzpbmTkKPygNDnextxehL
JJKs6cQ1hQoyB/XnqLRRRSUg1v0sJWQ06VYL/zytxo8XvUmx7/cA2kIn2Gz+6bYM
NxJod7yIFdTsuQRu3m0D4m0tTjzA0ubd93IiQ65BQddxKot4GFmlbnuPy5CghQ4Q
r+lPrEN3k9WGtM1fd8nPT6sSrbQfEeEljZPyNIPI/L6r7+z35UElLM1ldIPbtOA0
Wm5vJcuYvz8QxASZfLEjQy82zaBV7RyzREFsrkGjbp+bcUF8oRX4mF5Sf5YoOEcq
0+Iz+Exxjjt1aw84egZs6JoDyDjsdyWWuVqMduOulJdo47SVKooVuG7oP2IJbg0u
2Pp9oLchWrxTz3UwisVsU172rHmFR9rurJeX8Shzf65OLAbKQPsIwhvTKwZj1B17
XgUvN5nPf0vhhzZT2zC2ur4QnqVyjeGPFWcgSvrMerX31hNKqR2r0Wxm8FenpWpK
HrEQ1jt+A71M8bhnYtsSIlLSvkOLrY6ptpwRQhEKFSU1L3YuuKW5ORFoXXpA4D+6
i9tlUYphmFGw9VRiYHp4TRjpTChU9spTcB+fvDcn50BqpytvV9stx4J9lQf4ptJv
gYsuvUPJX8oq4nsFxsUzYWXjXOk+ion2GRyNkZpd6mUmkwjHw5bRkL2g94Ivv80l
bSLSFvMyaonUGIVKABw6ppLRXO3G8/6viFztux8jyqJgKr9Z8fIhzU6daqhhQCyu
QMJTcmBWMegtqjBw7wqlZqWdP3WUzj4EIWGiR13rukuwVap+oBSW5o/N35YyiZ+a
+Gp3gNSPti34OB95oxOs92gw9cetRpHgK5/O0BPNnGPQKFFZq0J8nzz/5M4kaePJ
4A3mKyUA/3qzYrmDiAGORYHe6C5i8HH4TltD1ORIbtG4OMBf1igxqsEqi+MPYqtM
uZi0+RoAHUoFgi+6+d8ItR8ez0XP0uD2KaEEKk+N0460aJuQobVDh4eAAlzp8Cvg
N9M6Rj6JTlNdMX4hYcgiekakMIp71kYZN+ZSlYmF9L8owW9q0bt1W1yWUGPIALU5
Ncv2Zbg7WYOYflYEDFfr16g072oprze44OXHbr4aBb564/LKa9Z5zKge5qAZTyeB
BQd1B7pKYdFufJOblR1ZuDUxqT+U4V/xUSdRoI/hgVIPAbQjM4W+GOtspyUdgott
mh5DSOykMgvo8gODbNfGl1jhD6FESZnSuJo7xzDvZB5heWNkNpliu4udaWn0rBcL
9jaCHlaGrOV8VpE0UFEpAO0L3/Esdhsk9msCqa6Mw6OG0j8GYc7h8+jnUVvUyk/U
5k5g2iCbnp+TRL5p2sl0gWm/qPvE6hRAkAEIMYpGtJ0RUEsO8LlNb/jcwi3nixWw
p0TZmJcVeaexBXC6yznXvH8f4SfFYu6nZUvcrOTsAv6nS2ad4x4BIUCK/HiTkRTO
OvBI+4xK+KIbyTdX1bGC0wceuM1vb/5CgnXQhHr8vDYWW+BPIxKFEl9tftSQyCuR
7q/14tmeoS+/mv0fKVVIbYy8zM9bWAcM3/EwLZJCvZEPevMwt2v2TnDuHV95Q5Zz
vPYR+v43E7uhPbi8YmCjdKl/AwBVb5PD0pCTdZ6CsFXPjJWXXLB8BvQbwkTV1vhz
NkUS+8fNnkRuvZTDCK1le1PKPug2HZj5geskb2rYuSbg5Ma9euIxGscIrVLOUNcs
FSus9/igGFktU7etMaFZwBConTVAJMasRhIvP5Lyb0k08NEmvvMDMbsfa/iROiMX
pggUfOQI8Gi8CmnuZKn0TwnPQ3RD2R7D2eIgOD+SHOayyoTdquAhi0ol9z/utVnb
gb5cAJlgSCw71Bk6msU2MYVrpDz7C5HMNRoKJaCRjz8uvKl26xc4vEJP2cUldSjI
fDDyx/0yrN5b/TeeS4kkIwaVcB9+YKiEdQ3ju8cxAm5STBiEei9GY4KT1ItsI5as
3Y0Lq31KmBLzPoi742kwSQQZhGsCWuM0s7tkpdhPEbBQiJe6Uw0p5xuMxfIRb4Y/
qoOsOUBfH5FaubyU5We2Oo5i2MnJgI0hinnDpKlIJ91p8xFMVMlavwqn9U4GemUN
Jh0iHofIPoLkLqK0kxwmhHEyrI4T035p4xusCxbzd2wL4XXmi2GHggWg2+6/xyia
WwLsIatZ96lgH/wMzvIxJmxFRjFor48igp39gDiQ4IF+0ADr2Vk/klTXP+KqgkCt
1LVA+/MEoKCWcdb2lj17txjr5dW1W6BJ6rbieoT9ALNae6osj+rJIeM0H05tzEg8
amAi2XJDu1NC++mRulYK4UTGqf31Ebo73bD755oKbGjQtcUke30eMC01LZSnkzaJ
I4VzBHK0yXRSnGRcGsqx2FqUid5d3BWzlCXaobsl5CbSfcF/WSUZf5GoM8TmDq/9
NJUzJ+ObIijmAwy77tIHlCKUIHHjL7z/2YJof9zfxBVbG3FbkjOrsP8jClOxEWqJ
n5b4A87OWTlZTp0NA5mkpZsSpzhA9nDKJDFCSidWl3f1n05jgDU+4hfvPE1dZ6DX
GDLUn/c26CPubaDwn4u/t8Rs316mUYZyDRI1euN9WMFCpVf0gZbmCTwQ6iv0ADN2
mzLq9lFeweUmPFeeTOMwZ2sYIgybasaIoGKrIohuGjAlSlJiQsSoUjalI0VjRgz2
gJr8WO7MUogr1zoya+rzNnGdrrybITRamB5szZ6jfrWgJyZNwAVyqr5pqvaojadJ
yscQGiJJZhElOIH+2/dN9IkLYit6ozryyvwJTbURJ0ne3gN23JGAM91JjZG90Kqb
Y6q2iK+zZQ+mBhCIZk28dNjR1sSLe+ZgWhtmk4OWA8Dg6Bz0RTXgiAYFGlZ7cZvX
zjnty2HszC96+4+74uYZWtcBNroKkMJhYEFhe8Igqd4tZKYjpqI6JCrLLc37TQDr
tHgTvv7MBvJX2K+d1u9oP0CJR/mst+2ntwked/ZNDuZVKdW+e60F97mDGcWxHq+u
SDs3ZPn9V114d1AIca8KRIWARGBgBO55AORb71HugIB9Qia9cmlhnpOzPft6vECv
wBpsgqIGVQVK3lx1yklg7NTbFlH0B2pnHTSXaEtoEHsQ10WM83fFYMkNf1rObXA7
YlRbGbIYA7mVVAsMqOmGXxyFPKrIxIclDgwPzHvnFFwMLJsEFenEqhSQIFQzah9I
CPuRbcZkc3nR88D4ZKecW67ed36OKWVD0ggQYYuUzxRrwXXbjHRnb1gqC1uVUM9j
u84c4gi4DbgYFkPl1w5Tip25oSlPZyH0LE76bP8rqjafGrZDRayUuUEJ/FMxt8Yb
iEVqpgi3t3tXRXhu7taUp2IyEePf9ED84xrq53GDLs9ITw5JUPLrX8M7EWTKoYgk
JT/PHEtdxOVtc8thYVxvxTjw5wGuelD/4PtZu1yT/HVIDODSvfOtdXMc5dBa0t9V
18T8lpFPlec3+VScZbWj6awVoLkbbj9MlrxMWLzQ6ufmnOkhuhxPbgMvqUYkTszX
wPP/w152aMRdyzxeRLQHqDW+72hOM6UqwczEfaOdScDeWVfx0Es75URx/zJLmsBD
htQpMQs2p0+FJ3Ch1sYRbnf6Q0X5nmUGsdQEn7lgKR0XyMZwhjDGnBGZMerXgpdf
zeuVcPmlpDY9fUtGphj+WG+ZpFQdydrii5EaRxa/YiE+6JI8PWUNb2nUaAhb5SCl
Q6U3tr8eV+L4RutLCqloBXut9x8FDBnH/AAiUl4QmcFJ352m9tppbUwkyCzdQhnk
r9Jza7TP5gndOOJqiURxSmQE2fPI0hvrFJ81r7+g/1Y/mSENnVLZ0mbSXDA6OJD4
gz4jjFnt0XgI528I/ORusKowVLSQzo78Rz0OSzwuIETYbYv1W/FrZCBgzppg94Au
fazE47yc8+1TPVecMs0MW97WhmR0VK/K+kKL48vYoJK8TWKd5j5TgIzzM8i+18tx
21Whyp8JKNKlQJSCEgVIY1Qo47KbTDY3eWg6qXrokzRP/bNd2dQt5+JdWr+9U0EK
ikwGeQbIXlV61m3t5Col86OpTY340n2XHDrDx0TmE+lICQha190PZpmD0Ln0Y1Ey
kDTXLfPc7wPY1/ON0sh+Vilzw8XgEhJDmq3OIzc3Syt4xm01fwHyAKwpNVc+ue38
c0Rekw/mc0prioD8hMmqWvpJH1ttS6XgwUIQ9niFcpHBs9eUgdXicB/CDWGZCr8h
8FLlrHvFSrKS8rqqXc/UKAnIMbQoDbZwqTG3IHs51bE7XR/bc5lTi0hCPk13LJBa
oC6jMVUtgGWGQmJsAlKnqmuDsRFXEHErBOBhslc240TeLR2xqnkfyoFq0njUH5tV
Hv+RfTKzx+2nnNaJ/UFZMjH/PHMtvvaWb4CroQKL9LmCXiUXTViZ9CPJMRklpSa6
HFCQTQS8gv+PvbmvEerDnZ69+0yMZ6UzlyoE2vfy9GYRQ3qJi+9Lq/yIH9FeP0PQ
PVZZDJsXddMlYvccVuzAibG2287he2R8DKXACnRJKDHh+y91KUgExFwnyG+u5Ald
BCRTy7mnYq4BGnm+lHqn3Jd45wuVzQ7paUo7x3I4kQVv/VU57/VF4eT9NGC/vzQX
PXvs0ufFJDi9oXHvA4JZEQWWnaMdZ6WFI2y8ULhc5yqoB6ihbq1l7BQm5X1GE/4U
xPlLnNbXrwGh24UzB30OATyKmTJBZB9BZQiZelR08dHizICJjNLzKp64Vrhwsfr3
KHByrXH6vf6awljOmy6YU5FD/Iaes4X564N9gIb1HbJC78MBkAbQETj2uUsNge6s
rc3cbv/TwmJgjmhIlfv8WOVd5X2m7SKT7U0DC9ZbwE9QiabKVKN1/dE38vIYRbwP
bIOQEnHxORjXO6nMO0Q+TvL0ygx574r8CRrI2dWzdsXrPyg5Oxx2LgCg3uj0I8+/
fYThcEAD1sVTFXL46EJjr/sgO/C17/AU7IW08nXMbJi27hWVpPHNZHHxRj3AgcH8
WbyNnQvoE3OjHS5orODfEijZqTxzxy0Xtii7I7v2EKrTV9FH2o67htLRvECAU7WB
2v/qhTr52h/xiGEWQ60Z5NrAarKaEYOloJuB+wkizh8LUMdBxuPSvKidsUpYpjed
uXw0BZM58N0JnldcUgqFAtWqbWmCQlIDVdAN++F8UllLbG15SnyBMeqQcQXp2grQ
lSAvwHZ+ljFf05vCiBtvhw6cdaVpw8YjE2pADZ1amG4VIW7W8tFLceYKqaGHZ80g
alUr/RWGALrD3NpWefr4Boqbl4+NO7R2NRe60Lw6QbnX/gg4t3yTVbHAhhNU7qL7
yluIXtRVRNTZSr72sj0dTAaWA3LSP3S0u0ZHlDOONqXUMTLAK9rPsrGcWq7DecFd
yWfXzkHBQPj19Z6FY3dvlk5/ohvw1rDRi7v0XVsq9RtTRpwA5z/sL/whudkViH/o
x5L2qXZwgxSHsEJF4uNWMe4Z1SWyIqLwMkoOMMKptbjDwKxmEEynQYt+Tp0BcMpp
xYBl4/6ew1vqklGEhWKN7WLxggvUGX5FCvPcPbUfteF2q614tuzySdRWO3q59Jl0
7WaWf+oIJb1kNDNjWgVW1T4vwSNCCUBnzoTNBQGQavh64Bs+5/ErjbTXKtW1DTjz
sh0fwpykiKfqGoO+qcwqeC89XN89s2zyUrVMBoQOWKxQflbQ6qX43Z1m007FVjYJ
LScrd6XqfrhBhxOK+eyPmEZ04jWww/BSP+c/CbRFZq+TsqqL4fwmGbA2Ts/UOXez
47Tgrd60xGT0aZhvvTovC996EV/lTi+Cm+PaO0JBNuypF8guXsWtQwEUPmqSwslx
4W34oZnP6MQvsmR8qfwe0YZA4aqQIWz/YSIQRV6O9Q4ri/HFR9HNCP/ORJffSeji
ky1Npy72tejiVcxQCB/AAiePyu5d2ZDKIpDPzQ9l+sQJKrXX4JLioH4COml15SJ4
1qwwrdPdNi3ILsZv/pgmbrtTayBWGc95hd+ak13yZ45a/GP9stOmZfcFs76HfznK
PTHBmHpFueusutOop0aXanKp9xGl6UDYsz9fudy1L0roKUR4VNujBDGf3/cGzI+G
To+YgFnW67HmsTu7wytXJs8xe70qZFe7u8WAcTcrNDCPOUWzJ531lnN4BJBWeM80
ewf0VmnGnfipjfvT/TqizZn7bW8fF2UYZWkTnbJNBxUB4B4JDffby5wSGCoD+flY
7h3kN+maWoC/Ct269RpMG/8FaDl8lialV4Z4VaWEvrx3kBq9wKYlgP02hBdRuyot
t8uUoWTcuH1L37IzXWkfBvvy4NcoM9HbL2JWu3ZwQlVy802xRvBiVoZFQla2nwXa
aGqcF9OLYN7YrUyjmzjGrd+SX5QEcFJ+7Vwpg2Qdk67tpsvzBTVyTCJVkS5j36ct
IWcgThfaNZOVim8tnC+pCNrvcqhyZhe5y3fke1F9kZjlao+4PmUuBFNjJBpcJUot
ofw9PWlXUZtY2bIBz7inD91mSq4+J4L17MDvvNpcxp2OFNVlIm/u4jNZd4Bj2rI5
photYXB9yNMm3Aay6vtnM0xl54JGImJ45oeMw0F8c/RdDXcjF+ljLXVvkk3NwqV/
vDw+HhJ7v4449zPHsRh+4H882DZzz9/8msp+FGITquj9nhp+TalGbkkx0Z9353iT
1RGrUdOTHeSlv5B+CsUwCv3UbAc1oFunVvja4u1z8/NhWQgCh2ALTyP4foR1Qkyu
+VHH0aHPcb+zgdpJK1E9hSd98araiErYj14r/xOGNcQthRJNbUtCYAl32cpW5bQI
HiX7dOw6L/vITx1gJudJryjT0EN2vRBNhdNhpB01G5OFum2aKe2WqVVPuZs+OJ7A
lDV7m9oG/4OgpuAtRSh1R3V1ZJKOFn6GcKbCLo5g8gfFaIlYEjVJPiftKgnjzoIT
WktFj2Gr2XP0XD/gPQCnn7VZdu0SBbumPf1fCqJwPpfJU9E+jBp9NVwCZazzi27H
INDBEU1VCgFPYIiZ2hGeBE+ZERloJ3IL+jtQW5zYUiVjhVpQvINyCNCuupaSTcfR
ZaNYvjT3nHmcO0M2pU/Ismks86/t+bPzuwrvPVoszeNaaSPKn4tzsYU1wdmgB+FU
vmQdAadI2j4jX8SaPtP2Ult5rA0g+Dzgzd2Pbb/LX5jF6eU96TaBaPLCXAlg4Yr4
fXS2WNeVEct0l7UQ/kp6qDX03hLIahFE2h5b63cZatcQCD4bHcNW2s0wKJWRN85d
pCIt+XF9gCT1SSHtre0EVt3Mdp//Sv4ViF+qUxT0957SlQ2WKfoklmoznJMuAulm
eAs1th5rOFsxRM9JvlmCsO86rzxhoOPHzQgtUKC5i6CEYBkfBLvWGZmq1y9jEzeR
o6R64LseTNekIfXlD1+GJ7MVbgntqKFVpwJjGidJAwnMvG06T/v28/M453Va8gA/
tlzuij+MV1U9ZA4QF2ZePH2puK76x3PTRs8AvZK+ThfjwXsk/XjD05AuVhw+EmAH
4pl1uSMS+s0+NnCm9lR0XpwNP4J/lm3zF6h5vOe0DFmneajsoTssMEfqoJ4InsGT
95W/bBy6f8GKGHEXqhK5PHtwqrHEOuuH1HMdgDvUw6N+1HQk3BWd7M0Fuw857deD
xKJE+RJvel/ctdSrMlZxdvBhYoa7pmxB5VcOpE5rUrkMhAdt1gdXjfKQ0vnlOgkN
ttCcNPE4vpKX/jY+JAdIIX1R41wpBFG538uOnlmbtBFDlLHsz/fznUbDBVAsmp+O
rJY5J0p6pLnLIsw0xBQlmiKeKjcx989VymfzRnWv0R1JE0ScGArHMXiwMNXEPZ7J
GebFPCMSJGOFDb22DE5CWvWd+4+ZtUXoW0VWblocSp9DYolMuG37SGrf99u/Uc63
FL+z/QvSqIm1hDjss75dv4CltlQqS0MoGQISVdUY4tBMKGM2FaiPaMx5jF6UIK32
toQiYlpGVgLv+ujR50LCS/jgmg0NLIfBP65aoOhaP2RYdNLrgsOlGUFXbgW6qh1L
gT0sR5GNqcc+x+UefPpXuLRDauw5pW0antzaoSJMLSM5nA8XLHfvkSvC42+uz1cp
x1Nt7na+ksAPf69jg95EnsgSVjS/JtDKcxM3y3vQrCTITcjFh3EaPEh6qnjqqAaK
fNflBiZhLPNicoWuRuo65j2Yu+6Ru2LBS4auNevF6EuA5ShNQzQTPJANpO92IKCf
YDZXWHa6qoYUMP6ff8x5KVzfZZ19uYRbmp/GXj4SzrVSTshibefYirMtNkVUtW2O
GU5ZA0AKDiM90FzFzFvWyC8KEx9Rqt/DWgFe8+qUjBZscFIiA4Rta4cqOxdUdu+j
9AaCOrtrTVFnif1cSiimfySr2GRQ+sFhKlSqwDeyBLBFuh7td0YJQKNWna5hGMuo
do09LZqAl9N585ykQjsMdC79ZPxgnUlYCB+o06DgGRfu1tQr7HcMMcrP6reOaoeM
3N39gqUiNYnusRjomt2fCaEuZcDYXSGDfgE5+76tpuF1bU7Z8q0jjLrsDIvd7ylW
o2Fc/cIC+mfEO6P5DAjE0xT5/4CP9VIktIHXienUHb9FVqfE9OdrgudvWFFwSoyt
68iRHETG6UJHm4iDjNfnh0EbgJAwuzdCqkHwcpgzva9W0oObViRI4oakLs4YaEhE
8Fk0K+1JPcVe5BgslDVqgsSQFElxb/GmhzBSQ41mw769zK+yYt09a+4kArY32orD
Zhyvpqnko4qnnBvazFvp9yfuWh1glC2ZAuMvKNN+0/Ow1gw1gFgaslE91dAS+RHC
96ZNlM+IMIOs1nYGS/3+y7WjDW0MiiMOluYTgsIbBmwgm64ZXmebt0SNpmLHzU2a
ISDL0E9ojvxSyoxtKjxerhQiy8zrUUr1//WwJJv/vLT/YsWSHK9mrMPfLjVLOA7i
kOI0yeArYx2Boog4aFABTsLECZYaZQ2vLvR20RUULYq3VJw2zVENhkGBH3BvOZkD
SU9M256pOWVLOVcl/N2I1flOw2SMMfz/tRq+vhURgteG1y1tVTOwkwS+4/k0k1t3
mQ7R262p/DZ5s0xVYH1yRKVIyLHYzu6KpY+riCeX7bW/9pXJ4f4yExE0oBOCjByV
DxFHCdbO6I3nu5Z/M/QhsRHzeChGtS83sI81h9PvbPGQPm7zNMQJASqoC9iP+yu2
mERMdh+A3LPk2pN+AmjvHIPklxzO1eaDt9tW0g3nFL4qsIyjGE458FAMoma4o6cs
KHKmc5KHu4Vp97Fo8GERpXsDaf6D8hoymmG8MYKCwEQh4BogIud0hvbYtcDe86cO
MUoqW14XE16nRuSdeaVAzFYF9tLKh3cX33yAAQ9h55UoL6TlQ0+Q0Jpo7UaPYqOL
2Im6HszR/9O7excT65IAHnXV5kuBccBrKBPIFN5UEN81pPpXMY7Zw5r//NKu8g/t
rRBAJL9U9drXPFp+S7XeufVP5Mrap5qsK3Cc+rFBlMl0Fo5+AW4F2PHZq0j3wBv/
HGfAUyrGbFZvAte9A49h+OV4mqPxrMQlBvT71fQJXXgZJPAcPKCHdV+GtIjVwzz8
7lUI25FH78E6ORCK0b1UUcYp6Jmqc93Msv+mTOTHtpEgvzoPwVajWba0b84b2Me+
y9+AxxnxGYPb7diwjuUfnzQElR1HYIrqYrVhwr+Ne8l3SgqqsRnba9fXcvYL4hqN
4zBKy/LDKkqZ28r+9lncKfCM9W+9GtkQpcRaInxHkc+38/vu3TW/UTWSiPsKvfZ9
hG/b+uuPt9S/4CFJFjN5Iw8OHMLf+gINYBrbV1QYpy/6fQJYlNEGqexR3E3d72Yx
kTYQvkyK2LuQs3WdrY8GXtfixId+3S98uM5I3hsGZW7CKacj5CF4Up0KX2pIFNjJ
UlnmRANbD+run8vN196ZwnN5OkkhFhXrZZfolUsngktK6a1BQmGaRVn/NOOnYHXq
oDpZqV0w9GaxV3GA5JnFQLKWNoyTRrdtdtW9ajED2wHIAPr6MiL1CxRaq9NDNqt5
Juq45Fd5zijwy+TtFLcy40mwx4U1nbS+XbAcaN+SIzKHFFV/48QcuwhFpKbnAdxv
WsDqBRCSuNkaGXfa/go2u5XQ7vzW10VFcS8HFf/5evoWa9w537zWrIzBNiktbOQu
Sydlv7slQ2z171O5UTmuepshuiOo2lhTI8Kx9/LJpwJV+BKu7pedhJfRjQxJiPEw
YHX/spFnjJ/cKPSnlmLoN8DZmd4wVK5n7vqcKm8U9+L7GzF+oBJvgyG591iOd1X5
sOwoI3B/jGrzc6AnE/OtSdbifB1SkpSLioZKuC0jgfGuBN747moy2Cep5nLl/zYI
vvc2Y/8n+LUJhFA2AWgSsM4ieBf6HzHWPdn90cRdxH0QTT2gznhQyoy/FVeIdCRV
vEv/fhr8fC0+EKxdbRMg7Ln8tj6Nar2ruQqE2g0AxlTR1U0zx1VeAfbay36e3Emn
bIPzZe9w75qXfbFxM5HWHbXcW2zZHTTv20YxS932ZsqN9YPoCy2ZUJxsKfhsXZRy
ZOzvRfYA0Ckh2e29gMk4J8FHvY9OpzA/bO94lDZmy+MkC78tiDdUjntUD/V+YMPI
PdVvRJTgf8JJyWHTMj73NrosSVZ2VPSmdvp4m8mRjabQe7S9XQQmi4axgcHMeYGj
NkkbIa69fK69/eUmYUMZZBAWRIt3lg/TMPOyK82l0GyBE5v8QcnXQQnAO5CF+aLj
wQMrpi+NRmhVyavT0lL9RsMY1A29UGf1SGRYaDMssfMIo4yuA4P77y47QiY43Fcq
GLiyjsc8dMWvwrCa06D2G1DionsK3nfTVwP+zSDMa4xT2BbwaFoSiPw345IAyd6h
OIgw/CPIFIwcBrEYkc6jmNX0/Aux1rNwaK3lgL47FArHkTI9NqKGSY+TEX4IJT5s
sEGbzVhnhqtJVmWbc9L1AlKOp9BObJpHlvKUWm8z0FKRNTon5cK7ImfdPOql54pu
zFpbYMN5e8w2fZYyzziSImYbwUFC05qRp3DR48yYEsaFnyltb4PvZyvCzlRe7RkZ
d5s0SRw7tPBEe1hxtyLeMIY1Mz5knNP5eNjOf1iw56iBjsiA45rsfFYJbwKA6Om4
So47VsmUAiF33yf1apO1MNcKE+4iQu0yeZLLh9/1eDtey3o9w/f6Uk5LokN599R9
j79o5D7DUz3EigdXZ2qrfghWMV41AtpwlHoQYMznsQcfQwDIcZ2n4C2/woURWmoB
1K0hwMXRAuTUNIgAM0Qcp+O/7ngmI875xr75azZin6Q2Ti37ASNBfV3cOxhWLNaK
l2f0BMAvkEXw+X82SVM85FpUkKLEqWIz/XsR9Tl9GQRsfE54ALRGGEQ5Mir7dOHD
D9pJbPNJs9I6WdC9ypP46gScc2+9zA2YDusC5gl+fWih++Fsu4eiltFRYAfWaoFc
cfc+ctdxkBEkLKWrX88gkNTORYMtSdzPY3Lb2Hj5lVs91phMNGUvYNqJHlLjLUuk
szNdhyG/w8xgSkc6+RXf+8bZx6FHLwi+vXlHiPoehgy8wiWs6oCbo5/vXbyvimfA
wcoMUMr67rHHMRbg387/b2iX9hoTLP7/xDkenixsYMfS/zP13BOi2Te9vpCJgjGs
II5vdu+a8I0alKfz6ztY/0/VhrUI08h9YZUzUIfcqsxPdn1vjoZ5suyJyAO0DhCJ
AiqBhR7b8kWiep90V2HgFXUxi9LOIhXaNFDF6fLiatBaVKunYrHK0h9BX/1EotO+
zE1PNrsN1ZyLUORHyObNSOiE+x6a7RsH6ebNKd9CUMirLRwY5qzROKLn/rABBXFs
0GqiF6ZRswoQu5xkKUVygQ0KovG3hRRR8d/VKcBwVUlneEPK55mlE1xXnyhkYbwr
8AG36mTQIlOYey7yVNpS7sdz4LpHWCT9fI6toSSkkeheZM/OB69s/su0a8pH9Ckj
rplatJrQi4/DUn9ojIBNEvgIY0s7c8Cc9ih2eItDLLDp4E/VDm2cB4+6boYAXJAs
yYeWgjKmhrl4Z5vekWIvgx9rZxSwA786WhNdmukSW4lABEfb0OZ9F3YoYEDNDKHL
OB8sqsygi+A0IPydVoYSVTk45GrdmATokxRiNc3+vG1driGWzEidQLbFSSrL9HzG
JZopacmjlDcLJixdI9TmZ5o3qXNQitEatEU0DKnBS1xnIcRETsQZV0T5my4/1cd5
7a8lFAHHqu9jOOgE6ORCF803Fd+YNbO/NY9tWF1ZPqKBZr4cmeBr3osbWA9IJTOU
9S5kTLIk8DBoBLZc5DmnfVHba9TlDc9I+wqpFGZ4uYhF6hGfkebjLPAsk/ZLeOU2
+hZNYQzZsBXeiCzCrrpOm4l2cgjo7Z4QByKEmGkJKUYPHDh8qHq8UlEWx2naiWdJ
OBP9qVCy/KWrNPS/llDSVNapAAsnWgLkqOGBI5gtmXR4gvWjrecLp2xixOXZfgIX
sY65Tmib2EY61bzXGJwsmVKKXN4j2ABpORITmibziFEnOImH1qjt/R8Aiuex40hO
wokKzhFVO9ul1X8JK/PT35Rm3NfYFPruJRcXBCuAo1lHOCCK0Jo9bPiN3yoJeEpD
+GX2ZFZcThVojN2VTf1vcRQlIgbsnoRJDoUoaA2aTc6hMw7vgpjGxZvheBTrhJ7Q
BSMGJAC235ik5a7sgLJTV5UODTSPCJRb+40I9CxbL9LUjWRZNP6+YWv7rB61RUGc
y7du3ZWBqQepYGcFkQZcrHipDAI8yGHBjuQGqb1mBEU01vNqpmYDrr+b/O4C6Srh
Jp8s56YNWmbJ1te2eUA58P8z3p5bpNNelGZ5NW87L05jzTY2TYIOM6wIX9mZOBO7
EaFksMidboMzoi4afhBr0Yzt1kv2grHG244LSaO2ZGwzZmAqB7sDCkq4M6jKeg+M
bn0dRZ4ZkyNBoBhj4kWDH9RHh8DI9pjBsoTML6iqYB95ADN0nSDDYoZzdNXI0EV3
acQ4KVdcvi3y2ewFWrjC3Nd9WPVtKPXjiDMniG4BQySmeflJYgfWbTRMgNCVTHCs
IBiFbwINXSI89tOW6bGZ/q3GI9qMlc3EEwwclbmRQXiteOvMgz4MH0qptBQdt2Wx
6w0tEbbAKAH9TOT/rpzsHd4G45SxYllfZC3rCd7YoVg5RdqknReqflpXx49hJtEO
g1X2voRy8BU5t8m5u0tbbkqlZVdHSfdLe2dc2++eJsVqtjIDYzL9YvaJevo97ddQ
hoLtZLmBcD1ELRKbc4gbw0AUtdrt0eI6N93RvaQhDnYifNkrPbg8/caAZveLHAhi
qhwZndkJWw6rscL/LfzMh4KMQn7XfZ2UbeT70UB3xXi9V9mfgsQ5CAf55CYhPJBW
1fJ/dl0rVxin4frGYomp0XanJfwRHrpY7CJelFWaoa1QLBHElF9KvV3lmh307vDI
Gjc3xssPdlhuh+KyTZ9hrajlwS29PIi43KaTqgWeA/Fqh+W/2NQ3cnImeS5Qd2q0
yUc0vfvfODnGGKXQQBaXMR/xIdk8fqMu1cJ5ESFcX7nzGWf6H494F9y3RjWtp8Q9
PqUcDS5kflv51thiU2iB71t7PSWYJsepiQCBob4sJ/we/KWG0rEJn51HZMjIyPNG
I7KOLVoRJk/n11U96y2nqQz1cuXtFC5dbywzKiBDr/Y4JHmyAzkphf9r0GaBlC8Z
krUfgE/PNfyrSSdwKTuHZPp5gjKHuscvdqG22ZJeIJE4suMQMgAev7r7HHKwaBIA
f/sbS7hA2JgKzRZ6ESdhtDHN3NOYA/pWQ4+M88XfV5elM7FEA+CvHCKPkz4/wtQ7
sCCMmoH4xHei0iPMRpOlnxIBOG06Xd6QBVfJuIrkoMNr6iuRkAZ/8FqDjtZwpjZm
wxV94vq93BUvnyQYalJfnmaZjgrRbY6nSsGWCycV2pBjueDAXHSF5K+TAsM5Khkr
Q00KZrHeWj0/H1fuCRzxeI2nKQ6nUAA3S9viqonkdw/SdX6oHnSRqwI/F40owMXG
X6wqFnYpuwLYrjGgbYAiBkHwJFlIMqLBJ60CyEanPHoz7jCLHl92OvStH9WMJepU
J8mE5BNaBGncEAZn1aDx2gK9bE7Wevzev9bc8vekG8UdcdjATiDzjMlUMQPBMSon
SFySAzdxXatk/Us1QmDAkJazR1MqG7uY6Gz7/nDvPOOD/eY4CiknwLRhdBbigEfr
nsUJQaAKZbtYMdGLi3nSnStkvrS4MHjVXU6wFMx3j0jRBRWTzo8HKWJgq+CcwZf+
3QAMwf8YxgGecylnNGGCQzmRNVl+edfmFS0V2b4Mx25uubmIZoEz7Sv3gjrfOFWy
3f5T/qg0TE/jHhLKMCcKYFjHCDD6sIc0jmI1LhNnrdV/diJcpjfvv8XUakL8oSlX
oAJoP4HactFs0srVPF9PrVyXue88ynYsOGWL9J9taclTz8VXkx8/wjTxL7bsacJX
5sHSAHvUXccf66YyziQUorSq/Ug99vKJVmVc+rrvYm+eU1vJh2+5lnN7v/IUoExz
YeJAcUi6mtRbsuSlPxIe4i5D9HnFVsw4Y/Z2xZnUVMX1879zv7qjplrZ/60tZQGz
jZBezUFX9vLJtWBoYqiXgAVy2g/0V5R6dq9H7aHQaYtvHSiYo/h9CyaES2hE0qbQ
HIKIGzrx07SB57vHJK9SRwcGK1ibAusCi4wRuB07KCq4DZ6tAYiK40ocCzE0feI4
kFdZftUJdWt7JJXAhwk2KiryKFeQ67HqpZROMmzCJSwO4DQSQEEyQrIYS4lxAZLM
1jB5fM+FwU7f8jj5JBsjUJDv/1MtGdDHIPcxbJ2CEv2Mm+h5C2TNxDuIdeViXKRv
psRpMsRHjrehueJEMaYT99yt9sQUG6oH0+Z2Uasd2Zb90W12AatIU09tgt3ILvzg
9hyPNuly6HoUdzVWl2dO76cgCheQJb5lznZAf10fzc+4reL+631r/+7L/EnCpBsV
OHLeDk9zaD4BLzl/wSVWML2G0MvkT0JbkSeTrXEEhYSX6z5937VyNmLj+dTU34Ol
VdYVpBQJOo63bVGVS0BQ2batH227LRilSHJO4ERiChiHA/j59k/h5+vPAb2i6ol3
HfI+A1n7Bt41rx2UQvfddOeBWWYycUV/zsIdT0Qj9QC37TcqOG/XzIvoBRnqz8bx
/0TFbbgoE2lwaUX+Z5Vfk6WNSzZnt/gwS+qUOSiyYdhCsh68oiEV/hH8QRv3TBfD
awxD2kYemGmPVj64E+Frud+cXdQ9EgvX9wAcvtz+ehSuQW97lrfdJUOFSgFMxHUs
QnGGUaC/ivPE5ZaD7FCAckHoTo9E0X+yBWPAiEx3ZNl5RrA2HOsIxKCyl8ajJWrz
EcqB3nHRfL9loukgC9zZuegR8oZK/hfT+QD4H9U1/KuOH9lpdNaD0hFWS7Xc8t3v
v8kOPJL5SQGLsh+2q71vnkSlpRe8KXf5bG0rc2gxmy516V6vR9LhIbtq2RZi5bZA
DrTrul5B7wpqcyBwFHGfLvlO3EdDM9U5/mEq0FjpCSCySsu2y9Lv9jhSBCcU08jO
QT6cCnKZRU9htdbDW49i0QGjmdYoqA4Hv5vCpnhwFkQqKwH5XxvpSpa3Pi0NSTVm
KPjBriApJtMz4hljXQubIYlZ/rgGzwyZnXmIZ6AmVAWDr8bT8pywJI0G7hArQhH8
19k+WiCye44iNYfAphAJBWIWhJUHSoigwsJql/nHnklqUYnziLchPz1H0k/JIufI
Tot0dvx60uMqlZSxXotVn5uQfVDOp7GEQyUp3Voit7cazUoBNZrltBB6ShYD7XO2
Jb3M7iVfHJ/dPNj8KSgZ3dIK6PNIMUs/9FnzRp6aVMgXxwnoIxVOrh0PbqrirZba
TKipdySPyaTE2znvuUy9/fSVzXNzmRqK/hHRasPoUAQcIdE03JxIrCMZJrgZRRfP
ZNPlCVLLcCEMi+03fVcwVOdaAwtvEqgObsR8ARhaeEuUmFMOOW7Rd/LL4RaPbpJy
LR5ckbOmAj0qJutmZicSzoFYFsopyc+C5LCJ22nUT7+kA5+QRElTMI7XxhSazYBy
mcM/E048WZeYVojifLgFsg1q3hPP4OYckUiFYv93qVti3LW+Poi3KpX7LWZ7QOUv
djOcaZJyoFZbTX+u17TJ0FlBdELYZkJn5raVHl6bTCEgkl1xBGUqj+QinmgKwETb
09LqbiLD4zKeIG4rF6OuRmzxhZXcL8AFMRhh4D+cJWz2QbFFpRYNFbJAxCGpWBhP
jX3jw4QIVApZ3cmrLznm7BnM/9TRA9NrO2rxw21VnEqmPjH4Fw19O3erEStVckKt
E7DQbXu9ewzsCwnRMSEngJdvle3fgeoP4M8M6UBeFG9M9noX87pTPINRYgMbJ2GV
qadSPGC0t0tzkbfJrl0G9nKCe4ZKxjnhDAyBWr/j6q5poDKUZA14X7knNDZVbz86
xYE3SQWNgBe2ZqpDxDUMv85kG5GzeIoRgVhEx1hHmchXsDNgO99A9rz/rfdVopeR
rgIlYGJI6M7GN5Ed6b1IOqsY9tjFSWpvJyw7olamqofRup8V4Aqna3QYCxAuC5Lw
rWs6BVCC6ExoA1p9eEfMh7OmKNej8zljOTWd2KnXPHjxKziIY5KyV44yvya8mD3e
+Y6zjRyAHxyIUZUpL9Pfvse3glqpB4IYTM/M8BG9pR0BlsuXvvpHNi0I6lZJudST
xML5YoITNVvlA3DHQ4oPCUcjJ8efH18hY4WbDZdh5gSKy54AmoT6dmKFbdcU7/Y+
9MzXqyd2OiawuRJZD8IJCqhHgIgeEkXDKqecD1pPbduBfAB4tLthI5GNWLHW0RMF
uHfPnq2ojf1riWFO8oHni0LCU/85539LPlxQLOqX8ePsyPnK15ktigvMKTu0z6uo
dLZWjxgC1tgG0RQWSk7RY6Flti+SjH4V9fI/l/SD/uWYs/zCyKkVFmbCqI2fj5lJ
631wUNRF3lqzoS7w6no3Ix9JIZ8vhOu4qI9AJiC39cnsZUhC60VGG2j1Eitlvdx0
DUyEAwr57gjYpxYdf5KNMbM1wEhegjVh0DzWaX7r/kwRfuNq//hvfRpJCwjYI42A
8qZHyfW1xMSz43fh3xj+Wu6FbV3zJr7QcsoQAxXdzj3oMNFW3xonEDBhfdjkzdGH
r2aMJQ9xfTtcOWuS/EyqgC8nY2tEghue45rKYiC6V5OYySzsS7AicyHE9fpiv3HG
AYXFmggNbAmtD7ZJWxqqTQXh6Adxp2FHKEd4WUbp6tPkHev1eYtJNukHGNsqaXBy
fA5eK5U6GWgSq8YB4mNqSuaRgdFEKmrfCpw0umDfiu+IdfYKjVI+h6uM2H3wvfGY
z610oo8VOtCiBKMKcebv0/B274fugfUMIGBkfXTkJukXzLM0aks1GZyzPzv1upbL
WfC+gfQKlFQgA3Lzk83Eq7LsWgDmirAKRoLZQ91EuKmcGPzZxcFP7TaVjK8n59DA
iYdx2Dp56WKwsz60C4inxBMbCSAYEngWAM9byZBDssslcFQPEhzIb/+g8ajZM6n9
oWE9X6hVXza6u8QI8GrWTkXyJCldygGeHusXmERSQPs7pmfu97BZo0pj6LiTDmbo
l5a3xvkafngeMbA1cFAM8lDyLaB6v4Y32oG+SnRCUnRNJKYAvFrH+Pdx+1VALq6o
XfNM71XuQPPYc4Xj3nxLxCBoEhCZ/0RZheqIoC7QMjZ4WP9WZJq1fjJclqUg7JT7
+dfldFrAZffJSuAe9a48H3HB4t5SWpbAVK14Rwk11n/Ffb+zgX9rFBr+wHL1r4EX
Dgy4T15aBtvgtu5IxLv+K2zEb75cQpLV015xYeQC1zqAUiDtYWqqSD1MKJAMOcTd
zlInCAd6uBABXCCDo2eDlM6JQR110Z9ENNYYUfwsY9dkak4pWG7jaVKpswQFEqhJ
eoA6Yqfb1+CLBQttdSHV649ggqUCoyGqIjwYY0q60fVqkrZoT/9/Z8Mfb2nUu5eL
atspLb8S4gSHJmPcR82TfT5d7cAGTcKwydboVVe+6+ek9mcoAyGUSqt8i1RZTKcK
RS0ICuW/EaNtNUdoJfaUrIZkuffxlWsfieDbYynYskYQgBOPPlSzuq5LgaiQlA17
FzObLLH68Q2YVdapivTJw/uqCbkADQjDD1vmQea+EjGnXcI4M8VoiKAhPlaK+gUl
yyoCuu+auM06riFProMeGqJNc0hcqRQjQFk6bWRPuWR9Y96DSMv+wFF7uCeKRGuY
PnX1ZOPKEWG9uglQ6TbbV0o5IJfhnLiP5fu3aJ60sgoQB3OmdPvaKCq/LDTcYsNV
yz/hSHtqFcOm6NYAdAbJDpzOcAYpYEHMeF06mz2oLUdioGfnUwZm7Uvr4Qn9cRiO
ZOfaUathNz0hLVLxs7s4ZyrI1u8r7sJM4ARMdyLo5/guzkEOuLGFk1y0dKlDWKLc
xfxRrJojVd5NMLljnTbz+GVKExl2PKGOv4E5o7mj4bzqimmJNPmtZ/DOnszg8mY3
xQG/Vp79xb8OGhffQ5jQz1iES1NpC3hhqEKu4w+QHgvor+Pmg/awMzqRxt3dvXGh
WX/z7Gx6OoYddYE3HKGeY9hId4FLZ3PFY0cSYVoTgMf8BU5oWslEpHo4NXI98So9
xsZsTQ42XUc8o+YYkz8cHEjQUfpne6IWlD4FZdPhrSBvqIgPyXonkglJ02+ic9Ga
yLXB59NVYjbmh/EOZ7MmWdaRDXVDAFIohS5AwMVf3F33zionISEzn/or74v1HwMU
N28rj0ssqefwpZtOfnsoxKNP0namSGphbM+2gq1bhlqnMuJmrCRQCOR/NGBVXkEN
XWfQmDY6HU/oNWYXp4+mAsdhntx3H5NRyo6oxON+Rp1cYqru7AHXEkqL+IAQyQy5
uFX7+hJ3palN2FaEMNQXeiwK4ZD46lEIMtrHjXwxH7Ra6OlpqcPkEI32UiTW63zc
KHPC5wJZT7FNY3VnfTx6UUrFxfz0ujvBo+l4MXc+7rwi9lQXy/biuVcscu+CU+BD
Umv0oYayZrUzmhOZ/I2i+JeA7LAEuNi1cf3CeE6Cx5jnrW49JTuyVxPoFnU0iKMv
CTNVchUIh/+zrx6iATpO++eIo+dG7Lvummkg/TlLjmUHUDPbbmNLE/xHwcPoqmKY
2rXlDAJAT0HJ4BDZH3d5ocKCUoSeTDadXfnYoQqNaFPzR9BKNJtG5AwwUeliKngX
XUxi5Lv1JRknzzI2Siexc/g7odnt0rG4doyuNiDn5v3m65JpWBBQPteUCNVxrAiz
UJSsPuqJkjywhsEune8d5IPezC6HMl+NTGSInM1nfpMYctwDrGKT4r3p5fJxHw/i
0gOh0dYvLC7uZo4ZRJS8iX2AB845/WNy6uvMQVLjCQ3HeCchSsDwn7/VGJOFxmQV
NBzqpIawZ9RK81KzznQzm6vLRwaPcUZyp/L3kFTVWQPa4WabB6CBiwc+qSYJ1KIc
VFe1Y6VaAqctoFpRLt2xdGlBhi4X9pwgdUYikIOpdIHD+/vzSwZLosxL1k/cR95q
DcA3ZKLFXMHfWB+3/L3yhRWGpm7g9S2X12ez44dWzgnwt3VuPr3m/sTM9ZaKexo/
VidSqkveDqE5j361EnobD/Po8pGhmN+a67Gz7KMEc4FWRdrLu6sEfzAKOjGaH8qY
zXilxxiyLA2ecYLGlhe9cvdZuwUgFeUTvvLWEE0P3a437+kZvEAn194FdXSLtFCk
tQv3hleS7S3a8huzv6+iOd27R7jYDJjQ1qOQ2ORKnrsPThp8ENhTDYdu6VmevQ29
ckhb8BC+VvT0cBZyc5AaXpRAV4arEThMK5OHzBSoFpnRS8pVWrN2YLggbdLPLBmw
AWs78sq+XEO6faEOHL1xJ2472LtsCb4jfUFS50y6XLEZs/XgXUeyvMG1BG/c63xX
6RQb0YoGcSYekyy0LMU+gzISqpOdNTw1WMwWgYpuGckpTXMdvookH2c8yktiySHS
pfRMIiSMTSmtXxhXd04/LKo6fTEJtzCmWuV23rUj+AXMfCUhIAODon4Anx5NlqAd
mwEqhbHLHvNI9byeUQXhIhRRvEEKg73Mscex2Al/yGTcu1NHab0x56pD2L97CC29
odaDJb5u6B25R0bZkFxYVuj9afEJN61IqvBu3f8wvYWnajrWt6Vi4lTBZtxckfjg
yW7+99VQxZbaOZM57nK0m97ZIaOoL3fbqQfu0v+T1E5AqDwCNtmMm1PH/3vLBK1c
yqkryIWexAqlohuw2JjZMQL0bFaoRzlGnL/mKfGJdoBf5jyg17jm2eqmvw8eoaLb
AFhSxtSl2K9MuE+wsXQwo9OptutWpufh0T3l2TfQQ/liRyazdjfMrMDiftA8Hor0
eYqS01yEHnKRvYjqQN5K7JeHdT4lxXy8X8gNSltbCPfNW47n5xgFY8y4d33L7r3B
v4dpjujB2Mtpl7qtcvNgvEVnhAE8OV0R90pjcgPNM7FVAEDpe3vBUdyvPjyBKusC
TgMgVyJxRyBWaWj/GCebu6axFKBycZ+WR0ktKF3wA6a+FCq/JctdpaNI7UDuUGOR
vGkWoxhwZnSnKn4gAHy2GrXOLv58QfzdphY9EVwKzHQ0X/hM4N4Z33gTbkFqRq6q
x7X4FQqLbf1hlYlZVFzBEkBaHG4lCzJ+GpNCqIzsqCcnOmOlw7vtfvrl1Sp/R/7O
uIwzeJMZw69jL5uJUdW3cXZaFimuRxQ6w0rs0HJKyvvuOXqFv6gzhdaO/b8KE+zf
KiYYxq/1OV/AlcmivGhccR2zERB33WDdhOG9Cyeg61Lwhkh6y6l+X71NoSHtDIh0
YYxh8pNLrACO2ajELXgCNyyVZG/Uq+9/4Gl9Kt1T/x4C/x14w1yGd4ZNXJmnFScD
rqxXVzm57170KXXjpZtnUNYVT4lATs0OvDVeREjyeYhzdrD/ZlwLu7DJoZ6tu4tX
2Pne+l2ukOB8uNsIha8wSt13vM7yRmsty+xAbpV1kKBxhF4wNhhG1xte/YO1Mxoj
r6VxKDs0qRd+bdIKqN7PgkH5R80zZloljFhyurj4y8q8FD3rmNn8alNG3dRGMxkC
5fvcQSLANYr1GB6LI1D3JBJwm32DrEwAQSLIT14Clh7o1++Bz/J4g6UFt+d5RsBw
zvT5vs3JL9Nmb5Rg5EakFJtVasYSpRf/R1g8GDdk2kCawHMHS4Xz1VUYauB/M/L+
HAeJO2ipsz4nm9obiYb49lDbWN8qbDKm0oDx6g1r92yA8qlDyLyN6/lWH/sjdN/V
YYb1UoL94KDRznVJ9dfYdcmvxGDGqWI6PdtntREaZuM+a3dVpaMA45eiXdBVE0WI
Gbs58zQW5y7vmeFGYvi4gYh+6sCDdNRNjZotUPuoBhJC4TU3ex9zGLuZtBjVoUHn
qu25Q7+H0xaL2mUrTnW0+j9Kxgv0Z+/9jp6mQBTjzcw9aFwEw9rPUCgv+e8UhloF
g9NbxVjzbz8kuors7BcXrUwLkPl6obme0JZbelxWgLz3lOhVba3NfC4uhOzuVOA4
ru7AcZCM3iz2bTlSrfqlzxQ585+73vxLpgf4Mw4Z/Rod9E5aph/XI2axvQPjTPaM
RuyPbNJxxiw7p995hgNxxiX8Jmmb/Mmi3ouLbY9IrAKRzewBP6S2/ht6/zizmgXe
D/wVhdwM6xWuPll3osPysY/csofaG2xmvT2BC/indzBcZXfMA6Hr7yUzYZaJL8R8
2L56QwwVZgdH3PBU12DNxDBreCwoKWK/5UbtA3Jkmrpe0oPyUBGWZiWmYKnt0ji2
wJKNpxUGlq2yyU8P7M9WUmgymSGTSj5mqwNbNJ0sh2Q7K7y8XVeGCsvfLleWM+tu
77lkVxAewgpFWJv/yJ6Wxie1tBjh80hO8o8it3aFuPWoIEVQ0YkdNQA4amr6GFD1
gVsbGXNOJ576bAqrWfHPKkW0KFkdQa1ZzhX/TQH5KZd3buJ+pPaH8/YN4+LI/wwW
AXcBRmXpqbPHS7KBuzgQq/x2p2cEO8appTwmO8/xgoRLcOzs1KVlDLY6KxgRFq9g
d/olgVnFoZzzlnvzPCaXxOrCPj98E46ffB8a3UFweaDlHPfwf2gH0Fs4R04BAmrN
MOt3vHYVkhg/S/06HSQWpkhZ8YUhCSTy3oU4YreewXR0NqlewBRDNovBr0ryNe6y
S1K0rRJy/suqoNfDuylbFV9UgNnRif3em5uKIbG5qkRxQsAMvapdda56XH5s3d4u
9/eCAJQB4kfAZ1bb2pIp09dqML1z1Z+7gIw74+Ln4h17PGL5NHEdmczAt8jAg5cg
Hl8Y6uViEv+FPjfkoLtGnR+uEuU5/eD9dGoXLixz2x+KRUn1+NlSDm2NnGuh+4Hs
uE8Cd2NE+I+uTOkBb9ywm1dKQoorufi9OU/OWuLyYaGS7ne4YlPvgm+d5ieYcQCp
YhBbK+ePJjucQYmsVMwR7h77gBf6OEiPYzuCTBrSshBm2si+E8UFiFEXq+tzs1Vw
8tBUyLoeAebWTG0V2Bk1cs9pyG35BEeTe68JwO6RXlCsEIgn4jKOYHpCHRN9ligx
Pb85ZrkBlu7Ay3IeP7TnxGjFFQQb3esoSEX/Ya7Ya/L7HRf1vbFoKqOROblMbyii
GyTg4q41NqqsOjdd0IHziRNEgxdTgn76n4YCo9krw9N2BSLb0GhQcYIZrc7N7c51
MegIQIOXA0vU+uSJUoIv/05al2FykwC3GEF10y24Pw0rg/MRJmBPiHfM6RWTHjlq
2DhunWbIbR7LiKrweDgFGjM1Zu/0t09klQ19eXS6u8dsRcNBITTGfZDDHdbBC3ZO
oCBntlNH471PS4S/GLXpxQ1hBCzopxQo2oruF7VtLMgxDXbXDvkSlMC2E2nHOJ3H
DxhdTHLtKa2wN8Rz6zo8YaC3tRTJpUdOECDnQQC7eZLCVRe/PDEnZWE4VM0G/yA0
35DbaToqUQ4SAJLOstB1S7AI24X5yH4tWIdQVEH4NjWOKvg38Eor3qWKt6N/xCzV
X8O9VT7tLFJoBD/bDxFpz6Pb0BN3m37T/Mtids4KHTQZWT7HFMCrGZOLS/acXF+/
SCHbSSOUVYjN6w5/FyxJZeYK+v5ak9Ar1TKS2KxGGDsKniRIrUz4Q8UKp+W+0r2I
twfDE4Nxd+DgO7lCB0StcJoSYVeMD7/W+Jo16fwq910KDYoOvwk/bxveRtlYVdNW
JL5cX2QqCLBYqDUbZUi7WM7LFJf7yxadFcPmqIAd7OXrClfCtSQFSMTkPT0EU2qV
Pbg71esxow51/9NGMtYoHuK/oChsbXP27jK7Zb3IsW3RfNgffa2TzT2kHl0PPl4t
Z61/+ow8LPGZOOhPM6OvB0q5A1zj80G14l7CLTwiPfUXz3nKkuy1dvtVlIvAyMCY
P09Zpg0+4VMxpGetfMdeLY520zbseSFpNpf2gtlLiQi8uEu+RZz7ofIA/IANDKmc
yTCF9QqeKy1cG8ji0cgN3NPUo2so5W92m+VzSkOTgKZY+1N8egx/803n6Ax4yUm1
9xmkdoWYEJf6xM9Pf5uW+fxIxIrEHbei7VASWqmGN4J1PH3rddT0pTLznhLMhERF
7EN5JVZXcVf1nKnGE7UX7Ex0PhmB8mW8/69J0SM/V96DSA+2gAwJBglvcJ6kMZ6O
sABmkpxEljnJrKvqQWdbj32UckwQ/x4fpugQG1IP5ysyxHFLaKNJUcL5U4TNpXse
ApmWPsA8RYsvIcNjFA+qnnBXjl2MCWpaXH2sz1R7Qara+jSCpEMpwGmOJiNHF2SF
21kTY7bhOXKO6tOnwuoKhH/H9/RSLBLE08DRbmLswfH3TyJg8OcSLyMk2N++RuIm
qUJ12PMmVa8fbFHRlkiEMw+WJogSCiyp/q4fzmgz6jwlW3thPDaEwteOwh0jodFc
0DhJMyoitLJH7qkTRLmWrSUiYRvKEkc02FvcqGAUqd034mgmLX/DJ47EW3JF2q6E
3eV3ztN2yCBuJZx+Qcgntg0llcl8UjTbUyMK0IDEgIuTZ0Pv5Zj6VgeMJcqc6Gns
5g9vkMOY+9PduaS8CKV60y65dpDHaDVOIj9e4hYmum/lFVKtK/+5QbN+DA6ewHSU
MLQCY3AyARCuuAqMRjMYb6TWzfZNTPBrJhVp6U5dU0fDvwmVDS8UAU7EqwqCES42
er4+u0x12yqxjzKIke47enyQrLf9gNu3/MqYkLU7fGoNRDPWoK91kJ2Ia7MVV0GT
Eq4q92vaPYPDmBtG0QTNw1E9iHXvmi4gwDWbH418FzInhf88sLKA5M4gh4ZCPY4Z
7pJBvjUJtayUL5WeEN6BzdoKKmzLYZ6BGf3d8S/vp78//MBXkTmyKyR6NC7ZTpX/
JsIXG6V/oYx97tVH0QXMf5JmxvP8D8wwEugdg7W+K7IGF9TzDMQgFnSb4sky/xQc
r6IMVFfqDoW9Sq+aOyouvo22qHZVJ5rNjjYuA1/hjDocwy2i2aHQzaQ7W0naBOl1
9YCTUqSy/3wP9hTDST3DjeDxn4BmcB68iFrFYUN/PcoZoGYptxUMxEuMkf5PEPEy
RHzAAfQy2MILsX6a/OXYhxuzYEpqXSMhigQaInJa1DXZjK8GQs/HBNP8KFB/32y4
3Qo73VNn58S1NjwjYu5GRVNbHAOt3yNnolkFzXO5ST3NccguuDp/drTwhH0c0HKQ
GQ9Re0J8Z8frxfmPdliiZ8K1cMMkUwEbY041c7p1o4+g8tzDSH/qk9sVHXdCbsGM
doH6zF5dIp5o5i+zBzmb/RqQFi/YXKxhnEt6+czHRbXgXRdd+kh5WGvvFZEqbZYu
k+yO2RbcSi4mpdsPhBkOSLlVnmwuHhdDQYmYNOF8C9k1EDYk7RdRsgOLMpTpCiYv
FwTBHywe4dyU0qyH1qWxPG8iySkDpmbtgr9Q2MLD/KsllrjOxMEU5ZEe+STGy5bs
g76XGheM19IXCt0EN0KeCoFbDQI/InRlwrkXPWF4lIIj9qr4MCIwcVqy0M2hC5j/
laik7mJx9H1Lz+LKqE6iIUfyPp13+h8I8rI7FHQsXo+s869mkhtqMyJ0FDOa5zMV
UL35mh4hFBnsq49CjN/b//FmSsP293D6dYwFgutQqRcFPfZLkiIx2X5rkKv0KQB5
AhRNz7flcqmwiXZpN4aZz7W/VbjxUNnyrh+EO25VoXMrdYoJXadDZg/1VG6qAWAF
RM43B6tOia5MTGyOLG7dz42rjp5HiUvQwa1Hcry++oJ8O1ghVlVXPROBrIQec1Qv
TkXFaUvISVTc2pvQQ6z7MF5H/thBe1MkAsOt1CR4zvoKDfuJSOHoX0YhTBqYuFe1
0mKMCwL839edZuB/51/5acxKvhJHL2A51+g5928KaGGBvM/iayF5Q4GGtXSL7Nj2
qPGNdvWgJtH6czUaKhqVsSY7dYNwMr8C05E1+kowjGL4wJY+DCyNCrgbnN8H/CFr
o/XeJbvmAw5DG2FtpfBBZ2fDoKWl/uyersJ0aA7behh4ljVCWmAfiwB5AWkf8wm0
jIbLNNktMPLiKsBWm1Snw1e2Qvj3ZZfg2RZ1z891Qq0o5mRBwkQwUHAAKKUpNCoK
LJOzfUJ6Eg44VsfHt6O9hTT24J+lIvaHzBTKsVF9zlHmg30EAmrnAa2DqMAdS2q8
a4DL2hv3iYbpXWWWV2qMLTmVbxh7/+7kZ4TjzkgaJIgEVFekG+gU3cMcCOpxkrHG
33VhAv/8F0d2hm41NlCLNf74duLhCC/jEDUn12fZzvF+xmco4N/Bk0AzkJpY3qCx
LmhS354KB8PvBYVOd9Nn19ONPRSIYVwVtGKYhbL4Y44Qcfkpk+fx99q65xpZXQJS
ZGmpHba73i9ZH7fzR57bUJQ/46sQ5H/GeSlPi9wUSmqfNJgTXFLTXtBp+/ltcRdX
SQdpKDqi+aXmmwPpivzpTO4sQhkkAWvazBjzE4YUNPkpgL+JbzF8MtnHtBWgLQ2U
+aSnKr7a3mb4EEYY/Uilrc8bjB/QXSasrnUMU2bK/5Xgw3pzxOp83iHnwrg9oYSP
IvnrBfJWhofnxXNuxH7wL2ByAODbrsMUBp1au0W6EC/X5Aklx9HrLnfRqVt8e7tt
FEYjgJJGRcSv3c/DL5t5zeIQZ479sbmLoYb85+B30nZueowbWys9T0nwgY+2IPDc
1rQ/B7BmFvnxu4qESf37GwV6YjegFOkqWwTJevCzLGkNAH62iwHlvVNrhPJU0jdm
mj0dI06LQALJ1lYe9H1ta7MerNE5cEqVTpl9mZaRrlwKZCJa96SaGlemMsio9iXU
/evbFNCp8FtGo38yMBztqhT1UTALgOkbhTy58EB/gq12unqaiPr4SgVrn4SPW1qb
kGV4MmMnNz1D+dUutPO6NYFg/Np6EjZl4dbj/kYk9UUPfAl205dnq0HF4beaNBUO
lrACU/rFxL+56DikAP5srAbJjibkXqHjJTxHBebC1h5rLgPhGxhqX2L/at8HkZGG
u+UkA+0TSXnohSrlmc4qTsTHNlYSogyR8DZCkJkEfihiGnMMJvqkku+QhA8STFsK
RnmessbOHSMMZSFSHQAwDPDtL2upYDX7beQGiv6Vd0FenDkiLkqyanloCXJXlC6Z
zU1I3We8zogJN7vEqL9kcev3j+dST+Qio0z695RGe8xODTAUrniqsxJOGwHSy6+s
KCmUTDvtaov4lSwDfCXewCaEhyF5pPjdO0UZZ5muYrnyKMN7ax7XTJyfRfxD5ecf
Q8d7Jo1xtBN4foqqbdkPNUDe4ugmRN9O46GxYWAKPWEtDDa4RZZmcGq7LOc8c6O4
aMJBsbiOzIKAD8G491lIiMkzCAqBLJPDLxdz28dqTiKBw3sPRJ8f52IM+Z3jjbQv
HtaTLhxpb5tU0CxHF5FSe6VRu4OkTOR8WJcRNJkg5M5Hw6V+5Q14vL0opu82GJB7
HFzXMyDZtsU+461Y8VBpke1ixVZaZE9U71ufriYpfLQ7ADp1UcwZUsa/Vlz+ukxP
jLY6QAFipSqb8UVghGDHzKx9jhQH9ojSqpvo13sfJtg/BXFElKui7aD1Ml7GwVQ8
Qggrak0/emVDF3f3ElbuxqkvLADrjphRGARd/syUxiWSB9PCRORY6JfSoW9+6VWS
7CTrEXmqxAafUonmzI/cc/k1lVYSI1PxcoAf2nXK4lkByAqbByZ9uYb/okTpcPck
zwceHcssjzAKyxvFDgmqbHXcOKsSEsqlK0AmLFQXi5SLNbm6pJiQ1NGWt+vWD+Xn
We+BKswkLcbC4xNbTf7zKqurn5K15A36gTtihwYQTgfXfKyZMQ3+DJq3YbRol/F2
mZ2hJsV5xnAcDoIpe2+HM9itosVHgYTou6klYZgRkXXdseAz9YIHCGMubbo0JWRU
wLeiyf/yk18229dgv/UqFgTGCUj5aSeqO+bGFJDi6SA1tUtUiwRPgsSaeD8+Sbf7
Bry5Cu0frt5J32ZAhzr22JBrkRbOBfTXWrDuTD3WtVfGNdbAS7EfJpGqwxAXO6k0
YteLsLrdDpOP9h1NWYZp9EfUxGBFS34TEDCMvHaAGy3B8Wcummez4cM/IvtQJTxl
44lDf14liWpIXLMnYcl0WQgQlvlwSCh13XUGxJi1/PP3iiVaLbcmAMftPAdjM8If
Z7FImA7XbCECn4Fwmyo/VrDQ88/whltn/n3t3YrTULgK5vCPLTfBGA/RRFvcC4fs
EQdHPYb9Tv9QQFwmYsFeirY0oq4g0UQHmjbDrgBhuiL0xMezysevTiSDwP6TYWIR
KDbCmCCNZFrxCngylQXqzquNLqDTAUTncmT1koTyYKb3j73pFX9i5s3ePtLLGIDE
ftI0y6XMhdwFaGb1uFV5VYPeeV4jywuhGFK5aWuccOHu45Xf3ao0XZseVjXGWKKl
xYn0m1txw4sTjUJJBhLCzi5S92kcFRybBf5RMc4MnpLDnUk0gw/OQkCgIauARrBM
U4NLFIb02Yq8HMDsFvWpIoWimf2WCAUmVnTA+La/5zWgqJGr6sIpHZJD6yhteLb1
BBaAiiB4QFwOZgad3/Q+SFxAwvH7iGqOli5ue5x8EdMO6YiOpV/w+JYI+E5pStGl
kANFeeT0zKvUWubsFRjPnd7c4Pyax+VkAIPf17/3J1axePMqsvlA5MveyVsgAUNW
QCq8ga12eSdyamg5hpaw8WejyYm83dPRhyAMhD/teVnYgXtNLJrIf9GZpUp1a8eD
8jq75ynymxJmkP3tZaKNShGNjoDAPPLN1TOIaOnxDK4pUInt9lmNWbSTjnqutyKn
g66JazXki+y6etpcK+rqKPcGbx8ae8h/gf27vMyYEcO//xJtJFofu7rAqX6sRx4b
GMvqSyJ8GrPr9uq+q8O0V8VEh5k/a3leUbboLFZAy5PAq4vV6nA4+6j3uEODwd8T
rjOa5rOZy3QAtWmnR3w2OgTw5O2U63rm8DoaKksjWvN05UG+QE8+vojApW8WlucB
dSIwForH9esakYSRUFN2/d6ncnV7Q6r96EIQaXMpOW8Yg9bFoIVCWxCGLQKZLPOV
igay1tokznvA6mYCUP3lH/k3K5kuufo+s5yrTXvG5KJIubTK8gx5w8afZpZpKHAa
VjbLsvfBytKINQI4SbRUsgrobYJ8MNzs4vWd6bX49eQ5u6UiuJbN6amhDQK3THUl
60n9kEuLSUq18JuHBpCErqt0DQnxI9AhYMZhX67B1WE1vf2pNt7uezKk7KIyJUCU
huQa4pGpWr7SLrYN7tgxoZoEtg1IIuUfi8iYo03s3X1ZaMm3jfFV6lBFOBIYlP9L
/lNYPXwtlVZaer2JhAwop9db9F0YKWWeaYzZem2qTuTDg0o2CBPSDUYSFAdVz25E
wTKL+Et2OrDjSuBIVl7lphJKwK6F1xRDlZyW+2WvGH4EOaQl/JLCUnNWf1KwfNLU
b9mFTlDbPA7Of/bVenKt0iz4lFyLXAclABsu3LQ0+RezVUrxYPzVgGGsc0t/bhJG
pOsJrceNiuPvoJ4MiYQ2fpo48wlbhjTeWR7fe+9LNQqepHqIYsKp+2smiSAP4vS/
f2NudMqpIoK4gLrMa/5T8tp7//CrKYvD1kcGKn1YvXVOJAyj9GPJnONe4bOs9BrZ
7WrSDLb1gR/We5Dvp+Xe/L9CUxHwZ14YG01nf+k3KsIq7WCYHorU6K+3pTGJA06C
FX20xWr4TMY1aTRAvvS/Y5OfSS+FS+T9Ju+FyYqn9qhuB08jxrMUd0xGZN0GfRsb
BPcVfLPpaFRytc0AgULAQGCsvsFerNkLq5c+jo7jnbgZFU0MeHQ24NKgf0IoEcvo
Sw64S44bg6sAgaV4Gc/xVlPnNmpqgxnWR27n/gZgsPHP7K2/i+fZYPE/AYKw7YU3
TDKlnj99dJXt6QTEinzZBGoWyXvRiCNiG0pUABzU1C5a/ubuAdhWKGXJgG9WKh85
/+IgQZ2id1MIAw63p/UHC7SgMRMwSuBo5hPP/CxPq8sI31NQ3hXKH+pmohITa/AN
78UQKRElUx/YbdDUkuT32sB9zP9C3xhMnn4Mk2LCKSOrItc6rFd9G6KXAUOxSXAQ
7wZ/+/yFOnQ6fWPZEsq9qUXqBFwUpsxFVDHdyVAhlYvKZqT2K7Dwp+VRN+gaMLE1
u4t0YjO2Z41T13VLh3EZ2dptCd7/O+UGhTM043FGZdOe+hy7RYb6BCHWDcIaxmIt
srLb164X8k5EfD2j4TTQ+Rraho4C95y6v7K3f/9Yd8Hj0DGwoiUl28IqqMnKWjQK
4Np7r8is0s4DOPLVggzUyEZRJHMb9GxaIMUR9XcdEMZeIrfZNw2OeYsX2hFoP51c
JQX6yMgj+9U5g1Ezbcl1IsywtFWSDT4Ebc4epcDFs+x2BjvlUso5FbiFgcWbP1l0
DmPZKly0MlfEsv1nqZuXKIjPzT8v5xI5kwGA5a/WDnGKme1DVcOAx7AufIVYaf78
OoZenTferMiOl2JYtj1m/cB9kEEgRPwhOjDJO5az66otVDiOkQj1tM9lx1mkBfUs
Gz8GGMVfN++jrSQOuSll9KGP0J4lmstjp/urNjJ8J2/M/JZNffiltqxJOF8g8hJT
vOaod+Y5qV1hAmtDFs/vHEGVvbMYxLij+HMXI8Fyvcq/tDAOj4bSCQDcGsM4tPaW
6rrH0PGZ7m1vDm1euxkFi2GQhzc7dl+5a6J+QqPs8gcKFF/bj1ymdxMXT6xHmSLJ
p6zKhocHE7PTPkwj86gjTf02fFxfstCpXKCvzwKkR+wQxWkJImluV+Ncgd/vcueE
vAjVVRmXuJS5Vu3uDrAVB9SYMzAlx6xkpKL1zE782x9kx+K6dXfDiyCtx0j2p7IF
LWYhZdv5iefm8dGWc04FSjgqUZzROaU8pqE2xwNYvX469zLqH+aHlpqmko9sbzDJ
3wXsrNeQiNp4SA+k74FCbsnqvaWVbsKyzxUtkeAhSrs0Zy0LNvVIuOkrCYKJQzPt
OoPQaoBCQPxyFltHQJMq05GKsSqV7hJqcM63jF9tFaeU5FbHHTDuV8TSC5Qn96vs
8FdxE+oJZ6u0oDDCk3piz6MLDzyXBo+/oEccDnmeHIW8XjDjzkUfI6z7DmHkib/L
GsObcZo9pUHP55aJrnMWUaN1nhsOXO/m6CNOa6Xl1Zs4seTD1aCX6B32naTbOEkA
D2e+xc2Udy89VZ2bD/jEKZ0Ijh0KxgIowW4V7fM5DvlU/c7oi7Pnsv+qa1Zidl+z
Gr67e6t8xsV45l/ht6SOiV2/QKgAd4n6vJIg9IakighcI24X3LiUzRJAhj1r32jE
KWoybHQGHDU9x78f0iwC4s17tYMIEvbyZPlwih+ILHBBi3ZihVdHPxup5dxG1HfY
Sdu2sPZ4A6e0qnPjJlPn5mvpy92GMb8o6u5LL4mw7OplznlmzIRUhNSXDckA5Nto
ev29spKfU5EFrzLirjczatmagttdBG/3sUfBxZ+aUUTL1KpYa7pgsoWtyi5EPwTH
ui1eGHtEdtgKVfh21xeg33ytoAeRxwR8nGUhla31PD/lTZL9BnHc+C/xuuhUFdra
4Ey3JFElInTHsNZr3SDC+967vqQb+zi3x3JA/R/xPnb7NNpVLwAQsC8FbI6Lrq8P
znsYtPMuLmeUlWhHLoxTQ5DIhAAAOa2q9f+3ed2KwAzjuxDaPf84Zak3vaR92Nhc
OvFY1HfB6l/lYHceYOkOlmEIgkAbxW76p3umNEKlX6vIcjznZJRP8UQl7MjLOtgG
BewrsEDaZWPs6ZQadlXRRmRcl2zqTrMjbUmKbr7nw85pT5spZQt4mssiZQFH8cTX
R+ZLFIx+qCncVGx9SOJk6iJBTjqvu+GTy8vqFC2SPteT/KPxW66x6DIKdP/rHMlx
EbhhwCpmPJfqkAzJgFnroRiYUYfpSlhuaT40aVKVXihCY6iAk70yQvOAAtVqblSO
wsjNaAtVKHI0kSqiWA8wViLQTNXu11CB2fYh3N4+QapVcKLBCx6j33Hwt+zc24S0
HCGimS0CoUfmXpb8cLLqGeNIRCkcEkXOkJu/GWdP4wCjBWRp0+B7Cfepj1EXY6YP
QpU9L7FCrv3OPw2+cU/ZRvyJGTI3qdg2g+qD3n/I5Teo0K4XXvjNFB57zD6fIBuv
ogj3kzzj5Q3tmNYkt1nGWkAJCeN7vBQiHhRYGS+wX4XtIvBNu+EYAG0b8NC1vzsZ
QnFvhBK1Wi7ykNbeDM8dd+HDhcBMxyLFueHshBtAcv24rub5uVG4UfuO6CIfTGdn
ZWPGtEScZwxXTMaUexaceI/qIb7pnC/EkqYe+zPs8DNOq2gehUc6tU406yuyzGq0
jMu3UW+EprIq1EqOax0GsDhBTw5c7pGHTKUpIPNzhIvO7zq1lk5hz/ODRJagJKMg
pJ9d+b7r/x3on4Y+8wgS3hk0MptQVUMN/K/w3uRI0STMLZ6kuQgkHb7o2RP0lKQc
KuVgU9Z1l3HvPdc5LhQeHFAvD5qXZPjdj5z/C8cDf2d9GQ8NdOh//Ux10RTFS/HE
6zkKyg3RV1Q41VQLJ+aAw6ocgYdgi9QM7eUrIiGCwPb9mefAEKgQsA2M5pIfE0H3
QEsYb0VLgwEJK4LA7xrOESHul5Y4j4wwbEjAzTfZtvYNa+0AdW+REW+db1NI7meI
6Xl/bkvRLeFeHXoguANbqX+0g9+RXxb3G1IzxZWZiIED+n6F2W+tJV4AzLN70L34
c8df74L59s7aUOPTxpNWDXpEe/fCR6ZdNMfmsj5038BxuIWIt4b+zEQjwd8AhdjP
GSgCx4TueDmtY/PjCFQX9oaRapgV6auYy2hP4YSil7LUG0bUi0JzPlc5FL9b3Ktp
6/7iERoQSsi9EoCBc20lo3OH7C5RlUBuEHBvxKti3yCx8dQfyrw6nOKnOvm8Yj4v
0uTZ2SQ79weQiWRqlZ09FoChitIw1/Q8LOEAaPKC5Q2z3hXBx4JkdwMK+hXwj3na
tY6rwCrbhFgzvAJoEPavYi4d/rHcmGcdJJqm5boOEYBp8bG9SZtz1VEstygjKyem
x3O2gCqGoU3yQ5z4WV9LZZ6/5pdFiKJ0PxKi47PKOIZD4e/QwGNeT8drj2CTd/qI
TpkBFF7NcFin3h7atmE6qz5QKOOCCYZgdhLL44m0gKjhzDI32edEIMXd0wpdRvTl
igcpzPm4Y4OXwFRWh5zpIoP9NVoFWjDXe+bHzsQ2HDwy+obbW1JHyHZ+4BhFuezN
7wrbHFuiN8/J8BFWcyYqhwmiojYCfcJgsP2J92QSBT4T8X4P/bDC9BqlrtHt+Frp
66UjRPH9OkijO8b4R/8OzefX89w+85bukJkHXT4Jfd/67CqoooSbNjhRfVBC7pEu
BMLxJzS/gGXI437L8qOpBGPAcoFi6yxOviaHxiqQUQEqUO1nGmaJpKbLqKGik1LT
F640vsKGfKFa/s1dWdbWZrK+EE8x2u+ZiQ+ldbQ4+exppwmzmUtX5n5urZYgcBDF
9zsK8d1rMJ6cGSyn7LAZCu0BJeAyYgYZiJDBNRwTK2aDhYtGD6GsUGyNBGDjpSHv
g25lS/kRsgIMYiVP9rEFX6uapvB038oDMo8kd086BPr5axlJYHP1XqyBAchJ6OtW
EWi/kAqDdueDGJgE5pt3X6XpVoX1kVScmMzc6SrbIRDHZq92KZTlt/446trSiZMZ
x9HFYIDLIoYIpFxmecgyteF9Z81L+gp3G2mjYBpkBDnYdrjWB6mx0gcwSDKU0HDt
nMCauIM03AC6nRm93TMppjFiNrV1Wfuubeia4/Iyde6UZRxyPa5sJ9y/wem8thYe
4f/UytxBDDJFWc/bnZUarwd6ht1OXKYHd48ErsxKfplceLP4s3B7W4MtSVO0qsUx
f1cxKC/o8O1M4xLGdKqoP2K1uOXNH0OtuvdnjbhsHwCvvsf/PkgPrLG4/nn6l3G/
qi0lWOhX/fZotjQfe3HxKBrWPr4crc69wQJZBceFW6f4YkJknqJ9LsHutp4KkW+Q
rvaCdNrbC/mW67DxTUEaj66QpTF976aFKVItAKEQdxzQZcY3NVE9D/tdXmuFQg0P
RNtCv6RrciMgHQxGtFfUqvhvW66Z6xTwqrza5h+mMJwnJxUTfxOWmDE+Hel+GrSk
UaugKouqZb0TLrPN67CmDw88BEN7kuNIvVilLi6A9r4fcHTmB2mIz/AaT4l3gVKO
C+GFpDzpTAtX4r2jDypdSN/H/4j9XcE2glskb+U2j01pjGKd7OcBbdwAuogs4QAt
rY/yZOLHi7SX+Wz4ek2apCXUYRkn2dO8ojmUTxP/msnrdv5B+QAs34KTYq+cVaAE
FZyZJb6G1ELtrRKtYC23CGQzvlGpLytF5i6EEI4eLDlwB9KHACIZ5/kkRvCbR7Di
zFI2JCHsfd5HR7xLnfRYcS6vM9IEFRmpTBW8zIkH+4z+Tw1BjAA2moxr7v0abYI6
MC3zj2I+qf7IUDEA9NFIHzi6/EHYI8wIwWX+5dwU8iQzhl3BoE7BpI2TZnnDCChK
yzP/bKSfdJDv5n85G6gajPuKA6AdYxMHh/5YeItlU2X4RMObMehCDgZKwtfwuaTJ
wRhi+Y5xdOBAUMyRLsOhhNOBBIJ8U4IttgJydVmkUTIrEq/amb9M+XRPQzuZHIqV
NE6kuegHNTQI6jXsiHxHrqxNS4NFNNaUp0RdM7IjgBv039RfX89934byhes0mx5P
GK8WskAJ6aliNjXMz2AL0H46dY0BGtHGD+hZ6oEIFA20Rbe+vPeBtUkKj6+eFC1y
Wo5Vr24XYd/kzlqad2pUVajHlganw8ZKWBL/aE+JTq+/IweMCHMrO7IyzNfkbija
qchIDFJiUm5/YKkLubvjmgu1hW0QBDhGw4EI2NKBhSzfeMhkTyoTJ1+Q6LUT500d
h+4PFq55/llCpozmJO2bmpA6WiX+zU8xcQMa74ZyFexJjXz8KVghDtkiT3dxZpce
SCAio2CXJwSquB5TUfuywIrl+kLoNiRvU8a34BLE+GfnvRPeHfIiwqCUgZIkB0ej
xvDdXYhLnZECDjlCqWXMTAPXkY7B259hzSmExsTwaSmwG9OYBNpoQckZjNfIxy4i
qSLsyD/6ICL2lgNQoPcoCxCZLzYgDf+LOSYArkPf1KX5v+bucAzJQdSz7cnbVDNf
jsFvEqfjIAgCnozfiGwlB08QUKrAGW49mDI3rnQjFzF7sJC9aPZzfSqakExNPN8l
JsbRtV9XBL5ArlZ24iF3Wf/tlEAY7Uh1CF8pn4stq2MRwUpW6enPtFe00eRglIYz
jk+i3gU1rdOr5Km94vzZNT4KWKRUXPoiqrVgdiuMIdlamuY6VuVcSZzs21OGvMew
7XhI1zGkHuI6ch2GoHzQJpjwfMMUWjQAb8lTfTiz/K81iSWcx+1QGB7Qru+Suz7y
kosT+9QBySaxbGw4EQI/3D5u6xW/IdyCx2gY2BHUVbAL452oJ2CYGART6NpcxTww
wajwCYwZhQN5p1iWp1fzk/pbwkOPgwV+KB/RFYNMEmBH81cR8PCWPZsHTnp5IpEG
Ce9BBxNUY7RfrZ0MaWJhiKJV8KBYvNzy2+ajVcKlf09/E31W9iSoeshMrIJ8D+T7
LcevC/ZQUOMtnoUJkLF6zz4U1UPSGSd3JlSNyLqjMjg2+A8ifXzO+OFw8zvgNpki
qKFdyPrzuEL+qcNZgesNzV4jX7GB+/GicQGX857jdeHiapszz8mwqRPl6SZcN8y2
DLcq7FbjOgpmx4tir35V3v0f9j4aFJ5NguJjhiDfUYHNRH8AP4nOvnEGRc+cdNe6
rIOdkFQgrQMwb2ccsr/+f4zRzuYG/v7t5za6ivbFenlTXfH9ZKq+kf5MUL8ebLKR
VWxePhRF4S0KET78az2+lOXHocsxO5kZGj9EbwZ8jfktXQxvBLxZopU0yxzpPnL0
z0p5Cr/Qq5abKsCrfU4AjOMl0kgDNKHCK6bvf8Nx0QMjXDj19FwfTaf3muH+eg69
l+tP6ILeKb9Wybw/0WV1pcfudLNpkS6wOggl7r+1jVbCPMYRFKSZBhqM1ysVCm4s
wq6mZzu2oS1aT74t8n5Q4967TPN8Qm4HOUPSRM7X7VPlwvSO5zYeMr08n2TSa/0Z
dgMk23BDw/W9KlJE8zfsqrOBFa+3isJ0xuCfLB+mMVwaIW2r6CHJtnSZN9d6hHkL
5pxxy+43OCoe+Podxx7OesuEt3i7K2e2mKuGj4WPsbBhDC7jpgoJxA4uSv4nFCFz
RmtgYExYc2TdGtMJi1gIm1cK2/4L3fwZ7t6nNniFl08xa915m/UJK9p3aFd2B3+P
2tA27wefUIcXMkHhg67DGM7NRD5kW5hVMLxBb9C5cbmmn/BpOnatXtQRiZfAqPcT
6khldHEhk+iEbH9LD7fRRS/tMxucbgYWy2V7OVu6cnLZ1YjVMSANoHre8RW9dnWA
MsGDqsGEq6W0jOy+eS5LqNIfC6H1E6d9FdA6lcYNypz8cmi0z86rmbzajRSVPjPw
sV8KVZNk12g+cL1BshPvknxO+gi0U14TcMOJVOl5oatK2NvaRnD35WvvloWDWAsU
bdxMaebnIcOQz8ow63Ni6vjgtoTxE0pggD2+mZgIpVUEVph3V5J0DoCSh1nX483d
TtB0udcCJhyY6IeE5hagTyF/PFNGW0kS6Wb28uFlrkURwLZx8bxYRCTCoQGk65Cc
xwUunYXQ/POm6vBnBe7NzByyey+y09AbgzTIix/MiObCkKjydIjG/+40cPQpF5YD
QGwUpDTYKfr9G+9lNNdymN1TiPHcrhFxsMYAYEZVzSWYMo+DXahbNzyCj9Zit6aB
gd9LrXzB6/jGVfZB0YwKB/14jg+TfpV5BkupjfOQLXVJY8JYrBKPpchl7MxjRs2c
0tAJJu81/bWMv2IsLTXwDWbtg5lkoTDC0lLGtEdMVHaYp5cqK2FB3qjjKrsv8Hzh
A6LfIYTBZAlRkYusvhsf/CX3AdGuNjZPM37EbIl/vD86om5QXneh5ipTf/yszuqv
+b/+pLAF5q4BFX03bF3uXA8TXGVEabzmza53fqo+ugzCC8x8gqWMp9TdaEPBInHH
X3RjEcVbn7EnwfjhtLd/XgQr8V+NTSz/NWwhrSXerb5e02YIL9rqQb2waRMgm1Bc
OSD14EyD1dC6Eo9jKilRr6E9tzz+wKInYWM7wsrXH/eqnXs88xsc8T2XIbMOSbiI
z9qxE0M9/4+XQ9AJKq1jWDW62Dcqo+i41sDUDOJ2Xpq6MlBcRMe8ivzek1YzhIZ7
6PXuhCw5GlAbC5N9+IMES+5K+urEPTGJgesfky6JguSDBfhMbXbPZs7/Qly3cPcU
K468G7YCxEBbevdNvMF3OqaJkJSZZgsfkJi5q3NYFWGq8ev0NDERc7+4Ibwd59jz
V3KX1QHFi4VNq9NXWI+kVypB04c6MR31W1S3k/6md4WvS3of6RP6LgYY1NMxsfCm
fTMoUZIhgzJDeVaYjmeSy4C9oVxeStgrsexc71TxbTv6UPLhFTfF5RCNV6n5/IiE
f1t/ddvICzGzBBVloNidCtBNM4WTteV8BHmo9m+ZuFQOJ0P0PqBx7pHZmapVCaNi
6A8IHwgyRdZGgBNnt3sv4iHW8CyhlTSbMppDWEA7qo1ipIz/Ktt+2/lo1Q1lDZTr
gsoRwNMWxkSOe6YTlWTwecVoBs+fUHep+GIsCCN8Np3+Ij6yQFP7CbB1QHL/0UL4
CTPZryIZ9I7GYDMPhakbrezT+Uvh3iBr2sCfaZY7VW6x7eIisSeixN2/z/dDmE3U
jxbJipGbylCKOltusnLEnduOuXPuezgUbDLYKIe3N7B64sQramdaeOlV8wO73ldv
DB40iffJSviicK6gmP43mDPwSqf0oXqmr7mWSPq3y5fo95hL7fjntnzLXnisGsF5
qzsT1tNWrMk22m12sia4q+RA1xBaEYwPUTBhIUqxL5u5pHYVJ0Jlgk5w5kCCLWrL
zBEwPWMB1MI6WIjS//X1Rw13yilb21CDGCp5I8TN0WDmiorW/QO7Htf1kqkF9YIN
We0GPIsUSCIvpT2L6FR7Y7hjqtyQDTIn6930AMkPJzu44rou7uDOesQHu1Mm4u2C
erghyAqAZpyghrPcM5/ER4h1yKqPK5nJ6XnRy+U3uTz8ROHkMy+Cigxep07KG9RF
a/G8SGJ3FVFnax3cjDWaI/PbpoUdRYVL3RT4y8nHASogjle1P2JZ58P929GiHo7Q
8meeeKIE9FdM2nXR+t92XM5HAhDFQJYgVosBblCvjr3535O5H3FY1KvmO1Eig/Xa
AQlWSJgioEqRGBnXjO7zk9q9jLB3dDk1c1tfI20eHuqi1FYlmAgjA2nq0vRsYt5y
Hf8niirv6tksBvCAQ3ZmQN28Q+PoN4R2qm5SxqfkgIyVJcD2y+79Nx8Q080KukTY
5DjMa9mvRmDBpIsGYFRA8eRi9u24VkCkUr05nyXPqJEXhaJjqvV8rQVRW/6DbQT0
86Q62H6vxpyqn9cAbZ9sbcU8cE5qUGaKNTLYh3zySNmCxxqOCAqPWiZ8ZUJFA52b
eCrm6gau3pRtP8oOzemh0RBIZvWmvTL7sjWRXQ5pax1BlWI2xkHEQDhR/ADVlJbm
BN6usbAkxEmBemo9OwwMLCYN0/yCSSEzLjxQaHWJH4kSaMXQwu7UN7aq+U/nbwVO
1PoPahZ+OzQxoQhTX5nfMjOYvLWcR3dn/2XEKlnzo05rUO7RtKdhXI8IgoaCtW0L
edcLaCgagLfN0o/sImcUeHfIZGA2sjDoLbmZR8nmapmV7Sz7Z5g0j5Ie/BqBYx/l
dmeigYYoj+haHdQfRMa6/pOnkydA1M62DV2D5cqNlyXxOP5zBxgXvRvcFqlaHgj1
drLOfW/FVDfFdcabnZsCST12s+QkxcJnI38CfWBp/wS4N3sv81KFsbR6Co2zJmI2
+API302P9NpeHEKhrOETra4ZXsn8EsTVy4BCtKEOshxAPh13vI6sRhNSzAYeR9mY
+Lwki6P6WDtQZK4OucDmCodMFtPRcUYon4MIx3196f5yhht1LSnALD0JFvnQUwMQ
hv3wHlnJKF3VlpXbpsoXJxLPiEkMbbhV8J1ESBLjDApWt6CDYMdmx9gg8NseVofA
jhSvpC2G6QNSXsdQRUNS9QKfFTOPRay+2GfhAPYeZqaW+ZT0KMp1pg7DnxWjZf8T
FxvAfJl70sMJGibKTDWDuCosCpOBhbv1NNyJuevjXvZewrcxYl/3So8bb5h52Lti
LHWrMBHgK+wdm3CotxtZOMjCfNV98Nnsv2+SQBfJdQQlWD4y1hlbDgIczJj0/F2z
hq9Jf0hmNhMBpAMsuxf3wfMutM3YtMnhN6ffIhl/+QIKIY9KQlqRF7jojNTQp3hr
sDp5DmCwnup5VOWzfov/IbJi2yLg+FxrDsGXz6Sv0YaKUvHJ1YIiUs8cP1ZgZ5wk
83SFheQveqJ62Vyel9P9S7NDiq6NMgSTn4AkUPuU66Tg22J8yegtogUqAnUvXVBb
IuPCFU8IXk3VcFGhrFpYjqBVy+TjslHV00d2goifbN0b/F/fkzYekchiGuKa0IPA
wdIP5xwGboGhbWbniJ6bixaSJe0l1TwhsDa5D1MrOg8fnQ1MLuEnCR3KBsB2ianj
D2W4H3NjzsD0k8j049mnyqYt7MH8jYfIIYeF+Y4PI9dNzgH9VCZWRydXyVkRvBx2
7FdpHULdRs8LI1e6uEX2vbZwm8JsM7qnXg4S4lLsNqH9RUV8Ywd3Jor2sMZjT0SB
Fw68PTZLVE+llF+7uWFgTVA2NxNtqXNRCO60JX6QBuR2d0wne4cOU+56YbRRORCy
j9dpgl5NowEEjlhVTDH8tBr6H/dA7zirV+9STyaa2Sec0jNfUiYyT8z3RVLYKnQo
3iE/1cpzAbvXqEScOfKzAa3D/yoSjyDG78v0eipaODk5fdvL//xJV5eA2WdLJfIK
IxHvPjDGHhkBNyvFRNy2ZrgNoVt5CZCwltRPQc3ySgfi7J/b2SdBFuzS82SKVuyI
r6cQMz3TsZX/ePG0Bpc22Plcam4uy0qrk9gaPojiuxGI2Kb2k/uGfYHhaz79lPu5
7ESipKFga3xLECarqj1wufEUDDHPr4oy6CPQOKPpI3NjYqLNyY4HX777WwNZLbUJ
u+5V1XZ6drHOOev13HywtpnIz4gffWKZjsgva+ERN3VSA0CcN+2f/pTmdykjpw2a
96jBHzB9osvGrux8P6veJASvQyhw65VY3bMeCuHpva86r3M2MlEUlBRkSu+29v//
VoWTWf3UqGwCytRg5fSS0oUjODmmmKs2/Rq3A+ql1zQXKQ9aNi+u6eHlTPS0jiTL
1frBiLQSx5fHl3dRlLi3RiXedSg0pkPbwaN+lJXNpyYSwwjrqOTlIZyS2uPg+BpM
APc6TfaYdpO0ihrLE9/pHLXKg6xpF7UGFEnVv/pkb4QX9LRMdDTs9oLS5y2Vw+A1
S7ACt19UhqOIGhdV+maRQGoqGgDSfKirZwBCBx94l0D0zTB11bpzF/R79UqPnvwR
7YnNjABRyUZnYr94dLmi5RLPXRGhh/8kc4vTCA7cdxFF0mm10BK92yVt+QR3yKoh
dHpElJsTrKIKICv2Ey1eHohAdWyv6oZHwZX4nHZ+d4NKRZH524XnFasqFIbdY1Sq
0zor3OG4m1TveGoI+A4i0AeKFnYPShc/cx4q1IKOud/2NgisM9cCRtuntqE8xrCf
x3S20kWlwXMHO4NIf6Uw+7BYD8GR4egcVJ9DADJrqtr5ciAwGCBWJd8ArimWi5Ah
rx1gcxopGhJHCY5UQsdckFr11A33OhjW25nezrwn58utU2AYPEKGR8vJhVqe+5Tg
pGdNvExa1Yq/5sPYfpv0+oz4IP12gqqPuAsHma9cckJKDcez1rF86IVWOyE1uHU9
EReN1ANsbBjzYPn/sLx7KEeZ5ykc3DLIdPlWtowmHY0uj5Klpxm4FThpHLxCH5ot
Z1hzXxdzN6YXTTTFG5pjgj9s+rkt3PPquy2x7SmSjH90nQPVe3CWCsmsmW8YjSQU
IIbsl7JxsBXejmhIiCUAW+rwJycF4q1ID38QUTgSUgOsG3AxMDRoEfS6+Zwe4YMC
D9WuL8yrha1+hvoBhFe53i/7N9ZjQGks0KHU3YxIy1BCuIsKhjaDFR38Q9oQtLk7
AxPARdv4kh2H0uC4vUoqLFJCgOUaZgefh5PMrvR4iW0c7LB03FMFS0aXhf0bDPsb
ATR/YfLIvhzjjUNGGc2FcNco0vDUPWdx2G210bHwKMMcYzcm24TRFyGk7CX9vLIo
uSChNgd8WzUOYaYO8Tm5N5bnEossLR99LrQSOd6dM6tVvnGABEaJ5fiEzdjXwnRX
9IVvWP56b7Jemziptd/AdoOemJl8H5qc+9I4ldRYO1rhYW3cIE7y2gQS22D9Qxjq
AWL6cXWO3P3JJpjgr5vYqWV7j+PPALBasX6VCjpbbsjw1ry6MZ5sFfhkgrrMdH77
4kNOWTihMJ7Mg5jd7e/Es5H06DkDg+92waPPATvYcqkxRhT/BpR7G0RAMIE3vVOY
NmDo4G1m0lk/jsFjGCyDnc8ult3iw15s+CenLOjo5hNzOpLmp+nklShfozKFrqrK
rCViuzIcS9FrZHrpn3YOOtnxOP8rou5qK7NTjxbIzawgpnzqEjsJWd2/C4pBY7WU
beStzvE5DnIdqKv0T4K0GZ3w3mMamkR1l4kngGbsN1wWOGRtNtmQVfaFStvovuuV
kg0Qs6dWmt591CzrVSOQbPwm6ucJbHNGyY375l7hSYyKbqabG28uwhXEj0usKzFj
xkZx0uaqNP/qczx+TJZ0j0ntcJJew629uug9i8NBOVnKh3pwNcboVoKcmz0v+gfa
9wIzF/s5Vlb/JGyw5sagLQ+15eb/P0dLanXghOQ1cAG+zrCgieRC7fv2l07EygT2
1DmFW3ytr4RvTLR64l8E7FybqishhIc32tVezZz/6YlAHuAKhvVfikks9J0WfvSO
Ic27sE59fPUhb/7Zi2y4PCcLtPHXg8Khgyk4iBaymWHlf+odO8kJr3P5fQoy0rtK
u0sB7FfCfvfpYfaNvXJEVv7nIlj2IV3ddqX0Fsa7d45+lV2xU5owbmjYlMXpqQru
ZwUzgN6cCag9G+H+0SyF/E68oI/ZWqitgfpJRTZELtN9JHDdMpm/y56Wl2X37Dz5
FBZkFS5wQD2L8karFBM/A3ikgM+uXH6N3iI73gla8ISVtmhgPvo4tUo1g3QQff0p
GAwSkxYgAhHswHXA577TURpdlFW5S4u4oJzUexleyy2lXbYbIrptlEouoWXsY1eE
0sAa+KCyNy0ZL1eOgrKDaUQT/caCxQDOWgWNsRYmQmoHWOMW02eDVT1/Ty0zhsyA
UoVmcCNYq25UT7nlY4Gch8R0O9QDGAsy8GKSsREALgPdo2ZOox0m+jsYAZRt88lO
H96mGpThWGnDazTmavTISN8zpqj/2d4AH/sN6bBq0A2Mlqi1gZ/FjJo4GRxWfQjH
wPjXZpb7l1t3niV9jGmrfYvWo5elY+UeiMAYa6y3Wu56AW0srk/KnIqYuiMKEb2e
XiEr+dpAuq4gRlINeMiLgFeV4eD7PHcBq7Tvd5Ij3H5w1jKfa3Afkj/ZEE4eqHVe
aPBQivc/6MsqOBtgc0F5v92GY+ISV4UyYal6BTI1koMq6yboLiUuMgerzrAwEqjS
mUsRgy46CtIH4JsKWcPkLuDvckpQV33kfdQE8A2bcjtr2rE+IXDyH7mdLAZ/VskY
lVbmtm5cpBWaylH04tnXs6MfYIpk+Z+FjTerGGX4OzCXcyX7u4QgZXFFR1cvmC1+
3/qC7F631nI4h58sZlC3s0QM603ktzgbIYobGOOzNTBT0WhqU8XqFk6keZrxVyEw
a2pEoKIgrfgTG/Bn/8mhQg8qgnjtqi7irKildEaM514x2RHZy7pnSahO6hdQoz27
JfKX9UweCliZI5APy/ODSc+McdcKmj8afSx8YFnxpUqq0VRbCEDeK9xCJnqgHQsH
A8Q87qtokxoKgu3jrrgcif1zPDYsNRDYPm0CtNOoEijzWNfrnMKsaTtpW851zNFb
ZdyQ1UerDqquTbw/Y6JI5vgnf9Nyyl1OIKz8SMLD6GvfDy5o5Kt9evd+GHoleltz
9XnjVNxw77ATOIncUMPhKKyrlTsEGGAdNeJ/zvWHdOgRnDBSzZxMf8Vv3hqWemJc
ZwL1adeFpH9Jv65D4QKfr259t37Pl8aXJkvke/bGOcQE76AA0LHuWBeZpjTYEDmb
EqOfseo0rDMORLSUsOfA9lkdUf831QidoYyQZoQc6WlC7RXehtzCi243el8rfAHF
tRmSMmhKKf/dulvToRyRSxnV4JfI3rhPYTKtxbbYRXlNurBCpzfu6FcbFxOQ1pgI
XCm0mk/N7Usl966Pe8LrGJJQ5O7EMSjdR5ZYtzi6xksLJ69LQPC1yswKCcupfyV9
FPsGd9duow6t9+WFr3SzBZnBwquMB/dB0Za0x8j1zggHAv9PJccniSOFCaKZeSAa
Xj/QHmtlYA3g/+LAbu9HTYlC3GB4PyaMX70mVX+w858+mCH/N9EoQrCkQRQy2GLX
WsoZCBM/76dDypW7QtjlcRBaRLPd0+cXU965EPurkYtI0xm6NvrQI/A/tZuEuvbm
6BonX82mppxsyXTN563U/KG9Fnjkro4ADVHlhT4Al9y/ePo1cOVE40oTB6FSoD01
ICnpKSnQRG9VYAI0fzQuacG0zYztsUTPoBRhcKlbU1B3CJHH9Xi6vjznYvxoa8k5
/CtJoe3Si5Lr+I5p/tv+v8nSotnWm/bGMOlm6u0lY2pBNFFGeOIu8OTQ4r4JeZvA
8YkxtZIupsffaVTd4CcpoFq+hxvzoxZGMfrj8XRMTLsk8Hpy4VahnwYKDQZnFPBa
KHZYk9xccQInZE01nv8S7TQNjWlHITta/1nBCBuAomNmScdcqYI9ozAR1xAXs3PX
3qnjdIXW14lBx4acObh9urkCQoN9WsBB2lOAVYOtl+4YDGrDbzfIqsrtE6GuYsno
MTTNeK1R8RTzYYGa8bE3UOiqxQroW7rBpJvwIu+XJbsXLhDbIwLVwfQBIjXJ00Dp
IPnq+JpUesz8gn8zcxyjJOfXQve6Qopvl+chd8uon+jnS3wdtRiU0eWtU9XUQqCo
MQUmu6DFSj8IAgT3tv4P43Wc+R5JaeRI93X5/cAQdFBkVjON7XhVJr1LIMgb4543
v5lqKK8HWTxi8bOcn1oZzDDvJ007Ntl3vpUryltF3c+0uHjcpvMZTUewmnRB+7ET
imQl+lqVAaiGqnJ0zFIJavyPmcAJL9Q+8rgBVzcqKdRptmWBk3GJubwDx2SHXKqb
AiXzOXw+F/2AuasMVgTd932se2sEgxXNz2L6bT9NUpwClFfLLh7OQXvNbGwXLJlu
J04LBRGsJa/Y8A42JOX17BMS6XRBQh83kP14CyFDDDYTG1fT6UfKTyRc6SLXQbGb
zlNh4TSH2C+vvsNKqKbPHmLu5TNIQOd7+dS5qHHqKH+ISPFC9DPktv3147Adjid7
qvbOrVbCQZMZbzCmFoNODu0aZFbrs8Lol6a8wU/S4YvYBjb2lZVp64WfeKDh8rVV
ZT2pDMzaKx+681dZXXc8E5ofFhqvIgzHCzjHdsmDFXrOl6gGPMCiGpJVEPmcXOeT
PWobtrUMzziuFZ3OW3mXhMb2gI+ILZosx2ERTrFpPCxg6Qo0AyJoCwtJVp0JG5pv
YqO+/FRnsu732bfkLMzJ2Baxq5jaYCRcQznAE5zGToGwChCzEFm9thcnlIyjoWSF
reN5QIJN2KOWeadBkI1wYcqZ0mT28tDU4QFXKb86Pv6bhMwFMibKRrGVE14ojRms
CU6ELIJDzBjiP8qBQpWiL11Of6NhGe6aeJTVSJhE6q1MuvPHPqeL0JyF27hvUb+k
RpXYjCQEn+4p3iV/pPm8PW5+Q5A1pUCEtDhaUntkeyEdNXpayn5Z6ik8j+iadmhw
gbqAXzq5kIPzXAKaHc5XneI5FEB0et82usnelgn4/EVOObOu5X/iPHDLwl/fJAje
yb9kWAImjPgu0NS+prw1o3fkVSICLEwI2fFd7hodOW/kuWyO9WVcDtkoTE6DocTg
hF9eB9iqKcm7q1t0/fRQuj2VQHLDzTZNnqFft9FNzNsEGJtLWGq5pqDNzXMvE5kR
3C5/Iu/IK0wLFqCwyb7GlCY/wvgKkQ6SlITHwIU7PdN9oaATgrNyV/+YWlScf8r3
TFaQQn0xUYztECzmD3sidZMJfygHhJBrFNPysLF/RkDIWSY1x8E8rnWLDuc8I35v
r2azqfqQv0b0vN+x5NUVGYg+fSsa78S27BSDctyjIFiYDXNtJQXj5iCPW6DQcgxf
47fLz95yEHWttVX13Mh2c6pcJtnatP5HPWfBCAu1+8nlhXx+RSKscUlN8m5K9mEE
sStoHLSVWd2wLvu9yFSY6WAYczvkZ/+gVGU7YarDvG0Fa/CEp3CIItWU49MEn/0L
Iym9bz69brKBQh/067PZLo4ANU2TevtehZEVx44i5sfZv7gkbDdJV8UJvSp+6SGy
QJ01kR7ZhcSCnZ3guypAnhycQYi8Y4Gi22JgsF4EuR7uoOYFDeDxfRh0wwYAO6T2
AZ4I8qOmZYLoKFGxaVAtEMJc82je/MgJCigofQeV5q6+P4Y9/dLY/H/Fyr2vdKSR
CHEQtGTGl7UvtoWSPIojC/Gn3n9iAUvFqQVGlDavrQkmohQtNhLz+1psBkby05EK
aza9AHOSnCXUecCr675LJx1+bIZRRdIDf27q6mwdxKfyMxU04xh8POVM1vXPdX9d
Dw+pBV+68fqpkjbeiIeT4YO02VhBYb/LDCX5VPJVm5UjoLDCkONQCzZSpgAbaBRy
4Pgd4GxccCrN2BoHN3u7llox/WqhFUhGUtTP6umGiAHRqqR95BckRfWoLXxq3env
WMfyiOK8jd9kmpZUnHbhL4IDxbH7mESOg2j7upQNFTHfXt6ftD2G6mGDv4s+OPiZ
mGQ/hzwy0i0JdMH+C7cA/xk5BVM4rgwL9hIVvh4kv3FUJPbqo8n5TNVCE+6Ir89X
8F+M5dtBDR/SJFq1PhWGIWkO8rLgZxPdtIoQAHEa+PAFQxnz4VFTRj8e3Jfm4PLS
XK1epCGC8XZ6J7L+NPY1U8YrVbkMG5EmTQGPo2UqNKC9B4LuHF9Nlv6uOnJoBcVZ
gBNUn3lrZnrkjEj0K0oGgYdwwM2096i0pvlAQ2CRzx9z1O+T6Lb8AX8Mu63NwAkH
hKwyFS6r1Ryi3FhfPcEQxoHQvuezCNHTyapqmpsNkKz3ht2ywaf6myiORhuTbgXu
vMrvu/lBQ3vo0vMLvnlhA6Iwl+BDSWChI1L6BbmkrAqEsZeuA89yYDzifCI8GOqJ
MRH/gMhdjGwOVoUaIXcJRi3iYEA3jq+WeRG144KmTJMBBqj5QXEEZC0JQF4cyBCG
g3+P5pP5z9KxcBQLCdnr4PzEBdKeoEHEtzuVkvJB2Tw85XbPA3NivYlBu+Bg4KxR
mQUDBHxe/OgQ9ClmIy3ZfFD6lQzqOJZaLr6sCCsx4u3lChBR90fmFY99uQRQlnA7
oynGWZ32vYWvagV6m4RhcruPpuR8+M+hROlTkvRbVzr/BgbjUFcisFf/wUgMnHHp
aO5Y6KAoo8yJaPCo76QoGjGnoAmNSOahxN6ZJiJaADEjxaOHzv9l1f94Rtmt32gX
629fMcy4txTOTwzS/RQOXm63Zi/3g2TfKu4JpBmKSul///nMjQ8cU2QPeQlzKoxm
Taysju83Isz1HqX058VqZW/nKx9NKg0ba2NW7FxH6UJia40715BMoRmLIv59P7dx
MAeLHW4eb6hAKk4hxvbVrag3RxhXqiHBlGZ5xLSNXV6zM+Yz8j9pou0UTlfT02wP
fl7cuPda8C3jZKohHFVQBtl+nb4lvrDWdsdR0jAOXFbHYcjGn+/8WMdTSlnOCPkt
1HA9M3WEDFB+ZXwtcCbJDUZr/06DuhlW3ynG0yPYVt8OZthyNBtufWDp1H5RFdVA
JDE9kLoFe2ATGsTlbmU7eo9BF72sV7iBYG0E0dT+G4DMYAxvc5XDcDucviwQ2sHI
nQU+pzAW9VAE4fGFJ0JvIN4vGYMiJNYWK80YgY8DSnqmT/E2VLHAjt53XGHITSbB
ShGAkaOxI9nWoEfXoIU47XFkA35ZkbETvMtY4xjayarz2NFtAdPiygMG5gNRE2hP
Y/+Tm2w1kHETu1jdOfO2ajCZ6dTSZeIQGb9Ex4zoZSY3sDdm4jcByHaCCF1MaMcp
dmawfUGnKcBUybvGzNfpaZN1xgVl/Reib2N6vvx23lTGj+xVd1xhaJH3yTkEJNjf
JmkrxbatqTATEZdLU+J8pnaNm+1R3nDf0ul2VTyf7l7EhGmvdwmODbwrMvynPS82
TLFfLcwXNRyj2pREU0S74kgdHoBIqtly7pbrMWjUrtjVwKhvdpwtdh0d/aFCnRRC
PChr5HTfSuBtAammidhJlrPRkxDSNKSP8ttZIGlbvB65oJjfg5yLmRTTIx8b0es7
k+iA3ftocaJth33SbCJtc7RV9lKLNCaPV2pUbxkv/quEZlwEZuKx1l+QlfFXLLVB
yXW0+5n/KYj1bJFnTY3gEYZHLbfoWQ4WM4+BvY1XrBkRPjWe7fTJ62NzSGSkhxL5
vGpT0FJ02MvbxN/aK8AHTIrGRkM+Uqrl1jJGG2H9fSUBlyajrTa4onKn5hl8HQw6
epJPw9Lb1m0VZAon1tBWGJiJqofDyzhog8Ke2KeT8xOXBAmEpWVHtrONy3tcLiSL
6WkLMYLtHLG4P+nihnkryQoF0klB2QNmUh0Bi7gaELTxsr3O/5hYLeeQsVGr2asW
vTd0XXAUM8G1bMKM1ToH8EExsB7BJFjAM/V6wFhfQGRmzAPHsyY9J51PzasZNATK
Www/mW68KkpiE/BUvIJt1PD6WhRWsvqQQLmuZpbRkTrIRBs1SaCAx5XA2tn+8djM
rHzfMNqYrI0s7pZumNaHfgbDceRU3wMi21qlCcCeoaucNANCbtwwcPRlGpf0NzBY
wQxNd6H7WS+eufZUMLMhZ5GThZAC6udFMKY/QzGxW4uSSvJED0EWPcSWwY+zGmTt
xnY57Nm+NIJIGEB5dLdtoEoBqvpS7la2wI77YlBKTb14MmgxpTWlh9Iczyrdx8Oy
WMgyJJZHRvgiYE2xciINbq6DaWjWYEdTBkXyrTORgk10QnXLsog7OptYSqTshf19
uEXVXmEiAQw1UiOTBCJUEbFRfkrEFz2/fqCSwEO8CX0FxhIEyrzbl+CCBJIcrnLN
pzqmBT+jS2/t7gEBzE4ka1ZodLHi9dm3YfiZ6FaBuN7dskoeDh+54+1uKhfrwczK
zMWESDBanNszvVaitSDx6L8cOa1tBKYYOxaDkEmJv4rssNQ7sMWGmD6kl9xAgN87
VvXHUBGmcfIXw8bY04BzQaWiLrlrrGmlAZ/IZqFO1ADLOWWxQBtATWCVrrhxuy+e
ImNXGnd1+J/efJJc4tRNM3STmVnZJ/9Wqn4Jagevokm0DFaKW6TXMbRFT9A2FJ5K
Hk9+F9jFSQP+BGfBph/G+duh2eTW4KpDZzUSMeMhlM9xcuX+K7bDCbGHMIIhYWRB
hhT/Mrl11mw/lqZnaH/QQR+7rCx1/UJ9zJKZVFE/64QRd+82RMBZ9JjHJIF5e0tq
gh8drB0cd9cIhfaL0h2KdbW9wHxWOcSHpcei0vXe37TGxB/ciaRjK4MveSNCleya
sy273LQWmUY7lo/8d8OG8+EdcG9yQTXxu0CyFlEO26Qt1NAPpJfOxXqMw+AMkMTv
Ru2zhTXyEhyVT5X+z5hfc6ds/bN6FrwsmAkab9XFFRN+7vy1yNDhzLv71DQ3zWwW
kpbRGkGgYLrAfQePtKgiwf58axqcdOlTvhODoLPT44aCyLQyQZH7yAR09OT4bTJo
0huqSXoVjTOyTc/u526jyxNUzjLNkeGwFS36g5EDH9hdTGrSeoLM4C4JkOecL7+/
uxvy56i4JGdIqRiXmTskZeeSt8QrYUAyVCnzrCsW3By96LlOMiLGgDuKrMhZcPaa
QtOQ21nBKM7dFpa9pYksYELyVQ2x9ZY8Ydfb0QZ65Hixg81uzTvgM7Id5tHqmDJR
bYefYULiuAiCEHBM8jL/3/W3qIoDP4DF/nJK+NJddynO7ca/jVinfcRToWTpKQUY
UdRYlxJlCLZX4c/bEUFzidSTEKTBbde/e+9917zi7kLqgHBtmRQuVM8aIT4ijuHs
miGna59gXDeESFkjQva6eTxxhBxgZpxqz/P9YaGhuY8n5W1jvvazVOOIlV3EnZfy
yuzgTnP8r5PNmgkWu+j8aOTOe/HYeSAdJAFLeWr8g78lqLkLcN56ZsRh0tCjDmaP
HZe/MQlEutpKXV7p1paosnjzMX4WWKZxuVqvvgxm4c+QMIPiXOFUbRbEJy0k6JVy
Gj3VBtpU+qPGFEf/JqQvPrSOVYQ8TWZ4CVkBNajAvkhblCdQLoerW++Hwd5DJKbg
Z5efn+eUDqfbG3p8EwMzENUGklqLV/122kDAJOWREYqQhJRAYFXxn2PO0tf0/u3b
LFN9AElXJPxChBOYfRxcwaox0fE3Z4x7s7o7gNI05qsvjp2/1mW+iGpXNKbEKRPT
atBP0W6AIAE4OKFWoIsDEF7g3lTtXCX007w4evfutt7gbw3iUMrPbrrbYne3vZ9+
dKu1XFN46OEn3B2xIiaQ96ypm3hkRHFuRFM82U8SE2XtKiwGznBE974KOH9nTjS9
Hfy2HajYO7BiuGwiGp4+tEiBf/RYJOSt7UsKgPbrajz0LfEtRsQ93qvRYSXKTj0C
RUF7niyFCdbilUWoqMKjLjfelivUTB4phqPDZbc0h9fICe1ffn0F6zR3FAhl1/f7
kE/f+GMZTX22MCdvFd2nfvn/GHbBelzzA5F1veLFq0DLAz9p6OAEKxMwhdwyhnks
3kLD35rzCfvaIHroP0BMCzW0nKHy5AtTT5SomCPeG0ew6lUou49UhUZMlFr5JiIW
0dlmaMCIFf1S41ZxJmweZLXlUHZQ/Zv57ThLuxQZSVybuwf0gM2B0rSsX/fVtDlO
W/JR1sJAXI2R+zrtsWDmumLGS9+6Rj6pkiR4VEQsDd6L6SD8OskMFutnQqVxFBqp
bCPj2fu7HRruVoqpcuhboJNl2kuPfV97Y8A2+JS6TuF8SGsxRvZaBox1zcI/WTZ5
7X86PIv45ZrguVPwoadfL99FtQ//mKOENboBk6QF/1vZkW6pV4waeuotdvmkTjqt
odeCQkv+P0sWTSaj+9ZRUtYdO+iU6RMXClBGT1hX31iOtjwFro3BeP6qbleziEl5
VinnfFKM17Dfvp0OOfIObf8BiDOq0++PRFcqP3YNRmdGgtGRpMzhVyCvXm/L+gW5
GWohcwxUoWdx5oZ5J+pOjGdckQGSy3LYN5/TbCk8KG4ixcKi1UX4OwyW13RbGZf2
RMN2sgkPqWrbXJAxA1pRRtt6hjBnXBROiLzZUJ5G6ig8/yzHga/Zcm3BKHqxaKDv
YZm0Qo88RhgUxBZWN9TpROmqgK61hnTZaZ481ZV4HsnF8tlvChzy1XELsDk5Zj/N
Lgs+IsUcuMKoTeGB5XCvxhQX1puwEgUduznUidczBeh8+CgH9noS0vNnePkA/lGN
m4n5Z4/A5S/9ypBhSRgdcsyaWep6Dy9KaK7nPGkccYKpEMr9vFeVw4EozD/nT/kS
os5fKjRxII/k6B7TBDY2731ekK9ecaUgqRh7JdI6EMDex1ie+EXncVBm0ofPSzNz
0wpN8kWs2sQb2E98upSnj75b6L2O7hDFan3S8dyeVyimkV4LE54gEBZ6e8rdYJnF
14WFPifNvyAjg/WGpPdAmsVO1+SJYqD8X+1jK9LP00FRmc+PSseJ7z9icedcbGqQ
7HRMBhOljm5MBDgQK1bOZcbLp5n64uw+JbbUVnVig0vjJwTuc77zUuNOArwouaCk
V2Un0YIOWath5qAVuY2TcSdrOkIS1cflEhRMwHHsSSZ7v//FuuT6KhlYYA+vMn2z
6TOgROEWjueipZ/ihqXH2SHbaFrm0lViiwa/7JwTRb6Lq0vr5QSHFG9o8JJGyugA
M/JOT473/Z/u+8DH7T9HbWcPF695vOY2ZsivN6Cftxis8d4sFxGBAGkxNQE74opz
eC3y3DQRIli7Nb5Ns96NAfQ0G4KXpj1UpnYTFcFmbiVJJWk7isLedDDQ9RY9qCYz
MJi0TTdgAAMDjBBlUtLHFUM+dURgxSH52LLpwcPD9FmZpawxNWE9Zaw5WTb6fTl+
tHFVvVIuXuJaF1o6aF622zlxbrNFk2oTdzL6dC/kNUauuH8lmtryw6cC4bZGu4g4
NG0SfQUxFwtfK7FNLSeAUfRNwtuGjPaVKGRZBq0bRrXWH0nocVdNUdYtWuYRh29o
VJnuqxwlzpup2I0sTjoab+Er/EBwyzOMpSARmUzdJSHy719J1pVtzkf4K7xTSu7a
xefq3YMR5UJIztqN+CIt7r1VEAK74F48gZPgSCpnpb8+tQF/g736H+V2OY7oLBbx
NOFUx9VFkoYhWQ/HZXsRRZ3QOv+M0HdCfC98634MzK7Q0+kSjyidZjZbzOg5GQy8
jg8JdfCNVODYeoYjTFZkxnbmXJs540UqnWkLCSNYAzQQqE8YJsAXdD/8xN0HopFW
7Gv/MXGzmZIVPLVuuQG88FKhwhb/blCumgr0MIeI6Ub5tOshUY7c1PkKYPoRD4OM
qiqyQgGdtakcfFVE4Kf0R5t1aHV3bEVC986mbnJLTLgNDZID0rWHYpX0bWSZYcSu
cgHeeeKQ3G6CD0z68HBzq0+MO1+9/7oFUOYQ2rlVQFQS6CVooTRJM+wgaWhgqzcw
aNd5Y6cK6GnGAYHCHpLA8PQ3In2kWZW4Ld3cAgEa5gn2t5bU3dh7vbAeLUSDPtGb
Bd68aWMAJ7C8fd0OujZhjdGaVKWoT3QuP1ghwEWwHzdLxt+Tc8bm4eqWNGGYgQ3/
R+Xl2yWLrCSM2hZrZNU36yhlxPPnlB7Vv9OG5C7jECk2/Zbjcn9vMo61pxlHEEgG
K/zbVlM92CF3z941DAkuEBgidn7O9nN19hxMTyg+jv5kvjWwHaNwigNB0YfoXp8d
PDpDytDBo+G5WLSghY2LjfTn7Bz4R00ivI959HbOU3sodyb8qQstI+39nqW4J7mH
/v6y0bacPA+zTBav6lyxbQe/6Vxux1uYlT6xnP5+YEWeFUeH/bQZaPuuee4zHEza
QGUboXkJWwkRj1gobfirBlYRPDHV/Vp7ZjhLBtGcNi7dhV0imH8/SlknBUvOkEbu
WK4SKWRjIj48/WTbcTTTdac2U1bfFM+TeCFNDLMyM+c5qrnjG7Z6JJvy8/kQ12DI
UFmJyunJ+lEtYgSgfiB1m2Gdm0SqIf7Ld0JTxEGV7Um32LFPWH1JOvFepNUgOP06
zWMH20lTrZyGY//iNTwKZPEQl7I+FmNxxg2bkwL9rNphlXdBCOh2/0uj3zlRUMUn
wBNkAiviXwSdpnAqQhVTHBabkDMupJSzBeQJMR/g0/2yuQ5DNSNm3iVWGmgUkXg2
MQIsM3JvcIFjMnodRfmpb2sjTmYvyNqUkS8Jsvxk6LyysrmT/ybpQqK5cWnz8wtU
TotUnx8LQ8ZDrJIYYn/ahN0Pe6oAi4gbHBJp7zcc8rnaDL1Vb2k/ytyoMJDG9aS2
syHAdkDmOpXSqjy+PsLDpPG9Oxe7lI54Bbuh763dz8toMn+ywcwABV3TPyJ47z1a
8BOVGb+7EJPZwn2kQk+XFIwmSYvkh4jDcyjQ7ukU8ilsD5P5N30vOVSfoWKJsSEk
/OQaeQb+uPYt1rXi/AaqDSe1o+oCwMntSKvEY9gsQacOSq25Wr41TUx+KwvnLxYQ
UmweYIGe7zznfVdtC3PdXv8yazDmjMez7YcDOgBrViLZxInXtPY5Wu5gWaehgbzd
KkmB68M3I0UAGvIF6XsDYfCYIahu7/+qxAC80HLIXefnPKyP1AD68lhwIdO8aKyX
MWjsHB/yP1BgUzNNhuS/0DRRQWCwhAfBKuU/bzCHwF0jCmNvtMDCzoZx/QfuDhXf
jfC8kXZLcxXWF5+2Dxa7KsW2xGQNIg7qKaad0GOk9yybczVo3Fq4LQqN8B1L5HhO
mir977U2ztqJbFLEG8NUBQLlP5JoqY99nx/tkDUXJioY3ALOrv3kIJqq+kIbHD5D
YVtK667IGPmb68O/wDmkLNiVeSfeQ0Appsux9nuftRUzQNjif68qhDqTiLtvqedB
A/VzL2d6Rnss8H4zkJEifogemwsvrSwMM87gLh2YCUkywcsIf1HAT9s/3k/CtOYZ
8y1oxjCTBaCW3juYq4GrGcjYKA8/3FaCxzKAgj9NqXhW3jXtkGI0nU5PhcZIJYd1
5IcMM2IkbxxcoRCP3wCmnTrxXS49iJ3Mw+uy2NfAosAEMnC0QoEKizyby+cIJgpE
dx6FYsXOru1polpY9oAQKrCsU3ffRdwyyHOeBJNJ/V76P//U3WEpdz8MZL9ml6U6
sPw/CV13QqZ/5dx/v+fEaZT3aZD3w//3e2pLGJ7ixajuVd5+VXdocTRJXsgtszsi
aHuFEX1ZRh+nFYM6B9VdeGS+1xGD2F8XI6oco2cHocWFaBL3Q5YmXbpbZcWZqyPc
SX2716R04Dx5dwQp4UdnnFJGcvToKwY0x9R062b1urzKmkWbBjkw5yHjVGf53vrs
QLUTOMw+Z6Ls5H2A8+5ZY3/n0K8ea3lH6t7qiFXvymVCWxPF770HImWXmgsDjmCJ
aE0rJZUkWkePlVKDngWkLQz4Low5BDOZAHcXoTzhnIJVTgSZ1jYuBIMtF12ZBgd/
hq1W6VnSFOzGSTarbQHmF0sga+rQSIibIG3JkHrKu0eHhkAbGJFT+i4f2YQvSG38
IbRwAh91KTP7WPxAXBRPU7eky1jmWNjQ++oimJ46i5bGl7FSmY8bWx220M4m9Flb
9z2BEOu4XiCtpmYNA0PZxGhTBFwjG/JLRAnMz2I/upKXLaMe1wgZtIWmfiilTsQZ
O5UZVPdVtcjvX32LGMrTlkgbGXSviylJpnU21iW9Gua2+4qJ7bnmR7yU9+H27eJ+
PDlqywdaM39cJAjxCDSCH0T3bfnaP2HZLNmPF/YC2nY3fpsHkFr6FoDO4F/6YfVc
wV6ug1k/YGa19Bue810k3yG5iqI/8Q1HzCX+Y0lcIt08GLfRA62/zsMv3LpWRaxm
nAS1W02MzR0ydmZKUYeUFZ3ix78srDh2eiMzvYwLo5k1Qf27+ynDR1wE8OKR62DM
XwPO2+/koYDnMmWeH0lAmNM1V/yFMOh7/IYfjCiCqSoXHBfvmb17sHKqGoeFYkH/
iIkUphStKVHlxN00TVtNB3ycX3HHoqjGBdEbAol1Jx0Gg7ywiM900BOEadX6pU9m
uO6hA2ZDRpvnBt9moidC1pwexv34m98L0/JIKX4mxRccik9+7xqOQC23RZNTbZ14
aVIYPpMtRHjYsElY/UnHorvqBF+GAKD0aWq8U/ImF4jF6Jq0a/X9Sv/dtfZsZv/i
h5snjmgkrRCpOe2Vi4uEanu5WRbh+vIh8GVismFoBmyX3tSOJE8WV5NWldeS9xIj
RFfJUbXahHth4KFp3mg8eJseu3ElXr21yWV6R5+01eJYt/RYPlttwDwcTeaH3NR4
hx2fltkQUOvqf+inKP/U9Ua/0Mpwjy/rad3f93IZARtanb9l5Jm3BvuaMN2K9AjN
iotLzyfUcBFh2OwQeV8KkZuVBi8eaL+TbupiV4mOUHhmjOmYAmBBjuy52/5IwJbY
PbTXaotuZmAwMUUrabC8ckYPX/nNUO3c3ZgbMAv3CA86NkUXbYINEMVMPo6DpYHO
dCoh+o82sc+xtLBxQ/OIc2CR7SPdVBOMB5qiOyafV40+MBcF5QJn0GgXfuMAZdWt
Dws+C80Y0i9O0tkHWQubdnukCtECGiyxok0s+xhuPDX8SnEgxxgGFIc45/qYmpQd
cmzCmxqK35AOnSoa+NnkE95zgWlurGvLXFzWiUoKgpJ8wkXY5okKu3Zc5diBjlY2
bZdNRLte+bGjPzIS97yngvBT3ZDSYvoh2yTbBbfMqvSr4k7+Io0QcG1KakuYU9k1
BQw5tNLgOIav7o85JtVBXOtw9YxCk9QzCIafHZRBR6Cm9Vja4WdTHGOpKOyXGXTy
phqVoddIXA9+VQsdwV1wtvXyE4jyBzH4aJK0i/jsoKDvI2/CK6i2eUEzF2i0aoIa
doltJ2AFP/LdczfTuV0l2zgSTx6ZXTbGXc03Epm2nWiLj6Qx13GySGyRM+L/LTUz
CYp29xuhSbUAEmUfl1yUHpVXgCtOkm3zr0kowjDuABwq4JlcrfHwlR6giKLLQsFf
m4/YU79/VyCflbyHLpr2oRhvRGgCL3na8V822yHYHVkPlqTmB2SfwMQY+nUnwrI2
rZF6ClJg1xdYr/jthdr5M2O6fI7Okw5cPuwQbcTVXt4D6YC5lIMaJYgC6/Sx9ZFx
yGnk59gcBJfGWf8vr+talyLrzz7cpUrYjnCN0KgKd+zc/J7Oc0GQrSEQpMU7S9Sl
TBvkfxgrJ4qaXbqYf+U03Bk7XnESv3n0bg2JuPtx6ZFOnVFCSmVs69uIgpa7TOSG
9/KCdSEhc/dZHZxO+a9UXN1BRvbVStB7hjR1zIL6FHSmUYQXEM+mG59tEnIzrFPY
y+9tT7cKldqLZaBYg6MujfQ9j/EvCNWaRcGfFPs5TLHsgb/eHSIzXfPACBM9Y/CV
3P5uXbRDxrn3DBp7lWRR/3BWopfCNvGCnwGBZlxjTbZGrr5Nrrxps2I0yAt2Eozt
jOucGBcB/vaAR8axv2xAFAIBIucN5mnmdYaLDvyJC/5izfCKCHqY0Z+avXQDtlt3
mZQq1DJ6xiE4hR2ieEIUaP87TEVQLALdu1zJbYgnnthlfVt7EdhaMEvxkMwXZc16
X9f8HzfBRrKZOyNkBNIXt3CGtg+gS6/8e55SZGZ3AkDBQN1XW71Oou1kohzZkhUN
kdvSo+ZCPY6Mc5rLpAydyghEXsPRWP9egpcunKsKEtLK9fkqbTmNXUIUCZcqDZJP
uP47aLVISk7rBN11cv1wt44vWFtrCv+qCgxDrlxRCDNh/ahPKIh3mDOYeDXWmZ3z
GGJ/EJY+P1h944fo6scCaBPpxirO8zYApwOg+ir9qjwfSbL9pFufcoUoANeav/cl
HUZJ1DZCXQyZDmk10YHw9g3dSEA+VfGbEVeDVLDNFByqqHWGiDK72+XJUOiQa06Q
4+4vLXN2/MKAh02AwlTz0F0QVyP+7fcWDGwjycT30U7b4twg8PRFE3uA2XkRO0dU
J6sodOf2hpq5W04k6AxqreylL+7jCnxH0k83dLbzkRAzaMYNVPyf/DmE856x1Lv5
e/16I7C6DD3v4FfbTzOxRzJO8YMdAW9maLzLxIxT3IpkwmUb3040wPQbNfYP3dwr
eR/BE+BV3HGrQjAh5ynVSxV/d0nLX2Bks8hCf59O/FKaZUgUVvPDljmPxCo45pG9
tz4hXYM7EI0RselDBlZlfoTl7H0ACNpJKPZ2aiNNn7n6kpTGvMesk6LSqZ5TOb+q
Y1ODBx5uRWOfP9etvhyBIHDesHvnhqWATf0vVCVH7aQz9Zt8j2dm9bZe3AGl/0w+
YwG1EZ+qTGrNmh3MXCyISq1WJTndNSU6xq86+EnvHLk58bUzKWJ2+gP9fXeFF5QP
5Z55uH1wYap5OeAZ7BXHodFF+cDDccFFTN8UG2OmmmzwOMo2YnHZAJusb2bT5odR
kfr8UgLv0PwtNSR64RhpIVLpJiKexGMYfyfUXS6XeG3mE69xksU455gjlx1rPSc/
Nb03GqU5y3DN1arsxvq4p0B/YOgr1kKMFQOMklzfIqU6OjEJ3cPfPfbc8+L7kcy3
LLSQBiSl8mMoWF1hi755+h9/Zhl9/J5t5qhs+/+/oAdBgiDle2B18YKRzR4P5e6r
dP+8RLxyCPnUT8/EKHMlt17DnwAGPOKZMFiS7WbJpt3ONTjs0Ilm5rd5bxXzNeMj
zRsOGsqQhePQ8InNNHs9V8zdpEigpytQPQs8Lrz0/O266cLCd8WfQ+LTvBWHeKGK
X4e1S3LOnz6a3F6MLXMoeG2Yfxn8/5Lu8Val2qWbBs3UUiLGJqE9GXgwOL+qTQ8/
QpGWgnzjU7GegGMnNvZtR8IZ6eU9zPp7izlS4HuouCQ1myY73j9ei9fjSaZfJtDK
4ap2YAC+Tjn53QdfOG2PZROUv96Y5nWfmQKHD7jBQ2mqsNwyyeowpVcCnog9XkXA
WOEIHKCC+SEQFIo807DC6s1qRu57ISPc0tC/pnm5s9ajILsnX0f9dNUE1UFqQs4b
UtsTNkePPVj2ARUmjrpRRcw74c0FIfgGtZ38y/1LUU0xIMoAvUBabpObl2AH4U5p
043pgnb7br7Q4AmIUyLZYU5Ue6OnDMgYMdsEZDo5rWs6++LbqFpxipKX/Up/MMSJ
4Tht7H9NCHzWEjD7xol0o+iK2B9I4HXaC0ygLOssJyAdfKyl+2CBfTD3aDv3xmPi
vbvxe2Ux+hPqqXr4y2uxrNNIQdk6PrgTBThByVCKwd+gUXfdosJcSRLhBib0JSos
UL10/bq143VVMQHuJrzG/6lwBn0c7LhujhAdZ0qxrjYxeqL9Djdvz4T50XvAXvjD
UsxnKlPN6KzOo5vAOzNrmbRnYfmeNC89Ag/kjYeYqPUfmmVRsDXdCUkIX+ts5141
6lq0Z7RdGchGt74V3+kSpoQf7eFjR4ZD6mbI9gQSAUz0tEaVYWP2gvoQocaodQoN
Gvk0HsG9ncHzazs2bU/664q6bJXjXukh2PgM2JYOEE0gsYKYt8hEIEetyK4x8CAy
SgwJa3fRimbJr5FftyqBEwfaKc8ShBwd3qMUV2fXIFTghW5t3ks6j4FzMctcBQpm
LC9Ngz2NqxnT6MphyR6DOqZ/ySomI73zIV7BDFQxUkuyFsLrXY95so3dZBwYfjMC
R47ljA+vf4+pghUIWSWnFUFEJqGWebJBc2aC+Svh6S2tBHgudmRL79BwaA2lbEX6
64nzLMM1hb6UVOG2aa9Fd+tkhGtm0R/QDIo8yPiWg9c1I5Hm3bUcgOXEWF7EkHBC
byfpLhhTYq8ghW0ZB94Esl7n3nHY5DU3D3rv6whb22a5vRPGtDrzpec4dm8YrWlb
bYEaMCn/6xgeQkPwsIg2purPAwvZ7klrXKbzvi6x8sRYlw2aP0DUE31EQNfizGaE
8eO+h+p85OKdWuYLP3kQVQSJlDnDO4Z0O07+xBknPMkh5J2TezEEsE+P2RbS5Wbf
qhnK/QR4dPiG38vokYwbBZlHIdlqTM+bSw1QSSFF3FUtTMeLJwOyO0Hx9Q/hWr/N
gCO+HmVhCXF1KG2h2aS4Vh7rR83zAaPxAV7keOdwYhwr23k4epfuUErBhHyk+gDV
5+yvT9SBqmaA6bdyjuipL2SAzLs9EoT+0pRYkocgEIbN+HsJlMs3emh66tmVY9GI
XCZs8eMgCKKWA2lbEMYQhJhzama9giqQ0Z+nTA/VV5Iu25+F5pFNtaz4iRuXz3yo
BZcdtubo72MOaiM4ixFMWURJ/kHB7GsuS127VmAAtNmGzlIcfrDwYrDlS1iFLJhY
MNN48HpNX9hRwFTUI/NwZIfNftIqE+0Glc/leEyrhM2hjRPNEVuo9SH9e4NbPCzh
nimMTUiTfpV+RP4jOJcpmR3zvpXcTjS8LkoHbOsC87i/TDb7yxqb/D+7nnR12NET
b2KIItEOf+p4zHj8OgIT3XtYV2Ci9Uoc6OmIj8Oy2iMka7hQO2u4JXwvgTJ4guOB
gMpCMhXALPx6wInjMjaLFbBo2mwiI47MUbXOEJyuY8KfTBuJ+sAw+T/zo8R/3LaE
2kAzI8LUSayiUVgcNX9sZZkSnIv+q/zpclW7jYV+gxOOti2k1yTsVjI+ixWmAKrs
xtxriFJZu9DgiRT8gaJe5Zd/tnlnV23SqJIRlyRNzGfQojvjNdZIgFaSTzfZRFNi
ZOn2X+XyfygQsb52WCtwGYS4JMR/ZG/fYpRVsykVcPYUH3aFVYSx4eSy4PqtLino
dhAMAOjBdwyqK0kXsbKk6hxRCpm7Yp1DLHXMtagEMs9ewdW59vtSXWHkgoGWtBnK
sa/tzLCOQ/E058UBBDOh+6TpJsYhxqrXaNZsqUJNjlOHkQEdUR3vZjjbu/JJbNZE
S2to0wFHDRKjdX3xwI1Y0yYnRtyc9F54Hh/PmF3iLZ+20UcrrrQucdywMGh/CseY
HHpINxgKkVxrDhfOEvvRmiNCxVb9/aC68cIbQLiJS3tf+BF40rExwIk2ZNW8lYAt
FklRZQtdEKz2HUpGWUym0FWKmz6wdJdPDZ6UKhxaFC8Km0XEChO8PJyXp1hZxISl
LL7yYhIyZLHevK6JsU/zTuZ6XCaCNXmW2wGgpIfULIygCSuRW2k2TbKYyhzwy5Kt
adwHTHUk6d8MgU0IKp0wZitHXCdCwuz9BImZJcAmEs67bWt8BcLrN/j2v4eN6g3U
jMgf7gPokJ1jG/aulRN1+HQ2yNKmLX3iIXtXkoYRH073zgRycMunMvuQBhHVz2nQ
CAqZj5uFM/pxwSoo6NQZVbQMjdcZQv/FG/aoIyvPG8sIiPdgX9j/TXoysUeWeskT
tTho+0Sp/DuwgAhU5mD9EhoTfSvIxj5p27Q6E876xwG7T4YNWP90VPHpq0vBxiUp
GkUvG7RX6w1yhlvf3CiilmYjINdNy/uDLIKgX8FPGsz7yivgX/1UCePH3k1J1daZ
qYL82LjvTQH5DsoRhQXez3c4zD2BApx+2t9Vr8NhhCo0FsHbW7tLBl1nbFROZ6sk
2YMjLEOpfLV83VpBXYAgScSZ43XobodlWGsFfmK99tb9J1fwC3+369jPI3tCu7ty
gx5R+P8VFNsb91Mawda8n//ouY8DUS6BUCQJVCn/oDO2zcmiFaybsUyhfPnbV9H1
z6aMEhWE9EwSC+qkwVAcfhgUths21k7JD2h4eN8g+ED3S1lKlyQn8krOzNS4InBo
72Lt8XJ+REejb4caWLTE0uj/xoF6YJNNU9xIqzm2ji3coZwTq/9FCpZcfj+iNN99
3xbU8YG/+a4fiqQZl/DNqzgOaffzsF0LXW7v5jk1jo3M3S5unBccxhTDZ3Ih8M1z
DZvr18qCy38ZtscrtXmG5Rn1i0QH9aNsMykoNw9EwCXWWjdim0YCOF3hfMCYaJzB
OACrieUMXCXPaODFrwYP+b9yVanu6TPPF+L+MureHF+hnGYpcJCjA9JOgWGNLLp1
eIcRaa2+bf0EA0sCsVlZG2P/5ZvvxomLTOhCeK2LINPU/ibb6cU/kGF0NLT6dVzv
NJYVS6pu21bo7Xa0VMym1MTNT3vGuSoPYRvObP/jy9+ZOIRdVRePjQTEUibzv5V9
k1f4oE97MKrm/ASIFL1q8ugGrQ21yLCrxlmcejyBAv/q8RfCJBq9CMmmtX+pgb0C
D6MW7HnXA/g/9DtqjeFSXLpwDmxAI/RVp3g0hmAO1+A95CUc9DnB7PKGwOJBQ3LI
N8jSFhfyy09AD6LzErpQBrwOmTGzhlXG6F/bY045VSq/svb44CQU0oHY6gBA/5mm
0XA8F+vlMvBGhooHza7ZXEwF+Z9cBol9XqYrBKmvgHZmauyMSSVdN415XvDjtCCs
TQCzBP0iwt9PxZUroXxFNtO8S8ZL1T9HiV83SS1juNDmsBAasSUJ0EiLyd7Em7ub
jpvQaoqo/K8GyLYzmXTp60oQh1JPlcl1UkzrHRAXCFNHoF2xhK0ig2niYNPhMgie
+LLtnRaERnn2eSBUCSJxZMhSUwcgwFbwd/GQoaSJioXZ2xtadVe+6dS8XdJeGHhM
pdQ/ZU3D46w7N24IhQck8fIK2cq28oo8sSOIht30Tmv1CaFyY74o4dS48AEdTNpf
3tlc/SRUP/4valZpreuuIGYxy6Pmy+xbWNlW3YIdaLkA9q0lH+Tu8XKgof1qFiec
Dv5RcAJV5yNtMsUj5eQzHbzf/+I9HOaabHSfx9A3auhXCqgTSdIbLl+Ne8934PCQ
LIOffpEWLB8LY3ILGp0DKYnzkk5sfMLLnNE3SYBBfdwdqhSBkERmf/LH0/r8/Z2O
X7FcCMJlGK9+Stxhhp1IpglYHb3bWpR6iIkVhYHZ6c5T2e06n7jk040zwKVEnUMg
7z8Kpo8Vf0Tbg/2ILsMcEnO1EwgnRUZS5hcwLgJ0J96FI/i6OMxNaFp46YLx5OZR
xnjM0McNqPQcIBpCWAgvwNGIuTa+UpFcdOfGfwxULZh3IUWaB6YRVy0BlpTotXNN
ZZzmoDNkGzaln36oUT8XpVC25z4dsJl38VmNpp4qVzZkG/Hk3bLKT2RFCwGwAmJK
hX5zPlF5RzmOGYCiE9fP4ngRpc5vvRBDt1bdx4MRQYRX18AtDHDOA+WEHED2GK47
APPz8jtpbk5N2y+X8dEhWR5Y1oRz7EqXs2h79nEbE2fwj1sMb+Tk2/zzcPwrKBW0
OPh2RnXeiZlY5ZET35Witjbv/PjphJLJ46fhAMtOdCgHBsVJ1qOrXQuf/wCkLx3H
6sm7Qn7Vk6fS5HPrx+7+mvH8D8Mh7JXZSwjbOBokRakUOzFhAeJsSfvk9ERR6qs0
qUqMiZtOfGAJrEp95HUuJfYJgFSirP+DhLY9/4Dc8z0Y2l+ACvI9V4iUq3rFOUIx
QkPqG+bzMzr59fpFAyzcr1lzp2LcL2+yjebTUgIs/fklee6y72o8CnbD++pyVePB
t7wiiuolcbb9qNiW6wqNj/TMzm0+bTwewGU3Im3yISaoe42ppDr1erg/bnVKOKHu
iEs+C3u395od9ZoHC3zYSfBSg4tMx4gMd8XMyP222gKdNpYV1Of93+O3tyjEvMI/
AaJiOcrrA2CqZH0yYmHg3Op91HGVbbeWEqNm9VVI64BhRFb90EdxBX95F6dNegSb
W5azvxCbtQDUd6tkLLg443H0n9ua1EMikuHFu3RMztF3MB8VHyyKz9etFzQKVhAj
Tp98UgMdofQSsbKY6t6jzJx+qDgBLdiw3AgkbcvmiySavBxDyZ+zIf7bFdb/zsgR
k225UEE3yWaUAdW/TPkt149BPFu2/8skBCK2JhlU8JCLTOG1nktdpKuRLV7PteiS
zG5OqgfaJnKpt3DQu53k98iPkgziCxj2xvn+j3wr7p8foECCaO8dHdQuCFrS/PvB
DDdX8Xwg0WDX8SaSW0aWXsttDfwbT4YZMA6tIr2zmwT0D1wBwX5pIzjMkuULWBMX
sh42vOgrBYrVJHvBnrgXwBc3qy3vj9jHqD2WSgT2QjCOoXtSiGX/zY9N17RqJYAQ
5iOFMY4LBxo5uI+VfmbOKBV9fxjAscBSq9YBRGX7JKRSvQyfRZmZBSf1drvaiJ51
oyGC1YXZamTGa19lVGoeiE/krQeuNsUFuhn3hOEek8HX7UvyqrMimcbcDDNrEXVD
Gqie6a+OU/HO/30HD5E7RG25rJDLtk8j71Agss+Kd9WY2UHcCuoFBKpGCuT96jan
g3f6msoDlEnMMkpFFzL7nk3Q+3Td3XkodGXgYikhNgaAgU6o0D6outkzLTbZi4bz
4RPtwV9gF/vlkS5t5joJ/1W4e/7zz7rWj3k76yxySo/tzec/sUsGWkNfYsXU9F1k
o/2s6TYBEAiT87UHMmxhHECZemHbMY/+e5Au2VWDTD39QqBF7446gYrXImwb+aDj
n4barch8SrRg6t6d7092JddURdC0lKfJgJtcXC1jAeEwP9c4/TK1TCi68josPnFZ
EY2Lvnqj6Y0FM4rPyARNIxUATgP+Y2RCcsQ+iUj/kKA1JR0ADgh3+QHf7rbJff3z
ZYYfQfkS+c8BiyCP1mpI7osZqnDUIOf1p/NM56sl1dNfb/+hEP4ZhrNQRVDUAzOG
YnXciLX+KzZe5+uwNo2M2C5enFvjYEEZCY9VUhg2tEQa2oKOoGyGcQMA0zHpUGOk
mrmMaMhEoCiSR8ZePNwwXeZqpNzCGp/CoLJzu7tYOIBmqOeKTydmnnkqR845cURU
aX3o7zRqMU/rteoy+yrTZ8DDPwDwOyTdStPfy2QBVP/3Lp/7qR/l6DmzI9noXcGp
6AcL8jSDyRtD8/l7+pg15wJsTPOEKJ8fHHbkoyac5YyAM2UFKIgorxjr1X/NFlrl
2d0eZhLTKHPBPe1d55rq/2vfa6Ld5wx0UIb5hwE4pozpohfh5s5NMMgOtHhcw0w6
9cfptmukNMdq8qN0Eb/5uJ9DwNL5sXynlUjbgHMMJVb88UIOLQtoV1mejlrRc97q
0Rd9w3o2hXMyt4f22NGUd1t7O6+p5ZW5WROiyhjnxTbZKJcmI4GkJ5qgYXx3vcCT
vQuxlawa4L5agZs/96rgi44DhD+Y1jwGB6klh1cjWXy/5NK+K7GN+llfwm/3Cbf1
4Tkquyni2d+wu7ZdxqyNavoHA2D5qc8QqaT0EFg7B5VLZSbWngbvkiikcA0eBerU
s0W5iDJiPiZrf3z48i6/kno5vUatRDvRUPeYGTcp6HP0+UbgF7NUiE3aZGO0Ey6G
u6WAnMxhBRGe321X7xggdDhIZLk2PESZC/MzVetlgzGqW2ACg2YUmKRI9YPUvS+E
EC18OB1m9COJYXjuCJVX4CKbR9a+wgflmfw1pFM1gf6q7/0CBdC0RzhOjnD2k709
Pjle7dt6vHcCoxkiV0oQ74cRgyBbY5ouOQX9xOfOMTQlcA1O83gZaZMip4T2Pe3c
GSvhT2dh2o9Zx9FD4N1OIozBWs0tc69e4kERFDk9K4c+b7FD9JjqeT0O9VQEYHP3
GxcUPPtDGXpXxQTce/z0eHLzxhYjJIoNfi3kM/S/wOHlITKlAw4eCxyJx/DOWZV1
Q3PfwYtB+J/rBBBgps31n6moO8vY8Z58JMUHRKgaeNPQCKiym+8vdajU/MZMq7Oa
63shNft53DxMBo1nNhNaMqXT1NMdkYgd8Ak9IMHg+leBgRzdIJM5H9NeFzvJGm1c
N93n0phE+Hj1mbMPjCOxbqB79QxoKfUjAamXoMpkkuCdic1QIgcZil9LR4NHLrmd
WwmFn7BJ1uqM+8puTozgSBVglmD+mvaraMVtkl8Y1/AItmAem5S6fnTlLKU0U1e7
jMxmqMaM3QalFlpz1TGrRxg9nBdjI8ptH8UQGCqZoN3caOyn7F1vH3JMIDt7q9jb
xL0oY2oCVhyHJqALNpXeLFpAl6ZixNYYSRNU8fIbptAin/e3hgilAC7Jj8bxoz3n
3M9JdnRiMNPC2iVDFEK/ki2Y80ERnQhekx0l8HDWjGQ5wtQwIIO5ck7IH4h17ubY
5mPBhEEyGWE7i7qL/Hky55T5/+Qe/eSRCns4QhkC+gpmKsBkIHpyzeVT7lDAqEsq
pw6I80ai2VWjxC2xdjO7VOE4D4OAqQMqDfRgR9IeoE53mB2+2EaFiXvbBdyKGOxE
IDW4/xUy0ji0noPFgzwIt06wDLgROeXfluBCYh3rLGjVGsEOSkdZtzlIN4plnYIr
Dw52rdNtvRa8oy3cWUSkUQtse1C7z7xyyu01gzxxj9TyZxkhv+QyGffxVOtlGZR2
WEeUDZZI+5PfiN+QHb3hWObns1HkS7mGeqDlAVqTNeHKNRf+yIGSh0WYtKYEvCJ3
JXnGuW3f6kqbsBOZfHS3oZf1GBdv25h0LpSagnbaNBfyUTQ7gVOZTZRmVvVI5uLF
MbhimNzxbjzYEsyGYmW7RJha7ZC2gJnqOBnCVaVcZoFXeo+nU8R1a2KV5SO7XLZx
ArrVbu/0lVkm52jTyC+N3ds87H9YB0EVQCP344kOJuTDip6yaZYs+Ww8RfxjYBPg
H5Ry2Uev+biY157ojok/H3iPxn792Q9DHlgKk1ZJzU8CA6wui1Doym+8IeLPXuPN
EMgAyZFeswDfZQAtdjd2OyQUb/oYInPBpwWTI1bWDROvEVs5By4pjfkRjv6VHrib
LgLH6IoXBI2Bvg33tyl+OHynnxXz4WRiLvrurYLeNjz9ynQCRs2LGS6ZhNkQwsjd
CscMeuQln8wYKXRCJ/zfm0blisEOvh17VEXTWU2qd3XR3J3QcV2sAXaAXZbPdd0D
W9K3RuS43wbCytZWH31SPg7DmLEbz4qwngvsdOMoMN2sh+j61rUTKyJTvFEaHxih
1gmTQcI3sLlYJSDP+N8U25Ty1PXC3zqqqDWZ3J9+az4gAfzwghBWQrxLaybNZmHO
1u6LbRwENt6yFk+yENP9PwXZcX6SYSL9E8DGGDb5TUBlq7GskLjCUY36ozPnoKTL
/abc+8FM9qGNETTW6NwormZQk629oxjDHtCNU0CYpMLGl9ltd3LU2gEY/kbMYPp8
1IGyCguW+jN+SmCEWFgXbCI77xxH+y+6Rb8qUzez/jOkTt4fAvJ8WfbZk0/AdgN8
acOA1GBl4yB9j6xn524ouKGsLQ/F/+144LONQIix7YjIdJY2UGFXE/22D5EdOBzw
mdgnXIlH79ApOvJbSPsIdhj6bNn1NVwKMl4tD8d6It12ozgXI0gyE4kG4Hb/0V3U
23ZCF+9kXB4S+qERGYnFxv4CYx2F/SB9GfkiAHlwyvFZAcUjGD7ApK2dQdRokw2X
VlvNMnQbLqSAK13C7NFvAPyyPVVr+pgbuipev4Cv9LUlVnBP90gpQmU3AIq0RIIm
638ZnLAYryS1HW6K+oybLijq0TcNOGp3lwRv8hA8dTMY3GE1cegEw1hQBYaCjeFA
mTiRo53VRk48xnG+hcmWPv2IjnaVHd4Pc2KS1VLr/jdNkfm+H5AeVf2POIl754nr
wlBOQospfxeyx43DxDRFZnIsY4ugYf6CVkb4T5MelD32j7cnKqpYbnWJFir+33+P
xQzEyyqQ/6AjvXpk5ZnHjV8f55G9TLLsR/y9tDnisCUKBlsS373+Tj1RwXmnLr5J
nhLZMBaqHtYSla7LIttBaPn/1OfnhLbnE7a+RaHzwuhqI8jQCpbPlP6D3vgkFFYS
ArBrqHMhCElP35U39z5psX5fJuOWWZykPQoVndTg54NtXB+NVXb6lM0prKZTS5Uq
0nAaBAXU4xJ4q5/zSaxt5WGI9TaAZjucvl3VxP14gLrAUvwaQ75qa+JjqNSa/DAV
RvUoUu+tV3hW749ms8P3o7ojSFuPUSKt+wo4On80CtH71cVX5CqVCWMUuxFS99Rw
SfyA/Yi0c945cRKsFe/3QB4EPRCtmGQ9Ti3vF2iCP/SigWKIIXzMzmxz8TpMQNBA
b+ela/DDbjcYataQoaNG0CluoYDEnDUUGP8ecCAPQSI2FpPrkXUFS5zDdzakXXBs
WWcbfd1k/pFVUBM7PCIyU8S0bjfbwispgtzkoVv2vgEmPM46F6+z3DS3weYsjz9c
jS9hmX+jxhTnsnBPLJeRKlryInNMKf+cW0ho2odHZY5Qe375ERlRLzELgHOdErzD
x1S5p8RJEZ+MTxGrAG05aTNjezGiUKRsv0DnM8oTsyNu6qB9y/osNe52t64cvjdp
9iXAjjFq16xE9XksBzN3XgjSGhyM17LW37VpdIBbCozCEdVF0ipp6IqnDozyEBF2
n+nFOZ3lUfe0lh77yHa56QVQW1+/PgDyTF0BqGBr9d/oddruMAaHabalIDF+Tn+q
Wv4QteQQ7Vd14NYB0ghw1sZiWCr5rQRzqQ88Kf46gVYjVi6rbdYUqjJkKQfiMKgp
bZpohm8ud181gAh5kcBxkMEKu+zuqb3DWxIGDfOBdKBs4qbBnZuc+o1Y2i7//GbI
1MNvAs/URPloVXfm91gOqqdQ+CW7uQ0kF2G87AhPNE9U8+cHgjPs8RRbB+kI0gPz
2gRU1723DvXgKG21zuWp6eeawyQm+a7jqD1YenwDYfoyYKDXKiEzA3vTP2PdcjJr
nLBiHCrF+EfRg7mNgN4Ufb2H9n62+zJobXlFMJCVpUWbdka8dtSCedAYdJz5s6pB
4jEJDfwZ6dv/ON5qpnraaoFX4y1n/889FTTy2bfIfpRHFV96khR8dOqrXlTlbvQm
FOdRBVl+vJtpbwsLls3F30EJ89JKj7cUxnbKvu4GOttbRgH8GgK+LDqtLQ28SUmq
lFGXvIeRHaljqp+tmvflmiEC1nPj8N2aRU7JZ8+2G01qOFUowZr4GoYP6Akg1+ap
SEpSINltB4Q7p8pbndpFgikSJr2+bbmnotRNq72Y8JsEluBkTTCGQ6eOqwcpRkUp
1oyuGSBk1jJ9nJncVvYtbI+CtGDKjYnA0z1yBKJogNPidje0mQTL7BdlgI/GZ6P1
C7gZiVQ8KJjiTprfmAjnqO/Nz34tSLJ97F5C2vDRVeZdJLqjK2wHNTPkf9GMl5k0
ctxHZdNYiYPIonOX2oZIW+MllD7uSSp1QzOSIgqfNF7LDKj4GsgGmiBwIdQbMpyq
eLNoYeQvRgy8IcxIz9aC5dBVyIYfkBRHy1BFLpKWZV0RVy2Ao2HW3lJJXEh/ZOMo
oelHxIAh3Ih3GPlq4su5OzrRI2saq6Hm5ma8PbS6trPK6mfy5tfvSLS0uyQHmm+R
QUXopMBruQXraTlKqBCFihw7ye7M350Tn55UrpctjbuXdovI+U01UN8wOooCSgAf
q0HJ3ws5HKR7+sEPyfcZJ43pot5BYK6SSh2ExTpvnd0jgdG1xHyKz8AYlLxygkc6
3gRmMR8Ah13upRztRKhzIWUb1ncGSfin8II8tJmiCphfPRCYZXr8j/atuILTpIws
Ua5bptWBG/o4ZYAuIdKwX8GSJePNO/wy+WzhXGtD4DMOuN4kztC8tqya2/WCR9Ks
80WMdFgpCKUKReC7k3ggBxH/aIoobAYQubEFSlGMeQnmAG7hos6IkXzSf147kEHl
Q4glvyoqnl9xnvSvcsIXPszi+4I6sPl6jEOuLN+avOOK9ujTKiA4KhYHcUqOfOln
MRp435270Nna6Hdzkesh4p4JDj1MstdntLupmz5y9GzxPnqO4d8dit7zcwBko3ol
0KmvIgVtTlt7HLLjTNZLzQwiUDFWjotJ7yL0+oWc/25ScX9EVYR5HLj2pHiGoItj
fAKWfgvbtuSFXviRRUszxmtpVJAjWlz2YPqSVCNjP+3ztTzO6ZOuaj8lSJoAQk8I
1MIA3WIjgn8Cu2Zunou/MWsgg+IAMKWp/EgDeUZ29tz/TUSV7lQZ5Kby3wNtAT5P
Kj7mH7konG1ByTiHhawIjl60/pebrth3tShvOaH2gEr8jGG9vgPZPz45JOnGOkLc
K5UR4cp7Qt626Uht0QO1bBsBS+GfcDndIY/dYo7l+D6JIed9TeYFgRs7HaRpGtVO
14ELtM+NTU8NetYDjIBr7kAZfCxpEOJAzC3tDr7WoXYSaKNF42pb8wxfccvquhhH
6nspkPROQq2xu0VH/W2nFh0IU7s4Hilrm+yOYWwmREdokAKNnpYM3R+vkcmm/Uq3
/HIw+8BQ0//h55YUgvElZO9oPRYafgKh8MZ56O69fagkeLYBdXmX4mr1xTfS4X/T
X30TINyAq/wDWvzoarqmoLzeSkvJgTeV4zs++Bv4vTqdhc7kKDbuETZ1II3VfRRH
LeP30kejjZcWRDnQKY1QsQZQzVtmjRlvcdrxhom1cTbd8qrvvZP3t0Rvv4xgB2fY
33aeqeMrXGLB9CNX2nFC8XHEAMQZ3yKzDCpjZZA9sV120KIr10fmsYoLtO9NFFmY
HrwN8wrfE9yieNf5jQxCn7VUxKZQnDLAaur8iKbOpmEBPzpQxut1XT03CPcY7US9
47pEPsrQBdA0voP9LLPVH8We8IVBumiSq+RJQSKr/5I4wJmMOQ5FCa1bfDBehWQN
kmiWN+0UBfqammsXwrDeaFssMRoD/tiOtrn2mmWuStSOqEp1nJ6hMl0mPmKEEFLI
jz1VERhWYT5QCAnO5Od+LybUDQlqUjitDpb1MWIT0YlbJZVXptmnLpASTgh9kLbF
WSODgzZRbfcc59ve//8A8fWyeJGvtATsO+3G4IfEb9f6uztx26n3HhdxDb/vFcit
x0KEJ+aeQ01Wbt6oADN5ICbxdq+am66ZJjm/y09X882Gqq7NVciPfTTU79WJFR92
ymwMk1A20FvJT/VeCwNfV/mEuCdLLKVDTKiQHNueY32WR4u3vJUdZnouEKxIs0ZV
3kfrl7qMNPqwU5ENTwn4+Fp3ebj76rJS/hnLnhk96tUWCJC+MLvmjJiXhqOkOsXJ
UrD00JXxlx+niVffP9hHK9r/XlzRPHKGwSJ9DIjwJC6n8LjsACtFCWPpjThqzcSd
aSrK/WmvhncM+BqX3JpocCJ5dxq7ZSVDjYHKAsDTznB3GQcMvks5t0okre5miW8u
aEkmS+fdMQ2t1N7sHx9vbnaCruCLY+09gpk+Tz+DDtMq6NppYeLOlNiu67CXEs89
aSdfVmv0a8oKbShSVavP6Z79pEhYo4NzE9CKlPPCQTQl6EJZuv59YEbJBXWJJXRH
ThTT2Mp9823ts84xL3WkApg7GTARiKRmXTaXt27BuytvnpKbQ57jfARpEGga/OE8
N9nnowYb/hwfAD7isRDTov87VMT2/U1aap4jLEqXTbxSuzjpfTcMh5pJ6KTWtbPU
GSpMFUqOr/dQmSeKDgQeNo4HYQKNtD0oR3+kuAZfFTCL/gAGyZEnzTGpG7f1RBXm
TB684Z3BafRAMOPS5ROdEK4aBeYgzqmuHv4bXYZtZaN7Xijy2imGlcvzGt7YCvPv
fS4bXdtTjfVnz68p89SRpQ7KJzIG11s3dAeQM5qQzXw6bICLpaefOlUw9MQwgXhX
a+fW0ElY8Tft8OCA50KtbubRqpK4h0bBJwzpHYDY4S5eolKCsYag1eF0QH5QVPul
X2MlrbxVBOdyfc5zHtjcoq4JBCurmb6qcjIiEHNsqh0s/40a9asFVfePjaFRcGIV
WQ6U8C1eQTfBT8I9LkobNDhuSxTsCQmh0tN5lNkAddzMaRZ0FQ/W/3Wk5r0mGcue
vzIltjl5WqxbVGfrDKH5uOAp6Znhe7/uxD/mSmwNNZiY2PJ43XLCWlSHLPOFHLYD
ZenEymw1Z2KHA+HWUui8RqCdOca/NvhpS8S4rZyk5LxHxPLKbOCU0HuMNs02ZjMI
PrucBDRaXhOfJ6D1dTxfMBYwDVxgJOS06riVKtyC+8NdouMKowtmmAlsdh/JGlXQ
W92WZ3fnMIeHFFpE8MhY6H+Fve6/VG1edcN9RYLd4wTUqUgp1Lo5UjUb2fNXjyA5
IznTa65lrc72AcW69H5VkC/BcOyJGfDo+7icjQI3vWThuiBBnBwWGaQtM6Z37PBl
F32mwccNKZqTqL+y98Hzy5cwgAiAqWelPStNVPOR5s9DrlpzKsbxDQCthuFrfjKA
LzaWVKO21E1E11QfuS6RuU85D8Pi71sV2/7YqyMBuA5qGGAwScCRzKpEniPHi4d4
UkP5gaj4BzhCYoW1bz+N6jpTfdaxLJTXRSsJdobG/kM2ADXXgB1KjyubQhWto0g6
Wy5qOUI/EaR3B4F3BR9CiOFFNARQduqiqDmKtCpSmTvAneR9fZgAl+WO5D4NWrEm
GY+oYh6/oBU/+wJu5RMvpbI2Glb+ML4bgnZ1O5cK/hRKV18Z8axzIhhJWiaLxS3a
kQ/MR5mplvboZcLsAYn8dxS2dHZ+otC56K4c4n/Qj2/1BbDjUcOOViocmp/S2K27
b3i0N+5V+xD+JZYRpabZXoJ615G5ZLMMl6Ef7iSonIumCB75ksmNJH87fS0YD76J
X94p27Pd1bjzFkUT6Ar/jEr10yRQ0qh7LmeljtB95gJ7i04zXlUbGdbBNkyoGhPX
tB0S4IIfQ9SAd+i8xyzjFpGTbCMVH/yWz0nUVxcUT6k8sKyVhadCwXMD6IMGFtg/
O8ZUZVd9xrlMA7YGrb6NI6nmiwCpzKqLizSzTFL9suTMmLy0xIBbXZfufXpqAD3b
HKIH1r7qUsEPiySAMGzgxlWIhK7dFsmrIK3y0xdfFc1EDu+T/iDJoXI+Wa20Uaps
afY/iU34c9vGwgYwCjWYGiHWzW2qW2zKCcP0Jmy+zcTGq4GHpxL3Ol9gsFsA+Jm6
OErggXzb9dvToWF90wtYUlMnoLuUqqKe4R4Vws8oYE74L+JeY1ODvPJlTBoAcytE
YgevFAWOJPm8IOuKFIomqPYOU4pa3ej0Ty5f6pMzpms8HmPEnny0DoF/UOcocCVG
LPKxL+JaEmvOFg1uvwV7oN1pJLKBr4wGet8XnKM5/pk95qfjoDRMlSg+Xj11hfir
Cdx/P1nO7afs5Gr9Y4QJbfo1n7RANPUakt2His4C8rBociAvGk3yKOAJJ0b+txZD
HLAwOSRqmOwh0u6S55aMqFXCXWbfMDKEVjz2MBrhXBHh0JwVlMw9sNT2oXyXmer1
WeVz2SeM6MJrZ/Wpr39LHRJOwKvkad1ZPI9XDfhkZPQ3AlnD19ovB+dtMuXe4IHY
qGhFp6ZPQZdsx3hYA48uNXvOOnYplAfxQ/LZunNoIB5tl4Rio3kBQLIDqAgAwmaa
n8CMmxZ1Cg+lPtzuxyL3YYSv4aD7i8Ca94I3LBqM5xeSodn11iJ+tFJuq8cu9Vhx
oihJ0tH5VxJMKgRk19GuRfUwslziDHu8Fxf0QvPLZeCmGEbFF9i4EMlwdwP97BSJ
bdvafeJfxkKzRP3o+yQIHUPWMn/CDCVJGNGuE/mGKi5Pq2ymh9PBV+HEOxAKVFdB
vHM4UxlpX3LkFO9iTg+kkEEHue5MlnOHID/Fs40pCJSUg7GwdA5/XMMaFo7Z/c1z
YBdgi7g5iOQEoh6TOBc/2+5eL/68Pg9hgO/LT10a+IOpFyxIOg19rOzwgLrs1N6m
n7vp7/78sR6dM/dqj8rYSlLYksCNxUURsne16M7gg4sY85S2TgOnIBqFaIuVfZ2D
UduwHcZ44x4xVBtUJSorbiBlDT8Vs1IZe3d5xGUeQB3IP3rIxfsURkW1Pz+bXcqD
arTb6JmrI2G4Ia0WjAGEvySUFCNp90KELRxE65Rl1HpnhLgz4IjV3BdPlxGdqlGT
J0AHmLvRbP3gy+duTW0Oj/81w5SbpjvsdYvN+lsQrgCZu9AQ5I0fTlYWTVC0Vul3
84sPUDAq/B3RL2kio8VttJ5kxIFeYJ4tXhw6LJ52kEQlRg0+jx6uTPX5kN+pVObK
nOrOAY42RfVj9s7jMivKOanA1HnPK9NJ1KrAtrT9cQt5UEf+jw82eNMskHdMC5IV
3FBcco/U3ZzPOSWUa4YloGYl8G+7wgcpJKRnsw4QPQuR6V0qlJBBf3KwSI1Kmhi4
LMkrbekeD6M+F8F2vvW9gZIrWhV4fbkVgOaeERTm7kXsbWxQcGf9814b5t4lS3pE
gIUwZmlOEf0OsZfSKsd+/6SFdc2qhehnTWSqMko2xK8na1PdUT2OiqCsSAZZeS4X
sq+zcNzhZVTtv8Fq1ERte7XFC9bXr+p9uiJpq/q9fckPr4v/FMd4sJX+BZAN6itL
MNGzy8npNCA96cwUxBcOojOngYs8qoARz1ym+o7iDo0LYOyLpOrmbuPbxXTLQRAP
T1UdSgkJ0ZWBq3SqFVOwF2TtjypaOvQv3fHx9PknvsXM9YpFTWYYzASDY19J8lrk
MhKjhYVKucIyTPv6pl9KO9uCzNRi6bgF5L37HIjt1UEVYBRKK0xUT1v4SYFn7oJC
ZeTCEFqgQXlmXbyKWLSZrUGt+IPZeJjt+ZGqEP4cmVa4Cz7pYRSV0WFKuWBbwiwM
UzWcMB/8wv/eP1xIlcULmoEsRhMJcBD6fh9yIHUU2uRTEy0CW86DD0oO4doZHc9A
7daAL+UmzwjZIt/XtKTh6oQ7Tu/vHCPVcqlUwZc6Itx//g5srB7g1anPX+eYNeH9
IZHbs6+g/apEt6ExB+hUE5HN6eQmjuRgz6vKNW+ZpWHmRhBTVliYPrFF0j5t+lTm
iSqkzNBU+nowtQw47eWSyKf9tUPyBS9oXKW0DUcwagFzE7LGC+YR70wNqZITwjq5
+hf5M/y/hZw9RDsegWyO+mu8r6losvnvYCbrgpU4TxumnWuVBQsGF0NH//LyoHj9
v53XglhK/FTS2D7LpFvKzn4oYEfVj8B3FEORc6eSPlpA5867eDWWhJMvOT2IME9M
uhjbQuD6KERMoYNSvjQue0xlMy5FRQvtqGZumBn7Cbv0lWIXwzTu3qz2QWWIndH+
uH+7JWI/6I8E0X0D6Iw4TtzPW/6W3Wn70lwpWbZOqVDr9uVcQO1WFvbcJr3t6iUs
DNOwc+LgZtbKwOPtnh3EFUv2xV3cqSGLY4e3OPvNE4cdp1M7BUES+chi+uXaE/D2
etBgt1ZEFSS8C8YO8rH/xiLesquomtSPrV0n4Pzq9igAQBukbfCPbcLqDXWsX5/n
e33FT6NdhRCcubvqQfwN/+TJpjQ9bD9t36XW/OJRTnUm5PNtFOvKjYvh0DBuSgFK
SrXufzA7TiMOsp9dBRuLgv3pV3sA8hi1cJB+778YUKO4J9qtcg/Keu+aM6wMcjyT
FW65yG/8RQL7YqUdk15RaSWCRCqor1sMRMAHNMRM3KudQQFgQBtZWCSXViAjSTBS
7dcHz4Kj4VW2HZkHJW6k4jbWK76cTWujflQgK9FpRLVh/qtBT8QDxnEOa118r1Vi
HwyebyJi92VfZwvZO9Zun0s/h7he0tsOPXIu/d8acge+rpG5JQbtIswKV4ct8dMD
bNT+P8ML6GXCHPy5/eSPV1/bByTVowtDS1WvWlhgGC7zduM8zHHkp+oqQI7hVNfU
3X3i8ZT5kkvxwuAndNquDx6Upaoh5XPthnzUif6nvHZJ5J7f/pqqOE6pzBGQKlHA
XZIge/TMG6qnSr9XFs4roVqbxwo++rhHwg+dCx/qhDg5yIpG/4tPEuK8Y0uy89+O
qmu8cZwv0cVp5uWc9QKzu/S3RLTVm0gG70ns4rensDti6EeKE8Zmr6HPiip/p38r
G8ys6xNKBaUH2EInAiKpJz/QdaDD8nHzJBtR/rXPkfeMoI9sauNir9Bc3Lchqs4J
e23ZrAxBta3/G4CjCI2lIVHh9Nj/TKkqYQ+dAs87j6ozarBXjBo+ihV24lkeZdXq
I5V6gAgn/pQDM9cfPDGm308MOmmPen7WFUi690qgMqOZhL7Uk+VmNTFHS1iRpNo7
AeC6lgQCpMWj83/YBvH8O1QzsjpICS3/UYyC9bctx5vuPugMgs2odhoz6VBjaud/
tvEZBMwhY/rVbgY5wdSBMMkwLSEzTG9gMd/KDVlRjASURj9c9wVcumcWnuJNQT5S
iNQ00vtBgzLnHmbqMic0wDnthv9J5XsJu34nHPN5DAlevS5nPZyoWCxLy0CzFz/u
UDb3tgdD45ZhWdGeX3LVNmdBcTMLc6c20lAQi7MDR1bLWYBwxOMrLDJuAvZSvlNs
EJHWFIdVHwIm0Ai2CpqU2UVlsHrWsmWwoTSgFo6dBWa/8LYsoVsvUhH8s2/jw0Ub
8/zh5gwrSFV8Z5KL9k0DyWwCD/F5bNcC2f+2H3f4aN/6M+lD1y15FeFkKYNpPS9U
csArzdDa7kRr+3+yeZK+fU0LdoImd7x4A+zH3Ao/hXrtwlklFtoV4T+ZoPrDOZU7
jR+k+C4S7lanieG/ZtykXBBPCO+HrOmvCwwuX4glCFMYVTyTfUHm60aPIUObyPy2
MDXrRpdjDHZvP128GmrEtorYEMK4TKq5wfYvydcnfN1z4C1k9iOxEagtRaXxjEpG
jc9pip5xCvq3JG86OU80IvzKyyhPMSckj9PE6g2wHlwUKc1lkfaatgr6q4aY5REO
q92COblINN58lvVA/tjwPVUnj6Mc+hlnV+tIxBxrkRe4l4Rrugg4QLwwhC/LSreP
ha/qwn0AM0IJoicXvUPx/en/1UktSxRkoS8WUEda+9IS5H/omIHBvwxXZYGrD9jU
vS8KnAVsTOBPG1OUS0AmmNT1q+gWNJKbDpwfu+snSkuqwOTdcO0OpUZVYx5uzX14
lbZ0ChIgIabbC6LK67TP9+27s6qTKPSy/zh5hjRWeHZi4TVmf9I1sQtLS7O6+Y+g
uFjVX/dgjt2BdVA6hW5pPcjQiTZabwQk/MH4dTQ+RSEgdJ0pyq67BQ6tk5vfpPjb
8VSXhOtvPD8DcAYoL3KgLTIUkS5qZSIbYbCTlhS06ZUpSsu5OEJjGvO2bIkL/kaK
yyX7E+uQUwyqS6xlEuVIdRRyXjm9JMFxA6GIxsWxz+KnesmhRCD/H95zonqqCzdY
Bt30cNAh2Iojwje0D2oKO+an4+54NbhP54H5wViVg0U4oY6pAc5VUWeXBZYW8vGB
ZknSs7PyxFoYEH/16V00SRN3SWwfuyPwhfD66dGF1bAqt2xRfSJcyJIVAcBrPv7S
/RRF1kDjUdyj2ts7UsKSPdTNOeAAaWyy4EE5ggCNXL1/weZ9K6yGGhYtvNzi+gcs
1s6BHgG52pI+8hMOpNGuWZJ4Co+oH8bsmU//YZFWHcE7SZxdudZJ43L+anElYK//
1wi9j0feqlZrApJlUV13dCzjFG8mDMyOJkV8DfLMIVIn+d+d54XQr16e99FMAv1a
UDG3vVJZyE6V+mdx1aniYvUe3zr930c6mxrTB2BpgidYhBfc0UMFc2dzQuMC/YQR
aGiNgRpGK76IXSMHORq8d+51CgTCzJEsRAFkCvpgbZiT3Tf9aV26vQUIJYtOFYz+
QTcuO2+IGLELJPT949mnndi4tdr40EZLrNwYeR8ZJyObG3loIfsBfeIIAyGLLSwr
uFmnPCK1zYjH63dcAK0u0/DitWI8aFApf/3t6B+L6GFlsXX76sh2cMvIZ5oqucKU
Z28+MVhjHAS2uCnXbX53Z5TYIR/n9y4Am2yDx6LUXTTk5POjKivL7Z+ZoU0CT1iL
KyjAiPuQlYvQlixHo65A6M6RApwcjaIN8mvzJ+TEXDJkY2qkA/zrnTNBfJ5gc9r7
mD5IDrXCw48lQbIjh+dozQX8yN6vm3arFg5frKTiD4wdie3dC2nMZu9dDrlCf3RC
JS0d1yU4e1CKwEAxj31ZQyXXDujEngcc2KDX5kdvLTexZLoe+9xyAau3nPm/gsjz
37NTvUfyIUoAMqAWe5HuOZDKObolX8z7WQST/dx52sEsjncm8mN1PL8HdugtzXMV
FPT2a/r+kQUeLR0WlW41LB4r2BKx6kcndNVufCeogtG1RMyzy1rCuI74KqUX3c8q
JdQpJiQrUrv9GqVvshTfu3ci2NgeYS/wUf/wuZKQG60dYXIGJj9WnxGJkQp0UmOA
JmwYdT14ZT1JoQgo5D26zDMXPLsg3m4Jn/sI270qOXzA3IS9dUTI8qnDflHkkVT4
9pleQR6j/WblPC2p6u2Dx9fZ33OhNiXf4b49QtOFbN7/cY9Xnch0aCCzI4ruU+Nx
hrJsiCFEsxIOXU5kPNfias/Bany65JfskF3/+EHaWEV0anEv+AMS00etYSN0S3UC
jDFj5cWVqiuOWfexPLz1yynKsLYBda1AGO8Jho8sym5yxol8ZM8Pb5msFsZP0Lid
/YUbvlhdFhqPOUJSXIX51PyY34IL1dOTUaDos0BIUs5e0b5cwl1Hd4gp16f7VhD3
JYWtGoiTpI715GkK/d9WOoFLehaK8kQphGR/wFQsmAHKLRP63W2r3UD7WihvQiiv
GAWJHjs7ufzRNSiiVcL5A5E36fycPfeO8Go66K4fwDQcq10OBbwEieX8931upCIM
DU4QVsIYiaQu38DAvtLDkRYg6bmLR72/7KCsYLMOCV3s7rwT8kaneyo50GWDPlU3
6OE4KzkBqnRziMuvjpnQikFqkBGJ10xPR+BT8LyO/c+Ts1V0ROIm9u6Ls/9YMXA/
UPF1U09jmd69eN6XQ4zAthwOrhZ1IArpngyoXVljweHRmG0VeewCOd2ukWY/Ug6s
cEJ4qVZv4lE1lz+ocU8JGmY+cZpC9TH+RQ1QR/YLydS6EHcn7NRG0mMzOYchBqO4
b/lB4LFsEhmPD9kd/z6H5IuxO4+SgXLVZuQ946MznHA8H3twljurlGJSmUz8k4mt
AvGUV9LsuPS/7BzT2+hsSjC2hnB0SxItCNTR5evxopPrvtIj41mzmeWPiRievwXE
TxesiF+h6D2cwkznl7NuGTrlFhndyaW8L37Zm1l7YP4EtzQa0Iw7H0dX3zJehqKh
PPXLhyTyMwY5uzeZtELUK6pG8yHid0wECBZ1lxKabD0+JLDXVIm2LUE8TpWwpMb+
KKDk9R000JlZ3KnV5QIt4IHc/7sWk2rH1OZkTEfBxSLzU+G8MIrwwO70Y1elR6Ql
WE1pQ4yMPCZYTmEHT1b1Px/LfVuQYFNVY6XkNfwkY1tPEGn64U2cKhSCxgHqpMMU
D8e5Ll1SAeBVOPkHwIYNHlUXgb29CGFClxnJQ6VP9SrGxWUT1P4GSa+4u+FUUCc1
/kuKCbQpqtzq0MfssxJm3YUV8T4GcJug6PlP34hLLSK+9P4ot8aZ6sjqNKhFx9/o
KyPkrj3skMjwDg7nomCVFEtkMzopHfwLQfLuwqf9DiRUpDy2gzlY0MWkmcgoR50Z
Etd9V8IcQQjexVjXdCfS89YBKyGbWJGjx3JDXvX47tn7f64O3X76ay4pr4dnG4Js
jxRTJHzNmzb2QGEAXlZ27IbxIoPfksmN5pvSQ42OaZR8x/pileuOZGhKSWM66/UQ
rKyBbolcjBcT3/OUI8Jktp/UvApKyU5Zo+Dor1VH/sb2p0qqP7JhUwvZYFDGu8BQ
owwQXJb7o57taPE48RgyOLmuu+usaox9SxDQBvjbrLHPgHZY3vnC8fETbGQ3i8TJ
suJoSgqBmbjriwAFK2bYUl9OxVlMXi7Inp0AX7K1kAQhWEe2xOgZotFMHmq019pA
3Bpw4frRyLB/OnFLaen7WUYmZvOyML+T4aR/Z7n0BYRordVCzY9Mf9SEnHa1TngM
KXE7iahT2YyhOQnhR2+l4GMg/rVWG/+LpYN6+VCgy8eWTlXPIPwlrvER2XkrVGYe
mMaY4+hEs0HZbYZk6l3EbhpSfRfw4mpS01E3Ct3pjQQ9xm66uBW7SW+mDVfxtbHW
ai44cBmhPgUX3nnM5lcGEYYykrZRI/NcOskoBhj7fRCb51C9xvHfpOYh7Mkgm/gh
ZM2s/eKYLcUGF7jvqt3ZO4IQb5ae7UxcO7d4R39ohR2cQrqXQFhMmhwQ2G9GYsXl
FNh8QNBPrHrzij+58L2dOuTLksPGEVUf5BJmJbgnDukjOyn2L5c0Bj3+aMof2uvu
UT6vKpLkpbceFiTTHKAmMBoyY6gez+Aj/fCyeHcrV6NRUz5RRAYIdxIVG9zvvfnL
UwSlbWUJI4O9GV2rItcMhaUALkO9MF6hs0+09Z7ZPesa3TsWtTkTHa8k8WoL3YBi
w2n4g+fdjGzlrsMogVfrmKjxfJUrbQwUwGGml36AR8vwOsuik96zchnHjoOjHkxh
EXfJ1cJoAlDUEQl5xKN+WfuJFMQtInu/pmMns2FSkB8PzbfrGCLMr+cIDc+6ZwDa
yR+UDoddXPMaWftxEPQMynM97RcW70mXkmXfBTeg9LklzQR7QAnogqFtdpBSFp2L
ajN/7NMG5NTyNM/WLTOBZE6OrEKFo4qBiXiOzjmVz/zbEoCHqidOroxD/wHPer6a
mRmvO3wtKajvyYUdL20KeRvdoGBc2849mGxE/QZ8CHxLSN9llOA4qqwp/0i2JahX
L8el5J34Fh1puedOxO5Eulgl1t/11Mq7NElw6R/kv49b3urx36b2Vj9KOfzD8GmX
4VoBvemMYGPjFLH2c+2A1oTtn14NFMdK4z5VdCIUIUf7L9pqLBkah4CeeSTXJGZp
oD85vwror3USqp49z0Yt9PvWZXVSBXB0wSAErT/r8yA7Nc/EDwA1Q+QDP+1HVzum
QicZXJyYxbeq4y12MQNYkjeSyY4lqBUMgUsPUQPqi3T++zyTmzognF9SpHxtIcvo
yr5iE1NxkWuW/5JxUDaLhXq+YUfG5Nsv2yArQTTs97aimG0hIomF+pOQ9WKiYooo
xVIkxW5DbK25vTNiX+oAXJ58O1zH7MKUORq1MmEIPqgF/T+rU3v5kjyEG+AOCbt9
PnQFGj09NXRoggVdE+IRp3617LhcIAMtyTPKQ3/qXWv7p7c0ghOJ+wxVDaqxPQIP
ebLX9Cn07kMr9JCiVvqK3D8cGBI5xpzgTJam8XaZlYsc4cKxUZhe16LWk9ZkMfTa
6yNLu7Uat15JfSxtS8eB33obidrQA3Ki6FAnk673JwPM4KMH7jgZ+CuYwRD3GlHW
VizPTEE14KagBDFoSAML096JVdd7Zqe9sdFEu92ziEoH6jW2XmruDbWgglLKzRP4
8NAmc4fMPHzt5uGGHJkrKt6iAy2vXMp+qkV6SqWJKYwjwCaR3LSCd4/EGWmnlBiD
9ncQKjTj0YSwAV6ZHjtdrWcIxuXeBqTin3rqNIJHFNL//cbv2GmclF+5GGQcnt+x
jR+ESMgjJRfCQOPqg1tkarXo+4PilmsAArGN2V0kZIWV6ezMpJPDfpMb8wrQsid8
ZtUbrMPCa5rIaOy8wykzUGdVeH/nQg3/moLDbNrGyuuOydihFd4AKVxH2oYV75Tq
QXN0IgNk4vzyIMV3H2zj6w+4pP9NZZvGbJmDvjeY9N1olzIt+3LwNZmEJhuh32xX
cKa55ZD8M/iVDGp8HlPJjKesYHjrUoJ8/m4ChGxrkMMx5GO3SZnPp4sBAzd2/7d6
zXVijz7h0MD6eJ/cvuAWKZ9Hgp1td/sAZqv2s3zt1Imx3k1YOZeULL1b6Ng4g5PS
+0EKvFTxnE/FrECIjlKkHc4YepJUQK+pETAc5Fb/vbuSvO49xKSeCFRX/u39UGOo
fdLkQ9jm3w+vh5xqQaPA7YQ7ZJ9OUdxy32a6CwwwNbey2tXs+SQcjfh38VPdduER
nxRfHUo/lnMRHjpbk4XjZhDgSQ4uvGsudC3dFDSNyoUtJB6XNKizqSG8o+9/2kTR
z+mqKkrwZzVoV0dImFj255vH0n9w0a54e+VVNFhMCBNaggkKQ3vmIm0MbNGQx7cV
AkxvxqXX1aOYfofMK0n/Gbyu1JsPGrCQpgi9lRN1sE3IJqEzO/zKT2haqbhIl7qV
bxjG5HgHICiAGFTQe6omRcy+jiCn1yHEPTz3B8v1qotY83/hgnjtOjhqeuEEv9or
uAGnvj1O+EtevmPBGE630OLj97t2cq8/qsZV3Z1dSZGKONTOgf4jnnqLmdFuDgT0
Vc9Ys5BDeIjKDjfHV+ZA/nlBrhr7OuUQYJ8mrTHvy2SNxiObUxAwiCYJTfngLdO9
KaRY4obpU4wEO/u3angjS0WxxTNRSSEeh1QjQRynfK8Sz5EbzzVs9px/MMrkfX4p
RV8rromYFTB9H7wLlISTWLBi1bQUBHGi3QyVHA1oVrTBy1TzCk80hFGt09mLDXaE
BJJafGxQ0QJye4Ooz0yIWKl2hCeu9wqD3AJf7t6aZ2+i8o4yqqyQ8DFhB3sk4DZp
qAV2LTLlv+1GC/F0Jb2j97GMQjC2F0xYiv8efeJSiSd9aGKkHJh2H6p5dHX7LkHK
fpmaH8GkQN20C3+CENBpMMD8XcrCSG+PT8P9S/3cc3qdG5y28RzUc7eMada9yFM+
VOHyCnW19s1rZzhADf7btDmpZUacMScOeDasN8WNYam+0R+VIWmot5qmuJvH+i0g
eXvsrlbakAMbb/zCpicIPGv2qCssTwwZGcsyESKV4gRUnmfN8RjQi3ugJXzE620T
pO/Uk2UCN4jE8HLbBHmCjzOy2BUg7mV2KeZTEUd2giQMj4ZHT9oaWq5TZRQ5o0Kn
VjCoJKLP8N1Y8UsBZLJB4UMtE67Tk9vcRKkIfodO2d5DCuMoX9gaRZH40AMD73CY
G6b6GhDAeAFbbaAtE7S1HUBMTNmgFDFCYmq6VEBYGqMVmShF4onucqqzt6b0uIpW
ylls7Zbr4lyBZK8ZGaW/P3Vi6EJvvUQJuxUiAZPiyfZNEHXrwW07uzeHWLYZ3/Fj
iSDICOGJ7IKsbeA0UCqwAfCSrJYekAfqqjPrHtFwSahPY29vHg+ROiabnPtsDdcV
nGliijHDFP7EKEwXot6U2AkAbKWCQ3HdTPP3XIdFn0aIvzLgYljqMhjZZ4kRxjMH
nH8ozu9FmUjyZ7j8TclHVBK5gQSXkOnKQlOxyT4tLVV4m7tzJnd+oLJ8k7tcr83l
wN3w2hiF678+UpeXFCcK+bjeuVnTKBXO6z6osTnUmSvVCNiZExt+9i74P5m0repp
oGAlVJs2mm73zHexhDKzYCiuU8yhG5LrZiaz9ngnN3i3I/yuu4JUFXxrtste+WVG
cWbaluQRPkMucrCl9RMTw++9kVaCSsSclGnxPxHV/3wASs+3HBXEEyPuXCw0Zp4c
S2+tLxYD/cacpy1YFZgxcRtPCqyabnlhQdOCC2UPxa3sMElNdwMFR+pip38eT+wc
7kREh7g+/+nHhR9vuAzhtfdr3kJAeKaPGLkfTn1jeUAEadbRKAI8CuV4GeqH3xzD
YqtSs4/BhauK836R63a+9s2rW5T9rSYSWYFJ9X/s26GUKgkSUrOmpXaKaln3Dt/N
xH8dxe1U0ymm1rkNuSZFh6Mj0rqNeCcMH6mfAlMgL+U/JYtddxzSkZKx3xhXg+lc
25wj4QuvUDbEj4rGfQQlhIXRHzEU+wPVHl99k7hq3/wbzXwVKEfGyMkAffruIHsO
XzfrM0X6o6cOUi4NvhV2gLa88AYy/UkipYdmJF+2EwaVC77P6ywrRGdMIziQF1tC
bBUpAiMujK3dO9TJz+d2Pibc326VTbjfbppbx3IbwtiuInuSKxe5mJ3gtrNaAVk7
6I+ye3SvAB8aBK/artr3DfJSod4C3cYy1XhDTEiIsaKa6g05MfNJOfvC768m4DtZ
t2yotfVFvrYR+jlPu891yuaMrPFDF3omPRcN8g72VQPpG1+vr1TNpMxE0BdGQH52
/sRq8C71fKtHKSQiMd0owLT2SusDyYZqHzKXXX0faGDDFeRpS6VkSFfA1fIeR4xl
VJzopW/uEjEq3ozHcC5tBoihNj5gw0y9NqzwQshedfV/AQB918IO+9yvKPpamAJ1
vdGzquSqMYsseYhXM//YMabqlhhC4EQ8y7AqCZR8rSeLslAvRF77sIuuOMRvvt6t
MQOttx8ZaLcU0MYDpBHTAbHFWofoYo98N2AUueJ7lGikWWYh6Rqfc0xdaaGR+V7k
1ioOaQ8VxPbwEQENquYdCnWfbPZP0XILso2NAHDGkbva5Qpltwo+DwmQB0kyGRCe
iGhX8ScohMYjJ2jkMLnLYyRKHmJORCpFtdRStdGsZjT/I1jx/R1UUaw+XuqadFUJ
pMvK/uQ0jc+gWxs9cJd5Adtj8fiVTkRHL8OTiK5/5yUrIfLrWvsZTdchl76GRqB0
v+26IdSUjJOxTUAoc0xWOcRbIWy2LyKdGLLR0MKHObrM4ywlasKYUQ3GTcXVcHLQ
oTUdjal/gXWxo6LphOhsqG8IpxmTCPig6pfZr6tKnV+aGtCiR+jFg54hh9HMLEeB
BukuIbggp+uoSwnQSONd/v791ibiS3x9TVCSQBI6SXxRpqHw0zCMyIMIepaQnFL4
1TxJIFR77CBL9PTRUulcr8inFiLsFa5ucc+hR9T9n8CA1M7jbdPeo+XSiYmwWr2N
w5m8YwafzpeSDlVBBpB300n60mVX4gKDZauFasHXYws3UUZ0Ym86WvG9nBMG5VAO
a9yN/b6x9t8pfnnYzwe1D++z3lZJ22VsQot+dEelZqzLBmKamfBNLCm9GNECZnHI
wkgplHepMmJ+VDdZ2nVPcgCNESD3PXgnPtMbdU8Gj2AFW//XS4euCPhd7azbEB1h
kZ9yl8kwiE2AyDisVaY4I72vt+c9gkoERWE5MWziVXyTG2V5dgSAFLp0QIQT3OOK
ISauwiOMlGJLgj19BUxIaNIE7by8YPxvnmrca5+iVn5jiXRyDRW3fRb4kWfL5aq7
h6KqONIecd7ZySWUxotOWKqKHzgNpz+mmUyUmAMhhVGsBdquN/XT2UlqiODhI2B9
RYKBfJqDamrkc5VKMTJWiuYtuAcch/JXNQRIi9tcELPWsB86QP8wktCs71Ee/X9a
D8UQBOGha6qBZUUPIt7c3J6uV5vMxXVvNXWXS9iwc4X4SC3twNdvioiciKemCPus
u4SMFq3e7FXFdM4f656RC0YOHsHNRODTlfRN6m30j7bj1LbKHLKcLipSsSmXIbV9
woixQa8Q6I/Hx+/+majmK2l7S8pSrmZCo1+ucPQTQRta4OD3i/HYXKzXZnYDH1yf
8jTVBjdWKkzRW4y9k4aG++pMQVxZQfQ40PFhhevKqsnvZY/jmVSO+6YGlOvAUmQV
AuoqVXlnjpMRZP8VNNN0KPnUVbwpVX5qKTrZso/n6KEV1nmil5th3m8pZWIpKb2s
zkaXDs1L49qGm3GQOIsVMA/SQLEc74sDw8wHt+9Q5dUw0jNsapLy9rrIZGWefYwW
/h6pwNsIYIayy58BufF6B0YXIOMB9+Fbz+fcskOcZi2BV8pvxGuioErYBiaFyrHv
zxGXPdPauoDmcdtJBzJ8ZvQoSZ1J32gmlm7n5C/XGuJ0nx9qdeKL9odw2i7/h20q
WrHjEbEuhLqGn/SEo3iBW9sCINnxhWknMDfRJy+4owHXOl7f1Dv4cIzjCScThPMx
9In+GVYFASX57szrn4Cj1BFqQ1v4e5A8Y3h0X5/e3MNslqY2YYMG2hrnQK0FdIhQ
6BbjPbsq/dpY5JUYi4pCFjkVD6ZIg1c2MZO4LYxIkx+laIiJwlS0okyUGTx4991R
U67oGZylQUubSJ2sXHpfK+Wa32ROky8ty13rY5oduuLSJkgBhBlGEu2royTRpjRG
6U9iP0dhFMaXSxdfwBAOR90L70EODNXKkPdn5xEGU0Pv2ISE3HwM2WAhSUS30P6r
AlKHmK7dXlCbLJiOsXo8YspuXKc8Te/V9h13LNPib7IFJo/dIUZrNeTlDJomDpBc
NIH8/rY+9TvP4hByxcEUyvpx+et+MrANRLqMHTWyuOerFD9M+P5o67ShN1y2qMH7
pMU198r2G6hC2FHYV6ZTTkSpCZrLH0dWTEyN7NeGBH4RqNd4vdXoXLNKDwyLXqt3
+PA3jOgRfrf857rlZH1F5Ba3n1bFibuSK9XkO2kJB3ifKXZblnj0nss06Up3xZd4
UGiPl2C/iA+lSf1fqPK0NHEa81cl2uIVEDrPUUvgd3j8yThdcpzECRcNqGismN+z
QBzayt2Nuh3ngMW9veDK2GaflRwBttxJXKvwM4YoGDuvZFsvb3n+LYmf/ihaj0EX
MgbliWli2Okf9FEI6cwTjGG7YKODcuAfnct2xWeJmqhRaQoz28eCpzuUj2RLkh5q
0DbzJaTNQuv1vVYZ+B+bSz/NtjW9o8JJQOkmrHN9W+klnNm/06HhhvS7tLZst8hg
987e6zu61Xg74t0dJ2q8H6mkTuw3cbxJFCvj/23gqTqQbLfxh0kbH3Uhsv6q8NEY
/Kl0HruLvfWLpMIWT4q674VMDjK+ou9bUbJph1MiAfvm9+KbQlUZkdmnT6S/EtnZ
omLn0dPsZiGEzgOYiM7o0xu26//4MCNEc9q4frzHBrjach2j8c/qOr1nlhWqywni
VZdFROT2FowwEFS26Fa7nUJ/3pevbOZSnRPfhJoycZzgtJuSXN5tuSo8zbdI4wKa
dMD3RTCXVWLd9iCi800VCCAWT4OQ7lWCubbjJEQ9YmcKT05Ef/5S8xqgQl08rCWs
n35/dQbbUQRwTpuz8hquJBpzvQcryY/H1mDIVS2NWyEYV8oq38+Xtl18wSAo/cqW
5vM9NAJSSByd8aJw8E8w8KB3u/1kKheVw/NcCH1qfoq8No5CEriyS/a5FiweN6X5
qaCT40uGbRsIKpe8/swsk/QBo90kyRdbstp6+fFM1iNeDwiCc+botFCWHL9Qk88a
xzSX8G9Eqvg7GKTYyVJ3G3jHOJ3fOfRAlj5k8UyfCTmRI5XDixIe8+b2qVhu6wdy
pSE9zGnK+LfcemWaXlDVqEda3A4zTYLlC2jLoJjZ02LBtrD0uIr3Ui5d1g8JlnBt
ja3QUPSTLoZGEXc1kL2RJ3mktNeQWeOd0x3liUcwcsf2OrQCCQsoq5vuhZrgMrna
jJGaz6qZS3nKLmFeDoEI2ikcmM2c7DMS3wdhxetTn8yXUFq14FH8MOf4hXxRHSp6
VdP1ooGriKIEqRuXXibedwiXytJFrsowZOgZH8QTbC6Em9tZGoAal9WRITXmrniZ
exEv/oNrUi32JrZNsJn/7cpg9u3WiO6UXHm4YoWMiJfWICV8WozSimGbH3M3j24O
Gk3YrXM4h0pB3g9TqrgtXwHq8rO4mbMaLPhlPM2qlghNu0n5my6vTa5me3d1RcbE
CV5uaYJvDe4Bj+mEsWEtiMg+hrrIpohpHUCEPLtl6qFs4HITPhTvXMEZwQ/YAUPN
4QPBSh6Vn0Lfa/10prAEMuoauJ2Bgw94ZVHNibe2AlnjqN07/sUH9zsQ63Yqik3V
2HWRnkSPgpXkvHVDr74art4ornts67uhRDm/g53kIKbrXUcsQDCtdErie87hPRfz
xyIbwJu8E8oDUjpGA/+66P1mMxuGU0H4+SqP7c1P6EPRPjdAfSu9tFBs6oZajVIh
rOa8nNb8Rcd35gTOsACsoFQJZ5d+/La9xhIPaodtWHq0ERJFlRcDgPXIdly2SJc2
EeBpAZXlT4G7zXD11EkpfDlJllT4LwSAhOa55hBmg1Z/WJhwhawNOkjgUYubY7+P
NrzHc2bigopR0Ackmw6SKhcome5/9sqeus8LZYM8Fy1w+oL5uqNgjlcPLqu24d68
cHPnScvFk22LP+4diUnErISw8ELX0NDKEghRAt1PdrJKD4BA6iIiqDSeeuvzoiA3
xNM5Kk6TKySS7RMsepTRgaRYGQ020V19QSSWEzmRhF128TD16PakEMU8XbQoTlsx
f12wVfyKEneDTxH3CnXVkjpZNdV75MkTPdlAoJuV4LiL1oZY3p90v7P4gSD64UHw
LIRTbBiJuQp/tiZB2H97mxotYleTVStnUelQqpYsw0yS3TvJKFlJTjoTeliChqZc
0zX1suVgUDaC3X1J523LDI54eANJejGFCi4UonS1ka6z63/pGKvx2w1rYMwyDZcA
4A0wRj+hOEJE+estr1nRCHnEldhBnG+BXT6a8vZo66vTkqfREY/eyvTBU283AvNo
7NaAaxyvWxrR6kYtFHDLV5E/ATywTfCam7dZ+6TNmDsVkc0CD0bmPnNjV9UqiFTK
gjF7FUp0tV6qYW1O6DhVX2v1aaT+FmCf/j2/Wo9lZreUt5Nz6S1C5XF2AmCygvRF
eN13GUMg10XZiWJW0I6ysi11mQmfnpZi7IZMdtbSKdi9mH99QDZ9uu/jaQMeBp24
SoP2B7TTW6D5r9CdSO73+o3ocs6oZlBmajaQtte2G6KHUBAB5TZRbg3vB0DHCGws
nCxMZrlIqXfyEMl70tNfgMK60kL5jtu6nKc/rrPwaH4nIv5sWMfmIlVlFYl902yU
QJij0F7jGlR2Hq1MUZDrPZxVBldKkHKHr9rx6LFGViGp3Dj3DMfqOrj1qxR7MjGI
WgNGHOs+C89lbV3ID8Ku1wgj7Iq6qMvi6rrLXPVvQ6IBos5hiXxtdNOcYohB+DHt
BDCY1g27oIwVB8Vf+xXAAqIx5nHuglJ7EvZDnU3EzhbSQB4d5GH3FlyPGPSBpLqC
ckjdJJx41OouT4yetKhaUwC7IfI2SEVN/1I/+MuMZjaW+/h4kockAwfySj8AJc3N
u4i1zMSYQt+7Chr88e7UDP52sOKztn+XJAl7URLpX9TUXyKOtUY+kAl6pQchklSO
wgHnKYMqpk6Y1kBka9803a8kZu0exoxgCPEwSlVKIhRSJSRGuYflLhv9znQyf3uV
7kkj7dZgDLRMa67vW6bBpK72oV53+HnhDRbfAL1a1g9U5tP7pKzwrOQ7ZZVlznJ7
4fRt43i2ikklCQndyiX7Vt1L+SuSdsV8lBIrsbAwDqRh8/uV4lemj67T7Tt7n25M
r12Wz0T3nkzofi0CdiF7DpPX8O83dJu7BxU18p6Vv0h/sVF/ZBx3ATnanspeQo7v
nqbVH03aWwgnLSVs97aLGcFBa+41SEI5LPeLkFI7mRJ0O14TSLLiclbcZFFyuSHH
qzjDDAUs/VfW+g9tEXRU1vNXDEnA1CEOabsEIXfELNvU+gfOpUpTUAEzrazFQN97
U4aJnumdOA2dQKmzv4ZO31ASyLTz/Rwp17SbiVk+o9beEnK2XVE1r8xvfatv9gF4
x4QK+o+84BZnhwQA2sKU9VDO5EBY8xiPZ7ACKpOu7EkKYL/kVe1wHP1Pzsu01UDT
zK4J7WcexEnYWoHxa9QVZMNrOuKUA4wI0N0G27216GXz3dYg0r/nwvrFdv2aghIi
8/Ix4SNs8yO1Rizc5dy18REu8CkEzLWrcGwiwDHZYTpBwzb2mtV/E/+/pqmtfM6S
8ExpJYlg70U8cU3vtsn/XzfI38rx5PUvfqqji6fEzyqsbi1p8OuktUOVKP7zG6Fi
HuGoj1GvcwrzAV58dY6+FIGEYEr+7egShMIKIjYRM5F5AXMnYmE4XDGqiTquBVQE
MxzmXOku8xeywnmefEme+AbSKjgouwU5bCIOeFJvW7m4E98PIkXqaO/DtlI4MHb7
oTAY1Bf28xA9J6G80ZvO4F1gBz5tgj1wGsWcgFWERPlKl5Ap9Gf1C0yC/tJixbV6
Q0Ca++qvRH6sT1qCUgMZ1zbgsEq3HhXho+1K+PEMSRLKRH4kKR7jEdBjJWAKloB8
prxBK7Sa4SufiePbwEgi5s5SMwBSmctdcfaL6dgX5rZstEr6QdHXDutNYK0nmmiA
NGOFxD1RY8PJ+OwgCd8kMRdIdAq1Cc00awSKMnslM1MyHejucEHW//MMc1LEa2wL
PZZ1cjGex2caytH7MUQvXB6s8qhFoVCIQ5v97fH4nrFjLHDt5BhB3CkJSiaUWQMI
cFrRRiRdHCIWDnfKIyHy26r/7GBjBJcz+bFhMVCVa/jNyakFEQqqPxrh5/WqSDTl
B8BUy7Tm6KfzgBQxMAdZTHcTfhe4MI1y51IZ3cT6qRzN960en03m8lnZeH3njVCC
o429Xfd3khbT9c6Vqq9tHa7G8pkvbTkXYqFWJnqg+XA0pO71pjZSLc0QqenV2lwh
DYO158goVx2CwQuaEoVkkklq7+mjWJfB0R+dF2WE0pXuesldoZPD73zbRMFpwGx0
jwDcQhbchDwKXBNuU1dUtn2UwFD578YUu82h3Phw9XxkWWvh0G28Pyf7fEPiQDkB
tAKtbwisJd96u/GI9yEpgpi4ETmyMHrEaGvnagVMvZovdF/9H8mg7P8Bl8EaVBpc
4sHreNtDDNH5KhRR7ZjpvCj25RMgGfP2FTXFRwba5bnm5oUuqcuf/GC46XouvuaN
QW+0+eFke3QJctcOL1tjYvk2ueQ0IJfw5q3brGWNrQLkW/qJtoJQZaDKOwcd/XVs
V5QVfU1B05TCbZZySmSx/WD2Y3pbjiRHJUuchfLnzLdsItRMPYlRjY1LVIKPpgar
IovmhP5qbvcfyzU/L5DKJ1ryyB2ab1z1JHGCZA2uCyeuHqKxp6Fx3g1ug9fK5OiE
dbo6NDbAph0qvX8kcq5PNjSbJxWRppTah7QtdRfhPA406kpXjTFHCI/M0/PBkVQV
ZSA2ilW7n3YVovNLF99iFAHCxI+6ES99yfaG3cKaIUwcoo1tkyDWXa108sPRGkuK
x56VEzZhspY/WRWqpaPQf1p1yPBAGe/uls42huhk0RYTZRfn2BK0eNSPORAZ0AD6
E+oj0sloquekkS5shW6GEgvZYgE3WbGGFF/rMIm6y/4YNlUBVDX4J36cL4NcowmO
jDuqdya3W8jTWB4zHGukibStH/gghgmLucOAo3F7mBwv8Ojey7KsulWV4AFsoRr5
uIHGA1/zGsjsza/d0Ab5LKmU5+6nmE4NfpNCEgxykqjrxwciSvimTaWqILwl44U6
DpQ1tu0GRLuM1s/q7izLVspk1LXNjSqURqO3ABEsPoIAgAwEimingluhqM5zm6hH
j2/Qg8ohaXPPJ6HgU87MC0PC8/ahdKaWAGZ64cEQ5Xcp+ESaXYdENe6nRk/byYFt
lKufHuCvypAhxZsxBuMjdAQb8PDrsKgkwfxgYbGArVJ0jBJ9+rweWm/Dpwn0KVAJ
UPGA0Sq/RNBRhDF7CJKUWFjVBDST8hLw8DvQ5KR8uKW/Sni+cVD2Glzay7P/6zXF
mNuCYnaxHmOFp0PJyvZJigHvrhmUXgBkER6C/eanGqXVkBxT9JxolGPOto3eFblR
1HIP21ABbIriVc7mqsHyiwGAlYwiwrWvZxEQiGnE09aTap48iJ3tH5MV8X+1Guz6
Hj4aZ3NnhGnojWyD4R5Ii8mFy5q6qC1uugkiUu8zg8UNGWKR4yjKgpUYeKwknUdA
1aHaMw93A+fsoo8TlRtZar2/kt4BRynArXQWi1nTqIcjr9cemBNmRNFMayA3U+v7
gXORRjKoj2/EErhIZzHMTFnP1+5jDU4zuIse1wahC3Dx9/Glmvbx5vXyiVvOQ2Qt
TUzpGmBGsh6SjONBMNHUSgH0vFYKqO2MzSDgsJ1pCkEO7p4V77Y81vsU1TIBDPod
Ij6dvKFCgt7pPbzFt1Yu6L9dKdGM6fMMvKd+3Dmys3783xcMRug0za2EvO95CPVJ
OLXNodjVhYZXYf6C0ddlDOcUtE6vW9pPXp9WewcGa/ooYgznX/jLvZCk5OvdwrF1
Nx3uxpMgRHs1l+y/5TxiuMgrX7zcnaNAUiRP4X+lc3MrOCnQsJ3VZLymYLI0m52J
qLYzycC0Q1CVUs0b20C3+s35k4mLDhGshkoovxug3BvkzHfwcmbnFynbirvEu6wK
U/iK0qe2gU7PxP4xBFeenjFpHRtFX++O0pIJLNB9EJnNCSD9CEJbY9ozyAh51P5k
p7z00hfeFLgwXtEQUSrS5J8rSmyZMhlyVdXYfO0U48kI7eOiq4htX7XeY03rlJim
aWfC4V1K0IBFXe0z+PeU2Ieha1VeJw/FG9dGwQvHje+ZAbbQ3TqQqSWipCU31DZr
f5+OA1mqUDLxdb6F2QVdFmKMWeIVjyYcI0oSzZvCIqoA/WRTiswLZKE2edzAjhfy
ai1H1ZVFaXZFWjCBjSA9XroWagCi11gKeixD2Lb+S9SVoz+B3fifSRgai82tSEsv
6Dd6ZzgOZYyXlvIXOlNeHsKkmOts88gSqBH1cKtBRLbf/xr2+iUw3B6qjHPyHeli
C4nrDt2rvQvsgFwW35eeTE4q6yP1MxcbwovOZqazHGZg0qGGwEbvfLXpAWSnU4LM
FZoo7sy09ZGc+I49xwUJqHlBRwhgi56VPy8eqUWs6ypVDzAl92+lUUZ9X14I3BsD
DgaWv8L4IV6NJ9XzlQI7qyHni8/4+1ZLzuYISU3/XFe0IexU5ZRgGdUjc4ioxknM
xC3PwMCqI21d0psEkcpbaiUGjJoRfhhsNZj5wsDpclRAAkOsTZfuC8Cf1UhHFA8Y
mLmg2WT+9T4trnumah614MdMvD5bVPcHyX8v80HeY0I5+k5GF3Rj+tbEpudKF2kc
8PHITFAcC6eKSxzyf5nhog8XXZAwMJTR12VVqHujGp4vfijuoag2Yr+AK6vMOHQX
3MwyBBBmZrxu9CBpmV+PcrizcPhzkNlgcQLT51dkhHwgsfgLttM3l9qaT85PSS/t
yC9tWJ7+AoNJIWcTa2Kbe2a3Cy3eLwdp01FQ9FZrmzO5VoHbw/ELrY3mO7FPYH1b
ENATWcLxRuM8QPkmQcKjNncUp/QgjdfTJQBVHooMhB+zepBNgYF2hkOxrm3X6kZf
RDrR70wB9d3bzkwq8pLpPViwAhxmsyQ+wUJ0wqPC4GNUnrHoDpjqq7en1hzWeTPB
u8T3UBgQ/bE6fT4Xt87Cx9Sf4gafW0QNX/a4LAt1uImmIM/wXBl8illTlHKxeR5m
Z1lNv6ev8o2SUDHXyuQqamfxmh1eygVvSEjwZy1uzEM3cKFtdod8qf5/qEIX4NoK
ZHO1UUnqUr94lhXM2ZSwNHjewW2dYPwCjT8MnNB39Q0l7DRsvARpw01JZLdgA2fi
DdXtkwch8n2DrbP0NEfgeR855fu0Bk6KtjzjTzHzAPzMa5hSF8ZHA0b8qScXgHKY
rdkGWYrLesl9cb1fN7IJT4n+hqzoAUx3wXmbvSxkYn4V/xzpisoybcpUVhttUi/E
luPh60BELobAlvdqkBsMoSe4bBQ8lZ3lin342f6d08MCkTMREdD3+9YSoocAyU+z
bG2eIgtIcIXYNk/Xor6lYJxX64rSpmovNtv+LJo6HfS3ewz7kxwX1Be3pkOYcGvm
sUOQtIXJB4Wm67NKyKtIq/SEgggEuXFL+hfFuHW8sgoTUt2oBWOqUfjpcWG3oFpW
6gZSaBykEZWfMeZqWGyGP7ZLpAtS0pUcxlw8h2mCXdw0va+0T+w0mk0yWS12q45F
yb1UzKynK94c2M2C1SOvHbpccO760w4OpO5QHU+CgtIg1+Cs8FuHoZ277tzZHy7r
fc0HBFEQYt/hJd/1xaOsi2xnGpjsVZfjELt84yRDmD7gfJ1kNLJifl+fw7DZdNS8
MhRipx1/z4HBmqh3RzdCw3rueys5JabxXwRTk9CIHwgLTcXc/CsMFUq1o/WgAt6Q
RTyIi5K6F1BKEaHQrifmIIO+YmDsycJ2P6cwCxK8VOE8h6/aGTL3vq40i/o/rK5T
cue19Uz3SS5uHb2aFu99mjAXIKuR/Bpo77mwCZftvyuPZFndkv9sw/AC8yS36Lx9
Kk+rINDCCXYeIE+bfodMix1GrnLHb+4RELDiMqsqNFU8E5J2lu5lwaOYcI8G190u
ncvIAb93++bHW9mxHE+fUrmxbWSQfBovsEIFzKhgeBvzPxlV5hbWahLQSeJB1Sa3
+KgMNKgMMWWMu8gIdKPyZ+m4Pv2xaGpJkRlUbJjRGyJWh1N2KOI+JhrMPrS1Lxn0
D4t7ThDniUL89lKRkbXalSliAFqq2ooyBOt7rYppaxsJYLx+TEnbiIfunmrqJNKD
LlJRZ8O+4bhTpJqMDdvwxrbRk+7QJCy+b4GknDFLHOpBiQxLOIvOB8wOHiHfoHdR
gLzyIXngpUpiOwTcZRf7kEQU4HPXQlOL3Ol718oKpfTVDhAXqjLL/9b0xgjOEtMW
Ksfls+gkrS8PBYIkzdptp1T/eYDU3tnUsh7CuvgFD+SWgTdd+caBoi7EZLhQnGvR
uTpdRQDsVZ03O6uftesnGMQgmmo/S0kdJ22LiSNYi3dzdw0M2hnM511RF0V06BMs
uHnOdEDnyZpfQKL5gxmRJ5p1KVU9AK8T//T3GsGCWTd3wPYi9z6KK7Bxj8QNkYur
+/vSkfPXqigpwYywOTsPH72GfS6BTGZ9dWMcrIm07Uw8apWjFNjHFtdIhmEbqNlA
T5MoSwz20QAKAdFwppHRlZcCJvZ1Ynhdr576pnGJ1NLm3/l3N9bEavMmz1Ca04zi
Y08G37Fac/ab75ZH5hTEwjR2apjSMIlRuGcrvNIXJAiTJUNqvCx2WIWW05seXTDU
VPyqXT0bIw03atwmbuvtXELcT8A/fP1LqRUYdkAu1m/Ri2R8KiQfs2O10krO+Oks
7GpLFrL3mw0jR3Ke/zB/Xp88kYTmgJ2WsLbEN1L9Jr/VZHq9IwlgmJIm9vFZ6oZB
Fbgn17B3+RsCG0TihZa0v/7ehKC2OagMqyHqFdwWFy7Tfmc1+X0Kf4rz7/O9bYLO
0TnGNmMQAhJLPVjvPTdxuiYSQRd5RucmNjwPdZ7erKsrp5hWR+OgjFTlBe8Uyqkp
DYoj2jZMGYp1j2rpHpAJh3pEIpNCglpX1yX3Ox9YA49BXRTYVf3JCQ0AcTIlRGlY
25i8moszrCL+Ae24zKKhg9vm3zeqzCLEjDigUGec6cn0TUvcaB8gYnyA3sSs+sDg
i6E9P+J+J/0PmMYQF/B3n0zoQGJrfvSiBsL5m1IOprkTXmP/pChRwcFJqldfSAG5
Nbi73HQ5mfUmHYJLhfKcAMzsexUokAs4RmX70ziO2YkSWWuJR4kLkNg4Dbb5oppR
/wMjL7wuX3iCLvcXvI/bLJWQQQ8seed3TijTFBQpeETX7hHjwB4sOkpC4KOnVTw9
yoyr7tDjEWC/+ccW/e038VqmsQ6nvfzHG7rcBxECOJxrYsX37KWefWSgOa+WGbsz
JTcYkZm8pwhYzbQ+BrF4/Yu8tWjOqJlZfzObZMfS6/gu+48bpICPTroJfMVumzgE
bTp7NZy5RJWmv/edHL679i+uOaFsCzQuDErqlKhpoNVTZww7HYrxs6/cyO4qeEru
8CJ30twdyYDbj1qAqr/k7qYMQgTyuoZUA2by+HQAgAFgMw6iYbcnUah5JfFbFgGx
Wu+H68onWDIBtw4oyACbnGDrbeDheDOswaIsiClNpo+HDqcvofq3BjG+nX9tLWZQ
kxS6Sr/c8Kwv41mwMrmAmatfM0TjVBVUssurYM4LCVt3COKy6PRUr0ncPaaWdv7W
DOcwO212IY/1JrJgkocSPhgM3/eOvgCOkMDTrbk2z6F89vUtydZ0TNmRLK/1VFT7
EFla0sAxbB2pLlQVeA1UZtsK3grVuIu8BfSzuWkaj/hLp8FnaU1wEtv+1JrImSQ7
RQ0BaBxPsl+KeCFhTGuOTGHrTbZ1AkOMjp8/QRYMAoaR9YzIBArM7rZoRPTV6pBS
TMzLLFpUkrLe4ZZwdjqMmKj16anvky0scTlvSBp1t9J3Q/zIgKkAsDth0HQDVaaG
njfMKdep9WM2ggzmPbu8NKHoxTFL7mgJEG6kZGU+6qWl2prWH9MCQPwWBBHmJWkZ
+ZwP6hxMjbDSppAlpDkT3zowHcJXpYd1zDEXE7xv6ufF2DBrk6r/Wff/V2ZsLrwk
qO6/P03iNeRdkw6UDDrSD4SdcPi8I4d9jfglFQIbBovZFQOrUeEsZ4KYgiYNpZDr
64I5DzttYy8jafJwMsS85GVjpFg1wEjXvtJjTaXHYghBTqC79SXybXwXkqbkr+0x
qyS5pGvGLZO/V30bPtuDnVgClcfNcwMP7oyzxP1M2/MwhgkkP3eZ1gim1zysDHEY
3YryzHkSof61jBjL2IzJbV3El8i8adPeWTC6juK7Mz/zNj0Z36pEpt4jsUSX28rW
0OtrALaW3RjHbOdt6+9Qs1xO8qyPZBHV+sdxnJ6GizLm1Pqcvzm816tagsVTWQ/2
7Vtga8BURIWrRnV6JcYtc4fj7oH50u8yJ5I+z91SUJgKk0lVDMJO1VSY7myNQ+Cx
QzoplyXvNmm7VFC2bAWhepIWBN3MMAVM/Sl307wCWVwHpgHMDDd+L7pJ8woGTB9V
TmfRTfTYM8YYc42x3NjYUbyNGBFaVRMos56Ae8Ovaf8qmvcY2+rodMtLgHuV8w0v
lMX8F58s1t+T1dFVB/1ppMmD6y6XVxvV7i/LkebkKxasKeDRhJzgO31l2Ti0lLSR
L5Lmd9Jb1I225MABmsVnYdIcjhObY58Ap3z7WOpSy8/rdh+P5HKAOM0R1pcMdYFX
17AmXS+WTfzh6cf69LU4N+EIgn5f12JSMOfL06oUDGbJN2ltVwPqqL53IWExB7Dv
pAwZOAz/NyNShJ7/FykRFbwUuOfwWZzLneP6KS+imOduvO9YYz6IuAn0Ua0dyN9T
EYddTV8CX2uxhRPWxqEQZj4GMRiIpPv5u8lNpbWBSu4q2o0FdqK9FFJL5vItMyLJ
MHJIrQ5Cq6rpfapuElwe30y5RiWQeOj7rJTQRfRDAybLhYg/gge8txWI0IcNKSui
Gkc3ZdR++D8qqo6bHnRNboygPmww7e+fqVJ5kZpkCY9L8SG5pOftHDi++q5Sd+K3
5IqNPEyMU/lFpSAJAGdsBym/0x3O3IFRkSZDuhj/hDfgD/EsQ/bZfm/am5N4RHRK
5+CLhoaRYPSPGu0CRL49vQYrjKSSPJS/F/ALGKh4igmk7d7jpohtyI8pEWbNJT6e
hFAXMW3dMM8eA+dsFpAi/VUERBJjeSixCyBsIQbsDqhnmK7nvroavVOliU0QkqZA
kfRmScmV3cAR4hkfH8hoJSJUn9uIogaq97MZHtaQmGj//0T5ju0hw0jKO0W2ns3U
nPRhgRWIpT8Ax8kbFzKTQMnSEmjJb7wE1/cYTuUuL87Fvq1tihk5aI9l97UP4nSu
Yf+dyQrfMWv3LBa0r8687X4cEiVNmn1G1V5FDB3DfImnfY19/or/8+z3lakl3GGm
1QgsBCmY8D3fr6HO9NFY7tcYrt/CTQJ1wMOs9P+pyxpxLPh6cpWGmlAUfCpkUPER
u/WRbqywvsLRmpyOmzLjtBFUf1G/+peIHg4rfyxzfRi6/0pziwY7cPUv6NwRhyRL
/Dtlml9kzDSb9kBM+xsOu3xqodn8PAq3WUSBsbP9QE9WENWGtSczwVKX791uSnW1
lLcCyxLnA7Cs3/4Wypsv3QW1dI9GqJRg8pPyYwnkvbaYvAFUndjaJru+5BqkfpM2
DxvnFWRK8kyTDXQpLv0tFTxuhvyBKIRu12BaP1Aw4kjSEosnGW28Mw8JWg9a9Mu2
CKlDhFPOq7LRm76RUT31Go82Kx4V4rrOT5l6MrjihyVEfllzCTwBUGOzcFw7ulon
2ePOPIooelKre/ez12zeFnBZwwa7BD3fW0owrdOs8O7ul9QQDsDELSdkjwZDhKqX
z4IHPRoxfBmETatHKqIhx/CrpY23ouVrpydgG6rKSsfK1ZZzQiKPBY9hJViqv5j+
QxSgtehrJ3EGmdbRkYO7bM64vH0zNDYZGsiW1x52kC5FLO2RM11MZOe9KO+EQhWP
sBHlg/WMCegzw5p6uInDKH6qT5xVp0Y+81sAPLMN+qG4sFmy4FEOfAHSCq6K8uVE
uF4bg8E7KZOIMMfUPsNTFJKm7DxsR9dioB+r7N2/LnOBhexqbbX/Q6DZTF0Q9gkA
OWQykksXJccUVoTB1BHyOzyAejIxudSG4ivCkDHB8oxsUHvZeLpFrpVD/LDVDLdi
8oRFstygkzjdeO+pxGdX5KNOclA4YxUQFC9ErQqwLSpKKar+1j2GYWH1WwfhMwsR
PMQGg6kr8hbSJmRAPf8AhGigM2ajvxW7lgg0hPvxjj1MIYf49wSRnPOHHWEtanNV
Z68ql2g5GPyNs2GQVkC+8+VEvH2ZX/viVd1rVVvJy0u/CehP02+ngp0L+z19eFVg
zrzOLPcsy9ITneuv3mJBNwcE6LwpynzIjXqQ/PhPp5T886/OXSSpXZGmobIg8ikK
mQv2gzInXqS16s1p4DdHX/grhzEQ8rLzfQcZ6seX7Y/YT7AYDt2WZEfs7cYNrFlY
4H6nJp03xIwsBx06QrndQllOTIFDpsb9I7FNDZgfXVx56qiyp2B3S3eYkua8BSl8
kxAAZyj6Rmkl9Wa4INkk11RpmHyORDm9k03DrJBfaiVwRAGpLAPtjFEuiohaSUTY
a45UBNr6pnPHBG0Ygna1NpFV65ylzaBLz6k1nJ2lqzFvCXptg1/Lq1cr+L29jLkb
J6sv1/Io5bQtJPryfHsFLe6rOqsRPZH1NBiJyxtnf/pe5zdexRgQ2mk9mDFTWDD+
QxzPeVW/M0tgmNqm77B6ZW485zHiPpxIoa7W2UE3VORqmDA6Bt8n0ftENgE6RPPB
r7AsGvtc0bLkLY7hj/EXeuKbS/Kdx6dERQKN6EoI5tN75DmpPtYDB94Wdt6UvPvB
ZJJQXOb9sDKptfj6huB+fnXstwGNv7JuYIrTtrKOzvlSty+VqzF5GpjYTTi7ddpZ
Z7aXwsoBiJVr8bZ1EW5WsULQwJ7LxkolsVtl+U5BXQjFEnrK0igmL5/ZMWCREd1f
25Jq/RAKwArznVAAcnFYFOsAYseArP+Y3MKWMABJEsx7HG/SHQ2hro2Dfl+PJYYr
FjaGqDeHM6hLMpQoNZNBp13Sfg9frbH/CZ1/V4Bhri2VtqrA8ZnAvEu9qRXnf2zr
R22GYIceloSWAsTHB3Qbk5dk2V1UhbhlNlSbSu7xYGGm3tFI0lai4rag23jkeAv/
8w2JMgAxxnlqdt+6cVGvp0GVVyypt1m7m+nLUYkEJNbU83smazKVrSS/fcUy4l2C
1TgzeyosXXMteUH+YnOvsORQ3JnAnHJeIoT+Nt5h9r8MQHiSCqoytARfP4RGzdaW
fxpaih0bDC1enOvQ3B6mWKaSH0KuGnDVi6j8MCJjArXkEdFrJA9T/+6b7PfLkzQd
47kTHoA531NsyRMgv/kCBWPk486XdcdAEXee7XmWjzsjzwIBCOGYyY0qrP8uS/gY
AZFqhI3XgpLYbz2B4G5lq+HTn3RklOIPN7kjRbIJL1GpC68rc26zYdXHtgQo3COE
1IHR0SGqXDdyDVCB77yc0D5Idfd5PmYI3kRadUjtzoW/VPC3Uw11DWszsAjuyPiB
uC52fs2XzzqkYYcYtE1CW+6KB9Q5xkbG09LWsOpP62vuViqoMfJZEyE8ZkZepUx9
wQQ/pdAP1ZpSYjiureBLEjSRR01I0eOZMyJXPERNy718R4c+Z++35JYNBQdURrK1
I0vpCygs2EnLyfcXo43AdCxiQouPduDRWQ+kkpC6NXyeerZorgTFtKFAbOGie/lF
6cIMmKWdQcj9hSl0Q0Iyxe20wGFt8OTbDPMCOmCqeHtyYWddmEMn9ZiuhZLXPhgc
caQIon4ODBbdvFWsDio7cC/UIEP1iq8ESwNDSKRPWEyWw7r8wWAG4sYXEkMlvX/3
vJAlMoacvoxgFDDrB3MiRUYnkddVWg+W87A7eJU20hyBZUcPvWcWXq7B3OPX5ABO
VoO2Z3zTL3kYhMKGWhnk7ewqgSdlIWEHcvZAaM3WeRpKMbyTMHWRgq/Od9Llrr1S
gBJcT8UwfRRcNCAhxvEQmuL2Jeeki9tVZRbnGPggY79kUOCeg2l5zPwKxZeWk4IK
9CcIrBEuyDvZJCcF+XDuePpiy9P8FhX1CKZtMMzwgQMtZ3HU1rzeehWuV9Ddyl8e
INWeQsSy6qaeOaRqtpxLvHAzz2KhpPdq6kACeAXM49WkEyIQRMaf4ZpDMoZcEtcv
YZfxeQ5wNbY8KuGFw8gNSP+G+BXOErYiAnxdfNKHPGjUxcyTQ4H0RX+Ghdl48FXu
3r395tNHNFrnOfsPCYCgKSYkPPxY7a8oNKqMU53DYUXHybr2xv2Y3We0pGnXA2zM
xH2l/UCKgFzvydebP2Ppk0OfBYQ2MHhfvoUmJcMRDWsaRANmzX+im0qhAfZo7GdH
GHPF45E2vHMNOJaD1g1qU0TMNxMbW1IkTbq2/e7SoV4fSvrh2QoYJGjRz2L9UGBQ
m775Ln8y4+YNxYNyC5grLf91vofPm8ZcxGxj0hyuWlBD86qgYv9YeqV90hx+LY0d
StRxVdNDhuqlRIhaQjabOSxPrzToqHPxQw9oZ1gvXZtRN+WNIr19ptjS17GLXTaM
qY5ALlO7XYawmhIgattA7FipJNRMUlCo6GSaS+BCudmMTvglRoLp8rqYMtobz/QS
o/XljzvJascAl+WQ5VGJrLBYOze/zfFkxCF5ITewINImuBQLXg6hAGrQLEcKnnop
z78yh/uJG3rk9yIqmd2qMR4aVH0bK7m3voG65OrFDjBNhnXNDrKEvD0ebVqlNEWW
VEhYja2a0nOjNg8NxMyOTOGmVSK3IDJ204k8ARo38EQ6AsQhrPdyyu2ZTTzVb9GZ
GDxItAps2617LOMwpCAa756aynLIF0acZbyGtAjiNqR9lHF3Z+6ZY+v0tBCNYHTb
2ZdvYRYHdpsiviLg2cVOWKEfRzpJ6mu60E0bR+ebddCxspHkhnxPLk/vOVv/Tku8
ff4diG94kRvh7UjUvpFl2kVnZDTw+wjyTCUXETWtsijmyafKHu4/WABPnWwkL0IX
sidQ9UxMM22DyiwH7ytcxAnn0t+fqjpwNXO6byhYcto05A6tHHfwCC9UrvGjjnbU
G+gZbelTOKndkjLxyF06/cZHywLsz19QP03QD000mJ3IUrVadfErVeGL82Aq8NKZ
Nf8TSVl6KIjbX1mAf3EDm1WFvxpdU2pmq8etzqYhLKJuYKssjqHc9C76EN8VJQzZ
87AI+Ci8F3qwKrmoh0rNaZhOZ4on0Phpplf4YMGZ6KyhvVgUCNsY7RyUuXHphSLU
9780lR7ayVfTCSXYX1oDs/WEAGXheruBqRay+n0bRtz6jWT583/SF/B/VBaz5STq
aTUGvSD/hreFna0Z3/ayL6AhF+OdQ29d7zVtifQzPt4Z2Q+D9XERYj9EPsWyOoFk
Dy5IJvXTl8lDOUysVMHZcK88EHVVtUs9diJKJkN6JlgyDlAjU+bAeu0hdzm0A/B2
3MHeGRnUCtnFXbhg4F5VTidqViTykGURY1q5XlS4fvJnD0G25BFZJKMWV/e3a8sd
2q2rJL0O9Nw3xp0w6oWD8nm6SAjoO1xw/YC0WxS9iToyb2VplEewmxrdpartZL82
DHQtPkfqRJlyg8B4yPz6Kz6L0LWbb8nwZ7nP40nodfRGMK62TdNvPxtgwesF46su
9YzB73NjdWvxh97mEKmbuNipBIeGUV4g7+DqWZcCBnfFaO5unNqy6GUGBC7cSDiP
FGWx/H7n13YcCoc6dgEpSd9uvsHuNUNElpui4ezPgcMTtGFlAg9NGN/YSejF8xrS
e5uyHq9R5kgrVNzPIhuWQwrGbTa0Mz1KIS1jdhDTWd/08yLGRf2NX4lBGeJ638P0
v5AOSW/C2LmvXyQA+WarhvOq1Uv5TFndI2bEWpHo1eO6Mhk43FQ690zOIcBuSfzk
Ch0UwK972lFwWGmumzyiGlU7vrcyHxeBTTu5HuubuXEbSh3wCvAyfoh/p0IA5CNz
C4wXoXtpzlQMob64b/ALbPfMWjnzi7fCquLSZr/x5fkpZkJMg3Uruh2s+7jh+Vhq
8rkajGsURJt+FTZBgIaZBb998ILB5ElJuAigRgvsf5DIbNJSw/v93b29Kx0/yM4+
BZmCdNkLczaZixZgm43OYHIHLsASetXYeyDma8NcYzxd1QJKSvQfgfcuvUt0k6u3
IgPg8sNKEyY5K83uwcNOb2Ssb5XyDO9LnhLqh9pgoo607vxWcdjs5qHv2ISzSF8v
1NFR41Nt0A5pyno8OncbIlvFCXQAX0eBgw2/GEtynCo1fhGgS15QuDoOFfqtTfWg
VgFcoB0eFssEpF9J4FEf56WOvoUURwX4NNsUA6vkjobm4QyXT7TwkNEhSBFGailS
dk9FxJeHSFCpvLuE6T7zOTX3eah2mbSnEYEWtfkLyVAdXVqYb8DychyU7SW/03T3
3jdXcdCoRO69m0OlW8jwdbvTvx10rDKg48Ipg2xcgG8crkjreQJZJ8Wo98uJB72k
HvB2H2t9dWcxiXaPboDeKynS0x9cKsjz6MBfHO6ak+Rm+RjJAks2T7oe+RlGqhuJ
CoEsTT9fEXYszKQ5kyMZBkpLGX9KVesB6GBNxS5x0n0fpaNCklqwLWhTLNhrsYc3
lAz9Tv6F3hKXWIW0LNYVnC4gPHtdNxIOZBWsWXsU9SKo7viBRhUzFeDyE5Kmztw8
eFCL8G5dJg0aLWDGvt1VVcb2YjZprG+br281eWl9NjTDco1enCjST6aLZWBBnbe9
myjQV1L9lbs2RCXR0POgu77BWQ3cvhSeWjPsxiwXhob9lMDOlRbYE43U1P9niZ19
FrNUXbBUT9UCc/zD4KmDbAZ+cpgiKbTOPCXhzxMdqd/HKxlQF962jztqz7QnGLkU
0rgXzaXZ32Osfmb3giyWDZuEXOndjuoKe1r2oAgaYgVtbXiQrdPo9qfBGSIr+SrA
4NLhm0IUUxvjqSUt5QMOuEH9og38XsuLv/zv/oLuFr8DDnlopd23Qh7W6FtyvFRi
V4BhpBlbqZaCe3XxPLO7LuFs3FhfSwSq9Sh9uVz8Y6u8Qz0pSerf2SDUqgwhnjfm
ECEjCR1kEep+TgVedseukM/FP39p3NbliK1VaL0S5xYYWTjg1nlRzkudHkdFstcg
qzeROn57uNBmnQghOxZ1M4wYd3JTkmvqS23pdvHDlGqJquN/lp4ZPAHFmhCGUKUO
zF4fba42zmAdlzpZTgvC439FJwfuVWRAMdQ5glftNQUQY/wgg6ndseuoIv76QMwH
Dy9N49niiCWVTHBTaOHax/kO2muxBli1A/mFLC+7XV/Daw2XY0hIDkDj1KfxTrHy
xKq5gtex1U+wEhWA6e/PgomBoqCwCUuGgA2zoe/KJEts4I9pkEG9fXCfYH45IrWM
lIDbVvIW+pBHlNDARqfyOVxPTHLpz+qll6KTi1qVw3qdr+ySMNEVPG1AubqAuL7E
fgYZzU/oqq8IBl2nhtqAZIuwZDghGoNALy2XPeR6QQEffjy52to1zslZaVe6116E
8TRk0I/8OyooH9vA62Jawk2mBSVG1cu0LfIgPx4Bi58lC7/kxUMoUAzJWzbzrQVy
QukA2VbI5gwg8ZD8ulmSyj0lADRJY+gzMXLIbYs0L40ceBFB2eQ5vwpAZlLyfDq+
jTp3aUo+Enr5p4Jzw5BZAJcYB0iIBo4CJkjnOur7FCiHK86ejJymGdQ0DDriOoly
0LyT5qf889/eA/tPjkNOUmaztsUWylIUlW1XzrOMnDx9MeaQf2Bb8llWz5nkxnnB
Z6LvuGqBUpeHF7BcDaiOFXs4872YTekOxww1gGBfCgsQQB53ZJSo4DGU1S5gGjvQ
67kvlN2b2mqWw7tnJhThH69uaplpKYSxryyEi8Lsp6lB2l2bJjdwDzgfNIDgxrTl
OvpxT8XiiYZymQuI1gz5sqocCNCSOEG8OwxCygCOTslgxBb11DjkOKT4d9QQQ4I1
2ek/XRcZqUjWYzt3wk68+RmLjbpzgDr8vWrhNjwB6oquwie4uS3rntabezPguGgn
6nh//EcejQiLP4Uemn3DzkWB0k7NWb64NsOtaNOo+2QbLL/oQlF8xtSxOpK+6CCn
V6El3FwldOGf3cb5Q/Ss5wl1kCYDokncX1Iek4qwMCD091RBsDeYVojI0iRtiHXH
qml0ppYenquCGxpVrsyoN5otnq3OJ1G3LYtHcTPKPp9Q5SThsmNRqjUv7MKYKUFr
Oqd9s3Rm4EIfxEUnPR0OSWcYb6jyX63obeJE7bQtFX9MzYM7W7Dod2hy2nCWRJxC
IMF7Z6PnqB6LlSFvwVcOz3FYRWz0epl0xNSv9t5PAfSYLXjbqF+s1YednXb4r2cF
90H+l6zd4lcNOIDknEgnpSrZAfbAAyaYxEwayqwmi+oKLpG0UajoIvAxsYakA9+n
7aThsqBgB/o7CepgdmeuT5PbDQX8MLYpl2Iwif12cumrjEB7gX49/D7wq8RtQNWp
hytZoarxFlTGT54Hdo4rM1rr+AisTdoDbfqh9Ci3En5jcbUXiEcfTfj3KuTv6Zfk
BQZieUBCNG2wpEAVtzyZypgoXgy9oJaffEW76lqeg/qtcrFz8rvph2pmmyEKjHCA
NozZIyjQjEZ96vcyu5Vkvq46mfS/lIZ7vOAT5AKS1I85sthlcADbxDSZhJVz+PC9
eVg9o25AmTy1XnyVXWv97NaG+O5s8d5Ki3wpDd2xWpjcY15GrPf74pKtrJRV4ZAX
/Eqa4LsZyupFXJa/CEq6uQ6TW+9z9INbDZ3H/I2eBLJdm+LK4v/dbiPlBD0iuSoJ
vf2QyYO4PqyghPY8IoUTvXuNGG02YDktDO/snbr12qOjJJrZHyQoGswqx/l56qN5
sM2+LfG6L3v/Ksa7mPuckyTgIdAvQMcsiUuxOmwtBdGhxfyUxXyEBIUyXDtq75t/
AxvqHzc8SPqrAN/4aITDX8XcgeKGZ8RKrN7IKQU8uNWYc3wJAukMJ3gnjUW6Qhlb
ifaPVHZgFwwX2oYbvaatvfi7fT0R1uwmUZDgbFk5C0d+9RSmEjYPYJ3mftkX13kx
MqzPU7tIDXTvYIHw5wHHD1S9Nx/sOn3ty49cAzmha9nftHxp85xPaXj7WGY8iVfP
iKarT2eOsmMuJgsJ5DOSeoQiEiynGxV4sAHtmTFyupF1pdvkU2XNdZxj2HlsE7YX
NdPp9JEMNNIMLXR+xAR6HPPTOZBij7wxtDNKlmcOPA75/pGsHDj5NhIUrft/4qTG
pnn7ybqOouUt3TrpruFtbvEd+6dW3Zk07YG0SIEFQFfaTypUeHnHqSun4gyxxfrx
XVULZ33Zz7/bIxTdyJjPrx8xZKlEG20fg/4tdyLLQGRtUtlnLa78eJztvQ4UM5bE
lp10qSLyCbecqr7g1tM76xptpyM5sE+AD0MwdeqH8aUDdZGF/eoFb/4C1kgJIcO1
N/5UewDtVLgCQ59dTcl1QY8zy96Yzih6JJms1uBKOSn9aTPVGzv841U3MWn6XY1I
0LV/Xv/obtMvEs4VJiwlvBqWh6mG4IiDtwIkEMvMIDV38ZnkBeLftxZiQaBfc7sl
KTlAgmioyhK+EUIl6mpDDNxJK8Y6+5cxWmAHKd8QMqP78GAfhgaF/C/m74873gF+
nNYgPjLL5k2AYQRqLTRIxDsqCUFG/vfXvJqTKKZy9+97vZ5JHnOAV/Eez8JEnBGJ
qaMD02+ZjwGah+WtZb0r2owadZJBDCHln2t16SetD54cPnXrIuLcaa1R/hdTx83q
x4D14THdlANQtwmZB7IF0AXMRlArEMq/YmfE1ZUw2st0YDF12pU1PXF/igwJugAi
grg6sYcBDfBjKrzq75/Ec1AjddyqPfiloLe6m0PAl2wT4cCEL47HoDVYMx8ds52C
LP27PePqLZed8HGYEbVOz+OAcY0oeJeR1q0kcTQwC+w687mkKMYDJeOM21D59ipO
S3WHNVkTYMo4BrgEHLllBBEQ2Bi4QHj5gPmd72Crs6nC80jBWLyubuy7pRbMKBAR
1kbJJEd0KRXkM4Kp1JF0jsfQFYZDUR4sNHxCbGe+2noA/eWfOk+lz2pjfhpjtWYV
STxXCliRdImFaTP9uGDynXOAMjq2kSjxQku222eZwWV7zbqsvbM8aoo5RcTsimph
1By0NvIDOVnUzm4UhisPPEBQZOOaoOe0c64wNBNQmJqxGcaEbX0WIBAEFl9kk1eO
pqFnLgGIBdj85yDczNK9oejy4ZJR2Xy40iho1Qwn4H0A1jujxoEDy460+wsbhbcX
i+ZSArKNMLQdU5GuGbXw9UOsXmtYsHPwlWWBXWp3Ib+TdXygLXSZI+3g6CqhfIjc
MTIe7atqLX9OSwUvp8m9a/fBj4oQosuM7hsNE+63pKhgO90xBCQ2YdP7QGDZ9HDS
FZ28l5VW2iDzbtrxElsvNaisaXCjqOBaHOg9UtX6ZD0orQp+1rsGU9haI6rMv5k2
G7laptR01JSU5XR/NgIx9Kx4dc7Q+iBrUp/OUh8iDo613qsQxoppjsPqJPa5ugtB
ylNi0Qqw6uu95FGCiHXQPNkwnLu8ubvGWvoUEzvwQxk978zugCWULhqTrRSEvQ6M
suUb6Wk3L+n9DxGMluzuokx2ySbLttHHKQ0sOozJg4bBgb37urVT0dP8zPR+Deb+
SYg8hYRSAWjL/QLpX8suvpjU6llnegXD2YmMcBRuuZBKWsvo2hRwqgLQUEQxGw2L
RbHa8CcCC8meJRIvS5pJXuXeMunMcJg0U+pwSTZAT88I3sx4+jBlW8waZaf8nKzJ
uHx2vxM2/f1aMiqlctJUQcZAcZwVNrCxYmu56u8JpVzXuEs2tlYI96taPv3cD/8Z
802u+/aHHgbSpjWoibDWAqYM/6Vpf64KlgeTG4PYsNpnegPLl356/3mrXpBrlhIB
/zSRucAYOjiD1tJVl18YDC3PtR0zNmtpm1VNUqo3DDkS/b1AxjB2Szsdgq+N1YOB
tPRZ7l3Ifel9MxmAkAwuVjpN7lazvT8onDByenCNvOPrCfhZ2zSMyHFn7btf3Fth
4BVOAf6nDjvSuc1U4iz96HzeIREoE2E97u3zFOBQasAmqANNPE9oyf9Lc0kAt9JA
PpVxyFwrh6JejdnqoH5mcIYrhVyY/vyKFxf0hKaWyaqrALwEJR+gaGStA/VG6XsY
KfiD7IiVxrYO5pqjHR0Gr3axyuPgxWJt7OAx0JQNYKhtJ6b5MlSxiijSuVUQ1Bfh
buyW+VMB7SCOuLD2nXu/UE9fBQvyrapqWVZmKVkwnEH2KfkkNQcPsu8MtFZUTXaH
Vcd+/sjZGoeql+U5ouZ/bPjKiu12ALXqz+Z1YGCMdsETqNoUjIz1AVhZQX1U7l5b
hSZ3hD3UeYKrkJYMh2AyXknfM3qTcmg3uQKZF9SmBws9gxaU8OPRV1m/TWCw+otU
ydKxhQi8zTnMpWVhSFBDFcQtFXpLtfnKHrIcw0lQV11voQzJtIO82Vu1DJfBPLb7
KI4KAPlhvHbOEjjx3P8Z9sfe7lM6OC8kkq86yAnjWhV8yADTQi/5S76apVqag37Y
WYp9iqEvnGMag5yZXOwIQ0l9I0mMjSJxaqi+FwcA/CjIybA15+eLifBgXDZs0KR9
+qB/Yra0G8woBtrAdXoc0zNjkV+IZvHCqNCbYfcfIZwGXayE6RdhFGmXH+9PDvqX
E2bPkEvRMMq00CcJASyP3o0SvzAiVRUJE4gGZxF1pkh0g3nD1t5ZGkEo4LKQjTbX
jsVGeGaTWBgBtGM89QSCz3/q3RDSTC4S7+AIAzcnkfb15IhxZ4uIqxIQdoXNm2LN
3J4VIFvhDVl7W7WPaKa1Y1QXP+qO60Y0KanirsltvD/3TFkTP6vqULAVjMUwgYya
jeQVBUv9O9ONnSxGFVeJ1dWUtPwz+qIC7/vT8S3FyJKk3rS6X2af11+SRT1DWzy2
X1e6Q47+1V6AI81vks3BUQ6BdjKSx+f8T/E4IeLTpn77Z1lmnhU9MPYm24Dv6/3K
r26ZVXKxBevMML243QTxY5PeuMOOSQ869QafYhne5OfkkZOz07Td52MgaVSDhUqm
Y99nvhiCUU5NsyUbI2Y99nBQh5E/1vg9mKjLhLzgWc15WIMe29X3CBIIRRf+UuWG
YyoPJEOtS2Vn+7Y/XRffPSgU7LiHB5ZV+UFw2ckuTQR3yLSluUE+4E4QoyXzLf3h
yCNkNNwJvcpipcvubsaHEBJ+qvU+qI10GURyAmck40JMOUp1SPHBe9JO00BL/xPk
+QQTvK85rWXIbPnZq4q/vFsa6KYa5JIcpDx5BO5KyTZbkBkdMUTVSktg3b6cg2r/
WwtLAPQdJYTRnr4uD6yrioLPY+nD9AY0oyjFuvvXEM5PtRxiOAGcTC8VBDkTbyS4
Jk1DHTyT5Pnb5eR77PmlBB5G5Y+MBD02O0pTihbpboM/DLanol226qU1fcjmsgtP
3b++9tPyF066dhrTMKFh6PSueZ18/G7vlQuwLi6FNtWDLBTE8zICiKQyTvpXWGDp
jSm0F3Fz2tOra3tu3pLHch0GD2dqsYIEJsEFDxywliwZHohLjdrgWEsonZHaQAmC
mxmB2QVFTNT4ZcCqNXPJ2tilEo1vYlj3/YRr8WSP6vPeasea3fJc5aAr/Zfb89lK
Mq/xvN6yfrMm0nkR5BEJNkhmRj4FuaGebMEUOreDLHLm7R5PD9bo0a2zkuY9EMal
8RY/+B2a0MVhIyR1EXXu4atKw86ilc84S142QPcfZhnT+o8AaVGPJhtwZbFLUd51
BB/RxEeGPjsO+RR1yuA7IqUj4nU12QmorhM88KhnGF9Rxa4BkxSrXaMJxXYDrxd4
jF+U6/BrRUCbWVcoHb3ZFmElosMRCCMTeQ09wC/d53g9ZnZPxATDw0qyZCH9ldB3
cnD76dIGq9hiDRJXUP5wx6LVJqZe6AVs/Soi3IDinHy7YbbrRJOUWnI4gEk5b7b7
nykRjiOPjAHRmR+bOO20Av4fGUhtZpTPGRtbsh3ixn2GTrdivEmX7YJ1gg6OjLzF
SUm6pjyTsWF8bzs60RtouWpB/XrDLcwy8R8fHtS5U3Dn34NeGKIuqQGzoAQGZiv7
XTBnlz7jhBiAi296rJ4SLoBP1lI3f5E3WUa9iBKbRBkCtLgD8REJmKDOFdSB4YlP
K6V85fN4TjbpU4T9EMPKAWP6juX705pHYCvDOyaGuYWeeO5qxEjs8SGUEhxO+INA
NLmfVVLu4TBJ/bopbOUQcRduYLrA8hmNklVlJJs35O6+a+xTIhD0Ahutwfk+Zuhi
/50sEiB9KnU3LkNB80FX1pvLjP9cYB0hTQKqTSc16YbHa+FCjU2TM5ZUf9V8jsaT
WhvDHlqBNABQoUKLmkSIIJCZoZOp2BHb9T8OGxK8muBt+cvllkgsRrXb6L6QIo6o
utULKBm8PxRe+fNkhdeXtVb3r6nS+tz+U3BCvmKDl4g6iW+dLqMS/qG+/HYXtYfq
IftqMkF39Rcb1NUKwAU1jyz2xMN+beP4kGGIkbxyWtLmZO1w/cuya54M7JdqhP6J
8voP/Jb/mqCpAzfMR5JiY4+8Oj18iqIaH3InjjiEZcCCekknvVwdGKWVhMH+YBEu
Aaix67k0+SUlCu+X16y9S+KCWR12n2Cxhm104ql7w++qY1Vy3qF1lm0dtQzayk1x
wETyuycgd4jHxcIAcGJsXPGk9lN8WQ10XOspS5ec6jpo1kkvWpP/YuHUYDR1V1AJ
CwTMiwBiiGz5x3BLRInBGs+mLn6fkpN82+yD+NKbrheMZOJMXAhdXwMQBU0xJGL2
jaIE7jEel+Daj7dvqVQjGH6VHA828hAQ+cpV4/77s8ildc0Zu8cdLinCN0G/nhIs
ird/KMh84gpBhnQ/2kQfGxffcbdAVgUey+jUjkSyTAuG8hUuMOVumR5jDXnmydtf
4a9lATH2PBAFWBEeKW+JSpfAqOTi33wSTUSYlz5BYfwb+02athBqkrq6MXyHOeDn
lCyugpR9v+TcwD0e0mDnowJzAWhZM9ITsYmm7oAhqG/VmNdEPoQOBYLLwZpsYk9J
ubysGU4mdlcRmeeS8T9TrA5hUrICOIQaToQI5RMHTvb0ANbGQ40fxwix39VyXycl
90KWYfLk7E35PXIajjJBf/28T1v6VMT6ek46lqNyupGxGnHFFqsltRk9JWq/Ymlm
Kgf/SO53F+xW4ygB9FRAYkySBtFjWw1zVw47MegTQGa2VgAfdhSXryN69XJ06sJB
mdR8tVHnMYf0Vj2ymp21iOKxteLdHIPI+yNxpgyH+aqFmCVyLtkmYs1xtjoF+Pjv
c6vLgpanL7/ZsSSr1eFWYi57lvGa6sD5WaJXOZxe8MI0gWryph1hCJoz0yUiNcIn
zAeUBumg61eYCvMh4Adims6qiCauBhCIbD1ci0JJknFyAF6BpXdcgB5smb+TF6sn
xLlcFa2ZZHJG4LPerMZzvT4RJj9ckzT9ik2alStNNIaNFFB5gwLZmxjGF37rqFNi
9DQh+Prc3kJ2HfnlXBImrkCmaDBNdGvHUKq12nJlajin4Nn/qeOjf7BlvFwAKIF4
UCmBzMBBPaUBFplMYD9GTFibR7zxOY+PBLnuAubYywc8FQq8bvq60bB1FDLEqCkp
y7GW2IWHfoJhfTLmoX4L/oxgz1aRiWQXWyfITgsDDBg2akR8g6jBHOUlSBreRLeq
pBiqANvdkcS+bQU3LuG3Ipp3ejvoXy/CEOiO3+ryNaHSf51lDbiwYyqGwlis5z7F
V4MMUc3Sct7C7f2XKtSEVDbSOt/Y8m9JXTcYXkuGDhb6NNAWGkNvy+ZTz4L1bMlI
GJimuWpfKA6a9OIaf/60NZHw8eM/Llg0RZoLNwSL9hY1cXxobCbVymrrWTSn9qF0
l0TX8JzHq4Ps4KSC0U8LWJMzte1/pjBpn6mypsj0dOq2kqCySjS95vlwifTn/HAi
fJcosIMxy5RPQwTQ+yBNM4+17GDvbFPsqFguB4nNSugy4koRVs4GXOIT0QZDcw2E
zmr9Y4v6j3Mo8cCeq1ab5HM8amB32wDNt/GGdsX+UnWVPKn3VDlikLZ8MHEOXaLP
OcXgqQWma+FjckTEWRkx3cCuIxi7v4xHVmxWKxx1haykT+u+2n7cSEhfjLNNnhIi
5fqSrwhw6eyG+RYObaJkxvAf+T4pwoh7Oid2jaRlQ9UVx7Oqh/0Qm8EK3zp/zhfT
ETcor0T2EtDTg6Yo0ZgmyH4hNiVWRlOMuxkpzo+Xoe8fxQf9paARcPNvvf54Tvda
jakQXFyAcbUTv5cxaJ4pzF9hjx921dhEoznG2GvhmRvjb6hH7+0xgjrnpjYbvtRO
6PQGhRY0OGiGEtNnoEfT4IFCzGvTyji4dww9w4hYWRvRp11a7g2bO4t/HvMW0w0d
0hzOgA03CwIm9jBTFIBUi89IQTFKjLbE+mwZSjhu/UsXJiXmNDrPD9lJxcwdOm5P
xASaRoJfNOAYFPCuhAT00AP0GfkQrWO/y6CEduT8NLObOJLGZXacX6ko+MNfwGpv
NvooM+3zuzL/R2JVWknCDAi9oGZ83TR/GkzJ93nHoSlQXKcwh9thcde9UM+LYBxV
AqxwPT9fCPvP9Yn8299NeLvTiesXfTW6Bqc6OkUzSECOg9GKm1EXc0pYthfktDnj
1JK63D/ZG688a8N82ph3xKG9tTWTUD6X3rVC9sRwJ4D5cAFbVp0sPU0j0xxY9rab
HjMEnVuvye6E6WmTuUPyme71Xj1fKxlWp3xxumwtQZ9kYPcZE2uXJI9507V+OSxY
hDHBz2Wlvn7i1bzTprzl9oJ59sYu/a1ONxicQTSmTzPYD2l6bR+LDWvCOT4Pa3ga
LiDAY4SV2I8KOep+I9Rmo47lxgKbgB6ezABl8ykuGc1EuuMqFJxVVoAJ4CS6C3VP
cQ099i+sr8dl/adAKUFtGp1lFjyPad9QdSfKcCgefd8vtVLqLz44kXoBw3QgLuOT
zLlghyVWbLWBmQskVnTxqcDnth7ARg0Z+CxWdngZefT9160LhOvQLwy3xzOmrb2O
7R8JUeTWm7zrHGKoK9gQxG6I11C6l/QzPl8qXnj2t10ZXfj3ZdmGceiLbuKN7X4A
c3M3+0VpylLtqjqRGDWmejONqIdoAzpceZxFj3syn6+W2vJxg46DcpeHhPkl7on4
rC8kN7gj+WMJZE3Culs4O4SXe8ncxzoTp0YsrETti9NXYEiW36iTuP5qQZ8VPREr
h4S8GAnMSL7DpNXY+qyPlSXiwsAkSeJkNXsaNV5Aa7Ct5kqs3wemPAA/MhqImUji
K/Z9OjDVWGcjWm9fUb09lz/i6Zt56IQNzRfv2xF4UncbLlWqznsdRjJhZ1RowIol
0YrUYiyXlf3nZR9+OxoOZHWVZ2fMLTgHPxDZFKKOJ4g4kYPmLwi+LKPVHoLdHiw3
cTNnIa9QddyFFSyJS0pPSHJ7a2wZI+cQ6CREIw+QFscdmLtA6H9FyXnyy2YwJxRc
sZ/ZF9Mbr9YUADg87rWiDCy6GxdIFUFQEbPdfjLRFBY0AG40WAfza2+WVF59atbr
aBu6k7kjxiNpk2NmgLKtW3uxaZdFJqrDCAjkFq8UwUCqDcABUsg4hd/QcbKQv/KT
HERAU4DljjFYdMlaBMP43O+Sre0rdyPmwYXypQYOOEFMuHKzrkaGboSjhRP2zVuo
1k7kPbXzP436ECCXPHKRNdCWFG7RHlkXkTX6HHHwN8TaS+3/g9wVzTAaTeMGuqrr
B3+Z/RYbEvf5n+pkaj8vpKs/d+kMcwKizS05VArH6ekGqBagewQQWwi8bgm+Grv5
KmhFKThdoD3/rWpaRbecp/odPKaUK9AVLr9tGohN60Iz7lUAxEaUAtxPIjk0NoHJ
RN8fNweVKBykF+x6UacksG2bJ4bBSl1qoarmTeCB+aePtmbB6B4B3asuwQv7oLNx
AfdqTvVN05haf+s8qYW+jgoQcIMUyE/UDllvPEb8O9LNOC8Zhh5J0cmlaHcCmEDg
mp87YHteu3hw0kAemMiN38LpdHk92KgnHLKeUJYSCLYXaKGET87H3bb09GyWyT6V
lmAkYVwZkdGG8iDJsan+h+5hRojauOQK6X1GnVas3PKphhD0W4X3vqlut9yxz6u0
7YhUu+5MeWy5r0j0gvEuDWES/w1SBEq5we/T50+MI4d2KXS01gCMywDbRrAuDOIJ
QRDazLM3G62JhAX1A83JAPXUlN/Y8VlgJqjVOxEKvj5GHx0NXRTlmW5r3aIb+yeW
H2dme5xP/YEi0MRVONqg+O7G/1bdK4H4xfF4sXOcS0gLkjLcnjFIMnwBCn7MSPrD
f4ycuSTmZUySZZcQIe+PX9nZc8g5heWFdINspcs5mxOwUH8IUW6DAh1EtRGgYqke
qY+klVdEj2yVtndaJUZZe+VyM3m0k75Wg4AUWtVQA0AwwZUzY28IqDVXkLavtaIS
WPdipuDJouP6h6OTInBNzA+SLKdA+/AVDPp6sMXyxUhDCk1epzQjRKwE7phtWMLg
8G8QZPSOQ7KojJ9WTSroSKcjvHrAka4nsI2WNgkbY+FIaFPO3/tXArRDf75IsAJY
SLXINj5D7tSy4K/2YdxlI0PLPt6Z1YVk2Ja8Px74LnM1kEwkIYWZbkqCs2l4YB6x
QnyV5nLmqVrZ3mJugpcIune8baarufMBigtZkCFxTmStjcGB9LOcnxHiZaJRJ5xg
o1tvhPQHJ++15ilkShYxzNcJQrmE8487zCo44L+WfstFxmHlS7wzFp57NhoLx8Do
3plLp4ZGqTWr5mok0FLSmFxMxCUqHLkyz+lDnD9HkCJYICIpApde8u+T4jlUvjqf
deR0VclCYsyY88rnoG6EwdV7aPRDtTOK0uJYHhTSoATuVptTkBkZz4i+pghuY0L3
wZX2usu3MfwNSwr7rDlT5LjjwUbqiLxANl/o+a9BxrTgjL1HWCi/HW6gsGdSX1EQ
dFkKsXkDXywuXBH5bcNqCcCw/iVNBJBq36CLLAd7AOeSLizKvm6VrGL93Ro/pWVU
VRGWwiY9yvCNGewISYIIpvkZbEwqlvrmiqg9XED5fdw355oodST8mXIlHYPXJqpr
oTtT0d6IVgLfdZRt4xLge8SPHLdVq2OcO3TdwWoX+8xcpQFpyaSMwa6SA8RCfw4p
sFPowV1amvaUzsXXkgBruOhmfnoKwGUDiKMLzrsxaTMPYjPA30VoDWvMEj9JmVRs
13rXcPSATY+UJ1MmRDcYYF68q9EgEC3LfGalirTSOLGJJ55d6WEJClMBmDWvhJ95
EM2MLblj+CrkVg05dcy2/lMM+PP8NpEkusqEDI8I6XF4EeWBd/qho1yIe77um8Vs
rzpBcBHdEU140ndXjn+4sh4qxrruj/xYI1FIxv9UBiDhiufBs/WhYiZbWxMomJ9S
n/uhx+GrUWraHasV2dylAkwtq2PZEALAKWjozAIgjoQmitliv3P3FFVfL7JexBEL
om8p/H3iu2bJ1zQFbVWg4tga9CUa3nSS+0KrYTtW4yVgzvesjGvl1wZs9n05QGn7
WaBl+TLhuxjBkEF4eTZlh/MEvFkeEk9YSSjLlftfUCni0a3O/SFuTYbBf02Fvn+5
wp55pjmLTiOcJ1xeO+EvpJ+2mLM46MBw1ff6CJlwbZs5aimF/GdewVlYvrja24P4
Zb9zSYcrG6Rr2wfqfRxMzHyIQTrAjkB4PC2Asu1qSkwC89luKQtH8OTWFMcTIwcZ
TLx7SXJnl/O9J0kVh0B6/VtieGLz6qZr2N/znyS6EsM3+33HEwiozRaRoevT09az
WqdXbheEue9KnRdziEN7pHSObr2xmbOyItsOTLXiYI+up7NL3Y1Jb+ZnvdJ0HrlK
Z0MI6HrnTKTu3Znykqzt8+O2IqS5HLWafIzXhcvpR3vUYMoxiBUNm2TuVWJsUSIR
Wa0W+u5Uyea+OYc4sED444M0yQhwkjP/guK4YOixOtA3aPyPKeTT8N0TE35ePegQ
SXAJhOclNDl8+q5nAXudwvuGSmcZLIGoFlIjB8e9l5tkKegDrr+Qtpbwa7AWCqWG
ZX+OLEfM+WZkMywhQIgJN/DE9+MdRM563hCc+rPfQSBDdjuXIWpZfhnI0pWCuKi/
enA5s4ovu0C7pRBV4RjuP4rzYkxJoA4h+gEHyqzmVYzD+pTu7Nd/v/jpsptXIzGc
xUZ6Y6pYJJz7vdgdWDh9gw/LsSvwJnE9d+sIs6boSSXLono68rd7GHSQzGjJW4c5
CFkPgQOvkpPQVIMEmfBMGP3DbG+eVzSgV9Z9RGH6I2YF4EiRWM/MkBonpk3qTjT7
pHSKNWe/AqgvJPe7eOyqGaLZRJjZOsQvijS5A8/agcoV/o+Wa5txcZF46u837wYd
y3LcI76cSi1GEjiAylynHF4SLUzIJtRc2OZYmlblIoFE63SG19eQxkfnpGK87Yqz
2CNyPJahVR4cLRipaqzZCOKzvdpnNLuj5DRqbl8KZEBcnz0AsicKGii+wIXiW2iY
aCzxNtmDcas2zXQoxUPuIcbrDWwe4t3kpqP7qtJtSXUy8IoqH0X66ntpKC9N18qD
vDxoVRFkVhHS1qjvT+JkAj4X0JH0w4ciOWIKxJG/ELsQDGygb1JSq/ADbT4CY+5x
hXtf4gaCl5nOFBjds3ncr5KRStLVl2Aty4TX2u2Y4zJJzDBXOIP8uIzkHbmBsbAg
8gQeVX9X8rcizNAhBpbDQQA8SUt/DSQgZSCyYas5of80yO5g1DNIrkY86FfFlI5d
GMwOfTuMQcbJ1fMTWGrN54blDG1VjYtEkjwIOhzYRaksB89bpMOQUSRKizVreSaa
N7iD9mCugdRrBLUt2/0XuSS5jPH+yDSm9IB3xGzEv58SE7JzlIU5aIaeujP/7O6K
X9n5z3UJOX3wDfWhMunA+UhEosYivQL7EBdP6v6id5PiBREkH8luN+jPYUXLxAIO
DOjC4cpF1td8eqNMJKSATfBU179sZJX2rehSh3B/uA7woXg3nsO8SCTCoeI4eHpH
x0SOtRHPukHnRUxjA2gGJI7xuu1bY3jitQrRYg5BZcTt40/lXhvLAnhgqCgk9dPn
9wZ08G6+BQeBoiTbLTA4va7DPWVehmCKUbcFEj0SNfAA26WT6mY9A2qvhrs3tIRx
mOgi+b7xylIQ5+9mUrFV3JItGoVG60dvLwYo1B1M1T1TC3PX7I/e5CgKuNNhOH1E
3X2A7niqYCIX9aCYzRReTuHBiuJKtXNCFPWcnwykDEVv5t9EKJ/Fdza71dcOzQq7
73VaAm7b2NIeAYiiNotcLnSlgG/6MAM6D4jQXtJP8KskaaUrPIKMv4EwdnCTK9of
5MkyQ7HOJAXpQNOVK674QxlWcsKj+WET8K7MZwf+uJqHKSw//mBXS8rkMXXL+/bV
NS6WYDD9KjXVXxiMyOADDyOPUHOdhBWIXfMHy9kGYWiQAoA/C5Zqu7F6eMU4scO8
i+Cb+B01qcJzUWDGwEGc5LzoAwKP719EOTJeKn7JjUoHHqdQHEb+j2MQ93/KoGC9
q6OGF4jaGSWXhfgHLUlyyk7iXCCoBwM7Q/HxO5E7rcLxVzmMxscMpTZ0n/J/Nh+/
6YmceXB77DQEOzDgq4wSM825uiInks68KC7XoSMTZl+nsJqRsPGG+ulZi+0mHJhw
oW48iXxjkf8t26/QnUoXmnJTi4KjDwd137PqoynIjckZEbt2/AkXvfn6vxKfe/fR
9EpeIztucZxCtjeah7YNBplRWt1TqjUbtVh6RLbSK9obPo8HrV03lnXts0UkY5cM
GosBO831a8sAnwygYITXDkjyesb2F7/6SzDnOLtG8f/J0xd6cOOy+X7UpoGpIeTx
a2C1bY+DXSRvJA+/w/NSRjwQeAEWXK5jtQMNbo2zKdVCO/Oc1NHiLhLsjwbrznK4
1KMTHdaFJzPShekQJPexJOcznxxkwnSWIj1ONDQOOW8ZVIN+JC+3HR8UwMT1jPnl
6Z6cBGe45ltoaa4Voc8NkW26ShCcPg615y8A+z9VZKylj5mJu385SpNueOEJlc8u
ooW+8QBZdLoLRHeo+8e8qWdDhvUDN+SEluKF7uRRT/5J7Wxfx052zKfKc2eUTkFy
ESHd0zsgNELrqIDFSgF1D9/pa+oSRjLteaAXOoua9FzM/fno+oaNM5vzWn9SIryS
y+NaG4qzPt5un2Yb8fFzjeuUTRslQGJZ8b4HL62r/YP5yXh/4XJi990k3RUQr4OE
HwwSvv7kouPyG8kk6ZtT7jMTPhzKryNf0sBzkUMB+bPY9sDXFiBr0zFSwq0wElSn
Cp63syy/zo0r/wlAxLSGuJqLPAHAA66AOFuyfjjv0oTDoEnhot73AtVeW0/Q23Y+
RRfMx1UdhXpQnCl6wPSjJ2+6qEzLqR9ObrYISk2GKgdZaNzK7RQD7M9Rb+IfLp6H
Abiy3N/j406vF95Nf88/X8u6a9QPGMmsI8Gky92cFs0mq7NazsddlBuYIf8Eq16O
bXmhJdlAAVPCHoPPW3mlbgIzUCs5rGhBvmBLnyKLb5zwy+j6p0brvl3y9TrNWIjm
YuhnNML4aF85GGxbFOTAomeUmZeXSgUa1j0NYqiTpxEfxKsr9AcIeofTy9RAUVLB
d4fsI9/gIRDiPCPaPSXPkCyYjg+cJ0nFJURzXKNIvnh24c8wjED0KSSxEEjSMR6/
sXj0YrbvJqvzqh7ov2VXLPJs+jR1wgXc/kB9aBDKkA4XpbubkijZ05XZiBes+tNL
AmA1ETQZMkaDT6tXrxHmD9VuMcmTStGAyrUuBUXRLfwAXMMF6b9+4W4m709IeRiK
RZmfL48hMHel5u0Nx9KAp8EDO1+doQUexuHY6UfOi0gweYWPk5r3FNHPt9RKfyH+
vWoso//g78ilObb1HefiUqtYm7D94WlwsoPr4B4bYMeLiP9wiPsZtvTEGNRxBS3v
wAvDUglM9QRqphzty1SxmTGDYFO8uz8gAuKPwGsmOwClcPh73H9HgllXoqYxRLg4
ALwxRSDVFTc7K3nJg4yqXG+DXxRqIAD8Z+QnFNLYZm0lzqXbMR9OGuoIu5b1iTO4
9ALuOOrF2DoNUThA7zhpXdMpdADODAk1B7R0YYuNU+PMh4G33tzXqjsGMIIzTcwU
jPHJpTzN5SKJAesNR/25KhTt+G79WL5g8Dv7z4oZzxA3i9CumeFrBv3xTCATgExP
Pg241kK6hUpz5CEqfd5CMSmUWf6FdXQPw6qgxJNfcv+Lr9H5wH/SXZfbJ1wg/zjX
sTdR9NSIKkEQfN1RYQ8asckAt/2KqLerljvFetvQ4xrS9hKXcQ4MDidD1y4Xt319
X0YLf7AiipkjkCCR3vCXaNwgPzviqhOfEwiYsHrnl/KxEWuCsuGbZZX+JlpIePO4
Ku1OzAPJZ6xMzEitsTAFv7/z3bt4K++gGTVY7GXkoVg91Iwi6Wa6vWVB7Uazi5pD
wyc0LLh5pq2tFSA64D8aIQU/v5zC3cPwK5NAIHI/gNuuGDLs/uwV5z99yq7BzYXl
YoWH+/dKIdxTAc2S4JG/9GHLiyGs15TOhC+n25QByMZLOMrJDg0yxvg1UXFSW34n
DAQxkTssNFWK2I0TlG9j5jr3DsC+2fLcrcO93aKvQYQRjjI5/4i9sccftmTeCjXv
OgSnm9jKM1B9x2B6lBQ9zmIKwDOaC4l5Y9fKCSYGHYycyQPUY66R135xe0/emDTv
EG0ftwub4UsFcfcXQARo3aSR0T5+cDHg4cwySxv/dYjXJ1LafjhDA0ahKwzFIP54
nE48pE3TpxZEagUuXpPiu9+XgIBc6AChjVFU96kTrzC43Al/+CMZA8oBlEnqgRvE
imW1QcOkkQw1Iaf8I+BHo5p6DriEnAodhtaVSffeNdcHX2cxcH6aewOube0EbvQU
ZYoILerOAK/+0d+amBQuN/rFNFd4+tB1iRuon12MwjQNx+wBwXhAlsdCEDI5BF8w
CYY1xOKDpsTbd6H+4rydVOliXrq3KgTHrhH+R1GtIC6wYTDCiZRkkdzNdCo9Y2gk
Tc2TAxDF3E+NqHkXYPdEX2gjPo45LnEsrqlAwXWhCpmGdFa0a6mtGsmSxaL/E/l3
S81DR+r8JQf/fY9pZXU/YU/K4znY5KcQAjGqUfKXb6ZoWXdw/B8lIcl2Mfs0+4nw
93NlGIAGmia0pB9BQ5MYK8LoCJblt3/RBka913f724wwD25L9Z5/iXktygKU0arT
JbulU+BhFqThwtprET6gCbzC3KHZA2uhZIwLftmaEjiVRtZpTpNbe0Vdu/KOyHHF
PDk58E+aeAOKroEYwcJLYZEozXTVP2I9IgwGxtc7SSR1egOvTYddAuByvRaHrz0Y
PUVIYsvJTHRJWcg8fbwvi34mEyjY8Y6luuAxCO5oMoV4TwjyZU7GYnHfSR7AWmHY
8iK2SIqkllExnihC88uVoaIrEagTKmVQOtO1R8p25HtLH9R+P/3z9ijKURGi40WP
5okgEgNgeRcJB/M0J493jiOslVQhgGc02skoClBwY3l+QFrtG+iCkDGHk4Fhqkzm
0R+iGxaD9ziCd1Ecd+Dw0ZWXBC4rIbSLV6Tx+tKowSkHHfUsxjL2+V70lVPORRbe
8dZ39xs4SmBaE0Nx9knw/JPe3yGeaMrIK4alZ+gfUHCEcunqSDePiZH8nkgkpnyJ
xsYbIT1ffTXOgB8+WN/04hqlksHMkeEHl8cQX2PT0SVIHYymivth7zDc4VLbQgkW
9cTESqbN40757DtrDv5mIrwwW2YJ4IVJmqTsSTiXIXb9KQjJE7yav5u8Q3daOFQ0
FS046ZPvqVQuCmsOCkERieOWmfq1yncZ7K/yyTgrFhom7XUk7lNRc9hTquAbI/jl
h3V5jT4wEShDdddUg20MSfjeflMO+nO/GCmdW4QKonylBvc+QnTkcpXywvKtrByV
Y+5eOXXxnfFHaGppReR3f6qqCy7VITgnigEulDcQycjGPDRYxx4TYvacrhFTA0/+
Tu97/d/4emvp0aYaMBD/AWxGFSllv9x7wOSzB0NfNgDEbM8Dk6GRzEfe1RjQrkCA
y15icv8V8B+UeTyxQNVmruhecOrI7lc4TZzvfb39/NHm72pmGeQZN9JAFnYoCJdk
v53zc14cCOss4EQqPx3Hzp92EXT0Laexw8W5MTivJ6+NrRJKw04lUlvj0lfaZCbo
slC22kl79IWcNtH5tm6bZubeiCN9VY79Qu608vUKsKaR8pImDFbDl5o+KEMXJj3H
o/pQ47gorAm98mn54DdgXGCv63hC5ThwbnZpm03hPGoo6TgJ4MKM6gJs8h+Nvq9E
NAkBxZfbVY7mlpvC9fOUiD8N1qKYOZRHqErORrSrrg6xA6p1PgozPprACmCi+msk
FFsGWutfIPRiz3YvQXvZy6EVYXQuzH4hgPNICz/QHOGedJ66t35B13ofvPTzTS0O
Rhl83IPM3pCuNgWC29aLjjAKuXwVcDYuovTCnU9qs/RLfdtJylwgFLDJCpGtsK6j
X053VjUb0ExLMm62T7zrGNbAc5swDKm18T5CT4Lthmhf49VxF6XUVLJhoLlur5c4
LqS6CAN7xK7eqypYdFG3clZN70/ZuMKalDvduPscnUQyUEzAFHfq0qTxNN9fHBxW
hXcet0JHcORGSWlhDe6VSHAFZJzBd4I36JfGAedmuoeK8ZeWh+6QFR7OFyh3SkoI
kqIIudpPYE55TYBU9yxHNCi4ScRYAmLcITIAoEFYYJq6jgdlT8Yfmfu5yWAR6YLN
cUp4892nEqS0pnkbjt/3eJGRJQ5H2A0D0ZFwbXmwpCj5HrR3OZ8HcQgBOuhTcjM7
J7gO9AWGwMdHl44J6VNCSS+HdTUFfCo8iQe2lNH4e+rUcOuVtgf983ZDlnYiyghL
P5+1gQ5IFLdOjvXOuH7b73RbwEoQfuaFIMy5PkvQhP7g4P1yXfpTaW88xwpzGX8n
lVQzTWo5DvifQueubwnMR9o1jxniBr1LZRAtqhJLngdsO+pd6sHEadfa1hs9ZOy0
P3CR8yAGodZbQI+kYMcUK8cxdfoY/E20ixN79ZvD5vdJgv6AlfiwjTeYryQyKy3Q
eKsfwjci4LJqrmhwnHsAFOBFAv1wlhhHRCfhnDI3DkJ6U3KItfNw0S77uXkYBtdo
5PHEJzPL8wW+oo55r3Pyxw/dcgjZRmdu+D9SIoGR3y1g7RCkwYmpTg9LFducoytF
uOFyPt+5PcJiT9oOmq9LfUksJvjOaoLPkUAgdYSrkgEk4TZe0QtJE0qJdq2gjD1H
+9Nw52VMMLIn6tF9xxjl7oc5qOopv7bENpUTMV9ifPL9/q4e7u6PkNAE3Jf1RP52
pE9j5PCudkXzn3jD9YkZY1dHxb8X21uhEvYtswVKmhYUMNqobNrbinzaltIdtDL1
+3akygOopm8JVGPzj6bpNNH2zfs9OSS+XgqUE4rhncVjYbO21Vo9DgZy3z7HkpNy
9hvh2GlLV7a8RfGMM0BDZYqVkvx++D4zBGyKuaOcf3o/KVd6u7rpnAtFVdbo36zW
AT9j8BqB8SH+13un6IWzO7q/YORgMmMd3UyZx036cWTkXaSQb7ecFes6KBJo40VH
/1YHhw8PdMJkjNLQovlGfBwm0pZ+wnG1cnchR6LGzgji3K9LeLGoHb7td0R4f9ie
CGyRdiZpGO+AJHFuxgoZjKZJNmsg8zMM2FmnoYdQb6FYFfa30fbQHURXo8koyHCF
9dx+cJIMpOTjrG54je2eYfO5YY+6cSmIHFKZf+ke9AeMI9k8Hecdb5gPVFETTGBV
KLgDoY3oMgVgQBxLUJKERk8vPQjiyHndgR1w8OJf30y97tFUxGu+iHGz5Gty5uUd
2lyo+jOMrAc7WgKl6HDbBBPMyWqKqRorc0hflGtX1MDgAPWRFwHDHHtKGmhLRDSl
yFFU5c38zyLjWRltVkw6MsOghzLeP3FP3H4ohPo2Q4RcFIgE4p41Kq9lGQf4gIZJ
2agXM9YW3Ry9uyTOOmBqKCKTiqcTdxYlzBpbtt+2iKL2yp7gNIGnjRArvGzMlXZ3
rInr0wyCvW+V6ZrfT+eX+8rYSEDXdqEjXU0bqAa8SvzenK1wTLU/qXnl6gaK0Rtq
yH0eG7fr2UVs5aQ9F8bKPUzqXOUUjI6tlt6nX54ifwGiswO11XmFkiF8js4Io1eb
HmfM3PI5Xnz/CSgYyYqJO8ykZHfsnSIwYuMg1J0VGIbyXiNo+rr2gYij/fPTFmwn
PZC0dGfdT7bNK2etZgT1IQysT830+mdky1LiX0tIvpKm5VLrIMrjma1EFQMrtTRe
fP0of2foAqSHZJ646vq3br9IXjCGkKqKaJcDIuSdLdc1ASD8XuMgXT13NCov+kbR
JAHk1jU9agLrgGZTZsrvgoYKGVzbu7KO0g8bTtp0r9A6vqxjYd/U87Av3QqiUdtN
GD1jkwjpoWtcVo/62uF+UMgf/mh38VOYNQarRdmt3DH2fG3wqRSncaYVlBS6U0u6
mxZ8Na9/zRbGX5AqNmC38nUZkLFL59HqovqzJvDpL/UrA9N16EEqAwwfrGSkAfjE
EVKNGwpmcY+XESqflA+KzXEZm9r4JFP+3ZJGk/l3IlaUiqQJNM9WTp1CRmpbyiZF
4ekO57Apj8/d+DyW3icERVa5kTS/+rOKwxdKLeSiX42LK5bAxW4/IqfYTvCXoHZ0
7BZH81yn7fdQW+I3WEHiycPeaqkX+o1+W8ZSXhxt8fE9IzUFB0QI2T0p+pNoVCEh
46PkL9TgHmxU/HRdtWCkblckiRXy7XaSlbzh3623/czmcvfeLEI63oexQtAsLU06
mQKk8Vyiv3EHsbNCI5KLAK3zIjEQKLlITUWMBE6GFPbCGI3SO79HV0egm8nU45hh
c9p48Qa5GoX2ZC1hYzM/+V0zxRXscfsMet/Oy6fArMDohy0dwgNeqi9XC/wCVwKt
0KLQWqGLJTL51R58WTck4pI81qoq2Bo+L/bWQ/PkdunOerwxCUyFkdwsWmUA6PQ2
E+146bw+BSOGvzByghfBeNvXiTSZ6fvgmumhKjWcYOnplrwN3HMh2ktLvjqbqo2+
TAXF1dtGpG9DTY26fK2GqDngqdkDroDhmKYa/AhpULTaMcLlgA7wfee7RjpfSKH/
9mc/t4/bm/vYNjXW/eiPaV4nyJ1aJ4bSs3EDzmuD9E/luX+H/DZiS4rLH0ulj9O8
iZUJCIVgYVZYKWFVQz0zjmbwmny4EZfdHpmcNa1yS2pi78JYCg92BmzkjfIYOm+Z
WnLWKMDhcA47JUtozyuV+c5wllTbJSGGuhXhbIwte5dFdOu8DL1zCQyEcmi2Lm3O
/OnvLdAR5yccDHaveACW34+QVFoI7h9IRe+IrINGR3RKKElUhDEJOO5KUSOdGqgS
z3kzBVp/1A3WyT0Ei5dblTyuHg1OGuAdYiAkB6mSHxYscEH7cfHPOQVVhwtnimt0
p8XldUxfJCRieUXYSURqEaSW2RYwKk3eDbXgBwCaFYe2fx86eoVIUL6Awz0zGJ7N
nNosHzTIQeJjkXUf6IdtBxYJXyaeGHkaXJbcEui92fOGALK6kiVz9WiKKnKflt2D
SqdYnq8DKS5trgCCUH41L511JLQvI5oXcmAtqZ6PzAGncQI5VdGPQbMNbGsZIOyM
YKbfuRjAmqD8hmGqx/z3500E3XOZhvaMAvV+GTbXlX1Z9rPEnauK/CzeU/PXW7iF
1q7z14pxj8DubIml05g9Fhc2GiUSYxK6FlRw3f3CQLbskI2UNPGPLd9R/SVGDOQ/
0Ay/CKAC1s9Sp/7Fi7Wn7lq1f+qSmDACGJZPNG5u5CRiqW73JXNLe74o77x+8LPr
tUnMspWnCo9M9pqzw8otAqNT+jN4+pllEiBMU+dbxfQVU0frmGJk/m56EXfvcJD7
Cfl+/u6agCqXqGdi465cRmhiVaKOGV+aNFq5ZzNok9i2DsIRt1anC1Wo0HBaJBc6
YknXeAglY0wM0aK6uvMAVIZlbmQSwvGEdSm5kWBrsnfC+CfmQ9pJUZSCyTfFAsXO
l/ERb9eS60YnYKH7+lpQl1h9l6K0bULwdBYxysNA6PZ7Gl4+ZG8oByk0V/aOx2O0
E7FwqbLI51E6NiqAgkBOBR2eqA+VYnKxYS9mnOEpKQzQzFwZhUwj4au7AGD60y7l
JNFXcRpsrc4HjkwsW6WBnIErwlofUAlBJXMc9pg+WjJ/jkH4HrR1lZ2GKiv8vhvK
vV2tzYfk2mZ1aXSazfax44kMVVptSkdMN1huURrsoiQeVB/YdRiR55yV/Da+fHEz
defzvPm+G2CpWTCymOKI6Shbf9IJeNM+2CwWxDHjnXAHeOVIG3f/V51dVkUfRNnP
38VU95JvRSLnQ5R+E2Bfkpc3Op3733boI8UljQ6Ogh4rXM6LEaLzXhn44/QBQkWT
qVu81LQNQRE0ZHKMLEzWP6Z7jMFPjGSmgUNQVepdFgnt+b0GnEf2++pwCexFfY4V
AaZ5zTKck2NUdh/yhddhDIBRKktDNuiGLuF5PUkAStA9TXU2uN+AluQvjHdvm+Xm
NftUNoFp2Q9AmGZtC/U8/M+KQHYLYtQSWhui2CVmsqjK2ydq29cyB2i1NPGCfoDC
4IxfOsIdrV9bDjxS2yEJ4ppfTyE7D0klctg0983hWpYlqiAlsueALgDbIuz3X0Cb
r4d2zMaIRUOkR+0KZXQim6PQweQi9V8qztIVjxR1dfwZbnpwR/SYj89RTaLvd6Sl
RswzhSv0If370wbrfOovMHyz3gS/hL05nDUbLV1dXi4RkUfAsugy96zyBFeIthk0
gWWdgyHi7E8LocX2rWxugkdCnr11aJorzdiXX3+mplrlIUpLzP4FHxm6S536gjfX
hOuON2iDxf5ShyvvRi31SbEz+zXewrap0RZ1F/4Zp5NSJtVMJNUEeRvCGdP+mbMJ
F6VpAEEoAlj8cE42VVlSzxvUBDpPNFw2l6YpqMFPQH9McD4MxyO8fT+1eAgSANGQ
5/l2X1cZ+KoPGddMl+vYTip/Nmg//8Q0a17R9kA5Uw7kNG37dMQ6Zl+aEux6XoZH
/DPRhOMIY2tJAhHo/lsL3yGQlrmamR0d47jX/epOVrpSS+TBOwQ4b4z2KwQ/4F0w
4Ems+Y8iNGZDd22LYaRzjooxKyBC1E10E8ewLFj7jZi1T8BaCuNLBsbAb33rieV8
CO7wiAWhHE1ndJP710hNIy7Klc1X6tGee4lNNBpZ8HotVliDbumRm+uA5wB4zxXQ
nkNdjRvJYoL3r/uJZn9/zED8guX/91RDRjnUQ4JzNEJdNmSiXds/Yj5d9jR1YjbW
QdEUaUYHD5jiaTUzp3oLZ/3sP+dkT/ifqNqYws+qI8vaggC+O8/e/J5Zw6kZj+so
q7i4PkSEJdTHd+cdNYZEmnbIcR4aGiFjLX2Jl5C+W/HAx+bM3E74zVtwePX80pwi
p/G8sZyYawBnDujstgExKnsRCyRbMhcoTzsGg78ZC59EhI/i9V9CmQgZK5VQJ72G
OIfX6aDZB2dzXzSJQU5FTIfQy/b9HTmrkBxPFNwV+3bb71OQ1FCb/vJtQni/U7bY
fdX0keym5h5wQgeLnqnMuF8p/dDBvlpu6JOudAKhKRFQYOVgkEfXn/tgdGiaqwYZ
JE7oD5Gz/4XO71GWAieruYFV4gkHecQi+gBaQGCcnHZK1bHQca7BgMcVsIqN69w9
RmGXSM4UsDAHKGV6ca7nh2sCpnMgrNWept7FjVMa3ndo3aFw9CosTbT7u3LAXFAM
pnr1me4fLsLdweWhv9WruXoPRvX3rSde15IA6f8G3gQ4Ru25kfzJJxy4crmH//Gd
3GCMiFYzotNNTfpxI4Op0/5eNrdy8wJSLsLDx+OfurtWVwi1x95fEiJvQXMSTQH7
I+3fEXCSqhQLkNJlZHEoYvbF76CTcVEGdG7JEwC+uNLs296Hgbx1kIxTU2YvouxB
gvwlGC4QiZO6p9pHgGZlV8Z9g2nF3SDkBc6UTyk2C3LHrRTOd5vOscHXhyCTjw/W
Rj3agbgKw3Un766gXh3yyaP/5Rs9GFxvHs70BDjxB8AR0fdl85aH0YQJ7z3W/mk0
+LxnXkd1AX6TcZFQJA0tmpr4EmhqDXTRdw7itBQCO3D8IYqxxa/vDn/uTBm1if5G
z2w7ClMC+RNDa66GYGuHVIDLzr2cdhGUx/kZ7i4UFEiA2DMZVRE+yshQUN5Is6ue
ihyczAbkdGGKcg+Oq1bt9X9efKPzQbHEgHFBjBKiM7l7Sd0i33IcC6+3x3xhdzbq
psrbb2FCA1jOthLxE1mtnMIVE8QDEMrn/35vHKYHEOOk5uYjHNz3RKZ3criiphAR
1umm+f6DnN1XecwUQihyKxvXASh1/wbBak/K5gVC6iLRfbNqWnAXMdQa6vzguA7c
9h784s07LkGzZoAs0ZfX/OJ1kdEV8Z+66iU+5tYFNd0ikJBg/yNH0kdtbRx505mK
+gyGPOFHp6YTOaNh8/upF1btg0uSCAeIO8s+Zn866BJVOagXNWcXP2zhL4ig4Gb/
YZZCroqj0gZgamw2tdVG1vA58F7qJhbSxfby4dSSS8ii5FSVQlP7/yRJL5CMr0Us
WiCu6sxAozoR8p1xI72iBCoXZBPOudC/3AHsxgXW7eeB72WKW1kQAt/5M5ub78L2
XlvXJ7QGGvKWEhWTouXbAJsdvRz7KyMWaIp/D4xnMXcBwfiVVReVTmd0mHTkslh5
X9QaqMjPwov/xaOINuI+3ML36LmVcoJnFod7QpuLn2kYBEzen5JOdCkWZJTyfoly
cgv2lKomAAlDTclUWXBKj2Cqg3SDg5TW3AdPKbHQIIYPHer6doVE+DqPt1Shbl3w
BzNkZn7t+bFfyw8A102M+U9qoYZm8LHtynHLgZQAHvdW2V0n6lwZ9qJ18oqsWW0z
FuAPbrVZsf6Mn3wpvLgeytNHkx0oXeqLDw9El5TZFwFlREmj/pGM8oweJw3RFji3
Dyc7j9ooMVi5/2shHzjd5weGdwkI7iHI6bBcLmdJUdgjzu6yxtxsJ965D7STHcsT
k8XN/hMP1jLjm8V7wP5A7pu8xVY5cHZWvO3avT2L4p712P4X9aGRF3iNzWukxuj1
xKjeEgDGbI+WvzVuCJznPapw09s+S++QPUMET8epBWMlXf7mp2JzLqVI457qNiGX
tUJPk/QuoVjDe60AtecKTdqSh1PRhOXy0xbecIIPTDDjJVZ6UZ+ClOXKSHNwW2Mx
KrYt1HzzT4ci31AjMGdeuzWArqVsi936lZfRlu/OaNDLIB4HsEQJWThr3S5WLYzg
9UZl9G8YljRRsVQNfSmPfP84dwbdyH0t1ng9cbzqgxqtYEDA4u/9n31xj5uulFjG
Jl6ceb4dQzn8InO0eh0O2sT6wZSEQPGFKVzRxrskTtjcJfnPTWpp/XNdRDqe68dI
lR+wnOJgDavSXssnlN75hTT8NQfL9v0ano39i3KHqHzB9EY3EyCpmAbMeT5uJPCz
P9U83NjiEM6E5QTdFSbcOULzlLsyz40e+bkQyHsN4K0Drj6J1drshEIFNQjnJ1a1
MnZL7wDU0fLpL72S6eg+wPp0RF85mamzr6HM9Aq6ghE0NQmhtB2AKmrmIIUk/8wM
dQwuvhcjgj3KWg6dexonLUUbTLABlkm7llRqeNEaeGeAIyUs+yalcCRwTdBhKG1/
Ea9nWtWtt+5qxvHL5J/+wlMQqeqwNOyqxlL6TjgHi3ZCT4BQyAYkLSQFCM3uRmVN
El4yGHrIq/kQNV0CB0bmInTM6kPyDsCgqx/TWjilzCoMMVzIjQX2gcFI9R5JViz5
EKHiDA3dP5Qv4HjvrbPVEyEy9pfg6NzxGgZDyiTBLWuEpwAr+/2whiMDpQZ+vFyp
zqMyvJrZWKtcpiXhJ/rwO6xqSEBAlKl+Q7k3octpqMFaUlXybDH3JLhVjfHOJdbw
kPXYKZTTOg6uaI6O+Q6nqKJXF9LOdwvDA4XMAXAoB7OzI3L93goUU7m/7rJiYFTE
npdfQonGmv7L3Khq3fs+VoiHn3aGDYLm4ANuMlcaBd2vgkoasSLyORx3MPWK/bTt
dLm5VyVXbx48hpou83eGEeZicaJN5EBYtatsjVRhCucBoFkwhmEO4NeeZTLOUie0
tljlE8N3lFyKTxb4z6h47K5BeJgujgY3bAkNumFmCWxdQKUdCqlHz/reOUX7B5pk
EjJJwgfKl3bWGPMZqTiXIY3dqEvfDfjGMy5KYx+cIhf0zsSotcLto3qgwBszm3+2
A/HbGBvao0ocRU5wHlPoAh2jwrW/e7NPxv2Ocr5kEWFSpG4iH2sqiZ2+BqL+zIBg
22inDeL8nT3HxWynRLM2/PeGt6zlyvztBPyT0vPC5iM+8B8R1EzhAFQN3egzLjoV
tjaSwbgR/94nNfauyD8DUrmHKU8zWkO/bf2MHVXqWELA9HNEfGMkULBd4UL0XxAH
mkzyFZ2Q3LjATEpdCWb12k3VogtQSD6yVNwZ/oMoRpIqtVaZu/+0uFXpK1GyQVGp
i9PTscDq1rkAFSCeAc9G0TuE/kGjUoU1v+bu4OQHF4eU0KQAtHe2nfknH6+Ca314
8XG0oe1lc3pCKZa/lcRjC5h+oOevcNtqYcRwsKrSwpdtx8n6yGmATL8jnRmbJC/I
AW4B2cVbzNG5bLYOyobXiP1Zz6wM1dzx2MRCKhyJ/Sp4EUwIjisOYD7FU4Fneeoc
t+tETdq2auD9WlyMbQTjJc2sCRsUEl/68E4cCNcQ4CfRljRQfw8hsvUhaiEF12Dz
wd87DFzcZpM2riD0ggLDhnoS7Y7qfx8FhXvh9Deh/ND/Qsyb+aNfW5eO6B31cOKe
FTUHKtkK5NgHoMb1ZbfuVQ32dW5o2n4yeMeyL108eERUM8wA4E9npDqXp8yCitVY
JYMkuofnBu3hwzt4m0uqPbItZ7FGIzntWOgoPm89raC2WqPiQGF1m7GbB5BfmvnH
v78Vxfz0Squ8WXfrO5uvERpY+0omEKgIEgFtN5NjqiafQwLu9AAGCfb4huupBf0k
3+PxyaDmSQeKEWhtW72zyNxphWqnnBvNifGs70F0tcgU2RiZVX2tcunyVPiHE0HH
J4ZOYuYgups+FgPdZlxwS97p8D3DyYFf1A8ag1BJyhOXJMoni1d+SSSKBcfp9NWw
k5Sr4W5K4hxwtGYmSjaSw58p6ZVBKDN1LmwJE+DwA+SupeSI1yEezlX3YudIl9ZY
ZtH7O8VDjfUpgRCwIfE7kR3ffPtLoYXvkl84Rig7chyfcyyZN6fTlmtTzfK8ESmw
PwUcaI7jAQvIycOtFZ5XhIEgAc819YLm59hzOeZ8sFUlA6DHXzqDqYU7htAC6G+I
zuuhwvfkR5DhUJB5/D3yGlCL3F7dmezLl5to/L/HACZmKL9NH/igncXjlUbFJImK
AnEdQ8++AFqgoKKMszB1q6h/05salJOnV2wjiZOp78sGlQ7ZTPbS8og9x9k9adQc
mCFh1GMVgHfB4gl7XEB5vbyw1w8/byq1zT8b3wWrSfghIn22oPC4duYwYromX05R
cF23nxgoMCXduSwyzGn6NOtNHc1wkqgzsznihVScjghQlBsHRIbI5QmGp7B4gZAY
l9TbZICHhi4MTaIeK/htvMfNSiw56iNbVLEDSBfpkiiKusN2NBtd5G/HGo6UvFJ0
eDsY5MsxrrXrZjLdBbV6xwgcg4hunuJw1bNg86zDScRZEoJY99JgsZCu1/Me9IC+
Nh0FTL7guuzQ5T0u1wGSNvSsVrnawlfS0p07FGtBwA99eK4Hn2UEsQGnD/SJN4Nq
KwtBUD1xCV3H3mg2SRQqwdfX8j0yjHeDlBNma1IHtssBuYAOlx/g3p8vcEe5LDgx
NEwx0wF1z63Ctbb9mcPIyEw4VgNb0QXp9rflDVcwdDPTKReP9496sP0F0L6OrOZ2
+u+QigCIDCdFs8jiQMhkxz9S/Av/M60QSVhmT+5zRRu+jpf7kZQOKFrEThUkhe+S
vJcwb9ix1uOltl11w7Fkf1l9YceF8vvEdCGKuKajHIftYDIsZjNn2/PVNs32D1nG
VAh5O9ZqHcfm1VGgcAWdPq2BavC/bpZAEmpqLjAN5m05VZhStWvNkC1Og8X7dSt7
qeJmpa9JXPghr6m/k3XxqNXqWjlErwLtXL6gqRRaIy0yqVJ05Y+n8VNsf59PysRe
FnwQ2A6Y8HGpjw9nccSCpmrlLcPaSjOfEy7o4Sswrz87fNitFtWZWmkk+hOF0tMD
QU/NVWcnpZXMkt+fHV/f75FZ8awFKZJ9t2ELZENNKETPxuqITmjMJ8BLiK2Nb1Dg
8EpjlXJn+9U0yP8Iq/A8l6iNiMHQxwDrAsGWSzrvdcUYRoP3fMnvYdqndHas7B9Q
2MXBnZqFqyjelM9j9UtsYpXe68LOB2gR7caa7CLD/Yupbk5swZiS+zReBR396G4/
cyKVNEwlrc/6JyC9whZEF+uASxhc3uNWXI6iLpl6Zgne7sNbJ992Mh4ghPSVDBIM
yL6Hnpjj0Lw2ANaA2fhtUvVo6Ss4eZNlNtBiH2iutyHaiPXXaQADG8Rw6ru2iuC/
x1PkofZBJPSucpbbkZWZKpVLYoWSy/NVjfnC/rJNdDF8ZLbSi6nPackhj6I4/4Mr
r1o3JjFqbdYsQjqw8dPmKMaoieYaA/cOsJpn9dv9EKmX0PnRSde5VAJN7DqY2Xjr
6mL0gpZcyqzhvgiVzYEmEhAAwT6moQW5aneei9wYpbjOH1jgAimS2VJLq8oZArxM
2tXZJgY9ejvU22zrZIZlLNFFEztJzCdHTrN9NKYVrawu4wk5WVl1cR07ubWiLawt
QAtgA75LnH32AH6TPzg+po4+GhNdZ9KrXLPDAYPgBHPcPRpl/v6QaIaqNT3DB5O9
f8DwqUfH2079yUfAQcvYcRfX9GzKnNOzYuGsoGbZy9g3DZbgsPWYt2DUzFQXQZfh
mBEtGwhVOhVS5uxGMD1fK+DkmqxWcVPWhjXPY9TBN9HoO4KiwE+21kP+l0fkcqWR
lj1rTqweqs00mrZr9Ohweld8K15chRaDyTP+/bIYRYSSIdw0/qhj9wsJabUSZ5XT
I+VHSCLgodt8pZ92+sfZ/yPmDmWrXw2eJxQ2IbsLxG1rNLrFPvgi26+iL/tnkU0L
/2WRsDwbsNL2TrHVzvHVfgx9eCWdwrb1ljB9SsgONmQO4hRgNmgz4H+h4Znh1+37
wTDPwNjLvVAtkTWeIUO92n7iF+q+gk/hSNITrU7XglCoWeD2cGXaubYwrATiEkBa
Nr0cwJvMEJqdqYMCRQsQC4AtwOy2yqTg6UT5ZTy/OuLjb589jHXfleQNsCkJFzFG
agZ8Uem6QQFfCkaK8IAT3eelVSHaMOx0UAauqoxZNyaH7otTg7WoCXUTE7wzLRHH
3SIEvAnbi1egM4FcI5Z1vlmZO6grjNDtmQonmXBbSMOitGKldoaMWKRKGxhKnjZS
T9k6NL1D/St2iRp2/89OpacQuWBvuzud38XVa1rlSIcl/w5evlbveapIc6jrXXVA
9Y9DWoIMj8PDV4IAGa8YsmydiYuf/hfdTjGWyoOzWp61GCCLkwCQwn9esBYDY3d4
FzyaUFH81eaHKoRQpTGX4oykdootcr6i7l1tuOsMytyxWUNgCX/bsU6ZO8AVrprS
jXZF1Lp5qBu9iLs9YgldtUjDGpiujkUBpu+eHFchxGAmdC6psPNhKBpH10uAxisv
7iDmc62TU7oP3SmV5HfSJXQ0ppiZ7N2vX35V0LoubpbibRKgSukOPAL89NhPaBRQ
ntI1u7FIqXI1Q69m1Bjs2/DI2yrBMMa0SezLWfoqj2yLX5sELW25if6s06pu/lGm
sm0uLwyILTl52LXsey5qVZytipeKHVJUYR6tzT8EYoYbCvbS1WHx6L2JbAI5uJVt
GH0XR7h6Ip1yEwbHED69ae0I/SMRfTCBM3gHWyAzIwqKmkEs++7w8Etm2if9vRA/
afZGpL9EE10omu4ddJbBP3pRUmlAWnnSOWKUWZVf7dbVUFdOhgf2oa9m0mkZ5/u2
FNSVgBiXgY8AWzMdfk8dkwFotZt6tJzxBYlK9bLUAOgzW6wS5BOq0o5O6ax/1JU2
e+ur2FJ7IfYSa4gq1H0In4uSO9SXgBlah7PPUTIT8uvkvSJqhZ73VG+3DAeuB+BF
OkBLVe0jIVECRbbrh6VvARjxd7F1fGCFtMtZS0jPnpU7hw5PE6R8bfTaoDokYt2d
EPbSWyGGekcm6l8IH5g/vTrIk91vRWjyS3om3M2BEkZJxxz0q3UBi3RxaOlAfC8n
kqJUcC6sHSgHBPegUtw2TzQis3pidam02npwJagx1j/baIJrYUcCPE6TdybZjU45
dkrgYPEgQkGAh7plUx+vf/h2E7sKrZQzWRJvrfFDpk+Vg+VLObZDnBAvZ9R1nRpV
51FdygUkySk3okEyHByo9+MT0hWZtDCe5RKZbdXtjeo9utJM5CR7FI14Qwp6p3B4
R7evo0AfIMYgutk8p/KeqQN7KBlmFRTcejUY4grGz3g3TgaldtLEGX+fjyUwU5qz
qQFVckOQTTHFYgD9met0w0ET0FHdn2oc/1Ww6YJXgCre8IuyDqxV2LNGfktkxwXM
8hJneVsfN6rGhkJtmXLwykuJNys5Jpd6LETyThZW1NGIYues3/5HBmOcSVAgSJNa
ufCu7PuFcQG99CHtLQpmPcG9fhrxmeja+0W3uB/X9S5RQxB7e3tedVxAeGCLfIic
2rBsz+Xuw5CX0qtaGtb00IQJbgzgxDw7MAdaBUh3fMBslgxlICYvadj9ZJM7WyiU
8r8JNIItQXTh1XMfjXTYRKrRxai6YcqyCn0/jl9osXs2+1HRnXxyRDSU0yuIodCB
E9F89S2ZyOFTyU9VwVcniAI6u9u8TAmOCMFB90CqVxqpncYh2onnLzjDhPCmmklO
b9vvombXyXhDrSBq3ryrtlwxF+4+YnpEMhyol/pY/v1qCRd374gaOpSLHZq9xSRH
jT+a3WrTmXW0S7pDpRKPfA//99ZEtBztyA3bjw0AieDC1oJUL5xn8zDL8T4pLnLt
CggEdXN3nduZuIeBPl11JSKFhm77zPOCNN8yIwvLkikabCXitIMKOruhgwJTJcCT
0asJ2R345B22ZeKD7Efp2ikFHFNqutwUIoPS/2yFEPcuN5Bl58eImQAH9EzsPWYA
1KtgGT2k1vtjFpp/gULr/+6hOy0W6OWlHrJ1EMJk8vQQWZusJTg+jSq0FwFZFdh0
FqVku+vQzP+zfmcceG/5PVDoeFBjgZFx9PTRAHbndxkWDY3ASpYWcrglBYUh0XpO
OfuhORMhQltw8Dpb1WFNvKZNcy+s8vY2m0rH1g9NJfaTcpW5ybDEBskEYBSWMoTZ
gLAVh2hTvcfHrPvcmdHbVz5NB543BoGrOCz9Yk9BvY5aM+M5E3Y7CAxmDbHGZQdq
57iyMbZ44h9R0JyXip3tgkhAt5eb69K8Qf/+kT99P1vGmaLexRX9gQTGPjbar2PW
CYulIrNzUo/4bn6NNXsa0JWKg7IKLRDmcIyj24499x1vk8o1OGZba+dHdA80Rgkb
udfRdcE0cra+uKq2ljk92JX6vUXLQkqcKCR44OcKP0imtJe0E8aQCReLglawhLrn
0AsVnYEiCNrbqbEcqHqYzblM7hmvF4fzwZeW3LNepUkH7kG/fV4puPorNmoQUj1t
SkbhDM0quRbr8R3IvEvFwTTlY0X20b+2QXaooCCpOkNPlH3qyoL2RcaSUp1c1xr4
E/HVCyngl2RBTHU7i/IQDuQy6Yt4ioZTYCIfxLP1+VO8xzFBLnL9vqRrdn7Zka0I
ky70nggnM9i5aCnB3M8ZglWeK4vLuebhlvQnLgwVITIRSjkr6/gdRJ5+MnFVwdqN
4YL84z2CAG6VX4ymn0TLoQ3b1P1nQrw62HOtQctvyaposJ/1ON2GFXc7PngU8AVy
aQ1UlvAb4piigTUrurH94Z4aPR+tDgkLYk17wX441T2WPtgMHzhCU3pD/Ir/QXsM
r3p0KGGk9WvzNKqne/+tILBxxVsX0Wn2WnJYZihZvjGGWxcJZFttBpHQ7pbhk6L+
xs7NOuhkLcWW7svOdGpoyD7IEosFkHZRyxp2dhIq3C0Crv3GXyVvaEoAcdzb+DWW
tYagOAW3scZtH9ArnTrYLxWKLYFJQ6yp5mlYspFpTHB/X0CtgaqKaRzcMqproP2m
5Bg17kXPaRHZyAqpVNd5dOdk/UJ2tvJNeky3uKcLH+ixu1SWUBEcbVeZJBttg/2z
paAJnZcMUk5CQsbRhOjgOyZpQAcvudyAOmklfFGkodLZV7bCfr5cV/9FxPqFURoM
mSUEC93zPLSjJEgteY9cy7u/JvytAwO3nyfW/QVUWIaKHOhjB+7vJGBzuW9rn7JB
k2iYRYvXcfHkevT/fJWABhezjw4++CKezoXnzcLgtAKLzDPOxas/w/wsbq6A8P9f
uWPifm6y9HsU+62HKx5zHOMUIH2Z4mJSlv7+c5juKMMgyEsd4u1g+o/KaNiCDxN+
4EDIOsz61N2mMuDAG1Tm4Uz5pKXwTNAulcEUt7OIze8wYhndE48shBEd3s+sHgYb
BDlV5kXyIiIRWHtxQzYzrLlRI7oaWAwIfoadch2ZuJ25fdOw8lKLu/VI/vGjYuf1
E/LV0G+CiFoUzuBWV5EIOCo1YwjmZGjHupk17kJ6svWjqFF5/pZI4m4bmP4FfBnf
dqYfZ0CeeFhNAw7Tbrv7J+t4ezDSjxcyq/p9NRvmhIq08QUWgfyq1qZyy/LSyfq+
FmPMpus74C/OzQwCjdVOVl67R7lQ3r9gYDVoOErFsPQAKfpOEF3xj5b+rfX2Hn3E
ox5tIYSgzm9gbkbNdanTBcRiU+GpJW+ds4yiJX1C3QCeeHMijYGAOtUxxEv1rkmm
sE3sLAP+S0Dp7lsep95ttr/fEZ4FtMazU2OR9ByAaSMvFFAV6s8i+sAgGdBohBZ5
nfs1f+C5G1VNGkwNPdYdRNnxKwAgpJoOmPT40RU3ck0bc2KtFgzpnhSLQr7HmGfm
52GEve5Pf1J/7tIc65DPT/bu8f2TDOUJmvSjLKUI+Q8jk1jrrtW02OTC+Ij8k/NR
b9Es6QaNLKNUwgNu+5vrW3BeeD2AxFaq7VOi1HjPDy005ah2X6E3MLYT0rtHyuBQ
hOdpr3kzxSKUdKSpFk4tbIDCCKsK4UmmJ78jUa1OKh8lwyGA/73sY+VZolGHADGa
WeNvy6XXp4UrqOhbnGGoVZ3uvPtAFIn4LOEL6vGIo6d/f0LUZvsTYSS1c28bsuFD
fgIa6X3Qe0CGjkOO2a5dCF4MHt5V4B4s7kj8Xfdo+KrCLUPylVPPpVl5z8BgfNJR
fiwFqK+/GF0yOCydBVOJySREZGRNijT6HH7s+j6Va0qa8NvKWVcrsIZr29WAiivH
QmHSn8HjIh2LaK4w8pRXhaBW+75HwRa6+Qqou3KRIChRUdcl/u+Nr+k7YStJtWIW
By52LzmAB7DZ0wsm9+k0GOmVSO6bp2Ox6z41YR/q6oCJj01Bmim2kVfI7t8W52SP
4g/XdrX5LxWiw8/bCMpxkkI6VYGgwvySSDnKpFqjUQIi+URXalal+UxAXfXqcv8r
fHDUs2lDNJrkYPYVwZBortxcTEc6t6/elWoo8o5pduk98VksyGtQDzLOTlscIbMN
A9wf9CaaxF/Ihz01q5oIZFj5stCTXMneXxCvnAT5aCYmaXOUJ06UjYUElML7qMkv
H/wxczYsuZGgGRB+mKOfjy+5Ucu/IcjMHRETEyWrshtmSFqzPL8h23+In9kha44e
SicQUWb2Fh9j8XP8eLI3RH+VOzxNv7pm6PhEzCav4B+dvMhtZdWfyrD3qUU0Iocl
rFQ3Pm1z7X2rbvMSOVc6kQi/DQbTNBcx0o8BR5c/ZJII8neJWZ6xoElCGYFg/NtG
Xyt+5gjwGHqO0EYaFTMyRsVE2HfdjU4LJj8vkQPfWHiHIx1zmPF9hmnS73p2sCdH
SVxQeevPVK2YIAB3NPBj5ml9+LsyJVLBlNT9cYa1S8JL6FauGXY+f5rGK3tZQNOO
Fsc4kG3qIGLQj7hlAehuy0FtiY/O5a5TqmqaeOGNkBWZzaP8yNBG4GNl0ZataN1O
OABQIf8qmU2JXNb1M2oiSifQgNODX7dqSKsNYo7cuiNBlrjkqx37spd3LJlZTrDU
I+HGyJOBrOFi5HWIrSUqVn7OvedPB7nAsnydYl3d5gPTFLtEbzNA/L1XYFuZqJEP
1Qz9oyRZC/KDC2N7/cHvu4IPNu12b2RJh+gVekL8i96n3KXa77yIGC2DUr6LhAB8
sLLF1kxnPW+mHIH7Fdkkaj2OcZp5wkH0gCM7CSepBWMf8Y/Qpxz8Q6VcCvSY3jZQ
h155qlnEtCgOWdtGjjOYsfVY1fn/dJUh3FmNOXkOd5tiKtwiMKj42nBZrUINkMH9
Zt91qkgI68brqWq5gRg2ih4DYiMu4YMBHRo3hnMztfU0e9zXmGCCS6iNAxXDoKDv
nVqDtAIntw4zMQuZW5BMD0TomiNs86Xu8FRc21rtL3uOIUwaF2kC5REW6DBw3pFe
PYbnGjABiQLggKE9kszFFDWl2VDwZw2EfIucPAZ7LP4bP1aOGzhk/j4bxArj0c4Z
pvvTlErNx/JpzXUb4SN5mz2ghWwSy3/a9Dx3k8vnOSe0vITKWPYsBHAZ4V2hrV1/
qwx/WBZa5fNDl/lQD6EoW+oiM0XJvHFlgqo5/CN3mIrTkWtSui4s2HNKqL1pu5tD
LEss3AZqzvhO0e7Auys9PUK3pgqQ+/XUthU0ietbQoK6ehZgi5uWhBsz6NqH9xZN
3hApxmojYMQT0Ndmz6pi8T5ORNp+t7LkJbFGYQrU1CecW7pt1NQagmi6pJXjlLnP
sus6J5yEsUs/CPgpDJckfzuTgxpJbgkZ16+HiMAsAnjkYzNl0gNd+4RYPucKys73
kp5XmyWmJ9C4xMaG7YvUwZgumkZ40J+gsYZguCDB2KjMbmeNdM2SqvjmNzVg7Fpd
JEdhYrrz+zRCp06CcJaT2JVTrnDSindpIkA7mUI+NdVco0s9d+Uwjnt+tBh579pD
A5y5u8HfJK9vfzn65LEkWVOhgQ/KY5hkiUdQP5VpyvAEvhyC7mqldvmgM/KB3OK9
X6+QV2HnwHZGkv8ZhP7hYj740uzaCzyH2PTSz4j5lp0du/h/kxQBRF/U1QhpyNyZ
NyJtfoVSkNnCJuFBlA+Uwgq1nAK7rnKFpbj2c9wMYQ14sP9ONE2VuDjjS0oRSRpj
zH0qfdzcOh0mUbWjkBcn26D9RzxWlNl2unkgS7YnNeXsc4zPzfWBTZwSMzXj0k2W
/1LLbLBR2znwihaTFjHbGlhN2nTCkJDSDMfkngNpaXwEyx705upHZ14uH2GcETEo
GGA86anXnaWjLlqLgsUtkcnjFMLvQ9ORHA6Oo07KrgaDm2pfHhJguYUYWA5J8BL9
EBQFsGoIGZaCNOSbIsywYOl2igmXBSsQf3qW1yDEF+knTRc+Xf177b0s/zISnPbi
rg/xdHANMux/4FhTJqS8AxhkNvNa/AOFIP75mJ5C7RE3VxN4wHwpoJhpjFGFNQNm
QxenPulRPmc3u/k8lM1y1KnvxMfpThTMlvXBjd7PuYl8cYDQ4BCF6CgHetSkPEwl
J4VjHZEkid98DXLmnmKwnp52b/UJggK8e3kVqZx+2FAQ9pm6lXR7VI0M3x2RluZh
Q0eWxFWJaR+AcVSeBMg5TkJo2osjnk4d3VwGhKK3Qh2e9BMEWxqNf0tNvKuCGuQS
vm21THrruGWc4rdPOwnNvI5Tn4aSkwJlzUS6LCh1fjoe6I0KEuIiWN9+MA5ARYMj
p2fnH2ffqkjVVXpq9cKK2z7SKcsAnoRgtKVDf2raNq2msDkHO66AXIVM721pkijb
srsvWzrvAf5e4M0kl9B1vDvrQpcewbdJc9o9FX+JF1G5eWPctXDYktGwpjNZ6PFD
pD46c5z4EvlAj2/iKE/Y7jO6U6F1OM6BRgD0xBkq2SbHefiTaWX/thyMiNXO1O84
xlsDH+idVfs23z+7cH+FRp/hygydpjpAMBRU8beqj2f5kc/IuE3yE0F17sszSk6M
Z2WElguuxDNPMApdOPdA8AT3y/hZN/D0B2b1zlZnSzHkwPn1We9Vy50Hid9aYTAR
dQ1oHD1JIEt0zkH4kPbkN0jdqZijwlEUP+lcHtzmd25aL1E5H2nlt8zWFQHPNdCv
uGJAZtjXHoNrINj6pN7JqQiysC5/xSD1QOS7O/ClMsgH0GT57WWwtV4vjl75hmrW
uDbzrEYB6rL6hA/8B3UtNXxIVm32+mrnbc2YIHsIGpSN9iNnQaEbFFYDYQAcJxJE
FKdpi7U+KPGyAoEAUU63ACN/Xp5GI+PMFr5tVsizNVKGnktqvKZ2AQWLSam7I9uA
0VyJegwppv1u7BIaS4rKS8a8ZKpyXOQGAj6td3WJ0GMd77gpBuVtbPedZxdX0xtZ
1TJ8OdNAQHhZxTg3B+owGL4BxV+2dFvUF9MbjxI+Br8igb/AqVfjAbtCbqAp9CdC
oCPxPv9WGE0kgb1AA/1KtZlYCFVhfwUFLFSbbZSfJzkBD8R8KyZjPi8ZoMuxUyQs
SK/oLQYN/oo8TICK0XJXOvIZEtOcf5dQkVtZ5hk2C4BVXnYZlnhcoBDwr3f55N4u
K10wM+/3HLm+AvsFx9KFI688OVl8IapOI4hSe2R/XqvMnPjM6g8JgY1aPnHYMhBW
KVy3GbU7d+S//lwo2CAZyalzXtQ0lJbIfQiFpZPuDb/O4SIOqep3Q89htkzZk/nD
MVt5i5jEplwpV5o1FAav4MM5mZYeOkiLCyzs4MQn2V2tWzuHvMXHp70F7E6eewQ/
d7L92aHahP3s8x0PJbV54QXBWcmQvr2Qc9CfvFggDMuTmhps/aAZQXpIvTyEbGDt
tppLcf1Pd3A5lAHAgQnI/6Aot7c930QeNAwtanN6E6aCfCCnSVim/wFsnZQiNCRJ
+4ewfIQggfSMny6A5qp9CFI5/QJ1huhOcCjfiJZM8cNb7uxq+95nGN0o1KtaLrdK
7T38xhYBra/zIegXoNCSMpMsmvjsek2tixH5LXwqJFM8coE4BQrfH9NlDqDTYwOb
Uihg3dTC9HAaisSgUzQb6TeVK4qIkpaAdovYqSkAE2b40+CZZY0qO3U85IwbdIxE
TQg9LINScryFVqPv1xh4BaNK0oK4sHCykWMXtwJll+GkTWpRXC4qREPaxeg/2ajH
jP6eFstpxKtfoMrNPgFep/vDLaU66Rl0DDq6BV7K0LCsqGjgxGKsf9DSQIH5VWdD
Dn/vtbAmXkB7D3MARtnXNJ1uNCwEvwzz1xZA8EGiMRvPvfQSuzVhuZIvDOzWwsgq
6a6nUZahe5qFmpkD9n70QOiviNr2V3OPsqjkUH7KFd8nVUn3ngYGEKPEbJzGLSaz
cFD8XwmmYmn+76s28ShcjaGP/vrXWeKsp869leOJHT1I1wt4shR6sOq7wCq6mQGO
nscF9zTr2UDPfudtwHkeKgUPJwbOYc0OmJHk67LM8jHsFlR00IX9ACbHKqdAfhAA
3mpsG/yoVkXKhqmL4NiIoyindlxRbJDJLEsJxBK5wbVdS2K1DM1FwfwMCFCvKccA
GrCaSGnem54zimpsPrugzGIaUhlnRwkxV7wOn+S0V4ScteE3k6AgRINVuqQlPZFe
j2ak/AWwv8jiXzir9QZOtAYQlDFUS6WU3Heq+9JD+9ZHl+ZfALH0rwCOBxd0omlL
XAC+zJzLpG484fEKGZzh7JK7wuTozWsoO/bGKxVHRXnWkBdvUssMlSAi/iPxNH6S
p/O5AR4Kur4yo0IQkER2rC6Q+zIEeLw3nIvLZ2DPFUaWrpfgSSBkZKMJ8SmU78nY
JsL1Bk/5BHJjeHAGDjD0MtMfS6pTuxXPjZ3h9OK5EhZJTVSB9c3LhFDFfjlJ9BaC
+qwUz4Ox6NBwZUFo99pZ1i+fFITU76MpdcBnOJ/ugv6TJQ9v9dHXFLdtrSr/TTZe
5eU75c69HSDPZhoNiE4OlluuHaX+TxGrW3pVnGwbj9dqcnYhyUs06jK276iAQUGl
hBFbTBsQ9ei7c6bgSV6J4MFFH/KW/lOcKxiO5LjBc/xlWiCx6w45/Pn8KtPccvy4
b7hQ+sSZQzKGWgd1TOw6VWgBslCKtAlpVn7djbXgTKQ5M2IEQnLY3lOQTwMwZwow
2ZS1b3YSj+tvBquYhcRSu23heUk9cCMYFLYjbzH1SbU4aBGdReXPfqk3zHObrw2C
jfA2iL77MgqixXUZBdq/EXsmrTYIuKFGmqpPuXLuYaXisDIG4oEFgBkV9W7eHTys
u4xfjAIkAhczfUHhDXyr0V787FtUt5r33MXC+mr7c9xcnRIc0mx5lKY8nnxZVzSK
gES9l3JbFZsnaxF2sG6lysSF+uhX7luAkfFTecO8D4z1ELkK7U/CqBTLvQtgvOpZ
TV/u8/E+KmFI3tp+bL7lSht0YkwXmitsRIdxyrnnPBC/mhS0WVMe685XXuSKkJZI
b6kTfqsZOq1Thrg04s346LZTWyLAoWm2RdXIUBzCvaK07wvE/0iwg4KccRUD1kDN
4GXhDLZjR023qkuHOVLm9fHQD6qfgLU5nspSvefUW294qVRM0gc9upTpEX+dylfA
CPfyp0p1tiqDwOnErQPxIRtbrl/C9+uMFY4T0hbRyXzExOvyHb9qKpa105XWgrRu
Y/4bgMRkjlIO+IJtERpWO/WbzYCvF1As4oq8XfpqiVhhl2T5U51jFeU9VjayU+89
1JdbApmEkc+zH6+gCCPxudZxpsROA1swqss4jKu6ygsvMl50zAar/mqb7aoSZs4t
aYWGBBWsNBXg7Qt3+CqOa6OrqWvdJ9jKFfPefWUiIMkmc1z661NrrDgb68urU5Hq
RLicmnp+BCZxCP5ZcDPmviHY5E8sW4oDbxe9I9U3mm4vcMm8Dkm0+u+XLU9AL47v
3wWVJKd4JA6Npxm0ynw5YDV8XRtVWQoLpvpo7Oj6OMK6dMFvdJpg9HrxwrXK4fE3
ieyF6mMf4p0qUsKhDbBD/Nf7qNrQGRaUwSep3AvhsNsYh0mB5SylwDTghRk9PrG0
jnBnYqpTAYJ1XtbGX57yF5kXtwrmH89Dz/IcqkClkA/et6KJO/c6bXjBYDSZcfFr
U0LrMpKTMqmgKjyyu3gnXqGV6prZR9g3tH8XYPQf317cQeFOnph0V5cD4fytrk/S
sv9LceaOAHN4BZE14pk/P+3ycuXsG0/8ZKbhk+kDliJpEkGbPvYMMmXKqZa7D9Jp
0tow3qMpVuy6SmKg6xrGs49dCaE3Y1rjV61vFWXnOvZsHQZKtRpEygXNbthCM4vX
DRAOdeUTCqVWGGUgSw4+UMmyMtam161JUlFgGxjhNAstSFOqS5MznyklCeH1/Zvg
2xJjswh0pEMYMYhtLw6DzOlyzIl4xNqmEvScKZVKPhjnVdA/6bCPzlApEdreWVL/
8jOchbuEWz+RsFVwVwCjEv6/cgH3bjN0jPFRf1SRZgnpV/pZw7rRbxmwYfN/dU+B
jn1Wwbv5WovuOQbT/WGb9/tdEMn19t7QoC8qyt4Eywq+IhQjVQCU8OyLdq9e/7Al
4GcVCnMO3cIMaoNJpcfTerM928c7bCEImldp29HX8d5w0tKMbm+TxLUb5a0NaiYk
Bb8B2cO4ng2g6Xj7KbBrlscxP0xHAzCvK6Uf+M3ZHtAcQkfN/dZk111wP6SLNc8Q
r9I1TLHf+7eFr2VtZug4w58URLLameo4Ah4hOkQNwROZRhOa1NbXQLm4s5/uXzrr
NWDo76sXRxzQIfz/RJUFIV78yq+2v6ku8TQDynwYK3ZtVJW38VG4d1OEsxV7MGHS
Nnj/Gdi/8ThgGdJ0aK1k4f03gRnq/teibJRtEF4t/sQogJYO2BBzcYS4LOhIQXL3
eb/46ZyW9aBV0iW7xwp3Uj/7Apn4LW+1x2h881E6dUS6T6+8y9cA8glXch9JniV5
DDlYbhx/3N2n1VDfFiM5IV6jvSDfVzSHcad85ohQnuCt2CSLjA6Hw7EGteKdwDuM
5TBjaeDRcB+Ze1fPs/CKPCRUnQuQ8yvnrNudHrvzNBGbxK+bJOnD1YDsPk2DbJvV
nZMpYa9UoU9QUldgf5f4DUnQdxIqYuucD9VrhajzZbRKb8o3gWnun0T3V2yKJjua
KtySEENmSsdIGJ9p69Az9ej8e+EfSWfcUeF6ztnJ9J/IHt/lAvDiBq2XlMzjI80d
JGfu0EmtFOKa+5lntztBBROhXemv9IR9CRE3+QNFdp+U5yU6qeaXVxnv+pcnln8C
uIgEeh1OSTCU7iLfLhYHo2K6t0qtiliGSbwx0RVsFK4UfIxrDHKbtuBCIpJddPVX
pOYIX0sBJ2fL9oIStXHoCtG+CXk5tXoFeYTt5E3yMUlSuozdOQ2vEWpS32FPVx+t
CM0geYo38u2dbCIN3YtE5b0Sq/YaGgjoZkaxllD6W8sz1pj6pfi4q1iBHAf9UrGE
YcdL21JVoMlY3thmbOcPrPLrNsubryOUS5xOGLXmHwPdAq7o2x3EExUYuKeRBaFX
K4wXfFrbKOrsdXgSvVFV+u/7xjObTW09AUlh9pF1hM2EoN9ZQ3ftZRZZSKugTOzc
IyUR4RTrHCPTdd5qndspB8PRkHWLKIbteImjjvZd5MnFbFy3DaA+gIXT10Q2BORd
0VrCE3EwtWzvrfk/z5j1+zD5DSPQBcT3PqyEdL3oJJC/it3v6uYruJrUIKxu3h7F
278iraXhsXCrqNTrCdtED+cszW3L0RIJl/TA9UdBAjwFsy/jjFQJeSZgFQNqH6+R
6+udt2uO0d5yQd8reL9CefdjoqXv8JyXPBot2LTAfGAzu+xUUF7lMo+AcdKoXkLr
4WdUHkwdcu2/lxC9KJe6fPd3OjnfyNrrpUMeB5+Nm+RVzJ6W04SyhLV9vH4hDnU2
g8SZhrkL2bR+ER+UN+44baX+GdDAsmaeZIvYzy/qatRMxbOErbSzcvQV7sSvKdIJ
lq20Y96OyRwPOLJZMvwne/lHd//LZiTHl8STTIIJPCTuLRVlE+nIXsCbf5wgD34B
QTelGwhsGbpW1m0gGySBjCP6M7pxos5DMu2NQ+dgiIUJ6a4fElVJWqOC9mf6S8fW
v30oc7W4YmlvfZEyOgkEmFbsZzil+6iL1L7I3xO1KOzyZ6n1ut4PwSIUvDzwpUJT
9s4KSyKCuoPQIJXQ7ssgnzPZRLMwljsoR32TVLG4pN+H4ElQVjmDiQCdL/wx2xBJ
P7wLscDzAx9MyOkWJF2V1EuD37c/8QIeVy8zbsq/x5G1PRAWmyYSzD+Iqht3iB6Z
x50DF579Ns7egW5qiLLp+iyZvoKdyqyH8v6y3YCh92FguBj1PoJfklyVI8XMe64t
2S/+wFN9JTKx4LNnvA1IYRm3jmidq+rggOyORYp8A7O8qnCnOHqbjgd4klBWG1j2
xS9dnY78f2V140iDWMnwOzBheAsm7VgUjHuGLyQSldZD7K0toGCTtLbMAlSrYvv8
7Uxec62LJ1XcM7wsuHRSpHnunfX81UjVXYyFaLTNe8t/nDi72GXjblBEM65Ku96Y
TCTZ/Xr25GgNyOpi42dNeHwyHj2327x3FL26EVTvvxEXQyhS7y5Xl6rjnkpoSJ7f
GoopzU0OdcSY/ZrXhqXh0Ii2iQ+Qr4dpUyrVVgWftVgHGe5m2QqOc+S3DympQ3AY
wsDVsP9AGwDgVfDjXQJbQT6wEzanDeoTunV1XjSbEqq29rPX7OfEsBakVLc+RjS4
1Efu80eFqfi2zShndG8o7gdyUjlmX1o8p3//kbNm/Az4n4aZpy/XzSV4jX8CYy+8
8IGAnDobzFist09ggqfeaIl3QWA+tLEUrAsCzSL9PGM9863ziE9oP7+KWo/r8Tjw
m/XTZU2Jyj4cRPlR6pMNNqLEITeCt7pk/ptDiGFIJZo7s834nFuBx2IO4j1zyzkk
YkZZN+1BlMQXfYTo+zToEQWeEGH/Fr1PvRIKDp9qhoGjjaWhlhXJ8FdVjdbi1JhI
1Cuoo5E1pTkh9T7LWIflWpy7hkjFJEXeBXbug9IySl0EE4WC+TJpDOLyY61nj9gi
oA870q2dh3utG4cxmnuy0nECWVbbwP8zvO6HbjhIRHtmINq1MZZa8W9EM2B9QiHk
gimxlY/CJIV3mHj3uWTYtA86TWW0nAGxgz6cx3OJR8/4jOsBFibKnhIF0htDvhGo
vpXBgKct3X5jc8MjcmkwDQcXx9HkFxWmXXeEAg1Fr/M9qSJ3Ly3gAYu9gKlC6e98
5l0lGZ/GLMyQCdVOKxIRInywM7nKvbqUoodWlUmvb2JsTPcHwdCFiBz0jkn6KCmN
wzo/We8p3CrZ4v78e1N4OEqzCBRP/nCL8tctd/qP8QXJef2lCJLRgpLU82m121jv
UR+3MNRbyOdyTs3N/hixymgoTWQvdtkX64s/4ZVxZn+8a/gvrRnENr2/Z3OoF027
OogRLWG/chtyg+HF7/J7+XvNMNFhwSgPAr1q8mXxAZ9b+1bBYZC2EvDa1cALcfxc
RNtHyS/gqwleQ3dw0kVLcieBow3zhaHTtQitCgZ9n18CEo3uCvYc4CvCWaQVpPis
z/mCjTVbKzVjmRfEi0vqAqqXdT55/yBe2L5JcxpbTXd63Y1Xv+/G+CNZZ+9i4mYT
WKXMvcF75M9gALhxnnLQHhKWuB3UQMYrLFwih+BQWAkCXkYqJ8TyGIdyEcI1twSe
GcaMHNgD9z9AM0UL6geUPkUpz07qgjMNLKf1NB4smaPGbhYKaAep+Sslr4sUOmO0
FF20iwRXHy8Cfk/FAC2k7wLgsYwkQk+JRuXZy+keOV62V0/HULSMpsBjDKVtCDtI
oVE3aKLsMYMaD8CQXA4TUdW56zgLtzvTOhc/kn5FH6DS+9+UQEjxFZsQ92OayuoZ
AT9tOSfwLM1n93HdJk7snfl7ACuIvizYrv57ANP06LIGzcZzUCdLw5nhZUxaM5im
2FNtj5cyCMMxcKloVCo6wsyV+We36Ykk9owk8alUO8roxxMRe5p1qcXz1ZCPn3zH
G/Cg1zDpRdxMFkunS+KUkICFq9s/ptlCzzgy1juTrKFZAHmNmojrJaRftvLVNmZB
zCWzGdoTYJdO2ZKIiKyjmETx5N7kwUQGwBHYyE42ywS/XMJ4tJJxisQlApuZTLuW
vmqYsJBkU4pzGL2wj+0v82thCPrUt5Px8swSaavZwhjTYue1L/AqwaH7S5mhsu2u
8ckqcnB599P/ZAtmBVjphRCQMJyRcVJWRQVfPagOJmlRZ7IZvvJn/7dL8AMPNoN1
5heSOxArOKfc7zhBz9Nftt44NzGpLQnmVCdEdQP2TH7W/efdibNLG0nZQfmVrqhK
JY0ZG1IBAUaUnoXqYYtjFKfCrLfl1WYKUXvK7wecSo8eCKOwg8aSk+o3miD0MPCh
blqIxa+HqIAlBWArdiL3QY1xbW1OT4FjSS2uTDNAhuEZ149OuFC4Yiq/I+JhzOEh
a/9hSwSEwhq49wmgTR2buPZlNe2rWO/fy9h9uhLSzcE/+a/kAWMnSoDuWPhH4qUl
6fFGnaXhhGHZ7Kt9hxHcHSBgdAmmU4f06Cz5oXgbXn+dMDUejxs+3T7cH74Dwhie
No997ZwH9r49UPCdrp8HWuvxzw1R8b5U5pVrcUPolN2ZkR/4XRFbsoByMDIFNUcP
tACzRuv31fJhMZvcmy1/SPoh9dV8Sdud9FxSIcz4SkEtDu3UyINUxD2QXqV0MYm+
sxHLTp5BN7w7Ug1pcM4NtDVqY8VeOU5i6SgWkhZdo/KY39kgGItI7s0TmE3wkjsL
/bAFGqyqx0v8uRyVdgkTga5vcJaWGjwRYoMKlgGumzUqvjPkpbbgyNkx02ESIpO4
GvlPHTwf9JmZ9AB7sED0yKwQMpiQnxkQCVMczeh2+19aNfsU/hugkpRkCo+yVFFw
qdFt9K7funJvbEtMxnCNM8qO2pFAc0xJ3w1CUYHmwL4OKSJKLV9KjbgbZ8/jj3Bq
SLojZX4Uu3m6Yt238VU7RPWvv+clPqkFaVY+kTiW/9z7MjPhKJErJhvSmdltPZ9U
0rx14v4YpxxCTOxR1Hy1wO8cPjK/rKclxHqXWQm6U08+O3/vqWza72uAUMyItPnt
oWcmIu7Vwz6Df4hxbJ+TYzwonMxHKjGIghiM5rohQEHwSkSSowcVonfzxtT36bs1
RfnhmiYASFBkoU7ahlUWUUH3SOGyXbNeIdW4CWKPXcaa5sxrTL69C9WvFnrpsNwf
4TzCXjKP4gcywGRye/aHJL4wkVw5y3kUsP/if0vYLxq2AbmzWILvJgWBhEiAl58E
BORYmO3ofESKa+TCTw4LTkh9efkfSZ9bUe1MAYK1/XcvYR8AJ5kptOpDUY/I/Dx4
8NpvtXa87xcRrHAteXszeW8/tq9RjsULLnUCF4cDKku08gOjNuDhETTSWoet9euF
MjnsUVhUUm8+LuZL3Wnkvc8/PwuegguVd4w8yoiNbZPmB6e+W1nwP2w8CV5pqTOF
UGVAo6FlS2wbOPFKRsArS9x+6sPZiHaBcTHzDe/3lbBgIK/SH+2lgrKPAUF6HA9d
0h95jUUJPnYXh8A8+px5Rg1+t44P0igTz13bUcm5DrDsFrx/M2y60n8mBU4Tdn97
Vd4sKOJqxeKBhBo0pwPLgQvTAndJK9tM34LW09U6c2MuwMvpe4sSgxqwPR2aqUb6
P8pK9COjODjjFg1PoXkgTvzoP7S8gxJUbuV2YUQ3Gd/IUL7DKEHy0qVeGlNKfcuh
AVYH0+fTFpnXSKszKLsPU3u6PO+msoRsMQfOCKVD8zBogL7Pl4upwAR1dqwNbxeC
Ti7vtwpt6DsqAWOP6lNT/8cwu4ASuNhqHAHaAXn4hc/m0+KlvtwLQHa3VAY3aE4k
yrhNUOp/0/Uf7NMZI9yYbML13DRvj8L5k/lNr2DcVXtHPGR6mew1yvxpJ+cooqNP
EHnH0MTUhSYpLZUYZJgEWT92wln5VhNf+/EhQU98NPSI6EmV0TOCrmERvDTZ89B9
iObbak0iFpRYmo3CoHe54Y11gcDUN5SPDk6BQCvOcLvVBc2hFJ5VpQa9AOVRsLWv
2z1BbwPR6We48FmAk8U95xH8wUIZ92F1XCv0tSprcoPnvWFuRsYk7tcrXxeiiztW
GMTbN5vuJaULj9FrrKgjvJ/tp81n7uTf9Vb1pWgRPtGPa3XCrAxlV3HT3P+lQYJN
E7oOm3xrYFcwKIU2DvABoQJ7gJ48NO0eKNm9uWfY8VYtUJ0d5icJbwQOgb03D0Qv
hEmjYcNWMKLKpvFa4ps0+DS/jMtxP99uAFrYGb3gOtZBrHKDPCKKAHFWGHLkLK2n
hNZoFZiN35MW4QTi9q6NtmoLGn6dWsxwuXuUf0ROLzObPaH5OQBqTxp1gNvYOeV2
4EayIn5Z+ehlE7xtqoldC0kb+eynCJ6oCH/urur0/4xSKLNE//CE3mvkpH4qhkc8
xQqwPxJemiRs4l0de+NwsSMc2gnLTQvkbFpX6xFIEm/TfQWiPFPFOcyEvGHE90CP
C/RI1ktM92ezgIhXtFmNRJ6xWYveuIRnzIvP6jJtsmro6DaEhB2UwYdqRWDDuX6D
06oyFMvQCu4ZNBS5QPwzesoxx2tghLc5teMGmRrb0O7iQeK64v2r3fhYiL12ZSZU
ImM5iF61efdc5gzqyNoZqYVyrlbMqNqHL7wqk0mfpW6qOMXeyZ8JomDYdt0BkcIP
iBnRll5wzTX4rqz8sJlaO4MaqbVyKmSGmhsl6SIyBmSKPHMthTt731TSukraS/+1
MtAkVe2cYakjXCFZ5SdfJ7WlMmkD0cvSyfj6wSIEMmbIuo5ubaQ/LuNSfHIjFAT9
6FgYapRRqlVhZoO3CGL2TR5vM/lScToMeyjM+65XfFsr+veczjzZPL16T2ttAAcI
TFF4WAHHHcJVgyxAUgP6xWXciM/2eKmFYDqMi7icPZcZ0OX3UEr6FAZYI5ZWfkse
o22a72KYz7iAgFqiOeTTJ15r5P69h+//FlI1Gl7xM9k3vThYOp9uHReAb2PYyK3b
PBTZ+ek8PD1AmEN3ajk9gbOBHdl58Ya9aCXw6nanBa1hYWZFZ3sLsFTPk0Pscc72
Mf39acjFSTBJvJVkSNQzjvgixvpoX+B3C9mXgWwCwwm+GkinxrX07kNrD1Sw1V+w
wRY4uBc8RIUJXNHAXIzni1/Rq8ieg/7gLIRLH72Up4TIvXpEnunfMMkfI+GeD184
2VYIkLaI3A5o4IZ1+OfT0jvdslNK1F7mjJVB5Z2AyZtfazNwx95S1pCtKD3hUJNP
ntPWwxldP0sDZc28l/YJQQfY8iMUBUBcA/W1rg8DhZBfK4vxOiDwABHhR5cPr8Ra
aQ35IXrhmxpLGuyTkkSvg3ETIbYvPh5efA+yGiZK4sqyBnj/00y3Ru+BHjg3zFtb
ei0OXjmg/j3Eq/meMgUDEew15phUCqVOUIugixdeH4MiKfdzXU2c6I6tvziAJ5xI
erBGa/09jpMHUxeR2slKVQYBUie+SRskj7HlfkgbBibCuIqKQP99oPmyUUyzRbdB
5BZC77LgM67THpGd1DL1ndL0ZTiN07hIMxMRy/wt1at23opnST4Gke80wqyV2lpt
wgXkgfla5PdLr20gHwNY7Tk+RTHUgOBfJODOTSzEt5MF4d8zSdd6gFehqXl+14B4
V249H8sWHwejBj30UqUnoIazEUDSGr1TOBjKtnhBEkGFX6uTlalSfdtXNH3QhUWw
rKcRPkB9kRKuxCVlQD4kFA+z3JI0ufPvw7uZ3rCa30fDYBLbE2ecfrgRpQ9Kh3Kh
2hTsCrU7Xz7rd4vmqI/QOD0YSN2WU3QpREH5BoRscn1Vqe3l1PVM1vgwWRhO90ZZ
ps25+BzwDaiJYPkR3gQk6+bNqBA1uzCo/xnNOIqVXWSMRPGZzSJkvp+Sk4kLoYI6
86dshVQZ+pIQqtase8xq0cQ7ZS+Byxasg0+sN8F3923hfABzErWOnlGngLd8J/vl
rOPFno7hCQcsYQwadhQILFyyBw1Si0EFUm6sKokhqr6qRqb6sVk9a7Yoz3y8Un+9
CY1N+cx+UB0kcwJSlWVvjGppBYwO+BB5tyRhxGO2WZ4D1oA+/BMmt1SJV8qz1Mf6
iR3qxwEsootqSKGKM89ax4boY2ZHRWtyA6ROxWJZeG6xx/R567fWz/uwQoC0aHem
cdFFQBD2jDadVSgJA2H+HokXhlb+06P3Qk/WR00bDP4Nw0m+5LgeF5Ue+z/FP1lG
m8BAMmG4vDUMIoyFF+XdPx2vN/goGjNxZNJEA3afhSJtYWHg+oABfd9C5YagciDw
cUqdAHD5EionwePhtVdv+CHD7/6xvGIlQKDxvgU0i2P7+4eN+PAynsEjIu/GmLVw
sGtHpsHIjP9kEMEqrqupaQQjhoG4q89ooHs+DOUfpq1UhgPAHi2LBj2/j75FCoDN
vWOwIx8pW9soz2dGb3Gv6WPJ0SoQqL0qcZmhP4qpttAJ1AVIAwVnY9fZ9sfvJzTG
ZMHMQ9PzrSFnHZNqqLkxvqqsazMw/KhvKI2tpCscUK7U3dUElu2LQrPnGgevBUDy
OX1RiooioBvFyeZlPai7DvfSmwvPC8XTM9O2moB6eJH8klTdTWjbTBWyPjmFMJKn
Xxv972Nv0Id0TV4PYK4VKwcWO3RI5winecf2ewXiMpN8fampMcX4Z8EKWaoFXx61
x4E6zi+RNv8Nooq7ClmAMsr4AmOd7EKsGAzC3oB8LQjSruTDwkUw4h/zf44cDJKq
z9hACXKzx9tATOnpVO/dXB7rZJ9RGXmDyG+wMjtTasfNttq7ejJGCI+RjELBQ8+/
fjYjDCUNBTJmc4dOzUJkbxy6QLhQfhJyUu/5YBJB5SYkSs/R/SOtztWNwJUSQ+lp
CYlQnxEX0if3jYY6HxiIrVMZGUTRoeclUx19Foglzz7JxJKY55Z25qvP59NCexZx
l+chOLCL+eNJSFySI+sn56nKkXrXbfeWIe9ULcmHmw83KW/JLJ6UJjQmU19Xy6op
O5d9J7MLlIC6jzk9KoLCyFnSq9huVkOSoU6DuSlnD63h55z2ruUSXXd1XXBPgkcL
QrjaUbxIAkRJ7TCOnbFv1T3iNZ7NfMceexC/Fo9INnVJChKagcCnDyvH26ExnAV7
5HpdtoFvuj/6Hix/D/RAEhYelabruw1MSfcR65KdeEIRHArzQr98Q67YIqV195wk
Hxwk6Si2tbO1+a6j6uQYwZycMEDph7GxEZfFAdq71u2aVTb/4V21DOxa+K5wPYiX
NiSedG/3/9dAmGXweh6cE7q/RIUcZFRNaxVi0jOLrvgiCiWL3Jk6B3Ds66FWi2P9
YPJDfal2a8eesKYEQBYgishdQLw0uuPtXBV59ggJf0RfVbQwgwr1ePlRTMRxg652
yq0qWMtdZLt9P5ZsLKB9bKlymdNi0SW8VpkkKsUXVhq1brEmfwN4IVCuWZo8o+gw
I+P/Q0flvrK3xsDvbRz465fB2M9EZ/dlz/2i0bFzwZFVyPJ29VREnKjU6ZZO6ioD
h0WuhMrAy22Ikh6JPwN7sTJzTeXnCuqJkZKXXb5uYiOxek2TYpRn/MnWoyDulkqN
1Ve+PQja27vJUJDXgET181RHqAV8dSJS0pq6dlOAAYtXIl8hVUVAO2RBc/J1Tx6q
6DOwImRdd+0Vb488KijLPRiTShXyq2GswQguK8y8XCV4vIcjP0m74bKXJeMt3RfK
Q2HCGYmgbu2qaeC0eiU5N3cz+gFnb8e1TLJtLztQz5Pf35OiKijyHm1i6wfpi2te
LAoivvnosDpIkTfwuLSSj47bFFH6ztO3CxnXAcTZlcVeBLFFhpQRFq8qsZJPbOGQ
fYBvEBKIRWZCzmohxy/7SvkwcT8Hvfu+YD9oxkAtZ75eZNhjUkXCLafyy1FkdbVC
gYPZLV7q9k2gfClYsKwPRHunQJ4hxviP2V2r1fOFz6PbwU9oi3+SrpVMepzKDjCp
cUdl5B9j6UOBN5B3NWfbJsrMgjUqeNYKpv2+VbcM7EzH5d8MK0ML7xpochLfwcAD
ru7hXhC92zHudc/Y3E8P8SSjvssDW2w9BjaGZlWtnQdLEAeJyJQV7IqMA50IHJgf
/eYmOkMlNruzfWiHQq5YBNdH/HHYckM1f4dxD5sbnlCxFlxZmKuIjHFnSw/vVIR1
e+Wt3AJ49j7kBYpXbTbuZwSX6+aFskob3fEBSXndif7133YsEbcp4eYQmNEmvwXN
buCywmbbsjtVeuQQU++2Ft/5bSagK0Hl1VmSahkp8A93C81PjXUYMKB/HuSIFJDJ
2vZQuktdhwlKZKVf3Q2zLa+bCdd1/ViWh16bhW/lFcip/9kQDNGUQ0UbIyacQII1
spZDhz8EtH6++Zf9n6N/5kc1qKTtTE33nXjBHpOWL5ctojY4gb+AD9J1LttsXSrM
b19zLU92+FOHhmnam2kMQSz6fNQt291J3bbuA6XkiCebxX79OZSb8pgqDaLQUvJq
F7gjD9yyGFrqAK9QUCsS5FMjrMSc4G6FG9OdvgIStlkpTIai4Xs68PAWSRWhVDui
dr3m9STVrqVB4GfE6OJarwzd5TGYuL4wmV3ziYHN239QRzlRlz90mOWnyxbK3qM+
tbzUDcJUYEoREba9ss1h8y8B6GiLE5FpyxTda1diGdpi3Puj+Y4qWXI/bMi/uz2J
sZIKv/NgoSXNBpi5j0N7aQbjsxQVCK5XzhCLQpuPH7ayePnlHVeykh56pAuepj6h
KsF0vVI7Gbhqsa1zqQx7gnjnvpjSXnVpPzbpQ/z1QmnxgHlIZ5y8hiHtqfpuOcIT
yBkaxThUV0PrMTMsi5RGdeYkUArBbrvwHBQbKAWt0cijpmBDHy7nlzVUkHVPeiLG
FaGexexP+/oHE26id/i7vv6cMKxHaIiOr50w64TSTganUPGbVcXjb8zJb7BVA5QB
2Wsg8I3YzV+GKPxK75dTlw5hu8qwHmq2g+O/Y8wNfq7SQMAjxsdCrqrkJ9GmUqnP
Fhtaxq0s0NE+mqsepVOCqr9VqTH2/GC04sRHg255dqNnBdn8I8OOG0Gg1NuzsNyh
xDo+ozpn9xg8kVz72EK2OpSXOjf51ZVSpI1Kg2fzAgIGX+H0tiXhLePWt5S2eN0d
TkW/SjH8gZAKbkfGHj8e8ske9x/nQQhBy6ulnFeAnT4gd859KGj8Amen59+K1uIx
T2vMJ9sklUR8L57TvHmjnWYNJBSKnDUZYzkArmM8UNWb0FPcx4O02ey5alRwMIEO
IHCXSMoKhXLYZC3p73mrDJJ5aVHnC8LeDfFbLfvPKgXvelmUpOoroOlyWlnzOzXh
iynoDp2NB5AYzJ+of53Lq1Ze0g0/I3uWR1eqxf2CIYnbWkM4uFwV+2qDGMa4n0FQ
N6joCU63FPnprJnf0DzOudZ84nxg08GBSzaI+PFDdgyBS96EU005G2aVRPxMCCPh
nPhQSiuIOnSUFzhcogv54amPt4+/7Eexe8tOHe3Ghy72lrQgF0JsSwVhBkIDrtGS
O1xhNzc3+z0EDLueYxugIt5XGuhGcVF5HvGJtT/Myr0SW69zkJSc8CWlEpOk9oHT
UJgZKZ8t32Ef79iV0fcUK4r8h55Dm2hy57kU7DtHJfr+C6543ZxXAmPXIrDPlWyU
wQQlaJoBEtDxbD1WeDOj/kz9+nPVK58fHUo6+ohGtn0kza+5K1J0ok7yFodF+TCX
3AP1ABcJS7r7UuukrYmpf1gNnvF2axFjWcESD/+p8Dpb/1CsYDgaLlm8i+xBJ3Zu
Ras4P/xfGL15vgGxHj4rqd3XnU4BiknjFiYePZ/Reukns0S0pqvSI8v2VhGmI/Yw
NtVULJGunQyQ1MwolZSqvQyFcPGQLzM4Zd0hVbMR+A+h9/IoYQBmgtwUwzt1OkPF
Q/xqUgbXVy0hbtrN+YUGT/Lf6Qju7xIgSboAkV/65eJGnC+S43itgBpfcPKg5hgr
QW/BXqu6FC+waxzGh1nFXx5eVbD88OhQJDRpgS+6EicWSxHrG1I6O2iqikdHs5lL
fb5CUjNF+xWndXHxq3eQMegmCx3JhOwWzq4GGDT6KDAAUIYahGvFc1J1LBpmlibW
m4hrIwBUyKlhC7bdp84IpigIksq9nkreieeIzhnLe5gTI4cFGO7pNyNNeK/DWdz+
tg2K5ftJxdiQ7Ts3IqQRwfWg3uL+mrwXfSn0a4x7ANJ3KvqN8YOuLdUfzor8pRrk
i8Qk4UI3pLQJvyhfmUTBugNl/pg9gBFoUWOduUOts9Jm9YLTnRx6RtRwKMyhOXyT
wgrsk4UXJmaaBviQlJ3OginRatU349P2MoBoIpzECTc+9DGF/9vLqx74144l16VX
R10Fbk4z20PbBByUZZJN0Q/3izn1pYzM0/SkxEZfpzD6KrsuSjrIsQQ8jm1yNTmA
BFaDAkYkIFY7NZpdu22rFfhWqzul7CqX+LXYGeGv/HWe3VSVlhcBVYgk/e64Z6lc
Ly11fp6pK8ubm4iA5YpgjoE0EeFsIpx/TVD1zHzDwFdlP2JeXkY+eEBXPqdbSUao
8fKSlzXtrH72ZBt1PLDzmDlYSzAPmp5gdUf0XtzO8NFQfvmPRbVBUcOJnXbyRWrM
gr3yv20hUgDZjYupRqUeLc71Qrc8OWGF/fFQ2Dc6XTAQl3oQTNLXh1yWQGp/A+2B
pDNpZjr47voyt1l5pWYDYV3IA9W8T0F9NJXpowpgPftl4FWsN42AWlTkbyA02AoK
HsHabc4RgyXak9rq91N4wfx0BNOla4WJxhF8Go8SGcFbLZfldrhn21V4wqf3AVbI
+ECW784L2PDyisUfL7ISdFfHkqn7Ps7wDtz6pNL7wPK4qsjYNDhXl4nu+1eTpyPD
iEm0LU/BM43pc6gJSsjCjQ/8LySFzSUA+VpZzYA9nk8Gs478zDoRYfuRg2eKvD/f
KW2mKFZVduNxwuSDm+u6GVYp2DMAfJBafwQBJDTbZRpONhJ0wOWXWntvpEXenNPi
+BXMsgFmnkP7kyJn2WHQ0ycU3aRfYpCEiRE/fg5cW5ZAUSeU090aDpUi/pLrqFyc
6IOxnSLBdoTqE6GH7xfim1Ibg9WWxEQ6BxZK+n6nmo1s+OVljcEcjiNJRA0EMiky
JufUedrgNVPs5TizYjbpkTKaSFfkcD8oj8+rhZ7JCGoTRVwRw2q+drxS3i80tjTs
9Fanb4P6Zw2s01E46uk8quKlu+Kwdftg6XX3g+QUu5tF2JrLQPsEgsey08MKbssh
SQPCc+Vq5nw2yEiSQr2wi6sek9VCkwCfpZlu8c4ma4CbsHtafHb5xbriZjLOhlbJ
r0v8uRGLU9UuJ3CHI1il1+Gn3ltp73cfBfFBOvElm0Fy0wGqhX7RzqZ3Rn3N+ifK
EfQcq++LObNtkqIN8nDopq4fOnxWnknm3UGOHx3pYuQjM/HdyMzHYicb5lbXs7I/
uL8Z91hhILoPNKu5WS4HB5ePsYeM8LNJCD+CQ/522krv+CZuRWvVRiA1vinWNXCF
OsKlXZTZ2dD86GRsg4VOidSBSS8rG/XK18GFzY2oPx+gqLefZmDUWH2iFJ0/6iWZ
pjkKL0t9bTbMA2up1v1duPlgZtKubpOil2B5g2p22N3qzQRYO/2EUX8Lhv2lK7PR
pxOTIYahn74Pm52vaOajSVem5e5WGncqc6iwWs/5BZFpNDtBJIpbhx9Vr+BoLzEG
VXZ1DiY+Jjp5Rf2YztMcZgHlhVyw5oRoUefMbTxxn+r9DmyUjKWH2nfMHBfZr7ID
B/rEnZN1IM1Dzb4vl174iE/RL/ihS8nsfaVhbpA5JK1+/NIImB608uHIvjn8wd/F
qrGeP2KvB8XiCdWWBIHPz5eiDjpDO37eWd3TGtQdEbl8rV1dDKey31uwGrZLh3B+
mD+O7ZBTajzrDUNTETuPKXTnbD8D1P+FqFDM10RaGa9p1iVjmpF+pOnHeBb3/7Nx
w4ZF94JMjKAKBCVJP+E9wh7sULD0K0DxfZ/ERiZZ0zxERg0OTD8YSAG6gLL5b6KG
AwVeFwNbsq6uuZz9u1KEjI1jU+zMDyj1cwStMAGHb0ruo5GfXfosJU7KTm9eQ8ju
/amiqcDZnpKMnI7yuyBAIqcpZ8sEx78zWNBvXdZGAlg40oR6ZJDyuYow5KPDfqmE
9LIXUCqDwW77BmeMAIqbqtr70daxO0E/mXObaiHVyACUVXcdcHcymVIvoNRc/HO6
Ht0UOki6OvG4uaM7q+jVswYeXRrZO/Pg5LNlSrNItgA9x5oSNO8ELd6c9Ah/DJGg
Z3QiWkzSxsuCu5xb4PcTm0PRkbYPIzgyZYKrTC3yoo4/L6Re5rb9GD/erWbtTDrJ
Krdm2k1Ivi9r15XkAGLLf6S21i+oO70plp7kJwNznxsO6SyxQnerkkUtzsYbKzBR
ObT0x7Uk9BGqXQ0BKIVXD/4WaTl7EugP/4waMkwyn1EfOmz/SVPI2MINdA489KoW
MWNkA/quMkYi8O3teuJerO3E143itIOvkXAhFTThOV09sXVnGhMH8kT2l5rFOJKH
UvonqM71jb5Gv24yjNS9nqJEuyrfkKeX/nVnkOy/ydpJ5aKatNBTEVSS5G42yQMe
zQI7e7W6H0lInjcnODZ/29K5clKzrtVFKyNBGo3Nscvm8bpJd1TMw50+kPpCDZrB
bOgMRqL21PI8vwQFrFy9rcayYgFUjUtdeEVuLEZVA3cDNTGnCt8tr9tYsRFp1ieY
umeeQB9yDCVVDIYTSzXnZHQJ/8/rwiZPR+L8/vXFRKlMgiXQRP2Dt3/uIg91gV0z
1YLjTmXhyYY65Uh+KGffL4z6gkUJWi0z0OlysCSAj53fmP/AsPAqT3Y6yhLu71zC
ji6d/2Y9EmVMy6w3MCL0QSoSp2u3nPacgMxGEki2Xn2sjwoQKgNq4e/fWOO73//h
GGf6f0roHGVDX3eeUIWGPuawnu+peEuu93Nl9u9XTrcSW4XYGMeEhUQy5qhbnKMQ
exjkc73bKRmtJoCcWZAmcrETiMr8X/O1ijvVRxGF/0oQ1XpfFl0syDOwd+btBg5t
2p9aR3kwA+YUNtwoHxRaVEycQ+NXdLp9+Oyulj8rlXL63BYVjO23gPAhJaKjD/1i
/phFrAm+nHnsX092q6383owLY4geeAtb2IpsEZrMPxyWVIdyxMAxVFPQAP28vlsg
KcLhLYMzz410oe+SEy1fV3dd7P7k34BYZsbUIBWNUUGfIfVSNx/8ZUp6N2OSqFqu
ZZXGU9Rb26bS5LUjz93LqIrjm3/EbfVGhFLX7jJRjJ1W3l/PlZhl0Kj4fWkPVKOX
QzrrFdSjYcqC/jjHg201VREeK6yo2M80YDWZXAogVdLW7fIlNoR0tlP59scANqqS
vWGEG6n47QQc2uG7lymysMVcSjMmNZusJxkfXe3cswHdClC/rlpZm0Vjz400E4tD
uomjOC9I7Kc2G7XAFXbrxJ4qJHPFZpLfM5bm+y1txcN92fpfQOOrd3wxBeP7F1ka
kCZMBGMONA1RFWkz36j18hRk46j16xk8WCqMLLkrrMqpfinpjq2AMe6nZXzwFjPZ
0jF1HQV/Evski8brYfJiHzqqWRpnHXSCQEOfk0qJHKTG61xZPn96yi24FTHH61Mx
pDfkHBrM3hZnsHvK96N8YuVO8m9xT5b7O3H+IMpbi0k/cg0NOZUFdGTm2NmVsZav
q5O6kuyerPTCAq7UNLplhxn31PSeYBUC2tTVlisExNRoNyyH4kbx1NSh5/OohCNY
m17D/j8+m+xnsRxvFvIh+gFfKIYjCCdwkn+6e+CwajtLcr0glo3Vy2YAM+fN+lyU
jB6IxXQ322ASjnHyS9Y+nSUPRNpy4BtKsqozzrjRM3NMhhdKpfj7YUPwQSdZopYf
FUhxWpd5QM9u5f/4Fww3wba2cOSuoBIkakm7o8S23Gmqeokfh/YaHm2y9u7g2w6x
qc2uqZRRBoR94GabAbYf9BLWpKkhx2k0RgLRE3ug8OsMEKaD/0DxYBjMF1Z00ueO
AFatU2/cu1ydVpUka2FUbqLGWF9FMtA+squLEDdnfskaqGFhKICfQsgvfut0KtMH
rq2G5sEFmEwDApP4LmHm6jyKEPtMeQklmYcW9CcGWgfcnQk9liskJJaeIDOnN9pS
llNmcIjENY4kFDfDE5W2UX1+hNd/6Hh66M50RaNfLDHMym2+sOv1oFdHwQc/o/Ta
foanLYsr3oBWa+8DUIAT4eimsiDTe1H2q6EWJdxS3U7/2719IvKv62bJ1xY8E+CG
oY+7MEn9uFDXWrZhrNaHiNfgzryt9g2XRmcboJEIZ9ysMixudh9CJNbLR+KKKo3s
WvwHnUs79fo5dMGRKGYGFImepAHxOGOO0I0RC678AJIBxmG1IVRa1VXDxWvrpLEq
+xSlo2Xo10eW17V1D//RT5juCkp9vsLNiH6Fg/j8E6exkmHv55Nu8yN/l9JUnBu8
14l9F6tcuGLLqd7ToZYsXSB8av08fZsTALCDKPXIaO9A+TH0FwGN8GZIfeW9Iovp
k7l5fTtEh3XXmKD7dZzu2+LXLdwTTVF0IT9mhBlVmgmOqaQvX7s/n2CN76eMXEpz
wD7Jr42yq0eHUd7vrE0wbK/GvLSaPg2odzY2j38CL7Sd8cNbwiJmmCeekMTSJe3c
0Hf1msLodqOSjoJM5DD1iVdqQVDuKEfo73jVzIK+Qgyp5az/taTbNX6Q/42IELDi
qFWqq6rGbIzOHr+O1J48gesFkj+LQFzJX+9GZbyexBlM9xZbtWinGQEfN9eq3wCe
6oCgoL3oa/4cU1nkzO0LeGJdQhsB7CGfn3M1zCUTMDBrQQ09ORd8dcmohfRQ6aHU
4JJcF7+QwhR9ZH0v50mkRHmc2YbQNCcF5k4JN7GQLum0VhA/zRmCfeUOu20fbLhx
2YG8c6NIR46o/H3nipjDV6UpnbG8yJP9xafSkSdHjg0TmQsyxCNhD2dr/FwgSIH4
xXNvEfRtSBtgqbiofE+n2EKjVu1bGwpKjysBOgIj1PYYXY8uOg41583io/z4CXB6
TG+dm4lch887u9f3vOU92N/vicrj7HMToEB5KfijhKV7x5whAzVRr0FPu8/UmJGT
+g338RPT1zLbNeRlvwAa7/CnR4zoVnA23PdIpR1m6wa94mt5gek2LYV4TVfon970
T+20Mm5lUgKDEKTLiSvel9VhCtjdZfBN3EvLqtIVwtySqbc4+MMcg1g+hoJS+hrC
Cm2+4Eek4+rpbmDeFDLrFdCV0cAK1Myl/ATPYBLfQsxeC1W7t98SAW67TcRol0r4
/Ae2bAs/Q42vV7bttwx4cMkckv7uBJdQWX1HXyaaEIXQWu95qzN4+tOJuvmjEvNz
3IyCLrSzDjOmaxndn6k9TEGPfHls4iHT51yz4QXG4ctCnMB6sXP/7TZD9KHKd3Ok
dND20X3pF81fhBSsZZHT1OeSqaZULfFZ0HdrNrKo/4l4LsuUil7MrhmKcCnB2cIo
i8HRCvBJaiHoD0RvhF8hE6fRTATb8Yiq9tJ24wWSxqAZ4AgnKDmd19VJy6O39+EV
zawC5+zTjwa4bfIP6XKdJEk0zDmE+66jN9sYQMpb72qNRoxa2pX7HNjyoks5oOo2
MtufNN4IZgLr8rNRYZOA1AIAO05DgdNzBqJEQa4FQQFXDc/Jo+pOR2nwNU1UHLTf
cF14xU1ABgaDC5y5Tn6uCVxdo9f57oDSlLf1l80bD/+cWTIdM+Fvtp2aNYIK0COk
rX+9p39V7mvkykiGC4LCIxj2DPk3JN5C7kcfV7q04pFqkbkeWOP5QlylR67uhnsd
GRBhwSOftH8tJpj1IBBq2LqVwcMtsCO691Ctq7b5Yjtn+cJ5a6oO/UqFZcxnQCKR
5TvcgLP32r+XtL0m3T/P2nc3f+qeJTnrktsNT7v6CmxJkgvw91ETreljbz1lpP6A
vbup7+g+n7vz4AAhH8hCyaXPpRgRIQef/3XOO8P7CzsCYKsqrZushhIFIu4utWhd
qctlFWTx5ucwN73Fm8ooN+jqsmx9Xu+8qHjGyQTuWAygSdCk02fzeI5M6WdwlwQ0
DUd6JJ+GS379AyGSXBww8z0uA0tkelyh8c5Fv2H1iamCRksB1lptwAjW8c+97lWV
IYxIJHIA9GkecUVh6En/xqnwDp7vDGE8Bux1V6bqveT+j4viRf0v65jOhfJA1sV2
cZtX9c9OmU5J6t5wTcCEtlE3qiiGNS0sKzPX2HCgXnkQ9iOOOPMINOjVe5SBawfv
+nrFOz51jR5R7J33aIw7RZ+R9HBObiy5xmNPYskcIMr//KK8tt9pfoj5fqT+QXUg
nUHKzQyrRsgJnyjTPPmB3tm+BRONB5BKv+jacFE5RKMDLvYKoLGDCdX+DEkFlDgb
Bhg2XAJIo21GoCdJEL38eXIz2WFFv4QdX5vNO4F9BANqi70cawcesIDDIWm+jnpl
Hum8iEYJDL/qzDuSjlWETd5sS1l/u5QSFEvwSTRbYvFHARCp7Up5RlcWoCKDdbk+
wFOesa6zRAL9rFPZzJuQhIlwlYkQ/AJiYpugr1jVQnYfXdQ1Kzi0KJA06vCGzMpu
VSX9eJCaBOrDebYMEF6Qrtd5AeaMsyDwuHG64uslpDtxcpPQP2EpZiITFFnPF1gc
CPjPWUR+3LTv4pMuTX1b3+02HeEng1PxUELKRMdH2ydj1IL3zoUCPxP3PsDQ/zGz
Rz+9AQA1OG5SFH8jDJltNl3JNvG95LJ15ztCUaqiNHTI2y0XIcNdFQxnidZsiId0
1KS2D/pLageBf7hX6Xt/nDf+qA1NbtUbYFQJu1R72qTkZ0GDAcpin6awyU5SR3FB
Tdj2y27GKRbnLkWLNJCJxRXIjRtI8711ddJ65CAVWBUTg5lISa/crRKn+T6D3AGE
2J/ggL0PtKOJJ2fNJk66E9WGW6xMPkcPyP7VN63nSbYDbLGZv4bHbad3lEC1q+A0
lkIZN5Nliuah5mtlQvzzSUku5y3o6ctBb5NB0yBa+yoDpL841u/WiRObB7iRJ1Jq
hFky0xzPGoPEl4t7MneCRd3dgDDmrncbT2hQfvJc+y9Vqcr5IFeIIm/lHuoDqcEp
wbd8BTc7pnmIzJ1QIr0X/OtqYSZdL7l4DWLNOw1HMFYMshAwtkz04Tu4OzQrCI/o
7GiQsO0zv0ScqY8A3eeupVHCbOLeIMzNW1EhDIKxFSaU+iTo+hNLBndeYMWXSuLi
RmG56vRN04Ud0EbuLEx2NgfaKxHU/iZpXIvcuCHcAVSsGoP2quuU4r1z9JftAaP3
ogfrquWuMqAtMRlsoomLfxlD3364+YJUTNkuV0sX9oSw1dpFk97lyfxv3r51r0RU
a7RIIr2vAOrLmEqzEHxKEgNSsb9r8NZxIaC7zM7ENPvL9sxUwdrzBBG0gSIR99ky
GM7ZCu5BGpp0DHEC4pMSL8+sumt0FSXXyc5uSsAEtKhLXpdYnwLIXqr1M6zgJ4ZI
eZV4EqlAygqrCuhbAgFsTu1/qV9rpilCd6V3N44Jz9ILRH6OGpWHw8RMcaoQPC21
s9pdAw334Er6nBp35SFmDBHE/CJj2wKrU/KFPk634H/lZz+8X15ygdKLPN96hFpQ
sOelDK0Y/ngvAIonkN/3hLWN3yGghlXvz/BedoVeDemSKV+kh+gGqhRD2ow6qktz
eQRbw9XSo4Z/W10jKaXDf5pkKMgzT1AejXngO2Wm7O46G7V12W6NBxK7dRh7ewbu
3kr448focjO+jBAKOUT9LS/5Fewm+ay1HvlueMCKmT+AmGakXhQOYVpzn2aGlzJ5
z6EGrJbEw826IAoFQH7IiOKpKT0qmFkHpfoGb2WjI5+6LT6Iaod2lrH0FajbLzZ2
knKcm+Z+wfu/ywm2Irvz/vHIZ7Jz2nOGZ7wqDoAXzwFkS20CXDAH3VtHs4958Y2h
om09P2WRDsGkeLfJk9blEHwmYDD2iXkXT8UrP9bmxtXgtEfB3cRqtKMMpX8LYk/S
tGA48wpv4LUIIlPsiLlGQMB2+UYHFILh+XIuoCkbtDnNLXu9/Mu2yqIh7yxt507H
oEiUDejeVNBehnr6wfZyfWBNi9UWgZ3WVSrDQdd2rfcbm39Zi+n4sb22Pz7XMOVG
4/7aoPrXHmieRsvzChUtw0X2mPIqUKpyVy5FSW414s8IFYxJBi31heZsemWTWlZ5
JZqm2b0kmIUiNjRiJiCtyXemzwuQkbIFJqzrufGaRI//J1engFJAJXqaEoilEmKa
LB1dW6OJjXnYuB6B/BVWyRgny6vN3yekGUeaGW6FOMKjdFUuM4daP1K6f/zBpWzv
em0bb2Su5vtW1uBtBFVqm7NhZTPliSQhWts2QD+guWLTORxrEMrjKQdEUk4h0pDi
7w7hRNABCVzkLr5/sIHGXVuDP2s7th3uj7KTRjv/CfBWHtBxOpaioD57J0AU63bm
7JLmaDuqCR9ns+Mvyf/wqb9+AtQKjyBGnljTKoyXU3w/JNSg26Ed7xBRokQcW3zR
PlPS9nhwhCfnar1x76mjSngXPxPBDU0GNbxcHjE8QYBzT7pyGZefNlvAvYEVyOtr
ylWIMHU504QExCZqedQyTuhjxEUh1r1P+fxVLDrYnANeIcIZ3Pa+NXu/9OQ0w0gz
CI+6tbRyBHB/BRY+NHqKwQromrvtULrhfH2xgtDYC3vkdVYAl5u2zBI6D0gemgxZ
al21YUL1hO3hnfU8S2NqZP/+I8cUR7/nsoWkIC5yX+qeTglIGRYYDsLpnrkJfxpw
wxn666R38etJJXlYiz/xuxJ2y9V8tvTGCPO1ESCzZTNbUQoEdN9SkOVDMb3ZVbnE
TvC1iutcmM3ot15zKKOpLIHwXXpKovwQU1FSb4mrdzRWTikp3753uy/VvA9bJolP
lAOMeE6oAFVryIvIVX/1D8cnbnElUdaa4BMaYAm8ZAJzxTnsVkiSp3CEkjFX++jq
ltT6bh++daa5NAYVaQ2DgF0dgMnK5gsVFszQvympf8769mRedDyKT+cMLGFUulwX
+XHVumvWxFwnRe+tblAww75UQtmou5OjrGVT0nH23HSvCQ7XWoMe5+jeK4denxvH
5ShzqIWLUf6/7cQXyiDCZgoV4v7Yl2+Tc0VyjqXdUPadvuLLcUdzsfTtka7cb6Ii
r17dhBHCHOaOQbqFFrBmZ72aTcbDyWrxvLxowZlBaXLzDwBU539MyNUDlJYhchZ5
GFhrWDJ5LS+G4WkPrtfZRjJClEKPyUsuSTaGolzpWVGqf71bN0EXDHmYDrxyapij
mZtoX11uAItXJc58hNYLQt2xAORsYePZuYHxXJlg2AIPvBGm9mzC29Jhozb0H3lI
SeDCQjia+VUEf/A4+bRd8KVrpJ00xCt6IFpfdAmj/IOr36amIs60mq5ArkKVosQq
Db22q1zk1SrXG0bkKU2hV80+5idc60FjMQCtcbZEzpTZLOd2DV+vNgRHrjYHGVnN
sRZ8A/2bXP2YLnbBlGDFcUfRuap1zM1+OGPOtNAnFYhseNhf6+cJM+KjhREQbZQr
ul+cyjXyCGUdjtrjWvRw3NEPPBP844JocKkLIAiQkci+bJLnT56XOsa0Xr1sYEQ8
i6SLxAL2B/+q/pWPLL72ygD/XS4XWge39NDZTJCh7wuz7GE9/QLD/EWLkadXspPT
7PuDSWXLDZ6i6IfQ1KAY61v6puorhocgPCFUfppxRjrgMYIGHwtmHOtBmlAJPi1E
/gliG/dYwA/zxoDkEfjCJHwHwf46Ct6gP+yuMsNtXymFn8Qn0l8gMJN6a8vrvvqz
OVpyrTqUAmm+6OmBDbeutJga8Ok0uttE2oUjd2IPgTaEQ0yb7ZvGDHT7mcqeu6jb
gWios4qu/tfnYQH7mfC2ArOXsS9+2IyWv6Q+j1LEfDgCbD2KXxHDjEMlM2snHWo4
b6bPXcNQe0Y+9LgcRdWJITV/Y/RbgSi9mr7Aa103wWJwy940RL64mRK8tb/sortc
yvLrxeyc3778C95srRVEb7IN/fCmO18Jl9ZfIlNcqKnD+gBDvzWJLLeKErXvyFOb
I1xqCvkGOimoV85CBhy+/8+ABdgpsyY0AbTc7uX/3q0PFGojJ7nQyRjPg42/Zd/e
3FbTirs6jYdOjJNfZE30b5Wbx7YH+aBhgCDguJ7IwseRDYNgndaQ3rHv2zP7R+cv
sDvKKWEgkiT50imHR+bco3n2m72eJ7Pyxdw3lfQeiaYQ0BTheObXpmJqs66LlFk+
jCLXJhgSZzTszWI25nALkflDFYoZZjTHIi5WwDtLlh1/VMuijm5+svFJ0ONifD8i
9BtHFoxka8820gkOOwdbgJyCq5OW7HjzIzQrRfNvnz4qK9+Y1bQX/6NLwYB/RHYV
01HAWZ5pWDC7EFHIOvyH6O9XGjEtTI9dHl+X0yHPPR7RsCvN11es+XJi0TznQXbw
Im2Xh/PyA+7qFcvd+36WuCLiLb7f9xyVWvI0a6ilziSDNEXVl4NmuihxUP0h3Sy1
3WBSF476gBx27ibcj4E/vN13tDd722kKwIjFFw7GoLRja3zonokr+eWGdFoyguyo
USIQ0T831wPNN97G60zB8mlIMZm4pmdlreCQu5mQP/7mcXX4YSqH1Nso3LhQrXND
oVwaL5o2vsBi5ibUoULIT9L/bqBhurK21nWW1hVy6ddjURIwDybkL/1E58ULnU3+
A3PH4JiCoS1jped/3hXlbirJdXQ1clMY83Vu9f7175m693qne2Q9ejlFSVRhKm+5
UryUKR5BC+SqHUaL9jeLq1Lv4IQY/TuPtNm+fLJL7nJNUHGJl6QnngPGLbtvut4l
dynA4xOveUAFXK9XCc0UPJL6/sLBKlsc/FW14BNWEQWBvh9CYxUwi7D/UxFs2xxV
fNSc2q6KuhCQmz9NPuQMsQhCQJHYerMQfyxMyCl4QdkkHizPi7poHl9y7074C7m6
WOmVVKJw896sIf4+lIpqLNcNaE78jOnn4+ddsFqZrRH8w/IjDEJftbwkMcu82IbI
PE1HiJ5ePJBROde2BEH0+OM+KN0mdjHU3MRWRO6vGuChHnQaWQsWw8xsSFSZe+bN
VrMj/YW8vJqArOAWmISujH0Ix557cf6IyD7VR2zIZZEt6ZnHk2q5fFMsMjoXiIQL
DIfV/6adgLN+GCMG9pJUX0r1rz8nFe6upolzePIamw/im+tVCBZfOjZnfEg0CpgI
WQTDsdA2ZgDbwMbwQ5elhQd52Io42j/aqdomSvHfLEjvHtKRUHmgWE/E2CK7c/TQ
cHo02uvKXU09RSglf7mWb1s8aJGEmeMCZbYhhg9+bjNsaEbsC4IgbFKWm5gZGTQn
C1BK8Nbs1jEK6EVlsfYWWsl8Er2puN1txLD7UvW3p4y6Xr5DuKgAaFtN1a3Vd4bi
o/NffT6EGCPL1JMG91cJ9kWB9oYx+Os4UQtWW2tv2+C13S0mcCmpLHcWCN+ciAwE
2T71DpZw6g0a9JXLSKtnC2ee7zzEwnpKa5NpO7mJEMxD133V330igBvX8/QSxOp3
F/VNQX8P1KZVb4fwL5DZWM7gYdKnXbzJ/urCXMf7FBQBTPBOOQHIVMnuUELh8hom
6KvPxEbhMsNVx5n04tV+84jRWr70xfDG9xxhMAGiYHg3lB3YbeZBt28qB2Ur+bA9
cE6Ic+xsW8Ms9AINjU5xF7U2/MS+RypOc0zej+sJAV6WSXU7Qnw7sDYZlxJB2Lq3
DJAxz0BLnWkqVq/KdviaABHl64pKskjfCTAeiTKl+S+4/Kix/gDUOnA4pT+67JoD
p8gBQA+PlGiJfl1kP22gtqMCbStgKmViXWuCbtk4ZweB5r1sAtBGpY45QLOTb2o7
PgDnpiZpWAq0dG6FgLkoCvpUuCKVf4UnpcySXwjJH0HFWWF4Yuh9E797xZnsow3U
kalWHc3V932vRRmqEsbHdQTNtClkRyOF+kf/0hlF8v/CiKBMAFX257rQFQrX8BnB
nFVnAP+EI8JsYX2mQ4AxZ1MKrV4nkWHAYSDvRHlU7XP7YJsqQhUafHPCb505iTsq
cvZ/Fml7xffkT8VaySAdjIgxInzTMEIW2bbusWlVm3ZTHVcCZuSMZeag59sJzUve
23T5rJxVfHWRBUfeZY7O4eQPXlkDULApQJdPkIggd+TWJblfCE6rIDdqw9yOoTQP
u/4NoJEPj5qDYjKSK3KtEV848Ev1uC4uvnCI+AWi3CE+08YdbSamFh8pNxutQkuJ
dtqFoWUZ7hgCFmqQ9rBOOpUkw9RtxS7k/0bRvuFqNzE/2yYVHpTTRyy1hOVK2Ong
JOTaekpf1wLzmfNjSOHRWO8JY+TMJqL1GDsAXbB47v+oLQlwA44AlOPc60HR276S
WS+94vGAE/GcRWlVFIGlyWoeNKYQbgLjrvJVPqN39M3VBo+aufmNx8E38kENBZ85
SEetqcYh4LD/mJwE3YSwbJ3sv3Vxw5nhUK1ogaqgDKYqAuMvp8T3eN1Aq1WVzrCq
Qx4nZuqS2XHdn8K6Zbe5xjT0xmNtU4v6s/yiFv7T697hGDZS4fTuh5J3ZKK+Tb1i
DfFJdYQgceBxoWGTzxU0D/uwEQ7NZyfYge6+43OXJi/LfDdMzmNBepsC/qqRBU7m
5v4j9oTUulsUOkzULgGTq1MDCcfquL+WP0wugNrPjmxakdoONTcGno5/7k7OCZ7/
/mcBJZ05W6r54+kEzuA8EaOe9upG7R/fXSEIEmjNU7NTP4KFM71HvJqqOsnmyjdV
NIhyVEzMpv7ySCTxSSGDaWxa8TEXwH+CQoqlwYiBJOVU0YeTyCDHCAG/YPjZLMok
Aj71Uw1oQ6Vh7owxuwHLYuL2V9Pgy6qIG2tOl88aD/yU82L1fk0ShOXC2DMOE5ir
HB0iXES+VftMrMl4yDjc+PQfJ7Z9E5mc0J4bo4nlmmE24TRytBm9MjELI0enQmV0
fyIE/2dZtyqt6AVrZdNoTgDOHn+ZYG5YDiPF+Jf2HX1aLxDlkD/Ds+zM0G2cmKSN
YSKAmk1vME92daRUe58kfeMxJ6yhDXe/luJErSBRv27rt8G8y0zesZFDg8EvQyIH
UAOzeR7XFH8PJq7p8vni8xmHbh8UXq56hDaA9ixWL0k85MNtNomlWUVGaLHqiyzZ
n1+yVrdINMvR7zES9s7VSF5cF9Bn7t8ZmOxengFDO3qmQdkgL0fa8RZJzRzocbQc
cZMNAAMLqgrY/p78qu3ig4aujIzgqtjNXXblUpjxJ3SZYCjLaRIRgqJPN5E1vWtE
OpKxWXaBBwJBsWRhqokvzGhgUmXiqSqZFRAJG01te0YX7x/UXo/R+p0IWyB7OMR8
kyA/jXVPfClaxFZDwwXNroB3jBBjRB8dU6jMGzdADEng28/VHENAm/wM+bJPMtL1
5AcAng1Cse3vVA+6aARQNg9COiODcnXNnt/8ScZbxCExBTgzQQpD+t7ODdRNLAJi
rkDCQLOHCG9hT/zgrxXQApJqt64X82nFOcG6WTg5AV+p7ofAvlcmaEJOQtJZv60J
vbyXRx5eZy8PPyTZFWuLFABiokfJbbDCl0zsbAW9GDB5FBb+Q/Oy0pNHTee++3i1
qx31g8rVNU7bTpI3QiKC86HcA3DfrA+2OLwhISs9RQEIRg70MmElPiz6swJUBxZW
3kK0+AlTu9d6C3ojOg7gYQSGAenxi/gIvHDHnbfneZlBj7OeOxa98YsOVNvBnb5C
DCN5WC9YSDs+AZP7Ia3uJIo3VC2lGEuBjj0UCU5VoPJghr+b27cPWrt+ilXP3KPm
GYVrbXM08zl5n4Sx/IAqUxenif8bbRut8Wlu4fispfoNvbmG1uariEtPI1NsMhv9
lMnVzZrkQ4nLRoY//1izxGx/5jZG2ZlbYMdX38ghdzztG9saQDq/vUhVDjGl1dsf
szaHTMDui0fGnDxiUTOoKSWFlJY/AewX9YgGgsEyDdS2PF43sgc/L/cMGGdgEkox
gerFay8F4n55jo+hSsrWU+qIR4wTBzuX3LuLo67MgjtXt+JVet28QJ5Y9QPq3aXb
VNGHxnMXQvUe07pAEHyWPr1e0HUZy2XSJt8WVC9V5oIO8dtyPzzfx6e55x7hwt/c
cWSIjBqEVrW7wZnt9GOk6KQJ/F6DhtkHRQ8m+VzIqbdU+kV8XVBmOjNynXyO3+Qr
zC4Uv3tFrh5EPkZLUzLrxm7IxbXMfGgeo9W3alKYYOrs2BOiq8uND4Xwaluo+9Ts
cRdSY3f/IoMxNlDsHd57W+qkUqpSXdNA0COParG16BD1ZRFfRLHd13Zvc8kry/xy
maRHUO6u8MeePAJ+dUzOcPSepFctu1a1JAGf5+1aFN9ocCigs7x5m4NTAXy6Xi62
4S1SRn5HAhl7j7dnUeAFKzgMjfJyqS3cV3ogFDaraQh8vIxE9R+XgbZiz+rYLt6y
4AiUa6fMv1PgcWXzqkK/pIJo9+WRkTqNpg1J+DFC9hwnUpdu8t1t2MO0pSsCne4D
UN+7Poge6w1OPvZZwppDOYpy9tLImZ1Zujw93axP1XlMWwfscR4DeyYPGEJ4dOT6
vEMxjf9LSm2OIRgf2IddMGPjc4HV3oQvAZkiHPJBGpyheqoQSxzGDy5h4W/WmZPL
BunXC5H4xIvAuEg031hkldLM6FkXr++DvZFnRaducCZNSSnHO8nu26Klu3xawp7i
d19ZFkXWvBp81+RzVpGP0fgKyyQGUVdydpCod2jvVmx+fPfz8Rhs26XCAOU/EJmI
rFyxdcaT5SDxM5hQttm+7XCpvNTE3qGwSciMZtpuq2chXYjnQNiBOxhk4m8Xnlf6
8WOaiZ4j5wacniGo/iPBe/8xfypVvImdeG0Slc1cBOvbvPQrDef3UznAJ21e4ioS
N0kpIMVX/S5gTPh0O3IubX5Z7JnTNXcdkkJxpsz7rgZmtpnjFYjdFRwTwGupoWOc
GQfmUPMYZkjA1WmtTdk9hGMWoYfU08l/oHX3LY3E+CQR1WNfpOBDRXXCmAbSzKGn
vu+GXrteFlB28KaQiC45DIp8U8pG2Ffxu6OgQ/K8r4GnEegEfjgLyVeMsGZdiXRt
FDo33q3UQx4QYRrR7Q4SGsQvDJPyUhP1GhCtTR/ynypljJIfBvWTLZSdcQX0zlXV
hrxMAv2K876vUxhbIGHlQOBtNJMpWR+hC+VnbplWPJf6Y7+If4p3ocEmdUK1tKzG
z21Ma2zfxSTc1XrhE+yG/3uVDpQ213poROmpnrrSZPhHgos1fkwMKQu4eIX0B+bL
MkDMlpKiZD1x1ljZBfMK0+u2MOuyT+c+CKUUTXaQYSDbXQUtXFmnvxQoDCTpByEH
IHvZoxHndE8SG7LInVX3kj66RURAp4VIwJrpUhESoT332q8zNmxcJTc+S50dMeiY
oNpbd94OvsCKabvNjcMTr8RzcmfCM8vTfi1EeGgq5RTOx8HTaqwPA3aWxyfWQ5Cw
AtagxZHDXK5OLL0WY0s02iNeoiRvOtf44QV2vNDtsBG1+z95Cu2n6yKY+6J5zMCY
j88ZMekFa+OaqD2rpSEJGhmj9DXNsyEuTZedzM4sWzNVcAyydYU8h9ebR6uT8W38
p0lDlpZlyTjtGAm5LeVgPw+I/gZIuYUVdVBxwIErwtsXjPuh4JspElaM0uJZsc9C
JXIgvdcC73t8Nxts1qYOmptvMh4IBQJ0Xj5Q7P/12qN2rRsiuzvRK5DbuqFuvhhd
nFey8I9XbSRpD39ayWgbCpYkCCC/IwHdd7zJOf2Pz0Fa6AsaG2XwU2aOVtPjlJgF
oz1kliVgoramYxiLBkI9C5nIigC8BTLXfba1CDLG3jw0K7DM7xomfpO4tq0h+s+b
/IHLBxq/sanil6WwkKKidaSgWWhQCjMk18t6hr0AtjRYckTwWdxjR9R+2H1Lm0r6
/HKP4coGn8Ey9qHaQkziEXJ49keT/7uoLYk7l7YRL89/0ACaMQmua3tLmdUywIIe
H/80Q82qZw1LXbiVYJUFiA5cvIRC6XeyrQYpMj/DyoGr25aa87NfFYLVZo+X3RtF
wdrFgxqcwUwzUoZmR7SHuUWJtjJRzCxjTiFfbgEAqH7VOcGDZ2xWILthfaA9VCCE
QZrV43DSjxEa2Zd4VMg0lAPQupi4Nap11YZ/1nlh/SHwm2p6VXkY5IopUlw2VnO7
7Hby2HCbNTJ9qpdG2XFEUMrL5VJGRz1NaX1y1IiglDjg37RV0iWDscoGkOyNkv3w
X40b8mzzQmKEeO6YCpTToIkSQBHvGdJCVerk1htnBYthnmp1Q6IQDCEh3hwXHkg4
ocSiNL1lm1YDVNyahMxefiULMmSY3DjM+puims6npRuNA0g/oG/4ZSlI4BNHPIDv
Enh2Llrj7bhFRG0judZh1QEJPZAyPsbFN4ntMLFmLv4oyr0z0rlB1IC0ldGguZqA
BKEsrx7rDnA72Nx9CNjwBi1HLzYIOrqG7HzxJawGAAPCQpH2B+WJI8s8XMw6jBEn
lI75R7tlmmqP2WlVMJegHOPm9In6+jt+Bqcyeun9Xb1xJBeDOWklqD7sHZEN0JgJ
jtEwsFHrtwkGCjMlF89+SyKV6KISr5mS8Et72kSEZ4g4xscY7J65qcdoZCce/jzy
Kr+xU9BMLdcQVRIMdo7brBPsw2Ff66bPUvvQhjVTASyEPGyaXmac1zbqdF3ZwP37
YYOW4KXVCHpOtvYAHjSiUkt8scPO5Y06ISQuca0ZLD4AfRTpx8oz9vkWD8wqGoEE
T3ez/nktePp9Rq1F1rLNAlbOWTh3R1oDGdlbvlAgx7mnCRiYGcrqsh7KTpsHI4dq
h/3YOYFKttIAOEl8Z/seWkiIjQRMKx35ISBMRQqIfZM/NsHi5ALwa0nBx2Mh8qw3
prNaOJZ00LS1AuFhk1DJgWpCIlOAwIajsvOxUvOTS2inNEoow9SnvwvMK2f16ogd
7y5HHXnNvfeflW5pz9MS4cApucdPlTOxQc1Kn49yy4H3nBrbyJsQ9opaJo9CGeAS
vqZwQbcQFxCzm5SwLP3fmDOnGPw9bWBK5PCa8e37Cnyxa/MEsiEXzQNF7JlSW4Yi
Po1CxGUasTBylPeX+94NXgVV+Im0NLRtWPEvnmRo5E4e/o8iFVc5iFjQ+czRhJsn
JTnNMiZ361dMPi6tfJer9nsg3vxDl4aUL7YI7PQS1ql9fyRoNqosG91IOFbU9Zwe
Rl4mljsMVlqvqrll43cAXLtuFMnCJCLkHzLCDgnwmo6QOT8upKWaCS1fZUzkqJx6
FrN6MxLdUXro5usc63OxP1u+pJUQh9J3T51czgUk1GQWCFJDhJGNCaQwvKg4PxAf
597oGfB14lPv01s3SW4sQUxTi41/pWYKS2LeblK9oAT4d7uoLWrhP52yzG0rRdR8
xQhxA04nyzbo3Q6hICC9BcRWHVTHeibHStfbW7pklq0i6ZutyCrPT5aTMQU20QeO
2tM30uU3Q5RQw7Das/N5BfrOXeySf5MI9P2x/onPtmcgf0Z2fX+QsMHE5yf2lPJr
LXQ3dpX6qQu/xRPjxMeOAlXmnLJGBcoJk3ee+PczMDY4ozZv9i8kh1IE2SObWXkf
a8DwQpcj/5fBaGGEv0QUDAfAevo1F210cs+J2OeWhjDyaJYoQmcNmFMsNe/QCSzl
KadKzIqDoTOXPGZX462eMK0+4YWdakCTEtuYeOIIFXy5zwOgJ6QfQkLW/toNpdCG
jjAlxTTx9ssV/aaJNZ1VYpP7v5TT/6x9kGVtX0owIayXrNn8Tt6kTMH4O8+fx/9+
QsLhOkqfDabtzSv4s98Ud6AOSs5JOckUYXkO0Q0zh7jyid7YUy/6otXDPKHE0pQj
DT0x0+CbObpKMYCFy78f9OnFObtK4OMCqns838CqbaaVSJFZccy9Lb3C7M01rDfG
u2mXiImAUU2HQs7pu8T9z5qNtCX6XrrVB6aDDMe0I9AxSkhXR8F4wf9iCsCRr2WY
UHITtOUkQ1xov/cXRm8i/NQ24im3VHUg4A02k7YPB9hSHjlpkpBGCW2s2BYi+W35
L4FWqaEj4d2Vl5zD7HFT/Punpav045s6/1ANRtBVHJuVU3U3k6GPxVldaiMeSd0v
+9XMbMu+mNRYaRiw1bgNUtk36gDL42RvA+C3kTOMOFyfDZSVaOjQCO5rBGyp7iEo
z2EaN5dnbfEYW0t9yjQVwS9fQUT2f8XagKqI2VKX8oZVI4b5hGG5EDippRSGJ2Lz
1QOksCBDZ+Fzze5qJcvb/FaOm+cmfVF+ZdFEsRxC20ZjUVgjXO+tzfcFXO/ykxHe
ETJAJ4RU1spC+a4gZvJBqMBhLwyPNQWwx7vDHAdR6F8QeqnFuNfgk85KEqhMXe0+
XbgFdtVVbV/SUSfL/tt042B8TJXbLvGjgevgcwEEvGuAYRI21HavGWhArS/jOQjP
J8+clXfL2nnmugFZth2xB7yWXoHCxmzLwa6jflmb8snrB6CWKIBHJv5WZiLJN44R
VlfUqet05nzfJixml+R5tWDa2Sjxj8HxqgiGyPZLrX38nIwDgKA6DWs0fTPpLJf3
VXSMF/h+UjxAK4QeYLiaufheENO1Mhvv5PVsiObsn1EXKS0Mom8aJ1NtIQlxitHU
Wgr+bNpAoFT1/MY6o77D1N0cn0gqBEtq4poh0Dzhem8DEpPcasZ798Floy9Z02mZ
vGhPS7V+smCLq4qPT/knXMhlhu3m9R6fxe5pI9A5FyyeFRaKkGysy8XOMK0dlZXE
dcTNhDQAFv0D1v5YnlTcEUJxNcObub0Om4F2vWOmk6abHJRLwtnXbPrID/CtCVUy
EPY6v+SiY+LuTq4wm3JZDacTo0sjoOb0X3Dro+RsBGlKjTEjCo2Rf9mLURdOSwbt
t7jo4Q0FSQgLdSrm5+4QpsTuKrmhV/JsNl9r8RQrasJYqnSr1bGbgyMv0HAeDQJJ
bgoq+XE8Yeif+Ivp2dSKh8jvYv8rlWgARQ4Lj8S72Lucl3uzeF+PMsetrDN2fDLy
o+JmrgzU91ubIUobGObKytw7135WN+6if2NF5fPgpdtL9cS4bzIqGEZwQSmvEYlG
nrU8ob2zc6wcIYEAziYG2YqcsevEJwJ/mlBVOyLYaPfR+X/R4rhEiwkXfEGFznHF
troYO7rd8tXNDDlHkFQ2PTdc2cW3PmvVRnP5Qj6SgHERzlwHi3AGQJxUpHJk79eT
qOi7WybFzprksBh9SYKHvIK3xokq1yUYioWfVeRfGgZDHFmub0GgCXhzwneg6pDT
R4TmhZCLZ8R4hKCwK273lS9//cclYEmC6hPV2naLTtcHAzUEfGkkWzBKMV/VdYMb
BAkFXxykbXxMImd47DEpO7pgARe5Yl5FVLaMh7WMVfCsSH+UdncRaqOfkMvqxkoW
qmL948/vcbduOr4lc2ghEpFKFSjw2QOjfOUm2Rv6Y6kye65VX8j9Jr2jpCPdHVmg
0R8RMqew1KjG/35Gd+Edb80s0gn2WeW+zzfKaNYwrsXFjRrA1qGgeAGCOI/QKJ2j
iluPPlK0cvjmPD0wpfqIYkciADT4L315DD8F1YSYa1yR3Hx2kgB04m00eJSvsp/a
cEPhMKTN7o922GaMbvTEjZAcDZqhCBFRCDKYJFdgVvhQHC0EC/BE9ndvOzsNb50N
uW2/eMwfOYOiXM3S8RK1rxMJtnkpalsFBBlVW/y6voAfSxoNq1fMBy2QoKzxidaq
ZPq39DQIkqDaQ0FnlDaakHblcABBBOXdgzRzZkCIYqD3y+OmzBMOOeuuqpO2ohpB
OaRa8GjjbDqA6LYT+ly3cDXtN70EaXLq1iXH8rJcfwrodob2XXgjDztxEICSIRAV
eHUwqg3TVXznIDJTxBt84LhPzClg7ymWsSNzBujnxBF1oVu9X3C+BeWYxMip8cXk
qvcCuommEne/3NrZEkVeJPs9zsHFqrr3OcmZC9inJk2n38STzbQ9aVThgBjkH9hu
H2rZFxyNY/3+Uyq+46UKHKPWMcqKffFgNkRvVo8GTI3po0pZtkniBa5ikx17KjNk
i2lvLOlaqKNXQ0oxWnUlUJeqmUs/P+aQ6cTL9fZ2lyY3OrtGFvCdLAlhMTdK63L9
HDX9uCZ16y2JMMGnsNRppwQ3gMuB3e7WwXGxc2kdfBCIOc3lhD5VXkjvSv1Kmwzn
z7/NO/1SM2s49oY28VE3j63xIO2SOB9X93JS4diW+4YcjDaF7WvjYG0yJOsru7+x
ynsAM2SoPF7jdt4QLk8CDX/ApHDQQSUyXwJ09k1btvICCRrNWo108EczLoR6w5Xt
A0EvN3FXD3lbOySj3e6aEQApbUuBPAj5L+J32z2f/5sdhDzA7uPo14Rgppp2BA4g
0xVAV7CQsXyWCzEAWK6ftg5Hw+g68dULEl8uEt8GJg6ByBpqZXLUi1wM7jypwLbG
Z6c1dt38KN1FD+B5ONGfllfSq/gctLUNr3jvLQ8+aW8/aGxu7RjYs9cXN9eRhRt2
tULIkmYw1dfuIaqq7RRGjFuDQUwbwRyplsxtr6Q+N43V/CJdxUI6627NlCvAtyAK
vGbl2B51GKDaB8ci+BNd1APKy9JCjjf5ugSW9oyxvz1p88FewUIQp65FT/WTFLM5
plTK7FBI76T9GO7C6UX5u2anFya14KBoFUrwZKWUeysQvu5d1IM+t+OA70QOKqiH
b+pflLhbleaz1gPO1pL8EGOLUhz4TwhMDo3iyKpSqLKyn2PYD5m+iZpZM4vugSOc
3Kd9nvLvKil58O1iwJ0n9KCoIA9s/RlQSt177dnjcGD82yLvpjutUVYCuJoF6gJe
fYiMwlpOFsV9i7K0ZF5LyXOaFKlAl9L5xAPwKwbvxbYjJiKkTU+JiRzE0IgmtEGA
o6apjvtXCf8GkfxUQUifAp+Uw/A/CtgTGv9mrh1QZeWCvSAISvKzMlyh7eZBnZTh
BySsJaSSNH2e64/cOI27zj0TV7dcZGtTnTyanJpkza5g0Ak/DCI3g48Jd4K0B3RF
/G5Yb6TuS7FLgJovZua9zzmRoCkIMWWNUQVnopiFbuzi+47/dgzJlL4lIRwTxJEL
tfnVtZqYymnjo70QDzo1SZI/s7Rj7jNABZcvGLY7kh7cDLqvgX9kFwfLeZ+5eXms
eSDLTgqJqlf/fRiivYoN/eiJ9p3ziU2OQ+dpP6j3ci8DHnupoILyJaci8MoM36ZA
DbIdxaYGN7nd0oLPTyhNz38Vz4b2OBNSuARiYnIl3O4Stz4I3k2xJFeyL5vLouBD
l2dyjGCJCsO2/JEltdb7VqY+Yrgen5ppdUP0/4nsuBBUtN41s5wfLPJFV1nlVhMR
lzhoXQA0F0ZpxiWlqj3NKC8y3Iubq+Iievzi6JY7AaJOCzzJ3shmag2IA3PhFy7D
v1XAd+dyxQzgCZSWptt+LW0yR4fCkZ2HArTbpzJ4+rF0FxWNMtMkXEyvkHWQADak
epFeU47A991d3mYmszyovhwT8Nvu90Z3uUbbRfC6Q1rfSLykSpgUBJqHNpUOSWBs
6zZYL/TnHWYMHGNiBkweud2OmmCA8u9yxu93G+7pkrmdF+OdLEKDnIx3UH+ZunPz
pJRATaMkyXZ1o+5xp31PGKsWCMVG1KNkqj4K1kp36ToKY0E3v0NFKBvxWS8N8Nxr
jJMdMiH+AKTeNc62EidyqrDToig18+evHwIjHeY4h8626mtYV/q4nqPk1VarJk9F
A5oUsf2Q87Iem/Tm/5Chk/o3PZ+rtYFu6AXbyNSZRtCodJV6bb7xsNXHKYgT8gMK
u4hGELEMgqiHHYHz+eGn2vHgCYIhBkys04NzkaqWB839oinFTFqQsAJ9W4Tck+A2
3iLqyGqnL9aCgJ+i7kwBpuRd8/u2TVfmU3NJGQzBxzqUUtRZ0/qdBDo08hhtAO/q
mpmNEAHSxxd8t8pbvQVWH77m/iloQDF2tV6/K2vqj9S05mV2fiwz8b6wvJ7kKgHZ
CPCOuKKWFSbeh/YjbUOISk0uGoOnObuAoY5/1C9NViix2pawUHgFu2xtlK46Zeju
YiUqrXNQ+eeAOgfXBXpz2vposMhIEBddjCzG/dJGr1v5BvKzYqbnhdQaoZmUiluo
I9dGpu7OJ9TTd7I2/pKrJXGQ1claubbzS/FQRIAwy6DlTLYCDCm8spUJUwb5uArI
dTR28QocV2ivmfZJ8JwC+TjM2Jh81G0T1J3TLzEhcl566fyVRIhWqAJGezHRgb3i
q5xTDayxODwlZe8n2ikyUVkWfEdCpq+urTmUtcyYq8ySwL8/lfbXVttdT/TZwB8D
ojJXmtUeu33U2mC54NdkgbLspdm/WLv15VWP/VM3UuO3RWufn5OK7I2NxbRUbJPi
X+Z6pIIEjWFiFMej6p7qwsq7cZMTD3XHN8zo7TcYoMd79oy+j0gvfE4j1J9IMPVR
A60PaYizj2qo/adMvYtaOHdzoiRjEeLIjyNDl2X7Zkjyqwlia6ZZ5JSj8OYC+fWR
/4csACdXWJITe9GMXzAvbZOW2HX7iXFGBB5EOEzqr7o/omXDUpbv1cdCPOPF2esY
ZuCB+NlOIzwO6lgRINKttWt2gB7uOOITGOIpspk1+Y0Y4OHey5BXPdk0YTIOBsuF
c/mTONwNRwSkeaXhWCqzfV1eKfM+BGFjAe60oZmOIju4zR5/sFw+9j+bC16b9tIU
+W3/EHNgaOqf1Ko74ICqj1qkBNjAUxMemWlPwUqzRqX4ugy8nywGQ26ZkSGuAQfc
VRWvvaiuZG7qGpWOI7XfMvxNoVQQ7nmqtH29ORfi7VORc2RulI+hx8Hbiq1R+3pY
MrsJCdELFtxURMqshJbg4CQTWXJcRVf+jk1yieXJYboQHaRjy+/QlCdK1s4jl0A4
X7ReVEpfCzysKF+062HRTACw+Lz2TwMmQDKPqhGFN5Oz4jG4ThRyd1JLJoJp73Ny
cH0/ZWTk3pvsXOf9FRLAApcMSr2pMBktxvOxPgeyiLhbeYlfz7FmQ/OJSwC65i1N
BM6lQSzGqq4uvt2Qha4YT18/81zTQsklAMVQEcPv0tAWKjRd5UOng+6J41rR7juy
gZmzMMwhfW/zmEF5XlrCldEc5bdd1nDZ1xMeN/zDLYv3+vtkwmd/CtZBgKnzDBUL
qbQuaUnrENl0q6q7GqXLKknCa2SoCUGak2b1mT+5Peh2oFPtycViVf1OcqBLD/Vp
uwfFZ4a0yHQT3zQxaD3CBSL5E8iyOY+q9aZuhSErGV5tViMe6Czs6O0X4zhX6z1v
ko2eGlqlFO506/EK7hg1JwxeEWwGFl643jQRRwS9mAewG83lqhpk7fgnK8adVU96
85TJ3oEO9LLY6P6LPOXHrjoxgNlMN6ffmKkoWec/TJFugCNLt5LWgLz+SFzTMbdz
kMrMbH/a0Uu7n7DV85BSZMUn8BhialapzCm1gPFOyjubGgUvykQqygaH5uq0AJPS
n1kKNVnvnWMaPPOdZQNEkPZsHY/RerN1s8lHK/zeqasa174QeXVxu2IsWimF3g7h
/QbHFUrCqYWkEiEuTh+Z2is1rgHAGdc9JZ7a55Ui+w9uOkNJNRChqxLth/JhN5j8
GV7MNacTMIq0hbxlvTQen0A1hz7UQvMKcCOP6QB2MdYmrFL3TZNn9dxWTimmsa9D
Q+KuKbLCRTZEWn8lAZrRIU1CX7+K5OmNa+ST9phMsGBXQkkNlxLJ2xC58gX/aoyw
UUr+0n10cDEx8PyaV1Pto+fsj7S2SPCd1//rDlsc5laRPU/4BXTTAnu7ZTtoY99C
E3hVV6zEfRr35DqpzTjMTqxGb1+O6p5sX0wC7mAFAzeoTRPOF+Dr8eDGnshQNOzp
o6W5HU+eNqsYAgqRrGCbv55QSzT77/SCqeBaihE07Q5bPdSldR3lpcEil4AEXdDc
ttQPvUbi2VijzoAQr8YheldgJ7ev+yAIil/bzSP9prSLWpbKchvZ8k+4IlGvgwxk
GcO0xWdRhxr0y2LHepzWNzUz229puSXdXRsO7oVlj/7Fw48ML3xPH2LOk0xqfIx5
U1/Qr7mhs+5Z/rhsk/LY9364KwgE0DtglD4obp2ZVj6uo5PNOOoT2AeveJ58MIeb
2wkdZahKLwYKs9lzAFRXfiJaDp6fCkjED6nleJTCai9d5O536ueUkWdG5mDTmzKg
EI7VnswsU4hBsN8Qn/s2FN4ToHMhVeEkq7nD+sG5UvyEZnBSZCdSahxEosEU/Msp
qiCwZ+IhNX6k0x/LJ07mV+3A2JJmFOMd44ZGJNIaXEqKj1DRRiJUcIlvWMov/NAa
qxN34JWS/fUndNUpIaFVI14ZKScTyWVdHzSywd0tjh8CdkxDnJVY6/ANZ2ePZBrC
ibf0wdTu/iALP04xkUZ19GSuQf0fqJIkLno+7i6KARoqljYQQGzU7ltYdMkDa4x/
LhrQ0qFTfDF6rI26en69JdldvKdMcL8XdfelepTEQSHvJiNgYOIViF66wZnK/DU0
NM8A2Y6tLwhcJYlkjRXPRBR9L7p21F4XtVaPFQ0DrHXuobSUD7u1MzsYtcQy3vZa
JUn1eMLin31y98Ymant9XaGArnm5VfRu1WbemqhHBNRp2tc3fwVSNbOe95q8jUdc
2zRednvjKvUQmFxYiIhMzHMwv7Z/qtv59gSVsvVuFqY02ZFCSS5DSbtMu+wHsu8/
AyqX3uTc4sFDfhxwlc1FeaXCNPzHY1V+GW5zX3FB6b/4wYuJLlw6C5hwwgRfQ0dF
aV+IVbuO8X+LZuoYDofNGBKse+wb0w8TmNildQce5wI/5Lo2dBB8PZpmv+JS4Fea
jgXz0vNYns9sir16XsOFwi9VfiYF5LvzV69H3TVJuZiBXFNDREmS9JZjKNlHBj8q
P6CDAHyuJ3jrlgMeBdxvOOMOlLykxquq5IzXWv6N56HCSMd3dyz2Xr8xg5/veX6v
ynQ6+M0hLmJ9Dpgx8j0yAm/AfExfz6bJUko/QqRq7Na9TfbdNRLOh2U0ncuHoDb0
mzQz4fGc6J3tHItIyTqiqxSl68voPu0UMCQYfGwjuG3oYtYaXUm/LdRD/JHCj8n6
Nvospmz6TUERsiT6JB6f3aNNlOAuyATM1bSrqje8X2LVf4wRLBV3ESuaiT6nBlnd
lODVKReGOoLgSaIE50wIYT746+fs9Tq0XZH58dnaAENk6rS4OLyHcOPhhOs0tiOK
T2kIPCoLqYS9p9g1jWEQT2rr7uSdE2+9eTcvBlxAOEASx49FRfpuClqmG30fRkXk
C+k2Vp3gaSrfk9xNTVTc8rNFDo281XED45KiripiPl79k1G2LDJjtt+VE0/53Xna
kLY6DpNB4Yqo1mer7WuovyJCieHGHbirok5LVjr+qAwoDmfsJRTcrg4Tu11Jm8uu
TeFIc9ZSa5GSG9ESnPyNSM2Un6LtMsXzYaBWv1IK7fzWd8Ui5I9/B0kcYqFsl5yn
Ue/UatWYZVpp29PKcikMfWOS0mh+m5an+pYeLEjMA4ERN1aWn5022jPeA/7nzAL1
dlIprTB3QUdabo4WX4PxYcRpesxfjt27nE5WTvfHGq7H9C3DJjTEsMUcSQ4ux3T1
Bs/dskOph4KW2SWvQVvdBw8qzs/cBWjahkvxNTBHJfAWdaM2V7DR5d1MePejXYyA
FCZaH8M2AipRbLmj98WyHYKhq0yx+8Sj6xzdVCaAGR0J+qI3GVEk2PtaysTvZFDP
m6k8L9ycb2aVJAMMCW7GtfB2u01z8Vu85wYi46dQhW8y/ZvI3jOMDg73jVfaiufU
JaTqkcxtrKRa94UiHryZ4ATHjr8nkCY2u41His7AjzLPmZiasGy8FHYhinst4f0q
wlKjynAqHqpVATSY70EaOGmjEUGevZmtYZMrxIygfpz5e0IhhzE/6mYdF/oEi24L
xrpqwhoCcltAY7qN3wPAOfqPb31QmoDD81R4LgePAu/nI7GwtqBmRuVTDn205Vwf
NVvtaf+DoyATUmEAmV/HUabM5NM1DZWwKp4CLLOepk2DFNM1KW1Ilq6pT2A7XMwO
VdvncaRXS4hMVs6a9MNdL7lwz+6O6sgbMJxr+7mMEnAHX9taFnuzm625lEqX/s9t
cPVj5Jmh2BRSv6xE8rY+QfIUJMDrFrc17Jl9UT0MX+T4L1s+qfpDqBzrYCvSwSoW
fLA/ukKJwde+MDDrMhcA03WI1CObkPZhemDFaiJeG1ilNYGf+V+BEK8XYSSPj/sL
+x2XffqmlW5z85Xn4R7A+hllr765ySoa5eW+nyhRZoqCalKfXvmVE4CBZapWDvYz
4gIdTZaWi0azs+fqM0EaHKrG1xQ2Sm7PZm6bS3WZdapgEA8074/6KS+zLCHGlcb1
hM57nwJ1b5uN1ZnMgsrQrZIA9jmhwO6WIQrqxtMAgg3i/k9tYEQY4Xw8hRb1QqTv
8sTDalBoIWoGd3ynmAFdfgebx2WAcO/YEuP2ytydTiyliE9BeKMGg1wR8+bdmqJb
uYkypkJJ+PyOU33tGfNfvAQ3cnCpCkuYWIwg/ZLRyDo4OSNzvhycchncDlhudWFv
fhLDHcyU8GvII3o6W3QGjaAWUqwDXe9lAbJONxvcWImkqVMAHZW89g8euPgjTFzS
QKCn031Bhwy4UOvRyhF8rfJXK5ecJLjOKkcBCIEDDetnLwuvGoMPw0OeDw401rmV
YkhqKMpcECxO0H+AcAu9EL9bpZXUoUm2rRKFaw52HB73XNCqH93VeiyS8ZybGThl
dMfjVVjb7qYrqaFsmNMsmxOu1FF2l/iS0wW2Rr+70zqTLvs6Szy+CiI4XiakG0dV
7tpVt9GY3W/bbJXIefFxaezeLMu/Z1KGz97vaPuFtxeiGAvoRJ5wxBuy7iXvKBeg
RBGo9TO0dua/tbf26u8PZo/1XNg8FrFg1cAQZAY45V4fabonzXiA0z/3yJ7Qx2iK
YSYxZ+Ac2gApf9Xm1lAFVnbm3BKG/MAsH3RoIxbqDHI/2sLXeW4QEkk5x6kbQvOT
kXRCxjwjKPlBYSNJUnd5O1XJPIug/n6+NV1b2VG05naH+vCYSYNa5409dfM4Huj+
CcJWkx9Ouj2JVY4J1nZdBDX3TU9e3uDcTVHKxwISygle2UGPHbW4mUcvYLiUr5I7
DVbNu8enFmfMIUilrdi26TlR1BJws3N6BpqzNDunU3knk6r7jMnQRWU3EyXbAmN3
Cwf3YAIZKhrLNM7WdxSJSdNG2clOPIdrwoCPtr8V8vaB5gTFe5UngDF8oFj5fVeZ
SLiblOpjGu+HA5BkxBLWmH0VdeXnGfPeEKUkt2wkJkZ7pdGu2eAm9qnxDpvztJFD
VQmsOT20M7uXUAM8I3Y/97G6+vNIIhEhmAzgMWkxOxEXsZ3JQ0X+QRcNr7Omc4gU
fjND2yskvIpLz5v9yDXgIFUzUizBQjYp8S1e5h0DqhQkZT3gHs3PlfabSP7eu0b+
8fInbqGPJaSS8TsgXnTXuuLnnQERwiJGY4TR7bYMvhbfTKQv06Spv3fNF8Qgs+Ze
1SmJsBQOS2xr1iNnwxanudr2D1+tbGKlP14OvnAfXx1pn/mT6izauHplknts/Ds9
VldEfUbfcINGHC2PVf/+vq0JJpGmnf7C3IW2RgT9vLhjR/CZd8rc4JwOiz1IzGID
arql3RpeP4pZ4Uwif3Yq3N5HYvRrbXN/3d9bkbv1IeWrXpHHvUJ9V1IU6ks3FqKv
E3ao+ManSmiT556yhqJ91vvYmFI4wm6EcGeZP/+sPCiekYZWsMD5RyZeO5x66YDP
5LReVa7B4ew13o3eGERk2VH84IWcj58k3s//67g4gGJ23rgm5xQlNhX79r/d+96f
CQaPmQ9un3fm8Dx3fARKQuaJ7Aiy3Z8PMKPkVKIScV4xIf6+inkQCzIHO5PykiDi
ZEP+dxiCHR1aLBN4W2PXrGXRWarz4lbUAXRm+4BBksfqqD5cPCa1QOO0BlieRtYB
Ya2FYNZpTD2kOqVsz5ELDyPdesUIHpjMxIs2adSTGdBFAnI9ROEK5TscHIRfgkJ2
70RYcYUnBOX6H04Kjc6a4lukpTyuSTtyssGibXC0oHhn1i1Bem5WppVhZWT1YRN5
3QlsE1pAz9U5OOvQMNUyVPHe9MQITYVg/XbRKbydV15yToWn8Q6G2XWXFdxk0VIm
7pkP9AfZI6oC6UaqJ82CAMx1ebN6A+eTT7k4eBeOrj8jtwGl4y4bhQ6atGJwK2FH
PNT179jmaWCEhRnPG2CCKhfGOEpNXHrTzGPTru7F08d3oUjMMuC1HHfFXoqlYUdm
Qtcl0i4nNTOw7ISIziZvg/Sswh7zQxW5L2CAL0UERswaEcsM+t5M2jtXlhIn+GzR
vHanQGeifKRWHXtk6RwzSYMpulL7E3xwJlHKXsib7rJmQ9MzxGq4fjC2xnU2y9s3
o1o8KoetZE/CgHwounNRycEWMbYidjJGarkjaAXMSI7PIZt7v7p50Prc2dySuRvg
ZaGn0TgSH1kdoWX3YXe9ZknI/Gjq57CwpXIbLzOyFzwyxIa60IZ7L0wZ1ymRunBr
8A0ELY5j41D8ajdiJDCoVLcrgG5nVBO1z70SufuYEmq+2AvDh6ddmn+dh0D4fU0g
/izp+ELujlYUe3OOsVy64xoZSjc+e11rWl5UwQ4SdSpvIWq3+/fxwydyuHW9fvoN
5N/OVAVRaKRwVnyumQJvID5gaK91EZRHm9HCwVF4t3GBPP5fvpVUyLpqzQCfg2Aq
ufMBZbGvPMT5dc6kAAcgZ+fy41lg87oJ2V2Dg5asoh+K+9Dbc4j8iRI5lfWtPZ5W
0x8G7/Xc8erot4YYwbPA5WCl39TWx+/M5RrGRd+VK8vbH1dH833mjWlb2qtmsSus
WJ7N7Pvj9EjyR44UWH21nYrnScUx5JYdyFzH1oQNscpCDlbgxjcukd2+4jMgQfBU
1ExF+qod6AWiyB8TJzrgMWMt5xoFduTByexoYGDRvfIBxHqHImaeFCA5FI/ujUEL
/dc1hEolv/5dhDmTDwwR7DR/SXe8mC2Ej/uuFevXjNTaTdUvEzQoF0MHWCiu2kmi
fzfIxf14+4aavOUGmWfsgCb4ZXz1rFrDEDbfCwmgUjMC6SfBKNwqxcri1I7KIk1R
oV7WiR6V2hV0+HV53Hvw3vWf5iBoxjLJ19YEDDVhiDTdMfZxZEBfArtVe6JEbJWs
qhXnf3poKq7NRuRtbZrtvTMauWgzZVnBJJM9EfJSXaEaIcsn0TQjZMc0rN5J8/x8
nXRbAEvG5Z6sddHENU4DoeIPp4lw/w+U0UlXNG5/zwtiqpvc9Q1mHRxjHrvKYN3y
wpOT0rDpX9iYTitxmnOL+BbxDKjAIVCZV6KWYuFsMp7wrP7lL3xzFDFoGBP59bXo
dRkykpd6PwHPEXMMxsE16Z383C6E6I6jhlhe5LNL1oSRWQLZUkUzxZP/HyBFvj7f
fmF449zjijAlMo3VWMmMLuU9Lu7yxwpoixXi7PODe5P8PdtfyBtQBBxa4Alx3P+A
+TmIT5/fhFvqTc6uod2ntCAIqGnMvi08QF7SUzSm2ZdxaF6bcOAqHKuPNEF1Ifkp
YdwDvzzUND5H1gE1Rco93Ft7t7gtSqxcJqJZQefsGUuUGQcXWYzkcLT53GPMg++Z
GClSy1dcjxCDvs/4isN9tv2dMOJrs18nQhruPhSl8vkVLcHwLEaB8RVclTbf7PQH
Rm+ItDAGkiNDLMTIs3hzweCGCms25XknogO6x1ePQjdoKQwshRoeun+ht8x59rvs
xEODXY8krKBgl0+iIAJLLfIAKAHwx5g/kooLydat3QLkZo5kXZoUdqszrLMUVFXA
1P60zTAfoeabOxnSYQVQIXR81cvIKFt8XwQ42JX6wjMZgSsEtJgpZaW4xE6lNgM6
4mO7wCwam2E5ntQrA7TrrslbcHq83VpLmGCp/BCpVjnNffBhcS/xbwYec3VGrgHK
KnyJyGrRwhdnxSFoUIA/BIFTK8B65gyqWEUZ/ytjk/kiBk37GKbvUgcbBnauKf5t
4cd3vXScjHj6c4nmz4htE6aA1CdKpZvKPgmZHd/uvPgB06hxTEAccLhWfXaBaZ/k
3vqqvTgMQSWk2nbYZuRCRd7cSRGe49jAiGIFOesBKxYBjtQf8ggca/rWUXV7gXU4
1DIiKoO96Y3OS9evaMDhhYK2tKLLPWUxNi/N9ZNRTgGVTPfGtuM+BTopkJT3m1JE
CuvoOMKdDUHbml9SlXbvTmqw2Zbd01+PdNRK8cQRYgOdHNAHh7uqvRhFkqYteVxy
GfLWgQBe5iwrmfEkGtDykYuYNI18pZRr1noSi3pj4jenjoCO3yMCH/uniWr6es9F
hZrMKeNCQQUpNzRsdo+UUwFP/wK+u3csmTIdkXmBY0Oyw94ncEr/nUunqVj4MhhU
haLTAgGS84iI/UiaNX9DgSOBe/4Pe95n82WLBInFjg6jz6vwJaOhwbsAMPgPxFdy
pdAA8ki9TWgC9sFlWsNw0R1z78ThqkIJUNM1vAv2TtTjfgaE98k3mVM5pZBygDbx
AKgtxZLUGdeIzDeYse8NCjWHXjQ2b4rxAHnzqwQnvUMK0vByGqCaAb0PIcK9kDR3
n38N+cs9e9/KSnJkYfkRdTiNq37+yNt1paQiTwjHC6jBUbx5wbE2DH0+lonijq3v
4cBKHZB2nkC9kp75/ZXx3LeNMu7B2uojy+oNC6RSxjc0YquYR4n6u7SlZ+UfLq/Q
MHe0LqXavO6xT4nkUtV42dd2IGAV3Vlrdt7Vt204BCsY0CsJcuB+VALRv9AXH7S2
S5tBL1raxHoFTKhhUb8YukGONSPz6t1poulNWV5lfypTeIGq6JHumHsPlPbyV13C
i3VaYiPRGz0jsxBCjVburYVdUYhL+KrrnPJrLewZCMStRH8sOyboz/lesWI/RSSQ
sPEiVkX8Oy8cj45y1GYNfJWTw6PjgG8ifh7YRmG6G+lGQxg9hWoEpcu1fh9MKwbx
q7ltU4JcUxJALJtvRQwmhrRvmkWcM0mehzguwO3xnQPXW40Sw8kA10xu6SqiTxax
6Zm2RrDCYzWIfcZYQ4e3RgtExrsXLc0mr/A9ZZsqkCVksP2YOjfhv/PTRgjA71qs
z9aT2PyFFzltH5Tjd1zzKjbAZZDbLb6amvfwASoS0Oe6ar1KWj2Q0DQSJPfx/FqI
vxJs0czAhfPBo+JuCFhNfbSBEdQHH+urYNvGBvHjXC/mTbApURJdo2ah1A0jAAJM
psDU7b/bQfi0IIipMXZkCe15v73kpR91sdxgoBG3c4xMDrdpMvVA5RJ0iWSPUnk3
8n4Sp0koRquOp5B7rBCXLoCGkTgOz4iyGqsuNySQanO3ePfVBujgOSiZQWo7RzAR
y13hIXAG+I88V+xHMDSrbOXpB2cr6U7JwTlz3tQsS73yf0fP9mfCGOV//SuQkyXL
H0FqDr0XNsReqrVIhK2ziDRnKXstl4pTvzon68/+y6tiIjLRoHtx5vVgKlJumeq3
bBK8fvDhzkmBY1VboN5skXllyKTrNw7QtqJyxLTvaRncwTF/zQprk583RnqRcZ+4
z65imVP7OL0bx9LflB2ArgIBIQL9hU+pgznAX/9GNBLALexpV0Kcav3by+LGYjJZ
P53+a1lMU06gqcTl3pQTzh4VkWNG/NtfW8v+Ra65q+3gRuu/tSYhWH1nav094HIZ
Y4ejscT7/I5piAta9qvT8PoJQlDNDjXgYj70zkiYmKttCf/RJ6A65k1DxSACqa7z
fhmrwC2o47ZttXaVVcTGjC4Z/dlBLpFel3B3hhBnnPF36r5sHaDPHVkS+kXQrrMt
NDWldUBxafmdUcvallG6Zb8z9eFMpe7XeoSpI/8gKVMagozhQOl2fjouAAe4enJu
AAVmadY7vwxDNAHRYZBIbJRLFfkeBupbOFlQjbhj4JBJT50JwOYFQG4st7OI2+9j
2w/gxYLvaNEjFpAE1QqjrNzNr5V2W1xGo+lhtlsbhI9UN6sSCOwCmUB9fOp8cmZS
j3sWsTAn/Ahg7EEw9QMZPyPyZzRrHS2ABMgX8eDI7B4uDLH6GNwkhdU2h8CDGrdP
kD3xTWMzVc2lsi6L085tvN/Cg+KPBXc2e/x9Rz1DwvFrFdsFZSJ7ToPpvQbJJ4ws
G43Ojvzn9xmnrO0Iv7QU0pMEJbGAVx8ThipBhOhukCZWKFL66WBNlB/kMn+gGnJr
dx3Y5SsUEVjvuYTX3iCCMZl15Zg+5ipQ5Lj/tHkopykQiEVfPPop1aXITi5Wm/lk
2lHB+NGmvaVxWDVsc60J1CKPKnkenRZ4Q7NBBXgLpZRb3FWaRI73kaoAgCz102Sl
MrCDqXKE/fQdKXKpQ1pbUkW1bjAhMbmk+DCD/6w8qLGVceENCOM6xzMZ+9Bt/20n
oy874ATyLgwx1fIfPnyRGN2UX3VenYRjsarWLL2dJ9tRgF4NzqUbYv/bZWZ0w32r
ZBThizMRC2XqrvB2PHR1K8epNSjxbaNz5Z0szmfaL/NN4O3+yNxBvDyTGqw0R7Z7
03Xa25KYiD4KNGzFuYypS/lR10NslkiOgTi7wwnkjSHrj05VAs/j2tS13aofnNcB
m47kflZtjYlsMQDuyyFkgSt94YDGVpwgKMWjERdSrnliqmgLFfPsj6b67Zg0KDKQ
tOuI1Y3zXBYM9Xrz/bD6tgpU+7Ny6IXy7GTprs8Pv4tcGwcFDaLhk1PWruR3sPDR
Mf7K+25NSjvdCsyw2BurB55+H8AlhwdPfXvMN3S0Pyzp8Wdl+rz+GCD9Nqp+Y4lz
aLrP2x0RdQAjlQTXJx1VytwAOsmuVn9UcZK/uWn9qkZHbn/e3k9B6y/EUkoMzv1r
PZTao89z+VfwIUFIGe6MQ00T2E63jfMDL39cflsmwwq5D/w1TzClciCN5OHic7zm
O8ztXYKRMEF6dASN3Co1cXsRsZ9rx1McYSKF35Zot0JuNjPZgerNcO0e5o84o9FB
IeBY2bXe18l6QaXgutfS5/zpBmBl3zyiuBrOAhfggUJx8gAHRpPnFthBu8TXLJLr
KHIDC+h4eX3FYQBz1iN5Yt88y5QN3XoIyzj+irnMrHgonxK+YkX+9pn+/L8L5tIg
sHQ6v51fskFPnyatjITWRKB/kt8Wf8jo5oJCDzmveQdppcOAwcSwGrtqQnevPoDH
98ZBj7sxIlgkuZ2Mi/HPJzpXUUFmuHwIso/Q+Jz1VIAY34euxyFZVC7LLkzjr4Yx
inHl3LmCvMIWFUr9xy/BgHlXUgwwbxMxZ5zJScY7j9giP87JXPkN7w1QQ/6aov52
NLPkBaULfMn8iWn8+NeagMYQMmmBoxTpRP1HoMV6qQ6qW5dnmYLn1w8KGmeFFMTL
NeAdSu3QnGtujbBEQYz+Uxp8Cq/D/YNMWjsmBwGa9y4tDZJKohefcUcJhodWtlSa
cwlmzyYa5yhlIKrXYD5AFQ1iI3opgDGYkOYFJwWwo7Kui6WJ82OK6naRriT5F29G
G26catX4jwKorWJMojvOLoOOiG+c9hibP10eXpKpsI1NLn6iCnMQZ2xVhsem+jr5
/KsVtfWGXEGfr8/01q0l5vJBJ1zqYWDA9wzazzBwHMGtRjG4873rkMuDuy/JyPr8
QbkMqgEBcGcBmfF1OMLQ32r55x4ujXb+BMFNyqiFjoJ3r1g3tMnO2Y2+tf2Dzava
H71BlFMxrAm/2U3tGQ9Tju+t581bsY5rNARbCmlfLEzEn5Rf/gTdGStPJs2ogwMb
oNqmmD8legfkTp2nmuyDhGnifRqkg75dbwL56POvh5KPA6R6g7qDGR8YtS/QX+25
oVjC0M20mD2SaV2d8uqiFLgq9ZoYZsEh1sezHYn6EfBgRjOdLcPw8llL1TN1PdfE
HrBpz40Tt6eKwdYjWVIUPu3fxupoJYTRfhqrnVXa37MYy7qVJxRx18zoWFSikyOq
5Cc+p6jqs9lFCfHr7kThTA1Fh8S35CDpPhekjhZjDRJjDsIAMfiB++2kksk1Udo2
PWeufchf27RwTs9UAUbAHug6Jii+FKuyDxxLKipmjqd/3u4COoQRC0y9nLqYFkN8
rs+lmE15E5TLH85q7xcvF+STHmG9pJuWS+JJDjjsu2a3qHegdDLLpJDtR2IcjJ/g
1GJxfJPlE7v8vSkaUYC8CD9Mv06DOuVoX5Dx40U9mGZ1hdh/xYaMOjHaw+aUWak9
MOjEo4G1uFBVPthzC0+BVYVhivRouaCP1NhCHB+efi8eg8tnkhyV8H+4Iiw5FRho
6X4lhc7cR905AiS1wp9EVTkMwsz65Kn94KGsfxg19ERmE9v+vRUG9wGLyYhksfXx
ql7ERFJDu980gJHf++r04kg9AikP2VTvXUSnssFvv0MsX5z0TPIplyIq9mXkEXPo
OBoe8k7PZRazJN99IniOr7yID/4+UgjisHxaksWKu+8jwxS3OHGv8n+SnwDL7rog
TGls+ezYhKu7YPpjCApBi3cj6AY9HQscJfEmFOwy8bPLRkivEezhjdm7x2O+1Flh
SB+32j3i49yk9sHMHTdUmF3ouHzqlFmU86JZMcx4EFwzYJc4fpWgR5JXpa0MPTXG
gPYTLRuq+cXb4KnBV12KJsMAgxc9DVnA+YYCGkluPe24ARLPiGamzjNbKEBbRjzC
TBbIBdXkbTSOMS1MTibcElH13ErSkWPmmoKEZkhBXjuBsMQt5LxlnetX6oDWNUIh
JwdXmBkxwRVObDcdADffLTMq150hMpQmzQ0HTHYfNh7vzJUCpcNA9sCrQ6NV+rvx
rwYFla5TFQOduigvsB9euuvhYbXHRGp95s7x7B/t8XL/d8GeJK1CLSiodAivmzXq
iHzmmMftXLWQ7QfIM5oOZb7uq7DAJMsT0+DjGEb8mm75yMi5ori0yy1bzkwxniUR
aKvxFJjkvbRsivFHciH+QSIGWBxD3X1jU90fyJEQMSU8sGzT2o7yK5E5BUb55jYI
COcGsWdl6rxgckcFJRHHdWIGNRBCNxHtJmHd8bvt17vt35+Rin3XfT6jMwc71z8P
qVffvZ9fSO8A2QcmTnjMTKpbUlaFuyvf4vDpx56xGIVsRXwgnHP4mqAwYS97tJWK
utd/NVzGeN7HyGhvofar1OHqP7asfhV2anpHt4E+nB/MnmQIUMVek68m7dAb4ppw
HxqwddZ9DiJMDk5U4BYzR0z+fisNEiLZblhHdutpq+sBUsOwU18+0m7QeNto50Gl
IZlb1hQHZeTbdkKOEJCbbkkEF+RbqXq8whb7uVqLBv7dsG/a+7X3ixSW4d9+xMpx
oikfsHgzT16FHUpi+R4foDVytRW1SFcG8zbOh8yDxbS6f2ZshljubUmHncXIrYtG
TseQNgRQMT9S7A1U6YJ3KV58lFceTkIAry2+ymhfNGAe81e6hyviyCwzDb+hBaro
BFYigiE8V92yipgE0E48Wr6efghhKfufrI2BiDyzjGm7dplonuljwBE6r335HfWJ
6EdqWpHA60fvS3d4UJYw7xssTHcw8z+ZiwdfBqNjprzozCYYVDtfGq9VZalymEan
JqpHuGCxYgDnIBIY/kl44uxISdJtkyRXAOk89pBTixHxKD+ElBU+M6ojU00NGA52
MEUPouupSbo03ZjzAPFyCzH6qJvxQr780S5YkTDmykKhF7DvoVMX/DSimZtockz/
ZAZk80mV1cpl3129WrDl5sFXJ5W1o6NNA3gJpXtpEGmWXyPRWDHuDEpyXiPdtcCH
1zKsCjWpTs6LbuqThBWkzgJmaNMWTrJSoophHqeHpdRUWagsyauNY1nTDXFlU3W3
zf91r9BkO5cXEeeIG6n5tt0tMW2UGHsVsE72NKu86i9RUJkiOmKW4BmoF7WdeucB
i/vBtxIFb3qmVEbAzyDAS/5jSkKIjOpxqqmZ3fZ2sj3SgmLJGOOrrlEGkanewIuU
VkdiBiLFuPvZJrImANozvz7DfTOfSKShfbqcJJqgdj5pXdq9boFOWxCYfTUAdJUJ
nmULXns0gYOUEhY/yrYmpYU66THN6hfY3ZE1p7nmQMGm4bmkmUeYl1dx9FFcqdb6
g7OR+Ia5rNqXyvLIZBbxcBZ50VfpA/9iCsddXeYaJo67XhM5csO5x7eIQTEHFUYg
BRdU7jjJ76upfb0DL9lPeA2nXJTJ5sLaIsSKb2vieJeGDXPUiS/IAeiUWuBvjZVn
NRzXnPpI4DHUWrg1Rv0NnJY+uPDwOYQ08yAzs9gkzrr7dRRpz61qFQ/d4zV28wjq
qzM2IGX1fxXLZosYhg1K6Wckh+SiGrszjX7dgBJ4nLtkndt6AeXZnjJRw+JB5ohm
+gPiGHxHfbkOLiXUOCRYJaZOMtX3QrdCIjmrR8tpzdzVEBC+bgFLKO22a96q1+i4
oh55KsZEG5uvVoo/BlTro5skMg3HO2g15nftfJBmp3wbzc4oml5JXup2y6JmyJfq
PsPPRuGRoTt2kF5IuZzfN4gC25rqSw7TYypPhvtLwY2DHNJxqizD95T3UQG5Kjfa
mFsA6v1ItZiCLVs/eF4GX+DHN3Bt4V7tqyLl9R9e/VsKuCfXv+EocF6Dys3ZJm5Q
3ERi0d2xgEZpxn6D4KgxV2sdKcArGD2IAZ7VgLESCzE4pvaaehWyBj7O9nYnq8bE
Npwa08+QvaElHLNoXrcjb872eXaZpSANUFUAeFmOFsBPtA8U4T++YWITp02yS9Uu
7Lf+EkFew0X8jWzYHleD9+Hxvtc6G5CnmyE2YDO7WoS4lgMx+diAURxYcQCTKb6E
+V9Gy1ZL/AE8PPLri/2Huvg8HFDNC0OcxMiWMyZmIdZKYw7X0Fw2hBeGWVgxg3J7
XreRaIbMyAUypH9o+FpnkpmzM3R3MpFC1HHkdblS0NAEUY6QWuRE/E4rjcnEmuFV
TPbifqjMHSr9WmDVQnHzTUlhRYs28GFB7L/tGsDG4Ise14xH90uZGKgq+XovMTXB
cAeaoPF/gHHjo8UcxKBnUEJrCNe4Ck0MwDmccZuHDI/Js+rlCTb3pobzSuxK11J0
xIPnY1Q6WFUg22wGieZh3eQwz2WlDJhaH9w7mVVlwwnTlnVOich635su7m7YLqP+
/zOr5Q78ZG1NLrest7LFFXdvncrwQ8xRr/GblyW84cm7kyK0RbKF8W7eaal9VbeD
NNZvlIiMchToAmGaUtCXEKiOfijs4SDuc7gM2BMj9gV7IwEuc1chVTTGKKot2eK2
LuF1qOS/6zk3DvXoogpPKneLimHySsGkn8Ono1Lm/Y6kgoLToKqAmPrcbaha0Wv1
zXGfjCLI2iChKxSiLyLCNBc/pipeybK+FVW11TNCJ7PIw7aK8PW3a9OKgNv3FBbs
nubLINGPrSgKx1f/cY2s+TN8CSmnfrxlHU3Tmpw4kST+y0Z+oDe0Wb1sIdtPYZnw
S8xBw4htexiuLbrqBpXijag6YsA9/on+IPYXRHEGeKcDAbXKCaALd1pi6vvQGaPY
gCG/lCK+pJ05itFPp/PJRLeyow648MdA4yyLZ6D/UO8F1rTqrhxa42rWFy4ySyBu
54SGyoeg2JyXyAyVC9vS9OGc5b/nEW7BOOuNz2WYveQ0ounRhGPsn9k33FowU5xk
FjUM5dsu/D+VqrZkFEBHsGvsOsj2BkYwqfdIUn9jRZ1qEIZoa1H0x8LqS0pJjGvn
0S+pUA5NHNY83JBza8V6cSVLBWUR1/+96i54fehsKjeRF8cwlGHfhllw1NlqkGQi
GSPR6w7fH2F5AkrrHGxvOd/XGzYgJ/q8cqOSEyk0aDBb2FmFriU8eb+ql/lp1uPr
qW++c0QsHE6mBTJAkvmdyodJKEzhnnb9LmzrgMtCBz0DcZ0U24VaCg1YcFltGMxL
SV/XXLk4P1ysayu+CV2M62Aibbpda5S/CYZ+qT2PvYcznNyfSKRoun0Qa1THDlt7
3/GSqNNzE1eXOaS+a7n18krttXSviAjPYWNu7V3GIfgzmZu8AVvSOveNtqDZ8rTo
67wKUYn9GBhUkhq+jotJSo7hun30OeWFuduY4mq5mvOmpb5diyqsT2YHTIQAF6GB
1H5RUZaJDidbqkm9Ycc4ueVTa/gA7S/tyxY8jozgnU9yS8CvycO7WqwsJ2GB78+a
LFBpqKiozvTBJqBkg45yRywaBmffp3YKP5UKkivyCRtwmnE7fpQSEpcXyEevMkzZ
vnn60g4lpEg00Oa1qZcG7EP6lXST2Dn+R/F7Z0UBeuNYC9Ywwmp49ah4qpP2Bv7O
37FrX6qSiDc6c0cVknT/oFZi79GSjBPFEA633Oy6LUrbyqhov4ueogICCVCR/tJi
I9ZFbKHmZ1E9c0wQqABSgXhn6K5LkVngCbqdUA07umYePSCc2fFuQnmXQrwqY7Pd
GQdYKSVUhfMqA6Oc0+xu4I+HUbBEyES2dWyaPMzC4PNNO8qWZfg/6cKjukoQ5Jxk
vpoXCFOX76Np8NWUP5cI93q7zCC6tKokmisLwgZHRtnQ1OHwLqY/WhpBctT+6NbU
etXnCpbwIfte5sEZCBhRGXb7rBGdOPgrqblIMvy/dsb9mCraQ/tid1wfQ91Wvlr+
DR3r76YuMaMEfvAOaiCy5DK/tCaZ2LrNl40mOpP3wIhU9yFXzTM4fQl9Uz5t6zIM
Hqp8N4rPzlq8cO6WFjZ3GrFeUCJJQpW9eW3jhUgBqAeygUx7fpUkuiy+zzir3jzF
koCxaPYUD79shMY7j5yIvgOMghVQ8AE3BOIOH/5OzBr1UGSqR+JfOoX6q0Aj3Ftg
ndcd74Rqbmx+doksLoZmIc4I01/Sp/fp9I0aS/tBLDZUy+nMXb3QErEHOWsf1TzB
3vgGryHsx9j0nuPwYbKmMC6DAA+Rb6YeG2/CGrJwMWLHXWqQ4d7y1MoWKSea5xex
PRvCxFiwHqdyZ0lUGkhmlW0/5wFV0oXid3kozyxuwQ7Morb3jLwvAY6zZfTkhNlw
iFKxFkKSUBugIw6LjTRe9RvY01+FbawSVc5bRnOrw2cT/MrAW8Rfgz5DHMAqfLSl
4ZDzQNKUZOECNpmOolf6Jh7PIr42jd/bd9tgpY1cIR6QOBpDMWGbABfwJndEeZFs
sKco493YXlheagd6qHi+wCzooA23Zwj4UERtD/wMtYEiIYeZNla962oivnWvIjXO
POyMnaqPfqY00681GMB6IQzjDECGhD67kPkCYqdnYDntxlG5F4CiglNS6f5QivLg
ixmib+wVb65LLpXGcdfV7visEk+azRtmUiNJ2vKe6n7WsTvPrnpLOcV9oqn29bSe
g8DNd8kxCMjvos+L8mA9hs2Zjg3pllqrCIQ88BEIBKAbm3RctBWZERNom0BgBYXf
ws75YS5l0uhb1FsBPwchV7s1QlyvhT083fRZ3Bn9Cm3wRzKzpbf9dGPgg7a748tY
MQCjUz9/D1k8ggpfflcsd1yQTOHCULPGVxgZPKT3oJQqYnUA9nXd4dV3+nRF8l5w
siCKwaFmf3njhxbqjTxYe51fnv3/yVxwP1lAvDvcWTG+GjKCoBKVRvbU2SMPndk3
JZfgbQLy1D5KGNgGso1P4HGkseNIhO6fI9+asu2yCy75/+WJynrDABZ/vkvdAlSA
epB9P0TUqztLnUTn8fN5xhr+6z9p7/KrxZnQE4vAkuBZhJJI2ZzXiWj3iA7hHqxX
YFcf2p8Gz/k7d2KoCSH1EQyIUvSQFXkNtSuSy9cMwa5Iy8wpqGWwXcxYRdct0SnX
t+kifZOLuY4hyEW5C9KNWkv+rV7Nnf2xr4GXVqsph0GZ5J3uagOrOJG+B/Jgebyf
elktfdZLCYZHIcS8UnBcGa/ORUi7KTvDOmrqGTEMJQLAM3OeWe9uWP0y8ca55HWd
4AtRIuHYRJj2zQGOY0Jg/Gr6Bx7vvUHPNU+RJc83xisTh0hpl0hOYXDGrRKlgMTR
1si0Me92lG6DD53oje++XRJL+8Rjix5QCDRiuFq/CSAIYxHci/SV2y/mNFlYsPUJ
cXkMmRBusTJPQuYOM+o5INtuMWCDfW0+DErw1HuNjo8tLgJUjlyiyS8XNGuvQ8dl
zTZ0jWnWh1hYNKo73QTb17J2Y8sE2DxBT5tjqZCL+oURp/+FMEMbndJwW8z/zoBf
gFFNjdIK8ssJGmS5qVcgtHXaOL7cfUvdMLMrkwPbD1HMMRSmZWt74OkUXJ7gYJY1
iHN2hr6vSNbFHPlne5tGfsoxRv9WX2LoKoDr+cFAr+vkUkWPaKulcWIuHeCHuChk
bSz8tlgJ4uANR1BtTSxFPY8SsKGCQuXAz6XJ1ccL7kVUNgKavj9MIACID6qjQjVI
YqSSkaDqqWYDp+EpQvstngpvrDvpCNuv9PzLtd/kGPhSqKtnWCLyH/L9/XKoVHPQ
YBlqGpJgSeaWgZeb/uMn85WySe5m9vLB4bL/NbwE9OPLiECpB8Ry6ezwvSdMMP6/
fg7EHN++UQy3ct7Enw7Se3l4FbJ5nIloa44gb48jDbORsrcbs8uZ+cPZbhhif6Cz
X1bPGnlqnQD59iqGu3lEpDKabTZXD8jarvcDjCC2TESqdKi7cCP0EbbCpBQZc3FP
rwh1a/s0lwvmy584mRKZZ4WvaJt2cOEAL3RkutWJW7NwI93mbFZUwxQtRPmkJdVW
E8UwpwoMdIahXX2OKajGS4edOAG0PKPSHhNLL47ORgqyFqOhWk5T+5ZzYKmBFhy2
IBDOnEUQ2TjZxTcIU0D3Zh+YkPCXps8hItgP45CZxZfVzW+3Q5e5uVhp+SKwtj82
bgidWYMa7zS2fCWFjgq2PUgBpYL2gasg5RFdC2H3Uq3XS50pPMhtj1jbSesaGBnF
wnA6N3GnIZCI/MN0va6ZLsY2ic8fNkNxTOrNV+tRTbtSPjIqDIsj1AQmGEXFOdkX
F7ry7f/hU1Wy2bKUE03z4obH7ggUK1wUTEorgRmOAQPvRPcYiXB5h3gmHgcfYiBX
Jul0R7yyJ1fdIrMYoLUFpzu4/1DZnYjRSEIVjn/JgxvwyDNy/cV46Mdk6iOFfdK7
cNwV3hJVqm+/66EVcEQpjT4p1j7QJJMKP0gjs6JvmVL4GpfI1vXHmVb5lrvHMPpa
jGRE/aClYh3s49hkXMv4nWvp0iejH3ruYJiDgnLBYlzlsM2MSCWS1TOb33KhYa4x
0uvABzrZphtIKtDDGcg+gRat94rX9CN7sPTCiTdqkEZcigsh5DyYoI+BiMVrzfyu
qD8lWVyIm0EaQTfH5rxytA4yJK0zbIGmMXeqTCHm1KWUNktkIb+Vg3kdAO+XKVni
L134ka8kGon7zsKCchA8kOr6gFA2tl3GpGppCMUlHwMhRXYuLQ1dLhQerEcbCteM
hSX2JOTnYvGuCJc/1frT7sfrZIWsFk0FmW+63u7hTay+Yl9a5LtYxZF0i55XTMT6
2TbNLWv2owQmvfPLKlx9/sQDirWfclRh59X1pViJ+nWWuyxb5RAI2f0fqPonngpM
XoPZTPHX9BCLCo6A8+xSHrCp3TeAm8J1+WG+q2pMyuwT9WzIv6DreFH21NCHVAKn
GKQ1rzVkFCVvaDf4wSXxMi3uadBXFfn3Q5WZlwfER3DQLDmcf97ioPSo1HZE0K0e
QhjbPpA4vCpPOOuDmbpv44Q1BL6GRvIqHwMCKRQTIMMDwvyudqGFivBiszNAcJfo
9KjLFstMqnMAHaS8JKs3XBroxZNh2zHsjTzYgW8C5Khjzr3VA8O+PG3qc0nOa4WU
EUUIlhClSGGsy+NHKePL6O8mkab+2XDOI5xjWyJxM/y+Tg1Iw4N5SuWTpY/C98ie
F8HAWD0dr4xU4sc+jTSRGRKoAwAf7fCASDz6xHqekg6L9maJx9aadC73VbUXhGWp
ikWQOzh833Xk0IeHqioebn8jtM+ZHDTMuI5dKk7uEw3RwB2fNnSCEobwh6sgDX5w
6fuTL+7DZymG4iNqowMzW/L7DzWf1O28YCn3s0xSHrNglpcL38wk7JXvB90TmAYf
OKlEbtOKIOu46KYd5tS0Ed00bX/jnz/OL41Pt1AfanLQ3bP+gsduHiyJCpwQdl0J
Ur6/pl+zyA6Q552GrRCKPdkMZZy8psYb7BpOaQP2/CzpIhqMKlQ5brSg15qTqp+f
fvr+wcfa2Zy1N5+M89f4Sv2BDD4pVDOArhWYXeSu/wjvlt8DRHk3IlBMLBu4tKsh
x5iEg6zdUNmbirdG2XTW/WS7/QZObZf9tvvnrnjw3PBz9DAEUEuIG8YZKC/8sTCp
LbBr2dYMYK6q8aBboxaaT5/vlIthwKwe6GzdsXaFEvk8pFNHbuwyBwW3845O3m2O
TwEOkrDq2iGvBUTxNxtfw7bl/yraX+k1jgrYCimR79j7zfcbq7n9isZ/O5RpEbV0
6vBSn/Dwmx1Uo+u+KeXIjO0PC1OERsDbbwCqWaiQr2GqonJ7Po8a6kJQwb7ky19V
bYbUoy6FWDbdtCDG7AdbwIOm43KMfgAvOymzhMLAQFxc6ZIzNPEeRnwCkTx/cvTq
tjRYlXM3mm+RQfw1GqptTZoccI1Iclc7TawRpxK4mL+771zy+ewNFwAidUWHQkIE
zQAxNVhvQ+J9bD53KJXE8FSt9A5GesgCqynnd52yZQITc9VY/+/lGDpoJp9RylJl
LZnTPcKXZmvX4LH8s62mV5eQB5nFBwLROtVCHe0WH3Hx78L3cvgQyioFJjoFK8P3
nfBbDrHK4PkbNQlC0ZKtcNY8WxWPni0/GrW7Nf4t8yYPumF43pEomRUF03U8QlpR
Uq/QjYjgukqnW1foTEE2f9qOyFyFd2ibc1fiB1fr1un+71VXrctkY2DpTRtzcZt7
TEnrK1PUo8HKxr9zbAMsnURofyE33O/hMfta2lRmtKihe2CeJcnXBVflTCvzvitT
nOS2W20g7K6y3rBRBfz5ONTSZH1LN/Wea86+qLS3HcSLDlylW+gD/dL5GTiSgCjP
aWc9ufaOTkCVyhDHnOG6lXaevfLqhuY9v5hk/XTe+avgwBdcTr6h9oiH6TY1ZXCw
suDabg43jTDbE7doKuEJSBVBWvNYyttEk4y7Oon2O7AgN+86+OlKcgdnbAJCemd/
1tz53t0ZVI+lcfOkCp5msCsO2ReLHW58bUyJlyVV51z6w1E+b6bm7rY9OueDdPV7
x89r37Sym/4/iKyu47rtJCh/PNqKMrictOf0wGnqaUdzdeOk1yMtJmRYIBrR5CYf
+1c6dU6lzdm7pTIvZF93C9dzWk5p/3WEwhBtpWRTGNrBD5YBWMZosDlf3Zy2UIJa
4yEXwZGskguUqeXN0mbO1wPwIYq3qDJKqGIMPtRFI5rZP8R+q4l8rOBmO2UenrdL
kTJFJfup7DeRKDDdhCobtVtOjh28PSZpWNLJwvXZAauFrjzjhUB6QOBO4id9Ibrk
4x/2AM4BUlcUFEd2yEyVH9+Ly5YQ73dspHSGaVPWzWuRgcaHvl1rVEMuW3UTlIQx
y4BRHdl9MuhAcxLChxFVqX8rkSTtcUSgjF1tZrX7kW+rPCwORLnQztMe5aHQxIoB
3+aORGgIVcwgL0lDIQXYZAVHfUzOEex8nAKrHKgzUWImdmU7M7teWUXYYZdmwVRg
smmbzJmJ3Wm8QWui2jLwM0m+3qGoehIz2iSEUAwicEmnLO1M7d2Rk2GmzOANbIjo
NLpOVz8hK9z/JnMqrxlsIOOdSDyT0eOxsMLN/DAldOfwFOXNiP9+s3GzMwmOCj9y
NBEuNiyWB6rWV6QO60PDQFnC4j95MnwcvwiU1gkgkvdvBgT74NbrEoQWo0jcDios
BpwpEWPl05i3ngV2KoLBvbRoRy8ZSgYI5G4A1CtK2x+90AqrW5O3v7ZlCu36swUc
bKsP7fDSCAeyNkjIFZJ46AHA5csCbSvLZPOHgoPBCvNRndLZuvUofnca+9gnihCd
OcVLa54dSD5eZwzEgYbPPotS+LIg+POG2Vm7maE3tNMHGLFRVDvqt5kRRvQf6DER
4MKO81b/APd4SJHpbYYX1oxR72CMSVfeVC1qwDD5N+Nlw1Xx4QfTtakm5Kl191LX
QeEHWVDsNMAdvN6On6pf7lk66TphfjtGq3HkW5mSk45NrW30+hY5rRTuP89cFD+k
AXOSx3roQRYNo4K/FJmDS/n3FY1sGemBCZ1+FEkR7CzGyth/bnzO2QtLiv4/R6ZZ
fgcNvSXajPQjcAj/YCcD4hnrmq3xRNAJ2IyUR7PQHV6D4fPAaCytyuWNNANT88d2
0i6q4YqCbCkjKc8ZrETRt/g/MLogYVQxu2w/PSCjpes8IgUHzDmVgjuni1DSnI6C
pmOWpCx0JvosGrAV7/92cgKIT7Iy/5cuitF8kufdMQYMg9wSTUuXjdetRa3ekWbP
eIJ8y6v20LDw7osVyq+MrEmfRjzEAucnuTmqAUVRF4zurKu0gAtnpuyYt/+yH8Xl
JmI+UKQuBDd5noghMQrb9BmnlsXSpfZrXW5M44Z2C/ysI7Raha6ZRPDv16Ith3qr
5SRrgZnYvlcTYiygOtePkXthZ17ZD9TxvMeTaOcaXHRqiZh9xsCmDP6aqVIJ1YyH
HucaDoC8m3pM4vkYIn8atsxHryFuCUG5d2SktuXbchhcbJIUQMSZEToF2Xehr1M/
Bj+qSAiGwrllaReP3WrIOh23iSoWi+NEjIRoQqSnzaRcrte0UitPnOMvq2rNF/t0
waysFNwjVi6yCF+S7dkssP0GaYbdnJF+8DbSaz8MRHZvrIAWLQ6ISCOzzckiOZ2k
u+FAdO+W8OZc1+0oNDMZixr0Y+WQTERfbr3YCu+HL7HKjHClPT8JVtYsNY3UTYP8
wwF1DmbGc8eUmbOLbXlfn2mAtGwu0zl3CqBDFB8mcQV/olVqBfotWt9oLRbtBpCL
20hzdSeMjl+zzMdT23XQRR0kBOwhMBTWOXt66m3F6Ed6fyhz7Uda7pAn4NoH9SdJ
1qoSX00ZOlL0kXSiHOTuljQbu2Z01BjCPNe6JF50T56PMrSDlCR8Y6wTx+3TgaV0
D7jcuEyufn+cBh2lMpAGrdRv6sUIOMtS2d6T5G5hD7BSKhNIVmOH9Ig23vP8BwGq
LTI5kiWQMfqv3BWXad6muf8A+f3lqn6SlIvLBZN45mrTLhU0mqV4lulP2nY5XmKn
NEXjYKLO7fHOaP9LAfeqFx6Oi1HYC7wO4QxYouG45I6COeHqsLMoSX3IL5BApKHq
JSBWFS2Uaw+b7WMA3NDeQ/DwgqsnJU6sgmHg2tCx45nyOSASf7OBZe98a8aAC+n7
IT0seSwN2k3JxXo7ZFFJHk19uuKo4CqKdPKOlbVVxWG1v4tor5QKQU7u6BXvpGf4
yyDvi2hPUYI2IOZj0bXNMax+Y0ANgF86EUlRwVRDOkWA+/34GZXDfI8KL5i6O4HY
5lSZOhdrbbAMUiy/iW8sOYv7CRG4t9fAbM0zsxwRwnSUzE+YEMsrsugmpLys3Jid
LHFsgpxPLHn4LBq61DsdtbgYYregNep2iUFgueacm1qAj6ly32AyPNZLktz0YrOq
cklsi3Ro3eb5sj3l7rNgBl/lLCvG2xyQxrRNzlgbJuxUUMlGyCUcGEAGN4B9VmUe
tC12xN3scs+Zh7OyuqQTGVpgtLXiR/KzKaG06eZM3niXLb+M+39Y9aMUkzXamdSb
rDtQ4YAZnHUCVeOxuq/i1gr5q5M3FJtstIzeXQ9TpWwUlgp5luXmo9X/GazNkuXj
5EMivdQP5QIy8Fa2nsu1xj0ADdRvWYLzYGHLFCZoYOiKsxg7GeIiaGB4GUh0Uf03
hnH9rHekTIsa7pVHH1ToTsHmWvoLJ+UYAuzrPpzA/axus0X6iZ26TNPsU5fzCAvR
EohxjGwf926n69tShGrIEFAzdWN+tbKJy276d+9YA35E6F+brOliw8ZbwemgoYMw
kEz043hmAZbUEMRCcL3Jpg8UH4b0tE4zB+3pYkTc61cOuDN1m2VSpQFo9gC2aYq3
YQSW+4nfCQYw3Qp/B61/Ibi+bCRMTIUioL8Da70CP8KJl2K090wp8SuXpAUSwNH1
9MHcOVpTOsFT8RMqy2e8xOxxbB0cZ3xWRpjLkdhuxFmkdou94HQXQX1k/oz3bvNP
vrAGYMUjPBrEUArKalJfToLeST0q2QKj5mbpc9AhmJuGWBZsb2YaHu8sVA8QRrcy
VdxLsIwDPKPF6RgrpOUZiphGYvZ6kD6/XIhTZsWqfkt6c3XwJ7KdkR1EZvxb0jVo
Xm2KMr2WoAqIZO2x8vPVL7hHHa1u6TgQMc/t4Y5ANNuhsydeoS90gGK6+0j76pdS
9XqbxWqk93Fy1+V5ZXRrPU1YTmlQ1FBjCTSrqV8297E8cXvTV0KxZtrwR8QcX5nn
r7nzUdxGGvI3lwmxz8XDNivn9fjyGC8ILIY36N5F3Eaz6SBzkqEJeGdZOdhoEm21
aGtzTe5CY/nYI6ECsaJkoa4jXCpyD5EAZ6yRa3xAR3zBJSbJy0F02mmDJ/etvDTU
mizBaFQVxOtPuFjZ/14KfPOuGgo+1z1veVY8R/rUpRvuB3Mgnd957uKpyXwDKVmy
LDqlT44MAxnU0xzsjMkA5RkdgEUnVNROwSpbKeqFH7mVUiaBJezZmlZG1cf+65XP
Nb0L6UAmFZI3RUo4QvBIQCWaC5WZFvZ9zz4KMzu7CWl/HVLwbfaD86sPQEyPavby
n4EFLfZa+NXyO9wLZ7ZLZSPHtVb5MiBZIQ33QXzbOf4IuvkXe/ecg+uTrNK+FSsm
6e5OmAM+tjTQjj0BB2NG/8ebtylmyPOHyHJR1WOlEI/71R2RucEBcT1aIMwetyA9
cMObfgr/QvyVr/FiMHmNfuJmE089+9LhEz+unQIEOn/9nuyumFQj/D2/jQS/V3Bj
qiN2ho3TlYAF7sT0qdI3Sib3IodlSLvZcQuW+ZSQ6SQ2CcntE8Yvhh1bfjRmAMq0
BFAKEBjLiXvYS48yuHf5mFNBZyhTTGJIWQ1D/EJPkfeH8SRKxyDlVUc1cN1nIYoS
cRwwq5FPwWNm+fgWeSGpmwjmGnCnYXXJ5LUlX8SYexikYQmJG0noy3bGrXGkOoCq
4exTXgxnWiPqrIWImDwsFhqgzf00cEN78XxCxTeqo+D7eLn2pQn8AUJ8Vt9e8dIg
c2lnZsabAZyEf3qWZfvK12FJp0mkaZoN8ds+snNv7C8FstOh3REKbn/u/87yYgEj
LKNFVVcOqetvefDdkkwShJl5s+SrOm/J780nwO1eo6uBCZZQi/WIN5ndgSYVVFMT
c27GeoBNwdQct9uL2qq16c48OY+eLEj4Z6Lcn6xREQBknqnFL/Zcgpq7RdehCpuN
9Z7xHhYT7zG5wMDJe268JPCDT9PPrQDUpOvcUdfs8k+iICFl+7Q8XSHXr+uiPZZd
VIpbgwd8+24pGMHp2lnBzXLE5phDalLfz375uAidQ665+m5mpWl6P0/yCaJuVDg8
y6p94YYY49HU950kotZDWnSJPUwhrxVhWeOb4OtJ6T+sNxmbZPUM+L4ppeRYWXjk
mKCWH9X890OA/APYtXGxNkPmMdOpR7Oz/t2Y2w/Fq1UdQw6c+iqHVjbGCM6sqC8z
46d3gcXmU3kx8kYadv09962kM+6vEh6tlYKMDz2n9T0Q6jUJwexyD9u15nuALNrU
HPZxi41LMQmY1F6cI4ks2EG0X9gfU+ghmeiTA6eJk+GMSRNTHyD/ZOwFeNcWQLRJ
EE6zzuySBUWSiSZ6+wT369hk7yDdRzLuM35Y1ggPp94JsVvKxn1HGuNZOOZ9j9UT
8SP3/KTleTfnqPyc4xOg40OMAMsUGM4i/vCQjoxgoxcpSkiNWVILpqWOimTjhHyU
kiZ7HqXTE5csTqiM107Rd7YZyC81GjvDrsDz3tx6s7aH+AImxqD6ornblKepizX/
cAOgwhXpg5bdO4pVUz6NT9jrb9ZKnLyazWixJX26rWaO2BYcgMebSu6y6LV/cDE0
V2hjt9Px3nvdFecdF3LJp/9Sj0dy7E98lXajSU+9MbQM149ybBrdIaXP+DylRiNQ
CbjG8Gq0+GgXB1mEnUYRfVu370VzTVKjhHSy/Dq1CeXedf2gJzEb27bYhLkdgPts
KyMT48k+Q2Oae0SQCY5HWEjRNGXPAY1JGCBKnO73AkoJrhWh97644lq9DSCS4IP2
NrXOIabgu0dHcdUMDwaQzKr6LjCVFIu/yOqoH7WWdNXgRRZZycDmWhQsmMeboxTn
z4KgyW8S+x22MbEvbE0jsx5TrvJx6tsnG09xIJ7JejEChcvpVkx3mQGdmCRNNaOE
Q/GontZI44QTwj8McgDxCOmC0uaRARxthCBIwSbVWkJfxjXZaFT0Uy3J06Etpxmw
aHbq2jNaJnnvdYMHDu0Lw+6foPGS4AJi/IeXCb+HZK/JssDk5awALii+xcH0RCwM
b4mazrEXYFFvcLhB7IF9ATJ+rEMVXCKoTSg8YRP+tp+AWHlPWy2k5DHq5XGQfOk8
sZdbPMWRj2DFT5rGpjdcBpVvtJypdwHOfuWxyIZOdkC2C8/SZVHexFyiblqXhNdF
hU5aSUWOF1MiwmMX/26czVLquGGAjWIwino2PYZsKBA3LIXqEZbEF0vj2lXtnXtd
KNZQ9wWP0CTvUAnCHgb9IjD+BSFX2cm+3YTJ7B9roMFm/1BSgUWTh8XaBDFC4Wy7
NKhDMkRbWNkmrxz59I4KaWsx4bePs23SGCmptHoBvIfVNQfLFA/AP3fr+tNmVEix
qfdA03bd8y7OGgJ8+guzY02l3rxp6KHE/4p7ZAahD30mijf2NUUla5UwAyOp3dA0
vYHF4OdKfc2KtAbDqtkfkz8/h1k0nBMBPBjX9BhE6K7/xVt7A4QJsWf72SE9Vc24
9x46GvEk4KH7MkOObNYQ8cvGHReCXI0q07oI6qQKMiCri57ECO9W21WLFT9m+o38
YuqgrfmsI5Kb3T1HEa5J2prRar6T95VgwIOhOEZ/OZlx8Q/RRIJeSTJ5FwjUYXYT
TPg1ADciijtPGYG6utcHkw+cY4zlPFDiH8UU6QS/3zaVZ4Fq9uD6Ytz7Vmz9SsC6
Q5MZwWULKlDu6ZsPyNRPo6OhCBTiVvwVqF3mPLnthK2dSWJBtgAS1GxyM5AwopkO
OobtMAetuYPMelO7S+S3/bOc5AvSEjfEdnYK8rpqY7shcfrvzexQTJRKrmKLeQUL
xnwQh68ZuQKpxRSf6CHEMfDb1BppZwOXjKKn0jubUlT6xm7HSxoUtWZKCw31NyjV
vjXwMp0Xt8VXfkJZ6h9NG+lzka4pj0bdxkAxeSCdauEryKfwSH1D7meYPDSqaNow
Ea/MhKsFROQWeQ3WiLOv9G7Gh7T7WBDlQ4GL7QP2M/VBUaCik7HgJQHArb8QIKw+
inYEL2y0YisKC1RM0LJwoGAhQmbSHDVeYuasRy7YOWoSLD0IUuPPd2MPwfRaAqQU
jeKiAxrJPRZk3ukmBC8wL6vw0QLY5nwno12FnFr2GSwjXyGq2qRZXBrwgXZ0dDAv
u/LLzBZSCZW/sqEkzPr/xgi/Mm1GYEA0YHn0zaeh7GU7POTZqaHbceq2iI+5DQRV
L6qg3Sl0Iq3z4XQm0Huoeqt/ymCoifZ6Ia11XThTQ8Mpl5NeoEaw6xPf8cdyL4zZ
NS8sH3eCxoKv/9gfb6h37hC+54n+cBRc+92oHpmZ+U4AoR1A3KGcdDHP1VTZxl84
Adn/6dpIzsDylTtUzjdluXhSKYsMlLqXRAisArveH+ohAiGxxFYHKba1vac84Pxm
kM9FYpRxdQMhoKv4e+KwXOYwNrqbUZwl3gBlJ6aZnIcVbEx4+fKSWtSZlKSvFH+y
lE3Ko8o+GB15zxGlPwCcXJqXgnjW0/jXnK+FWnPI418+shCk+RcVbIoF4C/KKz5g
Vzp52wopfz6uXe0d9zsjwyldId4lH1k60u7YvzFa0ktltkeCvJ2O4I+TOF2HSTHF
nxziO3swjJy50lhcmd2sfrG8cgP1mSyT5plTkNihEYLMEptmt/lCNO7nMyJN2uuT
J3eO3d9xmnpJV9QMLThv+pEnoel6urO7L7QhhAdYEH3eteHeCdYe6h8th9nMgwKz
HfUjrQlLiiY15gwpLQHtQiBpFgzCUDCYkQEvJIXctctva3eTPftWilT5HFNma9Y5
KIErAO39g+tY2nyPdTitGaE/1+6fWdhOWvzceGtj5dWGX2Pf46KpSsOIKy2x6/7q
UaebMspyNpaplChnTiD1E3xhHjSY5lAygEZSdtgSn/oOq622gL3cIUc53aZq1PMR
1Pvv1T+FuL2DcvEAMcEFAjFlU7RoGpye5rhsjLSvkzP8DgbLoNDNpGGRn+D2j0GZ
VMDZ2xAZaleeEt4Hvuk6PQyFRqCoFw37LJgNjZuhbd/B948vY5KmAVSn3P8RhGvV
6TkvoTL3+Ltk2gwN0I64dbZ98sUFNCRNtx4ECMZaPxL7QFrRLJPZvs3yQazsAaaS
+FeFNNswkqCk1ID0P4OOXRdamd9GC8EZiBRuMvNJoGJpv+3Ho5EVD0RFXRHPcJ9I
F2RakkDlec23VBfd+BhxyIk7QPp0+LUwXcvN7b8nPUCqj3WeXzxO4Epj56cj026j
mGuqV2VtBcfxm3ancCtjju7nSUTjVpuNK9AmofSAX7VOZeQFiSNEdKjZpkcaWLco
7PsPl5ut0nyZ4W2GdblROutabobr0Ba6gmAH33BeOdHrFwZUFpiLQ/jH0J159L8S
9UymMJxRbfwaNafGwWt3TZjcESIsfUTAmAfnTm5N3NCs/KNBlJDUdUrDAymEEzUJ
JN0Nkrv01BJTZqvE1FVTKvDJfit54u69uWeTs4Py5vjDondXZgB8/IePwU8cdU/N
lsHqLar7z12btnJvwAeZRJj4hsSAZ3Xzx50GYqoKo2Bhwf8m96GswGo8K5MPttn0
f+JKJ0LSF3YBXbBToP6a/zGVW9YZHKkmlqhEh5ETJD+520bf7vsuhg0TwUjX+xTV
mRwmaNUU2R44Gm4mF9F4u4+Y0p+mMNaMXIg2Uk9ps8cJE0ON2TYG0qyt9Uc+JVvU
QJ43LRDl1Qrgso2qbVGLAEWAuI4GrPHebW5infcB0/RCru9vQIMmCUMPvdPDyCkT
TGxCkIIugAHOu5ledHqCWAS2ML4w4+5NkvoTvsUdHx7DslRVsPOruOHQVTi/2ZjY
Pc+MEF6oOnaFFzexwI8ogsiYAj0FUwJKjjQQZkEXaV0mPsYx3iFaM2UIeZAtuBPP
klmkCaNpgCVyjr+FF/l0ezbKgeKzXJ9ozABlp68lt1jF/bJXvr6+Xpb3vaHMIB3T
1j18q6A0ghBgSVZinZqOjSpHaVkxFTGbZmiBggSmTQM1tlis1BssjjJM/yklRcMj
CzojuueqpWFsWnnku/eU5rfGp1NtuQ5A1lm++R7VMghnuecwqP52sv10bNUqG3d2
yfkOTw8QLCIsVToiO4UM6VVTU62mv1dfldDQxBuqVjvS4KUhd5XzXnacNZeuy/T4
MOdL5MCQ98osQlhzfuQfeL/tK9K825MyJCpuV4R1eHxOGBsOrS/y0A3kRSRFTNKL
sgiHIr0kpZ5pYFP4VPjNMDs2orILK62rkmdT8JnNsdDdsFyAkkSFJXqWTUqWsyIg
FN3IMpi3SkOTdZygaIzk2oXe04mksjYuxRHHnzHXAlJnB3+oq8whb2k2278CAkTI
15QZHxlCK8SvJ2OBRWyr5QU0YFMQVgeqddFMNO7hJxKCvx/DCjR3haEMHuaIDmWs
8QnQM97/pwNoY5feHR6M6KsK8Msz6St4EpLgC6lyWpPmfi6/Mlmzt4wapFKmmPsf
de0BaygoAbmIdKc7VlOOsCnSthCKma01X2yUnBExguPUGInRyVDWSRKs10k71//l
a6/OvbMkdvtY2hTSqIl00GrTxlBG+D+B+MkVlJfaTUjXX0Oro2llJt1EQuXNTBkT
dqHe5LA3hzFI3DNf1GC4iF4vleLoaf2z5TfgDBrgbUbwdY7WiH67UVzT5nmca/Lv
8bikLC4m7rdHi0G27+FXNzhRzekOPM/MtNgMYfYC593rfaiNBXX6k4qjXCPhMwYX
IqC6vML2IoQOdbhtHaglyFhp+a2KMzuG/9deDaoFm4FtWylsJFIqUPTt521E59zi
A6CjXdjf9u6+S6X09qttOwfu7CxCZ4fdFNx7bQeBQCfnhZk9JF48wVXXEzgvNNjH
qo8ALiSbYrUf+5jHQyPwfwIaOYInyvrPcyIJS81V6uNp62N7YobdfCE+5TGGw/kJ
N+YeBnbPR2tMY+oMB0EK4knchcB1GqsA2o/n0umjWOihMZomcyiDztwAWcypOFxL
G2UKLKmrtyGbbkeW72cSOiZf10T6OMwQcUL8PGdhZPxovhishjrDn/r6GbBwNjrk
8By2Xu3DKUBr6zXqVLgEzyInO/JIRfqoy9buR+HSKAKF9FBGAmZBz3PoeDTerspS
EnhhszKoQbcvf8KIg7GA6KenuQlEEg87vffU6LS+jcqC8xfZ+0YLpX4D9F9qdmEB
vI3T7UnrvCGhanlPJtVYcbFk6gxzjlS58T0DcH26XVI3DX2eoBpU4eLS8NLqJLgG
a/j26zt1b7IZ+PsT3lhMiDscip7EVFLTMMn/fzEsN3AW2BBcr+6HbC+J8IAf5Ak3
+fmVJcR5Nr5vrY9Mq2VHD0Ckc4QTuUH41MoSgbcPYMULDWpq5SVvYJS4sItnOejL
t3kWmSqd/5dwerlgC25GDW8/mlcTcYK/U+BZbdT8ml7wOE5+EPJKAAC4sRWRjKon
k6bYcEBkVczPPGVYVapyUd/lQEU6hvnuQrV+bskz+Yda7fGMpQ+u7mC+rRQc4Drk
n1bHnR2t6CQsdcevl7+rrY2bUbaIWxHJuLQh7Eybj40ucVDpXx0AiST8IxYZeqgS
KBK6hNJNUFGpy9JQ3nbO8+T/53069jnyHF8ne+EIDU1bw704LnGeVsKWzV1Mp7g0
LHUrpB/cElYI4NXRY5kGh+ut5m21fNJsnUQUpuFGmyVZxQ4leDYpiBhdbi82wS91
xt1q1tm4qMb8QeL9uFU+cyUnr43EJVXW75fWQcX/ZLebnOvnqJqC0KC5hb5eB/It
qCcaM9/uFp5E9ANA31/qFXhWG/nHDHsXkABUwXg3KMhrG7gR3yRLL4BsrKSCvpbX
RAo+PeudQe5343uRcjCHM3v082NZUcuj1A7SuIvLaQeFaLgwoR+2clBJAc4kCWwW
dGDcrsbBE0tlaMxZG8e1I8N3GHNoY1rKW2ZWwp3MHaDq+Lmr4cRaegSZe7jBqoyP
LPqS51mCBPKSrNx9dUC4ZdUQEe1lp6t5MbdaL6ELqw6ULk9C8l0cEcmWXRsF4SGE
xuJ3ZlnSwdv5wCkZO+0nYjTPVFALO4yrpqK4VthIBjqdyhiATKwSkMfLghbj35zg
xGWw/vNaNW7KsTokc2TNsSItzPHNRBeT0Ax0EiPCljJjuhXKWOqGUyyKlZCiINym
RDDVq95iPjjuGsMxicm7jUoOp29tuRkyHbGWflrbsveEBJ1UfC8Xb1IxdRb4dWks
ZEpm2gQfxP1iYIIzhWVHb/wkcKEVkZMvXPt7K/UlmACh4bcrcZHRh7lxZemCYAXf
RA7Trhv/FgzZtxUm6kgNcB0Zv/4Yet/paFVRTVq32ejCS4/c7xIiq3Er2oioAfGM
FDqhOlyRbk83meAB0nqozMtRTM4PrcXpEbYuFAA/FODmA3Bm749yS3/ox4gUSnR5
iEZdu2l5/Ib0gcVVGK/ORVrMtuuoY/Ob4WsTlwX35yA/mu0z+BtHZ+tdA51h2+Mc
Yo75CGZRBfWps7+TQLwW0obWcxObDrKIcFdVvuzix2qaFde4mdfaXXlwFxsWBFYH
Ou417mS8We1KYipe+/LZ8zEAdlL1VLfrI1fO2KqLEjS9uSK/Lz534BLWA5/FA3qb
u9DJv5Grgm9UiqAE4HwffYPZnUY5vSEwjLvB+sRuWQ1/XMa03YDoEa+aoxypzFx3
gANBelMqRLJpYh0emogNJswRQVtxhPr3ZksMi7V1veRuyHIn9kpkD6ndrTql+0U6
A5cA4laspAiYr3GqxYCMPW9ltxT0vHctQKhQYTUzKiETMAkZbByk1ZUD97ErTrlM
x/nqCq+7rePpZzYErpvKwfgFtFw0BDZ2gD5EAQG9a4IU4RAfEMv8wbRt/O7XElbV
otNU3601TXKk9IwO6LGCyuG/37WFyxM0DKmdSsBzJZAkx7hptAtBX+MAZh9Uulux
PADFOr8kaOnpwMOAlQlsuMadPf5nahw2qUNwLysSnX/cxH9doMiQaoYVC+08FPnb
G8jyLHUlCjVeshZ/pR+eL54zEMf0wfBjZpqkLmrwzT3rpFPlC5wXlotHUelzi+Lj
y4LRu7LASoOj4cM2UrhOS1/e5iy2J43PF5CpKs+RvXMJU1BMKRpN5UK82PN99YTh
SpMH8AHCoujNcylkquHbkdmc1HRIof8X81h0Wx+0a7B0Rmw8agBNML8yG8cH8Zpy
Qj8cjCUa+o4+yw8B/aQTNl/HnmZRnAhVSoWYEYPDRTK2irgQlSxb8wqp5shB4cyq
Nau85IUwA+Yf4uh0QF8utNLQ47U0UfkN7o3zZ7w2kDLGJXhcGj/E2r1S53J/I3+3
AbmL42nonhFoGAX7ApWWgCVz6B1DnR8Iu8TwnkIFpmb6vR6BvHBCgClcE/s6fFUb
BszU2De13zSVetY50qFgYnuBxglSfqP0rMa29GGCKUFIbzZ9ZMx1VtNwu6nwsn6E
N5vDTz0byFaGaVSY17cum9MsjKXNkKT83gJXqE8yZLe59GcK09pkwo/B1CI1d2nd
K+d2Sjj43aCptfQdp57kltU/lKRryqs6iODeEAN6p8YwFgPCbQxDbjPQLTwTbOIe
QSPAjsx0hU+oDRzO2E1/aAdEY5/qmIolVo17X0CiKs+mOCSoQwXu17H89o9aKlyp
VMaPLCwDWOuZjDEg5g3PfjRywWWfvJSa5QlhlIR3i9uwVgg5KZZDIyinz20NWd9I
I64XawC8F6gQogKT12OImaSgNqHRYYWfIY4VLfhJ6A+YQPXr8JCuiQRbjRF+jino
1FjSwwx/bjeyxTkhlgxWa6uCOy96dK5I4WVD4VQNws7ZxVaNsRDsqRgMJnZuENGV
RDvT1keWMV4daA8SbLioC17bqnkBJQE7bqzxczO4cDQ6zXjPbEwqSicPVubrFnvx
i/lyuioYMRi8G7b4FkX7aytzoBFDip2mnKQoVaUxc+LSuyALgU/cxHVEoRfp3JvB
OOGsr7L6Xi+jAjTEo0x1CUJlMqjQpdv95o3FxlQFGvNYhnj23oJ92HspqKzKTCsI
baxHkfxzUbwW0u+5Wb8vZAvoNz3QByypJpI7RJLF1tmxVMNdt9Ba0zgyqVHkg2AH
8s8Unrp+pl6wGIdDil941xxEyYEoZjoRvsKhsiawiMSwbw5laTyuguF2v6+C+6F0
KedEw6YI6EsQVoP0SwpCn+NaJ63wphtuqofRF+X9XVVnxOqcSYUBD/qT0PC33HKs
euWJxPd4YVqohLmVYhYR7XVENhpCoxnpUVuW0oUwOJULxgu6skL0loGnMxBs6Dq6
RVoO4DUWc6YjuFZ9mxgrCLCZKGtLbjE0K41oxKEJ3ctioGbR8PxA40cmUF9YiABU
sNSkM1LkdvxkguwvHMKANBtiWfAqQURnoYHHos5lzxaRna9SnlptvoVUpOuzfIUS
SQvHaNSGFnOyFd6XUCKAEyxOFNqwIfKmuuipyYBXFDfehUYY7pSRYefwzunE5BV0
mB9GS8bBOXUVtbAr/zOK4YfKHLDARZw1+4+gqgobO2nzi+ux7+1Ijgi4/SbyyA7V
21Lhq5+WPF+ZZYDYS1a4qYg4HsZ0DaZovqstZr0kGrW37xAMyeiObkaPX50bTbzX
vYWQiSrN6gmacr9BnNPDqbmhgaKOE0rPtqYSvrk1xTPAeDPY4mQ6/9o/odYylmwp
FUM6ZSgXtox8ALIkEFsvnVPSa+ddNz0vFgZb0dRtRxj0GwrREkKCbrjiIba1+Hhu
MnELLaDVYNP3szg7Cmf4oqjwqxgM25v5wzycyi5ZujEgQ3sE9OalEOiU3TJDjSfn
6MCm7JOaqW4qjq64MM7u2KVjHIJxE1Ci4/kTAD1lUrC1WbyGkcs2BOFo7EYwnoh1
6I4uptMqZtXyWxEiCFPP4Z+tebPelZeImW3l5PwONaqzRNI5sAtFan/Bftt0MyRR
SsDOOeBqzGIRdGtIuXUZSapOhZgBFv0UH2QoJkRhT6NXu85Wv+z4OWFYn3h4zR9x
CHCuKJRi9UXz3iLHt3/FqFe2cgiyIfzNIpW5vJZ/+s6FEM3MLJ3X814/nYOPDpHe
tfHPG2lSvjvs4SnV4aC+Aw4Cx5Xw9uIl+7r3XF6fQcDBale5UDZac9WWKknzbRd3
G4gKA/gQgEg7C6zBzN9834gCbQkGLF0Z7qySDp67DkxxHSi2CARbOzEOAGO+kSsh
MGloFz7tjBZJFI/+qEiP36N/g99Bd7t0PgHAizBx0ZrHLItWsA9hhWPzL5cWv7/V
U5KLZkjI3dqpFhem+WwecURJXAxlAEcaBSgiNtxUUhji47aNdurUjzuCMqNSSHEu
6obcxaqTvhjvK41bPOM09N4hLFsX7j6lKcezAeb9G2crXQR1A5aJtN6pm+DvaUiy
8mymi1msn54Jq28mtWIy7zzajmF2NSM5NAJHE/oL+dHFAcQ9i1rg7Nxy5QbbIdPW
CguH45rQ8Bhim5I0xGy9ATOE2BXiJZ158Xj3jobyjjnAu9zoFDEe+VQYVftJeko3
SMFcfHNXDXqQ4FPZ0scNaSebblXKxA8xr8LLejDeu/3fmB1ARUZGDqSqc4SyN7DL
wuctLW5/vzQlWQgapRWASk3MACBJKi5NlLjjGzpoeAJjNlZvM4XJA2m0mZNtWvkQ
l4LOJ6MPo7MPuEr6uZp3FuoKUn1wmJyi2vJt0L05mV+V3K6pfWXtROJ8WA5z8sSp
CIeCNEdJqDV9ZH8AC9vb58pzETJI627Uyw845PSOMFSv7VgxqqiDFofFlIARGNgB
i+wKDy9HpVYo6fZwLCjZYKGwq76INg4LzGOCXZgFdssn7FUMIQJqExbuUeE7gSBf
8AljBC3yAh3c9VYxwCgZrZCaClPU+tOuZ8aUARs1NR8X06LEsNH+oaBQn05vhOSq
VE0SliYjsAA0m4+UGn2vYq19Nwv2ZKUwSdw+ueL7JQ0to/I/H8iK9M3FK/2ty0d6
CeccQTw2KUWMAOgYFrTydnA+7oXVMtnttL3KYppn854HZkLwRpTwosuxSEMJ4AhH
FbIhgyhliq+fYSu/kCeAu1hiq0edG5tMwGt4+e4c4TQbvJ8V6F6CffQyiG1Nqmen
G8cmcuRXT0umetQMZ2KGRYS6r7jIZE+TBwrXyn9+l9pNWRhHaxckVc+pOgc3EcM6
iHUzbF/S5Opek5zXh0LHXNDQWDVufgTrb7w3VNZEneqaJXtEViC36S1Ojnix4HYw
bJkS8ZY3Y5NxJ0X0XyGN4/SnyZJFzZev8szhqwJOUcHXe/8VQW/13nfBp4ctNbxp
yRxUxHSMEGYQP6/NXiWoVpmvslYlQsSnIAF0Ea2KFXTHqDeGqVfx34aMb8JESstZ
pPRXuL5f6U1SPPl3iNoz/yzk7SjW3TAfAtX8J4+0+l9GXlkFS5NDacqrbBPi9yir
+P2HZFzWJCO0LtYoPssLzTGJW2ITnLnc4FBT6xn2ssFQznRWgQrJ3EFZ7fKw9Wwl
hvOGz8irmQiMq5YPj1kL4leDL2rf4zusaRVc15XOxz84MR+IJh4zyMu6XHH+oPiS
13EN9YfSYz0aQ444s5VFAj/YhGmNDrPcc0U6/JbUH1+kRWhz9GKm3ji4B9cJQYQi
885xM7O1bdPIM3eTKuJYMhzr0/hMUHlgL7huT97HnkfqIn46kyfJvBtTBXgGGa+2
oHLl9eD0oGS+gYEeqL6ni5ITMPANGll8E94G8mn3LHqkbUZaRXIy+JWJsu3eCU27
r1YgiIz/SpOAu2dK3/R9mrjJAr16QQj55zmFVZ0KHBZFhe8IBDOo72BLsmKVkuox
88kwNp/e7E740xEGWkvblLPwefWoY47xt2Nm5kp8LDocNRrMdQqRjqTk+msMp7a4
vI4IIHt2LgJXGqHb2mBcO8w/sPLnhH0KDWiXBlJhr75H2yltdes31bqXFcs2dEVO
zcKdII4qnA9/6KpwO3FUUwmUoM4qGQeFNDAlaSRzATnW4PGzMrQZuTGfONQxx6gr
xDPGLwIz9blqHBnF4fiYD76Uf7v+gOom3YN9iE4+8K19ARG4gbud6nqeBxdiByv5
w3Q5t8AAlIiN6sCOFOHGvSwn346lOWCWdXVSEW+yiw8z5GQW+cr7wLqz9WsZhwZP
GHZaR1kDsVPY+b3JGz9F7QVia99ft8nIUI++OdQqWMixO2T7RgPDFMeziDfBzrtO
oVG5Q/TuPnAXNJwK4HcZtMd2RIt5Y6uagASj5dNmdEmwQEgWW7a6RHEVfLEV182k
3T+QgL+tA4EA5xy5XLvS65i30APtds3QE6zbG5ypqlQ5WcdhHSa7R32IJB4W+dfq
3xShRWCRH9YWJDPf+1eMPTDggz9OFARYoV5BIkQ1eQExsuaQE+XRW1h0U/Eo8sJo
OdbdalY5tDxY2wDVDhVa8XcCUoOU4/ClMUDj/hG17ybEKMuRE7IIVRebIFJivA8M
Ewt7fBGGv80QxGRYJvQnK7EcGzkwLyg0GteM1CQuPJmkciED4av1edE5XI49hGGK
zR0jadRb4sEjfDX/FjriqbUFnvF/Cv4qWTq/WkP04JB7oetKxDvJhFHfHFT6r2bZ
p7mKMeQKtJqAkI3/iR/AXNkEYF1c3Na+ZQ3Uj0qERMlVWGy8yRI5u5uiFJyvIatM
ruUb5FHeOXWS/qnsqkLiIQGYnzDitc8bVgy25xV3oUXXQ9Fkrhl9oIziF3ntbMwG
L7F+3336g93zSVA/kkUW2yure+EHEOlWkYxPHyim0GssuBnpcBdwfCNcSm4ypTQa
jS1stX0uWYJT0Mw04yJ7tlASTCBwwmo7x2EMR1JA+xWaepYJQOEgM7dK3q9OwvAB
oNTwnFej/pl8l9mCOktO4zhd7LJjEIpC9J7Itl9qAuhp4HYefcV3pAFMxmjOs6wg
gynN/nJuyg6a9MutcJdbasCPjvLYs9tLjsG3tn7G7Kr23916sgi2Rx1GE22y2xQO
GTMRYA4ccfwCaDgdDZ9mNXjWm3Mp99Kf4x4+8XxpvF1fz7JaZ5LRttY0P+c+y1XG
4+k+tK3Klu99Y0TK7tDpYDLzOFPY7mhOIkomDs6eeK6gH3FsFfi+QB0mo8zoDYr/
9l8Uu7CubFvhdxJdZo8rW4rkRqCLdZ3NoYPWI717kmy03dgfmfvrqDxOvFSkZ8cP
RTYFYRXlm0ghWG2oEIncwc5JVgNqeq1M++2LWpxlQtGoaX9WVHZQ8ne53PYOhrEG
3asJxzsRBgkU6IChbH5NRolH/c9NlfQhyDUvUobp1OMqCJ0PUgmeWF7w/Y5ieE9T
Ko52hwV2ce7p+eiBJVPf+wInoBT8scsv/uvJFKp2TJQ4wum1l6Ak+i27OYW4XIKq
BdR7jIgGiRbsUFz4Q9EpZs6BiBHRpNRrLl0cYWw4c4v++Bl+o1k6j9Th88+MuSsh
Pts9fiw67Faf5GMgWU5xWQdAyNK8jm6ezYL8PgQH30jCQUWPSgFxuYcPMEZRblxw
hnb1y6ktV/IdpiHVGlxq71N7L7t6mdOMxnT7L/03rGbM6KHIg/Q3jd+BOTDpLnVX
1EqTesBchI8ylc2ZbUEfjhYBlOo06zlUxl6UHoqSsbpW2Dh+PDuuI8Nce4HIzvTd
kCUD87N75yBWLl8S/jk21nbmLdrcyIvYASnsRxmvUHjr1xZe6q+vEjvGay76WAU5
4JtwPxA8feiwHCH3ikCqPleMZvmYZVhcKKTugY8/Lu2CR5jwt4EouqsHTVcfLIlR
xbvJCK1Xri3Laa7svsvMLh4NZscc+vRgEhkhN6PfqNXz26Amj+WmKrXDVvnlK0yz
9Isn6OfqcYDz3nYXzwFV4DO+XtqL1HyAsH89Sj1hEAE9sppMzWxjvajOUjjrB4Cs
3xC7TgFdK2IqIvUKBttR2EYUx2jBDYoUVvoXzPc1+B0mrDNeqEvlq9+NfHDAy0fl
v8uM3y3SKn/QlVH5AHLVPwpKzOUenk2K6fZh4S+F/R2Pg2VOx82+v2J8eFKXj3NU
dXJ87QEqxHqVdLtvTSMlv7i55hu3DaVA3getbQ3o71+dUPYvh442TOvdwLSnUOyA
eG+vDSQAZRLd3Z8CzBuW22qjpJMcWv+L1fG6U1EUxuAOm2+SSuBRpiZoZeYlO2mz
H81kk2bqOKJDW9nsuMqTZskzcO/aqaS6R7iyL658Kv6E6FaEpVDeiOZ04CovRkBU
VJOrWLx2AYkFZHRkLz0Bykr/SqmCjpqiPwmzGVj5Txpoy2VKlt7rr/4UN0ItCKhU
6p84EsN/ZYtgD3YII655lrLdvjIAaDv8FSHFaTB+GAMVbbw8sGHGdHYhIHUByuvt
IjR3FyoyMsr5qSVUUbU2CLnZ4uD/LTqk7NOdZmTyZQBA3kejF0QXEHh3e6mB0NyN
wG9dRYpeS2i2uUDEEJzcSunQIwCcPoA6UU1+jMtJVBENl9w4IEDBmr17LDvNDBBy
0uqCn2Lj5zlaQ8dww7lAPyFRfKeTKRFPlHbbxyQClX5/5CJENEmKXiqGhAqM0j//
LGj686Z5qNafzgiX/LNZ77zpkt/K48wuB6I+J7x7uqdtWQEmSci3LYfxBwce1S/e
j8qWA0u0JUe+V5qWMVJ1CBoy2/my1h5CfW+JnOj+oeHQMeZp9SGYpkE/P3ALyegM
YU1tbx1iY0TxQXhl2KRttfYuURkRdRMUvfEUh6BQFdK7DGcZLlUp8rKmvF7gFc9f
GwoDLGoMmoAorMld1lBID+YECjOntR6qs/pbR9V0FC2AhH3s3n25WyJLN8zzaxzV
0p+7JKyqdB3CKoHSToecD+M6FTutL3yY4NQe2iqHUFQBQ5AshkYcmQ8Qo56maWYz
jt0EYaMKdz2IkL7u2q0a0fR4zNGfgQR+/wcTAp7PJksZyyUdHCmmbhNWdxeVML4w
TMJFXh6x0aM2tPDqAeheoYsCGTr4D2p9XP58SSy/I2jkNj3GDxdbxbVYYUIFvfNG
Cng3bG+tUBz430lpKoNs15k/3CIK+WM335yacCPv33aNJzIdDvTTJbk7q/5EhLID
8qnyToODnmdakSJ6xsYBOAzYC8J10OPk3ZAxjLXZ70MBwLP2aS72g72qZI+lV6kR
mAoNvgCIL3ygwjdkYcNE2OQ7SvzBToNnmMU23tu+zPCUQIEqSiYs7FFeML1nOKP7
XcritvmNVY/IB8XTIqDTOnbYSeOIsMWggaapFheC5WaFbmlRXSZ1QbsfzaKvctun
IRtmsb8T2q2sfriLCS0GuXMo4CTZBSZSdXYmwu1pV5uYhjjWAqBxM7pFcdS+lcAm
/2DJxXj+KnnftRFtpi0a2nAHFoeYMNsEH9qEWtshRy/3dM7Qq+x1syyvuloJVdDU
cA1ZWqwS/dGYegEHn3vdrpqXZjCrV0qPfKv7hp7S5VZq2e5gMYmUan1JqMG+Oacw
SChvU7lJqUfS2W2tmn4rbxUx0i11JWRSuwawZbKxPpvIH9D8BhVGUD2ttUIv52xz
5jECkydydtxzP3A1b0CaUpkzlmCwhHUChB459xBo2loTO6Mr91ihisDhENTyLqvx
Gv+E1XoVnTFrPm3emcWaYcg6wcPcCeo79d0YX/BJPigQdHGcb11k8FcQNvcrBiDV
mgeRiIZZWt2qbhhHw2IE+fRZNjvpvUCQtlorQkiI6HJglril+pUIQj3eEysULRsm
koFmYAXGKvx/K8BW/u1P53EzzkMd0xZKdcN0kVEmN9jj1qy4zMUVC6Ltlt8w7Nff
sYXqO1WXZ6RSgjP8qKZ+Ops8K8WidWHFO4g0FbJjwNt99/SnRWCJ/GKosVOEyOQS
1Ili4DM8C3YNnLg12xJGONpb65VqMWXWIPiNFn9Yt7q7qY5yVP3+TsX2mYHE+USx
RI1g7oVAQ3FYdcLl+xn0+qwmE040CeIdRQeBLEqL5UCeM/gSz5/2EHseorappy+i
2k8kxbckfKfd9YYU8ISYMBVwVRHAluUwjKSMzPD+KRK/RMlgvNg975W0gI+wm/V7
327GK+l17jl5pIwZycw9k9RVVs83V6eeCzKf9WKytvl4AKx+qsptrmQlOdsFVZip
X8jIL5VpkzimPFa0P3eaofjQGuKNzGGUqsp6kV9or1ICNL8zs6YY6Y/V68F1x9ao
DXYwVhAbcXQ6MBTErnVjksRA3jDL9LWvOwngexfs3zSKeO1+aoBDqqtyYtfGC/jm
cy1kJ8hb5uG2jgImaYFmolL7QN2qynRRdh1MowRoI26+r1bz7oAnzism1KGJ/9cf
cquMbYWZLEErkNR3bjSBuiuQwgPsKC33oJZZQ8RSYpfJhx5Q9aZMPCtn7trpk+W2
hZyfsdtqTVUWxRTQE3uL9/8R+cFNfZqQ9XYHZeDalg+2P+8dqK1nxCQexJmd/6rO
Lk42zxH+NWXUrB0ET2A8KGgi8HhZSfcJBsi/fMl90MvM17d+v/G4ATx6SF/kEAP3
I6x1SEqRxIEqQXMOk3mLXcoyj+bQk/r4/XHDngduyTVdKlGg6kjKxXYnIQrismVz
eEeSkeVtZ3HeCQ9pADxQ8xXyGQJkIFSsqJyPvJvRp9al8DR4bIJ4gwgdmfMydIWo
a2eCP+agg5hGZB+BTKGMmOBlUBTQJM+HxyVnKg8tMPKauPeE9Sw2IovEoGEDfsDr
1W0YdhWqms0p/fxeBNhVHokiJjtTpjVR8IOzZ/0Pn/u/bTIm3LXsVE9l6OAZrI/M
lCi+njtowFfhgysN3pd9iO8h7lIueNkWv6XI/ES5gNXc+sLNML4yb+ilMet7bNXw
LmY4wZ+Fl+JOZD7MEULYikNN7SNcC74ClaYayAVplhhgBuYKxRS1pbkPSylrIqdM
RsVfvDWJ5yzWEibYIjUr32sW0cXz3argnixWsQKX/C3N1qhtWAe0ehcLcsQsVqMs
Bwl65rlhhvIl3pZ5VDjRnTM7DyAXGpxd/dt8o/vwrSYCefX2vOhf+vY5LYeyJ/Z5
x5uW4VO8PreaqWukQS5082J9eWE1oohsjiGfcAc2vljwcwF5IimPrrM+ryeaYfaK
5c+XyaBkzTddlM0GOt4DFqUcTFq5SuMyYb+Sf3VDOLvSARFs13sQsfQw7xBToZnY
b5V+Zmg5jBAXJccdysOJJk9d6qdtdzogsOignvooyba9kaMdrwtYGD/koHLZMKPI
gFr6lzFD7rWBcYcNX1Phq/nIdvr7cFq+qJ9xgJvwMQvo3DusDFjU/X1GeDDJFwzo
6l498++MqEszm0EAmKp06BL+xVObuLzbxok6dH2259xWXfPRpLtBpIIZQ6MzPn4m
GEjpUVcmGaFuoa7i4+KGTKolY9vEt8yRXjVcUTQ3ncCJ6OHm6Qkni4FCP3z21PZS
ta7kyaQRA1G4kl9g3/61kjuiDwFkRxB0QzHeZLyfEr//F1pjCZ8jiHg3iDjwuN/R
i5CTgs8D4p/ORZ5LKQkjzgJHq3naOmeQlN1YTyCOG5jwfrJkXyXUvcrOguS7qXsO
OfLa+F/jWn/5a1MIPF9ocOk7NimFnalKzFFrMjsdImyZDmpMfKbS4HQ36ecAkyLP
TH0Q8MLin2sI3EcVa3lOYr3g6ov2uzCIsAWLD+nxk2hYDy2SrNaYN9D5JpzW9nSo
7mjXXTvuB1Y9y2FkLaY2KBvRhZDe8uHcBVp1reFXSWMUSvTRtP2sRwDVFNo3WMaj
I9JT0GJeNIRPBlkY78usQSQg8ZKV9QlKl1PJKnEJv75o2iq25TAYUCTHTx3SrjUn
m/55QGdpU8l1I4vyy+TTAmxQn8ojthCKIJotGuZkCkLOGX1xzUjT5YImfsukOiwR
8u/UPmp4alOXponJD8n3AREg9FO6gLaNDGUhlp3PZqTD3LR8muAptKtmK9G4YonA
bOCEkk/Mvtc5aJc1ti2TblHvRWJUxotkLLu3wGb7CuMLyBSnUXD7lRObyjq7OpiV
p5/NOIvF75KTDW37lSUfu/O4tzu7uph/1Q6k0aQC7DBTpbeiEn4Lh4oSwftCUYf2
8xmU1iXDMg+M9wPxBdWPNgpF1YaBLBfqfHa0Cknwql9b6EEYd9p8qLiIp9R0jC4z
p9l3AE6rGW3mkqcWsb2eGVbA/Fuh4jVsHGhJRGVJNiC4uJxB+7ujeFbd1E/dtqdq
xhGXZ+HyNgpMITqlr5w+ILSUZXwGSfllXyVGylpSZLecv9+P4MDQf/2I5yYuHt3m
nn6vrqYiR+XtVPUw09NsARmIofW/WKfWi68PkoJgEK+9mDcOKvudaRornj8Ib6Wm
LE02IUt0xFgAgjgyPBI82RVrRnYdMxdeXdppoATFur3qnyMfno6QRPG8ZfZIclU2
Ys4YkozbRNGQ8qI8ll3c2rTPqy9iu7ISqAIm1+JS3nH4bovCj60TJKIO/R1KCtpE
0EBtjVOSIk2IqfGGAQ3Ah3+BxI99uYIv863EmnES6izdMpsVaWmjMG8VcF+jPidx
26fg1/kkdZIw4D1/wqt3Ppww4AyATXQTiYChfF6Q/shHFAAG7YkCp9bFLMrXEOGE
0IGPKISnxFgOW8Ou9yfw7Ka8P6x/VTZok722SEcJYaGJ6lQEGiDQY9fllJocT4cp
3x4dhQfUgd8ZJCP7V81kHknn+g+ztn7ZPO5313UWRbPoNkhNldz/kxfQtKZDU64X
mF616in5hXb3q+nb9+RAVbe5pCku9eC+omkKwMMD9NzsNZ+/ofaAzY/ti+gta4Jj
J5FPVZlA9AscEd8l2F4LMzT891yFdQwZrE9aFzQI2U9QSjg0B7JkoMWYDsAxvira
IzubMDOEMPD4VLfeYYJnhg29KZhDqYL0+Wli/M+Y/GQ1sfsW/66aFFsqJNgMe62G
+cTPjDDMiPm88CWqZYfMhehnYtJxnpoktSqWTjJC4rZQxIPTvK9CeP1DOCQd5PM2
UwNcEe8Sr4jmCcyVGRZjiREA4Ni51P5g3sZN+WyjcVv/FBQMrOoAIFQpLwvwicpa
rcQf53EYAMi1OI5tzjaGYtP1I3v3MektveKlhPThIAHTG7FI3QRRlaZzlg9HwaAO
zuX3A/3JAXQD6hQf+oNmufzCUoBgCrpd/59lKN4lyI+eLxox8SPoJfUdEf/OdOJh
Dmv/M4TRZkbFjTGOI11Ej2IrOAD0SGi7Rpxeq7RN7ReEVM8t+5Cnbn2RpuLsPKVi
vRE7XgEWiUY3wVVKFt94D1k66OrfiGmZQXnPuyWJ8D8pPnTfBrUG45HqpBwAvMtX
VpWE4OVaxr2WJ2Pc37pqj/T6T2VUkmW33hrt+a+zKRwsJllwrWz4js2UyGp9ORzi
jgrYR7J8zgT1ApYaRuKR2fhZo/T/nEAc2Eon7TRk56a9rVWQ1eUZP+RxXoXxPWO1
9FcSVqpaw0+ihLItWWlJL3jIG9NixXl4WeTSwaY+ce6c48MKiDLVZF/7J8m6oQ5Q
dkoHKwJQFSDcSLbfovDKLwGYWfMRlsJ/PSsNqk8ziBrtQmv0wWuli0ne5K5RCGAh
JTtDUZnDIZMY0GEDZ+T5n0+ij9sXBSBUhQ3QLdTXOKghYBcukE/2BZim0vGhq6KR
rprsoOdhy4RNXt933pQNEOZRG8L97WqZ4pttB/59s6CPfz9fej68J43R3cJM5UJl
i6YwATUDHbGYDEEJfOuMhIdwcZ1lN77fLQxeW+i2wBIytXJFAqYJC17IGzKQQ6zb
g7XBJ1WUjNTobdJNmIwlNDlKX8gm+IJCotZzFjzA50dq90q9ElNJhVOWw1v8yobE
0m3gLGLJTd9YRCW0jh+dlcbYL9FU8Nm4dzNY6J9LElyiQ5O87UGmvCuS0Ht28a64
U8TFU9jEPY5j/ks9Qrj0XIU5QCSrEbQmdROHrAR+r99N3asgae2OTgxDeZRT4FKc
BRs4r0xdaiN139MgCdwfrEbsLLabQtlxCUFtb79BG8165wwMmRsV4lA6ayVcM8HE
TJQ7J2OL+tKmIWnCKvYW+Pllh1AeFK4kyUmDzZ3cR0z9fvv5NQJ1lsh5AoqI2yan
Yv5Nc2MbQ/eHEzN8cwWueT3dcRctukutxj2bcg8N8wRFGbJVGpuZEzlgjRq2BojE
jGsihRpQnF56tp668HhZbQPgENxNMuwnspvfWeOxUwnx/iiQXIP3736w2VGqSpC9
mrCsz2DoIy81txa6XHUYk1AXPkiQDHyVTeyXICDXE+0g++lLuqGADF1ub1F4d3+u
2eHNHuAhIbftiG1eGdRp4W5qTWnY1as4HDZO4e+3FVJ2rB3FTfzNIFV7bHF3i/Y+
vHzaozOuD28+JmGouAMyNwTR0eNSoZIkgehWLTUY77FFvHic0CVm/iyl4RE9nWhU
eGgMZhInhk2xeIWHu6NRAuL27Y5iHWUnJi/0Rhkvc+KASQ4S532yjA2qJFt1ja3D
7oHza6vips96ZxvpHSUH1ZVo7h1Y5WfGWogj/zX1kCu4RyNoh5cHGWsgZzhhzcxN
krpRUQc31w3fXw81/ukrxl2gmXx/Q8YjdZhWG1COQV/u2uxEVjWnYgPgVRCd5KAP
vO9NT3iFSrFYOKQZg1FFQrzV8mmL3tSnT7UJdhXG2G/zbA2iy5IJTwccZEwxuQmD
Zm6p4rHiukwylK8M4IBFPv4mKuQao7d4KN17oZbJYPp5BMOnTkZxyw90tejiiZs6
yBIgMdTYtOW1hPdyfYK501Nc+UdRbKh5Ymveh5Zg24yByHIuZgSpLA8pG0rTrhxN
hg6Ik2jk31eD9gpqV7dMjyDsfQ+MlWzssWePonAvY3S0z6wMZZJERvnxvHw06qtX
U+ev4VfaxgsZHv5WDAeapVvGgQtRi37tFHB15J2TIQD8co4RMR896jW8ZGvOBl21
9TJDswv39O4mgvaUSlXusYD2RNvJjGMdpG625KKFStPE3vIr+apAcNegIBf00GJR
Ipp7iK73igROOG3rHqtPMM5wdQnpVIKYnY2O/MnoZ36zBBiuYM0PwucLcxOh0ixM
QOFzvjQNK8otz4zJU3joJX4iz1h+94qYkeFIAGGsQsDHeU5f1CZpkP3Sz9quC5HD
6lvlvYL+LepHf4iFVNykyhdp8v8vOitTKV5yTwmda7yR7E/05gDzQ56FdXagnqWl
k+dwsfJVfjyEYn2xEEuyWGa/xRXXUwGIQTe3OYXSEu+O0Tz1U3rO87rTkAdA59oW
xl449k5kV6a5Hxq4cMS2aXS5Ew64uOfUqZf/M+Ebkvw2MtS/6pH/uhPEpWE0BWUV
Le3LZdWrPn/BsBYyCHbNzaD0EgmELymWixhH61tpUYTTm4XGbJJCoLY1kekHIkCl
Vd7GMQbkToSjU7xVAmX5VBqEhZGYYyMpXV9ymMV0IsWJGjwr+vCVXxS4TjmdXqb0
PUEupdV4SCcci7M1oLTTcRNMVJT3VU2eZBlCkX/qd5nXJY+TdcTtf3Ce38KAmDOZ
Ht/OlE0Z+G7Gobf3l5p/+RzrbSW/hwOpLDVsHQiWmv4xHiGmYRQSa7iXFq9K65dD
yxhCGOFrA5J4FrODC2sat8NDNwZeYDFQgAFsTvxMT+mtsY38xSO3Xn+2nSi0pn7n
JBRNA0QLfRDKglu73HNpCaY/MZBpX21rLJsT8sVuqyap3BAEJsi/OuE/+/9gDrgx
UekqoHTpVJNyUIAo88TEI1M1tPgTo29X09NHmxVAAqMIaBnPJItjGESb8JvsX0MB
ROTpWmPK9BUeg7D8MehTstoiRQoKWsrXtE3lt8IegRFkw1fyOLmwtdNKs7Xo0JnY
N1My+nwWzNwgLY2YeOiiBDbD9wCqYyhvAYwNk7kBLvvwGjHOYtzcIzizq/t35zll
+Haz4RJCG8mHgbtc5Px5y+vVIIpEYcBbGGPsqpwsXhZjkhfTIbkC/wW5USZpvknh
rwmvOKZlWEYa0cYPU3snbowZd9m/hWZZOisDNo44yfHigZOjyKp+aMnFucoVcutm
CADIeFnuO16oVgUou6TrudIh56Yfk14IExfJjp/Y+Bb7ei6Jzi253xj5ivcVuuCQ
s4qtKPPOI7qP7o9xNMugR2RU8j3XmJp3ldWYbmWnNawIIRmuKE8Y3tD71MZaSH/a
RvsiqYz17vUNSwevE118ycdXEZnfVEjXVwHriAPHLwx2dnSziHYK0fk0gYKeXyNz
EQPLdK/+MoJLjtPBS3it42RwtdUlOd7PrWWJFTNuTLdoKosIDJZFb0iZOwa8h/q/
rSLctDd3CK54l1wpCtY1QD4UlcMKe7Eqo+HiY053EBiYL1lFnsL6i+esfmuVvwnp
ic50TLxnWnIQY+NATS/z+7Mds1H9bsnz80vEwRxwbAwtZAKlyNMd+4dJ5eYsuoQG
720CoXj0BiWF2rvS9ucs4KDtWZiQrFDPJEgoJUp2Z0KPL1kyDIhfDY80bbbfTpqT
d5lwUe1NGWblCBmALqmIuKzb0yqUZBQtnye7bfexH/bqTXjCpzQvQFQKR10QDraq
/LXOrqdoDpECjSqJThY3Ft+JLkXPHdaTESWZexKEpEYH+pNDcTWiG8uSjI8EafHk
5UtCDZAvi7njIYccIrxduuXBCKr+ah6yVtP33uDxD+1zA2rdLH7xEDsxT0ZJA7ZO
E2QipRL0xdwMDOxHu4lYY56dYlV0IPzXYbGxdXN6gkaOzJKtYFLUm1jt2Zu1w5DO
Bhqbp5sJ+faCUv3fFmtpCtDBkULNrk4v6Il9ONUIkIm8qo/M/Eok7iLgXZ6oDWcr
bmo1oOKfBDTzXk5TsxSSho/PWxb6jZgqKMqKvLuB0e/vAsvCdAYTB7KPnYkHN5jJ
3PKWDKhmFYcrQ+VOQ7EfmzbhFyRNtEgusJ2hSQEpfvYdCzKfcwQFUd+NtX/RMqd8
3uQketu0F6u2OZO8BriGKzDV5NLV8tItD1n1HB86OP2RicYlHf3yIsWFxDMxDNc5
eZtst04dMln29mKeMwnfJraC1LpQShm6UGIHW5m+9GDV2choao7nCPGmYcq9IpwH
c3idZn+M2pfgrltvW14TTSbKp4VWvaGmyHyZpWFZqQLKcbRqeh0/smWqzhY7k1MF
MWjHB3LE4bzu77nHYPpzIS/3PwnJizYIqrfkD/8RxAKPYCwLrmjHRq7sRzTLabgP
A6XfezpLMB6s9OmzKyMG8xR4/XeOWCxJcNuT7ZfiWlFRKUzgPx5vN2y55mFjDJ4t
1yzFSjDndLPzPUvfnHNe9vH3IfySzkPdQWCWSE6XZount2WTR3XXqd8s1snFaKPL
0eeLp5MyNhYiGfDEpnCyGeSsFd+M2ZGvzeAuMuOsZh9p/qggyze+9q+8NncMxkWC
eJ0D85IiJV/LMQa1oyclAmgry5OcGjkVldit6I+JbhpLSQKzlUDstvWmKs66u7gi
0p9wbNPfB2ZgaqBwThSDFl7L6ZejPXai6Cu9q0tVlYih306bRIXaxLAMGeSaehSs
jcx27Qw7792QVg4+fwFbdamEQ/rcqVR/el5ZbLo79/nVe9ViSPiXCiIX7qq+xSqk
Hx6v6n3/4bX9Ag3TcjrpHvOWYUizYsDQ5G86awKlf/SPeOmLe3mGyec5zCLvHgAv
p5f420XAp5oMTho2T19OXiLCH/fGG0Z5HG4GLMrqjOLZWFidsFkmrNg8MXmbgJ3Q
DspLJjW4UCXaXDZVd5rOAc4SouYF4mTb0HkeX5Rqg2lsEwcHJGNLQ+HMMGlkx5Vz
bC6myC7OG/Mhk4NhhYfrpLyZ3GOV3uEFhJMSxE93OYEtowWuq1/dKHi3bOQnyq+a
6Ib6w7b8I1uCE8ojGUZ4g2rT29v0cUlhzDT01A5bm186jDJMbVieFThsow6nvLvZ
XNCZq1gRCPYcsspSK/akyWYu0F7UpvJfLA7iquOuYz60SAcQzHHTvDQw6OGHO6sk
HS5+uHd3Ei9fcx8njwcnq6CiJPbpkxYrlXz8yBfvyl3xWo17+9TAy4Soely7PtfV
HWxm6pmejncMWs+20S0HIzjiF9CHZlrFjXbDr5cGfyJ0rn4LvkGgc3UeIzlPPVlc
tGxATiAZM8s9Ce0PI1/pRKMmEq92cBVy3/WnYZmksfHq49EpnO/9VjVhBOLo6n1Q
zQEvgeyiq8YwmJjgKaRumf4jRauTaQlvGUe/w/cvcw9rwbIj/T2Gl0qSK18C0TVj
0tI61DpJiKutEQseCg17dGy/U42zUNRCo5dvZulY9JATwsMgvGGOfDCL+T4JO4kx
hi0UdU95dl3g2YH2CZ6gcxyMPcJgOQ4rVp51uYTGUvL2pYTWdjdftWLnzycBaO4K
dpBtg7GVYVS1BowQdz57U6jCWoJ8ky3jCXttIMIAZKAGOM8NoorH7n8uP9z/jttk
5Ff15O0i0ffC/aswEe+2Nq4lWhsM0b5q487sI4QDSwVXARtt/1wjjnsNFQE2xo5m
86LWn+jazgDOR43QJCxZNkNzktMtf8bayGsidB7dy5IxEew5JukmB0CZqWkWjvoo
SE6hIbXUa3s6ZU6yAPMYTDx2SfCLjmyfMfDTiJ4WW/rwj/PTXMr7xdc8AWqv5Q0P
U476H/e5gylsSs0xKERXWIO1oDSRt6QIQO1Qyp0yNqWv6ZuvArIsYSyjp5tGarDH
qYId+13oUmvV+inp9D2VQZO8Kf4ej+NFWMp/QEOoEL+ueoP7ItXaXjNhy+fR8oeT
2YLxwAjzUTFhlKoqHOHJpsweslAXaUqT2/vcXZaz++IiKB8UDSWGB93sQlXA81oU
J0KsjwW+mNwXVYPgCjm7eKfw/2gTr1uZWmSl0gI0aDUNlTuGbXxfrllxS+4Fi66h
Vh9Zw8wkqQRB3BRX075pSNTpa8T4cmPh3IG//j6DrUO1LH9kMhj/xYV9yESFXfZZ
7qKL4QpJEtvrFvyDPJ1aV20wPB3q0iSrkOWmAyEdw7FvYoGUa0ScwTAoLZ9h2Y64
OsKMhb1jKHP0/OGMW1qYRXE3KZ42lkaP4Xj3o1hr10r0SBmp0QkjtKblvUN7rWcs
kDbnINgwgzkhP7SEEiw8GXeD6We9T2Ppji5dwJhNJIlI8pzDgRE6eSVdL44h1Ur9
zBgZRSOsEinwqdQ3CVcHrgKUXcqxvduH3vHUimFuxBgO3WYNX9Xfro+QlSmbBNoP
ngTd6aj//wD9zYYDjkvDVRiuNbD7rBU9xwfcRHmNt/o4AfBy4uZ6jEDEgBto6crw
5vEBdiytTuMjVOrOrZ7VgxbLh00MMMzMw1NNM6WvVOv73oO6DAJs+5f+pz9fHN/Z
GAEygDSumgAwRjW3WN3H407/H1Oc/PBkx4ELDQHeeQrM2/KpfNNhZijJFZ2cn3Ie
kN6H5T/GmSiGyv4AUQM+bzG/1GESf8laEmlicG+uM5A93ggk8ZypiJ0jnQQqQAkP
0L15PtH3OxXFYYpQdEMweFD6hYeZa7hpHnHDsHF5eS29RIhtSSV7ARLN6j4I2CYr
dwi7Cn/Msu57OgxlWPlPfebL0ZwwqkKHcgBjievdB1x/zHhI6/xO2mJtU2jB6Z6J
b5rg0VUXh54Fq4MFwQtiha0J4fyvqcGYphnMVTK0rJJy9F9G6jDr/ats7CZL35j8
Id1Tlk70OqYGGwPQ1KMWZ6uvf3QxQJZUvn8WyvLfkCxiUXF6PyxA280FR86wJA/y
IXwHVKPOJtUSCBwrbsRKXfURZ5iMMiZkaOXSawnk6zAOnj95aJ2rd1P85rvdfFxO
Fxk8LmINThEtdcsMTJIwhKN0rFTAgCuYt5KZO/L952o4UM//qYr0Tk1qTJVt+iqI
YHM3BvplyxL2lZJ8PEsEMAmNxE3Zm9obWtvKx5mwecOSOCfGC7TM8EiNFaCU9xJy
aTdgUoHR3TP+NcAPbd1yDrlcNWd1U1MXWNPDTX2lw0Q2doxElKcJzQFDm/APpIfE
w6NyAUZD3YpTUbvHC18CT4rNgjXSahSwCq9xVYp0mK6xBtvC2THAZW89EdwYm4LI
uh3jQYUODliSaecNoaKkiiPTqtXQxBzHMQt/o8vNMu/aOfzX/rkyd5D14ZZGiAFm
QGtvqa/jRY86GXfbLPoqY9Pnaiz2hDJPdjLkQkx94SP/zrpbazu54xpjNrNPkpKO
uscsyZO7TTu50Y8pCFOrWy0MgG31orr9ioee4BRYa3E73wZUqY+1fk5RS/Z5H6kY
JFM7s+hbYJzzu9JqfG74GOz4Rm28rj4kdNGODlIIi0HW10nNLuX5p089IRoHptvS
bnFgXsz711HtHQkXyTpNV7Lds3+DCYKNvewXEtFBai0+L8ylBnuiWRjm9ZkUvKut
4sHQ2sGLF9F37zXWLYrGhggykDKXALXXUcFGJ9giF92cevcDc/Q41LYLD5kgJ42l
z8zlGOHuPNpZV+BU74i3+03/27L+4mZwyFj9bRzpq2fUvihbK17KXW36EUZgbx3p
IcbnGUStZ0eFTGy/p22sKUGh/74uJcXX4XuuMHYY3/eQ9iO9JrejT0cJE65Av2/6
yYMsQ/17iRzrklGrr6mIgYLOJz2lkhsY7Bn4icOQ7nY7EIhkqGJQcFVRyZt99C6c
NZxuXjaVCeOnBWOE2rjnIdDPocDNASTdw9zCf4A8P4lsLGcirAfFF/Jt0H3ajCOj
VjjtLvBuN3LSmEZaFY3/FmbEZz37pMhhZ+8w6cSBtQESvJ+h7FYwXEtgzvZ/a67k
3Tty0VD8gADaivRiV0VrNZs2IGgIKiavjHQkKByKStzTw7xi3R77INwrOdulQnVe
uuwH9bzkdREw0JkDqtENATg7aoVtwSGtoasniMVPaHIZIdoyUzQe/5VWEb4JmL90
amX5u4P2pRd3xfm1jYlCFqtzU4n3Fsvg8FhHUeDxbGnnh4Jc2FuBXI6dNxjx813w
NRbmvsmtBtA73MWVICmd75cEPy9/iRySBPlvRwpGt9Lmmh/7LUstauLhlRrmxOHz
ee6gkkLIoImpyigis1otb6lfKRZMDF/f/gw3njdXet9G34T8TlAs0IlJguYM9llF
Z5jX64Wa/zCms5uIhzAVdSJIHrDG7dj9lH2hjAE873arkE3X4rNkhNdumYgTedkl
Lh7wOtk4NE0IZcncmDELBDWHFtQekhRuSt9Rk8Fqhw3Lw+7i985LhtNBfv5FbcF3
KXC1ko0B+lGhLQxtf5LF5GMHqEejEzg81NnMBP1iDFBUv0EwtPJdQnbbzt7aZwTp
h7yKaMtRTF48QC6+epDB1JT2YDK9FPFUA/jHUv2HJbmz+sAuB15LWrT5KSij4qqb
lQYGGOybyJ+/+jrAx7LytT42XNxpV07f9az4Wm96XT/mgH3xlmViinpVNrrLCf52
Th34++0WvUQhgEJNCll8eGA2A0hQPQT3f3t1Je/Z5BQk+5MWphL5jy+uElf/2vhN
Oa5hQuHMsGN2ERwpqlHon8gBPOmXgpJIslLGfLOudEEfaiT+oHn6itxdKceCu7+V
RsDQ0xhr71W73k6o7L5vg2CFKjILN63+gJ25dOZLGWi99pLxtIYKoNu4ZmpprYve
EB/1H41Q0wvXtND7FMhGIihz8ATtjMmgohGFH8r0YhXJrtQKqkEhgKrOwQZWfDX7
I7ixzI62YgezF9MHXnUWJZNoHrnxEQ9jiNLvcxKSX8N9pU9E06FyIT8qajPi6ET5
p/0A8MQ5BXljvGugkDfwb8BkuzDffro0imCu6cHgpaqt+l/8Ww6n0dCL7h8ZzFEO
i14GnOjsyY7yjoh89qKwUSZg09koRDpR20EG8FCN7j8W4X7fsxlEv4JSuKwRU0uN
QrnW1eyIW1XU3S57kVRUttREq/wFY19rg8A3/0/dvoZySWtcYudD2N/+Do9xLLWV
J8UACkzA32SFGwCSwqCNGluvwoIpv6VEGOhq8tElMe5gZ2YyfmoCtHkZuapvuIsZ
anKhGsJR9wDy/dO6obin7qUq78f2wBOvOlPMWm0916l62VeYYBEVY88s7UXgYhCF
PP6dcHrItm4JcEg6weHhJFa+bN24RI7oq01Jsl0vEEeyYOzweJ6Y+wC94xJKBJN9
0Pxi/FM72ZVc/Ie/4tb31vxWW7Xcb5ejSvg5ZEKd+zT2OVd/gLKGAAeS9KpILkG9
2LcPdZ1iT0c258AEqwIkesfG9uxlfz6V+zA0H5oMtFWsytiH20gR3eMdUNo/XDPg
PSD1RCQKtZN6/VtWjyjVO0JiEYEDUmNznC16JNLYEycAi3S00w5PIAgogHaFrh/Z
PJnNeiiytGrPV+KcYeTJ2P6cpcmaP7RlZbvZk/SM7WFj9WGgZgnhx9CsoX28nwGc
aqm0WGefujDJdc1+ohIfV3kga5N9JIfYM1/EmcWCRr+vR5BSwRn5gT/MdctmfUuc
5fT3M8COZOPXVb8C5AeaDe4uCvOV8BNgteVmft3Pqj6o6KKVuRQgeNl49dXn9pYE
uVQFiEJWOX9Qbu86KHMSqvZ+xZpv+zd8v17p1TKtFZFdr3CKanCOvM6kT9KhrGYX
wKNCOHEsBxek4vskNmPBjcM9IEH8ezcvqNdPng3HrYbeK5KUxD9y5m4xgRsEkPm2
+gtllDETqNpJZKKkVvaA49TcHzNfOeGuoxYcWJaFq/r0833qAiBcwQCQgZp7EezS
1JvlZQX4x1GqR2bt/dmikewock4tf1Bj2KGjdFHUEWpDGRnVH6eOBm8rELYWCq71
/3SW2P4W0kEXR0I2mnSnqtw6EdM3+XtV28zy+BuFXPqRh9D66j2Xa9u1DZKm7oda
3LSfmB9z3WhIqCE3hWAGm1lkDqPGzir2PhJ2WujadXGMIvokf2HCtiv00oxSH/AV
IQSmzcxjOBP+5s8J/IXV6GGP9Xyi7IM4EfezhfOQWPv/tv7V9djf6GJOsJLYmJo2
dSBpDwR9RTVqG1pBZMXek3qZKrD1NJ9FSqJF3BwYsblAQTvk0cDentke0ms2tvdy
AVLWmDnrVItQYKFreSmex5RcnhO+/TSPR9sOf/UvxjgJyPWtsC/WfwWR+BtkBSuR
gSTEZlo70T1Ao/OFE5giZFEdsfJAIZBZbPRFrgK7va6QtpSkCdXjCGPOuw7Pw8GA
pI3n+Taby/Cp4CqHerCOf0mQL+s5nKAmrBXEA3Aya+kChJ74eTShz2ls5OVFMe1R
ncc3sRPjQ51nBcjztvrIFRLCXKA+hk8FZSsvrS2fAKbAV7LVPAuRPtKad1/Gtdtp
Q+NhC1cFPlZTrfJw5UtEJSTkIuKTbXlROIVzB2x9YhlOeLt6Kok2JeF6c+jEw1Bj
5iUhSSGtWee8/PQZSl3pbIvFxWfAKEc4iYvhwPIUxBjRexwEhhWtdVlK5OkEf5pQ
ueSgGZB4xYsq5MkvPj/At2Qr9TDHml1euhIzPKnEL+pOTKJKerpR4TzEPOOVKgHR
NxKNPYKMu3eR85srKApGmAOvj6cTN7B7HnNya0VROteSH+QL1L/Qt2VkbeYDP+6G
YiN4BxbBxVaBhJEFD6npkFGrAartwO2HzlzDBbe2lvL/hYQM37nfaYh/FQZerrWe
MX0arBxSNdXnYQ6919gUocL5tGK3MPjSMRANhkNCSeY4PR3Mmg5waZ5sNh3tL1IO
HmSIVMHbPf97RQacKwwzZrLDTXmDCUtTlYAXoOnNPqyy/7BQhxAzLkLgS2B8TAqd
o7BJkk8TkYyq+ACgX3SwVg1YscmCT8hDMUoF/uo2JTZuIJC0RNfVGuQOMu2RutJ6
Nfn7Sfvx7kzxchRknkvggAFBL73J1i23RxAWiJo8nTljGq8sWK08JQk51cpUckzw
OXhzlbCE098qKvQhlcR4tA1x9JX78x0uoWSOquV5Hb08d0KtmNeNKj/aNSxJFRhV
yZQiefoRFBz9Va8s8k5VHjollyQeOL7XoRVS7wT0wWFq3L6VxT6qhQoUV+ecM08W
Mc40KHQM48uXkq3AJg2NU+9Bv17vnsDCS8aad0Lcc15HL5oCY9W7jTuyFabYXZ8T
q2PXxSGoDIJT+Lhmzc4csdtdgklhtKsGzadxauTki92haBS+EFHtWFm9XdMVMOxU
2i4e4Irf4k/yCOJWOPk1vpJbdgyXOMmnazvp5npnfEFTKKBEEde9uUc7zmAKFNio
wJU6Nn1BDFltUAgJIJ+BTARo5PKkUUvfQRSbN5AqmGQld9TlW6gFsMQQS89VVi7p
sybnhehgAXSvlML7KARuCjgxeN0NBHgqcgM/uqLb1zRte3A3HGe9NBfHr1WqIX1/
LJhymdQ2WY2QxoRsu99kTruGKo1pD+Znoj+oTeDSf+77LiAp+1qOaC6KQ2OExb00
2yKwMu1rUbS7t+to0Clra7rJHcLOIRi5hC/SZ5u+3341A6AOxR0//uEvciRBMjRt
hJxHvzEUkxogMfRxl9H5omrxOSFBhwy976YSVGm0rM+f+CfBjNgvH8Ta4d55FU2B
ClF24BTarxDKFexLl5zFPz+JiVW8QwhxzJ0oATDZ1JIC4Bmz7l8fkbp2pCBmGKFl
3MvXFrxZcrnENkPY6CsM+MwLDlrE94rJiWiIMCUp7qwHNzUt8JE/xuVhBf/n12ly
QXpuZzNYms6QjkD1qDNGCIco1LcvzbkddAfi0PuntgWKQZTuCf9ZD6opoSaCX5Xw
mp4Tt5UzS5JtYeJFzDOW00DmqPwd2cDkE3o4m//AKMD5TzbWNLKthOUD2eZQJsgX
nsi0vV9yNouSj6JdStqv2hq+aWo/llhzwYXGRMPtacqscna3jn4TJI0WZ9Nf1jEK
I4x06cx5Pg5qf5PptxX3WJi2pvSzXIUB3xkEw4GBqxtd/2zeW7wIr9zw1SQ8Ounc
K6Kt9uxpV/cs4JI9QGZAmWMjSjeOQ3jklK9AMbhwzECbIVLGEfqBbz+IyCrZM5Og
PBn/1oiXo6dv3zGVr1LrzRJhoVdkAd7af4ssmTaZkkFGv+UBe3+OiJRTXp1jYHUw
L7IXwJbf0Ann+XP0U1csLY7uwIDHCybcSdjWt+fkne/2fr7Ro/sFyYd8I3SZhkQ1
tQHGw7IQ3BAtPq7wqtHTqEJqjf8pRwoIr3/zSPissFvwGLzA3+Tw9lxCA+9HiIo9
dzlbZ8PohWrlD50rVcX5Jujp48wiK8gYHM/Cb4vnnyCHigk/1F432w9vRTA4BPet
aNTLgECbrMM4X7mFEmwzx2T2WNMqRyelhjSlZdNcRMXu29baUIuqm5jmsLy0aK98
QiiIy59gqMwrVU9iBsb7/Z4IGH9wZLiA5nUE0QpYcvNW4vB4IJTn6xzgvhjA5fBi
IbjEhvchmVm5IETqJyi4cEbeH6rZyk26x1HMakv2xtry7o8uhb0FzqWS82aCvlAK
7/FX3dyzDh6tMXKDsZsAJfXYTXkk9Eo6nAlAX2ndDccWgqnCM2SOIeMmU8Bdtwdm
/B0WOW6w/vLeAkOfN7XVdfSvpjOyedgcNMVfmTotJFmm+VbHpJGcbQqqBpIbnW/G
TUyf/YxzG20LCZNRFKAFTmAfuMbeLFOoMIRjP5ZAi2Yi9pAHgwjQhMBgvkCPJQ7G
FoTPNof6bTfdkiSRZrtBnaFkYm48OkNcdfVMepjJrOfiBpYIdkeRqx426wAAyL/m
rv7pNFilTAVtidcHfkMyayVco6Z6L2/bcTPNr0Ty6iT2B4poYXa5Q7OVCwpvUzyI
3dqc4x29adng0lrasqrBMZuFBBZTDibSrchFo6EeoNUabJDV/pOR55Yw1BLsTFc6
xF5BsDP3xCk2wqQ1wnjO7aksVNRg9o+elSK/nUrKfihXGgqxEvi7f2aAnyWyS+Gp
dx13nWduTvlPtO10HvG+unnRnyBa3h9qK/5CdcRIyRuPxFMxqIdMvG6d+qOU9r0b
1NowRNmV9M6a49AokLL5rzH6jdLikXdgKyGtiEVzDLwEb1MozvgUabEXele1VAr6
ZWjhdtC98LGaZSRi6Urd/vpJi+8A5mH8nN33ggzsBx194UkR6CI5ecU/9ovvvhRq
7InBveHUZILlhRG/zAO7Mxnjb8ahJoUiNuhDycM2B9bMyZtpyj3pU/5kDsI17i6V
66ocssw/ZIAKUM9USZdpktkOsPByYxOK6j8kU2SRT+HpSlI8lEU0iSko1X0tjrvi
p9Cyisx8IHVnWd60zx9hHhVktDkIfov2wCH4RIEqFN5KuGiv6IyNM/HBLHD+MmY2
AsqqYFV7lqUH9So7vXIpEaB8xn3wPOWBkMiLomDiqj3HO5RBR54OLtKprBSd+6rn
OsG4tfN8DcPSzURxr5Q+Xo0IDCMywKV6TKmSMHyGN+tfyGoT7awcEUOw5c61RdDq
aZhvcPEUfzW8sEGswIzJGClKvBk1TwTBJxTE/2UXdVVxB9cHW/do9XsP5Mm51E/D
8k5ZaXJK2uYNQ3U+LC/hQj9+mRaXtwMque6kj66dGLPvF2MbfuyXUcrtK+tuLcUD
SPZ0jvp/l595OixeKW5vj+hir8eVHVPyQDrssE66hLJQmcw27nRu4asde0485Inx
I48Fyg8gTWrUOLQYqYhCxdG8YA7Nr+b6FVgRHpYA9qasG8ADi9to3WDedACuc59H
PBnV4TU44orZ9C0RSo15F8PF8Kahmavx+7ZHvK0TudZf16oae8aNiyI6rUtK7fnt
U791G7sfpfZKI+4l7IxH8h0y1thkz8v88WKy1NJOKR53X/+k/ykJKXUYFk8glJq5
E7bVbjRsTvJtDzN45AJvCpl8E/p72xsyKZz9AfyYlwyU4GsULExLXu8Qr2XoeA5V
HgZmK+hbC3+wW0t/2mwSlcTEK9HdS2s2fSN1uCLiWolwusl8T805Lg+gNZac0UfU
dIxuDWztUIa1AeM23QNsDyVKPmJZRad89FzZayxSnjh7opqopDeyZQ4HbRlUVKw0
sJkY4y2mAyCqK7Yy/sORBrD3XUS9vGw2S2NT080RQbyyitZpcuvcX+m6M/n+RZ8V
qbSYF6/UIfCVDrUmsDxocpsnMQaNELWYINRUi8K4ewkTFhEXA0mPbATM4G2XBFT+
AnhVAUkAb92/1ZZ8zaOLpHknNBCKnV2oTOAhcf/wMIbRGCz3bg/yAqr7HbUZB8ih
AYhaxczBC+fJ4RK+1WNOCOQgNGVKw5bZCeYC5+4xLRZ0ggxneCxUDXfAx/X9Jb/c
2zML8grk4+q+b68fA/3pX8SUGZO3H+HRplWy2jC5+D4iKkYH6XLBN8lq9l4ONW6k
LtQLuh9NweTXDHJepg+bWAy2uw2/oqlEoCG5GdE1koCffee6DMr6OYYq6A7WQO4R
ys86p/5mYoXz2w8QEN5oxLe7uVAgUkjhEyxIik/A1/fBHJi9TAvSK9xs+jPLnuEW
Yfp3UgzVlc4S29v+8NVZRGnnzmRZZ6YnSu6M0pMFhmDEwuAWd5oa/E/MGpp4Szav
VBeLv4jSnxmuAjk9IFp3M7/n2LoYbqeC3BaU0d5Xlb4ESB0slhE5AsZLyJLYgOO5
ni9vQMuK/02NvWhMuNBcZ+kb4obZxaWqESz756JZX0m0PGz5WOCwngwrYyjn8zZi
Nrm/sjYJNP4MzvHDC3jVnVBCGpRDQdzzeeRfGJu17mWOtyVre2DPHMDuuHeRFeq3
zRNpZtyL0FxFeXIO/xE3PKO6OqPQZL86Yshp9FQA+y2WM/pShQmxWrYX2fXHnnpq
M3nmhAsaUjyOQ4Ffu5W8xQaU0zZgEY//SSWFpFYu02yYtrS8h73yLy50WaAgYKOI
N/ynSjyp7HEps/yel35bE76x8pGLonbdHx3CRyEfnYOc/lDpPFG8eyin9uSgmegx
jD7DM+PXyE+98/CneUxh+20cZhl3wSBWqq5FRTSxgfO1xvwgrpjUiuBY4iXOZ4Rq
nJUksG2MxH8vTzTxT9pYDjYMuvffcIxCZthDGooFn+AvIqnZmooqslRr9Pu5n069
z565owwgcYAD9LUwkNXzuh2Z6bXNQ8hVz1GetSokIwEDFX47lRUXvYuOgwCaGqBP
I0r3YaSuR7ERkvGFFxbTr9P0YtgGczE02Qab4vLk/URJ0zxoiJ2IRUp+pw3pHUrb
elmpBLX4hH+Ujk9txneFAsyTHcjjIZPXqx/tEgdgWSRU0d1Nc79Vt30oBuzUkNHB
hX8B4kZrOuuYM4ZEU4hVz5tjSyB5m9+IcMFXDczKwdK7B7mDryU5WHhSWDa9VXZ7
FNMm8iHK2RAsEPmMaBqjNQyRTqcB2aB7HlAg3sHuWUAA5W7dH+fr1DeZFDqDdZWA
EwLuDzCP7BhIrZCezATY/JZR6t/FGmy1KFJgJKo/9VVeRZuDPciuSRXKsbLSkqbX
3e84NKmtlHQCOaw1ETCu5p8xUH5EpEReMyA43BWYsGrtFiXmjyFg1H0tYbi9spn3
zLp9bGcilg5rMrMfdXgvoK6A9BkAb9GWPlw3NePR5lDJgrutg9wkYahsFLrdUhDP
6njij1wsb5zHzQGM6RlG/+KvZFvsfz+v5K3LUAYwXqpiMLhN5g7Jot2P4Rn7nGwy
iKdrNDWbZscO74ve/nQ/6JriYYf4OjvLdPG77h2WcQt4yLAWM0Gck/KQMzemzaqz
eyydZZcr/V/g2pX9Prv0chzOkUXddNC+otExDkpY1zoGk3tiXH+tG9lrZ3jnhmnD
ZlUAcbt5Z2sNvMPp7HFc08fHq8WSfNR4SbIO0k+jVidKs5r81gyiN1kesgn63e+M
XGHJpFBKa8T2Mdj98WqilWxeNDWfwtxE4YEAwwrRScQ7Oam0VsqRnQamIl1kQ8kO
qsVpAsX8u1DuvUOv7hmHjIBNyn/JJh34OKaL6wdl0wu1xULdYVj89lgyQX+1iCL+
531hxUjem6+eqJWddGyYLvInfJRlgVK+vdYs3QmP2szoP5DRzbrMNr/5EQF//+LR
nvOuacvuZxPGYQS5n+IWcttXbNDtwpKFB/8Mm3qX0ug1nhS2wkbjCpNKAU6dX6L4
YFiCgiLTF+SYGKp6WQhL1cuz93vIo8gft/slCxZHY121D/olMftV5DBvcvviOlpI
y7OOaJvF33FMeIZzS7Q152zHI826km5ByZlUyThv2LsxVSxZFtj0EX0fJpyn0f9i
vGbtXg3U1PBKH1LPODFTUy3MvTLzzw6/quctGCg2q0aYgs1pRQidTLfMFNV/5WX0
P75juoet3fNrx39QdSk/W6JbQ8wuKzYx5s1DS9FgQhtCxpz+8vXby4l47GoxAxRV
P90CNBsS99ejPFiufnIjlMz4GCE1KXkInlVlbDbvHd7Zg1z38SzyXWUfYuQ71dmo
sfaJByU530na88kmUaRzFOzOTjQuxe6litkpkMzn/dT8/PKonSmeUWTqEVENcj3F
nD+BsVJ5cLcRfMakB+wGQZL4TXRq9GWrdv/fmSB3G6tzrRHxklGb69O/IVkxOwsO
BnSfX61Gm4n9V9E7QXrSdmEuW8ZLEhfEwyJTJkTylT31MFH6lW5tlgjgnrUQX45Q
k6EwgkteiQ//WTdXHB4oGb09MIm0y0iCe5cd4+uAMA0BUPRt1JWzRavxfPgkZAM5
+8y2Bn61NPNcaLWmc/Nysuu9Rtq/zZWSPVM5o2cxQ3ZBSSkdY0xHQjNDMGxB2MZv
fVXuFi5GGYLrRlZ5NoEKDhk+qSkrVZorwl7coNhpw+GmUJF0v0FXokFLnux22jQw
CkEXkBuitJnmxpsI5O+24p+U+bv4SV71dcz90WngOjlycN453CcSH4RWzDwhQi2n
o92cIPSDZO2HHl/Dmz2vmr6Xur0Sv4pvTNjI3f7fpdUa42cDA7uVej7wWRi6G6b+
KS5y9Jwj1CfZW9xypQGO6KI2X3dN1SCUAfMd3v/B0LKZM3bE0nedoHYNU0Qmf3xS
w+wMaA8SHIzNK1iOr+4fx9p1hakpP87ojMM0I5fwdbmUc7179MIKGosJzPqxWJjF
dbzBkcOQmOq6txOdHp/pm4mVOWkgc3QwWOfic9MXH52mJ5rEKmuCp3TXZZU4Lb2k
ZwiffbcCXgrKIiw7tPxuoh6jf1289ogKBntPD+w8G3t6qu9No4UMJJ4ImO1NYpMC
s8XtFSGMobXzMykl1wHpUqIdu23yvumTD2dfu9lfr6kKvbYJxbXo8oJgjnyw2eR4
oDtCQa4vU9Xuns4mMZrax3wfFj89oj4r2LlKoEw5Oz5Rb2SemeB9/hyDfDe56g2N
2i75cVmhgucBAmk7Kk/CrdTqozF3ovy57mCZsQo286SwwNMKI+09ouFCt6jIafKr
SLTZmLXfg2g6uaoBtdk44sGEJvpRULpbZe9lCK5Zb6hQHsSE/pR2QOvkdXsbaEgf
/4y3jZR0xOSVfiKmGeZXCXk320oxqlQu/cMFuhVckIX/xieBA6Xp4cXSd604UUQz
V6xMPFqDKsEymJT7tQlkO4jDVpw6fgzX7GcuGp9NZYOYli3pF+kDoqWD+bzK0K5d
EYTBvqrW9RHjdzYqA8CtOllog5nfgQ1OAvqoitB05/2mhyteRUJEdL789YflQ+hV
oE9BjaVwY0H9gn8aGx6Dw3TwbdXeluo8tVBQyhw6zw0DMpg+NIqzCkMLTMEviPEY
vJUR1VV2dGLCsZSB9APMp61T8FSqZb1qqvRPxNdtuRnPa1A7VyRjqb17qf1mIe8r
K/XHy0g3JXM3Jmbd/8UXyZDQOgBVu18OvLCmtezr+WQ3kmNCFcvYhnQgpayNTK9R
kBRVLqDSafYj5cSbm9luOfhHZIgaTT8cooYSoQo/BgPVMi+ZzUnUzGXeOBrya+gm
/1G4FjjBDE74++Y/EYlo2Xo9B6wxyiVNMQBOA61HH0NQ2o/jhXnC7k6R8egeCzQ2
DirwqOyoubGKR2Z3u0bdvoXhQxd7bVvHesfmIhS6D67wUeBgGXDDVl0ZO2G5l6Nr
nQUx7pvXsAVq+zRafz797BvgjFfyhAdfBQgLSBHmrilhaWeybsOG4rLcy3QjFMjm
FsUw7Ce4mHoMcZe4gsa6/UkuCvTfNzkKJROe0p1OJTsUFfq8PIQCPBlwj2eh0NQi
pxIGyYOJk8X359zBy1XV1YGFFUXUk2xj+SzaLWTdmC1NIbpjPwBzIYWz7s6FgNu+
/CJ+g9hks4KPH7c6kGkS+apjiG4d9SZKYPKPQD8v3wy1u+BLWjKqqAnkOXlxF688
dsSxIFbrDxepgvpKi5smylBQwfPl+dzKPExsqzTH8GbUbRI6HB1YNkYgznepEAnK
WYevsT+PrzWjbgr3A7nVnJmNPC3CCYhIeT2I/PMtj280t6Ai8f3UyiaRc+tToYtZ
1p7nCX+sXH2Q7glmYZ2OrXiGX7uzDoN69ZfxxaNmCwpvoRwL4cLwhYi1XVcot1Ph
AC3Zc4J3Zo/I+3NR1bIQDsTglfL+ntLW8xXzN9Vih/jDoVT9/QNg95RmWN1k+Iss
UvYiqBsTTFIRDthLfPjUiZWLeT0SthhkjwJSVB8EspzH/sn8g6LHLtGsPnXfI6ac
1zodmrZAvgNFnHxUaqiVmsHg110MJ1MbDjyvhDPEL9O/QS9+00TFZi5+4DVj/UhE
CyOCGMjPzkqdEisKu2xDs+n3HQiIc6ASZMV/mmu1s3le4tVbAc1WHgl8YrldnI92
PYyTTdO7Fjk7Ut4YDL9A/pakHmDDMH8DgwJ6WonM+wFPmE2GmBR9whFux2RY+Pjb
POtqcS8m2WjZpxhWSR8ln3tiB2C0tA6S/8upbSfnpcUZt90neFymyxrua+LhqUah
cOymc6dFgN6tMPWnA1VzzSFK14emmZ/lOG+UbIgCWjVV7sBFJJ6VgUTHz0n7XLFZ
BonM/qEuuJiQCrcgfCXUqXdmlWAcprNJbUAREHRqPKO9+qa4fjoCxPN05u6rFUh0
+LBrlQADNhnalVyLLLANQy5wQZeieMYPknCW9gv1Yj9thHy2cKoRZroRpSHh/z1p
ABe9wdbiAs0hmUs1egvNK4hCHshzP/lJE++a9ahLsyCUEuni+Ukz7kBQQ4281Fjb
UUTdgvz/ADN11YmVkqS0HylULBPEnD/viGno4Y7wdxv0yDmQimP614N3fdYGaF5Y
veRdue8ZmmiAA9Z51EjxEGP0L+5/0ua6BSyfPccMeZfRLBSPNxqijpcOnVtNTuEY
9L9xjcAuBMOnyqQRP1hpgiy0lEErtVt2lmrGCujVa7uDt+FSUKV0Jv8jIjFFPRNy
O7jxAhgppgiBNUTqR6Bxfz7VXKJMZYzOJYkHaeiRKEzQ1+MLJNkVddgd1zix2VX8
e9cX7cYZC6Z4fPRXBK6UDhQNjRQrSwaWbW+gKBReIEXCvHuBU5m3NtGsiQwnSjwD
iyZYp6bPTJKe1mrSJK5bMbMGhSGQ25oU+LDJLBTC355puWalu3S37Wl770FFVif4
2JDI2vDx+E8rtvWV71CT2js6RvJ3wS269E6f25B83gFPdLApeAimXVyL5ooOV29T
k8F1K0seeWUqWFBiys42yx0iKo6HnF1ThzHhjyPILfcAiOTIJKMdtGxz9hPkg3ZH
UmzXKrVuWVj8cPe7gK63oHJOl4b2wGE2iMneO4ABmuaChfb71NNm/NwGb0ln6+QG
zdt+lS7+oLpvwmxNDvxx5nHfPK/7L4No1BuxwKudO3Pzlo2FcgWTG16bxww7pbjl
TYAWpGtB23gi2resd3KkZo5RCptBzlZS5GQSrwVLfbt3MmO5ZpkxBExsqUGhJjWX
eXeoa6wbXVupqo0NnUQsIezY00ryOKTU55eBhOgUMuJIFjsY37yQajYiYJHqdcwA
T1mJQmnzxQtiYMMKa+wlOMl54Pj7guwe0UywV9zir8Cx01qcr7DWzJM+0EoPoZIi
xZM8WdJlgpoKKgpBNnamg6XG5zangmbRbhqZSqtq2d5bFMXyW/A589C2ZvWcbgbH
N3phe4oah7md6f3Ls2KGEa8j20Jtkz6CuZysgBWaCN44PawhdnVbTt5pGPlziEM8
FYzjINBCz/YgUQbu6FpLtcw99SJ1Qr8Ah8hBnkaJOu+vhjqLRsvuCH5hd5E1yN7m
OqqpVOGRhJiQD4z7+DJ2KHOdL9LLzc3t+ZGQhoVXvb9nFhQJZjvkRStIGQc3M8O9
KeGXSNOUFeFGMzCWbvWblg+cA763i+kLi0+qgG3uc/8mkXRUdbIrRkHqvqYx1dCm
7+sHXuFo7qaSua+NM5m7jzdKTgLSaPdW2kmeSaUQf9g/4lyiioFLnYHzf1wpIUUo
Io+M7dHuGCYL3mO3MghQRcLd7fe09tdDvr9FX5JvX/Xv539GyWQDyioGb4jE9k41
6rJUs3SVK4JLxcEyZnR61vYaYJYANiqa0VI7yn7ehBvLpur9RlRL8LnJVfF9HO0t
1GBFekULV3l5yRqK0ppn5Bx/Z6vRt/Rw3dRVsSfaShmQiyzKAtPEgvpTcv5pytl8
txgnjgrOZQe6zOmRslu01FtPsXtJxvl25cF/ySA5G/78Th3VG9kxLfpvmLFJVozf
DuUyScgsGFBwePulio4PzXcmgBeeuCBTJbnJ5ir9xgV73cYVW/N7L/DGgOWrWc3Z
oN1GylQv78xX7x8GK43RmIIhiknSJ4XcIAaR8QvSY5ojmgOURZqnUS8Y3RbHRCsI
0erI8btXs29QC4rIdf5mLsCH/7xReTUQC+JsQXUBj9SaDqet041DwGIQPDbrT2ff
J0AIMFJTU2yGsg5TrKJY/do6k+Wr7M9EtVae9ZoawRUmDwmhUsxzDv4O2hl2M8jc
K1LBcEVbSQIsGEYtrkQE2pxcyPJslF0rTs+y1uZ1jRxdkbobkmEuABO/gRklwgOs
MqUooVbYevLNcl7zUVN8O/jRBNDU0YqTGzPL1CIP2Mzlq1SyKvX9fIajCXsPAWWM
3CcA2i6M0QkiEJsItH4kzMsXQgQhD3SvJ864QEhFrybKpmQVnFkDSM+dunPBohs4
xFFPEWOhd7iJAKjMhz0kG1+SUu1OnWb8L9EEqpRiksLaetuCRqtgnI7hLmEwGh/o
VjWNge1dgeQnpiR1hg+PwsvcQulKo9AfjvfDIAxYfdNehAC25EtIsK8sv2kg1n/b
539SMn41fP5LGRyq/BuDQGAbD1MXw9RuMCyVaaHNkuV/fb6eRCuVjUyEBjo3ax11
dEdxl0DHCQJzOhyaGed3/lKUTIy3fknKLTK4CG+UbdE/TeNwYIfdPj/ou0QkDMNH
CVr8wuNwduU1JWUJ7Kt7q47MY2ou/owEiCNINAvrKmwLMq4gz3KGsn4TEdP93Y/J
BSVqt+yfqhEegy4BvMR8WJUQx2ffxdo87Jz4D8mrQwK5oLeKj/w9UaAWgzuIv+5x
30V+WG8N6ePtKoL2X4wcMzfo/VbayEeA26s/HE6XJ0TmsVyWeVYtKajkAopC5N97
oKgUXP54ZlmH8TQMJ2/Z47enZ8mZA/Uk/k/H9/w3HVoZprLwzUe5kAyZxz4sv+vT
yoH6Ok55K0v+34oIXqil/hqYSYmaXW+M0CoLBP3IGgU9ynmikmOuSL0GAWaK7ThY
hwgDi79tTEtQQ016/o/E1reWqeX0pazgJQgnagT9NK3fRyrOH4H8ciXKowrUvbSq
N1uMUerafeQ5iiFL78s43Uq5gXieGuFTzH7MaKxpBYoWbMkB0seAt/WNXK21PDgv
H7wcypAxNkm3ZMGAEZYTqxAFLuqWZ9dm/sRnAWKrJA6lm/AS9zTn2XzdoDJtrBE6
aEreoCO0Ld876NpeMn9AKtsL53wQqsDslKYHjD0mHvlV1JqgRTGisx6H3xyR6xrQ
QT4meBs4ij4iCIR+ZbVk/1Mpu8usULrBcNS76APXlyK6D65xgRSPXFNT1B8iSS9J
VayMYXl2Jkg4QIBDh6m2UZzBvPemxp4W7q7UZOIUHof04NsIbZnfzkqvb2+ytI7q
7gNz+b0cIrmH9tCV/f+KDM/5MjhG2QTMBlEo8S1hfNZ3vKm4HHGT/T9tl8j/tDUi
JrMNHVi4zkNTeklcTvSM//LoX2I1ARTibTUonbiURyL0ZAxYJ1FUZY7/s++d60xz
MJI7Y/Rd43IFDeF2s1dZ1qYZ6rlDWt56B2Jw90b4GYrBN36K1eI29AJ7KvX6/koD
BYwqdzfT9LNG4fSEOQeQN1Be2cHjhXqIEaPVsxRGWsMLLt7aKuoBIJBJNwVdCqsU
t8q/32C7+XaUKL4NnBMugOvVIi6KI0gO8cG86eUX009iEDci7Ro9Qpa2nqcEv6Ik
5hqv24mxd2tTR7ZESyxVFkiZwWXZmgNx2ySFUzFe6tFWXa1WP3Ad7a2fUIqJd78s
aPRPePR+QzQL4NyDqSwIK/4uIbgCSeFdCwflKplOZEyRq/NT6geWkJjsIbjJsoKf
krLn2OO9TC7xlsvB26jwh8aeWWJLeKyXROksWZAxmkUffrKNJA3+N01MCVPZFVkT
fT1OUc94QjU7PE1+ZRaGrphXRnndBvV0Ru+f6felvB2ZB8c/h5SP8hSsb7J9cgf4
hG8qLPjspGafVHIirMrM2voa+I/oa+cna4D6m3b/vfmR6qTpV0iCk6KMHYHx+W0J
DxkEj6d4ObQP6qqmi2cuU3N7LHeEGni/Cmq4JzVcGiQibCB6xwPwBFRA95r2g5/9
kbCgT3o6Ka3CsEYTWcDZrQgc9Kg/SeU/G5xMMUKVrAknR9G9WNDmIXU4x9VwRsX6
O7qyzbxn6WcQv219KrH3NsdtCPJDDK91TEe/5UDbcE6qr5IaMgF5aFx+IB+QLcuJ
GsHkkvFSkK7cMg6c71zaArS50AaCti1MuZAG9niV+GbNDFGlnUPIRTO/ce79d/tH
ZHKH7ojzM2pWgJG1SkKe5Y3wXs3ma+EqQOAs++hTNYfneK3G49a5qFeTupB9L/TK
Deb83urFhBifhKroKH8NdVs+TElGOi43UkNTIVVLfoybwJoMdeFIvZvD7/x88DLe
4zB+Mb104j6MTkFt44lLKR98VE20WchoIVAe/yzYmHf9wJS1jxQ8YKnsgSmv4Qs4
O7ub5GIwMKdCpbpNMXIgunWjWnLkdXYbRoFPjBs7UTMMM9uOhLjU42MpbomDqW66
SjbilD8Xmco/zBErTQA8Rii5RlCEgIfy+YngoZZZUgSIiAiV9xOI12VuFEE273D1
34Usp42meHGaM9duVhAT0E07WmGvtKXN/JqleVLPRkrxEWOU++MskI+c4GCJWXQU
x9BvjURR8/tuT1LYn5VWslgI04TbECl1972vC3ZIz6SjRz36PyUnT4RGbkbXWCu0
tzEzCHwnPxNcRgg1v7fiBgjvZg589QIYSB0IsTS0jJYLAUmkEWPzodmfMuTKPuOA
vGNQJI71L0RovVX1Tqy6LriMM73NSsFaSmWTb6PT/sUKVMa9T2opEdEQsrKByzd/
Ca6/YKiZo9LmKQnpn046NlvyEnUcYTfTSeBpGhIhT0y9IVtHvp4JpAgBjvLifLJO
UXz9PRTxzzBbXwHMWzs6tTlw+31GF5zWPHCspRVIy5js1WJ7vlAdXDH8jDP2OKTA
QO0tJgz8L7tKZ0T6yCMSEhjNUpJAfB+y6k/lrpH9e/o12FB/whTMWv89UOv3s/Jx
oNXXJPFc+nQDV8rRf09j+JK7EJojjFAN6cuFoNPcTmyoDszhttg6IOHoWBqUObl2
yOyha5oaHt5GMPAy0zWl48RO1o0TUAIWzb/41OHgouN/dbhdVU8JjNRODAesE6Az
476dUNScLwVBaBk/MqbaU2swyQgW7Esik56A+hnCgincDDvuG+9W6CYzQCNQtxMA
ylFYflkC5pLnyXe3oXw6asLUhmqhprBQRpVvC2r76oakgkDSC+7FAXQZP+f9Ft4w
0abuvzq+4RdvZdO4snmaD7oC7NhXuoYHKcJO/gEWAe+K7J6zBWriVWmU1kcK5vl/
OiWRw6O1GT1Mifjk+oad4xF0cDPgJdEYRs70vjF7eO63aAYtFDsZwSlOS3ps15HV
hRLdCHW1hLSTcCptxxZaUs37nwNaCRY3Yo3eTxtGTtVANXbR4FRQk16yaK+iN+pO
oO24SfSM2PRw7Xtemt7LH+nP4eRlI7i2DyanIviKn8UR7rZd2ssMrLzQWD+f/2RI
CJQIDfbOWedgu2ZJ0IjAkWwAA/nW/PANDSm6yEuevz1/trwYAQNNk2taiwNN6+lz
O5DkvcCWhr6Rm5ERW3OODOHF8Q7+EUCmzIW89GyemMqk5WDFKvd0NrSV0XZ7wSsl
2quuJZyqfUSv7v1/KmCOfS9x0dZ1/Qws92rlsgjjcYaay2kG6qrl4ppwaCe3yeUg
i/DGwzWi+8GU+qYBnrEx3g75HrOXKg5pAlZXswFD0KTQFVCKGCjZ7Bu/W8IsVOa0
ML2Ev4Nm3JZsZ4ueMpBVZbAPJM3zPVozSYijkIaVuVoQEXRxciGJRz5GgpA9wEWT
ujBAkz1ebojV5dydRG3n/snx+jTkSAEKMJHzDT3Ooft/MKrAywAjTWAOsowTAfqG
dzibdeWz612EZEuD5LtmepmEwwJCUd9vDpqMsS6rv+W9WSRlhEF5Hc0A5qvyNfDq
1CW++rPb86yOYI4e3tt/rt4a/8BWuCOvcdkOSC/oPLCfXhUVbT6tIVDvpzp/byZo
eJ92xv/pijfhdgFJtan09HOnkSl5JXzYva9tgJ6QtwdrPZgJBKG0k2ZDVFdqDpwy
zEo9TQaLuh5YCi1lYZQtgklfD4XNpIeB2aQSY7/OqzIK/qQsXA43p18cVB26xGtZ
ebbmy9BCZdMdRJRIJtshsPnx6qix9DUr0e23N4hElZaP82YmQ1zHzvOyaYF9NhzR
LCRHVwZAYwbF0GfqWnfeHxWV1J5Y2juZ8bd+m8d/MnEL7uhTycZEo2N8JmLsXday
i3GL+2ExC31qXVn+MjHUD0wT5sy8x83vrCZs2YlNvgfnwvtjOH/MOMqG7SWn7jf4
Aa6l0Z43NuMZUPWr0RhnFXUKF8owXDFtNsSF3G6WwpmnpjwcZAvFZVtXhhUkqs4X
thmOE2/4CfcH7jS+gf1BzdurL+GussiL2yh4jVIyMy2FFd6NRfB3BvpS8oVtlO78
yVL7yGJZl3yvKhM1ObeUCUGB35PvZsbbW88Vab2Puimple9ZFwDy1XNl6fzAbXUp
HiwoFP+b0loZJISTyLWXq/42FoltBmCEP/Cm5PcuhCT8/IcgYKAUSgtvBecMfLEI
b6Vqrt/fvKiMqRg000vv4de8c258lAkOb4d75a4iIg94x8e4dXp5IXhGH9FRyglT
jjDk0PIZ2IokQNWmdajd66VPHach9Y2ZsBGhpER2T+xKmfo+dmlJ/jcJkVn++f8B
010bymTdD9d7t75ro3tUuyiUIJvaSDS8XIFKKwMnpTTJisABobLfCYrBzs91WXjs
NzFWLs1opY+1b3fBHjGQXRlQRiEYMNa4VOpWKhyvENPoonCJ6mYkQLKgEWh+nP+J
jdbCxfDJYq9U+oLFwV6f4pLaz/C/qPzvx2A+LoPKS02YJ2LfTgUfcwTvqqb0ccFz
KFtVEX329Qvzs+tVz6tIhi3WvpipqnUJ6CiVD0t7BHbwlh9gBjLAW+dV8MSGaqZr
DUKcV/buZgKXMblPElevN0KKd8NtBid5ecQ0leKQscquWA36O9jBVWuJeITgRib8
ZeSglXXfDMRoO5Oxa6eEp1H+qcmfyMQpmpA8LBmhSMhAAjDz0IBKJtBnMN2eTt64
pqGEdCihQgjMFORrZiYB1tBwedTgSVO4XwCg1wOSRbpb2YRjAGSaQ/Cw9SNcwhsp
TpbM3KTldkTK8TFwMJMNeRfBZlG/J07FN6+s6pkXcIXJN+hO27gIjGYS8hr+zEdq
MSZcZRtPkLytMU34k6Ya1dh4wjmQoTBJDr0x1m/OdohRIJ0tewVYRNecYyP1DoSp
emo+7akISI1pprLT/5frqY0ZN7OmcQ5xZUBP5FBQ4MT60LIhTTybiUxyaDvHpgtJ
V+wF7jRCtZO0ypSu0kI17u+yDEYgqohFEa1gW0WB4YDT6qIleO9+pQlHBeafLM+v
Xv6IAYGUtRvzkVtt2jahxHCCvfW1wm1xAYNcMNfIkmEJPq+8UZPVJeD9+qvr4QNL
KdZBblVYcheJnaVq3/1QLN/dm+FBioWLbNdHQdHFvMGL8+lCcJVXNMvI953f/iaw
Upfm5n/lfo3/ZswmcYlHJ+3kHmDmcr9+4eXtiTuUgMg7aWWYIOCUnzvGcnUDmyej
NhSyqp81Qevdk0ug68peJzjSglg+oLAhfmmuxY83E6dfOMCHVEkB8ucyJCH2kymG
DzkLyPuhlSiDUNrAGvxGkztPN8D8FePuptIxc2tllpEVa0VR01IctSznf9MU76Jf
7loqPtXtCLn018p257n/tzaTkEvl/tiplQcUiJ6lIocdajN+kefYO5LhY6B0a8Ct
s58pB4W/HUDHSqcLUEOxTbD362VVrbD72ZCKDJu0xI8VvRjiUlV5ybSrt9ipNNly
N2BYQfrY2fB6rPJBFDqjbk6h6CkNqwAsz8pp6EUL1DjbFT/aiJZg7v4YVoENm2wv
T4oOryMRON234C2hV1r3Y35NM348gBG5Vq0mjwszZaHtemgHYrdUjKTald0KnyEL
CSvD9Ri93gpVJL1LRjneZbX22cFSkdJvvUGHohpVXJ2sHwMtC4wOH9XgGnQj7q6E
op+rmE/M6j7sqtq+F3en7etqLJo1kShmYJ1Y6rumdXHzwEPM/gjdjpYisFPfXU6P
neuGlsS0BJlL3DS+dF4Xs7AudOTA5GPpjdVtmg8I4vyJpvr/2Yct/f19VBKih28w
/t8K2GxVxFOOjjRx6iETp6hny7ZKqZw9EKaLpE0qV+muXlw7WvMYtmWdvBvH3NKT
bgIWRjyZaFAPoYIXhv7RET5/Q25y5/gE86NF+3B1wa5I/UwJDPIezlCw7dqj2Vxl
TDx/WybqrviiKaWrbSgtTtWiPNtzxhsQFiTFH9h+txjeKjFDaL1XhOPy5vgC47rX
N4z4XrUh9mv8lcJvqbx9h+79YHz09MPkxI1IExgL3YYL7dvaBdOfZdp/ovg/4YyV
4pq/YsON+HbhpRMOzn9RRZ8V9iUXTlYqjHUMTZeKC+mtzQjAd1dra82Kczn1BchG
Yypp0f5Po5ZMDOMOnVy8iKVxdyvXym7/KWXGb29RzaJuSOr6IH5oGPNLrjGGaqNp
BHbNl4+JAE8BfD2FPrxO0vs2rr+8WHPnl9r+x9KzO8cxXruaFLodvPV5RO8LVUmX
/mqohi4tMFb1yldDofBRFkRSwboxLhfBvDHgsx/d7p9ZdbYmA/IlRKgnU+DPoY4j
MCevdKV1UUj4m36KSQihEw1Da6CJP2fx+iuzShaQbVmv6TeAXKaZpSl1NsECa/eH
0K+LclO2Qd6TjktvIql3TMcxdssqMTkZQNqiLxN7JN6wjbBrJf2n2FF2DAPiK7fS
rphroLAaEPyPojA5Vz43+MD/VrOS7noHAwbtdOaXksXi7P31HC/G/yCBkiKuzCw/
8TFKexuYNr3OgG23wzJZAou19VJAtUVEEtY2RGQDqsohsYG/T/sMz8IFeTBjGd+N
gjKaZVAnskL4jDKbJuOY3eohnem6seMjyQtoAg7XLr7cjAeMhu0eBjDn6fnz+yci
sGKJOGi97JpRLe+JvevSwvrV8I+hFwOakySN3o0tCw1kPJymoK094jrrZq0nwCEl
z5YQNwMv9JezoRA8KQu2TLqTs2DMiDKiNGIXxmzIJm7XlQx5tDMfp3GMJoJ73tpb
Jc2EsisRnzX72TJlsfA66GvE01CfRhuYhCJzz8aq1LLd9nWKgmNJEBolRLDlmgVH
u1qK5wWaKGkZqKOQ5hoIlgXvhWaTwYfrIAXvmk1dhSmm9N/lwXMTNrCfv3oYiGDi
fRQpFsOkgWq5zhVt15MceRRgy3TElHCGBa681juxJK6gG7Ro5gcqj29FTXwEEKZi
He477sl/tILznzMgIVEZhryjBp+9MgJ2Wn6bstaO2Djvx8qhv/0ovoCWnNrZo+54
aSyzqsHE1BD/RnZqH/e7KfEYc0Djro4zQYKUhgfz3sukgT7tac/L7OP4CdWsICzi
+A793xB7mA7A7WF5k359W860LQ7n5hCTG1pkrwnIF1Xb2vzs3RgwCeqmV9m5FFHu
kCKSIr2GTkGfIJyWwfMulqRwGlD2Y8Xs/H8rEdR+1+3i3U0NbY9xjxM1ob75Hxtb
czqzojWOJHn4px9cyT7J0lWERboXDpSUeVfMWQ+k6W4lo8utu+p+aQOVT8PDDmPh
felA8cq+lxmpo8CbMjz5z7Q4NvCB5u8x0YR/bRslKXMET5TWU/uq2pOdlkJkopJV
W/x0i1BQ7oZrxc1Usy35b/RB76EVLuD9hDX37Xhx4dQkNQCCjFCzO2RnIHa8VK1e
ZJteS1Y9M/R/LB+ZPJOr2//N6/NbrWtI1WsEnrBBL2uAjl7q44ycw+ntJOTrWozn
KpthWrNN73DzDnhZrn2o0wyaSSH91R7JJDcOkfg3ekLVTKTLPcDMLZJM33NjsOrT
82q9qiv3eTVzHjP5oDBLy7xi2BSZQrw8YErnBn1ao7K/MnyekpSqYTZhPHfBb4hI
mJNDj8wNCFxWEAvQ+5WK/GSbldJJTm9sRWy0b7WyY+TwiYxlZZGviJyuYOxAbebh
WS/8Pqvd7It0x4+mMtEp0mXu/nrkX+aaiLPm9xfXs1EyrBpTaiaCzcZEB1/w0VuA
OMEEiAmqNeNJFhc0BP73H+2wu6WlsTjcgOHxtfPzhD3VLHARsxFwU1Zwc80hgTnP
rrxff1hjEaPTUSAKy8a5tsckMM1jRTMe2qKRx6sVAhJ2Al9qzd0ACWJUBjBTCEVu
Lwlsu5d7NOajsQvwhOVdJ9Xxxo5o4bhSgUsp+8bW2BXCHrbZL70PdNi6jzkFiIaX
0jSjb/Da/5DaN9rIiw+q54UEbY+wjpm546N3llCWKEowxPbqhqmxT3LH9Loq7M5j
SrK5ZywuCQ875OjZxxL7fhbwRVZl3Equ9JuyvutPaprhLe0gngcJhrtLVoaIsGjb
cLoVCx7FioQGOm+bCHE1ahzUI/1zXkyJwBPBKZm9GzgiGx4dGpt4ZXtMEhXe5RIO
P5zjs387fpovct8YRzwlYZfxKsxmVf9mUAZ8Q3HI5pGtc7hyW5gpdLta0sVr+tYs
0u9+jKPZzNbjnUH66MyUw2jYyTfFw75rx4ql+XEvWJQ0XhTSejHIxC82s9DxjFKQ
ZLFwtT9MHTZvI1y+WgioAfXaYz9N+CpqeazIb1SNeMJLe9fZtvT8W6K3pAV3Yx+y
nAupx0pb+5J8tvh+/hzY1DhxY9z3CB4cREk8mx52tGOFSOGgznLfAm4MMO3JE1Cp
va8YHSdahiKmtg5vcxP3j8Fqjah4MmG4UpU3iQzcLsQobRG7fLNKCsGonhDpIPUM
3cRZtTs6CBHtcZ12naNa6i3/+XHp//g0nIzTzMURazFTR0lEqFb5XkJHzA+ad7FR
bDU+RECdxALq3htYKjNRkahAM+fCBWCy6Wn1XxI4jTGUTV2wU8IcRStJnlttDmGz
/gA9HZgLsY4J5LXI9y9nHOmkVhwIZsnpYdQSiTxgv56FZulW/+OCP7w7Ee04y/Fu
YTawsgelQsegvKWEOOVD6SOajw/x25R1Q7dxxQE2BOcAFLZ/VG0zmnYsCJ7bdnx6
VJ6uxoagZytW/4FNqd5kYtV8rz+f4/j+d5H1IBGp9hQLGPnMdupAdsfv+eCC0Eiu
/hbGR+BxLY+qOIHKXPI+WwY2tC7h+Bcd8dDxS+7CHVIPzeAQVHt+ZRwPYpq/2XNU
482IppJGow5jJ5V9D4/EJoYVgRsJ27YvPqod4r2rK2FzjeuIvk0huRGa5UXUw8Ms
NTKnxBRKi9pV292q+EHqIF3vWGEbcIMXOMPrNdmvZxCDIK2btxCV9qBBzhjAPn22
or1VbEhREVv9FkiyinrgKY/FGjbAs4eailghgRDf+Fbb0vEJJk9b1p+TucSOr8p+
B+d5VBMXwbfzreX2UCLXM2Clx6QekhcZlkXHCL08jCzccuQQsC+NtJN7WgSqUYcu
09tWTcltY6/AiLlfhk27B1zJB3NZo6W0zKYNZL3b0KnSForU5GDJMzfJl5nqVDxR
jkPeOLHxQcI7Qk4xhiP7nvTXkOJeNNME64sd8MyO9yGwN17OTxlyNxGbYUN5APwc
ou3sfezeW+dDKDOT/JWzR1HPEOd3aO4fCZCSUX/zdhKFxdE2f2Ef1yR/R47Fx40c
38hXLN+HFHkbLgQJJ76Ttu64o2jrsENNED8O81C/Jjz9bHGRmkKlyvWc2Ng73Lpt
Icf/t/9Iyqi6kHSJuv0vJSzAuAKOidwhubaCg2wkHX9d2gXKCuTLEKh2G96DkAPS
dx1PifoYkch9+9bwPPDJiUqgMAkY/m+cBs7fYy52dz5zaGHw90FryTUEEVn6MN8T
fnqbnrpmhYYwTL2O9Xj+AvIsQKzR3E1Ed2tUBwy1g0/1h3rmmm6eL9yi4YdrG0i3
gOXS2ouz44dv3XoewszupM32fIPj3imP7aguN3OrnkO3lmypOD/AIlUwL1tnV7g5
e5hMZPXwHEosKhithG8gmSbkMWzTgYOWej2Ls9i71fg3ZskpwcDTJMEBPoS9/Lfm
3+qiVdzy5Ih/EFzDIjmeLFq3ov0igswxEnTmlWWDTVzJ/Mca0W5a6hVsSZGiwoeN
lLTl/sMBqZzXWOGBaNbl6ssLKXA7EqKpa2Hs3Q6ERjU8ZIbDTKxVaop8aqdfk/FP
OEwGSvEBoooXjyeP0uiOIZ/akd1+7B4iKomQx5gwFYACm2QXC1f3OknNxLaOSeKr
iIDELj3gt23VJP8xXXwG6weWd0BJkKnJJcE2WyrCGOuTetWMI5FO/fJZ0XhbogGH
cTt054AGk2SdlLQpO3N8857RtpJIEI/g0TL1s7ROdZHPsUbZNggp3ChZWwxaTrrX
f4sH6ibYTczyhK0pHv9MI7NecvGijy3qZfR7lc8TrernQSv1bXgJZ/UOhyYRQym/
efjX/PFKgaoPMd4xJh2MAczKhRxlQ5BeWNIb9RVxMPyeL708R/0KnNCqJd35jmkl
B0KmqFRgqkcu3jOygEFbwLiEOJk3hO8pNrV6tD1h2ctU2gr8hfHvo3TwhTpMuu4T
INYP/bfhkLBK5kbFZUnqr84XxSDUcLL7gpuxgCBntcs7RFsXH6lk1kQ7sgKLCDid
tL6Pl4ImrJpNt+yP2fAiJ6O2zk5VyDYeCy1JLtl/CI0TCvif6Ca3hZh88atTQohh
3WswnBArbTd/CmpZyvh+9t7MRhtp04WQ1Ra8Antze+HouIFHQt5fEayqFzPHQA8q
NnUQnzfLdWMoaHWtMrq2eF9gGrDDWLUvj9/6QUGGy/2T02RCAeT4JndYmFammArJ
og8gOuMiR7xTXxCrS4E5Q8Wq8RPBvNWaGJQlzky/y+XI1xcA9zGUy6QNkvo347o5
KQL/Gwa9D2D1QjdKJJhdGk5IuDiVI7co7lsqsj8l1VPXpN5sAMYgtmH+lTH0N28H
7YCTPuiLcWLEbeKYv9oXHoKZAe6kWjklWiyTZPyeOoO89wMKCHI3gmZRmxqzha82
VIhABSmCIPZDRSoHR6hMDomywOl/zw37p3O/SrNPPb5ut8ztlZrTJeDj+QmzJjAB
MPohLXaTwjWVdHnX3onK24uv+iKJCsc38BaX359Zij4sYcum7iNyVlEijZb3nu+I
X7HGva0ZHm6/nh7ndbr2Bwa5gVxcpJB8I8MlmfqAQxHlhJ2j1oMyObd7l1Io/6zu
t30l0t3DaU1RAwqr60LaLXmP1WOL9jh70ksjQgwvfxebSsKvwRSGa8FwDmCkfwkZ
CQSl8cuhWbqlhoZMSdtt2p3cAjLYTJhApn7AK2qkn6pXU0/zgFFTyHABvAwE8ZUz
edp/ipzNryV7GoLdNE2+Y0syYHsO/EupMCVUawXTn3WKPs9qhTQiU41J/tV/2uRb
bM7Lk3UQV76qOCe1IoBM88QBG0K7EXC07EWfYtfBPQSGfXjaljwbSUo5g3wUxm/r
OVfuRmTv1QtEKKgGn7F0vpTypg57is4AX3R3pINmQBOrgCRj5SQqYNo7tZOYFVHE
OMk6SyC1+BpjKMPLDL3txNe7BRENarD4UHSGZr0PZGTMa/PKWyHDtNNu3cILKcfV
HsEr1tEPcKoeua6dB1QkqNfhm3rPTUCz0wde3GnlesCjeuGpra21J1K1LE/ZUtRe
sVH6pv9Nk/5vgj8pGI9LrzRYznSLdTcrM+DdMypz4aNgmOWrLGcxikc1grY7EQ6g
Q5cmDkmNJnPcmFDO6v+CytoIBbgjogxFRQJW5Pr9yNOYkqnS42GYrXkCwUfvOBQG
RMTAZS7wH5hsV5gbPEeOG0TZKZZtj0dKbkvA/dV6ksOvs/3o1w+IBl3Lwahve4DI
5o7GxkYoouJJznOLDsyCw0mCITDKwwBfu0pLGmmXNpXLCSb8usyHzhjA+bwaOQs/
gI+NuDLKm7p81+l9PCnl4vh1+/J5PDZnDPyTAYLgzWlFhn7KNP74ITWp2983TdU1
cYqJGrTu23MfUOylwNMaXvQCgzJ8Mqd9i/z0bXdfU4abUr7kIW2yxded8YAncLEg
/hbhIdrD1zrnpaXA34OFHgsNZZI5I54glHmy48i7q1dJ0sgSGtr1FZNBubE7+ueo
acvTiXC8Yg6KrjnN6c2fTHoNfgrF8W84NMnTyCpTlMBMYxQZ2JZrUiKZCACUBbSJ
57wewvufd9wq4W+ztiO46R8R1ilARqCIfXfhxWR4nro2FPBEI2X+AlsRWAFJEpGY
DbmbQkadFOVRic6o/Y1BCXD91gSmRBiMMuqFQSWi3KKUsERPx4DD2DZ5Li2m7cVx
Kcr9NFMFyPtdwZIPlJq6bsamM2UGwInemU9u27M1uKbPNhBC451qplpHhBkaF07O
mWKaeQpVbNrQw3GYQ6TaJ5iN3OnAYqjoGJfeQ6oBvFPQh3Si/Adv4AzJWYSUTnxC
cvvBgSdTaJpywyPAR7AlX6lBRDeLS1lv6j5JdYPLEx1golse3wQVfjMxaO1AEGF/
RIpcTgxvaQWDuebC9lI40bg2/Uj8FqYg4yxvzgj1YHJhcevzkS6pghl7n6xIVN7w
BwdpHnn2NIL70gkyD/xcxesv8d9fmduRmZjPbjgguyIwAmsHHK7SuAiCP6wcze2S
rzzPqWHvM1SPJWl41ZHd5y15xlwWbofidFX/rFf1ofUculfSGVFC/mprzB3KtwgM
QuDEpmXDTcZv5u2fht0IW7HMcteek5e2uiwxlxOjI4aoBQoH8Y77qws9gxRZOfQQ
HDXuWLfD7U9idgyZbzdxqWplJguGarAgchC/FSFJigk0Jplmdg2wUMsQn2AFMI9s
4brsL068ZmBllbzv0sw7k8hVSUICTQuW/HaaCqa70nQPbG+1+L0x6DSEqNvS70qX
ADpaNvZvZa7XLFvzYJ5NZWQJwvfBl8zvK3RWYzudAn2WG2XoBCINrQWUXoVXgnwR
7HVCvzvDhF2O9pY/j0TbubkLjdqb8dObp/j68+bPLHNxIeaWeL0iAzwFlHXl1qZf
d3DTgJ1F41sL1tEPT0nue9N28keLMgcX/Hyt6vxFZ59P8KDThIDEMlfYUCjsTUBB
aBgNuniACYL03629IP3yvAYOGFLLR2GORsDd2ZVV+k9O7OHMKZdp7ysfEXMiDzUS
CAKdQgQgkmd9H3NYMkBxkYzwY4w0f3KNlS/dKiVlAdUMqYynABV4Py1n11aeWrWJ
bLfcePXl+sAqU7VCCsrodtT8tcO/h5gDHnPMZ5BXV1n8Y0uvZJf7XOmev98wKuKr
JcErs+TkIPJlUDRMDQqwf4iVRiJSTYMbLFmkOY4OUhshFQKIegisRMsS3A5w4MvJ
THubYIgzIl5ETj7sDntWy1ds4OwrTrKmzSU08aUGmyOObTvMEU+uaPSVaKBx7g7p
stObxG5yENvcT6cjsB9p+J2OV6eQeE85JGSgby5tUoNdlDWIkolRtak5QVIhQyCX
7Zwp53LwgULRCxefPax1w+XAEsi3sJ5FUfxmohQlzyGuVDDM15oey9+WC9freHd+
gEmg/u2PuvlH8g00V8EcBgfcbsfu3fHiv24QEUyWiXIMMGbXfqjYhAcSGwPhfm8P
0CYv8emaRzJm/K1qBgy8J84e7X+cjAcs6xOVbtQc19+ynTFIp8xNkF3rTIZPSgUH
S08fCX4pRFJOoM4wTVDjp39yUkrLU80KLcT9OL43/gDppcTJMUHi+4mxXyD+Fdw6
pEBXCzTNmraJPtJiUGwOGvxIXpT2vE0X/rlAiuUyHzutZtkf5lWI7e15Tg8YbpDg
WWMhXCvZgEyx7HRQEFJYglLc+6QHzTzSdjs1I7OlIYq2w/eIU6luQO2lTvC8S+HC
JRcKSGiVo9+tvoEVCUEvVm2ZsL8/KigrknH3BJ1DjxpvpGG+heujczsTLPgDSL8o
HZsPxD9FzK1HqFyDjQ/MofPn3GE5BFaqzrW0YutkON19Dcv3gmvm5CevXZX4iuEw
lEbsMKt6xlUtRMwRfx8HQSVxROri6iUN/vsUwcSpr08TpqMje8iiCxD/yaxymhBP
iqksEjRiKEfyWAHqv6Eq3FbE5wrC5pQXgaYR2+z5AyU7RJ1bl+BSs+7GSxco1Yib
UyB+n9Xlzw0BcpTuzBBeVpwukEizyL9MDY1zzO4hcG5DbtO2EO8TWu2C5HlOswMP
Fo1YKQm3CxR2qEpwixAbSKfHdQ3kOnxbIDKcAw7xcVAoxWw/0+O1temSkS/DhYFU
8Gw7PuYtQojklrcFrDRADP77rLqE1sfoMY1gpC57dD74CnJg1IDKzZ22b9nb+Qrj
g9qlDxDqE4hE3chAhYqWhL1twUytmKZUl7ZIeeeS2rcy6AHsudu3nLlgXTmZYuZy
2OZLLima7bhzOYPJz6+x0pBnMbbZIOcyCEBvXK2PA4lmdY70/QFy7rJk5dOHH8jO
GTT8Jd9Jf7UBKJe4GBCsupqCt2OjtRTr+UX2RXZ12SvYXRRoRZYowc8LLx4euiwr
wmUWZsX7z2EI7B9l2TUhmjAwfTNh4gdTveyHFnxTsqjh5SSCk1PXWxgiePN2UHe+
O4WIf1AQtu4jqket5yo67v8za9zVkStfUb1h4T4s6rVUUbdjpV3y930ejHzjC+MX
ZMP8ogYSLic6SQrn3kOI/Oy1i41usZoakda9q5nROkiyMu/v4VaTCtYffvQDD+dA
rZNa6kdzqIg5vu0O8sYbzrO6D8nHJgSUJH3pwtA5eCd1zCWWAYTwiUR5rZb+auiM
r0POEvatuJCh+UTDZcASibBwPTxaEB52ooh7AUZWVJ07raNpgzyrzB8ik9vXBiGA
ancjmJe8YAMUqW5Oi0Nlvw00SC9PY5OJBsFI7dxaT4ttNR6JVoCCNp5MM6Bgwkbk
PL+RQM8tuA2gTfBtC+r3joldJk+6Kbd60IkRqyIe5Iych+2d8DzoSCJXHpXXO4ly
JEA9BzvuCDovz+7j7p5smSiWDuqBiaSkrTkHYiwk20RpfV12UQGnwPRYRTUMhLYe
Cae+uhkKU2LJsUN2yKW3sIUN9mYhjbfbNWaVYPl7IFB2Dhjtnpvae5kCrMuGmgn1
KS1C87gYAtBUISu38F6aGCY1ayBGt5/VLVtHdD93YVVUqT+Eyagf3Z4t1IV/hmHE
WResV0aHT6q5yL1YIqgQBc/KPa/u3HotXTX8uC038FkgM9yIM7NGZYN3L5E0Wdar
Hz6RIZE5xt19f3z32CrtgMyvkhip1hYe9JlbiLPeHdkTVnB3XOOEw58U+FP04rcq
GHrtS64HnP+mtEyAa3HY1y5ujkzo9T18Ah7avo6Ite3qiw330yF9LFNmMHhzPPmd
TZojnbCcVvG1xZ9rZg/qmv/LQo4ZbPPqqWIFRFAmAfaHkveqk1dzFVgCTJxSMUze
quZgqhfgWa8O7rYNuNERlqQGHv0bn33qXQigAS1hI03h0SE0S0qN/8cEk5hQt4Z8
mTfGEtiO2/T6b6P/gR6ssyUA6qPaqWnaw3D28NG+r7frZ+0JqmVmdGk7eguJxrdY
IXY+im+/Rejw8fQaGcjvyaqLW4J1gE6rQMTtLb611pYC5KG8glY4YJw/oY1KQcGx
s9WS7bxG9sk5a18slsasy+o+fRqCflG0u1rNBD3PU/da2zKh9pdWSC4dYKSGB420
vEKvhIBI0geMRLDDiHUV7x7QmBlSRecDEmJ+h0ojjMdQwkXsN02Axo4hxGCw6Go9
udbOAtHh1Ncn8WQOzal419bspe/dILsxca2oW5S2GDr7a+lEEKSm4XXNQsDBQCnG
ovlcRotbCJPBLk1RmN2rNkPJR03mVxtyGzi++T+OhKZImHNVwCLuVhMVkzOb3441
g/4YUEigrrZcxSOp43DOJ4VmPVHPEjEflYfDI3rOs7in+TjhCiAW5u+DqdG0N5wB
QgvMrDgKXgsNC4mtJH8gWR0KMjyYZ12Gewu2h5Qj+93LqWtwvY5amk8dez0lJwe7
NntLn3GHYvDtD/ldE1ZzCMgeYakfiVomHKzAHCUDoeLXREWdU4rxeOGotwRsZPYE
MdxxcaXePCwWT7ZPzkz9jhNEJiL+Lsod+KWq0CorkRRL0cXAbYTdFJ3+MGOLA5HD
oHipYontOAxXifv7P6RMjQQnDYdFLhtPpQhu5/rZ56uNszZW20SXxusSZWk20f0O
o5k/K2AfY95SEACce3sgiTd/jULxxVaiu/ECerS3Nkv4EPMeWDCr82xYHTgHnHKs
oWd7MCgzbh8BF0fXzDIyWdTOOefIe4hHfb/s39uEY5ZIvh5ZBhhpkuENeOL4P2hb
/Ug17h2mx0PTsofzv55Iv/3On45Etd+lIgYYt5H01Q25IYXUSBx9A6XV7vSjj41k
fvp07etmHpX4GuJNYz0Ad+Nwfb5i/1Kfmn5mGOWxPt7GLAmZCOQUB2/tPicWLGms
NZPzgiuwOsrFU5I54sz26yeA/fh7SDFbFOKrmvZHJplbG3cbAfu35qRXRBi8lPi9
rZN8izdGmxvrfdK0TIF4SwP09gTmmrkU1PQnYG/fP0doYMQHX8O/Ra9FSXXOCV5B
WFQETmaztteodJPnGwQoRbo/B1pyF7plMupZsjAbuHV0ueNeYJ7ejM6dGUE5mJv6
Cicitp2POnz63GXNRkQA++TNQkwVNylBGY6N2UTnCFC9uFrA0t/JzRew/HePukWj
aBpgZKvsuHmsSPjJFWnpd+xbNgtW9t/N3UUkA8AezX5GcxsbsKBlalzaOSXWjtYF
bkbIqH6bZJewVurdKKxxmceRrKV0dcUQN3cD6GDcaIarYhNhIuE3pjagt/mIWwZY
JW1ii+06UyuZonc6zjcgSFRbRWlBDkQze4/6P7yx9RfPsFVLkm+PhWaWX2WJLkWn
MtqVisarKg9TJQgwD+YJTvdgqv6yovRt05tRfEaGayGUo07i11GSVCKSsN89WKtL
0tYWw8xUyGxGSEtjE+OadXFx/kIuKvjdge6rrgg5OI4T0sl2v/0Y9Ko7PoiaJrU2
AMLWfHyxd1NiBUND4MPqZkZJfKfSQJx0swdURAgd7yBrdcswVRlOCc21c15AG0uJ
xq1ECP6tPbL2dJwRM+aRqpVwREPmDTTLvtdQYnx11M8+ZH8jFPqb0WftOSRsK+ol
KGZu5yDxKdg/oy4CYum1DPTFbXwPxA4nSDDsNUN16KF0l8cHrCAD9p6OcrWYcCGL
SPxUx5liX5K14333wK2KKw1eQmqJl24Uyu9syEvjKkQlDinUQrIleRokpPfO40QO
RpoF+yM96e4tNP0uOAIfPmCZgfs7zxsVB+Bk2+jRosDIcSrsHwdZDeRJZj0HZuIT
qaB2ii0V9IUg0YFeR+/xjn4o27KECte21UphWDP4p5AtAWKWTFeiLDvttORpU3Vd
gtTwad5O63C8JKBD2w2ibeolrRv05pv1z8K8N9PIuq4hb4XVh4nvCZ/bh1uov+/I
lEfKnPQSAS6Vn6hCgfhCnQ4fn4/u6/yBTllf+XDfYv+/9hYulJP8isyBYgoEMpbP
9Iiou8FwKAxMQ8jW1RY7dLAw15qq4hqRz89TpVfJ8fBRFg1CqLfpuGjxbu6qyDQw
rgkajdHaQipDqBd/PkFPL4iB27PwQULgYtjWC/yzpOrvrWKIYaxKTYUB3FcuRTqR
/zo9KlSDhlq4WKsJrZHE8r+OkP1pZfljmxv8+kWGgO5rH6NGEJcsU1Yq2jePxoqK
eqwTPGzy+HI1fxWQ627TFnkOQkP9TTGvDPHxhyyUreLvd8zvM/jEE99cTZmetl/w
BLctp21cN3p4QLGNS22M480O5nNiep+0zNhpWCweK3ibi69SR+YhG4sJs+nvWdIZ
uGrv7cQ5UktVX5yH7pp7F+pu1E0Ye8loKa0+wWi9/v2K5P4fKG9aNJtkqev0/FGK
HvVKjUUJq7h+WdzRu3iIwSyxPXMOiIpAu9XSKJ/6DAEumOP6HiHgML+EKCJAA7qD
KTfc+sUQRH8GtJowtVjy96roX81J8YyCiW1QYchuh4QAXlyTAkK2D0v25GPYVIwz
0WMCkxOAe07E4pwvpu+rJ4rUCeEszTSVsPMIH0SjbKCEHAfsOn0yBZsCZEKquNza
dw/b+DuObMwlH214L6GLnkg0kclblXm9PorOrlLWv/7nJ0tuiGfnCcobG4hhz4tI
l0lD4SE0JwlLWveDuQOFByw5HPXMhLe5UJj1L+/VC0/am1j13Gjv7bhy5kzCsWds
XgHF0lAbX6NmYbA8K+s5RW6J5fLcxmgnT+5pARwL5y9yyltQ6QcIfglf+VDcHMih
3WCLeXJP0U1ulwsma4YwLRANSmoQQRLjoLM9sDK1PsBQJfhvjeQmY52EWh1ZZRbw
VOdzTAAVCmW0Sy0MYQ8IlCvudzXsIeZkM2SUCDPOulbnj9LQQBbQqK458E1XJ18L
xWnK5uHLZsgk990kDMAbrGQMKmkG1z1lWobmMb+cFUVcoK8PeaiU1Rrat9Bx1UNB
povDjctxR2iE59EYmdJ72tmI6EVaMRvdAv9L2keuP5mLjCyuTEA1Txf8pvdaTNLj
Ck34cqQ6E7T991TCjHlXG5m+ZYkugja9GEFg6LJQ0eEfsS70MEZe7JB+fbVgr6K1
LdEe+9sHuwhALfQ2W9tAmUJR57+lnrH9Vf13z0kEeqF5etjZx3/WsgCcKMWOku1W
36XD6Nny7uXmPNPqOsOu5+BXUGrof3T1lpItGo21n83OL7HMvcHD8tVjGMNvgYFF
W2TYn4Gl+3sEE5izR/xLbqV04XOGWBxXk8U/dN9XdyaEwxkttka9APU5TpGf33j6
sdUseS3XZR+seVWEWklBvxO8V+kEpC/eX/srdMtMlu6raGGjOx9oDd2htRUAi4SU
GBLxlzUpPpfjKeper0RsJCccOz4bzH8ztr9xagH6C+1anA4Sq94EHCMEYqEtfkXz
v4mK4D6n7sEmseDVhr8zlsE3bF+P/c3IgutQN/u8uKCNuMyYoT0H9FKC1dBUmwtY
or+vVIUMZqj/qR/E+tLc5T0E/SogQk5KXtfjmvtyh9iJvZb9KLAHknJBtS0OGJsG
51XL2qxMWg9V1GXE8lfjC45D0Cima9zy6WMrh1gU2MNc3TskUZOPTuBbq/esgQGj
Dwaf+lg9u+D2gvrHKOJVhVZ4hgOQKto0B966yNd2OP0POZKHTuNJsYqV5Fq/HPRc
orgo+w/O4IyOng9HGV8X75cA7UuHK97BGGX0ALAvr38wYB5ncKsrhQJSGH/d6dtR
cm04pwtIQg9YyjGteKVlrPyqCU9fCzjmknYkC8P9q3qnnOGovcsi56uAn3J9uKAG
I3HcYSnYNnbBTo8bSOG/n4CHsTOVrEjwJ0ZKZRVPPsm1/2PnYO+bihLxIKwmnEr6
mbM6cSuqvwTmX/oVqxR9fwcSh0a+5HWM37bkCdrF2IPQFpaxYUQDODp0jGvFAC/J
WSDHhjgiSq/y7ZEVmXpY4Iw5Nq6rjGIrHnBIKzMR1JN8u7ESwV1dMlC87BjCZEfw
k+nBCYjvMMOA2ZaWBPb5df2s6LNgXlB03/5iP/AqU7agPFHC5Iq2boLJQqvA+dhi
rNgyyJCDFfeQ5E6rxohVch9+NLjCABdj6dGM89H2JvYD8KZ5vRGTGLbqtFf67HLM
msbDcE8VCPL09Emzfra/y/r50oB+0Ygi8SLRFgaU6cOXcXo6AW8wMLiaBnR7DjHY
8avasjpyb1RCq0Xm3WBKi5nUm70MzzaEE1eP5WJpLRGt4zhdf9Ol1F/mLyPGuk3c
MkLiyAlpTLk/Pa/U5zu1VarGo/icWub964Aa8mc6sbwD7+dwQIZPMxDk1seM6IwA
CPOjrdQVtHaRcfKguPRDRk8oxeFHt9sIHlUZxSiZW6Yqs/YmkIQ0BBn5JXMpXrqG
aOeiQvOFq4UROkznqT28srl4APTcqpA7qNEXCkMCNCUTYs5k1iDfQvIgrxr023YT
jYRzEu7WcZwPQVY17vLqQ7HD5bA/2nlveUGsWFHSlvBDdjYwQX/hmFrqGV/vcv9X
1ABxe7nvfvlkLGKvROU3g6zVpwo2UrgF1YkPPEA2fuIcSjRCT5++omrRPsuWNCcQ
8qHtD6EKzhR4ipHKC+jIQ4cIeUUyimoLCygKR94iL0D3VvcJsbNbkZCtgN7bkFSW
gXkyT0G3c6qanfGk2DyWevCBY6LgHiwz0HUFNygMBFEm9h5pJ6Vj5HdAN+u3b24f
0DCEzizfoNXsrWViZ+KI9fE0wk7bn35hNOxKUlc4Y2zYpPC26r80LINoijv4mZLa
55tiYGUzhJvz0bpkL1/TPpO2h3YuZNsL2hgQIun67HD3Y6EnGsqyP/fV0ObOj9vX
rpvdGzZXjgkvx/BzD9FCHqf7NpN2gIhev2hLjDs1dByScRThdh1u3dXgYM5lQKna
c6ls+s1KRcbrpqLQ8lpZDp2BEUxckuUKCPNQG/JyZueBPuKzkQh9ll5qc+Ee4sHr
JVyoIAXGfWymXs5ZD5PTCnsBfHStJX4coQhYktCEKwsItruRUvI19iyHHmxfdFqD
6gcdXs+OCqdDDRzedjgdfMlBIDa/AtL1yKjsWPw+byzuX5sMe6ul3gj+mfjnrfq5
VUqqQwDY+bfwX5EtgaLBYYhsk6k6vzHud5OaSl12MnvQ8aiZ8RuCZQz/ze1NNmnK
0+9hyT9jEgrZuyQ1hcJI6d6j/WidjOwMbc7jVaxt5Wz8gsC9X5suvtrX/uzV2B5E
RlbDpUv9RVEcTe28kmEs5xTeluHXrp+6Pc9ERWeJJUo0PeEtsVinHBn9aW66K00j
XFvHwTHtt4Hmi/q9zpEaHP+OLRHoUujbgwejZgZ5el4WlQYdaIUZ8qNtilPLbjSd
vMypzIQXj0bh+TBm1Gr7oa3z8vraYJ/zAz3F2VsfjWZkpVk66lKf7eC9ZtkDlv5/
dLTT/tM8khAjU0eB1P+o5n4ILoZib57kzJZ2aDyDC/Extyieq7UqRsxxeT3Wugq+
5sgdY8P7YGB9mIkoq/BCk25BpA+Y7vkPPn0HFPcqqJQRX4T2HQolPSKTVl9ypsWn
Ob/nnZtKkMUxsLCdghIEPU9w23suWrWYLpboktUET1s5UZcDva6E5SM5jaoRr/aJ
iyPLIVsD7Vf1RaCwGAcdkSF62DW7mvdbseOuXyBRGTswZ5mi9yd7PtH7+o5CbwfZ
m6s93OCDKR2k+TG9JnkMSz2fktm9sKCkVDotgiun+5kG1iZ7gXQiQh1dIeNQJ1ps
OnNIj7gDZomHf6aI5VAPCurqgptIxufT35R1nCMBxOLPUREcKkBOCbgk3NMVTpIU
wXxX2Y/n/zpWZthoQO64DojCltpkoIAAsgF6SNCpm8jRoUFsf+D0DhQ8riotNUqJ
DTEiWJlMOJ2+X02HjbR5uATB6mCwk5K6fsrdU44Zz1CAKgQyparbQ2dzbrQ3CMUL
JRqOc+I5Wzw/2rB4FSwFly+OH+A1guu8gvIfCBxt0Fm9sc0I5rJ/hljIbboikaOq
qGpqLPnL78BuytQGg2sxd4pciOSdmnFFhyOb8uNmC9qTx5n3fbw+zfjLQAJBBHus
kNuhm0q2drt3pbj+A59KlhN07jkhiiQ2Z0lWjCFDcC1nsOsaE/auAF17lGdokLbZ
IVGdkukS4IOa3up83+5DMVjfFwptnLOmn+SKGEked0AHze/x7ZbiKqIrUdnD3p7t
SoUZkyvL42JwDZ5w1VMcPl9k0lqvvgwKQTBXMKwR1lKeMf9rrfKEGJWquwFelh8F
G2nI7hUnZJzJlMf12+x3YPZZAS+AHRDAdPmPqi4UHU9Tdr3pGkAEi3UhaZbu4pxL
QTmljfCpHmQ2WmH31uOZxz8dHqWcCvdU78SxoOoiv2GSVra0Spw2oxtBo6akVgLj
64BnW/NhDcdNhptDrTliEoyZ/6BGgdc5QdmmrFJEgcRB0/mohTMGrImyV9FUeouU
DEkPSoSVKNTlqbsu8FT4OZLRW/ATb+aTjfv5zC49IrDLVC7dewRtcTraDC5zwYm6
478Ra2d4ZmShCfg7Az18AIybnUena3kxxpHOwqORZRWap3+ElEqUEw3fr17tRzbj
xaB1jgWFiz4Sq2vAs/s7SO2IqkqC71RQyxlN7yMuZi3DyHiBw8s/ULbTrNLKtLk4
32IKkpF/HoPMBYds0bjDJ1XoK77EJz3CExlss5/y/acjvNWBD28sWt0liMuBFFNX
TIgk5KpznxDS6QZH0JXv+4+edCxTh0uAEsWRy6uAJlD4QgN2Cmn3W8pEZBh0v9R/
oiWU2FQMSiSRxdTb7nwfdECo/yogmx+/A5iUsKU6JerOFw5SWXDy9CQXEgjPE8wG
KlqyfmWIB6qYKNXTPkbzQmG/j1o9W5e9bSgoQQ+DZPOtwmEau50gDOm+RsDJJyOz
9CF8nGK98CGSjV+l/krtZGn89+QDumG/Y9QzFTlXou4pv+RcGGAtiQYrLr++1pxK
mFTauj2klM94Kgi3jy3vP6rftJ9RXxZ2/6NRnBGGGVByMo8FpyZC1rd3+PwYOkpo
m9m5iimK4kkwM/ed+7YI/zhDKD2azkv2TLEUmXnK3POePLHn9WJDCh37u3qbE6jP
vH5uMzqK+FdfPi6tlm9Z9wdDf25+yM5eThSsvMPmmceQtt1Of2X8gCiu3Ca0/zeH
iLmh9O/R9FCg1eJ9348Qk7C+97x6lavkSh5wqB4KkD0YkRz9Rh4dqUfH8hMLYZHF
6kAaoJswqM8s/W0ac6BxMTX0lV1A3cZ/BCkLZgm64mj7i6RM/CQLdMre0q7bE3gy
MvgyiDDt6ZzlvpOvVVWUxNeeJvIsQco0L+v850JXeLnld8ip/YQh2EptPm4DXHKf
JuyUCjpMG/UeEgH6VpPuJn225IES1heI5A2MbxxmpCFJPcgZzaacJFeMAlHJFrQB
5K+3CKeST7Rxb7SED5rvP4TkEo1kwDMPypoPsl/VgTc5qnHJ2T0t1TtUHZTp84qd
pJmjV5AyT1KBomnHWRz7+1OUSM0TRTg6GGPrkIwHjUGOdsCQBHB6pUyHJys0+Y03
hIKpE7J4tmWgM9+fkfz8uSob10sUum56gS6UT19MDqir94DcKohrjkspQ5qUakxr
CdZMM+kjL1BwgYTnAbjQYE7Agw3Hy3HaJ4ZvUhMfBYK1Tz4aR3uBZ+n31FlxCgbk
gzAehPEFxWKHrg8rdZ8Z6T5nE3YrWAE266UsE7RvzW5h2rqoBPCiKGCUGYlq3JBg
JbRb1GLlnHUTW4lTZCdbU0yu1vBAe4urGIUVX3J2N9haowVC6ctDWjvpK6d+BSc/
dnwbOpGqNj7lYNNbGlPDsKMOdGt1L8Xjy7206dykESvENpFXe0pT3P8BQuzJMkN6
AEhw58zA1HqNIEkJIgWzS0VaQt46ci85aS5k2KUbeXUpgNd3DILbmE0dyNDhrafF
LR4zRuYNg1kOWWuKn0UUVK6L73NdlhHdm4ushGCb7VWgNp7e7qleDsJJVfTbPPWL
v3K13YBWZnHzKrUgAgBIkjQZcLGWMxHPKxJZIqsNuByhv9UCznB3HnFmEY9rKn6o
7GOUtTFBFFcN5E+39r8SfjjCgHGVsOidlHsr6gd7g8UYqhV+SSOGCrkgYkoZAKyI
QBNP+uTeZAfGil77BIC9QL+NgM+nEDWPBai8H9yGPwMLibNIxnXVU/1594HyNwFJ
3z2bQOtkVycJQAsQNfr8WRxiu+nWHxmX0wqw1hYoUK6VcDFopxfw1hpX8fK8rP8a
eBBwQgLG+I7XkCF3XHQ6dK+s6Glpl/VCMwtDoK3NglEXGRKgDQPD99IOdAL+8b2P
CRmg8qcyPtgXthNHZz9exCwf9fC+zA0G5a+eaKz+z4qMAvCJmRZ/T+AkA9MYLjvh
JqWDBjdRIUDxNc5drBHbNynpu+cHuQ8Jw1RJBQE8Tl77bSfKceqGxH751rkXhZDg
Dp1sOcUs9sG5U/LKrbUCHLoSrgAvUrN5OXeWmdKB62mJrSuIb+3S1gbxakk4F8df
6bmfQLwjOrortmlLMgDIBd2/y9UlMwKmC4CGXdl3c6BHzt7eoBuf9ZCtHjEV3fQq
1goPZPWFo/mGHWNuK3mgncinGSTkiTd5i08dR+6LRNk/oB+/KIa1mu3RJ9f0mFXW
BEOKYIYopvTj8VFxU6skwD7WYkV4mCos27uzNIv9JYl6DR8FoIEbsV8QvyIjBMyn
/ey7pVxMvadpVgGF0KA2xZGTtWQI5wXcbersU4Wg7Potwy+YkkYwDgdwwDadMuMU
wY/7VeXwXv1/iDA/FbjfNK6VdCU1qFneyCJX5jpO3tyPYt1zzkJsxDaj+yFzAmR5
FxiTxxfxko31zO/yMJLwwZ3rP5fA4fLHkW9Qt+PIuywGfHByyrwjknuud+AleW1y
1OrvqD3jdEnuPJ+rRopjIPfKMsVXxYhoF1KKsZRf4FwKx4XZmoHqqG9OWdl0KNQ4
PDjIUSbMnXTP1kMT/Q5QAVNsEL8pE/23gLzQ1CwHjARev45hQxqBqhA8BrCJi20L
jOyzPSij5QRCepqdfbtBvDwuma7AhciWLeJUg45qhkcf5KeZaGnDA6EE8Z7q/jBY
lLeRPC38HRkDfVEpRhSrKWLVLyRsWKioNTeP8Mce9N/PwsoQjJ5n7IGYk3WkwaEY
SNx9ga8B2Qn5tMkwxJBhbHxC9eYu6yo4ezSMqtvv0whYDtpESbRxDuzo0cYdBEDI
QAKJtVH1YptF+1lMjnZYrlyBZ4e8TJCgj4spj0ETK5dxWrhaN/Rx2EDfRV9lUIFJ
74ULZoxs/CZJXmm+8CDalmGqu3w4HiLdHmcq7qFHtDSmCz+XW53gfseAWvawmd/y
J7MC9XY+bgO2TB6PA05aLEFHZMyWT8k1ayBglEydUy0WyHpsuWLWIsHdtvOwCkLR
w6u//Htcxy8rW2D/35gZk8pdggmFW4JVxuPGqS1bEWFdUM6EO2dsWNSnd4Ig78Zm
LesYH32BYDtTBV7+VBypb4paHCLxzKtTDEF1PKcvZjM0//ChHSkn9ej9ipPPpii6
/3eaPAegPK11UwqIVJUoLI/b3U0ArtQxRTwdhtdBb5Wugboue2uy3qY3/8WnJ4lL
GhAdlFkx1zPnJM89lDp2zCY1c2fu5rghl5ROEx7s7lnpOotwQJayA7V9ClCEiIGI
NG65nR7tAVcjwAtwogytfkbR4UngI7935iWFKZOTshx8LRwJiAHHPtsqMG2ay/Pd
oy+0/hhksA3i3XCF/6R6SMAVnndM1llKU+Cx/4CrxvDGFVjF3z2qzIC2bV52+QbW
g51eBN25a82haGm1jPMPevSOdzuSGPYcP62UyNzBkp/Bm0A7KYckMl0vTuc8Kg68
yGHMz6WK7AB12HKU2aGpxRhcXgjXOewIxvbA5UyxJ+738nj4uigrtd4qZr0VeVkZ
GfhpnNjRt2IbBo2QkVk4UiSq2mGuY+dpgwA2ZHUNbCF2vCZOIm/ni9yj+itRxHwn
bplhVRkqjo0X3eKPIUHQvSPa7i+8kFOEWGE+BK8KcGfgFR8dzsAIuvLEFyfHlJ9u
NokJgVsO2aB3BYtTBmgtXjFo74euDBJDzkUYXO13DHlq2i9q7zvGVwgSqgrrxZZ6
b/iO7vFVW7UtNbUE1HVr3zAptZFrjSbfxZZr/y0taDLA25o6ZJGt+kXv1gV7LDdG
/sIUhGhRZvSSYJjhMZe4ADVr1Cu8W4DPxMVrb8WKLJKR0NbugteDTV+7gM0OvRi/
n9szuqzd4R8YiMGS9zMLn2RcexKTUUTvkye0GROP1trlf7COUNTZ5AHkTC8/fdDJ
N99eZzA66om1dleqg75bK/NIeoBwF7BQNiYrPgJG/26tlGR+mlYsz0v/tljTofhk
bLYuXyycRsvCwjtiVegccDwmmlDSvlymWqfVFfziQ4uX/ZHjMyFbLXuTWdjLIjKF
P61LffSQOclI2pu5HRIyqOtC0O5R/dF7ldkdLVhqP//uaXDJ8s/5gRT/WV1qdSF0
TxkzYs7jJ2M/IbmWJZ4WSBNOcZhZGFA4F5HWvCfYeqwK6KJceDpDHcK05ImLYveO
qZcuZ35UinQ4e+dllOV27cGSVaMquIv6cYJ0CHi8DPP7igRpHwJwek2PGZ+AjhsF
Uda4LcUAYK6y4/nHl2Z5O2Ie2s957vuPCgEgvE1+6E9OeruxysMVo6DVp01gX2Si
HtN6PmeSeIUYrIp7XP6Lr53NxdxT7jR+CmY6YOyMzqt+0xQK/8J6mfKARmQyLnq/
iA6iXDhevZFxN4qpy8iEfuo1z+VbvUFsZvLlaXv5KUJGfmOzHHpfqsVIGcoiUexo
FGcsATXngqhsCWLRvH2HTijLnNO+OTG614x0rWOwNGi3OYJhrLk6eiJUe0iD8RXY
YV91pCCJIPljsVHIlNg+mnlM/4R2dFOqMiJk6n9j0YHX+NPrZ/Gn21UvHqiH7NFU
SnQp7uAMVmS/Cd6MnTpInE/By+jxJKXV0ZK1mRg5ZmRKt4nhc7D/vvxUKjilKoA/
gWDNsAkadoeGCNWWX9AHTU2MD+Pc/xyO6pfE+oFm7I2BwBKyr51jpymM4xQTlnhf
7yjh8Lh753+8M0Ww6ssIFmq6pU/74XKkD5QV72AA7k2YfAz9BLsWpxeey5pSDKst
KcfrZWlQtUzKwgzr3JYn3CNPmItgO47ijL01Xdul02qXp8LN7bSapC9WTkmGB6Rc
1PxjZUbvf2/rh9PesVo5jEfZIMla/OBE8xfaho0ASSIurPwIKme9zbE96YITeqya
kRhUQWfRufGSaiaGX99Z+s0MV2fiEstY06wR/1Rcz5VuWs/m0JLcdPqNxnyWcDBC
LSCllIZAnu3ekKW/RLgFdhhRdCk0a5B4/MO3wBZO1gndX4yuH8C2ugFrfp9cFz8v
UcgS+UuGK2rpuhPEVutXYilCLg25qtWZ1W//RJdK0GyAsa7IYQMmMpeK1X0XpRUm
g0fQ0YvdPhw9LURb3JkATJt1vWEFx1Yg0yPy+hELfj9GF94R1F66hJj69eRi/v6l
64KCgB8DqBEoe0h/QzT25kzheZmIfEiJjubA3ZhFkZbieEe3IF34J6ymBK8soS+K
yVuV1LYbFeOx5g7D7Hw0aWBfemdrXmvfCggCKD/De5M8quUcs5MqaKfYjv58wrgS
lpNxzmEmCp/bmzYe3ns+8jSFoEcYrMbiUDk3mFtkpG3PDhM1BZpM0XivBWsnePkz
ECH1pBaZMSOvGNn9999VA+F9TqSGSIxJaXSbJyICQuvGBXR551w7Ru3de9D4POy7
q1fyBvlt0P52f6CYl75v/kWsBYohiIYuqYsyVyFo2w6v5g+y+nxNjNwY9dnmc3z6
3NvSSzm10awfkHUBbeEqtWShXXw7uamHGJaFWKQ/aVMraimMEAoBuE0UcRXeyVm/
96mItjrwQXgV0HmsR3MTVDyUztY3pHwMW7WWXvOtUafZ0AFRlimwEVZe97ogUvAg
jMGDT206WzR4mpQ3vB1Qq6p15zurH8hssMJoKXzhKKlZqwgSIj9KkUkozkNTRnQJ
6kxU9za9OXF9bgZV9IRV8mNgWeb3YsoglUCTLwFw9PntL4jKOk5K9UZ52vmJRaOj
DvZ+QlxYBe2iO2NHRPpTejE3vojUV8vnibR5JShceuGQ7U6XE2132qr+cCEmWhwz
CnYWoGHUZoeBP6gxNEyFnySNBVQLJwrFMdq/Bz3xQhZ50cgAvC3v+zmgX/VRU2nv
oxdaB2jM37oMIum9gNg1lt6hzeub7BzkF8GqpXOt2D3dBq3cPKlOQ+3mmwvGnK4X
8je5JnPnvH3T2oEioGAIeGXHAld2QdZdwf2hsxJUHXADovqLeRCwaNoadOdYmmXw
s+NCqIGCWyZqFnRaMvva6qsk7Qj0VXxdx9V+Xs+ZlSKwTO3x1A2JjrPfXm3jqY7X
x/yPz4RuRcfRkVJwgOlgHPVywYmMvZkLvIf9p6MfCMfQoMjUCbRZju2Enqv67WMk
sYBNC4RDsRX8FrGzxxAzzqhsrV71zEN8MG8/Tq9cwzJn0Cp2+iBfI7iXcYi+4aVl
tGh2RLOxTZDs8fqXJ1WuKvsxRDZzfYFXum/zxTh1XJAZXlSXCHiVF2mF8hzSPhyT
gf7RtZPrncGrLUjyM0WfcjR83f/KqWx/fX5jrUaiT2/QpJFbUNP/yMxX8Vi5kGLb
PWP7GaKite40PSofvO2paFazmeMLi62ha3dWDq7cDPZ8znwHTQeN39l06QvSPfx6
DcIoguLFdJA7VaWO8b5b6pTYrSNKwMlYCPUwjHE8owfCArl9eAt63gUU0K2sHSRN
l4n/nW8fqmeRvY+Wr3nQCNVq9gQRtkwt+xSi16x66k/WND0S4IOKQ7/guzdpRJmK
cISVNWOv5t+OIyBMo9b1DYTwk7GzS/7rRrDGgzBWgGH26LsIMjMIke5an/o5BniY
mpBRh76Yzcmb5xITpSztL7AeUWVRQyWMX7a4/7HpR/O1+Un9YTHks107H1zbq2kR
ReMNe0tMqZehSZ0PyuvNrWv8Hd6+lv+A4dcuI/ww2onm3GZadyj3Jl/OzSj/DPI3
kwV8hEERTvWKwiZFf/ymOu3v9z8crv7/HaVVnwJM7vABosFBPijcBwZDwxqswz9r
Z8WFO7h6AB6Cpdjy3D1yJ6hpFndLbORujNpP7ZHk5G6GupqIJxSv0gdYmPwtzPkJ
fQ3nLtF3jQOD3lo/MUkYJY7f1XKpBE7eaKTS22zs/37gCUcd5roQrcQVIzwg/3lH
Ya321A46PUxKNMJ0TmRSXc4Conz8xhGQWHDUnSl8oWMeoIKdelK/NevigwcnufdI
UYXCDtPtt5IyHeX2yQWZ+Qs8dDumPmz/EKaHQgGSGFV4K7IAbXs6ySZEneV3Rx34
4tvUq9yX04qbo+pW4/pAR/vsuSbKKAAAq5+E7OFLGBaU176ra+AVBqx51cWt+78Z
or9SvBaBfBxRtDi5OqDygO/DewWdkfviluyQfxBGNoPR6r+Cn4z4ns56Wi6kzelO
ESjUevTp4qE8kLdLrKcdjV9Vxe9wRR9gJTruILV/EAJnOywXiHkcQ1oQ2AJGxvTX
zI4sQi6/dFP0IC7jHeMZnAWuniPrvI0A41uHUoNWzTl5NWJQ+Igra4R2FC5rJOr+
jOMxRbkgYgWUGgwOxPPZt6jIpDxFGJrl/7YNJt2QiB2HKV0X33QhDuIqkJIxAtxs
YNT5WJ8TXSzRb+FYOlYilTMRTHuP74OBTY/vzK7G6BFAy9fA4RDHfcwjyksqqhMl
IUl7vOQFSi4F5zcvjCiQs+pVy4xcpmEeoG0vnRuY4F4finosHSX9Qk23bz7IUC6X
hoDqLu2FPmrpb0pO9W30ZxCXh3vmM4al68ac0CjbtJTpD99Rb302iScCqjxVuNge
+ckw9utzeiOmOYGE0edG5QZdAtMrmchyYv3srqJW17T17pIxD2dX1VNh8W92Tyzo
1zsFNSjObAJb7i5WJcrgbUe1ECOCfle7S7cqdFuhbcza6Vufe0AukjAe4X7Xza8C
6+9qrvwGwQEzK8Nf/k32hgStNYjKEoXaixjvM+kkiiSfpsmhQKv0a7QM+VHmJrdc
3IqJ8GhiKrbSZ80HnZMdCZ0xkkq4RWBIVhG7xbu+J0rrZgduSRJLGhbR6P7u110V
LJmgVnwtxMTqA/asDngbaPDmIACvRQbPiSFLVLka411fazlq10eg/PsNI1BirTE0
yIvSIXZWPn/viYQElQdV7c+Cn+SbTAWJGZhevEVsBxwZh1ClMx4x++r5aBYrPrEG
DwmKuzz+tAIO6zD7sJ6DeRMtVU2jDB8QDIeanW7YEVSYfYjusf3mUeUYLBLPIiwS
S4TrwBU/D3VuUq6r2S3gImUMW02wbEXm1oBgBY9dovv5XgzI/8ux+fXBE/irOsb8
DvHb2wYCDGRb9PTDeTPtQbdy8+jxrXEJ+AghmwNX0WqZK5mFEJO+1JxinDe/bTyo
i5qO37AIkPCFva4bJ12e7+Lh8i+5z/TzD0MwJqePVwl9BgAhAOERm0kv9DBhJ5TS
z2iptOvDDBVsKuvUn20aN3tRNV8Kg9zbDQERyt3Icg/Z+GonjFlOUOMWfKIJEM0u
7OCRlefB5MZmT7v4ncGEQ6PRjorwhQUongDMD7WYDGIwWKiICfWhlseIu66NiKik
XCgk5qbGsDIbBtARPGdnIA8KX1R9AtczsaxmRBFSzXB/zktl+Y5gcd6OybA3Yrp9
Oj3OCEG5dUsKkIPZQlZoGkQGAHfYo0l/2x6psmQF0krQ4M14s+VZOt5bF7y1anW/
3/Yl2x9JdrciG5Ul1GTYeG+1xZA4Il6SctdmOF41MjKh2pueJ1nATCzloWT9ZZfw
hQ+97yTCcMkd9teaUzq4+XKnoJKbzUe979+yPLZqrezZt3q+u2J5kInJmGRH1qgW
vho81ss1fBCeqzO0PjQtZcucrfEwlGjmbd3tREC4REF/ICZT3Tiuq0N+efYDIBTr
LclQIzjIeNOvrQsDbOXJ6ArmLKojKHeNIzt0+LN7q1khdSnxI7tELcAU6LCmQ65a
ciMdb8Y5RdDa1ZZar28sJqqww1fXCtO6mmZr0VvtYvF+rQASeU6AhUyYDMELZeXd
NtwcEF8sHxzmYdgj3DGvQRvEFSR5hXDqc6t6pD6MfUQA+y14/zJJbQu08fu3ODC0
vrYW54WmnGEtKTfCyMKGqMyldsfT6cqkNlhVqCzPL99hHrDmMh797zlNW/OPRELP
bk21p6iRl7iDU3hPw9wkWlCIOncNW6YCNuT0Z6RRMkPjlgMcG3uglOrNngVdJSFz
NqHL8zqJKiiXBjC1gtbLTkHNbF/Ri3qNiZS7W6rY6iJfhdr51/m0wpdeB2/OCu47
zuG3xZQlHboAwXxyAWrXwFitIpXavLi2bqVv2dAeqtW3wb80gyYLrHfqB4NCkvd+
r9pX3GRKh39QRPdGs8qvfX3jTFpd+Iosqj85Gt+/3Ns4Q+IllE9FE6R0u6Bnb82j
3KYzQiNMUaW5PQbau3/Lwf6NTtdBK5h3uqpS2nsbQoZqkdnnLuDNwvE495UDxaTe
3ECO3IdfcP3+C5zV7iI1HUPnSdQodDOaA2egrkR+CUcaF1u+P7MRTBnIpnC8SOGV
EIPjEOWx2ldaOY6CxRL8xBF0ZmoHsAfr4xqow9L9FpzizNdU5gdPbe7lJZSN42nT
2FLOSNEzTSXkwIqb/9NggqJTl+pMKKBZkNl2my9sN3oM52oK0jnBGI6jEOnPWQzH
glDmsWtQ7b0Hh2piMewjU93s39xFXuJS0FbuIMIv67fuwK1Uhr0W17ePqNcPjIcC
0gZDufSElrP4UThLNqHCrgoiVmxOqxgBB/iOEBKOTQqtZaj7hGCVc23MOmCdS9cG
QRJI9bClPDTsW9/rCBTF6q6ZD/W8HI54XbIQnOYIjbyFa3XiY1KbfgSjASh0dDjY
v9NqqTkkZdAoT095IEXAGQqEWa++OBKceWGYx+wY9RI3owHDH0L/9vr+c4cJn2GT
2TTFfChPAGzCYpHawQpoVh0Yd4jfAlJ46ZOFmemFBboZpv5Sy/xJ3pawKViAPNWa
Sv7WTdA5tQj2TUVoSym1zTwMVJQucW+REdxMZ5dnr8FFZyKE13WFZH/bQOWpjkaO
p1CV4m5MHBTy5pd5ofZKG2pBKdJklL554w4z1Prj2ORMob46xw2Lwz+IoUP/Ok9y
c6mBQRVEgmVUAJpgLyORYcdHR7I/NeiKkL08ZoMz7we5oHTUe/S8GEyzH06J9uSy
iMAAf6JQEgkbQIVoOP0EZfN+YRuDKDCoIWlum/9Zg7JvvtZmIYPIinwH+sdbQEMa
9nTH2czBxL+HiudTSa/n2R7oo/rGcyGHOLYlGq+EdELW104SnYWv7BpAWvzjy6qB
lKKGxOpofFIFKTDxBixJX2Ymzs2zVOif1UoT7HF3JXX6L17iikunSPeLWbKNh8JI
A60WUZ5Rngg6ePszscgU6xyPPm/wGnC9GMvFk792p1czzaJ5/EJ3El2ldzofviFu
D/u3BFeu59pvJ/hButDZ1+qlQcp81LUiYkQp4DuWJPB90y7sqdIv2fodEKVx3sX0
Kg+GKI8cSXXkuTXbu7NNOclaHM3RDWB9hgqxqteVu52al5PoD/XqjrwZuGmift/t
CSUSqfXYNoE20xhp12rkRPqeLYXIdt/gT+Vjoe4m/mPnPQeAK7nhijNJr7RJZTXY
1WLD8IQQ2I9VG4uV1W/r8s66hc+1tVvvZJf5VLkCtI7AQHZ+cuUIQJtmnUm1awwP
XNdsF0qXfHHMJZAbaBHwd10W3kDI9ycIg/oDXyZ+M6OvdedZgruGOfxvRRPBV0D3
qgNnMVjqQo5eJCM1kMnWfVlElZjpoyTVPQdxOuZzU1HHNERzFRE5jLfir/dXCMJi
u0Cpl7n5DeBiRHWWOMVilk0OvuREhufvigPknzY+U9rHLLcJtyzGxIT9QuzB3kn3
sRbjeRlNyEvYmqjn0PCjLlObbsjsmX8XN1C1qnuxdbdzz7udCVmOHHQUgfx1QPQz
FiMjJzFi5J564MfKkvy8TPRHnDS6+kizWh9Txa/3Q9bdiASZyIz4p2nN714TeJQV
LpcDyik6dGmjt3fmZLqgMmB/HkdRYXpJJt+tpax4YN43IgaCEXCMXwFaGOXtph+s
M4XHmF3i5EnB9jTqyYeNL1suhYTfamz1/PqBYg5i9scd9CL1ppf0/pLngxESmYop
OZSObK1CvFesDco3d/UbzCidxwleWekYrKXssJFUqddikLK4/hgciiUwAlIb36+m
uIyvKQw+i4kuhrPypvJq7Y11aBfmqX3gesTuBJSqcEFkL0D9BKsGPXz5oCdNn3oP
3bXCHFXnn0bxmpN9wq7BRyaglm2IJZr2RPd5nveAtAn9He9zd4GV/4VGpoFqASZn
mLZ94zK0joVplhT3XEgLjhOrSIvxZVsUnqw7KSKpVzfHUL8NkVpVXaCE954D3ZG9
s439n7Revyhn0NVdM1m2AANTpYlZEo6fjb+AQAq/Gh7LInEz11LQcy9Spboy2Emt
6VbJm376Pt2iOjMMNRXjpRywfwy+HdQolUylrZc4+uu9+Jy2eI1evVF6SLNpyBgz
lxG4FSzmg10zDm5n1IzvFY2n8SnyzjVkZ7PlePGz74uG3eNMFAhjfyproABCk/hY
8J6fW8udwCpI6bAYoL13sr9WR70G7vcqnTBsyFOmhiVm4ZPZdMxgLFtJoqVcC2Ka
ObdPWbXWdcBPMCLKK6BO1Pc5jMBZX0pDK8bCrIb5mzj9LvK1yUq8p34Qo7hx2mf6
kh0AxATj20AxS7mslcpPaXs2Z6ebhtHGIs3wZXwjU9M7OVzesSC4NCxHzQJY0YI+
UBxNUfXVZznlyYb2PFnipBtw9xyWo2+QKLF71YzLitBnpWvTutReq4KaWG3mLu8t
tUmwJ+dbiXdsw/et0UjcMa9YupmyYw1TxvahblMfzIZiucSElm0ykSNUqfAPM+Sh
zILON/zCaBOHHvUvBI3s5WVTPr4mTmeM4d2+4ftLKHjxt5jaqx29JSiDMHXYCJU1
DCvy2ssyp9pb3h5RfgkUv5Wc8KYv5rHsL/QKcoCHRABwlblHe1/IH+Px9QD3kUSI
gPJIsWIGSWVygyqBDO1JhOcUtw8iMbGXfedtrPTlE93DvPTHeyh6COTMAI4YXXDy
tYPSi72Hdvg7q6/DNwmbfUrU6331u7AyUJCwPlnKlkLXyT2n08wHqu33/Nr9fto/
fjBAYx3exDBXmuf19viNotYOmkphNzBGYSMBUqKS3K8b/cVJLneK+KTKccRB0oaM
B1BxeAW/FUl6NhNKCl8pp5NET/4GPZbLMluVJ4pf3grMP1jiU4P3i7iuNNzzPVAi
oSKQgd9uQKM7VkCTZJXvgeO9UNUQNWCC4bptsBLzRIYpFoNdSC3eIfl57bAK6pUL
+6U6A/Yo9rFr4PF3BRbUqxvmbSK0aFsZkx4wsGwaFyicE95H1Crey4MscYr+mNuS
heSoVjJHKIcVvV9EEXACg9vBoPAVId5rHTIDuv2ikoCHpmKPi68f5f6GxK9iT7UU
pKw7rz8R1R1VV51p01qHucoxcDrylZMeFVITYcdnruc91j9jh4l4IIX1Iw52cob6
IehjNY0aTBojc5NLbFSqeoSPRlssOpPxVwIIr0y8cHDkKfytC+Kgpfd80NCGnRc/
bWenG1IYFi9juNrDr7azfZbteVrOH/a2Vm8fsvbUQDsKS30SbG1ahGGK3fYToF6m
QU0zJaezVkobw36Hx9LM3ugMrPeJXs2ST57iweZs/6hnd1RjxoDCp2LaEcyDYNBQ
/mvV5aqNiPPvgNHoKiO4VvbqfU7gHks8nG1TPx3oXyb337Sgx9S8NwVCQZPnmOLW
zUZ3n5wB3i73zT0fdf789/lf11CWYYSLXaNaSv1Emrmt1/o2imyuh0XISmibYb+H
DkgwxRwLGDA8e8R+x0r2qHsP/Io4Ya7UtYvpKEqK0189O061NtdZtj4hNYIl+gIr
ILIl8fmtMrD2eoe+sK31Ux7+zkSB/iQjpqePUIbHuqMjyUerdEoGT5xB9AriHpMd
DwABOc9T6QnA6AkJ9B2pKDuevOSZuFMXXGEB7vZReK145exSdCrSVAgAakYdzS5e
CT/nfp+nhoC5LaohNio3MLJ0acIhLBTTtkHuwXs4ORiqLDiHbJ70zi2PX3p60gqf
WyWbfN0f4mgDbn2N5PIwPq4VxD1JMPq5t5598ypA679K0Gu/NO00Ea+pGt4mszfd
mSjblM53FTZqG+5MNvAeBJ1AsP6hOcwW0vYtxwkeRJfmgltBbsgj8LGvXK+GGwPy
UbIyQ/MQTL57RmVRCzWorWygPob/KQZR+ypE0N0qCUSMvXp4wh+f10MGs4xkQprA
+NazH3ogCaOGnuBGN3fXH5xUvBbN/KPfpiaQOf+YKRXJj/+t0B9QVRu9Z1pOaBeM
OiqaAeOlY9aakda82uDNKOfrOanidHPpx5OlQnNK+aoa0KUI7JNhlCOIqUm54KVV
FQXyU2r8R/tk6aqKXSYyfjoBSG+oQ4ecxCS6ine863s9QXseAgtt5Osce5l0dUCJ
8I2p77roU+9A7IvIl9q/0fjFpilbl5Vi7+O8K0cgXX75md7H+uUuycylOJ9fKAXH
tf/xZMrC7BKVJrqx3KBXrYFipIXnqCwhZ1z3w1+RhvggLyb1YUtxVSU/vj85Ez1p
Bsf3PcPXRPVS08ZioPvhIig/DQGRQ/Xl/KItmpPKkiBbpRdClPgEcNxlm/r5LxH9
JeEu4SM2V20/yBBAdwMVgYMd4pYSKa1H5OW1b10BI4HSN5p0oqKvA6Ply69kAm2U
aRFRz+qPUhTIecrJ4WRVnyOIc8oBsSTrKesU/0Qk6QpY1Nts/XK2Fl4TCJwsa1gF
qsnntUHYZjXTLszNicQupFFTjZbASwCsplxSKe9/0BFLnuH/1unbZhZWTHdmRG66
hE5ksffJMR86y3gh6sUUEuIHTAftP3kkfjkC7YICWKonmCyIRF/U+oNQXL9d4I8R
gABP3S8e28cWXwA/ykZobq8Yts+3P5MXgXfnQHLrfnXov0q/ObTnBBLXW0kRqW3q
PcEY2yP4yEZxvK1C7rbUMzrPiAHm8jjxvjvIzw0lMXkC9HsgmQ03ut2RS+svTXnd
eql6oazDb+naSolqq8CjENDa+8HfknlCnI3RdvAP6PzMqeDHOvMuo3m09Yp54o/J
Zhlj70DOy0/wOzPFcaGw1RRVtLkHRrHB9mnRWTAav0r9GgtbTU/wG/JunQIpg5Oh
g/87QKIMk3T8W29ZXn3UNKl6EPrNLAdAH0cZ2H65zZESFd0SIMQH6H87gxDZHaPi
z1Xt+4X3x62RO7Yi/N+rG6WSKmeyxMDztGAgfOfeLPTF9335PeqtTUCAadBtE0DQ
UY3ATjiaH7iiTSXNAE723UkizKawkVdL+g4lD7hSDKq8d4pIylchPFqzxfbPN87u
rw8S3L5d6ep04BmdZjpw8Y5S7RtNdUcnFClaUvY2YbamtUxe+KqPy5YtbM86uZwX
J8qtfyma1COmcOQ3+N8xM/0dNYmD1RNu4jSZy7rn79isvVeFa4cM1vJqlZMf9Pug
u9XbpJtrVnkdLC8ezj9Gd6Dlmkz4JexYvwPxsOnQdyah+4W/NsofMSfFfQQKN+r3
IHaBnC9Fv/Ehi18iR1HXudV2MUiI9X83bGVvbqtALcg5x+jBMdi94N0LHBXDe2SX
fKy9SY7hh1hrWV17MB+K0wP2FTVlFmlQ1NnIUgEQ7uNWzXoKGgYxPhGjc9IFNcMS
rrMRRs5taL9WHaUWNFS8VvGSrg5p3eCb3xs5jwq/QROF3VIP5zJc9N+ZT1JHjb44
Byy+GsVqFxV0iGDgwIcDoFMbok0w5SLOGZiMQPnQSNCxnA9LTF4b916xzm/D4SqP
SMQkQeAQiQC5dguCXoha8zm4gIBbeUhOJvGh+cM3FQQUyGzlGNsNARd1Qt20jLkS
g70cpmvjFbbsr8sehdg5xjlI5tAKnQwwS0oXPAbPHcwZpFoc33wI3HZHyS2p2shH
x7GD+tKnkVRRXK+pUznXkkat3ejAT/6FP+XctW6/v7N46ft1tuus+gPbRbOjpp8A
DYhT8JVnR2Yg9V+lGRTpeTX8z85/36PKXN+nOvFl+wpi9MaXqpDZHes2dmCBOTDc
/ijDr5cxzcdpkLxjIdCjjNFDOlJqCj6A7ifHcdsZjYALSxl4fUtZh1nXgOEKEwQO
4lVXf1e91VS+XpLL+WvsBcMQ3NFVqOpxeukhm1ixD4aOpsyuH4/j6pRTXJqTDekS
MP2NdYjZSNkWeyI6kQJPyWHRwG5OE0Jr0QuIDFaMkJUHvj/EoLqDug8D2IvTVqET
0P2P1iDtSkvG97rLUg6B8hCM8z7zIsY9zEXbuj4kPwXEZcNVTOx29bHiMkRbLMhN
dCqwpxSgXlInnNMdJkHD1+R+y9jx4ddHKEYV97c4x0nOXQu0C4YnNcUjTv2WkGSH
zHQ8PNxco4+p/6J6L3qbu246pgP/OV7OKNZuzWdchUSq+9tdouuQCL4eboNqsfKe
In+CVXldq+yZx4bYVZrBPNwPQk96XhD4zOGtggm0ceZLD1Ko3zIy5mP+dNx5IAZt
TpxZYDhHA4k2q0gk4KRwq1n1hqtzm/BieAFXq2cyF393rpoBsBfFydORlAK/sKFC
WQX9wpo1L9PtN4u5ChURJ/IFIBhKDmgJizsgoGXZdygO9ujJlDxQvfMe4k0sCP0R
FZuM1Dv5jIwIur+xgAfgEFugYM/n6k2bNDWml50YNlD0CnqGpSJdWGBCdMTjAkuk
aoeD0pW+gIEtJ/VOJiWdzsNjQABfntGSUzf744et0FyZHQj1oyM31w225cwZEF9y
ROCBel7LW6e15vA03i8bseh0Qmm8gU9+8x7ymhhFLQrDFyXH7PqZBAOrDLWC3L9t
bKQirk1S6IE8ox51qooUdXaKKwcnW3cr67NfXHI11wMhgDFqoqE58ErJuV+cJ+11
cJlO+2qvPV39bh0bMjwmCwxwPe4+DMvgET48+bUhyXFaCgucuZVE1rhGqGZAjW8Y
bv/6KPd9tcdLwq+VO1HzRDfh+bjS1Opr1zXDSSSX08XKwgeT1VrK4CAMAIF38Avm
QB+NB8Yu6D+Azg7S3gorsxLRB/aeN2LUQq2d+yOrZxLhBsUP0cOjepbLEwfR6d2W
md9dT3/aQfab7QUGvgNana1QGk+g9lJJ1tRmCsyokQfmWRicnyYRtdRsExuFZQrh
PYZG6rgw3Hilg+0PG7PHkGQlX8iTxJWGcn6hXnC/UD3KbIO/7OJ5Qszp+uvdpvAY
t/0TEs64CYdwg3RCBKfADH/oH6cvMERgE9TsRKT/TYbCS24kxak5p59/6xOBFVxj
P+IF6Ewhyk+80Dxu9y5EBtPBx+2AL7fCEMLcHJNBkK4R8NvZtBzuuj6P/eV5EspJ
HWW3AV8XJFRZHA1phaYy1yTo0bGOna+6NH816bV3yu65A34oUpi19NkUsbRXyDJJ
hinVKW5D2o5ZYgtQNHMPk9lnCjoSXHZ5JVWGVo5+z/aUBiUaevf0mIZMUgCMGg+n
Fm6slSE8sCmfU0N+4c4OkbQb8gtAaqsyPjXkqViTxnvNYS8FYwVW0zDHZWvXUukN
dYJPimdAyQHPm2Lq5iEmsZAP5eNPqh2EDWkl8eM46vvlZMiS2psFO93mfm+SVXR3
LJR1+O4BpDXLApG/s4asYOJc1Szq0q9N87KSYZ9B9BWXLpR4+o5DAE5t56iWsuiW
+XbC1x+JOUlgV3VDoiRNMMpdHE3EKbl8g2cWjJPyugs4CLjm5hJfe0mSyIpleHJQ
pPNNqs52Eoq0Pr1QnfvYE/Llwck9BMjGWoyAixgu0TmNWDH1eJ0+TRDpH296du7M
E0tZ64dviTErNMuQkWNnFinpj/PA7ssh4LipicSomZATjhDtxUu+TPSDIIXUJbOZ
e1GiRIyASLEC+28GVq5RVGFm4mSJTGGqbNh50w3snGaIsWop8QiCT53G9cdhQ2ze
uFJzywNBUCBmqKy/gbaEJLr11fMfUjlhhRL/A+PruQn4jrAkW34HlSHaQOtOA5Yj
A0FF/f96rejqt61yuMYOvU0jiny90BmLX7Jf+fL5crSCVh3eKaQrh3BLcHVP50Vh
XYDg3Uji74GmYz4UCsXw1rYrxavBnBZ4SN1dxpM6HvclKy7ZeQ1yDcq3KeZHG5Y2
KwMWwArBov/99UbWB2STeehD1PLP0TEcasnn8TzEUxTtVO0v1onONohKDPZ0IYpi
iTbyqBRlNhPPGm9Da0Xk7O/WjbvLQpeUVC03Wj5GwrQXGWeofoknWEmxx0EkaCHB
qHyHAQPzMXewxA1yJ/5H8h/Q5PAb62DYK2aRV17+UkMXIza1yffkB1eSLKM+x3+Z
vjJsmTvbwc93QlLHNvttuiv6rb9GzXnyRqmSnvRXL9gxgbaj4T3qeLynyOmfbXEz
Imj6ytDDgSUQOz5Dm/ruHOPB+JhVAYpTt8AoOdF1bShtjANfL49PgS6axpzK3r1n
i9WBb3ZHyt6dd9lTwDfqdXMaUQ/Jcx4nrepGFWdQRw1+nk4zo43nKR0gHhX4dM40
bG2kxMjTtd6Eo5z6IrfLvbWJuYV2EQHvppeQQkPKld9yPMrST4kQNbAWTJSlMT/P
cGtJIFwCNGRdt6/LYF4T7ICTp8dzvcY7zUhWGNFDteh6IdYuuIutwJYna662Kiou
ZUIQkotKgodnyMXKLCE0pDLjunrRGt8VlcAL1zyx5T/cusT5/UVQVCdG6VO9eP7P
qXwPl/elxLkjMH+K5Wp0as38Y6D0PPIuWPuZjSzfNQVd6qaw0TqPw6hhW0V4xEi9
qgL8C1LIaLaxm/N9NaOJ0OS97mLaydDX279A+ZjWRmtbVfJNJvsSXLdSpvrVgbVs
OTJ/fvdJUiK+cPKZfTY05/DKsS5fPpq35cgFBrJHHaJuxUu7+Qq+vIehv7f9M3xi
ppFM18TJukFshi/ZYqw14NQyU8X54C3INE4mS9EvnhZE4l4UYl2WYTeB3MNPts6H
F3fB8QicMZTTE4pBsauTdNfnciuLMVrywaMejEAUEi7/1QRzaT2PqyNO0YZq/cy+
iRs/HIZXOy+mXGiuTW9mtH83jmWj1SUjK/HU0V6VQKif2Rmw0A38giEjwkWfaok0
W1rGHkAEDmI10yTybSOny6W09LzolwbqMFS8P/VwZ6LBkuSqBbA0TkrVUzujCfuj
Ti9Ruo4DYk9ked8S3p1JCOBzPBYTFGZqNBiZ2xgjQXv4+ZGwBX6IPQFeqiovHLy8
fb+NyvwaOlv8Mu1/6wRapuoj6B4vGNuX5dnCak82u1QB/Q/b8LwTJmFfvRiHwOES
KCY2QNXnNzJR9J340CbXHwuPzBKZOSKgZYPe2KQBBQPUULoIebNl6AF0hwHJ1biG
Fi3pMCLHkbWkbojDuZdew5Vzt5sDjtIpN7H+rydv47JAkar7tzlM8KHqukQxmgVP
U0TW7M1q/uabNgaURY93lj6Sut+M2HV1s30FEiegt+w8pCqD5u+t/HG1OMjsP2ac
WU/TVc2paxWDLknrFqC4SmlFEOUuHao1oB0++lKFgSFU4nbxF7UEFAnyYT/tCwLb
fgSJ+Ucsda8hd8hiG7Ndh44ov57GXp7eE6N+KcxcKVC+u9oKDCeZfhJp7965xKI8
tk2QFuwsYuG6pTrJ2b18g4VCjJGmtydzwolo6OY56kOD8hW1Pg3T4/k7wnbWyPqU
E4fBmIOn2pSC1yqVIsyVyT9itKY5r8e6QWlJ+XQj5mYUQzSWjFPq0ZN3rn8G1LOX
UHDZ1ImemYZHknngHfJZxlLw3KwbJH6N5r7H/VVahDSWoZKbNQ7WgwTgUReiT7wD
Wl0XqgEm7I13NcI463GbXeIbSidHXB9hMo/4jsNA5NfiiLmD/GeNBSoga/AOWvyF
tTVa2TuYdXcdGRtqWEC9efwHWsQ3U14aujyTl/lrPe+CSnnFQNw4LS3384v9cD2T
qKCKCizxE8RqKBhc8vxR6G9jUzzYn+SVpLD6YvacPwXWhLtlk956T1MqIC8bvYwz
WFASC4DNA0wEfcBT/9GrdSr+yU41GQY0laGf8b9nDmGnNUtLDL77ZonGYlZiEQw0
KHzRjOC4atHg0MNnX8Y8RdyW2KCpNFvnU4CSTAnH16JfjUXm8+5chscYJZkjS2ZX
DOixZZK/Wuzbnlj3PnNp1xZhPvUZlWsn8P93mvuHXYnsxHo6mssAZ7KZiZd8GSsx
nPbt7YZezEh9ycGwbeGF1EDvRgPdVAevtNd2g7643WdalDZjJBLj2cgnnQR26XH8
/IF/5MDX6vTHqiFCbtoNyxFf+gzfXBpKolOKSZO657pQkRS8jWYY1zCyZAPOyjtg
zhtNCoGmZhWBLH6trH9g4FWrAMugudhiEsCIRNAvqAB8Ag4OBP2o4langolrlBBu
ewo4MvkMLgN4KtOOGVnBllTUCQJ7gk7j+RBTzLWkbtO5yykxhX0mr51Kd8gSC3ly
sS0vcdQoGJFqc11o8WDcyzr3Z83Qv/wvYvWkU90YWxLZnh3kaEYUH09F7hi5grZb
APn6SY32YqFLeHfQkI/2LeTp9CseciHq8BiZwoR2tHntDSMWaKVniTms4Gvl5XQ9
Vs2TEylL6yr0CQwE5/hPWgzIWLchL1i9kE9Gy3yVUPO/1OFuttXhDq+hGta8utcR
cC7ULmyVAB9MjTRiUIH5z0DoYcgI19Ulsmrk72D5u2/RBKoS9Kbc7n0WmaSiLvxS
ucg82Xl7NaVACTLBSHkBeLCaXof1UMIBGhlFuxdKwDkl0knN9WfY07X2lD0lRPNJ
Cie1KsTt0jG0hsgVYclsxGo6LxDEyrQg8ZHX4GR0qer2r6+B79kq1W6oJOQWlmw1
oicFvj38sZiVtCtTtRJVosBgU/kQdZNhF0VYywpX5P1UeWEFoRzvJlfsUQmQ0wIy
KRePruc0TjI/EBHO9K+xZfk1F65u/O4HSM+Wyhpcmp0usRIoLi2HdGQeuxAuiAee
zt/tpNTNZvg3i4yjXBRrLL+NMmD2qBd159IwdO6klMYxQj789h0nwjSovoqhVzRC
ODkrBNOVngNZx5r6HypDiDCBxAHFhT2k+XXtMulhF0KFBBcy9NdUgzTFA/z1z4yy
zhFvSZjKa0vOC+0Cvc4RB+nxIPDsdEyuTZh80JJRtSTacckDt+fIYUSfGSkDCVeF
9dIyUd0Igr4WD7BPHqeQjKVskN1AJGACSkMsZ3grC5d6scrOenDWvinVOme0ieCr
B49T8n/2mtu7BuUrzcoVKmH3y4tV/OjfF7IrxL62/YvbaOVh+I0KQ3G1Pg5T8Zao
xY+hUfCa2n74ISzsDn+qTA1PIwtW9K0eYb2+9AzzsPdw3dnjSM5r3fGjzoS5Zjoc
NrvUy0hHTDBc77WRvPyBR+A5lgH2EREhZe6nMZ5KXr8T796bFTX7L0JRsENuSUc3
Eks9yG1AvtDR7j79l3Bw23aCaJLj792K2baLjyw/HaZXmxAYUwYuZ0dR+SHCXbBp
FXpLY05AbHzhWaY0wfzbbFoW18MQWmpuuh8urSCW6qTV4lDTZHgwj72VziIDY6Ly
na1fIGhbcn6vgnbnBPZtYZvComuwtq1zbJAZ/l5Enx6RoZDNt1P8l4BiYdIpfhuJ
cNsngjU9mZNBO4LDaLFQwUSpDic2+l3OHAOXkepF29EmuCLm80MtDNDoHNa+aJ5R
lFh8K9P5x7B5ld0e3wULqZMRft8WR6aDVf0SGPw0wXaZjUjcGdB+bm9u0B9UdRZY
IELe0NOyn4yrLX0fz8kQH4e8nH+rF45xtPmPBLxxzfItAk4ANP+G0aeHivgOlBBx
05grstKrgKpxl4qHaAGZzHLrOGQhsx/44z6BvdU5D37swwik6sv+7BgNNE140Rsz
vY5qQPDDxzjEID1zDrHNklXp0vffafTwf+VGno2OJXREVMd1O4/OTmzFj9k5nZQv
oa3GWLrwnzO8B1B1j4oHEOwD1pIA5JDx6ZnRRuo/a5zwIOU/Q9N/4wJOBkIKvv2E
97OEauefxrhPjum9EHALshN/oQ9d2X6/CWWRKAoEV3C2DV5Z/THjK/uAepaZxztD
EiojIpJb0e7qWh3DP/A9r8u3dBx4C5BT5EIZyq6k54GtEfUorRu6qieJUkw0FYdY
YQ0b/dtyLEmTY3TNouBJx8YOOVqvKGkRHZbE5s2gD8do13/68LR26Wc8+PnChp4B
VhseLnvHrqX+oNhx1hqkRqUr3N9jwdtm90FExI56pJyaQy7ElB1b8m4lQu8Rg7Q1
ehAqX8yq0yPvbsMpwvDui6X8kDH7uCl4aV1zKBwnZ4q+GWXhHHnCAUr60QJEGuBI
9+izlLqqBEOfhoNepkFsWKa33sQloMUTWJNf6IrEE/gWwFLJTKnomPE+1JepNoKM
yBYKYr0NgYa3SM0pC3PImBYavoEqvfQCn0xFWEGqbWFgeIyCEROTn3rHGCfmwetz
pYV6Ntggxt6trgclDY/QI5vPCgqkIJJi8utvNNE9MnbY5g8PZpF0ramJ69/QJLYX
K5kXV15KU9R/1jDW1lAjfRzv6/QgAJUCXzQZORuScGqAe8ieG2I44T1UYvJRHgAD
otF7OjXDPBTB59+bxs2wCnLgVGfHhocJ3+xmpDwjA6Nt2jkJvoNQrZHBsOf7KkJP
E/8vnRRlnXFDP5tmdFPbvpp6DCjHPZP+LY0I3JfMForQw0sVKhxWHw5nMWRZF08z
lNOzZUFFCGNhKmBtaUiqKnxAGs3fNJo14VCF13wtN+oR+Jh53MWNBBMxodn90gIa
ToP2tVi/9rN1acOQOFdf0mxcsyTs5CN+JwXXUw42h9SznEsipB5uel97TpeJo6Vp
hLI5BzxOZnCoP9g7RfnVJaAS2F/HKHCCXi99Xhl+HRvh/3JnpEi1iW1XPOurw2me
gh7Dx7VjoDXZnKXx0icRglUkvBvRnBBDMafP727nV2xfQvKGJR6VFbChZvnpFvBe
EahNAiqmAg71miT4ldmm603TDHXEjgbhDObpgLxEKTjT/oAunHJDjxfdqakq8Mbt
HH7PC8pG2vY7yHxlbDMXaIjyBYqoKkdL6S9YA3K3x5P87SWkUGHQJNFW1NBmjgNd
2JqvPOTd1aIdoX8HbmBpJFDWE4/fZAfNrInVRfGxTFsA4GNZG4PoBxvW6XDsj/Cv
iX1TbSDQ7XD4SjxEpUMBnMozHUwKQrdy7fN/1w1WjTe/kGiwGsLCVUgefOCW05SG
BfF1qRT8F0jmUrK0q66eBCkHePOO1s9BSI3/yFVwzjgyMmGzsx4lkun4vLwjFAYE
/bqRyPh4yVTDZg6T7zfUc20zwCpovqvRdasF9pp8Fp0bwCSBwYOZWstB4o4MMboq
VPNEmgPRrEWvPVshzOdqvRarNBKRLW8zmgRUUUUN1s0nXcztYQTWCem+i6hNo+qg
XAhIQTGDfoz8O8TkmP0V46XcT5m8tWsqRu/URDz6MU/3nGQgBouTWfz+1OqBQRe6
+oRrQwiup2l2+xLFIgBG0/L7I0WoRyGZXWvM62DTEziaGdS4+gx+wnLo5rH+T28C
MzlIwX3/fo9fxp0Et4Gl9RY8a/dWTayyTuhG40Qk69Mq/YU3Twl+HdsZmVxF0DVI
UFUXsIBLWWCpMCqteoaySP9OBEgTzz5jK7Pz8NfSrq/QlbMJ+Bqd7l4CQr//Bk/5
dx1j7WnNwGnVBChY15SClYWsly9NqZY3IX3Sd1Vh88DhFheHGRtZ1TTifN68Gv2m
LEoiOYasiP3xfI+P58TtNyW8UBJJ0C9hWma4xn7yv6ezG6geCBy9z0VzXoJ1aSAo
hACEu2RVvHdsc4MloYrSqXZ51RQ5GRLASRM2fnRpOVC6WfPA8TXBkSMz/b6csjlj
Wfusjb1uDzkklORrRTO4kxCZrettKc4/0WxR7jXIcu6SdkACvF7l7wS1SRRU9YQU
r0zMzE34NvsStVxUmDlj9q29eBVBncvRkWwbR0dhk0iTMer682pw3K8uwIuxwIFO
MQokyDJVWlCjx79lFAX0bLqCqgTFw+lEykddQ9vnOVqzXxTFRvwMeP1gFVojjLDb
bJTtqf185+MB/Lirm5ZiznXB9ole6o2RcTgfv9cXOEPXg3+evC4TeYNSSkAF/l7L
v+YABLXKYO3pynLxJKAJxD2+JP7qfXNZkXYBhEKdXU/5jeRIzs+ydk9ZD3KK1Gct
K/mqaUMyipOFaanZpWTHg1w+p+sXJ6ghgK2dUnRVh8SIkbjVBvcnmwOKUiY2AxA+
cmRYBYJ6YQMwMkCUYjbCaPkIaL1SsrWx2z8odv3iBChmI9nflJyddIYkWVu/n8Lp
HD54l/dWhoADJimy29K9vIrNrmcUPOrb4K4650eMEaXgCwOwunm80l+54AwM/UiR
85ZZV9aMWnfkizD2Iqx35lfelwOkXe1YFNin9WXTyrh1ZqPA17vEeMleTpfOOyyr
kkZkKA4crYbLHJdIBEcRDvxjnhWk3RXWVrUzB7JsUy4BxzDRmEpO5HnfikZQMkbz
76NIALu3UnBRNfIdhFnZoR+6uA/IWh0xgBT7B80+VszwBaogytGjCzgD6v0/qSI+
HNnq4Q8mEun3wkxmWh6U51hHyYSRmiuGkElngWvSY0EmAE8Y024vtqPjTm9OcX8h
Q+Wy7FYEEd2gWgilIWAsEIKWRarTTc/1mnq7/eEJM1SyFk5/99N+ij/Fek5TUm3h
IGH4sQe2XMRY4mMtJKvB43pbTmgGPcXMeFgLN8ICtV5DxM9DUUbxCRP6+5FaprkX
UVjIt9GnsJTi75gZo05yewiz9EfvWJaavslvm7L/4Mk5WZUOEx89Ouuly4xQRbmW
Eub8baSWK40vkswjjavwK+LAvvf9T2TlLhBEPLng497Cl1zNE6Hpd66R/P7CGX6j
4CgrsWVK8FSwEs/tAIrBQYdDSmvqP7KwRC3I+kX+HZ7K0UrA3dGG/vfgR6MX0Z5g
Qo62QE+GySZ/7wFMHzVu6Z/vU40brNYI67R3gibrLSopjyt4s6Zw2v2Rg+A8oePn
yCySqOZWZngp+zXeUlWSuFr74py8IIE0Cle0Kndtp9ImbaBix9VSdwC3RI0iIcTk
CbNemxJoPD4TuKv/rTczP7rrRmNALmppdyT0Y0bWs9HGCWmYkm+k93hu4mQozA+i
vmlVSuP0Ubf3hwQ1Gtwd56Iebu+NrUwV04CgPaD3e/pZaZwPz7Xc9S0TOj37sxho
mSNma4jQ3qORRRsJHPSHL/3rhHoVf0HWHUsnEWt2HGlWIs9giVwpzYcDgv83ZU/E
uAuTkRYi6g4eICkZtD6MkQRoOYEMccPz0PyrFjJHTcXG8ZlSzK1YK5pZEwD2PGaI
M/HytSlAAZQZdKoqvBrKqc3A0LmpNfsYHPqZKEieWxysZvgWAcliQ4s1YZ2rAMXj
ewYHojOPkNuGBEk89RoGbu1pP/7CbB1CivaMnniWNWUKMdQ6I3vSBl+rkzWn9Gd/
aJVKQy2A2ozYoZT/7uh4sTX5G53/HRTQLmXGplUays2dITKupFja1Sq2xCeEUhc+
e8F3UnFYQhgd9Q2eZpnwkVcYxiOBctUqeDNW7x9m2hWvcLeZC9FaiCKyXEAe3Brg
FQrim0A4Ia9T6gKJctTr1W5hmzWLJ+bb10l2S9noCoXzpk0ItkoZg2qAHCzPg1PB
/qjl/YaoHSym4VexcefcDWzm91XbRRbcxLd1aTeZkDaJjUBYhggrZ/7UiMzV1fvg
tYJv9wOJfBFiydVh/eJFEAdXcoqlP4rxeNw7tgHw3qcJwMLd78lKrCy5XQZRxi8V
ULbIVPDKzaiJg8wXqQPElTprfqdmVoIAlLUBVhgfCqE8UIqi+pyfvVhpnHryDcDI
9mvOQdcaIaT5i2gAAC4neewBgz8oDQJpCc8gpfkxIjNMJuN8TBmdA4jAznz/iidO
+1vjnJnBNZI45fKuEs0hAC7y3j465dWkY4uT8qNFnHTOJ8b/RdB2NIVlKKekKTXk
afmla+HWYGZkHete8QL41XPMBGptp3EbJGbvzvFb9PwkwfE+kyNzZ1aEHPGSIM0d
ezMVFYzUEi4NPcbPBm18ON2vo1ZD/SnnzO7lSXFixsVtsN0/xbpLrb7Ep0i2+b10
q6RUpMYKRaIyrlJeXwcSY1fooBeiw8/tqV7NrDc/Uvw9Sicaoc/EIdLb0rY582hd
5ADxmQxYO3iA6H0N+DWEuNXWYrNfDe0PUw4idbgUpaMQb2iKtvYUQxGG0JM8gjry
x+s8IFLWVQtQI3Y77pu1FDLcD7ERDwIuCzDBJocrbEyr10pBJuhdg3TUCzTkGQT4
KuR/XTwr2Ppf3XzIf2ne3fhV7wmWFtOd0mPAa34vyX6qNMexT5lpO8WjEqvPMTB0
3wq/tNufr+omuhbjDwHrrc8++rpYw9Tx0JaJ0w/HKzfUBco3H0dmbxeVClNaSXA6
5/E3LG/V7T+wYj5CA6DtBK/EmmyOkX6cjoXsGxxjLMqLX/XOy1MnSAG5+nTNEr+6
OR3GRL9HVndSPBZZXhlvlMCbZ5viI3AJIQp0ONHNyz9SYQH0aUuG8tpoKZdfbRLM
VzGU1TQc3CgV2h0UjT/hitPQQNMfFUcG3OvRpxsJ7PqN9TXNDTAd6rGAfwnDOyTw
RiOF2OFUWzgCNfefFF+AOkSO/yw2k8bylm69n+aw+4HRpYUTATgsE+01mTWjBBSF
B/wXej1nXetbmNCeJsqeoTMaiGBrcOw8d8rPRp1Y4ooJxVH665bb5wjjOY4xPQJG
okdMwCL4rbXvryI2jWhRZwoF70RxGryYlL39b7uRRWQ4Jmu0UCwa0UCWlsQ2HgSy
ivAJMUn7Fq/dpxhL+17trt8sbZtBawBt5r8s5GudLtMMtXW89gTRjN8eSahAVMFD
RYUzDj41pkdcxbr11cniwG8cMxMqLGPSCtWdQ2TCCdBR8QKnQ4bZAgUwzQE6DMVu
ZI3U7THcy9/pObMNPj5Le6lo0Via2vPXh3l+Bnabs9a25VvMPee+wPKDXviomFz0
0MKUWnddz687HHdeO4ib4kFgMyjEMLcK+3EAa7DkWDna8L2rUYmySFkEZRfH3rld
H3ZtOUszWEKypCPE4q27D082xcruZXb9/iokkNpIrWHx/XXj5Ob1DyTQfwowB+rR
yuDFGozm8k/9ZgbFuQ/um+2HAUqiv0mbnQ2Zr7Kio2KSDQ7bmndlVXyG5Zsf59uc
37/HRyOKTvQNDpTxnmVSReEzPexoz8N+/5afgUcyIm6HgVAKdWf5viB/qjE7lrGb
Cot1CTwtJ3lE1I/ELUQCZYaQ128LYIc7DAo+D6QyWVzzHVxXjcJesJbi7hk/bacZ
+XbkUWVme2xeAuNr/mqM2PFY38xhTwLYu4hSDVQsAprm/h9h5uWIFqJrqBzb0JzV
6LVQTAeR+tk9gJG8UpINq5ItbtAWyHeMSsiDtmCeQg9J1Ht19RhXNqrkzwZW8aqh
FIgV3qDMdqTv20aGN7yGmNewseiQxPSvgmG9JtF8q6VxA7y90OHw3Ez2hMNkVfAB
YOBdpZyeZAWIMAfzZdmDuptsvdG5pnv2QS7v8wOSc9mXYBMoXbaBGDFnY20+ap4l
+wCUjEsWfO/0UTgRNUuDStUP4c9ftww7wnQYanRjXzJCLELkKr6xPRkfXQCzsoD5
S48G384yIBNAjWyHQEIjWGRqO0Y3SpGeAt1Yv2KpBvIhTVkCPJk0ALhana7ECv+6
2KVNOH0htUnnQVUF3RirAkpFZRhTyUqVKXH7241gA/RZJuWIK7lfBdx3nmNHslbm
4RzQUVmeDxinahsTk4se/QvekafoPo1S75EZBNhL6qmGvQ3tsyAaVkJ0ETw/RsjV
/ZfATEyXEepnWJpgsM13wX+5Jde8m3sE8ORSapQv1gtElLbxiPYfmqGIUNnxsbhZ
AHUZSMj/WeJ4vxJ64tYD61skjnbPcAiI2YQRzSEkbz18BZQe+AnTq+X1qrb+cGty
akn0wiGuMWFS9YqUoBlcABMuQLK+ImSqQpBh2bxh0MtPYjr9B59iFJ+JqBxzGeAF
d3kCwFGA20vcqffP6exoc0L6IbmRtOzcPzGTTWFVhc7OeqN8yGsWpNzy/FWJOXW4
h4TMjq4eZTLCiKwdDkAVUuG3jHucHfuJJg+ptaYqWzhQE8fFqPmrdKkfQm/JQ77O
DGJb6qKH6ulJEUEl9UCcMGDcHoEUcswQwAcrzVpN2CstLcRlL0gV8QrzykKdGxFE
bklXvC4/7rl3vOmXnUejcHQN6aAALIdkpFqVeKahcCdNdFZ4xVPL/XlU64o2nyyx
FbMd2WWgatxDPFon9JQaJx3MDznW5Ev5W3oD6dlXRtrbv9/saKZokmn6FmQiuHCG
OX2j6T00cgG1onxM5Ou8nw2RIOpWJBLo2II04xeVUs0W9lkDNubt2l4ugUjljchn
W38ysMM1PasDSbV/1m3WYo/vdrjn3caPzVDpsI1Ytl4AqIOEsT2q9WXqdJxqaR5P
WFIHu1HrYWWdEtXQfDnUCd7hZcWZ8qErT9T051egC6PKtIe6DnO6vfDc6+Cq6bH5
RY7UwQ7wSsislwTkOmwmSpwLoil86LGyHwxQan+WbTKp+38CSI5BTsla5xNGBWxv
eUw9Zfa7Q5N8EsntUjNtT5BHnGAPQnMYWkocN0C9ejs7KIl/RUvJ76G9StKoHlgO
Ru4EjP/fGPgj+Ny/E0RI9UodYjlTsaHGsNjHvji0D+xUvDK5+s/vZ5vI4j3iYC83
Dpc4BiTbohQ2evMT+XXIZl5KLqcTvPVaM0h+JwZrraoxXRL79NZyOwUY7Sw8CefF
43eQb+6qoJI5Q0r1SAycoJMkVyD9tVAW1DzOF1POyG3WRteDLNdlkIFJxSGeIyIg
TAIsxpX7IRwVhAdKiEHRg18BULgOgBYxy30b7AjkvqKVJ2SuZZDVhK5f7MnHZ5n1
IGp8bfPTQgwshr7SWUm+j24eEjjZKoY5woOYnI9WLEgLj11DcCgRv+ZwoghmfrXF
fL7FWDYmfPoksXH0j3VJNy7WoFrtuVB+ggRDq0G46yhppxlEunbKtKowVaThY1LV
1/tnIPmA10lgijCC9RYX4TICwuhyvZjOPf7tfetISrGAwR6C5MLWjsqsJA/70/IJ
oaCoSVHe3lyai6IItfTlRfpX0eTmoV+sbMVXCpcE1doNcBuCjqUA5kzVb5IpJ/w3
jMCtnQE54MyBBaTYuFSFtGlSsxdNmfZ4tGOt81osTPkFLeWR2RZ/ik5N56mojAxz
wk4Osz7cIleUZDEAjBQO+jhh9LtYrXnxxprOkxSuVAXqylK+RbkrrYDdv5eSIwcU
YV0Zf4dHGyArCuJpnBtj/ct1lyxzw+swEeupwW5wf3jAV+IrkSAMuuj8tKMCd/vt
ziJ9ifDkq5X62MQJlIlr679aO9CZi6VxxTF1/CtSG6kFWaU/JqrTd9RPBYY8/v1c
y6Dr4dcrL1ge1OZs15RvI5hVg1l4sCiI20HizqRqhF5YIKlbGdtEDals5R0tlZUd
a6MX/LcLZ7CdheW++J65XEPpHH9por8vvNuW5U+b5fl5Yj8r24Jgjk4y7sjYxX/K
QrOe1pvR5yWIpXiNCoHlR/RqoWTGf2I9ht1zonvgYOgzIPTjF7Bd9lftcYOYArUa
GVdq6EkBNuK+RmJdmKttdsK1pP7YiD+0O5zeBKEZ9EQoV67y0IhMEjgL9Vj+jubI
XfY7M8QFCL3ZpyXkmBnMtzvHGnIghx5MX3jHOREI5SKXQ7OM09tWrKFdc5E9TW/y
XMvO4htRvinnp+Kf2tCmEyj5ku8WCmueSMWhKgYsu/xn83VdSCzl1N4i8T6h1h3D
vKJfts3BZenOoFiYOW9ktFIG79k13zT37ozn4V6eUkBap53OxWIJuFBU0uzwr2dl
SsJ5ZSw1UJJkWk8StLUGxzM9N6dF1ddU/lQe8h/S1Cy4tXfJp1rCB3LborCULCVe
rP3hrVuxIMTXYce+T89hLNIX9U0BP6N9L15DZzLoiyXP926A6O5c6nwAznSwSvbo
YmX/F4Xe98ieXdbfglPx+pHbMb6kAQl6LEEdXQnG5ptNkUOkrHkTZKYUD2GYo/Zm
JPg43ZHnr2BsI01Ckf+9xxSVTalF3lXy9Gyg+hG8ZaXIjZREl/K1DNsYIFOAF1x7
mTcnPNxgeZwVx4IsGdtdN+CmU/E9aXQNA9R2oRyT+1VFC0D9wO62f4Y1CZAIuoFq
DvBnz/Bm54TZN/i/AE3znawURECX/mFBrQphSKpJ7vwxqARV8fmAMBkShpyJWjzy
NLzFhub20yxgy9JQ6aO8Za2GFkXLVYM0hZMXhf9jT/e5BAeI06xr7zRma3FHq1Gn
E+sTNLwlkpsrrGlQSl3dj/f4NsT1nEXE7XHUERL8EzstZSj7nIH/OE8tZTDStOxc
C6krO3xTe1a9UMctVypAXqIbmDVa1/a/5SW1UUwvSZBWaXSccnqwiO943VFRdyBk
VPzoRC1RppbJQ3VH9bSheDJ1ElXMzyjPaCDUVE+J4dGD9MYJpZwuELr4mo6arCty
COHyXs9/kGRRQqwKEL2P5tXFVy3Awl+rH2jVXoioYf13ic89GxPN0ck9pPE/olHm
N58hG1Djb8xUJCBUrh8r6l5Dg6lbg4nF8yC+mMm/qgrDjRtTLcpLvJjC5wObL+vW
M5XaxcbST6B3XABkdaQ9xTFDFaIBe8XhNq8cZAeq39QqE6HN0ZXWpG4H4VaIZAKU
j3CGLzCFImuXvW6+hUz9IPcWCa+Rxn+KMgiFKkxDT+NhgTzOrXRzMP2Yj4oqh/L4
DZHCdAZPw/9Oi4gf4ESkJ7IKIVdTB06PT5GQOgeTWxydDkSQExQFP2we6DDuo060
uGWmd/XOwRFwAeg+IRpzAZxcX3CbfJdkONwkVCr0kig0qQGTHt013iXDSstXh1O3
e8W+apZVAicaovMF6KNJnswz5lBxg6PymK0F4dD4QYBv0KFzeIigAjuskPo5v6NO
A2p9jY30uzzUtEKUpxnRufnCvsOF7dD7tExc7T9gX2aynkhgSk6vluEGjaTs4FkT
TdnrgMl0+OAw6tZY/5hYt9l7qNJ8OPX8X4oO18lf4RKRa1ft3Nkfb4xg6OWVmOyI
BD2/BAgTrpdo9bBQneGT8CMUylRBfwJPlb6g5lESod8P7B6/ejGTxNI0+zfcw+CY
ToRLKgxmj6thm5kY5BYEUHN8qPYPeVO149AV58kQe4ng33DFt2ZQcwNpYrUjqQx6
AdXutzI7UQfKujdLLMnvb15Z1FvJpylfyE6CMbyUixc4RWSOah4ralHvyeajxvQ6
2n9dFdksEKSYDG22muMF2tRBI/GdY45iKr5mWOYqoub12FM3XF2bApLvoAlDIxcx
dfuYGzLL/AP+3BmipmtsX4dGcMwHDGIJ5vsjDMN/e8I4nZPeXahF00yzQNbPJfDG
XKQ9usFN+gaX+25jQvk79c4yetGXs5M5SrWzoUbGj8xNhRUbdqyA16krj8Jy9e9s
KU3UDprc0G89IKJD1fwxSyDC7nOIlNfPuBU2cHCrXbWd1GLgI9lSxJH307Wa8mKe
klgKN09FQPU3wLmqPzpGqnFpvhh6EH/Y8P6KafoPkJ5ngovrOGEkFDURCUCN8ekV
90tqPSZghKKRX455421Tn42j+ccxPVge0oe9moJVKJ4emcjxCitRxVVnaK1g6L1R
6aJIuZjBx5Lcg4lksNum2sp9peEhI/XzMyjZboKptfGDlWs+bHNORzceNEoihTMP
TbVRvKZ3iHm2DzawPEptwcBQHxUUIjUnksab6CeupULxJkh7ZAglnXt0pa5irMBG
7oNkBKzEaZHOQ6/nNrmEEwu0OL8VnfbJeZ6yxl4fo6sTkEk+rxBEO63IPhOlnaYF
asmXf6L07s1iJFaoixOxKtqMequkhGTFK30XUiHAtMqzwZnV37eY6F29JRWoPskl
uyq8d4RBRP8WPNChWRdjAvUfYkFgqObTl4AuceKOz/GOKKBJ+2b0yJ5b0jdWC1he
Hn+PLkOZlBOQ3qrpycb9cpz/h9t8lJ7poG2Ha+/Ue89Q2JqF5sxjaUwGEDujy11z
ja8v/sFXdCP8qeq9DSaSuiGaT5wSbbVbQ7gNQSDeh9DVv7Y9ngpnnkSlR957okcr
KWVeezRr8RM1ymzsX/bkmsHmnMqMWYEe8IBT/Qa43ic32Z9/W0MEwcUicP02pEyn
lS5qXG5ew4Y3YZHRUdQUKysrrrMFWhTEHCFXcXNujJCiSAtFPzqZ+5+lN8JytI0G
Ie8FXMJvab107GIeOi2mk2kVL+7WG3+/JI0piBfCFGIYq4ZZOugKvABu2B4uxCJl
06PnJIaSWudw2hTYPsEx5CR7KSAc+su9CIePltPQVktHwEhJGjB3Pv6hM/nvcSdx
pj4JDd6dh6vRPBKTcwReRENWOf8mru8GH9t5AHAMA2y+ux2FvcMjGbGrDUcIs1Bl
DWpdTCOK67/xb/hAGBmqhX40yUFGds9xVvSkL0DHT9bd0FpiLjOEnqy2WbWO5vLp
xJ+xx8lS5JbLBxfik2QNAarSaCcsqn0GolRYFb1pRC6+Gz8wQkGbsOQHExfmvI5R
lWNikdhzi/nb4zD4TsNxX9Wl/YpZ4rG9GVIoMuJk2EIMnahl7cbuJpTWfEro8+pa
Q5qsXZFN9GCRwS8p4eldzIgYztynKSD7bZVSP75Bm0aN9CoCB1frdPmGNuc1mtSR
FC9bxCq9vzpXu/A/i7Zth+AHY1tmwQlsPh/dVV3FanvWHdeG/eBBsEo1Co/8GcEg
9FuYDnAp37IJxu3/k1sH945hdgcMWcyuyQNhIOM2SjMsBGfl8J1yPFqmA0akis06
ZfBoLtZ4upOIUM6H0mgIW4TbmXKVT3YIFV32vH0swoT1h5GAemWfpjprJY14MPb7
pttT35vYE0XDHo0Fj9Ooj17ZNHg5LHfjJAkAGMPzCgTq8lNVsimnvmjz1lll1lQe
eM0S1thHgKaMy2Ub98IfC/+kOkLJKpzImTI394aFfKzWY/gDAOzyc7Uk8Sxz8WHX
a8reXucPzP3yrZWEHn5Pnrm3ERiu25dA8fA/C7YiVxHlHSUkvG1c+w5ebhmc//4+
E0d+NHrTYYsSDtKD2DZhKrDCW4VbGYgVD3go/ZRxS3Ce5h+4a7RIGogXhm0raWcm
pvtOm4kLqJ6We5kubXrdJkZSGcwGMyevB23A5C3e1BHrAVzDV/mPHcMzBDNZrKQw
56fH4DpOvWkp9nkJhDDZKEZlABueJDCV+yYy7hpqLQTnQLBDw7ual19eHZQKzP3M
hgIyyRBVQ5VmlAaob86MY6xmBtskdpWzzoQg1WsBNFjqaKAf/gobNx0m7cJYsCUu
T4b2DdJZ5wqpPAH0gJjdA5Aj3W1ZYOPA9t5OotA79p+3NN6aeVG1bCk6h2eJitQR
YfMHC4gxZ16z1aEaLV7oCNasMNWUOhBfafRS1wjv1/um+N75yIBpuubrnxxOvC6u
EGNAPJQS+dw8wOQAmZb+x6gm+btyN51gnnz1ldtw824HB5g5jm9Eplzldy/7fzYy
HTVmwZgaIhsNg3Ymc2IL7UhX7FTopvlSPs9sjMNbQ/kvOCk4z/qLE3RfuuNTvZQG
oG7jptkcVIWtRpk8fAd9Wt9p7t5oDfh37tmOmyV2VoyWbV9WVobM2icuOUnG8Ykq
ku7vmy08vqgLQKxwtCPHCvvh45ahNU62Wh0vuLLaN5Qe9gpRbihu95PgNyzEbQnc
sfz5wdTFZHLveAeSHToiQ4GZozubSizuViiUQNhg7m4qrTF2iDLkpY6G9mvXM4rF
+nVKWs70BfEPI9armB0SJICvLpU4KUKkz+zlySzjSvnES55ce5JPWdv/EehGLvq5
tqy4rgsFeEcKhyxOETnikdE/HgivJr90b+6ym3lgMQBhLyLDYl4FotzCeQmDln7W
ijVGvJ0I5TIESBhC5v3u7xwghixC+rN2tIPfGD8ISoXOd5NEE2dmaI1k2k+D275O
Uq5wcHfk+GfMng5/we6V13o8V3tsuQnp/mHEeEOzDK8U72XbReknclFibgpE8clB
N06wALS8/HDTIa6zOiDTesGlRCMni5aT46G8KO4z5712DzHoS5hnqGmLehyYCFxY
FLmfcAbhFUlARZlOWx6wS4F+/y7tSGnxALZ3hmrjPHTIyKJaxA+NH0Hcz/rxNLKN
atyH/rbqikW/9NmNgRQGUNr7UVz++EWaCSf1gAOxqZntepOyEYgdVNe32dJGXMLg
wFFh16vXOSZD5Y2Poavv9dTQe8sstQFc9Uzlqvz+aJ+Vl0+auHgPDd7rL0MZaePd
05vCKezw/n7xzQtd5Pg3CDDtC7v4NKj1zGoyEIRlOrl4xgsFWYYrlI0qT1zgkzGd
I1W/CAyy0NgsaJrY4QmdWVCTMO5ds+Lc6iBfxBA7LHijXEUJerlYzzoqz1LDLcjG
19yYT69usDrzDm4G4iJAK86BW/sTvtGsws2hahBSwwue35Xvq0jrRf12L5fhe5OQ
tPoylJppqaYME2DTR8YjOEvyOLNpmm8cUOcpcPRO/gO8XG15S/BbLQrZYyEOQLHQ
PJM6MEmTOeYeQSpGSC9+0bq/9PAnrQbjL2e9JNI5g6j/pP28EJkUI4GoB1zhXGmS
XkmfqEjjVO/g9O88E26wdkK4QFKWufmkLUlDLKT5XDkmZy4j61Ze0zMu+B1v2crg
tIppAuWrJbV/l5ypsuGtTOWZH9Fb9b8QarBRc+OpOE4sC/9ej1+QJ5qBXnXTSKyb
zYomGbYKam/gu56pGb1oJc3QI4lkNu5wf5ph/zlMOsUcOybDUGPKM4zkhmzim8F7
hgLYc0IRCkzmBaweFGNRzOUN6ld/kBY8yslz1t8v9fNxskFxK96B1Kqi8KPqx0N2
ZGi7FpY5HQ9n1jM8uy6a5wz4nORL3MhecwrflK3ULUic12CF5dApmasmtBMderSA
TvYs0AUDW/qXamxU1LwdHZeZj0q3oOri8XX5DLnqdFthGsSG0XPODWFUI2J3YAPv
dFT1BoEOd2vAZ9R2kHeXn2zygt3bfF/EjBRB6TtsLIBg+3ioS02qW1bH4baQUvYc
HVNq6sSgr4TT7pmQ4zNsaR7+U0nUSPnQUG+1JAIEdXBnuWAnsOyhSy6BTgyjnTv+
4AabdyvCuTLxd+A9YpjfzvIYilFr/2/UPcxxiQdUr83iCheeF90pI0gTFq3R5Akc
hK0Ic/53N7uEFvs2GM6LOzVNONFw8ZrJ2UFiCvyfRHr/s1C2K6C/iY2Wx/r5Odzg
xzeEeStmMouBobBJ/9T28FujJ76mkSYjOKdS7nOQPKWP+UbfxuPh12k3w1vfVly3
bEwPFzJqHdFEBSfCyqzUcRLx0CAoO71ai0nQlQ896HXYqAlKJyYqGyseXvRvIcyC
x6uOoWve5tMmuhGAaK/MH9mAJPHh09rB+k1/SK2Y6s/w855UNk+9ko/QRwv2DUzb
ESj1QHmxx/r44O458CZ5EexNBlIoTdtNTRSh21kQbDCubj8Kicb9w9A2pMhqv8fU
Gp+E4r4XotISboQLTuenutk4RrgIN7AKyYLr9kvSssCs9Rppo1yXtCltocgxQ6Nn
5psEdoeBadEVG0t29J24UFEPBLHF3GvrmYI/UNuTaB7gfX+w7jsJEokrSWgaHIEi
gx0al5ibEyOaYqktGshP5ub7aOVt0iZtdC8pgeotii5HaGQYBTvnKaDkNPDIZPGt
hlXXr/at0tlNKYQ2BWYsmE2kCwYFqNIyxpAil6c84LABGLdS6WJEggmftYdYfN9u
nA9DJnzww8s83/00eR4DPD0upkK102EixCvJRNoflHqQ8htqi0QQkFIgUN3BSGVF
Zgt/5C1ylO62cSF/xhpoM0g6K2Cy7GoPwFbdMKM0vUcgOSbKf+zTOiGmd0j5WWQK
EeJsUfM6Vee5UF9vGXHQBL1nVQ8qmdQxZ4G+tdAg28xBjOwRpkq2HvsqTZtpbwhb
KtVXAHy/ThgTQDBqaY/WEJYWzxcS5PPyOuUAA4n3uvSISqpwU4DkcEnbTGqmUFxu
+8MTElVRjYflhHZ/FY4YN79O2jntjrf5wZdfM91XFHt4BHn5PSrvfHj2LfLhvzPM
VBkbwvEyWxPr3u1MaoudcA6DF06zb/7FsePFsSMqXFg9a4Cl0zxQqd/psjSxtcDM
LO727iCR3IWUo+NQAIxrk/2Y3pAk2HA6YYNN0mrYzyzScmm8ml7fR+qK7LcH48fH
ju3l8EQqkGi82T6VUsMSY8f8cZCimRjS62FLfP4EwoRce9tTYXyBiwB9v3/0ODzz
EMyC9oj/6hroaC65sOYPlkIAWSK4+YOD31uGumWCIUMrGXx/qEIi6jRnNnMnq+U5
rzJdnh3M4SBD5tKf+D+QmhGweIadenhybdGGa9E726D4I5etV8V2Y1c+2IhotwGS
0LL17JiBI+646fj//KZtG+/AYknjFq8KW38RHu7zrq1i/VzDZkb3BIedesuIoBWp
XwvQg6o2KWOD/QLUkqRIxcEXAwJXgqWe4aiaD2wi2DI3tHzyQrnrp/k2ejMPXYtC
TzvAbAR7S0OcnbGGmLsumvOR5ARC5EPQM4QJJtZ4JbZ+njuSolzfd2tG6fPZjNt5
9HOd6Jdr8jUC4g6ON4MmgKqFrYi0SBAPwqhR+3BF8ZXQeIljmD0cqi72qdZF/tgY
ycoFMbWfZTdia52HXsvy45vqD9RmOKikuURzYHzphcvyecTPZDcQXkn0a+dsjcov
P6FPz5KermLt2dKxG1ms3TUXB/xxs2pdoIMPv3YyqS/fMlI2jaOazJ5zmhccasVm
Xl/NWhIowDxPpiDtw9xwWvnHq7htAgyTQ4uLOwCC/Lxmi7alJaPDz0dA91TvurM+
y1M16sGajCuZmT3aeJ7Kguod5N97Q2elFYfooR21DEVXmqzUmzEa3lcl7NJsUs/3
/D3ml7CIqV4BS5ACF9JgF2z45y5X+omKPUP5OB4jnxwPYxnn8ur9D0n4Reg6wq4e
gGfmBxE9SWNYWbb9ymFjfmnScCarzeVXRsQ8UVPNtGOHfDfdOg7WaNrsEHrjY44t
Jdhg+L4DesfjoxnVAre1P0ziNUFAm9NWVuBLicnFRXhrzWDeURwCAUR5IdZdBGru
9C8juW+h5sP/VFWb1eZ5nqiKIRv9j8ikjkJGIER6a9zAX41XuQfp62ReKI9IghR3
6WJrOj7F91wo7fBRSJxwHhZSoPpRwsxeQbaNVXIti+VpaR/YCgufxaA2DvuqwE2G
9xJsslQy2mNfnei2ij4+ChRuARQz8U1AbIOY17oMT4DpsM97dIKHgdNQXedwOPCD
cCZVL3afROM929i+9rDnE8j30I3Gc8BIhfcbnHZ2qU51AD0XN3wkbdXwR/or68MY
M8P03QsTMiKVjRuj7PZ+NUtlxqSloe2J5FIKteu8e25d+ZKb1F9KvRu0L/0k/ju9
wi5jqCBJgwAdAlYs0gYg0aj3/CVCZl7ZjDPZUbQRqh0BBpn3T6FUZ21gJv8C1JvL
t6h3G2GEq9RCjbbzFyyZ4JA0TMFNdYyg6f8h+A0ztxcMoAAcqALQNhN6/k26EsBz
7kdRtFp6s7b/8glIflz3ZMrbzRN8W/mh7JbyNIf7P1E7iLhlyE7UbCU197mMjJBO
5Tm6d27EodYMkbwiGA6d4iW2Znu3OJ3UWR0bA0i/4GaB2HN0spfw1SSkZ52cIf0P
5DBEqLNHHQEopq8rhRyfqSfxr64t9vN7+UgTwARJfhhRE6ms5xKk1F/3Xp6K3/78
UxLS0Ipa+C/hRfD8UkVgs4Yde0Ck9meRd6zYjv5h4ZTzEqWEPobdqdfAkEWmK69w
zu3O7GhElLVdyhIKu2U76q56KgxQc+s3eEmxJE05cPxsfJQPgHRGAjmJyq5HI1Lp
hNfTxyyp0T1M7PMVpP3OvKZfDyXx1Eb9pBYFnUVqcZZ2ge9YkDXxX3k8Nn+pHf7m
ApBm8vMt71TSP0mNJuQCodBU9V3iPhzydC77fFZKaeJFWUHMhq6yv0gCYrRvM15U
nYcKzqt8kDp4GV79NPABTECURR9l3xZHyko92h8Wuj06ruojs0SIEUxAj/z9AEWO
Mw+EWQBv4wHj2NnjE6D0niiKlrINCYP/XQSPJjkSBpXwkMIIoQlSFR3PFnli+tZ1
P/9aaaSAtgBuz50QfKeqoiD65QFCqzFkdsZZlt4uayioyzM/nFdejYtNC1k6OvmT
wcjgZliJcOmULBGayUmT5WAusa3pVRwxar5vhaZYWoZE6Y+Qco7zSpY8zUr+D8i3
Bbbhbo9AGABRjFBjnOqCezh8+pLivSMwWqH9SVYwSeCc/UcXSobBroC5oxKEBftY
tudfkrgQox7xW9uc6/o0JJJE8a47I/fiENn25BqNJh/ofDhZnUAoqGGdIlHm5Ws2
9XCfiaf6b1zmHxSPDrDe+irmL0gC5+8jlnUJiW8cYi6U5HZ7nTRc3PlFZdkx1NjY
AVWy5lzaFabmrMSNsSE+653NybCVMRLQUOsMsAH/TLsHHEeKaNqVeiBw2Zr2QoEQ
bTIklYHzmdPtu23DPKN9vVhsdJBzjly07gnmZx+KhhDjESmrkVudwVxqLOwtvhAR
zn6c1nyrNTXkZRBhA8/G0zFq4htoFPv0nwSKY9tYt7SzXOKXXZITA8d4LrdBteK9
vurSrRjrjcbI6xkv6BmQnhs3R0KnC0gL3SGxk6Ep675OwgRKiahPLIFTzKXO+kPv
UWmkUs4MWQjErMnPqH4ffw57ibR8gnpcZcmcHBvGTKZjAEypBHoA0STTIcW6Qvxn
iLpGNP2egs045+bCRQjEY1xjFmc2joDnY//r/7EaqnS97v4iff5ZT8zGbJXtuMQr
dwSr7Yt2me2huanqtkCv5nbxBgz3zNH+uLVlMPf06PGmk87mpeXo638ym63Lo44u
q90rDw4gBJoUL3OY3Nqe2PpBM4V4mxlc8/tEs9YAScFSs0E4txcilvDt7/fwQPSP
F87FuPfJ1z9lsaQxp6M19FH6sEQjjDgBmAd7e8xI7/FUjkOV/vgI9IQDzIprGDWN
Xa8S+R144Ojj2aX0GbiQMgaRMOoMGFia4JSXkQoIaW7f2hn19ChTtk7FvKK3ICtQ
VQAzQnGYpNhFvj4kj3CELiXPR22wOIV12ut0YrqTflT7xIoP4UH/Cn3OPum0Rpsn
QPqHmLAfaWvp8t3kzuFfTEbFIlqE2byj45QIZOMooOmfxQRsOzeI1MwdFTM8DASL
wdx6VdWyqxJoWqXpdwOvrtskK++kUrCcjfpLm64Ji85lkakebT5iQVAXtHW9GvtH
ZNSCv7lFsGfq3GuhmhGB4XfWOwKQ7KwzgUzTkCDf14RN0X/hk9gqm+Q/FrXbvFv0
WJweEf/AqkJUjOI0sLSUaxIQrttFP/quKf3Qb1huxJZtTIGrmboQ6Fs7dYBxaMhx
lDI9q6lPFhTNP9UQOPLZFa6xMkmNUwMDdGUrxNPqIlGAFTAn7s6fJLBeNRQ9qeQv
FoA/0tRSFrMdksHOPc/zT6Qv47mqKJkpphaQICJjivP9jNfkGnLtQH1ld5DTxIHw
DM8qPYmmyNsFtw3xBwIidS3Hgzxi+aFYyGVShv3CaZpWkHc0vrFx+2r8vzMJK/gJ
nUedejCqqzRWy3nHT4flBreuL362iJsYEGqRsSkYpoPDgo0tz27dqJfh+SskQcZs
gT9wakcX5vDG+KlKMlC0NoMRaIRNOlxoKFRmIBNoGL/+5FUc0yzl1UUPZ/QJFcx3
PyR/6dTJrDtQmUteSW4cL2sTPxxQXIiyQ5gZMP5WX44j2LIl3g93poh1hs/daM+4
UqBrGQ83cq6v5hp6aUvqGJLDK6Yx367xMSyKo5KGP0rna0EEdWWT/DODhYTCnxBa
UmMnlWIgE3UjaMu/umVAK/Efuyqq8JIjqG1aEt5j8najnmEwZoNX1+Y/c6rmmzgQ
u2V2vCAVlLmrCqM1NBww0dVs0WIAebvXs7/+ZOPM8hvMuZoGWmqsdJyU2t+nu2bj
xsOAfWwMH2Q369hQDQMQBr6wH/KNYYGz2NF+1ZTGDa3LdwbnKyxbRmlcb+0FFgJy
Wv6Ckw8u2bYVqfw1DUCtQ4SDL9+KZ6VQVGaEZs4lY6oV4ylG4YfuIIYF6ygiah6V
ng3KnGOY1l/K1qGbeC4Ia1nMlP5bn4AXWxWC5C+GNjsUVhIvp3izi9L2CUW/1GFg
hZJAlGLGUlffFSWbBLzO/Uq8f4ibrro/ZU43kwZQ6tmyZAw2yus80dhE42oQQKmd
v+u05AqUwVjZoZ8fO3GeUdebu8nXzl6n2JcQWpFylrpaE92SkCw8O1oUfydfGGHj
krTWt5sppf6NaZX5pRzYoAMK2Qf5yi7FZqWa58oSMP77whFvUuQDAvaS6+9UBdDg
nzbtNzHPUh3B8OXbAqWrgT/Vhb0tV9QS68kNUhhdgYkb9nxP8+E48HjFcENmsm5b
1Peky5sv26qR10cvigTLg4EUW8tsRvJ2wXB+un/QP52JRkTao4Jpy2Gp7ah+hXLt
BbcqlNpYzG2T8jmT8bNSRrgrKf96AOE1jELiGKPg029qKtI0+fg2yZbNrakHB3m2
dzb9UBNLtAPiMGq1uhzB79+7ESKxnW3OhSevxehGnITvo+o1puRksNkACLOCPQ4M
4IDiNE95w9kMjX0d2VF5jaMNP0SoUuwek9KkYUBY4GXaf6+991DJek6FvCFcQkIV
iBtv0CfIVrTO+xNbpX7f2X8aqMuwXVJxct7b2pQpgYZf/rEZdGqz04igo6sO8RLn
goautD7N0n5aoCjQRFMEYrFQo+QCzBF1bqnRiICB5RQcwly7Zs14c5W0WWuSArA2
yQYRM7wIOc0RZI11qcVv6t7pQthsWZR+IyzzZrCl07D3nivg9DOv6uGsXiBSGnq9
DITFk/bch9rqktYekSnzl4pvuBB7DhIRs2/q2rnDzUd8rfYyCVk/gKJk9vOsK7Th
maR95Jfg4DLflWZC3BNjJnCxYt9M50E7sk/sOJH1dXMOpw9EFFFD/12vS59x7/lB
H0zPGC34uEXwtPZ+taGUZ9jwrAwrXheuedKc26k4pzIQRLzXEE86o1qhD6oD1Lsv
gKqrSGM3iXFbkaUy/Z0hn+JiiqX7q9ogoxSjc6XwZ1m5lJvQa0tdm/LpK8tj8qsj
KED8AocxwIrsTisZczbc4d1EcIA4FfTA5xHsAU4/cxemAIsuv+z+fffyvqI6TgYQ
FJD9HRIfHkaiZqScZbi31RefkmGuR01KAOYLx/SnX1Up4Iwj9oVAeIG2qjJ0b6ua
45KwE5D1W+ohV5wq2vUTqOEOzipjZPVBFOEkvOlJeUC0xdce3h0gR56NpUICXvgj
Ngs76EQ5189NJRIK1XKBmO8dVgo9vQZKSq6V0Fr83hUo0IpXZJLn+vBPO3eHNr3L
Gko12j3xTCQhOcAz44djoDND0Adg0XfWX9WC7OOZhxkKbs5DhDj4HsnPe1idCukR
J1XByM/5CcbBZaAr/FFmpopBKc8QB2YIkVF0uM7zxFydCPVKxqI76PJ7pohJZc0B
EjO3nPqEHgDCgLjLtETOzb2D42eqTCi5/rREZhtAoPDAcYivMiuRG35uVv1Sv+D+
JMkiSj4mRThbaKL9Ym8qQFgvB72cK4FzUa3be6OZ4w5OttRCA5w6qdqPVy03Y7Pi
/oIMKPcb15GGvy6nAwES2ipf8f6phPll08UCSlb64JW+xhKei6AJLCpi0y7bYIQ3
fYftYC6Q61G2KgEpZYE703YiSZyZmYOSVmItr3DQ2rIEw7lAEvcOKIBaJUGbLu2N
2HUYSvK55CAFnS5DV4te4KvyXblwvD4gQLaS6O0jH3CRcBRtVQZuHV5uAolL//L4
bTtv+H9KbmR63S5xyf65A6dZIb0mucsd50gqNUwGpOO0Jt1aUl6FIDy/NqQyCnuF
bup3pL0iM9HRN+88ACOZvH2XyB7htA4JXoDBRm2JoO1eheE7nnna2E3p2Lu6NRrE
HWnmhsDep4oD1kV2rIUm50+ji92svm6m9WO5300XwjifBhxvRa59Hw+K/L7mY2oP
DDBclgHypZG4zqAODxxm/d15GWCBNMj5ZOD5IaI4bHyhswFctC/Y0wyP1CpuZ25K
dKxr35/rvB7+X+gK6IIstJiPAzJxuNfpGkyU728AuBIEmaNcYSSJunK5pTWqOz0R
YKtThYfg3sVFvEffxcJYqswrVTa9XH2g8eZI11JsH35o2YA5lbT83VK7mnANiA2q
9Vki9hTvT/g/9aqcG6uTFGsYH9d1bOjssgoSfg1cje9hXaZo6h5KM4IgWICxRNTq
lwVKagkrvKaMDO5bZGm/3nTemWouZpxkDI81FO4P12jv0p70BYdYbIhLI0ka0Ne0
10NMtKECvjAiWt/UeKi+dr2auwaMFElyXNZipOXt12COMX18OTNa9GT2k7dE9eDV
gBCzrS3bR5KG5iUYHZCmZeTTU8NWDrsxwi5RnoaTVVs6trz5oXj3BUJH6w4/35AL
VFhE/aUuQhUQpPn9nGoXVgh5kHzXS1aLmKv7GKDi0uP2q/1LBXGO1uQotTC9tgID
QMPfqpSjTtrO7/8rMv9QKTwyqJMqtRdxY545pHJ+/BAmhRpMGpg1+TtlZbz5mG9G
uI/Yo0lglRgd0HoKfM2lxbKH/Nk8iHyNOHvOzHCkMdOaW6c4aLUxsXkvipKV5pde
SvumlcOj6LXoQANP1gBD0JgAOc7+Ysu1QmHvvhii0Et10CMOvOV5qyruwCpN5bLf
gmFmQOR6FQ2idseCAbHytw4HnF7jmmmFUFxdy/HRHWWcml7Xwd4K068rxhJpBtIS
NSyXvYahk36SirDUSo74dMcjouxYbAALU6vVKj+eLmDizMLbviWW8oo+VBYyvduA
0sGmd0kNjhiwuZMBi5+HbvOu72u6w227IfRKnpctbrZw6f5IF74JiraaAuOycBAg
DhXw9eRQvbvTa8GUsGVzckVzoiyqHDQeapmNv9q2iot0VhKFg6BjpxOnnvagkCp5
GAuvA93cMe9a/6vWne3LEimRt/s/xLGaBSHLEZeqyOpusNuJcoNZE+ajvKJLvmuU
scwen9KiaoOrkwV/ogzFSl5NycJrZ37v2rWlO0Ha1KdDmzJ6/6dKWAY2J0M2Vjz9
Atoc0q49inweHJxiz/HSZjDGeyXl6A0nSPAB9tBVP5bBG3xNa1f5lJQ/3vaClqjf
RRRboenb8H9IOABbTgdgkgN0bJ5JpbIGKZhGe8rjUyBGjuT5HUtDQErpK0YNh+1M
xc4NLQhP1jEbeT8HeKiL0QTpidBpo1rLTJoaNJXp4FcmJZ8j9ebwklv0LkN7hJ3z
zZ8qfgg/pZyHJMFb11AgqWv6qXfQ8mfwjVkdAIjQ8UfVN9WsgDGUOiyyE1V+i55Z
oPygYu3Y8ysmAV8/9Kl5Y2zTAFO+hesJGE2fsNIFtGtrPRutCYMGHG2Ft1MMMS8T
fGyOjbQMm/a9tfZtOb7MANVkF3DpjpUFu/QFo6h2bzn1lv29xXstB754jy5ovgJF
+PlNYWh+8u0pGmoSXsq5wrnw2lKJt7P1lFgoFdSoyoZLLqL9ynG6G28ddx1zDZM2
MW3U1Q2s86XIAA3IYVTek37n6SMO5olX64OOVkQgEZnueCbfRfAlqHupNz1gRqoF
sqEp4oCkojqnu4NfnUgPYFhzSZz8aHryYS5eKg0HmpAGrJJFg6j8UVF6Q2igzbxw
OYew8GPvsGDWMIRJUp2S9M7CVg/3sx4whfsdZJ8Y5DZXlnP3JXUp00kE9l4csghN
zlhmmNNH4Cu3kr6kGiKRRJDuRtfvuuJA0wbfZLLtSOWhAG38AagPvxYCP8C/qx84
NDzq5KU15gdaU6BdJP0bI376o4hYf+VqAdFv0G1dwZZFZwrv1C92dYnbks2rvCeQ
lu2nnHNMzlNJdkIMQ9nBrAixHrMJQfJW80jLHWnSgGUhGVBzr351p/eQ1ukBKOHt
uMi1k6+VTZq7UqJ87KvCiM/UU/weBz/dNXRBQU0w0RkhgH5r1bKOjCushn7unPbW
wGMJ76M5mkfbtn0kMlJkPGLwiacXU0zsgtxyIaKySGLu4PE9CCDZ2+fTTKZ9jsWs
8mzfQbi0W1Ymz0ADH7GawQZ/77hP0LssOcKqdwA3rMGWB2XKivC8PD5DrmBwsrfQ
xwz/mC3xr85mAuzeN7FcXRLG9LsxosXPbruWk7Xo9ezR7aEo/68AOrbnZxPVSkM9
MequOpD6w8/jpQ2hpqEs/XeXofHsoeVYC3pZpizaQ6JiDcbzOBB3Hr54hN6YXLGQ
gU4/EBHCupGO2ew18nIiFUTGrlSmW0jARsOfL1UEPvt7XROSaBbw07Uv5WBo0G4z
n8/MTVvTwuJtnpS+d+dPsbZVt/8ARg6HIRTY00+UleGQqyFvwV5OmxF9dZbv11EF
XVtCWMOY1XhNKCVfciXwhYnpf5re51IJtLX28Yh4/Z9yt5J+aRpFbDBsN6a+kd2N
YLam/9wt+2mCGr3m/nED7rzeB9NofVYQYtTmF6q/itsle+5lDbMtzQjvyH0lhyhI
ZNV3Jfy+m3s16UrObSgCZP+dUl3sa1Rps5FJQERNtVibZ/+F4O6VmftT7QiMaXeU
DzIMJhqo9WmG1ebdue4odFmeuLJ+r7yNYYjHz7CI18D5rx1f/HFd+t7X/8z1DvaH
aGgXoR32Bbi5fUseCErPfLuWwPFXGpYa+xgqTeoqUYu+IKF2WuHzx7tQCb3ADN6V
ljzzMYfiobgDlyvA/06lT9l1XH2DG+VHYnWc7f2qzp2F+HZs/EV615JfvUBihKce
UWH18ZFdzidrnbFyfkY4WnjwqQzMWStj1Ogoo0R/BxbBqPlTiojZ86UpaPVgblJG
gUeqiMumYlS0tL9DtXkCu9pT+9Jy+ecd0oKBBVj/xbS7wTxb3K3IqeWNZF276aos
O3ele2vq5gnRZYE6dONmm4o1k2Q8uqlVeb63QpEUemXVQSdDXJdUNcMo7E4LwowI
1MoS9a+lUUcxj3NvOpVfBsjK3GI9Ved6IW2XF/N33OA2VLmNgvX3uiryIpsq78LY
dtOpPfmDlStsmyB4a4qzBspj4c73mOt/48doG9/wHqJqX2dIKMGUz+EL8dji7G1G
ijUArQCJIPZvIVVOa8AxiUCMX5XuTdIIH17V2OeW7WP2SwWhIJPtpOq6ZZYXJ7Ch
/W+AKW0EqBFWDUC7z/08blHjdLlSEeuCB022xFvQ9CvThWW74S2rKtxmRYqowg77
9B4eXPsnzpjA8bLFm0NdYSx1EiExUS/cMrVsfM7rDBdF5AfI1SdI9iybL5NzsX/k
WlXnlpUc8sC9tyEww6CCKHM+dLcrOLvQ1ErsvOGtpwHGdYJp23IdZaPXQK42bFGJ
CH+7HkY4w7/zPSN7MDtyxynERT+DWGJNNQmELpOgkTggpI3uYpeN3m/8yAVi9IIe
q3MqBbg2H0DSm10k8/ut58fhznSPjohT/7TXV/Pupesjq/R1MLRO/KOYqVYcNyPA
tvdMnJ7PSVZCuZ1DS6/RZTW7xsbBS91RSTfjrGAfye9wOklCFFDEYWW2Gh+JAZq+
cz7PWnSnrSYqDJNeFRDkY59uXrlAjLEtEjm/iyfa6VFMhJZ34dQArerZtKUjEhsG
ebMimV+GxpVI013f8pD2sTp+89VcCUwEJlqnuEbB0pfKiZN1H4hFiWbaNvbvgVwe
lz71K36qISPFGNaQPs5CNeGC5yx8CDFCEzuxsnNKJKQP0vMH2EyH97facLje2V33
G5HM3ZtDygTPPPnbqvWxQ7vB6jMcEojXX0p8IGqx/lthH52/Qan3jKasLut/ofdd
wvqpG3vuyFX89/8anC3LmWcFB8iF4FE6xQpYxxjsNl8heQYS/1YqtANUuQ94L4HA
CyowsF9tG25U7S8eKegazZZ4P59iZsOMGQdztBfojSm13h/cM0XOpeqYhJPSIFCt
HY3v8KzeKEwkQfaKvEvcDnd2H3FfH1m0da3FwgcJeE+OSFLWRBtBOH2mT3sSskv3
B0mC4bevmNFZlNl40K3be0oAcBzE7iFn4xJNxur9TF2Hxeabs8cUsTfvA7K8KqTs
2YlPxyh0T7XaFZhxwHqo7eQMoT/NZ7yovtybJwBgiCR4sx/lehs1oToAFgmS5sra
EBAC+BAtZGa14naJL1x8N6Y0MjfV3g2m1+3P73XJcrcs9raN2zrx/YK5H1peHjRV
e5DMfWvMHSKqG/CA2eYfGd8rD2hS5km+wDMolPRVlxem1hjQB+wNO5cR4AfSuf5b
PDQL4edlS6Uf66LC2Ih3FewlO5drGd8YQz9L5XNN4EvPe8vW98A8LJqLFJSH8oWr
bNY6TObx5lAQ/E5E3iMU3aHxDofiWiCPd2JdJpxt5WJQHvtjF8IcT+vYMvHpRbYj
HQk0xm9zHXH187l779SA4dKidvoTPbQFWaYQTG5M976PRADQuhkEnMN/ffaRKVuB
O2LLFXxBhHzNMjWRLDJy8xswB14cisx6BM8mFMxSojtTWis3YQQ5jfDNbbUy+q6I
IQe//TIeq3D08vgDtEMND0vHj2wMtfZ+UtQHOsOUb8VYJ1yK4h8Xh0S8tPaATAnI
+QT/kHwNelY/xGPrhmLYF6T6hEHVaXxNYqbrCDw+aAhoWoTMS5Bhf4fncRMt2Hkp
hxHlVchp9Hp7N5sJvtQ42/5O6UxjEsPE9EWJYfiJ0+7OOSkYMRNJ23sjXc7HAGHH
Q2HZw3J8/PpKfk+Mb8Ktvtss3m6q7/OcmkITrJvri+dCzAL4TQfNRAQrts53hmMo
XtxOh6vcc0bAt7vMBt28L1gVep4psYbW7i9QfewNC7WLoqdfbqSkI0mXYuzueTWX
Z45njtM4ZIOr+77J9odmiFxGNVV6E/FPSTBfW7bA+c7E59r0lzXXgdsIo69b/SKV
W8T7DUGBfA8/GtGI3PwezZxKtNo15j0rw2dmOQeK64fKQiVXlracRX/9at0ek+x6
Oi2iNmqOFSMFD1C2O+uYjhqYFHJ6I027BjS4+oPLzuuwljY6e9c9zbj6VyqI7Y0d
xYA3o6Psy3EUDLB2Q1M3/wvpOYc03Kiu8pPwhITdMcjjSUtSeY3/u+NvE1Q2k3zw
/vXgTCTYsWL7JHYO2FQ7lGaGenNNvEiCakAOMl5UsBpokf44mWQO3seoGGHQQah+
PwMFSsrb9mT2+YR9oWncP8lVHNcGw0wXYp9mK2J3wcvdgjzLPZHo3WS2j83rhAzK
LQ8IBLUM7yXgIhUcJ2tLCHHq2vqZewj2Z8KEne7ylhcsx6h1ue9x4dgK02hOYxEO
QnDsC1T5eLxnvk6sLSEOeJDOJozN4s1EHpZx6GNPIAAlEkqukrlTPJkxrBKiz+Zj
7/2O1ldqi9/LiUPNFU0mP1iOIyslmc2BzWOoQ1/QS16LfN8aV+g7NNx68l/3oHvk
YAhhCgTtNgrSdnVrMxa78Pl3lDO1s/LIxmI53Fq+NEFsmX9yS+DdUcYSfRjuNNvG
UhWcOFRFPQAUkevLS+vuP1L2YY4545ig2Nhensp4FsDifLP1iJyF5aK3fsZLCwd9
F4SEst8GZ01mQcLac8pHOffl0/LUnCFgqiy0kG1euWC5IgYsmn+bDjPU7PNEA6ZQ
IrSOj2cSFbXmK9X4zkk9oNlEzbPy50lidSWP7YnAh2kHxhVE8WsegUDZn24hFHCT
YrsxEw5hguh92UPl21YE2V8bgXwi6d1VDfbvlgFZ59MPupjEdu+r7ZZJQGeJ6h4G
E5eY5PD8SmDU6WtYvbg6AK7iAwSEmW7Y9DdI84ltUrksHdoB6MACkZFoQ8v7/+rf
ttlRlz6Bi5n3RHXkO+7zpxWCnDRUqbQgMCQFLdoz+UA5TX9Q2fGbjuHl2Vq2q6ig
FZMH2QGkJcvSmZBazbxcpuyIwKN+zaMe9i0r4qylU5fpyKCeV+8r/ykqZHNjnbzN
qmJw4nu0XUzreynSmBCagOOQ75/8IaK/JspZRXcpKWKmRFs8VNrhhSbWkqevmyxi
AUh+YSdm2mc2S253KnVZ60KzV+eED2R3I2PVeJeh1K7AJelC6pJU4BOgJezQPIO+
dIu6k204VSbiv6/gHxJj5v+YPAznagP/xegFS+KfnWoomOciJYTygU7gI2eg5wu/
sJdYAWEw1Rm59zYIdm2QCI+eH2Xwu6dfTclJw3rkw0QNjTQOPUN8UspLpseQJQbi
5bAVuBOd9RctygAgVJ55FW770Q0AvYUrZsU0fkMuSJG9By3+j6I71VY9VfF5SFUy
4lhsDXJGssOZ8s8mz8/s+y56MnCzj7925pQThayVycNM1DyZEQLq7XNQ4RVYU67+
Fo4CAAH2wDV3xFB47ah4kwowcUVLY6WFu+VsLF40pcXbrWtgxio8UdrmjG2+4P71
lMwwHjP3oOFM2KczRMuH+erMvh/kLxF5L04rByLjnX1ujnePqEV4O5n+sggpLjw4
k4WW2lJELWEfbJRIiyax5FjOKxpK1EFqIlwpwKwiKWCanLnOgd2d9w+z21j3e/1+
bcJekHX/NxbBUU1+qz0kXNzl9RI3OV/AF5el93+91VYsIFhMqLH+N4Byd40iX0e1
OlvxLGSwmzGmdSGEwxOlI7dBc5fNRFP5gWGMeuP8R1SxIzQa7R4h+R6J0cJYNZD4
kjWqlRhpd16b2lryC08XeMya9nfCfGOJFjrc0EM3rL1VaFIE4tI1Ozf0UUGBB6SR
yOKdM4yLFjIBHe3MMAQnO5JUSaSF8AHq9q5pd9DRguFuIIg+DfqKLdCdHkmcDpdR
MlLbaMaa2lB+o7SSmFfyS4ljFZev9T0Z2o8Up/Z4nR089Z8d/rotCUsC4GFYngss
muBZYMPx6wXuXLgCU0WNTjEQOZE8zXzIox9pV6QmVh6uwNff8TuRg04tW0NcofDw
ZrckXqt0M85kzIwwQGmwkUAzmboYUANFDld7XSYOSihTHF99NqGTl1SYByR/7my7
4dTMcYwiGXEKT8HpzweYc22BGM332bsCa5zjElSQagagkCBan7r2is+ZbMh7hkuz
6ksL3AbFgXeEXTE2DDZVuejE6/HZjPtYcbAohzJyG0ccDpwkOoMBN0ImRkpWGDO9
bZiILps4WupdUkRwNWEwj8Gxm1FGzSw+V55Hb/NOUx4Rwxjo9NWA07vsuQ3q2tyD
vNBTOTH4N1TcKqWRefCUxQt3f+bB+mEOHaxNqOkzjICuCLA51KjrzcAB426nfOwi
GrpY/QOMi1+zwGBazOF4DJvVsaMHHIo1MbFhEGDXdD9HigeQvQyZUpgJW0yh7Vbb
q0zQ1jQFuzN5hXpEfsV/F4okcunTCXzQSaklAWFly1R7z55FDi2uBc511e9a6R/D
GFh4FUJzMwLl8Oal2m92eD6pViWIQpzzRTaENwTD9aVQSNwgLjFt0z08rxfeXsHx
ThPExmzXiRO38SZVsJk2uaPKZjnNZ1jqMkPjSRMDUxha5oQ3XFDeyuIDy6EBth3x
xaaeh/7gzwoRxCG7MeLtBgdta54g+PoCJ5ZyYFAMmPWfmilfWphy6iJwQs2xdVAb
W/AlUUmRzJhogF6LFKz73Ne2pOt/fIIo85c0LpxEXJxfiHfFLBOlZrDT/0vEqyrP
B9R5oWkedFer2LHo24lUsrVkKG09fXegtYv2u+g9S8arME5fSh4+EJi6AX+QDF3r
dlbbuM/H8GePowOdkyvPs9W3MhUkvZ06gUpgKTs7P69LEBbclFfGHlf/dKILKC5z
E0RwDucCr4yJQvRaC8u9B1jK3nlHtTZltoBwI2ZNfbwhJpvjnJKlvtrPSva8hFDs
iq39DYQX1VsL3TlfQWOaFeosdPwdGw554A48JfdBs+zsr1HduN+vSjESJNEGiaiL
AVZWmEtnm14/WBxbCJmyQP4ixIbIbiGPvqDGIf0T6yrk4bxdiOT6OU5NXy3RgCIa
Wo1mJ2hfKSFcgOsC3tp5VIl1fkn6w1kvQux8Lo6V/mv8edaUdL3qYy6+W/QiCDb/
06AjRuU+4SZhXcOchjL8gCYRvvm9gXSP9obBspespheCwqEAFIz1sjNZwuuni6sf
bvoRnoCH9hriloNd+MhvpVB5FcI2TgSx5Dumq8lzFsnMHvGg764DEc+IeJ/5K1Ma
KFM9UUlv5a6j/OPl74lh1VD1pElE2xk62peoBtNhQ9eB//Cpvwzq8y/4W+aHPotZ
deGj3uK3TgPqww2F6/0wKfR3x7HUbZco9wuV/0CsaFBSERGcmSPN4PiooN339dcr
kXSvZ7eerxb+1/rrxqpL+YYZXtOkC9ffzMmx7P2TZ0FGoZN3aFIPoBvH47hwIRO6
u97CcxCMyijnIEvRGpbHKMMEyqEsSInvzmy8Sxb6SSyrbY4ThiYFUxoP5DF8uZoV
wtM0kQrkYL4qN7UexDkHvR9ZihCcgtAdCRdzZqdS5YH7IxgbmAc6cvED2H7zeQlD
myKLwMjL3QeX2gYlEnv2NrGBPy1e2+U5z6aQzjANcQwnq9eH6A9j6fUx+jHmBpp0
wgrNLPg2o0mOOlAsiSjA/lBkk6vuFFgD1Qw7WsXXBLuvuT5MpF40CVip3/UDqV1v
Kv8+njILl6Gc8w5gkrU/M3SkhNMCjI0wl31XZOZ4k6GzrDjnDiOH66DzutpxWEvr
x8dLP6rHS94IfTxm7f8RevR5ttDYbVjQ/uylM6aDVmWfWPxhNJOCcMLPyoJGl/VX
nsEImDQdH+hegDauzs31kfrdeeerzZUDmtpBip09x+S+f1hdmLWicbM3+3EZaLdX
9vL/CoRmA8UABVvHs9hT6oxHDisz+PlYE/Mb8oSBYdOF58LPPevWBH2PekT5PANw
E0HDmYL6TOy6qEuVeUbqxaOrJJOUm83nvobl8DJz3QCEJyXuu39XBdhio6npyQrW
vWHA03XDjhuRsiY7hymXOJ8P5k8eYdq0++fs+ZtGIoIYJqusqcMaQQynNT07b63U
ba0crd8oBZ6vcF2dQ6I3DzE4VPja8wxIY3WQkkXMuqz4k+jqfY5Tx3FiAYZUwGvP
CpdaQ6JJc7UP3z5pshC1ewtrEh42c4GbLBdhaZpQhIFZ41q3aFwwX5x0kW69lJGI
Q/pg/WRWxjutFaw9KaZUaykSK/OuZICmyDvL7+OLTfPmXJGog0kH3KayiNv3PafQ
MWQuOKwaDhLKD+d2vbH0sYdCOziTZpCSMpW51KL2DesXNGdMx0DZB8Arahwv2u9W
VBz0xQV2nb/DUuJ1i9lTBcy73bpbjrdsXGAtMTZvfV//EchmzXyPQ7gZtT7gh4T8
gV0JqBucuZQdbIAyJNBSomSS82+XARi/HeFh5wO7+1fDS/Y9tA4GoctDcbHb9pgE
gcsUB2LY1dSQANFbvFY67Av0fU6f3k4OBmZwlCrO9AXUM9uUURNRN7lyHdvc+dSJ
ve7qgxN2wUwHh5AodIR8GAawAjXuf7K6UedWhqN+6S4QePea5IaZcqxcLd6MlLwQ
jc4HIqZqnrZMCL2m7ZrpysTegbQzqqb0iCnyVyR81BThpW/Pg6a7wRUmiRm6suQg
pRKVLJ+xDViUt+ORwB36xWc1QD+yJnWmy3bJNbkCPn5hkzb214hmwqzS6asbsv9e
eoHKcRPgMy4l8rCTaCDBMydhjUpcW6FhaRSqvBFp512Fy5dBH3o0vwQyagiIw3kN
1xVCacy0BAjGOaXNITiin9YR16awpGxHucezW8GjcOqLj4JhdYI9EcEKdaPmGhJb
Ypz3+bu99AQ6XWjwHX4PASX8O02W8q6CVfh+MFDKdjX3CLiuaIoZO8fbB2kYDXFB
ufJ5Ho5DF0UxxhiwAFLC6QimiQjk03GvnKU1/ILyFdDA6rQzCSMA5gbpuHbafipy
Hs/rpoevCWna2+kFW0qqsJZK4qNONgX6E5DD8/UBlS5Cib7OdahU5geoqCjibndb
CXGQdATQhs93hE2DC/HPNJKygsqeCc68JnCDn/NSjFT35bzP1MoU1lAtk9ijc1Am
B3CsFYsNVGFRjijOpr6vPcJcqlkytz2LuZtZcTJeSoX+7vPpYENcxGNmjXzccXho
KLW5jdYm493cALChcrH8ur/GiBjy/u5/NKcfjRLd3ufE+MBYID+Io7kBnIoduH95
HoonI2JVTzYutfElIS3UeXSw+5JYVlt2588vyFjk3tjG2aO7J+bHMapVO0BkL88O
MEYtAKe5iUaANpNiAyp1csNmXckDuw3eKMauxGO6h5erEx9pdDdRdXvEaZVtqrrz
yZlaYMutwCq2TRImuOcKtwgjv4D5B0kTBovkr7OK004WAa5jjffYqBmbF2lvXC9U
pwzIpAqjUJdUnBys1JOkPHKebMyeQNEtXhGbztoWwWJZ8GpDdP3HViQBEfKmo2BN
DvhAj30RoUnqhmsahlE/QmfGPc6Q5T1sVblrOJUiYc4avBr1NZUgCxG8sR01aBXd
NqSarZaEJ1OzbMlCc5FzTEqWmaWl0GmzUiHo8SnmZZZM2IH3LGIAmg0kOjY0JqM1
TR61h+QiX6tiqpVljigQJ0ZAs8s2HpYQNrtppkIGZFfvR6VG+YdpesaG3oLn/3Hd
AExH1sgg4WC0bmvGCkOGRR379jL5kyLGlnSAHPje4DVuKG5FH2BlIctde+/U/e06
Cjoo2k1B0jHyxAefHyxcWsdzmgNw1cdQkVT3NabheV7Zy//qWjUIxd7P9yqDCEkJ
qBLKR4a6cRopPMI53+ZpYYVmEecMwIesc03uBAHJ5fb3qdHFeCoLc3qt6iNx1aEb
zS9ltPktvw0UUcshKM3ci7PnBnex3qUniy9gu16VM06dC0TxFP05clafp3NzXnvw
QL5GZhILUq6RHzYTdHGY5fNLqoyGRtN4cblbblQPEsem7NlrYxR1rGvtXr66xKwV
3FbdlBWq0rzuHQ1SFCQxpmGRDT4mGJGmpkRAd3b09ZZtK4uZXMESVg0X+npg3O5N
honXsdItoG1D32mCe6vguyddwTmZCc+KWVEjgj8HLis/BQFv9keZPcAvRdxED6kl
/Sq4TO0oajIss9R0Z1cZRN3OxwPQ+SVauwbol1T/3ZMNb5aT2+RJsdzNh2PH6oKY
Ddshi/Dh3Pk9ZTsLN4k30gGgEHiuaH+IZXFXVa5TmT5VIZUjcUZ6M6qnjhMaBbYi
G3z+qPh/wcBvealehGUyQEvhVOuc8p9wtnxTbDhOWdAAVVHoTNyjBVQIP6SeVxjg
mF7eauu95T9qYMpELhvQyc+8WLqB49WsBBU947+knc1DjkJEdyBmY845teQJK7SG
EuIPAcaiASL3FmFvCzgD1sttVhnTOWJFQjfpEoYpPQyPCoBOEpN/AukKQcBgvb+g
t+hw1ilhTxWVnBI7AWsik8Q771QPEbZqfGT1GR0Zm1ayQMSiAvp8Bv3w9BMdxBIW
BEOm0HL55RhhFP43H2QgsbqfAi4BK6IzFvy1ssJ4fTL5Az50X2meE3J6MiE/mj9p
Lj3refa9oW+S1teU7GwXbr9AQABDEBIpjAeHg0gzMrmqxHJBZ+/ORgVwJkn3kKA4
o0MF+P9mGxtVDmZjMB23yqeNZswDkDnVARf8ZAhP//17fMuuFXFXTV3DySxry4Cd
txgVIDmYzfLIUMgGmuC2lSmkT969MLk/tVI/yUgf/ZFBFM5K4n+67mpc0y3KOvjt
s2qwyNjqyW4+2f+ra26/oQvwIT3z++ESLjVAzKezDQzMMogUoNXR9bxmw4iK+eo2
IsSlels5gCWRZPpjufwzg0i5djqHqdxNgeJTFBuNs7SQvE+nOsayWzLyn33W0Cz1
a0M2MsDTH9pjOnfZm+n9ikV+lyaqh1y5Hsj10qAdKWYVeurWdSrodMh3d2I+P5xq
UXrHxcRhM/Ps8Hp8BtNyB1x9j6WvYFw2NqFqjhD69LEqYLJlT5zK9FAJPNvM8FSa
CVYC8S+2goQYcxQv5TT3ybms/dUYEFec2/jH2/UHIIeNIA99NkFApM2g/RVwhxoQ
wsMubi9Xi1PgQQi+6osUnRzn+AriWcnV0fSPVGQ2TXwBBMX1A08uWnGnHUvuELtu
+4MQwh60MGNodbEuIRB3Q9iYL8IGWd8FYipMw9rLNDNYzsl4FlRn4l4XlxYAo6mr
og5dK+tipDA11KaoH9O8bqf/l0MhlfSBjdd9zEQz/jRDFj2pLc10ZMtA+2+Ou4IG
VbJEz0StO/x1BJCDyKInMMnFB1mtGh0EKMfrsMNKOL6jmPWvz7ZgrK5ZdB7ceP38
GCblTvDJ/hQBb/QSQ1mwKyEV3tff62D/Pg3EDgrjwArJG14R5LN4wWQVLSw+5TMQ
JvhkDlcyLpVlqpxInr42sfQYhQuTi4OzY5sdUaYLHYB9taXcuF1hRyPF6cGQ6Vj9
mDKOriMtpjTiT648GanU6EOzCMUEVaY3ZtIKGTgQR/mqEQ5pokgwel6R632Ml8g3
t3olYvnzHTWC3AMHJDFXVV24LD0HQFKgHdTWpF8KJiboHhQ8PlpCHAx8Z4QwF5lP
Pmb1GpzDMCb7fUdeGcxDFfd/G3obqy6+m/zbmUE4L1Y9/FVFslT7tsPWg7Dvr8dy
9lFdylzzkjMcYl5MRbZzxdbbrmzSvHB0FF+DyCrzDsA7FXAL0RxTmqF4fSyb9Z/o
2WYH3lspJ+5Vio0kD1KbJTsftnTBM3BnXJPZEY6vYH6BwaR94r54bNtito5dGc8y
6DQVqAovh+mf1ASzJW7ll+JoXtf6JKCQc0PtvTyq2tzf5J38Vh1Ak+xosC8ssj1H
cjblSmYxVeLzMe9r8A00y8tU6si1SD37K/fwRWm2OETQyh++mrcP20kW/E/weSu6
0eIbUavuVzspFIR2RaSWTKpNRs1go5dW3ynJdkK39F20IBCgfQZDPNjwcd7qyfvj
IywSjJejZVEvO7kt0JyGMyAPCeZoY4ocftVuFhun0BE6LqmTEABX1NHG1eq3yjvy
w8c4Zj+w0QD+kK80WJRVqyASPl0suLt9nPUWM/YMkX6BSHuYxkRM6csx8PAukuR7
nKG5HMLB60aOKdfJxJ4jeAGb1QY4eCipjPrsfq6a9FJaDziyShHtTtBTCD72t7Uf
cxoA0L0YzAmfceOaFwQDYLT7t7ljS8tWqSg/Pxcqc7sawRgSXUeu+VtqQeIbq3Z0
LvHvgSfjWjLPfprMbuy5MdzSyvRb/srbb7wZX3RcAfcSH6aapewRm/ZXKNvno9Ld
XpjFZp9EVG66zH00DGbp5Nwe0kS6drjg9/0F/R7JP6bFwsql0Yb8INJDZ96Tb7o6
BCqirZTClTitlQ8aHliKCDfrkv6xELF1kGmaFvnlIM91772kTcdn/0DZZj45gmLf
cjfKGR7fl9ys8woknnQo/H7GsGvNLNRyruI9+1+RtjyfAnoYnz8VJl1wl0tG3WQj
ZFFDvAGM7Fnr8wl/lH8U01z5gosshXjFEtWt+McYWtePPSg9GqcwB8Aip54O7dEc
sNykQIaw6A613OKlGdB3vnd2cHgs8O72RHBliKina9ccZT378jEY4kk4ArAekTMq
mRGgctXmUXrXEroUiCriltcsNcO2kfoclBaqv9VU9Zpy+TdMMyrK2I3tF4aXu4aS
243rmyLb78aKYvgy4+PJndxU3ASfZTaub7+4CTRoXcdvR++NxMRGtS4xlatVC29U
+vCJX6gfs7mPAAb6NOPypgksvI2KmNzPGbAYgrVpyft9GfZJKAYCmj/SZowI8hTi
Gu2FdZ2KS9twmrT14YDpaugC3sr4z6DAj+dzRmtybVIyz74yhxy6hWJoWUnDmJnS
2bB2CVtwrZSoY5UUaJqz0/NdJJ6VZRo0M7uGXAnCu+ZRM1V9cbX7yLkt5VoOdeQy
4bx780bJjRuf/sSH69ZOJo67fOP8JzPyQf8A2oNAO61EiX6W5azxqv8KeURxrXtK
GFTcN0pAg7hC0SySTbgPvh1UAjlRM50+lLZzsWonQhOSOyB0U3LPRP9kL3lldBP3
5+FdGLQo2Z3WwmUi+sAF1O+VZ9uj1iYHnD0FRizMCXOF4q/fy5YBsG1lUqX8m+2i
V6aEC3KlA9AXfeJL7QtT5zM5NmzDdaea5hCUjl7ryrhcbYWaVfj2SxbOkMmtSVzL
kogA35xWEzZrI1KzdBhdob21p+TfL43K7O4PCnmIGdEHiyT9wMvPfAXa2SAAJzZN
cEPln/eFueqJGLIllk+BKwEwdIpeXSPDiCZigoB3fiyw2ZCAdTePRbB6QVEK6gYZ
oP1ZJuQemcK5Iokbsgod8FpyA7cLDEJILEk1cr8JZyWruzgR07zsPMgE3OFTOtXj
aSXvT5Rp5C25okC+lcTyCS8SnigaR+qRxhs2i9pA5666giqFLUDiLAqayByoJa9C
Oap+Y/FvHIXOqWxysxKPsQK3POb37+92vTIvECT16tYG+BbotP3vYh0OzfRszfmx
3VSYyg5QIPdyT2RrLVj8ZjG0gb+Ldli5tUj+pyanCRWWc4AYETjHI3F/WtT2ZMLY
bkcoXLKeglyAJZIR/+9rlFULv3mtRfuTL31UlnLseCceSS6E6s/tdZJ9CW+T8rF3
gbJtnW2RdvDftf7hl8Wp2QVaXZWcyRJu8AonQFRS1mbv8PI+7Dm7mbqqaBpXb7hd
EK8l2H+jcqhGvAV0c43+DEbrnH3jBfHyqkQekEZb5Omc3KSsB3P1xf4aTHFNNHhk
bJNLvny5OJVNpiDvBDjq9iEKePMLB09oXlKw39EJTbuGozoH/6kzqP+v+ndtRQvk
b2p5mnNHEBMoEvDtZZFjjJA5JFKg1OsskyUIcDAdau48uiMBH0U7wYXWISdTd5cg
ZsgKdn5HkQ5fnbUqlUUrLLBcVFBAHBUA3jia7/S4HZ+IzSdR+1/L+FXgcJWJe9j5
yyMChOu5IRX6XH/27tKmDgnNzrDNjUY/OJhxf8CZxHox58wALbxF1HMurnRPBFep
gJ7hlRKjl81HNUOdjTo2zPmR48IeSAXd5+nbZTzN9mr3aoi+D/LGsyMNV1jll4NL
vvN6tirSXHtC8EmKO+t8Y9RRLF7pi68kv1gGniJyN5PmUF1xGeKI5vdB2MbnFdk4
bUnchr+8TgiXVOG9kpC16haY2NunEhC4l2Vj3RI6WSi70MbI2G6EakOwWYi3Fgs+
KEEOB94JQZmVVVOSuO+xThd4sfuIGrjaKbwKL+M7TAsFcrEsf0eK/agzIirSLfd6
RU6koBj8QCtyiuuDZt/Tpy1X/nirVDWf+/L8ymefTwoVmX+11sLnbmP7ClMsAGJV
F1XplfqW04+XtyX616tTzEWHKP93ceSeAlW++DEVI+UNEpI4TE0JS6eg8sQZ/PWk
mpjWp9C0IJ0oaOFljBTOXPpM+BGz3EWb1cJLvoIZ/pBNjbLXVb6wtJDcpexiCrq3
tL1IZIaUhIkULF3yRJeGqzMYLu6E1udAA5ZzwV7+WHy6LYyg9JHUaKsuen3kQ4dX
9w6j+DyCswMpiddd719hndaCegzuO/zyngmwaYzjVl5ih94tcq2WR0KuvauSuTlE
WthZTYiwRnNKGI4VfGOLnO7osTq4XCJuUyi5Mks0l9oy/hldwOl55RPyfWy/ASsb
pJqMTlLovZ7FnZQ9ptyZAbOtGEA2uqR9oCpk2bq5Ow6mFVli0fAWD4GBoP3awBWK
sDmfpQ4f9cZgAJ9uZJOTbl8ckN3O9tnRLukqta0sG8SHSs4HCEmd1s3KUAJy56B4
DRVntJSENEXmX4SSsV4Frd6ZMpG88OMXYkltXpATC79DW/8S79gVonId13fG10AF
QUNbtLxKPknjrXqT29SqnJzvdiEOe1CshbtJF9Nu4GZmc0YFb43paAcehpnB1dWS
XuQAQHe9kA04ZkBafU+RxZ3RW6QZwXZxBsr/itDwfk4LREAkl5O+FjQoUSse6h52
xjZufmfa37f7nOLjv/sm4RO1bUvt3TduAZJltoe/clN9ReCvrjWoNZAzl7MhJ2j+
RMNGOvWhlVRMQ7gfXuZZUcrMGd5UZPNJpYPD63Jmb3jsnYFvPLi7jVWjFiDN9tx+
hcO9hLf9SnPRRfTcl3eqYUIy3vARbTCjyRDAyRxcpyWjgvKiImhP0TvzdH34bQG2
qzKIm2O6BhR30ZxQKcPahUQKE5S9gRJomam7zfdTsfYRrpYmi3vKEVeateGacbS9
ZeJf7L1SWYix5ZwQvRAYrCJqVWCNNI1CLETMl7RIwnvRy1CFe2Qk7V7XePl/Rnof
jOSMLz4bm5hQBaxSnz8yElyec5I+V83FjnFBO2oj2fr7iifz3UxOjEeMNfjZvXSK
oP7Dkcag5ihYbUdeEkVgxq24DOG1v/5eCFqiQr+wa2tF96h3JYY5nkJvSIhPt4Sw
aYwGe5kfmyPAMY8nbA6NGKnRPifWMzjED8NH0pbMzbzocEt0UU+hP5cI75Cr61Gg
o+vFR/jfteNtnrVLVQbI11Vz2qDVqgteifyWPxgf5B73BB9WJhVHLgTuhnirEeap
tifGHODX0md/kZxM3Ya3DYxU1tXx/1WLxgmSObLXHTaaDWQLtLvLgbPOoN3HNnCQ
zcXB/7+ELy6NOOOtmS02qxjdKtU76sidax0gL/nF30GotGd1R22KGH9ppMZfzWrl
J/Xo1R0dbt4Oyav6lone5qx98LE0ElLyGDWmR9XOPkQebhb2xTs7cOulpT9oQ2wu
uajCM6oOswUvJ++3Hyc1/cTtiGc4XS5Ju24lJvAJjHp0bHaAmhn75Nx1TqKUcwDp
Cs7KlEysXrFGmW4YP9DAEsWXNzDjj1xIFb5rHe8+JFzb8Ru5EkDaMHLihIplhpK8
QvNJZJ0vkn6PNj+H0bLacUe3b/96zOs9wHrK4NMm7bTnS62qSM7dUzzE6mORybU9
ZtX6r3BNGHExmabXBNYbxXOjOh6fALs8zDHk0qnM7Yp+5apWPZZUEFhUc9JufoAO
IGKtOqFqXVLXzLLRAHt07uAgFSn8Yaq0TeMCfTK0NiobC8xjFSIZJQdEmmteVJ7R
ohHWUkxBnCkl70OUB8xnD1iaAYHd1Slu1drgWfR2t77fzJBMbZOleCrVXVwjK5Ch
O5KJuDSISDc+AD1CgIW60m0GOAXy9pTc/HSAYxo92wRo3L9uml1MzivC+33B3ouR
4JeGckqFf8suH63xwZH7GQF13IZkTLtORNDA0RueK0UmHwADzcWQirvMsmoO8Z46
+AwuTW4W1bEtJPfYzr2uFRqjtfCO4u9xJ7ai+/Pzz2mhYHUrmNXI9zU+ktxnTNLp
grp1DbjoRIImKbwD8NDhghNB+Bb6tR9BRUCfkGf8xiDdQYE28Lv8DAvleFpztAjO
V3zjHDg4q1kpHm2RGsQ84mUlw+MRn9yTZxAOzg4kliH6gHv/4zuDdJGLd9G4RThI
V51VHt1BIh6nDZC1rF817vcX8VjL+OCiGRAUkN/mXkK4Iwl7rGZexlzHbEnAesIr
I/UmfRe+YiaPcSlfsyxJvMt5IQ3eLz7WZgbsas+V23A5NhSXbtnb8bpxhZ2dr+zd
4o81KFILIak4NhY4EBFu9GlMI3z8iyJ0awerygrFmDezerToVGGdS8bRQdKHWT5p
0V3IKYVJA7rNQ0uwJDe8fyjcLJshW/r+dznyjsBTqGnRnn24D9ZE9MfAK9aU42/F
atP32q9cYzPb3Jl3vtsRmCiDVvrqGIf/xYHiMF3ERUShS+PprRlXrbksAy6iD30l
u/vleSHTv46K4W43lH1SqLzuLg39KQozect4CGBTfNMaMNdA7MKew1bsdx0enSOu
yeRDGelEnttI63GrUbJoqhEKWrmB8HoxYCK4h+CDRyrtV1wrM2zbwgzrNqMCmef5
Mx+LbnchaOqv37Q+tHL3slgY/+5lJOGZUdsz56JWVUz9nBVeayRvGluiaobwy9x5
5V0q+GBYZj4l9vFA/+02ZodwX99hypfpvW0dRZsG1WGIbHjt2D0zVD5d0QBmBgps
V71Qedqr2+l2WD5CEe6GKGDza1Ooy1cmLNSvsRgr25s9maYgYHkXD34OvdX8VS3T
rv6zaJfP3fyCFvoZARMR3Iu357renuOaGPj/LYrSvT+4ScB26xY42ZNuENzjAhOk
TiCnSJzrZC7lXhWvctKC75U100yE68atPPlm+jI+cG9BDLAPW5i9wLiVquh7zCJN
A+wXrphFmrAcmPV5gWp7raVXJcVVkJq4zTAWBhMgBX2Y4WgV3X05jlfAjN8s1sWL
3vF5ePRtoGCt6XL5AwK4gy0iEwQ3A9PPJXzHSAqQrJ2mMLxLM1fRwtMuY/kb/x51
/dG95N+YjvdDkuhTa6jNfexRZsunBKe4F6972WQJucQbH/uJUyZ98kzj5dYDBaF8
cKgABU1FllkfC/sTjrlhu6lS39jPxduU4Tz+MpNia2NJhetJiIMLzM1D9fV1UYbg
erVT4Lm5pp6PpLjluV+t+roM9blHs9oOeB0hewdNzm96H0h3c87tSso7IrUgRwQ5
PLSuScv+uscx4uhJzUPVnRIl8EWFzp/rImRCzviQ+wxsdDbyVVdep0cbLwkY6Nec
oyIuHwKoUdCi1iNMbeAZpAmsCbeFJi99EfHKldp/ZtImVa+bqiV78YaVpX9+SsBT
TSMgu/JbwVon44Z308Pvza19oSWF53+0AI/NeEGkKgeiCysvqYFhtqYKYG/CQVRF
Jd1gKEZqX+gYBjRuJKmrzQwy2gnhL63ov9TfglZg62DkEI7dqXN8KETFcSMK9tI1
oYYIHfkrVR+bQ7VV+R1Ltff3dYKwZeKbVl+A/VjCafX50QFVTjv/ihLlfi4zVEyU
Y80R5NhSFLh3Z1sIgfnPNtN8XBrBW3KcZIqzsqJRkPGNSkL4DCMGequZF+GVy38K
slcobZiEQxkV6Xd/y2mZobPdP/7UMZse041145MsS02wMqAmd1xGXBuVqnlhqVBM
hCSOesTkd2+Rr1NFSKtHcGpLRa9OzZSw+7u+WhCH6Vbb8qWPsfShpKEj0zWgJMHf
pyUkG2gVuCCSmAjLsQN3WNDEL9zUJZOylzUhcC0z0ftytNXNpE3MldA+D+GD8Vv9
CQeC078dUydywV6Rarz3kyJFBkWSG5m8sczZoedEH3zBED8CJDGL+SAaEAuJpdej
unTEZeEJerB19VprDL2CARnw9EcSQm5iw0cTI8BkOaxqrD2rLRIZKnSGKShoiSal
E3ZaaKolfBK5AbGzCSUZv3OQQGwV6yLBPsW3M6Blj1nb20VS2Xf25vNqLL1x/NCd
IGb+cYaNER/2xXlfMVZxr+yJGM4TU8BwHh1W9UXmA4nYwpsAAOi5a5VL/PnLsjf7
JhRss8L+B7lsOcPXRYMVu09/YXIwqAPMBE0u1Ywq3xGK0ilNn5GZPTksyQETKksT
iM6Cj9MKFP46JnR2Om9vbkou9TdpM6yvoQtpW69sBSR4iRZ+pqKTCZmNW4JCv4SS
EWGMHAyNpS+mYUCk0ivcAIj8DGj0tpjcauYkLYsMkU+eyqqCZPDZ5qU+yI/aDihJ
Wv8G61TEGJYWb5QJQG7KETEOrEgiLFFnmZJEWI/hpqNPfm9vl/HYvI+nqnoSSz0r
qxUFkz3u1VpQSYgRcblWl/fgcmhZwniL8AwTHnQEgVp5IjfUVklRhqyEQuWNOprL
SZg0+8HL8/vAGJZ+9UmuukIkO641lxVXI1gKoQYrybPULlpDuOY7zVK5NvziZUlp
AP2Mai9KA7qFkKrv4Jd3OkheYOVegMgEW3BXHgpMPaDtqr6WNvJQ/+zthF0ej14q
sNn7J2JRKoSOLd2xdL4wsab8SZfQQrXiKTvEiLBwxZhTwXDKqcjRBQL59HAtC+ft
NrdNQjCDFw+tlNyRAPbEVenb51u/ivJ/VwTUtRmUTFsz9cknnhuyhWEDjs6FRS6w
ZOunGw/Dlw1QkqJ9CqT/95m5wwdy8qhCUrckzSh0t/sjy4OtKds2EOnDBHh6uayE
z9sSQmjtEAWfpKkQHDNTxVi442wuGjwuqmDD3MLD/qhIwtHHtpcWE0R5kQAspcj8
f8FDTVCTWCjhpE+rtHRcyLfWiGe3qH7HXGChFtsLhDbtPl9/exCdR9wcImqVYqoU
/KiAq2BJ/CLf47kG42ixpmHeNx9uMt14n0jwGVfbewf3TCWVE3M77a6I0CfESeF/
AeI2He8xeioIiCVQKBeqH+Ig2/DcrtANzp56+nb3tOi5JMUFQiidliffnvsm4UbZ
D0ZX0c562KcVGqyZragiv/kbgGNvRSqQaz+EjNQtqiI+Z2oVbJhLKDCA1bWS5lMB
/OXxGwFJNw1GmLY8CqnYOsJsqG/C1c83e5ZvyHwWe7IIGl30LAWDJEaRJF5cu+gM
KzPSYXfultEsZ63CBjXVK+ZpNUd9zkkzacFQ1ftardehWzhTMrIX1J8iW9JYqNdv
40pxkStvqN85a++3iDWimf1on3ONcrKhLGcFUZL3IfoNq0sZORJMVlpxsZzi82Ho
Z8OSTqllJHYuiolcM03Va4yHFWmr4xl3h8tPgAgyNao3Iu91/C86pdqNlfnUwEKy
PP8TQxoFNv5qHQ7SBMHRwsG2wW+uK+ZtCPZqaNMy7s7z/2hPuvAvM7g2JVETlbHF
4WwqtVbK7lI/oIZb0lTTOmk352zvWf0oPP2IaJmrFVCd4p1c3BuBQ9s2STkE6fn+
KGba4mt/abTWKXs+Cs4is+OrsaJLfq1yEFH/Lm2culsH5a41Cf3CqV7susTzml5w
XYYaa+0Qgdjc3VXeqGshaDNXH0Ja1vnAM2BsWhZTje0hHGbJYNCY3dmIULIi0ycY
TiKKSjqLjVlDWUXYF6GgYTEJa5nieeL7qMAS8hjO1nDkiS3TY5yV9FnK9h+isB2r
nzKszjqTPCMZLIsFoQSXKeridMPn+fCHGmGWMHdUSyLuBG14zC0f4ROeiBLjVwXM
I4ghLoKkD5FAnAflozleGzA3/RMcJ33FgmQtnmYtRaJ8sdlzUxzGWTL9j43J7mL8
GKwV7JA46evCG5QUuHBE4w0ATwKkOCbbCTTWKl/EUCj9KSqlIgU8qTL7VFTF5VhV
SaTZxaDSYXcu33xk7oTt+rL4ILtbTy3k4m102bq5uhU8vy98H8o/eMF4vJQcLDLc
EaNW6FMKvpD0d4cYDkVXn00LnIm18/r7Dx8QdHQ1mFA6tcJtlmjjYoq/iNyjGH5c
7fIlUs+6bE7niRVlApZ1AS5gsJH0TldCcSaR/54skgbgArOYXJH4MaNB1S1rOeYo
gPAa1aujja4H2F6QzNhiPrAg1bbx1lFn45LgCnCvPPVTTwX//eJd9nZeCRkgk3GH
B2npCJsAIFzTlU0wEuIiaX/JPgOJx7pG0tv7Z2UocmsedaTlCEKU4A9Oj5DCCW8z
xfWhuXveqMVqSx69LcCq6YlcKAgMYKE+qE3gR7HmnBbP30z8OEJPO6UjJMcQibgQ
5hcecrIPhIxfZKw22j5XVg9ofjdpk7ikhxdyAFhr14EHNPAkEdc3DXktUSU3xS9c
qqr2m6KFLLoAFgtEnfiBMPtACnHhma/6fFz1EBD087JE+yQG1pTUkyGtWmTnMSyW
HsPT6A7PXuU9geKK3IfZgKIgGmdsWeZ+4Upp9j1WPSh81O2uDP6sBdBb/X/sprkJ
wxSR07xts/tFN28lSnVSqE0L4VGleL8zEG2pK97we+8S3quFpvyR01LQXE+WnE6q
skXizt0ARSmCreV9MJKFrZIZ3Hs8FEj+gQyN+MlC9BVQ2ZP863MSEHF7iBLdQ33B
xl9hSA0Kiot+ji7pAOvpYWKvf8BHdbwlCWN0cVULCJo3aZR+vU9Nye3shLAjI0AL
1h49oo/YagtbG1EV/gwgKxsyEX5nTWizrjRzX0XQZse5Ngp+Zo2+0XjRASk6Qu5Q
VaJdLB4FVOUDiRoJLHFpQpaSwQxhExOPfm6T/Dc8DAMSCtcMzGfNPGTMntQybdop
pbGK5D3vu6bYgdMPG+hkx4KBf/x30zhZzPEj74S/FHFHE9ep/PuYN62GbX3pc+SF
5wtX+IMQR5Z02Ekd7lm45n/1mylvWhymHHtUvuMzq7SJV5d6BdvltYvZ8bop3tuE
CN1D49d+kO/vxE4Nus7Ev3nPeOj0Vbx0mPw8/lm7MqEE9FUnNf5C7xznH4UvEFv/
AJNBnvRhfl2RHlvylFu1wzEAabPniGmbjjwBDf7GBiDiDt1Pfug/6esQvR4IpK4R
0XjEdUCt2ictdc3657rkTSYF7VnlXgsz2jzdyjWCcBENY+yIcYvtcY1S5w09TiRw
WBpKCim/gSf0OUYJZ46U6qocIXTM6WqERx6yBcZxwe/aFYrE2xKffrD2gaFK5w1D
7imKmNBV90xXGEKiUnkRGh/n1MgZ0Zz3sObAazBBdIkanQrNiwW/K5lY6XdBKvuy
S7wEoVJmUzEvaj/rwxpHiucjHZDbLbdawFdaXXS8jOYLivqOgxSv3Ep1Zx8IFVgS
niaTcM2ytdXdl5LzuNVByhPVtwBFlm+UHMokNba2F9uv2CZzUCUU5ejdFw3PbHG9
nkMu1mUGUB42+MP+6UbGF7ZvkMsgIDZhXkjHmF8AcHrak4ew2ojPrORkX7/HiDTW
q67DCCj71crMNAAs4u4bKPbaaoVLEtg+T0ZS+hTUGGQL/XIu+m2njM25u/FuKarr
USQCsS0G7Ejz4R1UdaHG6Ha/TisiqW5Sq/CiKI2kBwEo4A/ddXM9JtVofPHgBn5G
cgqWTnSFw+VYMgIaNSWDtdq4aJ5QOcileUV/QhDrJVy5QZebRiXujTXhjIWHv8+i
WohJ0BTaQ2nXftKd3ZzOVHTLR65sknLQfFU8WdKEzXMpN/3X7kSvL2SGMUoxQB+c
6+HcMfLJjdRqd53KjKmm30waZxuxEjMS2wrKtKTWLLFqBNTpuHjSqMOl6VdBmESe
WEQmuzsJSXTxKcA+1ptEY1ojY8BVD1dMNUs2nXRTNj8efyzFnSb9xcCNBg6xXnGf
sM5FgMT2n69Ogy0QZ4RIoah4VTsUfIvAhakH/X7dFHCzi4BTv25UEHw0Umjolkfc
PvqrC9OJI0sHtjEF7gWGrmkDOa3EgeluEBOR6fPAqQCs9g61LZRmm8JFgRdl67lU
fIYYDep/xiphbzY4xQTg3R+YmFqoUGIdb3qeqZlWo7Fj31WqoNBBKkHpn7jy2HCW
M1+bBma3L6gTf+7DGHQnOa0ma55IrOJcO8jZz7YjNhXuGBkP6LqY7BIwGShbEfE4
/Wpvwu5LwKvpk4VRwxKUm+GfM9kiv39RYRAywpCMQUNSAOWnVI+7cFHFRgZkhIE4
ucMEFOYO+q8B012AtC+fFOaK0eODC1FdlxlOx39EkRN1USbPO+PxX9kkgp+EVxK3
0Ix68iVbrS059hJ/aZXzZVmwmEsCBqWFED0Hj49yu0k8YM/o9ELAvcNdAOUtnM4x
n3u5X1S4N6zTMLjZti0zkmoZ+DgoV0PPn9c637uPYDQMb2h51YzezpVKZM8DgYVm
dprFLviGpi4Gvw8nK+Fkblun1fpo5nPbVEng2fWY5OHql1gHr4iuyxf4SJbJyLBg
Lf/OXfoTwOort1YLtgbWiONMzhbUMlT2v5bN5jMCM2yyZmnCQL74lN04H74gWWGg
MpWgiVcBDzyHOYajDaVFO0mCwFmlGnNJOnPlRwnHGGIxbKZsJDLiTE0Bhf20MH+n
s1hMpaQiuVhT6WgvjEcolYg9/5eOSpE+IjSGBmJRcdjifLQ1tgGDQnnqFWxXw4QP
VTc2vC2oUeTmk2BmR0nOcKtwBj/uiLp1JbyqGhmFE12pHFqIvtLz/gjmesPJOhlD
6hw5UBCPbqe9fCjPoNiA+vkE9Qs9LPwljN5XykGOsocJP2ZoroWpBqeFkQR759oj
XKyrIB5VohOsEENQr9khdlbk2Ona68hR3HLxKj/DJSFhDvY1zjkl9bldjZZ32hIU
raGNIqUQQI1prlX+V2bFf3oVuXNHeOCvJfM0WXtvP6NSzEBddd6lbLeTr0AKZEo1
he9C7+6JBz5dKoPhYEmIPy7vyBSMF8lTdMS0NvwNd0uKxEFFCOWl+9X52WYdSkNG
aesTadOVSoCf5RRYZroZ2xhrGowb0OzjkBaUqn7zyC/P7oYboqNTA4WwAaAUYf+g
uEcIA1EhnzDwFmooc/AtSzBiuIsxHRB9H8Mb/sE0JBOnL4Fj2u3vy5SCqokJYWlU
Ukl3RPO84hEL6NWHDgCCUI3BT3sids3e+E4eLYAQ6vTBP5f3r5b5YbJwyxpskvFX
5OjBhH0RJhXwTxurqIYPj6lzGxg5BaEB8DavBLndfPKisArex+09sEj9RjS08kqD
CjwmhJr+6/Q5C76m8GVkZCCDltf1wTaYebId1Bknvbxhkh/JOmBy5cEodTb/W8fi
d9HDik9PP+I2bRxWuHbaB9yc2par7ufLBna2bC3JhJ6iQOz13oXKYXs8byjH8G/C
30a+9G0etq8t/2+/Xob0iwd1xLq5yZ/1avqnTD0lkIujts+uEnGoXOAWV0JcO9NR
Ha1OY1Q1+zVmqdMaGPvkJzj5LtcmtUaJtOlgu+g7/1T+9awsLZbxMS8lcBr0EdGb
Oa9bp+IHF+LEeUdp4Fr5X5JmZaDJjy6jY6z1Bs3WV9ZFY5uO/qRClbi4ieyQioUq
TWQy4dUWSvX4A+U5dFHP1zuM2NUs0yAs79htJ4aT0qMlvkgPZjzZoqTnh75rDN7t
7XvFZPy7y9ReS6Voy6M7K8tU/FLvm5qlgfe6X1J++sp18hHau9k2ObK2yIywVqJl
rxJJ2FiSCkJC6pkof2N267AbDh+0NA3eYSYWBmaLRgj82EHO8VFcGnVTZifR07+2
viHj2GdlvlgtkxdDLfavFeaH9TdENr1hdXwJZAR6OXgUggyf2eAKN5GffwYmO0K4
r3gxmYNS0Dls6R/WVQCO5zzjEeVOWJB3z+epFArXhrkyz6fA+Nb02WRHAufpl1i9
VdhBTc1N3Eoi/kjqvUrO8E6c1lIUbe2qUUI/1u34Th3rY3G8HgC4yKXFRgS0PjM4
Q4scrXQniMhOVNKXPwBVItuDMmL5D3cXxEX8zhx5GYIsihK048zBV08NAoO2N2c/
AmoLlqOfilDkeROrUJQkT7B67oJmP5z4/b8cbrSf/0Y/2JzHgDBL9fUc7Gc7jmgv
df1MsGExafEmbQEoE9AK3RskwHqf7o0Td8kV5n2py8n4n+REQmXAHq6UJ7xYpv06
EmOlxLrC8GvbwLtkwU+KCJWntC+2b1qtVAoJ9yPJnuD7bo4iBBv5hU1Avl8r0ygB
sCqTrllQYEqxiPdDqH2YE1/jniXim/2xhGWirp0EfmE8zyk8LaY6dCcllNVakfnW
knPDx9Z1aPc1fRb3XmAPuQyW4flgILLWbVgWs55GPkBwS2vIw8/OBwbkmccN5zu0
YGLoAtHGDLSmSGdhCrAiGD78Q5A1ZI1lSyWuDL1fe025Mxm01s70q/RB840Sv5B8
3lCmYcggOGpWuxG7wHk0n9e1BVN++B0JM+cnpQnXDsX15H1zXE04+UXP0p9uv6OX
905fv6pUrZKf1OIGAOUSdJoYkzY/XTGC/AEsnQiMDHPWvEErk9lgxHO9AjS9mN2p
pm+Wt/mKAjclnbpTBOps2G/hgUXYkJMXmZJFKONUswuX1HiXZb1/W2bSsgtgNkUU
C4Zav1HHOmxc2SIII+uXWNegyXse4gBzkt17Eb/qcrGAOKYdzG8T/1Y1t8sfxHCy
DyZNQM8UqEUwMpYxI9M45rncaGLfeUk7EfuorAcer88swaM9lQnTJzDV/CeHhxmE
eUAgGb42EquvIurNtv6CjBOFlRUYrp1fDr+QAvFy4vti3f1X5NGhMyQOP8WOfFlg
16ChIVumnJp3NUp8IPkc96g4QJ9l5LjAb3qMU8KxV8k63NMlBMr2aruyCfzgVoVd
cMRuITaMGh9ZTgjIye/GafTK4WDPNPsplADvDaFPzFL1XXi9I56ZZRSiDsICg4Cp
pPvbk8DrMFyFyNWCrNK/SCIJLPJmox7x1cgFtBzfatCwyF+EISUjWAsOwa1PzgNp
9AP/ndi2SJ/0VELMKAd5T2cCqUSgqWyStR5tW/WvA9WcB6Y2ISNjrU4rhznHtuRs
vBz9O5zCVvkzVxKmKf6m1OLvEDXKi3TCPP6nZeMHV/C4n4Nrs7mRJdIV7xzo5EHX
d5lY15P50OQOMXef8ztbn3DPOoAVWYi2L5k6OvE4NGP0ozhLgww3Fcsge5x4RnRv
EMMj1ajvQKR0cpimkrp8nCsCTdU7IRhZv7NgYHz/LYuhila2rn5L15mU1xOzK7NG
R/kEKZiOkMlnu9su/KjuqIo8CZ9pU/Egwbxba0a7vrGmmjVQjuPbgXhf7rXAtbRL
+rKCfyB5YuaGdV2He2YaISLbqN8kwtHoeFTZapFf4dryX1/Z8zcIIDat/CHq3LSi
2vTEXCSYb7kzfujV4YNeeR+FvuyzBNvEHsbajKtOlIuC1+W8tgwGDvrqJLkUIuxr
CdZylWZBXWajXqcIvwbugiDXqB/ndMqkunPI6G47X0AwFBLbSzapH/als4P6dIPA
v4wE5OkGCAdVx+zmlAnqFsimiIt/W+OVpCbRDN0An0f0Xt+Ph/N4qubhI7OKCkD8
NgM6tjjjlJN5++bHTjhbhc76iSD2rh4DhE8NyyMIwjjAfFv0AwmvacVGC5lFFBUZ
6gxTP5tqIGKigxAb1QupOINdsA+ASE74eteB9oKoF9hHStsAdwRFUNbIZj2vQGUJ
0dXB/nBfIfMNmzWDuaAW7CSQtDO+MWEqKEDVMKECIKwh/gE106/bf70t2sDxPkNk
SbuVqkIjOFylFgBl1NX5KmW175T1UMhzhzWyuBFaJjM/0tAEkALIowgC77ySplFg
uC4Lc7UTGCYlWuZ9p4/Ys6SrmBIJGcRR1P7iBmsVWXjvWWJqDoKC8T0xhu32gAMj
qXP4Pmzf7HjjmVD9vRe4mFyh0yL0byRrpwWUlbn6MQ3DkA8TXOa4gLfUINTX4eye
Ry279vixCQdK4Lb+3SHTu1i6owzkdLiquvT/cPttCPBJYIaJfY7a3pNrLVXnrvKo
2l2IyoReso0Pm8OFRoYnoRtUDa0AXsU0IhW59HbCa5TA0Rw0gPf+jgD+LaMwLByG
QYe1gy1Q+sr3VeoLbcQ+1Ux6jDIP/+3zrhNG7GYtEx/mgc3W3yYGm/2dsuMX3CsU
sNmeepio1sBItvdB5VucRCssy73CMjFoTt81yGSXgQMXVpmwVim/Ksh4IU3GUaRj
haqlbJS+8x8tRoHlh1buYNfEaXCqafLLQm5l3L+tQbNCdi8ZAyYHHJ5j1itXCtU9
ZMmYOM0zKOh4v6lyFcVEAycrGyKKn1ClwGsRiEg+8mxowF3UGOaHJsMxcFd0XmSh
9B6SSGHDe/AKCATQPekIhtRWbA33yXXv9h5EPIOls56y9z59qjSAgp3RuPR91KQV
rkncxxceRJS3WECPODO0PtsNLs2j6LzNdSJh17L4Puap/5upWDNxUvRFjUkMsI2z
iWJy9KQMUaKOwFkILfrywY8MQNMolz3BZGSM0DSuhroiIjXUb/PzQzoQ8KAWC1NT
n30vBAqI76EOOd2PGkIiDQPtVVsZ4Q4+UG4Zng8ymEjrTINrxmRkOelyA7gF5ypk
nBjZZxkOAh1HuvfRaEn9FW8HSg8tkH/miMO8pCophPswmi08aRBYqLKjIZhn5Tfs
3UOqfQVt0E5tpnV02BQ7AkzNd9yEe3CljjuBJI/ZJy65itFVyJZ7issbLiqLljLv
ELx62FQgW1Hqb1vXn4l8RWY9buPXFzlj4kZMK0XPlz5zsMscatH5twAbPXrmW1fy
FfnnPYMD9+iGBwxWX5xprtVKo/NYRgMTeLjt8eFKawmJqxCxXV8KnkpvIQ0ha2U4
6pqRK5m4/BwhQEew71EqaALdNt0SoTlnKLFBkKOZMQ5V0U7L2fa7ps2QSBfa+cDw
xGHKGm3Ek1AH0N0FqiUiBPV5Zhj2gPhcRvtzGBkuF/yZ+I+WU2XcAe00SSi1eTwP
4ByGuHxqA6ugP7w8GNV8dqS9Two4dA47q3Lh8dyzGb9np4mtCqMMW3GqKgJ6CSB9
V4ApyEyF+x5oM73h1vI+fU9tEM4v8ZpKsngJREKhKxMWjq6ctD93Flw9kVPadbev
rynqk5B+8yE2ZHyPS494QrJ/nsER9p/Tnr09R8xEx3li45HYeqBUYKgV52dz5MFt
Txeuq78dkbTBoXcs/PpO2iz8i/KGgK4C4hkeoMN5YuTa4DYuqvZIaZ/frSexY1JI
8dybVCN1eHv9U4urc+eA/m4lf8d9pvzp4gzovnM3muSyU5ySnIq005FFE8CJ5Oyb
pNfj3an1ipVkHV0cqE15iAo5+WekTWkRYTjcrBoboUrx1oMKSdyJHM59W5UtOxT+
MLhlXh67W2ul3m7I7dTjru5tSDozeDwCtI+AKmRoEgiFGZcG/sQ6nVDXxi0n79vk
FwO/O/n5prepx68CAZfZscTUuaxUuhxdJ+tDFrH/ZI98w+Pua/WpqkCiltg+ehku
4kUEi1RyO4TUV1vBzdxsc34EVQMqe7q5mHuAjGQmd+EsHI+RO4PkDrOVJcMFbXIk
9/gb9aj6Z1wVpqnGxI9y8+XAvmnt7nemH+nAT58gCTdU4p9n0j/N9GiymdDU8l8k
7KwblwCkz6lDBANzLXjuxoZNXc+/1dJT6+uZZi1EneOrWzx2NLaixfVcJ6eoxs2p
UQkJQkY/zOpkOaZSfH4emoaz2dVE8VSllIaX+i/x4YKfgPwEU95LpSwSs/vJpZTD
pIzbXUO42zqsqyuK9VMbv2RzVS214EKiqLU/hxGRFNJd+bxaH69Zr4B+CkQfhjr2
q4wOU9LaCSHb8t0pjNBEZgMR5AnGpG60FA3y8qMEkyshkrj60ks47lOQAzQEPrUP
g5fHh92UZmRaPw2Lw8En+iS8Lox9dzCKOKkYMom10masmLshjf7y5kpGucyeJNTi
gG8eeczEebuYs6z/a1OcfZ7eh16rZpL7yqiOyko8gxC7vPrAmz6unVxiAfB2a2i1
zmV7bPllmHJP+ftoYllAHu6byqX052ekQPevErrFDSVpDy3XW73QgUieTU5hXZ74
TQyLhV2Qhp+R3Yc0uG/ak4oQ3uue2DW1e7TOUssiYibXQf0lOqzexGLG1nBAtiSo
lBpyai2W3jy8NC2Q/+d3VTKuvr+qYQW/kf46sKoSWAHeEVfusvQVLgSCmPHLzDB3
wGNT5fYFZpw26gtwPSUg16iUPCPzaFvPQx4M9tso+FAksDuk3EyuAWU87W3+1/xe
6sQshH5BI0B+zAutLPsuUMYvKGD4zr7b7TztYCyRm8xSboVufMB3P4OGnW94o4Es
26PQ+nWpJfoNF9+g9pt9t30BqTiR1YXGdUM8cglQGTRA/nf0WKGiT9Wng3akVr29
paNJ5xx17EPlZyoMosiFJCWTm1BCqypY7uGHbuEk4MSOfiUMsmSzxPAoAAsw24mw
CBdqLWvv8Z+OqfKFJt6mzlxSmKxdSVLSwGGzKwcSIfvNJzAkhd1WN+6NJi7U+xBN
KW3+Fm5NCnlJQkkr54E2hmP1K8IsJbsTYXrhP06shpSivmGRcK7L3kc3vzKFbrFb
pPmofEfteI08lyc6Lu57GlcoPewFWlXhJXpUEpEvgK2ULmsGsIYYWMyI+upjPXam
0SdgnjvXyuxzguLmKypngzDVdrdMJ7SXEIlIBP88DJUyBsK5CJee4ALOAlOqSGm+
bqPj6Xz0SNHN2tYxW7SCh9KTiNRMav2b8ISrSfL6uNtrmWSu2QS6vP2px58lRgPa
S2LzfSnCN3P/QTI8INXwNb1U62HmKaTVu7nU6BWJVNBbWyTPcM7pXfsiJh/E0zp8
xvXd+9b5EMwX1/fDVdXLxdLUYDx59g/gQFGUpRdk2sWblT/Gx9A1mgy8dlP2afE1
NMAgEsPfDMarIzBaRmfyCL9BCjJe9paATm3obOFFGZZdFvDU+EbFo47kAphpkgIE
VYpWyKANvO6ru9xcnpZcFSIEZlHRKNZYuGlFhcRfkFx4SYzkD0n5IeFqsuRlhkcn
jzBOLOB60yy1AD+Uj+lKTfQDyY3g3jjKDYM4mA83VYR+KoaX/oVR6ta7aza51XF+
etyWMgsVxltKMjWH5CeK0RymE2axngIjJpjlMte3HoeN9Zzp0lrvcDZqXTn55gut
0imLvtio6UpnRF9iCXOaMCig6TPpsxu+WcOxrlESLT143BpyDEnqDQGaoygq2paR
1fPk9zgFdfU+mwiQcoh/8t35Akli6gCnZTFsfh2a5HvbygVwRL0LJVb+DadkPmOT
Z5lP8xrMEkPm+8PvPM2F6MlOhJSBLw9Y9GOBP+chZHQqvTAYWHSXOBG6cBatNBzk
CsSF6TpKK95TlcUhYpK/yywAVMHYq2aDUkqg5hL7KvLVxOzUvH9Hp900ApVOA68Z
pKXI1bFRTICaB7+gk1z9KLmNApQIzGkFwUZw2zhLXQcuEGoMd7tKGoEMrhBQTPQh
twDH/eWgVMRJ+baZFPSjlE8LrEVBSYWrE9UZ9BQ49A6vd1maukUQUFHNXqUCByC4
lHdPM7HB7Pk349N2MtWnq17b1Qgco+4EUXqUA0AvsLSHYk80O6+FkJpiFXDw2SHN
Wp6vk/yLREiEgId3fRVonPUqeSQ3fcDYgei57nvUGCrQMYBSxwqziZVjK2vze6WU
elS3DpE+0fVfDS+Fm4wJQHfpR1WtfC3B33bQUheU90/gJMld6Mv0/7hefZNMNZNe
fiaXL6dF5Bh3nYWJh44FS36quPPRzGCmInHRobKKEpfOHiKp3urxEN1GIKtFwKQ5
jLg550WWZX4bGcPR5ovh7W1/ddQTYu1H5c4NkiQkOuNZ+RjYPdzeEtoGSCW1Fsrv
xOvBZ948d2n90nyj7bJ5ZlOejRqI+V7jUdmgjE+t6rOp0P4Nah+j60p7JMaZ/b0E
CZrpLPDUAN8esiUx70HBjsZcsbbjkePnM+DA343EhZsyoD4Zza9tSqTvycx1BcjR
CXWGneMIyM+ZAiatCJlKS6AFf7/lRw7A/XsX5BGUwZos6DYemQg10eBVhCKEQH4h
wviOqSNAWTUfg6HdsrP1Wnx4Xi52j74m8CogWrKh/791Y8w7aBL6n91/G1f8oGb5
S/0V56+2aqeDMK86tZumwZPAMNYc6Nc08sKJmAUymCRdpWYbZMIYOnROICWUTBEQ
tW7XghZagN+k3EY1pHXghgukzv09/BcjSEAbJNVp2i3ks+Tvj6Twx7SDmzNydSnM
KqW70koMh8msJzd660n2FY3dghUkFZiuAQvnMqaTfG1oGYoMnb0Pd1mSrNEQqJf3
/uz5dT573eaCLemxvY4XWINItF0ow8Qd1Zqk+MVR1LHTcYTFwXrwX2cgzioYr8bi
w8FO1nbpChCdKxOU4oIjXkHpgmjo9PtJLFm+g5RH1xKUy8qFmYExULTyEeYEtZjh
x81NvK+DtniHrl4dVwy0QsA8BFhuD8T+OcFOgkBL9l6mOzj2Nw9iiJ+SIJ1ZL4gl
yXgVrbExKav9UwVjR38azxzMPW+U7joNSIjtTg/eN561PyqI59DkY8RPlcRbJgRZ
iDZLoNK8eT/iVYKf6kt3KZNfv01aK33LzY5EUHeje4K/964SYq3ldTsvMrh45KMk
c8ahUWrB5fzrKr9/IGmjmLhLLMJrOIkpw2h3AxlvkZ4SgOzE2b1E3oKxcPzSvyFk
tI0A7Roo2P5/nQVLIIaFn+YA8itixxNHc3Ds3cPyYFMqW31/XFoGyHybQNjofCo1
FB3nlp8E+7IyGOv0U7w3cQFkm1+nh3NluSq0ldSS+QL2g+dIb9RkjNdvRvEzRh4a
gE+FHMxC2YKd22lnAZVZXs2edk1mEirl1O3NGY6CcWpV7YwnKgWhvNJPfWRF14ud
kzbWH0faY5I4VBcgCD5SseJrU+LUK8KVB+C2tdIjMR82CCgOZear9R/vtr3NQ3mt
UMVgvZ6eO89Pkt02wDH0qXuKod6fDMrYq75Pddm2qEju0YTtpDCzy8JQupOQknH0
H4vm6PMDx4WKKwqF9VSWBk8ryjcID8eA5B4v/lVYGf39CwTGDUBEdhWNzmgsf4no
j0yBOS3NuBdIR2avpr2Xfisj/0ObhZXP53n8Rbh7WV5lUd3QSIhx905u9m5InKG6
dbfArvMwCcE7lnwK3mAAV+9PLwyUmJVIM+DF4OA6CBlmEXBm/R5HZYTRDVBFteut
o1fdUqkefYrKVV0BQ2BG33+aQtV/G4tZO8wlzAPnAxtn53IvIxDTeajDxW3yFa64
/ceY17OLv7y7igpF4aadBy91e+n6hdK91r4NbK4EYZd8gC/FCXifb2em0aoWlzQZ
5G6yzNvOSMbb6yYQHPCErCDJC0/tam1q7s2129USAjWsNR/9EygFNA/NjhFFCu23
9Mjen93CpzGvXPxXDsdMTyzjkYGsdhX/1WlZw91JljJQu+EcY4SNVGvmDVWrfTJI
XHeKHWyrvmR3q8d+Gv3A9K5uahjs6NCL2lyZGsh/LMbOe1WattkFz54X9aXo4bWQ
3/PN4QBMh47y0xillCPLNjbcit9i4USPb4NEgYLFRL1gQFjhsfxyzihyVWFsTH5f
+FGj9WOCg7lonqnf9J7YM/qEXihRcy8NMeEN4VWIjK1f4zPqCFNmfZA/lYe0jfHx
EiXohQ+ncCWaK118oDoG0lJ6pA0M6yhxlNMcokzjxLZ1oAKDS8G3uL9RrvGnoSLm
OOMYWkmCXKl1o2//ZxENZL5OpIVmPQcqlT0GSt4JR7EZmlf82LCMvuGPPppMd6Fy
uVJRNLFGFMZFbqdIZ6f8Y/pfXOKpFNC/tQg32VjbOt8rjOrg3oUYFXuxA3geS1WV
iUcX/GUdyHXzxXSFkP+1gI/WWjn+6jXgvCmXWjwaWrowCA4M22jjkAu3iUoKtImQ
B4EXdovVWbFNazB7P7exWsBtqIu+UG5cpB+Fd/48r+6hBKJR/Z6b+EyrWsbndG2t
PoH7FTkqVjeh1SXjal2B5uMpPFwINapY6+pg+jnygLfxvBow8aC/efh81GT2d+JR
K7JKVwFEIQIMRYNVjzGRzoqjTO76k9uL8LKFwFQssX54cwom1cKl+DFgWu9wPX47
bWlNs5/CB8GRl0TPREVlOQY9LTpJjsy/if/1EN/lHIiFPWG/TZkqnrDJwc50Y01t
y62E01hQvqcBsNYgO9i1gQThdqW5JyeIw8hYlbLH8G1N8uIAYOo5TKTT9Ikyup7x
oui2X7xrSaxojsACpgnlLfz6rDPmxnAdHEJeLlXaktt2xbrSu+OYhI6QdP/ituhX
e6ROB6xXkIOZAS6+nYHkdW98u/l57Uz1IbdX3IvDFOuFDfcNwtl1iqeO1NF42Xpo
eKS7yp4KJ11nCy0HMnFwYSfN6m5QCEybxgjuNBolH5vcnSkOFRP6vOiTctBazknc
a9/qjUmuWp1VoRiM1jO/zWBV5ykjZAJyzrupPM3YMenIHRs3AkDsyWwoTq6998jz
0jIU0rHCuLnlQPfyuE8IwVp9LqFXXuGgq35wnFVXPraNX2Z93TsMRaJLz51pNhi6
Er3h3/iRBIDc51PTzF/gOUIFlArQQHm0VJq7H6xkCH+2M7SNNJvUz7L1weh5oOPM
mhEZGdkthbAVAetAetdwLOEo9JZ9KIf72jArRFhP6vkfDFXCDMwILT3BOS19IL1r
m2U7R7OVWAjVHQOiVDmgMQ90Phm35YSL6I8E5YlfA/jPmMUCUioXlnRNLneG4lMg
9+c/qbkOPokBFTAOhv+NfTjpXErRLDZmKj+g3ZWprI1lM0+o/RDUt1oe/t2lWyZF
OIuWvYEHJwN2IgsP3oXR28DS64kIk1aL51CiNtH+zTL7UDOW4YiF6vgTV6oWPk+0
NBY/mE5XXJlyb+9xuAr+9HSfsdFifnq3kon0XmbKrn2ka1wMfVGsWsUrZSsPknJV
U7dT0Rc3GkHquxVqFkp6jw/slDBZxoMLa1NM3GfXNnTD4Oza4OxuplkjxeMog7C1
ou9/BFUUXp7wFrBt6LO5A/SHrH/W8ok4+4IUmqPK2GChRTY/X4nygqWt9SLJQPOU
wfmmXmxtx75vxtQi9nPpprt5qy407HAYkFhXhjLi97vg00CqQg/7ju1jqBtLAU7M
9DKOxbVccuWx4fJVLbte+5tnr8KQ5EKMLcDmBVRvLJWcPvILxWDqs0geELa2tmfj
F5K8NR4Cl71wFv6YM6kDLKhm6QbpFLxUS4vqvyqsvtxI8r/MhJMoF/ZzWRdv2Khj
DllAxQCa4Ikg0BHfIGtIHtFLN7/L48QtlNhshPnKPp4cIqVRF/4AQFkO7ikzSHeZ
O2qGdEnRCLjWCXbOY7j6UYlFtQfHC4fZoXQKxLpOLziXfAVrl7msfW8kDA7A6v9z
RqHY8BeHyULj0ifdrvIOqOUoX9TFovgKadSeWDSSAbCrzilTl59OpC3oNiLxBqcH
6NOX7kI7ldzH1GxMlTWpQD1DTixh+NYM39IrVbJ7UAcMSe82tLdaJ30xMKJqFCkL
/ge8pxAoKj5cSsaVM9t4bcaFZ+mxkv2V6b580uwgznuFtGi3DSToDrOeYiXs/eBc
5mCcPCm4psg4dI873BccSoPxpudRi26cA1ExmveNXFdjKgvxmoarw5Lhc7FmrLX0
hbkLatM9L6bJxeyejO83wT/oXfqL2u7NfAMPoQI9moyAr6oL09446ytNWkEt3sNi
q1323uNqGhB/1ao9jNA+k3bKs17tzO3WgTSksX+GAvrYRXwK3t6oz/SjkzE8hpu7
hfn+Glil1D/A1OLEjnwcUuDf4pNuXsuR/KSzgVf23+EQhZZXdXVowKHBoE6vgTF6
jsSadIqu1BTywn/kwyXgP4E2v3RVY50ohJI2q4ctrhPAolGGKV3pRsKLhv2UEnPp
PJo5tHSqQBAM/+kcPCmBO6OT5lcCvy5/CgyKtHodn3pGFrBvxBu/z+JAd/H2HvQI
ZrNeu28VGDWuamRfBtBlBixKp5EMgK/2CGpcJS3E7y8rPgraTAGc+8EpZtPbDhP7
BrofIK6WeepZP8c1bbAq2BoEdkFe80eYbXjLjXQWsx7pyKOoqXGlIzd8PnwIiGBE
HZh/oF/PT/Ty94JvqmDk9exFCb/2aGuOsCJ6Hnkdg21Tp4J1NvQbb195xx/8Jy5c
+0OUigZIIS0LlS7FaIZM8zIMoLBJT2/X5lnzB4XyvEu4yJNMH1jUKfgZpg98qEo7
qzYjGle8QW+pJf3czwG0kSaY2lkgM/xwsh3l23v/4MfSZRnv8kvvoQISBVFGHJjP
8wa5rEv1AuL7fMktRs63aZ5ndpQHeJ+ehmL7EQLrFUXVLD/F9YQ9+3RG3JdbDcPf
pxcjUwwu/wJqfPEarNhPTee6QdGHD35X8gvRVzAeayTzuEdXUF+Ra0qbuTKaut1Z
eMwW2v+48K8S5fylRQrjRmjYlAd6pNoVJGCmRC4gzhIk0Zi3Xnf2Xc11ugKw5Tf/
xZd2jm7aJcRzVaAvN272HTypzrW+uhMbnPOaI1GaSKkbYHCfovZG/YQt+vtFw5tR
lDjPly3VQGCM+aMR6nEYkzgAARIEG/u1U862pQoXkfFqjfn8UAzCuX8cak/pvYaR
refgEA4Ort0upFqa7unIWjuMb4NOV0Zg6Xp3C0/V+741m1CxAIfMBFWYrmDiqPbr
CGaF7eKAmDBIRpmA514q0SwfU5kehSw9yrvwL3dokZuAb/Upzv1RNimnNAZcUb8f
9kyMPrXDq6MMchT0ppEgnwouoM9b111OYFkuMJehcDXQqI/o2kYVK0VitmHR88cd
GFA/3Kf1AemIdxixTYbLx7SCN26tSfgbf/oQuKP9XGMbYMdCfUJ8wZNrfBZYxtyk
cuz5eMi/L2dHJzIcfK2gZ3gfLarxJj+T2DyxYNMn2a/vuRt60sijlJoqettoOess
NDpS5w9nXBPnh1dTzZiMgGCKIoarFkbXr3ouZEKX8gkHta+mkastqeVxIOG/EUiY
RwVlX1RzFx54jf5kReWANNTakNka8SwkoJfMgwAuZsV7OrnVSI8ocSVW6xTw8pZj
f0Ivpjt+1/9YFavdcJtRW1IdDcZySZ1XOI97QHN2iivffpId5eKwYEGTZq+/mKsu
Q9YHkpeOCLguFidWAFb9btyraY/VhJwXD+R2kfxfTT6/DrxVGHuPHrqYIZHso8Bj
2obIebne6x28YEkZMJCt57Sjn1S3cYdpcI1KsKf+LpWJOWPvEQCWkJmeBYmCy10o
8qZMrZXP9+YvoI4MrrEO1i2tSyMvse97lHBhiLpZBhN82FKK968csgcI/RjBnWZi
IR4elYACG405zmQHz5okOmJBOheqF8xZ9lUv7ijIntpOKv+ZYE3bgnId0DSChZaV
fiYk7N+L/Zz1B2DFivT4hQX9uzGrtfbo93LmFQv4G6wWZwmyysQGhjomTn2UlH2l
pVz3ShV4q115KyCW520/luJOXSlYWkK2g6b1BeR+Hd6PLrF8abepvwpqIVsXRi/e
5s0vczOr6rAXDK0eklvvL5tr/CyH2e9qnKszEU+roFJatmlY9A2Hxx1/29umYeU7
UG42550a2irzB+b58USvyC5vowWMX5/3rNR8do5ZMlEDV/ylXijWy4tWY/TeCf1g
SRzImWpipcZoAiZWXptHOZwajmhWtpXa1NCiFt1BQSScYrDIaakGm5pA0HYDXJxZ
Dwv1p8CVyPtOEIZlOB8xg6Dn+6EXnvuMtSSHPy2JALIh1VtgUeY9Ph8yB/x1asKb
N+9yjbNV2RxDsG+Cd7orugy6o7CV4nnVAMlNSGN9f7DQyl7QFruQ2zCCi3kR8BVu
opjlS+sqcGqEO0uX8AsrbjQkmpB6LeocRg2rMh9aCy5jQ5trC6a+aSZKUmSjB19v
JFaPetNadC2AZ6891p932zeQljS8WuqQ9gh45sKxOtMi4NlbL/LYUVnCN2OAWNej
WfiU5YD9aZyenIN+Ri/twom8zW+/jYBlVuuaEkJGt5wjsQnYY5bLNxIWLWMLPFYQ
Pflf13XZ9WZq3duwX7ujSVrsKf3mLKHc21VQu3oKA1/Mw9vYyUndPXngmq4Fw16U
tsPF4CTHLUdPPqb6dHwaQMu8KOFBEwQEQGSJPs2Pw2I0E6GcYPIuEe6LinH6b95R
XdyHgl9BG3KTu61e1s/PYs5lFsFTIX2G34WuSc6dgO8O+b8psfBA35fqqWUhqSI6
hA0yxb99xTBFCScuMJhwDfcDoSl1Sb+wbP7jvWbur6GgYOGbDlk3ss1Dc0jYOSys
h/+Pc1LLE0wHRcUHzOhP8ElAE4UhJuZ2z5wp2V6sT0dQNWps4DdYff/D5u/hxBJ8
WnodJpH0OqCcVhe8EWy1DZ0Z6IvxO0B+lfb8a2IOtPbRPbNSn5BA4NbGOyFMS8Mk
O3Ri0xenTng3SPU5dYQ+JYHLu47cM3lYwNhOuaNtxcomFrTc42MijDGM6SbPngSI
vc+Ev83DY0IpaMy0M4vUhA75yxTPi30v+Pg9xerOUjxBPTLS4/aYkTMzdSS8ejxZ
RWEWzZwXl63UDCCBWqfb67TktqMcMyJvxry/2NXqjabvkyfedPG7CuvTxDvE1ZYy
y0TO/Re7p4KamVJpERD29JuNGOJ1cG7tVJzGKBdNhsgmaFvjjWZcsU4U+3PGmJ/B
TZ6LXQMjuargtiWtubFN5p93tAmOhg0G4jXcC8PWMt/eWeUro7PBj5D4izqzwDfy
FztSG8LzZKTCryMz5Hzv60PVHmYWEoSq/dZeZrD4tM833kJv7cfG070ZWb30obd0
XTG3+CZCuHXvaCMxzI07XehNGQJH9umAZl1+8RLCzPu696zP2zXjfnlPfyjcDUoG
NTflT9zpLDOqTzNlO+NV53EaS6xtRMXuwG3P4MKMGBX824V+UCe/dzuJnZfcorv6
uXwNvZLM47cDlEG4dDesbHhlS1wbjAviHZULp+ZpduHS5pWTSRz9yzrJwRedWppH
IkpPSw1EKLIw36PYDBUNUPCSAFlwUhVpsqEQY3gpO2QOMgi6LE55PJoAnMBtsMZ1
7LWD+oMwLtCH/ZNs0Yq/L9OgBJ4/jC9zRpYN7XYweGXjdjs7vwjtwmtYm8OHw7IU
FmIPgylRugBuvDrn/yizbfSQjlEpoM5hkW3BbHpd0fm8qzlaRQIcLFWFFeZ38qFn
ynyB8u2QDDf9y/L7rfOU7nwYVs1359ODrMdUMra/EXqvI3zWfixl8oZHaBtutjNX
gdmw0eE7Flzp5DL7g2OsWkZJQMa2FykvbBsAiY1cyYIH4BSi2mCBcy0HT5nJXS0U
YOt+OPhK9I4YiWyP9BQyzOfagFuW59g9EYygNxcX3FGtTZXO1puz0LpsDUJvOS+W
2qCUV9vRpPRR/vDjrReG+te9iCld3pt3HNrhpwoxp0FfsIEJJ5LEj0e4zQUTjX9Z
B9qApcmfWWydotfBAvLIrxGVAFGXolN70N4CqCTIi9o4SZQTQlQ/sC29BP39gnaf
Amm0clx/1uB69HqICrqMJfy4zdEI0hZXs0tWWteeKU0cBQ7tAB1/nziaaKRm99Tf
7yRZNFzwDdP2v3nctjGfozBsrBqGszCbXuhCnJ4pT0JddO3ZDXgotCWBCDrIpV2Q
pbfo9NAOl6qpsThN936bKp5fj5LT2FDWMDkQeUtB2wL7XczpMKolDCg4gSfZkdWi
tcF7pKj6jwovBI/FX9U1fP34R00Noknch6HwDOA412+M1jVjopFhesHU8alj2gFG
EEL40oJ3YZqkTooob+UMGpPw/Amk8+JHJiG8af9ODiRKEIjbP0ogj8IIuq8DDJGo
og0IG7g1GGFPSMGpW0LxETfuFkur/YWNygb7Ljy0RiU00pJqCyu5TuFfb1kSqVD3
Z0zdawDjdHWSv6iavbRenGmptLchoU03j+5exlzQELnCBKkSY7ACDsrWFy8YDyXq
GQzHGhy94Z4eoZPfIvDZ5FY2GhjOOJcblDEbqPHcNJMfaEU8sLWedzQOwWWVOk7f
pDYD7xBQJgn2em2HMviB+k0uLxi4Iwf5PKQEPdxG1Q0dIGHPVAY6m4r0qYFQLdwC
DlF7u89xZyueehRDUNbKbdKlgD4rX8UwNh6R0fmco/MMaE6YIS8huKmK+iloxPF7
/+zDUruFnSuInpj8+Xz1X8n/ic5WAEkRkXlpDkDDbG8osfTVeG4B2MzqeTdO9279
Yp4QM3AuvnamtOGIkua1RZxB6pTbJeK8C9sz/hnJJ+7GzbYrJEHqfWujfkbeEf3h
l7Zr4mjgdEmu8cKIwiX/6TNqKmf5OB75p1a5LQGI8jMjrdUhBfLWE8VtkPx4oU0m
jOkNJ4/l0wtROcgRski84NcQUQZQLojvT6YKycogoZFtjHgh2KisEy4FFmjWY3vD
Chh8MpMz+a8/JRQNKPRF87YUzrwhbzk0EPHdO3sBldCnNkVTEaaY2djpSMQ0qHPH
9dmLxBO0xXt6uIsFxN2MWuSQMQAS4MRwwkzb0CYkkpQYmjyGep6mY9VdPHfaAC7+
EZ87huq0pMwWJ9RmJyz5yShtyNKjHFdICZhzbNqY8Al1C15NHsNt4RVWGazkwW7Z
As5OowG7GE0GKN0WKwApDKOU0/TFNWQkGjK4OQRfAAraKXtJyQfDgbsb0hS7mtJ2
YmY23rUVKnHQunYYEnO164/C05m40zb1dXdapHTd2S4pHc8L3dy1Mgshi/RIhNYd
w85LGOejHgSPwTx4yBzI0gDx5k3mzHByYREaGfNbcYTyDhiwW6SE5LrGFcEPKN4Y
+XxCX2q0x1qnLH+GTDPega4c2uWuPDnSU3OneeRXlaRqClFlnBTgkgzs0H+usr2v
MM0HkNtUSG1lUe09KWplJmp6gKU0AeveDE2HHVPeat2iWzUuLEQjRtgwQlk2d9tg
puDIRVV3z8e0at849HK3F1inDOctuVM+10qIyX1OXpJlDTJms/37cEpTFHawy+5R
qf7KA7qtlPMkAWTuLhA6Ff1YWVZSOhpJIa4zfbUjOjBQ7hap3vMIvKmymQ/Tw8dy
tA3phw4FDsBC0E0FVOQMnv0q//qJyXX+MU6SGcHFFy/V0oGjgFA6vPvgnkxpOIIi
6lLwCiRGhiviw9CAVtgPrN1zyzFgeMKBii8x6c4v42MH9RI3+LiggK8jN7rpUqp3
tmOa54+deQOYRpyeTNFqPGIIiaZCetw4xEy95cnq/+XVQckWs4JyRONIUn/sG3zM
EZs2LnBKVm/gmgdIEUvQtrQ+NuM0KzFlL4wyn6YmWGxA4Hk6SC1w0NpUHPsW6OMi
3WJ3EtbLaV45h/4dqAWes1XddnmrbNymVG3WVcwg8W7kdYcfcV2hVbTGRYEZFAuG
+3XB6I1EReREwZYHEG5dgbgdnUT/eSt+8V2MNlkfnDP1kRPrstF1motS9+W4nRoc
7ahfhkdDWp8YVx+XkgQPnsa1yPfVkIQSI+3yKivwDMtj0eAGBMquUqy0YROMRfpv
VJHMVVr8h7y0soacZVnSToeXOLYPmvkEyLY9AmFkCfUHdDRTdXheVN7LKwu6I8og
DWTsU8oV6hd/0NHl7fiPCE0sMdwKlgY09BDJo0++T8C4ssfc2A3LhjyVitP9cOu1
+cZsQ36q4X/siK/B84ldSMnX5AQ2e5VaI3n9IARn3DeGrhY9GcbJosgItv2qCVG7
U8vKRd5PG0DuHVV4h6qoA27m0pEF5sUr3vbQnEMZ4JAVN8KGeEcyNrdNLtZe5Wvo
nvQcWS9xmZ/2+zfmFTTnu9WSRGb6/N1j/XTIdkDooFzeGfkKq5RZZdRewkufNNrE
JPqC1yRWiOzgqQDAz2816c5BWswWRjc7Oh+xlzKJOQ/RJoyQwnB1DxNd9pkUll7u
q+6rbGJGSKVGlZs3cq8iB1nUXjTR4DnH4qGXbcZbkuB/gM7fl1vzs5Ql6+kTG7Ab
0HGpasNnE+fgkwd9iU4CWdBjUAhKxlzabpkKfa+YNpJlRfVV018orytLfWaTLiWe
szyhXDm6IluyADawEfKYgUT8Ers552/cE5Q7jx1n95z+2eIgeDLcO4E7IaprDjtU
jSIbueXku0Hv/iaN1vADoEkA1EK/3mqqeqCiQ+CetYphFyBXzRAcbhD3TC4fXMyO
kdBImuMXUbnE6QjhuQIKOiIJV8pKMYu6b4NNL9T+iv0n3XAzqE7fohU7yYKJlnsg
XJywkKrkHKOY71peog3CQfZkEzTkvC+MH2mJ6AbCGB/mnNgvHdVgXtJ67RL/cYzb
VCRnkit/jnDNC1RPdzrlf125N2vgG2nWw1lyvMGpsAnMGWf3nQ0HpnYbwnDhVJ9l
7Jmcg7WKQcoEfMVtMnXa8GSNB/I1/nJkyMf73wPEW7hi3qwJ/SaAlUxT2zi18O2Q
Yi/1sqg/IeHM72oS7TvEOL4+Msb58FeldAOM0ozh7zi/7zI3CbPAG9pemPPjm6sr
BJhxEXvEpeM11dfr1h1i2L+UPdidsGlt1cvpIddBPNQ+qGTUjBSENm9dTy2x67aJ
PVvrstKTvSFzm5dECERHCg0GGY4wBQuhX6joGveBH1naxOuXDxET74joRIsalU8h
zYlyM8tLzfs44lEWtt9Ajl9Al7gObYnrCL8+yOF57OGiCv4LLXxgY0mg5/id30qj
eV9Pb2r6vLlVlYQMAjE+6lR2lIMPeRE+f9sVukGHjWB7oWkaAJh2In0FPwM0prsz
j9ketbGyVEA78HkeO/fzRYbHXAxfBiQO3B+R1yObz0QlNPA4/JFRKsF4SC5yHUkU
OyBXxECjPvr0eC1zrc1BuX6n9+FtXq9vyALYZ8sfS5/XS/3Aj3bFdXxOUmHAYPj5
soikyTcsQxRMQJena5woAFNlruBdGfr0Vo8aQap1Mx2aHU6h9UUtnIa8gLmBjp/f
wRXSuDEAk4rIVdJ+XrOjr92E+t/KHsdLbtmO0qCuQ+NCewVzLs8p28U0G1mjPcm6
qce8Ak/ph8jjNKL6X+Y1qUvxuceXj6X/mkfz8HIodaxGKBddjD0pmMc5PzugHjvV
V0yysB91qMQvASd/rEF0r2fdOv3DdRtDbulNYn8K/U5RJNADD04T7qcl5dt67dvK
cMbaVDmRBfX3t/FxfMzg0QsVW0XjmEI6u8jpKfPuhqdMbXPzwF8ga138yuhqZRO9
5jLw3HABAocfPvCs1T2YrGCkF6KDjlrZhbd6xIOBtq61HQtk7mPdtko8HRxFIq57
CAAhAm0Vg9H5Z/ESg9hbefm7dENug2KBbS5vr6jbLoTG/t9WVD/IjNzaNItVXiyG
DKUlDNThwBfoNaYWR4XQ8RnGTzygWGCp2WID3dTtwSpe81E0yTseI/T4f1SsKR55
sNCpyPTqDhi9QXIR6ByvTtPv1kWin5ITeppxy1jZbz53Ezvvb5GoJE7q2i1g+PM6
h4u8zp5If7dLMQHmuIhu82pvvN3Ehwf5T1K1emO8PWRHmaiMbg6jsgzzliE/vz2b
ofHhYAg0/SHVlSSMPTBP/WLcoVR36yXfE/4v05yVBrlIeZo+HmbJp9Xl0j/GrPTO
TN23rWfKGQxysW5SNSqxeNn294osS4J5Ggcv4L93JOvZ06aDX0RUTFFRXfytB+9A
lQD9HEITVcNMyRB0xjq1npEUZEe3JJ4hSww09imvuME82MQz2Ype5uE0FBk+3KLA
WLAFVMtNdQJGCfCeOpqsKqg39u0g1AYrLkym+aSUkCvsdDRHGHWAHkX4AYBF/apZ
LyeuwvNp6tRZkNXdlH95v9HMixutk3S0O2X/9Zieia4flGBC2A1vBGv5wN4Zag1w
snjxVevU5Jt8OuI7vOnDx74hnirbR2X2e5vGqtmE6SthvXHNRfq/YYpkQGxM4PAI
SPJAg/3Ok0Z/D/1QSFDlROR70uGI9BESg7hnfrb6ikjqUFECeZEZBHwLm9lrZ16a
fEoMkIOWicNK3A7C7xpwKrhaaQC7V1/BYsMqNRW86PwkxU99ahN9YQJ6j55YjS0C
PIiB39nF49blFbIZ7txduNexgATuSWq9vLxrncMHgrXjUGpT/WWi7ebccXpMRtcF
vmTXrh3Hk74iCuJGTbZqUUGa71yjckPzW3UuxTNZZNc7guk+/Bb9Ry9+CljIossh
GsusC4jRCcg9nSeY8qpDH/WvYmeoxCzF4PcxatAKkSjcury+xP+pIwFyp6YmMOcM
XV8z4N24W7zEtgJQLpKgdWJ5IoFJu+0lfHNgoDb1oDZ9feEuZq2OfQjbIlvbr1/S
ERxRNrxOQEO4u8JmCQrLjl+3N0JQW6LnmA+rY4iSc8ANF2lt68QpNNo2ciXNYyZd
3FXrjfGIYMsBPK7mV/Mpqo7F4deNQZhWeYbQFFtpZs1wCj1lyR3x8Zq9gZc9KtDT
GtMF/0awlQ7kMVrxqAXF9HK4W2ZLtK82a/GWhMYz6oSXU68qhKqdFRX4GxITIW3D
CNwH89EmLrw0aTXcKP9ul6xd2D7DoDvyapar6yKSwSU6af7A19rf67YDjb6B3oVF
ZPV9dUkkpV7pRO/bgWQ+Craswzn/lRlliXlVnTdHbDR/QKK4329dBzXRDgvXexWm
Jy2uCYlRI0Qk2wcluOeJrq9PBn0v5gsTSVQ6wp8PrHkrEdu0t602LR1GYOFaHfqC
MpZseFsGjWTwTPLwJjArc7PgsO8jSoaMf8ZKycxgfZNIiJ5fJcxtGNy7lyaWlGVB
kUpgJsP+O6E/gVByb2jksGnhksPvjVsnww08mjy61Pk/c+g68BtEfye247Jg2Kor
r6/09juzZh7WRzvQ37mnw/0M3I2ACERQ+Any4zFe5WfGjBh6MSAWfxH+zKKR1Yn0
C6pgFCvCgwZsAF8ihdV4qGfT5p4kZML3mmBc3w7rGjIeS/pOU53D3hlKqP9QPZv0
u/De9PSupin9EbIcBUS20D3qcQ2SabykyiVpyExzLCDbDCMDVmwEQQRN5bgUDCq7
eYk8Bl317BaaiZ0hjCzd8x+BOjaWnezK3VMq2ZPBTenw0OBAHKO8BtW9ZUevii5I
f8mUt9YOerlGbxq06qsl+7T5jp5sumkpg6J7NnjZG/RLp4SzDLuK9XFGJm6M7LM0
aVrUH+8ORxwdXtZpD2QpkRTuckAg0sZtP+4ImjHKb2aw2UMpwAEa2KTWgph8FM+X
jCtEOWt6u3s26DomPEXSY1uE/5/7RqPLOPo8vnnMH4pFhHNMwXVO4kddzww9ZR7w
01NuarIZAGsVFW+AFolBB95TeaLBm+wZ1oazG6jkB345PMLLQv0eQnvF1a9PcJuZ
fyZjSscXlnBTf/5oow6HWiKnbmbCEKJcBkTjib8l+DwHjgSy/QW37XDenQSY91Qb
hQB6/GelvayKa5MxiqxxCI7KBafV1P0QZvLsAYU/ZQEss+jeAd2W3MYHRF8mDXMq
DhgOIEP8AEvmgX92/GTB26i4d0Fj8eIwQSkFnVtX1heWsAhOdMuPKzwhPsK9niOe
xJSg3HYRQ+QFQkU00PNt/yl6W7m3MtTehxXwqku9TJPr8C43Elt0px578iqDHsFR
ns+o7f4KnLkkJk0UwzFn1wUDDm6LFINR7Bz56SSU5qwApqEYem0ddivGr9vjsJT4
6/KOe5CCDMVyExNL2XNlr84j5GFwgsujSW1kluYptORXkKwdBDFAYRGLFAsIeJ5f
jRverRPLPTAU8SGnhB3fx49Cv1sfzskepSPbxAcxprEZnYs8xksu6TRAkNfvzxgM
wAD6J/dT9V1MkCKXMpfYp5qaWwV9Y4Jcjpxt32QYwNF7dboLGsyl0TYQBqc6nTht
cTSbZwbloAxMG54xdFSZPDSNGxaDE5REbw8bBmCnEXaUcgBWykNLOwHV4pFlwTvR
MGbEPqEAYXfJW5Kp5Q6ZFGzOvBKHTg6xLu4I5oipYudVc/gEc64/TzaRNh978hsX
nw+gdWTmBIaG91f53d5ZTTfg3OQ20E6hxLEaSGt6jlMfnNPR06jh6fNgrXKyfMvG
P/oVhfe5sP1aN88o5PY5KaafrSDPBbsbJQNIIc4tfOIV8yzx6RIAIQx+H4i4JenF
KRGyTFI6hd/ljYj1vVjxiq9n2Y6+T9FA3OpBfcr6/eyPtG3r0AR5GL1Su4OGDXpD
pwooDgIjZR8W341S4Y6o1/0kHmEF3EZ7aLB/Mu/sdGY5ckBJZVWTbs5xV28ddgCx
0nWhf91Z2JeotCDi3WYFD+8tsqCGWIApHrMW4skvXm7GCJUZFYRglYT3F3elvrrK
V3FjRDi4I6lI4BE1gw+NimZjaFvHFloh7jvGrTlKPpJusec04Ah1Sjt5k68errYc
ZAOMOijSzy063rWcSM2G+Z06tHx+TqXsUDxt+JjivhTnVNLuDybzEiKEpvmFKtWp
o/+f1YN0zWeGNTYT/m3rhfARMfdOgeZrWXIy1BSktadiHKP5yFn/4uPLWl6i7Fdf
DNF/jkG3DNuFK4Rv0U5h9mpMoKhl72gce8zRJLCyGztQ2ucpS/k5oykWRbrkoCZY
3tv852YBRCEae+OFDTve866GY/VoluMzYrBec+8h3d99eC86TNM8hcxrjphe8pZh
zqUUXKa1jMysZpRn37oCehn4gVYjzacj4CUxj2Osb3XiiYWrAdG3HzK+2yRHNQR7
vjamZnrMH/94RQ1jEIHOVJIUGJmIXgCNzNUSJbKLfvD8YTeDhsl4/NnS71svjpAY
/kJfNKa2zTLa9SH4q4Wdf7epmiRB/WvED9Bru2DnvWNnvqLwTeoOVzamfaTwwFxp
0eA00vwqjdQ5t15SC/rws42tCC3kJCXMMzU7q8FBxApfKW8iz/D825cUFghh3g8k
HM1UtNcj7vdMnVypDywx1cQE/KehSFL9sg+2YmIEH3JGNtHn7V/k6G10P7yldDbU
feJCrG0amBDxy8vmEHUfY+I0m9j4RFsA/Fn55eqJy749lAAntezkVERfJq5hFMGg
BeRQVGZSv2X9FplkgMrx6CfT3c9atyY7Njeu340T5nDPtlOa5rx52x8S+7efhaNQ
xWiGA+bYV6DvWGL4BFZOLDHkivzR/6cv6MCYtvGud7lklJ9SviB1cDtTLZCP6Rvf
ApIJqPmyULz2or4DTPcOUYNAExpVLGdOfdPLazXRTGYk6UoArHtnio5LdG+0l48M
wz4SUjaeerNY6pTUW1NsO/AAMZ4YfWvfkDjotdxbQMkjUFR7enANcIW3Six72yKA
sRXvLmib/jWxv1rLgsXX5H3+Rh/YOy3gYY2kDlJpBbhw5udWXfE0y9pLRKf+d+3X
XTHPr5wKznx8Zgtv+FjOjBwaAtl3v1jy9fdAwhdcHiQsiPq6UOVINTcuvSOxCJ0l
Y8C4wpQD4WdlEUiGnA+OPpmmEKjsu08HVuWs94n/UrduVOIdGxhkGmyZIOZCpu9f
tKub5SyNrH2s4tTbt+ZuXx1v+FEz6pMqRWzhfhgzLlrhlQ+4zY0rW1m3EQ9rpum/
fTpkvfXF/txsXSzl6G9sceB+upjdp9YAsjUpavEWx0Rs8yfRLyV8xBXl7Ykt88OA
y8yc7oYckO7z8Pofqx/jMiosZ1bGJincScpzGRvf5+eS6ce4CdTCQBGnLxheEFQk
f7i8bIE3MA1bEtYvMSLisocuyJ1DyBwjnNd+fkPE+Req9xhET5CVcBtKKdBcQsnU
5X/UKcsGL0Cjjod8FDKa+TyDX17A8PmcxsSAnSgA6xO1Ierok3OfhrTgKA0TEMzH
GLfCQnGKIavMxASX9xf3KogbAqI58+3tST8V9IiT/xUs5VD50/u3+ULM+cZdIw5O
nqo/x9y9HFlT0rj/YrL7Ff4vCe0lDinjSIeNkVxbJ1rGSDO33dP+9b1O7QqFzCcE
Cf1834y5WNb6aWp6hzXtDYuHVzHunt1R8ysxfOUmC+MRBjVDww4e8PJuU+kL+uEB
Kakdl/iUgYYtsI9LD1ZRpzag3235GjOWZCe7T8FjKB+lEWrv22HBMuH5xiUfa7PN
FrEIxuiI2cmE6EojyoozGfrrfPH3Tv0q4XquDrOay/6ZhmIcKeMgBzaOiBwrF3FH
3LvZcScdwxcZr5O8ZWyL/ghYLbxGHdAhHyJmcuD0Me+riC1KxYHTAVJxQP3i8zdI
CLlHOd8VAgMMzL+871cJTPDBJ5i9rXGZ8/k9OJAYwhtyp42v8Npmi9D+fQFGGpUH
9q0nlaUJTUnOVJRhwwfo47ngYoadTkgAO+0TItoa381mvgkjzhw9/D7tPZRF3SXB
ux/D9kqaUtI1oBlTI9ooysd2vlpTCSgMPCX/916trkx2oC71XiFYc37m/L4drhzC
nyp2oKWPDyKvmB2ErJi4XXUN3djX1KAnfssO4dHavt+/C0q0GKaxAhdLqNudis1+
1KvDsCQmd2HWP4h5PTm3Qz7wBsVR3TpK8AvX9Hkyz7If8ngsDiyFKSE9MHSiYBbH
JQX+efYJVGSAD0kaLztgOlmwxexWnTOleUwmJZud7GfWPmtGxSn3ZnN0+IYzilSY
93xZH6RaqDkgmEQBTGvSrnxCCkDWPMwnZUqypIs6c6w3TxBDJbE/tGYnOOhuLv+K
mSp7wiWkIaoYZ7RscFhkDr3QkmkRHOzbWbQz+ckyyCTc1tMy68NBg0uiyq5hj0Ch
m1Qh4bnUgWsSNc0UVes4r4RZN1X8gujV0+dAOs/2WI3XXJ1u6nGqZc5CWHhu8HkL
xrd3rRLIh0Wa+3H8aLr/SxJO1TMDbVpsakleV6I2FFvfsnPDdw2L9LM0RKj30ieZ
XGZW2ygI+rxJxTZdvz0mavb56J0CJDAaLDcsA6IcKGutPx9pgfUW0loUwWTf83oP
MWdyfQRmywEuDwJ4N4Mn3S32TwVvML702/5PTGwW1wnVT4azrtoFCQdRhM5iDrdQ
jftQ1Wn2dA+svhMEc80sAWwnti56/yo74rG/DZowFUrUhKUWw5fjSBPAdnJV2TFB
s8Jzyz5uZ5AVJ+JlKpf/XfpCrEZiULHVwmUE7OwbgILL7miX1Ycw3QlxejVpYs6C
bMs0Y7LSCRwGzPr3OW4TpWQrXvs2+35XgPSId9xElUvDYB7IO5f1HF86zSFZWI8K
HLSFHtHTdw/7uHjD/tf77iJy/UReN+k1nDqVm6CmXcWBhhbf4jGi0441DQCLvAn1
wtp/d7rom10lmGl74gYQ8dceTd3aq61mZWWRcmFBHyAIJUql00dh/wYkvtuGuUJ3
Jh9Kky86J2zBiQfOzuo3euXYO2ER+lNVC1JsLwnzCB9g55lhd2PiR9+gqzT2M1Kx
z7QIt0EB7O7QEXrSuB3dFbziz9aee6QNtAVaT2jRa50YmsBkHt+ZSi6jEC9T4nTR
D0QuGHsgl0TA9H1EZc8SyP5nYd/kuJ2wezg/ylcyfJC4dYWFYyakpyNL5E3xzZdO
Sxhdyp2ko4g9CfVZhaDu2AvwEpMMr5Oc7N6tylPJIj3RDHvTKYvXao9SfalYT2+d
A8/sE8YASviX4JDyNqJkwAhUZHXvLiU5p4n6gIwAbIr4m97QbvsQrzwYSRo2AjvE
dtuuBG3KxRKW2H3mKrZ192/0p+PzjY5bxNcegzNHdzjw+iIhPjPTi8aPFPWOMWnK
9W2R0QfNNLUwQp3EU6he9AytYdnxuA9AI3FYneTQalxC22h+dePVngEqkO+/PxcM
XsdSM+EphQEmAnOwlezeLRX5istOcVZoVIctvTTHJBd+Z6HU6sB3PvV7yA1xz2SE
GMtSm6gjbbItTdnGel6zXNF7kruU5kLgNMesirnsPJkLfArvP7XG6gO0579kVwzr
EgsvR8jySYTcWWLE4dO8cFu2BmTcfWwBVBIMxrtRwG7cIBMM9v9EWE2s/fxFWmzd
I9QWV+HvrOP+KufvtN60zWphnj1ynIK/szOn26fLxvWmHtvaTsjpXgas5x89lNHt
nBr3aOrbUUFbDN5jbyteBJghJCp/63NAoUMj1Hw9GGXfQoKWT8glzGAnOto5Cmw9
B2mcmqDHhjbhWRS804mJYC1vh1UxSDb5nQq2Vbb7DHw+O4R+5F0jzg+hyrVnAVBT
wedFI7WikvXxxGXNj4p6nhAv+qNn/2+cSUg1jyVpQIXM1cp3NaLrNjWNrnyGNjDa
xWSJjZUd3W1qtqXq4aGGQXzWynFdJV7HzQURaQlduXki65VE6zwBmDf3z0s6igjS
hIWKPTEA6cfCHqftd/2eDK/PNM+e99YJ6Msi3uVqz/4azV5ZA2qJWOhKO/9SVSao
vNH5dON9A6vgGKqMtVgepFtCs5XLT2Qp69lHLyttdxxv3OVao5ivl/+VD12QpmYm
NgAZlTG53Ogxz1TmXhJbhKgDlXAEkIzAbIxsfalm83K+JQU3FHYVeQKZX2idmj3d
NgngDChmfkIJh+/zlORHvpZCw2vuWMHID1ro1mYP8ob/BRpgggo3LjVf7/w82pVL
lwr2tBl+JTslRPUIrRdC4iKR6KPUYW/ikFJWACTRGGC/32RxiDObbEtWYa57j0Am
t5IlwmpguI813qZbeHmhSUSjVSfoN/e5LAP3vNNtTu+hloCtBek4o1ZOUxM0Og4A
NtF3BOH6VvZkCPPyjGVQG+c1LWK/GrMTl9qK6H8I01D5JBMb4Zx2pB5kDw59/l22
S4x55T1WMe/WyYKIQhf2DnWP80q0LLHQo2jLiiWvp0m01Iat4bLTT6rwcw/tKRGv
2XBuNvp3kTU5u9R2U9Su2NcrxDEp6Dr1/ySGhNImrmEQNKzrzcIIumXnvvYO8Cra
eLS6nVKbgVHTuSJxMxR3AtClL2+1qAPvs5Co3o2NqBEH5aOsqJ+4N/j4oZ7rjJY6
teZ6yPTYj8ObjLRcvqhaaooeIP1nCPmxisJLCIKRorG29SRmBqAwoc2Cr6Wva6wd
eNHQn3B9Mm1ngTkJMe9U5cD3zrGPIRBsUb+Y23WKOdqJMmo3rvt3fi97CuppzwDj
tQktSqeHBMUrpdKtHAEt2eDAvV5dVlzNrEuD78PcN1Or+jivMIPGe/1YPHUJtje6
5J58FmIYKwU8YepWGuwI9PVVRuk0CUun6eLhBgFfcYQbBbf6q7ZqaT8oQxEgaQNU
Qtq3UQ/hlYyfd+FzK3NOxpTreZMy/+NRUNHu+CARxaRbNIkBsuPnHql/6RICfu3p
nsX8IpUFG1w0rd/+lGiDfkn96LJRx/N3rz4KcGKQDJokkHuAfOWgfRKPcBNr+JSR
QJOqJiAKGW+dPVG2FzuLAiGpY5tds8rXMhmHn8mX2688Yxm2VV8P6uX0KJ+b3odT
F03tOhXsxy8TlKUNoooj/3xhc9pC84WbxIyifJ6VPfcZjYQfkUBKtEdPEQmPeVyW
meXYO6yKljlBl0TZrLzMuQdtY+abYs/B2so5xPCsv60TTtbR8j/iEhMwevwhi6ml
hSXNHtTmjSxE+zBAGxAioaT0L5NlT2+ox5o9wm6X7oMRSwgOeB9NzwvkgznpaWsZ
Fd6+5ocTlIgMSrf1sdmlA8rvd3PM/zPaUVdsPudvjct8FZIa4pmlPZE8w/pRSn1f
4nUk1ALpyI19ciEoUYBEkeSf6GnkqQZ7S1/f28jStgPX7YlCeOZSAz3RbtfP/UfE
yXJsF5iOx4Bfs7pDQA03gHSVIE8JijwbwMre+VPMhTiWGFH4fApe6tt1PCEkj63O
GkxP8WsG3v9VXgnux+/H/Y14DMAsdsUDrlr8ksc5VNN9EUr67Y3FONxj9Ntpzsf/
OdZVy8WI9ZklVV2a8j0ClflaJNpi8sv62SnOA4C189C+lWDYUnYn2/rQiz0SB4QR
MDyWswntu83OWFSpUJFVDj3wVQY0T1mXi7ySRZv8LeybMKtRsoFpJ8wRfLqP7cp7
+v2M2fNJXY+ZaQUMgeHQNsizgjjN/Qz4EtuP2n4GN+dGiUfrn0szHxeMW2wnvUe2
B9R7oL1qdIwlzt0vu570tet46dm8Mlp5a+VNdm0YuQyldyH72H3HW63Kp/juDprs
CScagddhf6bwVUUzysAABJoNPL5AD8yyKOQJsMVnzsg+3/UJDrhiKzL3qJPp0xI/
s5Pvo4MbLlOQAVxC9zWAd7dzRB4dc21MW6IR0prR+ZbK4H7pkO2Xs32SQ3H3YgWk
9AkbW2cMaUA9c0XEJtpF9saTcU0RAnb8c3Rvhz/iPZ08K2/gIaHVJoyixpUHu/Ba
GG7KxPL/3yuhbzEATLR/Ul8WltOpaJev9FikEQ2h8DaWp/l71PyjYAyicKsMa3+k
u37QGz0GShQXbfGbYtau577HvVsRnXsk3OqnE2cVQ6H0prvhSgDNT5KBcpaIhHqp
CmMl4lnAlni3nUIfUUDPs1x+EmUVMG10kNUq4iI7sMu1SbFow3NnKEO4qlthlUda
1PJrLonBoTyHKfM0mrgQXfdf64YMogGnifuNc0hkLVdQiKHfOUkQcYcmrZrR0D4m
ltgZ7EYm8GS13GkQwHxWZIFSHax7AyHoDFNPLOQ5buNqvwDXtXzyRcvE8OCiPJgJ
jTl7bJ9aZmJeM3uP/pM6wfuI/KGDfBPOesKaNCRUOL+Ie/mtCej8CLMan9rOuTqG
PgFIgzLMG+BXLUv/Yru278h6/Uu4CU0cXQh7ROw7ddy7XecCwhLGiSDNVeHqVyu9
n8FyRUjOZPkKcgdLIZJNG7vKBrfnK+hLTTRiNXSvz4JYuohy++rScxEh+rDx6hfs
Yy9aAPic28CE+23OGc8lG1hTr67maCQRUEUSMdNuoBmPWhpb9Z3Kf3Jq+P8bnbm9
DQDSyjsMbVQJ6u8XV0IkA1c71ytPv456U9g1+NXrxBrPP1V3gN7n0MGwTel5BOHd
uSq1ftCv2IHmJAYDV/7SYWg09FqtbBZByzln1zWckzJvpNyEeBDSgn/gViKtNMf1
DnUlUi09wsk5YahfWPvrlLpwEMSZHaucTgHoDn4/VIhpdw82PrkCuGn0wViJRcFN
JoPu+A+MiC8ouLLsch9Nd5UcFJGpTXYrxiFROLaQkw1jqYMruCX+loeszAbW2cg+
E6pT/Najm1kfSirHGwcgeYuy6dDcTOwI5fyMnndr/btAjppLNIoIWwHOH1YL+tfW
zMm8fG/0fo93gt1DFmFV8MBVQmIxPLhwUEKHhOQprCl8js/8oV/5uuk5c5LBG4up
WB7ofiSkPcDxXwDueLb9ANQGuVKvWbd1bOvHUNu4ulNcagvBL7QYgXbggGy0WCCc
Zw40MqFKJ/z2TPVx/JkCliCRtyKtCusDMgooKHO3gdO2F6g/8uW7dQg32s4Yt2Kk
eGUQOdOTefnLutWd2Yqh1RP6aX2D41wMIGwYHF2Z0SPBuqxpoL1qRCY+jU/ju9HK
UTHYUMT/6JbgRnunQxlVkaAz/+GVOXSNVN5sUIDk9el/YYFDsGphF7m2qL9JJe0n
RujPE7o8ySUi+WUCpEBs9py9D6U+CyVx/4kn9cYMIm/BhDuAhDsUhAFeWnd08x7w
nTTmZZPUuCNM8eaP9zzrIWdKil2JqzHV7iEIuFsK5ZUP5ZWpiP1rwHSs7sM3VCCt
Qy92xXnRUE9jsvAWy6gA3o1+srF4kOT2XMUaRnySr38b8LrpHdtHaB9ppWLt7We0
gs29D5L7JiEvwQbLGdDRsHV6Tc71J11d0Tnt/4CGW9SmzYvUuDUiHR6pitl2wSnK
LbfgPqhCIbAIdxeyciGzI61KmzPEvesNGCO5+nP2kHMAOSIRBe4pziZqIZjZ7b3Z
epjY3XSSo8cg+DITpGbaDSgVqE5AYb85LvjxRqCsIX+R5yyakw+So2jIeOJZ17mZ
ecbX6vEA9U6WFdPZNuv4BbI4uCZOLjRthX/tWeidg67kUylBjimWfXIGq/gW3iIb
lapyDXMG8n2F4anrleC+mooAefgfUseACA40UqB56CN4equfXpgq2lwgiJ/4SsRT
Y9PtEVIGK67IogJk6WTabnCVyYbgFbZ8NRNqqohAj6Mj0Elzj3GbkXlT6FbZxjiQ
TdZUC6+V6264+MyhqyzIq9CFUH0DfAkpyW/ttT1F66DAS8rsnEJRiPMhquVRgTjC
WucKrxGT2YcbbTexZdohyk4shyvZYTbNTAT3q+u63PiGVR21Am7fXjNFQLax21+f
KHZXyq/rGA7AMD6nzLbC46hqtApLm/dUnfUiv9D9MFxUXWIUzjizDmmNvJf1asjf
VRAHz6vwKhr+3xsorbx8w2Ui6GtypmcUHxBRpf4o7bxRjsPAVntlBJMkWjZuWRih
fBCa3AEn5+tppKpG9uMH4AlqAh8JxsPR8MwrvjPsr5Z3TPfdZtAmxNkKsVpjKcuI
+QpWStz/pHTjgm+VFf/VuTN/FWhrY5uwSdRWyA++F8WUXPOSKSygvVbRxYaaKRND
NcGUkCN69kRsBhN6LSTYToz4jXhgotmP2qxi13OZF7DFj770LSsnFI+Q5GhXFH5w
kr1f4d1NKYCY+KUSNIlJN2S94HkUnsKCzlYH310b8+4VM7oUeqDDX5gewQVy9FUU
4rFCIr1z2dEtJ8JcfVD4yxRrfdfZhma/EYFT1b3qG3ucr/HnP+OmZSGPHuNO5+X9
DfGUUocA4C+kCIk0HXSno9PcHjoJGG0IrqcUU5c+sp53PNNle5IYpn/S+Cg1BLhS
ldofPitQj1j7d6U0EgjHzZGKpCtVzJzVsQ9kcPSrw2vQSdjrF2f+1+2SjOohLtdU
Tk+niA7Rs2INOeXaEBA0rGB3gaB9KaUXpEoAMR7FMeHKAhoXe50JwCvrgYLQK3CN
HHokuOs2AUJBfMFFaizcWBPjI9sLW2SDlzlfsegj3pzdphu+/Txp4wYEz4SGFo1c
dbXYoc9JOmfjGuMYm94FoKyuk8qGTgygTGGINOT0q3LchZwl0hzzUEi9qd6N9SzO
OUyQdO0JBNUCT6s7DbfZa5KlVCDfzURThDwV08egcwBOxzlxdB9I/iblQFWZzduw
rzUxRdXbki++zuAx/qGgO9cMFzDacIT2yEqKMkRGFYnD0zAuMpYunBrrljJSjqnI
eFQLv2457DZqJaLAMyjAesNJCwtheRBzMWiCeUd0sJFkOZ3mvvhcZQqs9bXbEQde
aVpuXsIiPX327SpAqckdmQM42ZrJ1zYKVTlFUQhPjUASlKa4pkbkC+/2ntSKjtYc
uxl11F5HcBSrOAHcXhIu3mx3h84AwBYu0gqulXchCysXJJqSQ2zh3pzAaMagjxZu
55vvkGxRcavT0/5XU3lx1hJBfu9/AoiJs0IeRtBvA/cNusx3onL/CxOXbYjT6jp8
AEWROYKsXEYz8so8e8KQjS0hAqvcUGF2aDKXVEHkV+F21NEWZ3yMhf8meMK9z2DE
lS2GgAtMXu8NqFqiLIN86HPyj85vqZHDnpD80rpcrO7JpQkbpnOhCwTlwUa3xyhj
fzghgrdOw3pRvgxJd1VQntbXg/BZUn144ePkQoCQerm0GRhG0PuJNnYwx59twQ+L
6YqiXVbEPyuK4CCaYeFqikkuqLH6Y7vd+vmAK32+wMv16CS3FNptakrNgP3r5MrG
cC9j4t11vGOh2SzGhImFYRFo8mxR2YTNoR4W33s+t/46HUBVur0mZsQez7csjxYD
AiigjtqNTQ3DoUuZ6oNUvI4ebFXBL/InvVE6jIwYwyxzpE+dhZihQSXyNMxOHaDN
MxyhFTwn0b4J/0tAnrofZYFkHnormvJa6NPTUVPPVmvLIyWhYlkF6jYVn2oLwBbS
vINdIg9cJAunNfuyw9xoG9bEfuSDpdppWZfeaM/M1tWGpqQ09pbDehViX2aFGDcQ
JfsDW0w3HljZ3I0EKSav4Ieaz3+IB+er9wSDQ+SgeF9nWZqOWRYKoPzd3cDVtR+B
VMbtK+7sdx+uVIyD2L59dzLp58+sxe9QK671QM2uqWlOxJcYRx9s42V5zCP5GVX2
G+yAV2eIXzWT8/tC3KaPgUiQHEF02N5RQ853R2wRVyyjstWPNxvyXt+aZZBOL59C
YLndLrUqEA7WUmCUcIF1O42zW0QWKrd7mMyf81l5q5wFiaIL67hV2ume2r//VIXs
+9yge7Si2MOhIWU+OhF0843DUkJx/pl07EwmkFkVTvq5P54ADZiD61TEAWnJKzDi
9LH47iMaMG2kcKPHUNtu4tHBzWc75yIn0XkO0s/eFn+e4jQkyM7Kigudv8ymYkVZ
Ob9tdrve8DE2ICFQlrbJXyJje2JliGhteeWB2O/YJk7HTDaHKPAdAyrLYbcm/+lx
hFUaiQhXjl9e0mydU9t4NndZ4G4NG6SZahTHSiNtzeoBDv6ealZr3l81bt66Kk9b
Tf+OU3I9/8/1z9r9YIWhGv64g82LVkvBAlcPTjrnTXlaqPnS4fGVvsh925FmiKZz
AnqTubJKL3TIJjMBfPHamxY/vvgV8J2M2npr+eoDUohEIzMxLsf8c5jQjo6ualpD
7J0018jkUuete3u9OmWXsVJi2/iOYX3t2HWSJPztyPJ5dylXaC37bVKmxZgOxYfL
RurPX1zwXwhkSL74k2uAG61xsXLmrh0tzGduNs88swW7eI3+jAjI0VVJsWzeCNn0
hmoHOVptr+EnQJzcWqAIIGoZA9s6qesmJLRtq+tDXylosvHHXv29tihtU0Dyamvp
O4WM5Q2cFdjXFcF1ZSKKk1Ud0Xyqd1jAya7N5ypLnHdewPy1Cc1BdLRpeRfXWbZF
kFm20u1QKlszQElW1+WR2WmLs/56P5sPZM1eGSshTr9hkgJdAQQg0IDWtt5uVe9h
Rnsb29MXem14QDtk4mQaWCyE3G8I3ovA3D4+BMzSgcD4WyhPblzTLk+sDTXTOBTB
ymzPdud4xAiYycMpxrKdwdoDBj/krA8PETI4zMdgik7uLA3PmvkJhLWckmNEPpaA
4XdyMhx1y/7crcyJvcsObqarn4C74Dw10PJnIk8R57/zhcvQKyfT+JvUYBigae2C
wT3FgnPYzqEAP8DAys0q2Wfv7I30Bvw5+HpnIrGo9iymzSnNCbk4U1REtI2bJ0iX
w2igzpD5L1csorsHvsgSiU0uf7t5wxUbd7XW5dxrR4CcAGXVkcLzmRdlalkFpZlM
RrB6aINEEbCjcoLy9+uf8ICoyQ6Ph+eENyQtbEGPWRAhjo7d8mVPwjnlRoKmjuFP
B9P1bQD70lSIFqRmQUIwWzfP9r4uOdMjGbwK4StQjBnOwYwzYmjknsiIaDZXLmq5
tRmkOKvydmOEtyMduSINGPbrYQjwkAr3x90zT/O5usvfSgPtYh015CJdbsNw5LrU
8UMoDW4N3xtKH3G8Cbchm9ZuU11B/KqXDktpSPMS0CcAAwFQSRm7e4YC9Y9FXUS9
twDoJ6uCeI9LqWptFs5/8KXYfRmUbnhdLIPlQmLDB2VOY8jXgNF1vXAcDRghi7Hb
gcVj9n4VTkMYjus9JpzeIKt6EIPag7v6F57R1pM4Yhec+Tp7EDBgMm2y2pJ8eHHL
oLJUYA+B/ZswFYZhmEsF14ZKNnk0/vXZrjN4frsRJilVBbmE2e6AAW4OoQLgHJkw
eyXfpyAqTk6bi2hZ1WIRFuoDrNS4P0M1eELeBw45sbtWxoBr6SP+ZZEStxsR/IV6
kP4BhHZFYxkRvinm1RWPQgbyTa/NZ5hft4YizK7WkBGI0VM0P22qQFfO5Ahc1h/r
EzLqHo8yAriBzoIsDbCrzHw+0YgOhxxAC6xWwM2ZRWxW28p/LkrBgH+tNjPHSa8l
bBENTxw5bQTT77rpJ5VjDgbonyNgd8o14i/YMxUqIIpkH2PoKw6hJlawLL7auU/5
0gqQXwaozYzR73zWX/zstJyP7B+AVIxh4cf4P0nH6eAxYuM45u2QYxdOE7H5vG0q
NefbHbP+1j6zH0/3FEcDhwfrn0rengYG3BmWcXqfiDdd/Lp/TOPTNYk9jAPoDpc2
hM9CsZa0s3oiI9g71wkq7b1x/6XC2wN7XSGIE0JCKgFEwFwKbCb3+BXSS8fr4zUx
MeL8DZK9EaUH3Bl76DoXTfVHL+GTryv3+3thxo8XGb/yGWFCo2C+pON8Zd+WaqzB
vQnPpFe4GYXzu1UpV1z18InQa3S7sLjhqHqkIj2qe90RakWOB0fT4/i3PfXs0WSI
jaj5aHzW0i3PyFcweJWhyqWwqlbIdojpNhlINhnkBoK1mUZKRCEO5jT7J343sTAI
LZ2488vMVdSCPVNQY1r6+EdyLDE6Lk48yZBDbBEe6RneE9mE+d7QGV3UlbSWLrIO
kK0KAZONwdmjRM2rrABa8s6upa2GSmiv1k3XNRIamnuutT+Anua62084ewidP6h7
Uwzc8/EoPDvJ1wP3H4b5hlJbITf8Eui/Aq4FoqQqPO+1b5TabZ/yvMYehN30Tc4e
EdUvdjzx9rNP+bopG3SDuJbS6xoVLMCaVmdG9ETKOs+HROEvDr1FE3/uJRVrRSz+
xScz/n0OEEbfex1x7xH7bU0hINhIbOD/vVoq3KS2v56UEbs6sUZL3+UTQXsBpSCH
QNhmpN62YSXrI8MllhXtXFTBFYhbn7h06JIGs+tdYYnUusMo9tfeJTCVggJMpli/
vzuTq0T17tTYTSefDUqoHLZuxiuz4leEX2oexMY5AHQYAbUpkPCCkaySULOj+/L3
CdfQZvF0ck9hw9+/Vx0jxxAfY1Sh3VBo53PKL81sXUGOqkXgHT26RtQBESmalnWD
qJp52GUm2aFVTF+fZhWfh/07VeDdmkN+A2Xbw40v3P0CtK8jGju366bKpTMv85Vk
3/rrhuXk2tmn1qtioytceBAFTEEshjJQpFL8US/EhoZUvK97bDgMke8jqwIPGK2B
Gx1bs6rdb29kk6WvuaaVOYsrQcjSY1iD4Zt2blSv7pFQyhEgzZqxZnEghoNh066O
YZmvvOprBLwM8Z1RacOfNOO1vYO916lrSJ3d9oZp4OxyYPRHkW7x7TlR5z+MvMSG
FWAgs8uQLA75NPxHExFGjcEkG/m5AMpA9XMxs3NDroDNUOHmbOSR8nf/VP2V3yef
P0gkbRXSMcqdwhOSYtjz+PhVC/eGV9DH7uSzzcW0zO9IVY1xUXcD2a9RvYumnQKa
VmKrmuP7Wcdelcsa0EH9pOamog0q/8Y5l3LtyDtnkHL/UHXxVeEekcyMpnVUy0su
2X0GMymV55yGf6AXzBQRX7EVWs7NhAHChWjpzfYzu3mr1MjPO9ELSpLOLTo1GUaI
+RMxg6iceb3CsyiDf+HNRKNJPpuLUIjtsLT+uXcRzsG/1VCoO8nMQqhRxhqk99mr
O/sv+c4fEskTT2kW5ABXou68/8yBMRqZyzzgjPpmlSoBwBY+YGIJrt7EhvD9+XuP
0zpaQfxqQDaPLBx+9PFbod9BMfwatrJqhMdYkKk7xicXryfekfZ82YhrzX9aP4/l
kLvw0Roi9qAuN9Wf92l30niIxsIRhrooAUozXrL+JC+80Rti2Toas2kdzjJjiTcc
Bab3i5930XxYP34FWRUSpYQDxN785LMa/yTpzT9DFnHcxxICgSq5hJ0L07OA0eS8
iOxedbkVoqcOiKR1vRKP0XdPkl19R4yNRWSFIyDC1UX7bzoA45yPbof4FvQHLNL2
Fu0cWtXKkW69JrjvKCvhLE2Q2o8V7Yx5NL+u25pCRfmEbl8RpWeY1jUDTFtvv1nP
igUxZr4mI4/KJ/UAMxBCIf2fri6etwmv/oD7EkzbDa3xOQjHSgz07DieMnPz8n30
Zdpfw3C/SdO+HLi4aVe/pvF9vwM9wON9H6r+3d8Pcbt7qy4Ntn9WOBgmlFKfAZyO
BTlLaiw9qVzSwAg2N8mMk5fo01f5nNaj7XJsSHU7Z1fUZVY4HYaORi0OHVPTWEGX
nt4UZvorgbpn+ROcE5+sHHxk/ubyJNQRWXsF6uuWFRtgKCDcn6V4UiQ2pY/yG5ri
DKaGS5ibZ8LFCwoetEtMBnDZRxIaWVqfhzZu0J5O+fZk15AHVLMCXTKY1AqJ5/Jv
bAvUszELSSNdqZv6juA/o1KxhRdrqdpiqLR3y9XzDYz47r8pxuBhE6MK6X2lbR5B
zv1QiPnRcgAItVRBepijAxVTb/D4Vjfdlhr5EhAyYO+E4NFQoYjhHhJWV8Ogse1+
EToikA7OVUn3m3mT0ZCCqnhFCIr1odLGTm7UpdPBU8/an+GQBZvyP70NbNwou3iL
osrk5+lL+bk+2XQKwSwi1psqE0pO5EZCy1q0Gj/raSjxsM45aGinODTBYZKaD5c7
+cWxkQx+1K2LkF1bDynhEhGKXVbeduvem8FVN+/wy5gSkMHE1XW42gK6RCRjGKXI
9YCzEW4dzD7w/73q3skllQq+vYdu7xo6l5SRIwSWGz1Xog6Od9+uFB2bHcFRXe1S
OlqDJkZst6lKxki/nkX6iKJv9ZeqecevUDLkmfQz6pbP1xsrOOjMizdzn81pemB3
PP2GfwwfG1MxaDW79OccAGiooT/odkELfTz+feFTdSJTXoZdPm1F+WCh6WwHuLQn
5Do3C1LkinnQ69lrNFUgIqdP+YaLNSX0dljCLyylYgS8vzyfgR+U1UZ8XnHj9UPX
j2OMsFoJKiimOxE6UIyzfNv4LXkfZsHV7muflqP0I9oPsuVlrH+TvYL3S540ooH8
DOVhhfIOqYAyuLWXvhjaXXnoixCevNgGnf63MHMmaVwpGIJEZ7wi+svwv20R3j8Y
SUeU0t10HFnC9+u+CkYnv6iL/OPH7N9uoZyfoy2QydoFByd58zljPbrNIvEJeL5o
OFT5+p6nLsixGs1Mqa0IKpDZOGi9JdR0flxNjqofEk/NaoUNyu4QjLrPmmy6O3fV
I1IqgdktcgR4BxAqK+TtsBxghMWTWfqgF0NBPrY2s3nVSZkK+t0SjqTXm+3XQSkQ
hIYTyN6QdmQ0SxVcPAO0bxUOHXmyq6gwm8fzdkaTQwgSLn8PTI+S8qCHw8+qSKmb
LTeX6CUIin695F4RdFmlWO1FqlRZ/kgxYcbWUqIP0pIBD+8I8FP1PVXNz90O8hsG
DsuypYJ/+FJJ4jNb1Y3ERy1ChLXsqsqOOHYH47LHv5B/5z0Fq0Adf2sbUB2ptV3T
69lSeQpSe6JmKekPp92L5Pt5BFzzBN1SpfOUQUC+pGMDGF+umxRoovWGPCw9S/fT
LvLhBWOtumfgkvfeKP98Onf5PcMkUD+BOaJGOu/jJfncUfo8OY7jUHL8TnQLIpkJ
ybLVSggWzQzX2Gg1h4hB+AZh+QzGq4seS2ekymdFbU+yR1dZgsv/aIxruyVAADo7
YPM+BVyeeb9ZoWtYzHui63gJhv46FE7NOkdrsCmQ0R6fWXbEpOXRT92zigpXQ6Hd
ImpSM2GXS5Bu94w9uZPjMXU56NaY4MVCOeU2C1bE/r97YDOFIpmimBq0m0oxfFij
JxpKWRuQV9oxj1bQ+YF2ClXEqbfEgR59MjaudgJDcIdXm4WC0DBOzlxQWWGUwXwx
pQIjKQ3RYtf37hMpyNqYd3stGnxhrqeOnavZrSxQkVXieVkxX4VlPlcfkiDZ5r+V
R4v67uPo1wlA1d6huiHLC1RUwymocmrBldUxiMxhwLPDg34QkG9F0LLMj+chXX7N
Bp6GoOdM8SATbXO/l/gDNdKllDlkyi5lyUy9bm8ruPEZADPre+6NFduuAy97EqzE
et6d9Bh34NFxToGgGxc8gggFgrUooht4FWGgy3TI9BR+7kZeMHIPiuINFumpaIQF
0XpLkhkPEo2bPpycQZlBVURyS/0HsWrH5jzFqjC7FeZtDOb1dJWcNfgAtJ8R6gx5
AWK6Lf0ZiB18Bwsj1cB5Vb/zWKxQlka7aLMleQc6ljazbgtAL8hMU8YmKYgCRkvY
4Ftd7+/503Z+iDWQ5OF0xGh2Q/eiS/Wp5PyzFYV68A8BciSXJeZaErvWl4XHXVnv
0JpkI70UZFYnG4az5AexpOhUikaPK/fAK4Hm+yoCF0zetRUxBX4qj/HrHDsYcVhH
YKgBZgzQrYPaCkpCtHICNFogkpnwQnn0Plm+7u/FLdvQm5h62wwqyM4YOiuoklh8
UbaI/wldYErHQlEXsj1qhKmdgepvNLv/bGei9bFGUIaFicVewk9S9PnT2c6926xN
+oUzkWVTiCKWaTMD/nZhn0xUcRYtUM03ctBhskL5dKV21quqJCRMZRcFt8LpWAft
a6ylq9OZJwPpi0cZE/mGCYnTTM5jzEF6PIE9Gd/kzTbh5fijuNovF+HYY1g8X9zn
8i3oCFb2fCKlVAyotyV6tnKf/4WHklPYtJs9vYX/yl4dn1Gdf/C1fHvvJ2bnFVW+
K7/JXxEeEAHlVh/49AZJOR5JyXj/4KRkXQk+zI95V5yU/BpUI971UmeJ/SrM5VYY
iOCaI3HiZYKaPZoXAHv3BSyL7squEFXNFI4MTqQ/Cf122JQKZG9cWDnvXLZ+9ckM
7aBUrtT/wgcz8FDtvW5Nuv/f4hWKUB03wdoUe0wquaEVrJ9P8xfSb00lltepra0V
RDNM+iC7vOJnkAHJplHVScRy1wG6ps24isFV0z2M9TytRfUZmmQmCK5ZWcTvLswu
Dj/81zy83l0bmIIcM7moR33v0f4ltFiWuRqjKU2nhygPI7Hyq3qE5Lx3TV9G8KIw
++Axv3ZbzRyLOloXp2/FNwkZ02dBm3hwrYvp9Wfe7m5FB7g0Eu/uN4TL4cniD9t7
cQwB4GTqW1vj6TkEc+oO4U+jVU6FRaOf230zLZlC7tXyrGEIvjddyUvRtBA0RB7q
lRI2zuWhX1XYqTi5rJfPOtgTubhlumyv5+w9Ov5IVmxu/hs1JLLWIhqOedb2jikG
IZdbsSFd7WRXeV96fZIEG/1Gm3q727SlrBnQB+uPwJXtN1eqFt7kGU2xYhjT4Csn
7mRc19AuMbpTSf0KfAh1W8MmG9uk86QyQnzdsNxVp+2ZeiLPCR/ikAzIoUMH/tMc
sMFZofjgyA6VNxn2A15WHFTboaQv2A41eIAbNqY34osFw5LAdGBJY5FPZeS45uq2
PxPqdVB+CuHrNAWbOiJfYBl3N7q+RWY61GF7EFUNNPKsuI5gmMK5bLM5gEG3tjPj
TPaGv81NUQeysmVWyNKHVQBh0yUVIdDZ1Al+abFgF/Q3PAbtTZ79DJUKUc+m7UNz
U5x6qJUg4gwhPrz0fg7vPFr0qbUZAk3LdF/K/l74nB2nu9DM5Se1hqyANTvncc5z
nDbcu5/9xSpesVX+/iQMNLJJORi+mv1jD9Q8b9eEE2tPEHtrLlCl+423JnQimq+e
k5Ux/n/P4rgwccur0lWdRBBmJ+h5pdLhyQ6We1OIp69xurSFc6Dr0i3oQfLbBpIF
pR3J+Xlwqs9R8te6005Ip1+ec4hWdo42PQwdHXoQUfEnbiqx7+z4I8QluwTwngCK
Q/s59sEVc6qFc2uN8AB+WtbGcZY/X7mlAf3u5ySI05EArKM/yM/SAzmCUjPW9NJ4
GblqrfsICQ81RbGOjo+uhJjPkUY5yIK38d4Jf/NXnP7Zn5sU0VtJWRLeM0UHTfX5
hAy4MEF+n/ziWjlAQo6EOU6e2/ChBNK22iGRf5IJHLgWAKqcCZcGhNOjix6XgOTZ
4nlGc+oT+56298TcfjlFu0flGaVxlxvUDhbvcDtVJVmyG/uFb8RjZxU9+TznB+vi
oBH4cNQYxVJqDC02xBNMF72glxzZnKqt3xAQx6HPWsi9jDTsRE9P2YBvncUZXzRP
cDiBpjQ3GsZAaMO4XWyjUHeezj2JZSLrzs/DZimVjmGYjl5xWR7ehQnLo15iGYdG
U1yQfix5IS62rJYrRVRnvFkQKqfOPxfIN52eKWuKTAMwXeaujx5/pVL+wvHY82xv
95Iyt1bMqjXTORO/8pQpPkPKHhd6Ja9+SC+SHa7tdiD47yuXX9omfBDpd+etYvob
nHxtxKlxGdy/ooAOY5lGQqvCB5d/HyrkfO6jaJCA3DTnzIWx7/w0iCdxsueFLm+H
nvo0GzwBXfIVlax1/ibmHudkpzFOegRp5RrKygRUcz73S8luAqqsAQcu5KVFtTIQ
omHy9CTRl2ammHI0qsfoBYu0mZnlx6RuIMD2tMOkkD3aQ7h99mgwrN2dX5GqCjUu
Q7dR4d2W8fZYDvCrdb4/TlliWtUbCiaHgaFdOs1wrisUX6c1cG6BIlUPX2ap14tU
cDXHjkVtWk00NQ5WbdIAB5h5fdWNaNTLEeYpEuHcpLEGXT2OV6MYaBRCtzAY6Vob
mA92r/iEvAdKlpK/oIu1GFLwu6DjQWBWS3uQti964jYYuT/0vYIOEeF9N067Kg8k
rx9dUIwsLOEXLO5cZH7WeclAZi5HupLZlba1jrTGk3g76xqy/QQRiecrvAktCYyx
08WHZQoB8QXZEGVQUaGVEsesdw0FBe4n6/Qft1iQyii6mG44MjAQSKOwYZ0eABop
EEVvFYiGy0nZLhW958gUAv0ycc9egiu6uVBzeTjgdkxSk2xNDcn0gkOcR2Jjkze6
osUHXlIUcsX6IMtzFjFQJ9wHy+CEAC2SBWcBpdm920soJqAK/oPU3kR1K4ULpE7k
vlsmMZLtr5epLsCmHKIXWQXK1zotV54Tj7AW++bWIT7azkBi/WXQZsLLTjTYqNNM
4wKagAmhnsYXyLvfYgoUd1SKo2ZCRP127EntYXbXVEbl1btyPt+QDQGXaqUgb7II
c2Ni9V5f5RHJ7Cv/QEANxNqckWYqstsEJwQPqOScMRCMDQDlDo9zttwecfiHt/Y2
dELoBjt8YTi9bq6NpFWdJ/DI7+9yDMl9HzbS+mkPxw7OgAOER+qaraHQieBzwxTl
5c1VqDPLYEIGbXhEfpJ3vdlsg2DhfseUiolZg/J00eC2ysADkUrD/2GnUD5qj0uc
j1bj9hmSHtyuQpIVxW4qIFz1ye255UklSFPiO0ZHSUp/KsGdKKpPjGXnqwEw3lzv
sLGt8fHlbSOirLrFnVBdiCITjc76xB6xJ0dyJgFfvvfcHTp/P5j5A3VpfhK6ThFW
u3ZWdtJ2yEDSROcIJFi+TeFvebyIFm8RB5Gmu+40Ce5BITKtlAxz+MjLWbzcemKl
keM4bP6SoNUSLwso3LkR2zDPVpmAFqJ5VE7AO7UsMKLbAKe8+SCjpGxZb9DJjZy6
ucXBjSjTfigfUm9ri61tg0PCHOU+5KV7gR/a45QQC8rNTR/MsHIlYvfB08zucaUt
Yk1K81h15gywXxwWMWlMZqWFYDW9Vmy1uY06Bs0aJEXiTUfb1TB2QpxczlB0JpoD
EcC1be5mLTRq0BsJ6eJK3Xvshu8XDWMqkofFzP+wOn1qa7Sl3tS/1zz8hprbRCUt
nY+0deaEn0BVvkaPAaq50wqdNAdXJba/Jd7WiOg7D57GJDcSnViLa21jOvFL6tw8
Wl3KKnuHIvNBdsL+3VOz2O0FUQa11hkF9ymM91MeNqkFv31OWs0qFyjOLtFVdRji
TTzuZw4eV4VnY60I+ZMyU0QRMVKPsNd6/GHUJmbqEgLJ/+orcd1ppS6DZ86pTk6G
fUkyfxr7sJjvrpriRMWUCF69XdHtUuwmpcii0qZSTiiYGZJtrVpS58Fj5KLLoX7u
DtiE70ft8JUpgx+ANSblzRWtF+oatZDrw86JH/3OBq8csbU92/z7O+YpZ94vPW/C
oTZVxr46jOIHZvZ7qc5aKIRXkrvuvl2ZqohZ7xMTHbwPA/i99UrsSFqnrV073nmc
LhHHzuxCC9Q1LNsBiWtmJ0TDaA/ovn+NVwVi6a6ly10DjHI8PT8y09gsXukRcLHE
qyBBNVGBUuQmzoWAnv2LTleTE/c14xrGeysdrA/xLtuEcsEiagLHtuX219iEUze5
WgVIV+i86Tc8MZXqZ8UzOc2dAIiL/inQPgvVVfIvBfdhivyyFfCb4bPDuEcggfJZ
EjijWUp+kfCKFAIjL8zX/dy36zoya5BENSll0QEw7RnJJ/YwzVSx23P461lINOUz
C3UFqUWYBcki5Bj4FX89ZAqY08RvlhiAv+w9P2fEW8/ucfrGjM6GBtr+1AQJ5II3
f753sKmDp8cW/I1gHYS48Ouj17yaac0zcJpQVzToMRmvY35yqHBDKQtRfEdaDhCy
94VmRvW2r3T/Nz7+t+YlAfxC919p6VbiRG5ffB/DCYhgbZXWkUwl2XFRcp+BwdQ4
hM0h5/sKe7gwdpi7uY66bPmQYNFqGG8h5gegciPyxHYIf/TkkqG67/hhdFFxHhib
Kp7gb6G6MaFGXTxHmO3L4elHSGX/2VlMgEozDvKOVfs72FGJSyc7lKGLWtNwlMdE
gs5Gbp+B1Z17l7HpIJF/QXHgAgQvoWNkgF605yOgIDeXHtEm7IJEkffj30ytARzX
hpYfmPNdpBP/59Hw4daQ2g==
`pragma protect end_protected
