`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zt6cIiEauBrNaIVE7s4JoVy+Ewb0hoeuDPq7nZCwJUKcni+3W3tTRNfxTT4OknIe
Q1rnDfRBSjI8MB3ERVxowEM4XbUL5HgRXrHVjNEN6dJJNupYDngcr/rdDKDb4as7
YpS4W0TZTaGaVZBG7CXurY7AEUdVfNir7NwgW4IpUMs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
ZZHLZbRHj3VVJdg45ez5SVRb3ZB7q6R8IqgkY/rPRgaKbPrbd9jYqxZQDgLSU9m3
dyd4XotQ0fsXc6AOp9aMeo6tSdgyZU2Zr+8XhEGWW6EzkofuV7FKBRjKT/pKXrmo
XuidHcifeT67Wm2j2hyQBUj59fk2cGaI91yu74nY17NrH2A2FpLvuSnmNBQW0Lmr
dRK+F5+jNd0ED6sNIbab5INXDauLG/7AZ0HnokhotdiWYsr2N0K/dgAc5MTxu/WH
FWIDa/duV11L95dQj21R4aLVoSWsWh+0yjky7kUFi65yd1Rj+SuAESwWVvNdAx4O
k9UDwpUPNL1936vnRHH7R1bSRIBLcRFORexhJpxdF6I8/XjJTMunQbg8s+CKETY3
BTfX5e4wySvax5D7VRVZ464MuiTEWv7hF5lghrKoi5xCF2wjYKWXS8pD/JAZkzNt
B+ixlAso5eleP9iUyHd/q13T79JwZAejrk7FdMMBNQpYxL04QkVGb0RD2856+KFm
5Gja7B83rk6N12hGNG/c985yUJgi1rVBrsrU85j/cWv/dyH4OOHBB4LaEYioK1BW
AvTydW+/ch8pDup4yxVuppfkBYkUG391mtOmOcnM6qioyMt+19q1umGk8fdyezUl
pPEFRdxj0qnDGjCsGw/5Z8MnJvbORxp7+AMJvzotL9yZBAdWYYgNocANx21T/gn9
OwunPxQXXDSsBgWctR4IqZn69AFF6Oxvn6Re18Ql+pUf7D2Te6F91Ml9ZsqU9DM0
fTwSfe2hpAZc+7mKB5TGODVFgVP2O/tl9m5bVI1hecMbiE87TSyTPOvUCIzUoSfL
JK9KRW4K1p7m22d++/AZa2eJlfdPhKZC+NxVnB6oz+CaC4I/wGfDeH8AtASYaUHA
oAxHg0er0AEzlGghZp8CuNSnAyR3iJdadN3w/yL1V4gtDMh/XVaCxMWI6uPvEC9Q
IO+B6JDCcIENjSr9N5d+Xtplus7r/AjkHcNdFxQj5GjBourfo3R3+YbGPIbuyhDt
XdTGqXYd/YOD0lari437SFjcgLJspqYijAv6Pn6Xx95oXxfNSE/7imoKe0KIphiL
DC4NxDOybGi0engr57fEGmaTRoqsI5XU99suXwa5lFpRRaBBk9UJ9ljfaej9Eig+
8lofmBEVSZOm1sbFYaUU7VwR0Bn2DAdXznwStv9T+AvAzuo7NS4uGhfzoGVRERxv
NJf6K1pqGc6DBmM76JtIOW8GBujCwYGEvU0w+Ifz0FmZXTIrNcTUySnzQTqPxqHp
rxThR9grMOfjn+RWqreHryq4fX0ur2L+4UaP0X+2x58cUEK/lwHT/BqhkS/kPYt/
Hs4IUHtVmUGAFJo/s2qjyZCP9jQQfpP3Dp7l3qnVL1Ai0f0PxNThbMZVYlsRg+qf
PZJqAnDqJhxHJvRyuM42LKF1FC6y9zfklXl73msJG3nO7weHeRN/LjpZoc37YJA0
xsla58RtUsyRtALp0vQxNE/Q3KyqNHOIQh0niuMuiXAMgwNRmHBlTCIQqs5xJclN
YtHfdnyhYOWd+m1nYrHf1wKX8R9Uqp4QiBOWKaTF2bOwmimYFRZynE/Y5QooMdHd
qT3Ty9IM9AoK8Kw8uMKDkzI4kHVIOG1QK92IdP5/j2SVwmB53CbNAfekrQXSPsHt
nLAX9UOGY3Xoox7cq/0Iy0yUJeliLkX3+dIx1nBaDyDCKqBPaUP3XySeqrFHqgjY
M+EuL6twAzbJc19EftjcWxmSTb2MCHIirmYfr0e9wYvuoEuIt5VTlBrd4WU2jgdy
f2oFbkSDrBOBOMIiCAr27rGg7ljmFoUB7X6vYkH61ce7fcjWCZTkPeTSE2P4m4AY
xE8PYHcpzh56J/ajeDyf/+84OZzANZLJJNuYElERISsllKJn5O9owTVaaA0jsRM6
4h0ERRaMMf+oCStJBLDd3OO5cWfmrbz570SCKU/b9T5yHk9JXOnbrJZjzPfjRVqe
GUrZHxtFrV0axb+rwDdJim0CID2nTat3xxEUtZfSV5VBfZxPCCBAekWY/VPlDnu9
PCNnz460QtUZ8utueRNinVgjOYMSlgZl/1qO7D3mSuLlCb0sOBf0T374DIan/g4A
yPEBp3TE1wpTkx7BCR5slVD9Ep/w1OnrqCYpObrzSwQ0Dd8Lwk1Vbtp5kV41Zw26
eq1awJRwfBT+VDDPvkOd8UD1LO/OPpXLgF7ZKpHfrJbceJGw/BWm+7a5CHdm4O7/
llGtUL4khZj6PewqecPwtUVYsESVpNMcv65a56YGLOSSQHzG7OFGjbOQnwF3Hg/0
OeAt+HVH9fQQ1Ulitbz4iooSgNi8+rbJCA8MhIWSl5ugvjbpWPZznto6fKw82hnY
W51hdjWup4ZeoZvTEQZqdABuEKJJ4PBJCcFy/7wpuqDLwC75n26kavuxABcyHx0Y
IiZNmfGH/KletxRLW9P03Xh4kN9VLFHTxWAo/x64eIKeu3spuL4MkNv561aFUHQC
0Tf8cSn6UAZpWw0FCNdVOjJRAsnTYjV2ThZ3YbcydlMWgl7nRYXdOzS/TgO4z6Ue
vjdSijC1dbTCGvdQ8WyPwbBZYO3dbmAEh+77buEWABZXhc/atX/z9VzSjzoDGd/s
9MFpdWQtd/QzrJSLZS6J4HEovc8iuhZYpj5qFYsHoo2kv1bgswoTku22X2NpjTAX
iR1j7V7MAhxg5mK/dPoniEZyIKhjqZFvzSBAzsjiDjnT9FFi29/09lTNKMu6Ud50
e3/msvQag9n8MtJJYoJXyHM3bTScX5vi+lurZQgxPt08kG3tPsWk8IorEvQEFdn3
dde9zgjJBlU5POUGhDjP5x2ZHOaYZs4DGNrwmBV6zktYXczjymUEmkjha2Y65LP2
+cQYIeu83M8xM4WVTyTmfJkEgeKR07ZdM9vS0AuYB95EYObSo+m3Ok1psmm/5SyX
Ekwwhmwl0LdQBj1DSbpJn338Lr4xcs+x+8G8LWPTtUAeTfMPNsMFZV9GGu9SyZ2A
o6piJj1Z8mbvLRB+L7RmeuVxoZWI31NYRe93tVmkXY1QNyMGEg753y/jmve9D7US
rHz2su4ZOm2VQdtlz1rNf+/DqHLwDz/eVsE+TR/RSE7yIp6gIdEs2Y05tZ78WL2Q
NUTf2fpIrMwP+TmyJcqSOUnYWYvKGnnAfksWukN/K3HlSUoEL2HWRVkS/sqPNvk2
QLv+1wGkW8YbLBEfICFLKIpqZb6bDfe+QQ3QeUZL6pSE96ScWdjL8azHyMlQxMLM
SRNh+tyYeywNSkJHORVmkkZ5aCZWGPiWSVho9osiHlUHkE5EeQDCIcFQku8omYqJ
84efhrWDpUO12ACFbYBG88Yd49iREgjATUxTu8jOrZq7NUrjPziZxvuewRZh1vbp
bpbuTuEp6LM49NWYfoq1jqgXcBxNRRukB/xim+wB/FGgdZ+rKILW+nIeZTZ/c4t5
BdgH+HUhdN5VWSV+5WgRm7UNbvpB4lAuY8FTEHlHbR1dss34f2Z0BIdT8zymPpEf
+2FhLRM48wL3miQ92DuXhaBZ+baitGBfXDdCytDGojRs6j97tmkKBpiT6l/CZzNx
jq/kk9k6KciaL3xLp2dcvUrDiu3bXElopZbY8wnQt/zNIp7Unzb3F3On8lEbRqqk
OTthiGPjnK4OOb0bdmsyRx8VEp7v3WP68LIoksDGPipm7Ys/SIO57e4eGyeO6rmD
ltLaPrA9MpnJNzt7sCt0WbREDXsCwfdkUKegHKYXUoYM5ebIXj0kYaw6r8dzdt+9
K3vm7MtGEp74LtyUxcqFyafWuWnftdse4+incXBURjz7RPZTmpki04ztZFRz9v4A
g+V8katiE5eUWV1ruhzndgfbYS55u5fSPfegbnqlj3ByC6MsEPYVlQWQWa5V598U
VwG5gurgDJpTRmkgcIcVIbpItdy3XP0x/olxBYpCXbx3vLs10PhXP8q0CYSYf2dU
xeLeJbGjJ/nzuwD494ztLA==
`pragma protect end_protected
