// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// 4:1 MUX of 129 bit words.  Latency 0.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_mux4w129t0s0 #(
    parameter SIM_EMULATE = 1'b0
) (
    input [515:0] din,
    input [1:0] sel,
    output [128:0] dout
);

genvar i,k;
generate
    for (i=0; i<129; i=i+1) begin : g0
        wire [3:0] local_din;
        for (k=0; k<4; k=k+1) begin : g1
            assign local_din[k] = din[k*129+i];
        end

        alt_e100s10_mux4w1t0s0 mx0 (
            .din(local_din),
            .sel(sel),
            .dout(dout[i])
        );
        defparam mx0 .SIM_EMULATE = SIM_EMULATE;

    end
endgenerate

endmodule

