// req_C1TxRAM2PORT.v

// Generated using ACDS version 17.0 290

`timescale 1 ps / 1 ps
module req_C1TxRAM2PORT (
		input  wire [555:0] data,      //  ram_input.datain
		input  wire [8:0]   wraddress, //           .wraddress
		input  wire [8:0]   rdaddress, //           .rdaddress
		input  wire         wren,      //           .wren
		input  wire         clock,     //           .clock
		output wire [555:0] q          // ram_output.dataout
	);

	req_C1TxRAM2PORT_ram_2port_170_hecum7i ram_2port_0 (
		.data      (data),      //  ram_input.datain
		.wraddress (wraddress), //           .wraddress
		.rdaddress (rdaddress), //           .rdaddress
		.wren      (wren),      //           .wren
		.clock     (clock),     //           .clock
		.q         (q)          // ram_output.dataout
	);

endmodule
