// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// 2:1 MUX of 1 bit words.  Latency 0.  Select latency 1.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_mux2w1t0s1 #(
    parameter SIM_EMULATE = 1'b0
) (
    input clk,
    input [1:0] din,
    input sel,
    output dout
);

reg [0:0] sel_r = 1'b0 /* synthesis preserve_syn_only */;
always @(posedge clk) sel_r <= sel;

alt_e100s10_mux2w1t0s0 mx0 (
    .din(din),
    .sel(sel_r),
    .dout(dout)
);
defparam mx0 .SIM_EMULATE = SIM_EMULATE;

endmodule

