// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// Pulse stretch to 64 cycles.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_pulse64 #(
    parameter SIM_EMULATE = 1'b0
) (
    input clk,
    input din,
    output dout
);

wire [5:0] cntr;
alt_e100s10_cnt6c ct0 (
    .clk(clk),
    .sclr(din),
    .dout(cntr)
);
defparam ct0 .SIM_EMULATE = SIM_EMULATE;

reg expire_helper = 1'b0;
always @(posedge clk) begin
     expire_helper <= cntr[1] & cntr[2] & cntr[3] & cntr[4] & cntr[5];
end

wire cntr_expire = cntr[0] & expire_helper;

reg dout_r = 1'b0;
always @(posedge clk) begin
    if (din) dout_r <= 1'b1;
    else if (cntr_expire) dout_r <= 1'b0;
end

assign dout = dout_r;
endmodule

