// pll.v

// Generated using ACDS version 18.1 222

`timescale 1 ps / 1 ps
module pll (
		input  wire  pll_refclk0,  //  pll_refclk0.clk
		output wire  outclk_div1,  //  outclk_div1.clk
		output wire  outclk_div2,  //  outclk_div2.clk
		output wire  pll_locked,   //   pll_locked.pll_locked
		output wire  pll_cal_busy  // pll_cal_busy.pll_cal_busy
	);

	pll_altera_xcvr_fpll_s10_htile_181_3xznj3i #(
		.rcfg_enable                                                             (0),
		.rcfg_jtag_enable                                                        (0),
		.rcfg_separate_avmm_busy                                                 (0),
		.dbg_embedded_debug_enable                                               (0),
		.dbg_capability_reg_enable                                               (0),
		.dbg_user_identifier                                                     (0),
		.dbg_stat_soft_logic_enable                                              (0),
		.dbg_ctrl_soft_logic_enable                                              (0),
		.rcfg_emb_strm_enable                                                    (0),
		.rcfg_profile_cnt                                                        (2),
		.cmu_fpll_refclk_select_mux_clk_sel_override                             ("normal"),
		.cmu_fpll_refclk_select_mux_clk_sel_override_value                       ("select_clk0"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq0_scratch0_src       ("iq0_scratch0_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq0_scratch1_src       ("iq0_scratch1_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq0_scratch2_src       ("iq0_scratch2_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq0_scratch3_src       ("iq0_scratch3_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq0_scratch4_src       ("iq0_scratch4_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq1_scratch0_src       ("iq1_scratch0_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq1_scratch1_src       ("iq1_scratch1_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq1_scratch2_src       ("iq1_scratch2_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq1_scratch3_src       ("iq1_scratch3_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_fpll_iq1_scratch4_src       ("iq1_scratch4_power_down"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_0_scratch0_src    ("pll_clkin_0_scratch0_src_vss"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_0_scratch1_src    ("pll_clkin_0_scratch1_src_vss"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_0_scratch2_src    ("pll_clkin_0_scratch2_src_vss"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_0_scratch3_src    ("pll_clkin_0_scratch3_src_vss"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_0_scratch4_src    ("pll_clkin_0_scratch4_src_vss"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_1_scratch0_src    ("pll_clkin_1_scratch0_src_vss"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_1_scratch1_src    ("pll_clkin_1_scratch1_src_vss"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_1_scratch2_src    ("pll_clkin_1_scratch2_src_vss"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_1_scratch3_src    ("pll_clkin_1_scratch3_src_vss"),
		.cmu_fpll_refclk_select_mux_pm_cmu_fpll_atom_pll_clkin_1_scratch4_src    ("pll_clkin_1_scratch4_src_vss"),
		.cmu_fpll_refclk_select_mux_powerdown_mode                               ("powerup"),
		.cmu_fpll_refclk_select_mux_sup_mode                                     ("user_mode"),
		.cmu_fpll_refclk_select_mux_xpm_clkin_fpll_pll_clkin_0_src               ("pll_clkin_0_src_ref_clk"),
		.cmu_fpll_refclk_select_mux_xpm_clkin_fpll_pll_clkin_1_src               ("pll_clkin_1_src_ref_clk"),
		.cmu_fpll_refclk_select_mux_xpm_clkin_fpll_xpm_pll_so_pll_auto_clk_sw_en ("pll_auto_clk_sw_disabled"),
		.cmu_fpll_refclk_select_mux_xpm_clkin_fpll_xpm_pll_so_pll_clk_loss_edge  ("pll_clk_loss_rising_edge"),
		.cmu_fpll_refclk_select_mux_xpm_clkin_fpll_xpm_pll_so_pll_clk_loss_sw_en ("pll_clk_loss_sw_byps"),
		.cmu_fpll_refclk_select_mux_xpm_clkin_fpll_xpm_pll_so_pll_clk_sw_dly     (0),
		.cmu_fpll_refclk_select_mux_xpm_clkin_fpll_xpm_pll_so_pll_manu_clk_sw_en ("pll_manu_clk_sw_disabled"),
		.cmu_fpll_refclk_select_mux_xpm_clkin_fpll_xpm_pll_so_pll_sw_refclk_src  ("pll_sw_refclk_src_clk_0"),
		.cmu_fpll_refclk_select_mux_silicon_rev                                  ("14nm5bcr2eb"),
		.cmu_fpll_refclk_select_mux_refclk_select0                               ("ref_iqclk0"),
		.cmu_fpll_refclk_select_mux_refclk_select1                               ("ref_iqclk0"),
		.cmu_fpll_refclk_select_mux_mux0_inclk0_logical_to_physical_mapping      ("ref_iqclk0"),
		.cmu_fpll_refclk_select_mux_mux0_inclk1_logical_to_physical_mapping      ("power_down"),
		.cmu_fpll_refclk_select_mux_mux0_inclk2_logical_to_physical_mapping      ("power_down"),
		.cmu_fpll_refclk_select_mux_mux0_inclk3_logical_to_physical_mapping      ("power_down"),
		.cmu_fpll_refclk_select_mux_mux0_inclk4_logical_to_physical_mapping      ("power_down"),
		.cmu_fpll_refclk_select_mux_mux1_inclk0_logical_to_physical_mapping      ("ref_iqclk0"),
		.cmu_fpll_refclk_select_mux_mux1_inclk1_logical_to_physical_mapping      ("power_down"),
		.cmu_fpll_refclk_select_mux_mux1_inclk2_logical_to_physical_mapping      ("power_down"),
		.cmu_fpll_refclk_select_mux_mux1_inclk3_logical_to_physical_mapping      ("power_down"),
		.cmu_fpll_refclk_select_mux_mux1_inclk4_logical_to_physical_mapping      ("power_down"),
		.hssi_avmm2_if_pcs_arbiter_ctrl                                          ("avmm2_arbiter_uc_sel"),
		.hssi_avmm2_if_pcs_cal_done                                              ("avmm2_cal_done_deassert"),
		.hssi_avmm2_if_pcs_cal_reserved                                          (0),
		.hssi_avmm2_if_pcs_calibration_feature_en                                ("avmm2_pcs_calibration_en"),
		.hssi_avmm2_if_pldadapt_gate_dis                                         ("disable"),
		.hssi_avmm2_if_pcs_hip_cal_en                                            ("disable"),
		.hssi_avmm2_if_hssiadapt_avmm_osc_clock_setting                          ("osc_clk_div_by1"),
		.hssi_avmm2_if_pldadapt_avmm_osc_clock_setting                           ("osc_clk_div_by1"),
		.hssi_avmm2_if_hssiadapt_avmm_testbus_sel                                ("avmm1_transfer_testbus"),
		.hssi_avmm2_if_pldadapt_avmm_testbus_sel                                 ("avmm1_transfer_testbus"),
		.hssi_avmm2_if_hssiadapt_hip_mode                                        ("disable_hip"),
		.hssi_avmm2_if_pldadapt_hip_mode                                         ("disable_hip"),
		.hssi_avmm2_if_silicon_rev                                               ("14nm5bcr2eb"),
		.hssi_avmm2_if_calibration_type                                          ("one_time"),
		.cmu_fpll_analog_mode                                                    ("analog_off"),
		.cmu_fpll_bonding                                                        ("bond_off"),
		.cmu_fpll_bw_mode                                                        ("mid_bw"),
		.cmu_fpll_cali_ref_off                                                   ("ref_on"),
		.cmu_fpll_cali_vco_off                                                   ("vco_on"),
		.cmu_fpll_cgb_div                                                        (1),
		.cmu_fpll_chgpmp_testmode                                                ("cp_normal"),
		.cmu_fpll_datarate_bps                                                   ("0"),
		.cmu_fpll_device_variant                                                 ("device_off"),
		.cmu_fpll_enable_hclk                                                    ("false"),
		.cmu_fpll_f_max_band_0                                                   ("3861860000"),
		.cmu_fpll_f_max_band_1                                                   ("4287223000"),
		.cmu_fpll_f_max_band_2                                                   ("4688476000"),
		.cmu_fpll_f_max_band_3                                                   ("5072700000"),
		.cmu_fpll_f_max_band_4                                                   ("5423191000"),
		.cmu_fpll_f_max_band_5                                                   ("5762211000"),
		.cmu_fpll_f_max_band_6                                                   ("6075045000"),
		.cmu_fpll_f_max_band_7                                                   ("6374148000"),
		.cmu_fpll_f_max_band_8                                                   ("14025000000"),
		.cmu_fpll_f_max_band_9                                                   ("1"),
		.cmu_fpll_f_max_div_two_bypass                                           ("1"),
		.cmu_fpll_f_max_pfd                                                      ("350000000"),
		.cmu_fpll_f_max_pfd_bonded                                               ("600000000"),
		.cmu_fpll_f_max_pfd_fractional                                           ("800000000"),
		.cmu_fpll_f_max_pfd_integer                                              ("800000000"),
		.cmu_fpll_f_max_vco                                                      ("14150000000"),
		.cmu_fpll_f_max_vco_fractional                                           ("14025000000"),
		.cmu_fpll_f_min_band_0                                                   ("7000000000"),
		.cmu_fpll_f_min_band_1                                                   ("3861860000"),
		.cmu_fpll_f_min_band_2                                                   ("4287223000"),
		.cmu_fpll_f_min_band_3                                                   ("4688476000"),
		.cmu_fpll_f_min_band_4                                                   ("5072700000"),
		.cmu_fpll_f_min_band_5                                                   ("5423191000"),
		.cmu_fpll_f_min_band_6                                                   ("5762211000"),
		.cmu_fpll_f_min_band_7                                                   ("6075045000"),
		.cmu_fpll_f_min_band_8                                                   ("6374148000"),
		.cmu_fpll_f_min_band_9                                                   ("1"),
		.cmu_fpll_f_min_pfd                                                      ("29000000"),
		.cmu_fpll_f_min_vco                                                      ("6000000000"),
		.cmu_fpll_f_out_c0                                                       ("312500000"),
		.cmu_fpll_f_out_c0_hz                                                    ("312500000"),
		.cmu_fpll_f_out_c1                                                       ("0"),
		.cmu_fpll_f_out_c1_hz                                                    ("0"),
		.cmu_fpll_f_out_c2                                                       ("0"),
		.cmu_fpll_f_out_c2_hz                                                    ("0"),
		.cmu_fpll_f_out_c3                                                       ("1"),
		.cmu_fpll_f_out_c3_hz                                                    ("1"),
		.cmu_fpll_feedback                                                       ("normal"),
		.cmu_fpll_cal_reserved                                                   ("fpll_cal_reserved_off"),
		.cmu_fpll_cal_test_sel                                                   ("sel_cal_out_7_to_0"),
		.cmu_fpll_calibration                                                    ("fpll_cal_enable"),
		.cmu_fpll_cas_out_enable                                                 ("fpll_cas_out_disable"),
		.cmu_fpll_cmu_rstn_value                                                 ("cmu_normal"),
		.cmu_fpll_dyn_reconfig                                                   ("fpll_dyn_reconfig_off"),
		.cmu_fpll_hclk_out_enable                                                ("fpll_hclk_out_disable"),
		.cmu_fpll_iqtxrxclk_out_enable                                           ("fpll_iqtxrxclk_out_disable"),
		.cmu_fpll_lpf_rstn_value                                                 ("lpf_normal"),
		.cmu_fpll_ppm_clk0_src                                                   ("ppm_clk0_vss"),
		.cmu_fpll_ppm_clk1_src                                                   ("ppm_clk1_vss"),
		.cmu_fpll_rstn_override                                                  ("user_reset_normal"),
		.cmu_fpll_initial_settings                                               ("true"),
		.cmu_fpll_is_otn                                                         ("false"),
		.cmu_fpll_is_pa_core                                                     ("false"),
		.cmu_fpll_is_sdi                                                         ("false"),
		.cmu_fpll_l_counter                                                      (1),
		.cmu_fpll_m_counter                                                      (64),
		.cmu_fpll_m_counter_c0                                                   (0),
		.cmu_fpll_m_counter_c1                                                   (0),
		.cmu_fpll_m_counter_c2                                                   (0),
		.cmu_fpll_m_counter_c3                                                   (0),
		.cmu_fpll_max_fractional_percentage                                      (99),
		.cmu_fpll_min_fractional_percentage                                      (1),
		.cmu_fpll_n_counter                                                      (3),
		.cmu_fpll_optimal                                                        ("false"),
		.cmu_fpll_out_freq                                                       ("312500000"),
		.cmu_fpll_out_freq_hz                                                    ("312500000"),
		.cmu_fpll_pfd_freq                                                       ("107421875"),
		.cmu_fpll_phase_shift_c0                                                 ("0.0"),
		.cmu_fpll_phase_shift_c1                                                 ("0.0"),
		.cmu_fpll_phase_shift_c2                                                 ("0.0"),
		.cmu_fpll_phase_shift_c3                                                 ("0.0"),
		.cmu_fpll_pll_vco_freq_band_0_dyn_high_bits                              (2),
		.cmu_fpll_pll_vco_freq_band_0_dyn_low_bits                               (0),
		.cmu_fpll_pll_vco_freq_band_0_fix                                        (2),
		.cmu_fpll_pll_vco_freq_band_0_fix_high                                   ("pll_vco_freq_band_0_fix_high_0"),
		.cmu_fpll_pll_vco_freq_band_1_dyn_high_bits                              (2),
		.cmu_fpll_pll_vco_freq_band_1_dyn_low_bits                               (0),
		.cmu_fpll_pll_vco_freq_band_1_fix                                        (2),
		.cmu_fpll_pll_vco_freq_band_1_fix_high                                   ("pll_vco_freq_band_1_fix_high_0"),
		.cmu_fpll_pma_width                                                      (64),
		.cmu_fpll_power_mode                                                     ("mid_power"),
		.cmu_fpll_power_rail_et                                                  (0),
		.cmu_fpll_powerdown_mode                                                 ("powerup"),
		.cmu_fpll_powermode_ac_ccnt1                                             ("fpll_ccnt1_ac_off"),
		.cmu_fpll_powermode_ac_ccnt2                                             ("fpll_ccnt2_ac_off"),
		.cmu_fpll_powermode_ac_ccnt3                                             ("fpll_ccnt3_ac_off"),
		.cmu_fpll_powermode_dc_ccnt0                                             ("fpll_ccnt0_dc"),
		.cmu_fpll_powermode_dc_ccnt1                                             ("powerdown_fpll_ccnt1"),
		.cmu_fpll_powermode_dc_ccnt2                                             ("powerdown_fpll_ccnt2"),
		.cmu_fpll_powermode_dc_ccnt3                                             ("powerdown_fpll_ccnt3"),
		.cmu_fpll_primary_use                                                    ("core"),
		.cmu_fpll_prot_mode                                                      ("basic_tx"),
		.cmu_fpll_refclk                                                         ("322265625"),
		.cmu_fpll_set_input_freq_range                                           (0),
		.cmu_fpll_side                                                           ("side_unknown"),
		.cmu_fpll_bcm_silicon_rev                                                ("rev_off"),
		.cmu_fpll_speed_grade                                                    ("speed_off"),
		.cmu_fpll_sup_mode                                                       ("user_mode"),
		.cmu_fpll_top_or_bottom                                                  ("top_or_bot_off"),
		.cmu_fpll_vco_freq                                                       ("13750000000"),
		.cmu_fpll_vco_freq_hz                                                    ("13750000000"),
		.cmu_fpll_c0_pllcout_enable                                              ("pllcout_enable"),
		.cmu_fpll_c0_cnt_div                                                     (11),
		.cmu_fpll_c0_cnt_min_tco                                                 ("cnt_enable_dly"),
		.cmu_fpll_c0_m_cnt_in_src                                                ("m_cnt_in_src_ph_mux_clk"),
		.cmu_fpll_c0_m_cnt_ph_mux_prst                                           (0),
		.cmu_fpll_c0_m_cnt_prst                                                  (1),
		.cmu_fpll_c1_pllcout_enable                                              ("pllcout_disable"),
		.cmu_fpll_c1_cnt_div                                                     (1),
		.cmu_fpll_c1_cnt_min_tco                                                 ("cnt_enable_dly"),
		.cmu_fpll_c1_m_cnt_in_src                                                ("m_cnt_in_src_ph_mux_clk"),
		.cmu_fpll_c1_m_cnt_ph_mux_prst                                           (0),
		.cmu_fpll_c1_m_cnt_prst                                                  (1),
		.cmu_fpll_c2_pllcout_enable                                              ("pllcout_disable"),
		.cmu_fpll_c2_cnt_div                                                     (1),
		.cmu_fpll_c2_cnt_min_tco                                                 ("cnt_enable_dly"),
		.cmu_fpll_c2_m_cnt_in_src                                                ("m_cnt_in_src_ph_mux_clk"),
		.cmu_fpll_c2_m_cnt_ph_mux_prst                                           (0),
		.cmu_fpll_c2_m_cnt_prst                                                  (1),
		.cmu_fpll_c3_pllcout_enable                                              ("pllcout_disable"),
		.cmu_fpll_c3_cnt_div                                                     (1),
		.cmu_fpll_c3_cnt_min_tco                                                 ("cnt_enable_dly"),
		.cmu_fpll_c3_m_cnt_in_src                                                ("m_cnt_in_src_ph_mux_clk"),
		.cmu_fpll_c3_m_cnt_ph_mux_prst                                           (0),
		.cmu_fpll_c3_m_cnt_prst                                                  (1),
		.cmu_fpll_cal_vco_count_length                                           ("sel_8b_count"),
		.cmu_fpll_lckdet_sel                                                     ("lckdet_sel_analog"),
		.cmu_fpll_refclk_source                                                  ("normal_refclk"),
		.cmu_fpll_pfd_delay_compensation                                         ("normal_delay"),
		.cmu_fpll_pfd_pulse_width                                                ("pulse_width_setting0"),
		.cmu_fpll_ppmdtct_lock_thresld                                           ("ppmdtct_lock_0"),
		.cmu_fpll_ppmdtct_noclk_thresld                                          ("ppmdtct_noclk_0"),
		.cmu_fpll_ppmdtct_pll_sel                                                ("ppmdtct_sel_fpll"),
		.cmu_fpll_vccdreg_fb                                                     ("vreg_fb0"),
		.cmu_fpll_vccdreg_fw                                                     ("vreg_fw0"),
		.cmu_fpll_vreg0_atbsel                                                   ("atb_disabled"),
		.cmu_fpll_vreg1_atbsel                                                   ("atb_disabled1"),
		.cmu_fpll_atb_atb                                                        ("atb_selectdisable"),
		.cmu_fpll_fb_fbclk_mux_1                                                 ("pll_fbclk_mux_1_glb"),
		.cmu_fpll_fb_fbclk_mux_2                                                 ("pll_fbclk_mux_2_m_cnt"),
		.cmu_fpll_iqfb_mux_iqclk_sel                                             ("iqtxrxclk0"),
		.cmu_fpll_chgpmp_compensation                                            ("cp_mode_enable"),
		.cmu_fpll_chgpmp_current_setting                                         ("cp_current_setting25"),
		.cmu_fpll_cp_current_boost                                               ("normal_setting"),
		.cmu_fpll_lf_3rd_pole_freq                                               ("lf_3rd_pole_setting0"),
		.cmu_fpll_lf_cbig                                                        ("lf_cbig_setting4"),
		.cmu_fpll_lf_order                                                       ("lf_2nd_order"),
		.cmu_fpll_lf_resistance                                                  ("lf_res_setting1"),
		.cmu_fpll_lf_ripplecap                                                   ("lf_no_ripple"),
		.cmu_fpll_vco_ph0_en                                                     ("pll_vco_ph0_en"),
		.cmu_fpll_vco_ph0_value                                                  ("pll_vco_ph0_vss"),
		.cmu_fpll_vco_ph1_en                                                     ("pll_vco_ph1_en"),
		.cmu_fpll_vco_ph1_value                                                  ("pll_vco_ph1_vss"),
		.cmu_fpll_vco_ph2_en                                                     ("pll_vco_ph2_en"),
		.cmu_fpll_vco_ph2_value                                                  ("pll_vco_ph2_vss"),
		.cmu_fpll_vco_ph3_en                                                     ("pll_vco_ph3_en"),
		.cmu_fpll_vco_ph3_value                                                  ("pll_vco_ph3_vss"),
		.cmu_fpll_dsm_mode                                                       ("dsm_mode_integer"),
		.cmu_fpll_pll_dsm_out_sel                                                ("pll_dsm_disable"),
		.cmu_fpll_pll_ecn_bypass                                                 ("pll_ecn_bypass_disable"),
		.cmu_fpll_pll_ecn_test_en                                                ("pll_ecn_test_disable"),
		.cmu_fpll_pll_fractional_division                                        ("0"),
		.cmu_fpll_pll_fractional_value_ready                                     ("pll_k_ready"),
		.cmu_fpll_lcnt_l_cnt_bypass                                              ("lcnt_normal"),
		.cmu_fpll_pll_l_counter                                                  (1),
		.cmu_fpll_lcnt_l_cnt_enable                                              ("lcnt_dis"),
		.cmu_fpll_lockf_lock_fltr_cfg                                            (25),
		.cmu_fpll_lockf_lock_fltr_test                                           ("pll_lock_fltr_nrm"),
		.cmu_fpll_lockf_unlock_fltr_cfg                                          (2),
		.cmu_fpll_mcnt_cnt_div                                                   (64),
		.cmu_fpll_mcnt_cnt_min_tco                                               ("cnt_bypass_dly"),
		.cmu_fpll_mcnt_m_cnt_in_src                                              ("m_cnt_in_src_ph_mux_clk"),
		.cmu_fpll_mcnt_m_cnt_ph_mux_prst                                         (0),
		.cmu_fpll_mcnt_m_cnt_prst                                                (1),
		.cmu_fpll_mcnt_coarse_dly                                                ("pll_coarse_dly_setting0"),
		.cmu_fpll_mcnt_fine_dly                                                  ("pll_fine_dly_setting0"),
		.cmu_fpll_ncnt_ncnt_divide                                               (3),
		.cmu_fpll_ncnt_coarse_dly                                                ("pll_coarse_dly_setting0"),
		.cmu_fpll_ncnt_fine_dly                                                  ("pll_fine_dly_setting0"),
		.cmu_fpll_ref_ref_buf_dly                                                ("pll_ref_buf_dly_setting0"),
		.cmu_fpll_testmux_tclk_mux_en                                            ("pll_tclk_mux_disabled"),
		.cmu_fpll_testmux_tclk_sel                                               ("pll_tclk_m_src"),
		.cmu_fpll_dprio_base_addr                                                (256),
		.cmu_fpll_dprio_broadcast_en                                             ("dprio_dprio_broadcast_en_csr_ctrl_disable"),
		.cmu_fpll_dprio_cvp_inter_sel                                            ("dprio_cvp_inter_sel_csr_ctrl_disable"),
		.cmu_fpll_dprio_force_inter_sel                                          ("dprio_force_inter_sel_csr_ctrl_disable"),
		.cmu_fpll_dprio_power_iso_en                                             ("dprio_power_iso_en_csr_ctrl_disable"),
		.cmu_fpll_dprio_status_select                                            ("dprio_normal_status"),
		.cmu_fpll_extra_csr                                                      (0),
		.cmu_fpll_ctrl_nreset_prgmnvrt                                           ("nreset_noninv"),
		.cmu_fpll_ctrl_ctrl_override_setting                                     ("pll_ctrl_enable"),
		.cmu_fpll_ctrl_enable                                                    ("pll_enabled"),
		.cmu_fpll_ctrl_slf_rst                                                   ("pll_slf_rst_off"),
		.cmu_fpll_ctrl_test_enable                                               ("pll_testen_off"),
		.cmu_fpll_ctrl_plniotri_override                                         ("plniotri_ctrl_disable"),
		.cmu_fpll_ctrl_vccr_pd                                                   ("vccd_powerup"),
		.cmu_fpll_silicon_rev                                                    ("14nm5bcr2eb"),
		.cmu_fpll_pll_op_mode                                                    ("false"),
		.cmu_fpll_bw_sel                                                         ("auto"),
		.cmu_fpll_compensation_mode                                              ("direct"),
		.cmu_fpll_duty_cycle_0                                                   (50),
		.cmu_fpll_duty_cycle_1                                                   (50),
		.cmu_fpll_duty_cycle_2                                                   (50),
		.cmu_fpll_duty_cycle_3                                                   (50),
		.cmu_fpll_hssi_output_clock_frequency                                    ("312500000"),
		.cmu_fpll_is_cascaded_pll                                                ("false"),
		.cmu_fpll_output_clock_frequency_0                                       ("312500000"),
		.cmu_fpll_output_clock_frequency_1                                       ("312500000"),
		.cmu_fpll_output_clock_frequency_2                                       ("312500000"),
		.cmu_fpll_output_clock_frequency_3                                       ("312500000"),
		.cmu_fpll_reference_clock_frequency                                      ("322265625"),
		.cmu_fpll_vco_frequency                                                  ("13750000000"),
		.enable_clk_divider                                                      (1),
		.test_mode                                                               ("false"),
		.hip_cal_en                                                              ("disable"),
		.enable_dps                                                              (0),
		.direct_dps                                                              (1),
		.calibration_en                                                          ("enable"),
		.enable_pcie_hip_connectivity                                            (0),
		.enable_mcgb                                                             (0),
		.enable_mcgb_reset                                                       (0),
		.enable_mcgb_debug_ports_parameters                                      (0),
		.hssi_pma_cgb_master_prot_mode                                           ("basic_tx"),
		.hssi_pma_cgb_master_silicon_rev                                         ("14nm5bcr2eb"),
		.hssi_pma_cgb_master_x1_div_m_sel                                        ("divbypass"),
		.hssi_pma_cgb_master_cgb_enable_iqtxrxclk                                ("disable_iqtxrxclk"),
		.hssi_pma_cgb_master_ser_mode                                            ("sixty_four_bit"),
		.hssi_pma_cgb_master_datarate_bps                                        ("625000000"),
		.hssi_pma_cgb_master_cgb_power_down                                      ("normal_cgb"),
		.hssi_pma_cgb_master_observe_cgb_clocks                                  ("observe_nothing"),
		.hssi_pma_cgb_master_tx_ucontrol_reset_pcie                              ("pcscorehip_controls_mcgb"),
		.hssi_pma_cgb_master_vccdreg_output                                      ("vccdreg_nominal"),
		.hssi_pma_cgb_master_input_select                                        ("fpll_top"),
		.hssi_pma_cgb_master_input_select_gen3                                   ("not_used")
	) xcvr_fpll_s10_htile_0 (
		.pll_refclk0             (pll_refclk0),                          //   input,  width = 1,  pll_refclk0.clk
		.outclk_div1             (outclk_div1),                          //  output,  width = 1,  outclk_div1.clk
		.outclk_div2             (outclk_div2),                          //  output,  width = 1,  outclk_div2.clk
		.pll_locked              (pll_locked),                           //  output,  width = 1,   pll_locked.pll_locked
		.pll_cal_busy            (pll_cal_busy),                         //  output,  width = 1, pll_cal_busy.pll_cal_busy
		.pll_powerdown           (1'b0),                                 // (terminated),                          
		.pll_refclk1             (1'b0),                                 // (terminated),                          
		.pll_refclk2             (1'b0),                                 // (terminated),                          
		.pll_refclk3             (1'b0),                                 // (terminated),                          
		.pll_refclk4             (1'b0),                                 // (terminated),                          
		.tx_serial_clk           (),                                     // (terminated),                          
		.outclk                  (),                                     // (terminated),                          
		.unused_pllcout          (),                                     // (terminated),                          
		.outclk_div4             (),                                     // (terminated),                          
		.pll_locked_hip          (),                                     // (terminated),                          
		.pll_pcie_clk            (),                                     // (terminated),                          
		.pll_cascade_clk         (),                                     // (terminated),                          
		.atx_to_fpll_cascade_clk (1'b0),                                 // (terminated),                          
		.reconfig_clk0           (1'b0),                                 // (terminated),                          
		.reconfig_reset0         (1'b0),                                 // (terminated),                          
		.reconfig_write0         (1'b0),                                 // (terminated),                          
		.reconfig_read0          (1'b0),                                 // (terminated),                          
		.reconfig_address0       (11'b00000000000),                      // (terminated),                          
		.reconfig_writedata0     (32'b00000000000000000000000000000000), // (terminated),                          
		.reconfig_readdata0      (),                                     // (terminated),                          
		.reconfig_waitrequest0   (),                                     // (terminated),                          
		.avmm_busy0              (),                                     // (terminated),                          
		.phase_reset             (1'b0),                                 // (terminated),                          
		.phase_enable            (1'b0),                                 // (terminated),                          
		.updn                    (1'b0),                                 // (terminated),                          
		.cntsel                  (4'b0000),                              // (terminated),                          
		.num_phase_shifts        (3'b001),                               // (terminated),                          
		.phase_done              (),                                     // (terminated),                          
		.hip_cal_done            (),                                     // (terminated),                          
		.mcgb_hip_cal_done       (),                                     // (terminated),                          
		.clklow                  (),                                     // (terminated),                          
		.fref                    (),                                     // (terminated),                          
		.mcgb_rst                (1'b0),                                 // (terminated),                          
		.mcgb_rst_stat           (),                                     // (terminated),                          
		.mcgb_aux_clk0           (1'b0),                                 // (terminated),                          
		.mcgb_aux_clk1           (1'b0),                                 // (terminated),                          
		.mcgb_aux_clk2           (1'b0),                                 // (terminated),                          
		.tx_bonding_clocks       (),                                     // (terminated),                          
		.mcgb_serial_clk         (),                                     // (terminated),                          
		.pcie_sw                 (2'b00),                                // (terminated),                          
		.pcie_sw_done            (),                                     // (terminated),                          
		.reconfig_clk1           (1'b0),                                 // (terminated),                          
		.reconfig_reset1         (1'b0),                                 // (terminated),                          
		.reconfig_write1         (1'b0),                                 // (terminated),                          
		.reconfig_read1          (1'b0),                                 // (terminated),                          
		.reconfig_address1       (11'b00000000000),                      // (terminated),                          
		.reconfig_writedata1     (32'b00000000000000000000000000000000), // (terminated),                          
		.reconfig_readdata1      (),                                     // (terminated),                          
		.reconfig_waitrequest1   (),                                     // (terminated),                          
		.mcgb_cal_busy           ()                                      // (terminated),                          
	);

endmodule
